module algo(

);




endmodule