
`define W_size 16 // word size (PARAMETER)
`define K_size 128 // Key size (PARAMETER)
`define U 2 // W_size/2
`define T 26 // 2*(number of rounds + 1)
`define B 16 // key size in bytes
`define C 8 // c=b/u=16/2=8
`define P 16'hb7e1
`define Q 16'h9e37

// UNCOMMENT THIS DEFINE FOR ALL 10,000 TEST CASES!!!!
`define FULL

`timescale 1ns / 1ps
module key_tb;

logic start;
logic clk;
logic rst;
logic [128:0] key;
logic [`W_size-1:0] sub [0:`T-1];
logic [4:0] num_rounds;
logic ready;

assign num_rounds = 12;

keygen Keygen(.*);

default clocking ckb @(posedge clk);
    input sub, ready;
    output rst, key, start;
endclocking

always begin
    clk = 1'b0;
    #1;
    clk = 1'b1;
    #1;
end

task reset();
    rst <= 1;
    ##1;
    rst <= 0;
    ##1;
endtask

task test_expansion(logic[`K_size-1:0] test_key, logic [`W_size-1:0] test_subkey [0:`T-1]);
    key <= test_key;

    reset();

    start <= 1;
    ##1;

    start <= 0;

    while(~ready) begin
        ##1;
    end

    for(int i = 0; i < `T; i++) begin
        assert(test_subkey[i] == sub[i])
            else begin
                $error("Bad Subkey Value: 0x%x at position %0d, should be 0x%x", sub[i], i, test_subkey[i]);
                $finish;
            end
    end
endtask

initial begin
    $fsdbDumpfile("dump.fsdb");
	$fsdbDumpvars(0, "+all");
    key <= 0;
    rst <= 0;
    start <= 0;

    #2;

    reset();

    // Known Test Case
	test_expansion(128'hdeadbeefdeadbeefdeadbeefdeadbeef, {16'd55048, 16'd43744, 16'd48559, 16'd27403, 16'd20374, 16'd33387, 16'd2062, 16'd61013, 16'd49237, 16'd33709, 16'd16278, 16'd65452, 16'd9968, 16'd4572, 16'd34933, 16'd35205, 16'd37470, 16'd42119, 16'd21025, 16'd13567, 16'd19718, 16'd1446, 16'd11664, 16'd40137, 16'd19576, 16'd15720});

    // AUTO GENERATED TEST CASES
	`ifdef FULL

	test_expansion(128'h07014645bf03130bf49f4b5e604a73c9, {16'd17554, 16'd18837, 16'd48166, 16'd39244, 16'd54638, 16'd34209, 16'd51923, 16'd44059, 16'd46276, 16'd29300, 16'd33630, 16'd55271, 16'd50802, 16'd44101, 16'd47462, 16'd50269, 16'd58548, 16'd1688, 16'd5774, 16'd52070, 16'd35646, 16'd50687, 16'd59665, 16'd24324, 16'd63665, 16'd63953});
	test_expansion(128'h4bf54a829b0f8c9d5776d1542e40b63f, {16'd10499, 16'd992, 16'd54846, 16'd13080, 16'd16030, 16'd33955, 16'd9833, 16'd63388, 16'd12245, 16'd25517, 16'd35995, 16'd18812, 16'd61023, 16'd40232, 16'd59115, 16'd4579, 16'd3303, 16'd33517, 16'd35340, 16'd30172, 16'd35992, 16'd46490, 16'd27589, 16'd19366, 16'd5016, 16'd60400});
	test_expansion(128'hf8a8ab15710c92eae46887db83c43ed1, {16'd51937, 16'd14621, 16'd10176, 16'd52191, 16'd28655, 16'd48775, 16'd5426, 16'd24239, 16'd62420, 16'd29366, 16'd62586, 16'd5652, 16'd11744, 16'd16758, 16'd995, 16'd20527, 16'd21164, 16'd48981, 16'd43904, 16'd19991, 16'd17554, 16'd51465, 16'd49709, 16'd21765, 16'd16908, 16'd41788});
	test_expansion(128'h46a58d4280665b103d74cccb97c102ee, {16'd59435, 16'd63166, 16'd51349, 16'd55409, 16'd21708, 16'd10557, 16'd8332, 16'd59678, 16'd59757, 16'd44379, 16'd58341, 16'd45948, 16'd60307, 16'd42467, 16'd9115, 16'd22890, 16'd61130, 16'd22829, 16'd19230, 16'd11444, 16'd59924, 16'd58625, 16'd4175, 16'd55500, 16'd36912, 16'd11420});
	test_expansion(128'h75a416d4824ee271f4d9055901c6c5c8, {16'd20701, 16'd10951, 16'd50754, 16'd14471, 16'd36125, 16'd62293, 16'd4263, 16'd21982, 16'd41198, 16'd10148, 16'd33341, 16'd55347, 16'd60176, 16'd48728, 16'd12430, 16'd9325, 16'd38051, 16'd49235, 16'd51837, 16'd32418, 16'd20178, 16'd59547, 16'd18505, 16'd22240, 16'd22851, 16'd59852});
	test_expansion(128'h3405ba0f5aef5388bda3cf3187a81ede, {16'd52054, 16'd9302, 16'd18213, 16'd55570, 16'd13059, 16'd4908, 16'd8089, 16'd55102, 16'd23644, 16'd48406, 16'd15061, 16'd22543, 16'd2542, 16'd21807, 16'd59229, 16'd17995, 16'd55416, 16'd54443, 16'd56678, 16'd64945, 16'd62110, 16'd58381, 16'd23878, 16'd1759, 16'd16459, 16'd8031});
	test_expansion(128'h89e60bf9760e5317c174be0cd61eb9bb, {16'd53964, 16'd37499, 16'd32723, 16'd46928, 16'd26016, 16'd10082, 16'd60939, 16'd34996, 16'd16145, 16'd33568, 16'd8383, 16'd54242, 16'd38016, 16'd40827, 16'd16747, 16'd54333, 16'd57293, 16'd3195, 16'd41061, 16'd55702, 16'd51115, 16'd5767, 16'd35546, 16'd24723, 16'd26255, 16'd40177});
	test_expansion(128'h118b74e2f32119246c168c1612c6a290, {16'd58199, 16'd40670, 16'd58310, 16'd43984, 16'd14874, 16'd36011, 16'd25042, 16'd51808, 16'd33631, 16'd58042, 16'd63684, 16'd17559, 16'd43429, 16'd27631, 16'd49660, 16'd17409, 16'd64571, 16'd59743, 16'd23735, 16'd22802, 16'd48466, 16'd37086, 16'd23863, 16'd59895, 16'd65433, 16'd38463});
	test_expansion(128'h0d32e97a486ed25e6ed3d24662f370ce, {16'd44900, 16'd23443, 16'd43923, 16'd63904, 16'd32372, 16'd54854, 16'd9136, 16'd40231, 16'd11316, 16'd44880, 16'd33358, 16'd623, 16'd35391, 16'd55296, 16'd60741, 16'd53194, 16'd30487, 16'd8449, 16'd42906, 16'd5400, 16'd39471, 16'd6094, 16'd62759, 16'd50202, 16'd8449, 16'd65009});
	test_expansion(128'h8cf0ff9257610e36a09b67400f951e90, {16'd32080, 16'd49869, 16'd44560, 16'd15544, 16'd34168, 16'd53105, 16'd22528, 16'd63448, 16'd5880, 16'd39591, 16'd51298, 16'd59510, 16'd44263, 16'd59370, 16'd22668, 16'd35769, 16'd11380, 16'd49224, 16'd58016, 16'd20412, 16'd65039, 16'd1166, 16'd25892, 16'd15131, 16'd28915, 16'd8480});
	test_expansion(128'h8a9156e27d97f801be296b2b7d0510f7, {16'd41715, 16'd5729, 16'd36340, 16'd48280, 16'd14724, 16'd55671, 16'd55829, 16'd24498, 16'd50637, 16'd31633, 16'd19217, 16'd64036, 16'd58036, 16'd22080, 16'd14979, 16'd40560, 16'd12503, 16'd49139, 16'd8113, 16'd47505, 16'd32183, 16'd46704, 16'd5031, 16'd40883, 16'd38830, 16'd24241});
	test_expansion(128'h1b1ef695f3244a9956b310584a22fc59, {16'd50493, 16'd38184, 16'd55153, 16'd62344, 16'd1571, 16'd64473, 16'd33637, 16'd10602, 16'd1852, 16'd21987, 16'd22913, 16'd26793, 16'd54327, 16'd12519, 16'd18136, 16'd59204, 16'd2473, 16'd53539, 16'd2144, 16'd46673, 16'd1626, 16'd16709, 16'd53150, 16'd57322, 16'd42428, 16'd50382});
	test_expansion(128'h916f9324e50198d0c45a3177e244ac08, {16'd63350, 16'd56955, 16'd59872, 16'd25814, 16'd36938, 16'd12967, 16'd14349, 16'd34773, 16'd19265, 16'd39854, 16'd43557, 16'd24619, 16'd45045, 16'd2463, 16'd27096, 16'd28078, 16'd16423, 16'd7066, 16'd30777, 16'd48429, 16'd18764, 16'd4256, 16'd1561, 16'd42527, 16'd15301, 16'd48409});
	test_expansion(128'ha46d8c895a484753091ccb6b813f623a, {16'd59939, 16'd26055, 16'd51979, 16'd38451, 16'd34103, 16'd51386, 16'd595, 16'd17581, 16'd27023, 16'd58522, 16'd24400, 16'd52776, 16'd61755, 16'd25746, 16'd42669, 16'd50178, 16'd28965, 16'd26512, 16'd9569, 16'd6157, 16'd39940, 16'd16971, 16'd57738, 16'd6578, 16'd17185, 16'd6995});
	test_expansion(128'h326706bbe8c775bd5005aa10c785d4f0, {16'd55167, 16'd33541, 16'd46937, 16'd5441, 16'd18547, 16'd50150, 16'd1133, 16'd62869, 16'd6126, 16'd48860, 16'd49463, 16'd10014, 16'd16305, 16'd23019, 16'd51112, 16'd20250, 16'd60993, 16'd43965, 16'd50787, 16'd27384, 16'd3659, 16'd60220, 16'd45438, 16'd33928, 16'd23331, 16'd29472});
	test_expansion(128'hc6275b6cf9e4caef7eef409d6a58eb14, {16'd13227, 16'd44112, 16'd52560, 16'd36430, 16'd9184, 16'd3589, 16'd64327, 16'd45906, 16'd24179, 16'd28105, 16'd46977, 16'd2791, 16'd40022, 16'd36772, 16'd45113, 16'd8683, 16'd42824, 16'd22219, 16'd5954, 16'd63899, 16'd56078, 16'd21245, 16'd24426, 16'd4043, 16'd62202, 16'd57009});
	test_expansion(128'h6dc171332b8919ceed572d3122e8a00f, {16'd64680, 16'd16856, 16'd18994, 16'd31850, 16'd17769, 16'd63187, 16'd34641, 16'd55327, 16'd52421, 16'd48851, 16'd23385, 16'd15525, 16'd61122, 16'd59090, 16'd46902, 16'd36660, 16'd51772, 16'd8760, 16'd32107, 16'd63921, 16'd18328, 16'd17558, 16'd30384, 16'd47896, 16'd30051, 16'd29536});
	test_expansion(128'hf5da45265633c8271a498b141443a402, {16'd57296, 16'd10978, 16'd51527, 16'd47131, 16'd61052, 16'd22272, 16'd34616, 16'd51241, 16'd37509, 16'd26876, 16'd47613, 16'd47519, 16'd11846, 16'd26033, 16'd12525, 16'd33648, 16'd30979, 16'd43290, 16'd19201, 16'd3745, 16'd260, 16'd20476, 16'd63746, 16'd35009, 16'd8590, 16'd64931});
	test_expansion(128'h912c2509e9f680b381f12c95a12e4469, {16'd13496, 16'd1076, 16'd34213, 16'd20894, 16'd16407, 16'd10741, 16'd63468, 16'd49867, 16'd64401, 16'd54826, 16'd28742, 16'd20787, 16'd13777, 16'd30668, 16'd42950, 16'd61516, 16'd34690, 16'd17373, 16'd62550, 16'd57660, 16'd46962, 16'd13420, 16'd29210, 16'd2947, 16'd40352, 16'd61822});
	test_expansion(128'hf3ee38cd186cb15c669789cfabddd51c, {16'd55882, 16'd41091, 16'd12123, 16'd48007, 16'd53113, 16'd2960, 16'd52541, 16'd15050, 16'd26605, 16'd243, 16'd45788, 16'd19230, 16'd6678, 16'd23978, 16'd60736, 16'd29222, 16'd36570, 16'd52498, 16'd13593, 16'd34586, 16'd53026, 16'd16746, 16'd47114, 16'd20750, 16'd50970, 16'd64522});
	test_expansion(128'h47adab81a93c19f911d0059c7d7df375, {16'd9618, 16'd12214, 16'd30052, 16'd65232, 16'd32602, 16'd9032, 16'd58601, 16'd19429, 16'd26312, 16'd5745, 16'd21031, 16'd42734, 16'd5633, 16'd6776, 16'd2111, 16'd36032, 16'd47583, 16'd50624, 16'd19949, 16'd34800, 16'd44019, 16'd32402, 16'd51072, 16'd42081, 16'd24526, 16'd16706});
	test_expansion(128'h69e3a77bb3ddb7da00eaaf81aa307ce9, {16'd30306, 16'd53977, 16'd6508, 16'd47662, 16'd65361, 16'd28202, 16'd22779, 16'd32523, 16'd18408, 16'd8256, 16'd16386, 16'd43061, 16'd55088, 16'd19251, 16'd34710, 16'd62289, 16'd23415, 16'd28573, 16'd7934, 16'd23690, 16'd62774, 16'd39699, 16'd1509, 16'd56181, 16'd33194, 16'd29460});
	test_expansion(128'h710972a8c8d2e369fb27d29a4ea6f3c4, {16'd39030, 16'd53337, 16'd41639, 16'd53979, 16'd10185, 16'd46648, 16'd46239, 16'd44590, 16'd39265, 16'd18891, 16'd41501, 16'd60432, 16'd23586, 16'd24354, 16'd30296, 16'd16610, 16'd49005, 16'd33611, 16'd40549, 16'd25332, 16'd56973, 16'd56462, 16'd12374, 16'd49148, 16'd7714, 16'd47544});
	test_expansion(128'hb8563e8b41719672ef2f494c7d2d11d4, {16'd21750, 16'd55455, 16'd15286, 16'd10971, 16'd34914, 16'd40656, 16'd30836, 16'd29074, 16'd14215, 16'd12397, 16'd30898, 16'd39501, 16'd58391, 16'd13633, 16'd36529, 16'd31251, 16'd44468, 16'd60609, 16'd126, 16'd33888, 16'd46206, 16'd55614, 16'd38111, 16'd294, 16'd2191, 16'd47189});
	test_expansion(128'h0c25cbfe2fa9d6e75378756a4181b961, {16'd49769, 16'd64158, 16'd10392, 16'd59975, 16'd60179, 16'd2046, 16'd19987, 16'd15826, 16'd62683, 16'd15174, 16'd20607, 16'd39843, 16'd2497, 16'd12792, 16'd13501, 16'd28694, 16'd52221, 16'd34835, 16'd14626, 16'd7728, 16'd31642, 16'd1348, 16'd62554, 16'd39131, 16'd32357, 16'd34930});
	test_expansion(128'h97d16d66b421cabe14638b1a5ad49078, {16'd34495, 16'd19392, 16'd121, 16'd43178, 16'd65372, 16'd38220, 16'd18440, 16'd49424, 16'd30135, 16'd57739, 16'd61613, 16'd21802, 16'd7026, 16'd49110, 16'd5377, 16'd28185, 16'd48089, 16'd40503, 16'd58276, 16'd7797, 16'd49599, 16'd41834, 16'd21605, 16'd34960, 16'd26549, 16'd38856});
	test_expansion(128'ha3b7699c7e965aaa3b6f87a3b289e513, {16'd11428, 16'd57451, 16'd12702, 16'd258, 16'd41020, 16'd7782, 16'd53829, 16'd61036, 16'd59717, 16'd33488, 16'd34981, 16'd35790, 16'd14799, 16'd51870, 16'd6384, 16'd40375, 16'd31250, 16'd37772, 16'd8163, 16'd24725, 16'd22815, 16'd17225, 16'd2463, 16'd22850, 16'd9035, 16'd25882});
	test_expansion(128'hd1c287f250090e17cbec72b53b221122, {16'd44526, 16'd64527, 16'd59470, 16'd1203, 16'd40820, 16'd38988, 16'd59949, 16'd27208, 16'd61672, 16'd58457, 16'd64605, 16'd43033, 16'd45447, 16'd24869, 16'd35670, 16'd52491, 16'd7999, 16'd27499, 16'd12288, 16'd27822, 16'd55086, 16'd62415, 16'd12172, 16'd39916, 16'd8462, 16'd15685});
	test_expansion(128'h6ff7c5302b56d6fbda86c82c741bc901, {16'd40730, 16'd6276, 16'd58631, 16'd41171, 16'd14029, 16'd30039, 16'd61332, 16'd14212, 16'd35442, 16'd12880, 16'd34084, 16'd63424, 16'd24172, 16'd29855, 16'd63678, 16'd10971, 16'd5145, 16'd24290, 16'd57789, 16'd2211, 16'd18649, 16'd1726, 16'd22922, 16'd23084, 16'd61379, 16'd1615});
	test_expansion(128'h4dc819d115c7d3cfc680b9269806fc71, {16'd24747, 16'd40735, 16'd13895, 16'd61946, 16'd38644, 16'd5352, 16'd43468, 16'd8650, 16'd41045, 16'd6035, 16'd32640, 16'd6267, 16'd57365, 16'd3722, 16'd18872, 16'd63366, 16'd1035, 16'd57202, 16'd7221, 16'd5933, 16'd5502, 16'd50875, 16'd611, 16'd34945, 16'd32284, 16'd5869});
	test_expansion(128'h49096fe3152294c58c8bdbfeb5466024, {16'd17174, 16'd43927, 16'd16860, 16'd27099, 16'd17373, 16'd34730, 16'd62294, 16'd42439, 16'd11132, 16'd54381, 16'd17706, 16'd59171, 16'd47181, 16'd54489, 16'd39529, 16'd17618, 16'd60690, 16'd2189, 16'd49793, 16'd662, 16'd50405, 16'd37262, 16'd32894, 16'd49039, 16'd58244, 16'd31998});
	test_expansion(128'hcf23f83b972f911287e03e8bd40c50ca, {16'd42313, 16'd32947, 16'd57768, 16'd10189, 16'd21965, 16'd47314, 16'd60426, 16'd14724, 16'd24108, 16'd34539, 16'd25665, 16'd2889, 16'd15476, 16'd40669, 16'd9432, 16'd63615, 16'd30301, 16'd37860, 16'd32376, 16'd8774, 16'd1727, 16'd60456, 16'd4038, 16'd24257, 16'd19502, 16'd40436});
	test_expansion(128'hf6a59288946134244f59ada75a979939, {16'd20981, 16'd35316, 16'd911, 16'd56026, 16'd30186, 16'd23350, 16'd37402, 16'd20596, 16'd9996, 16'd46002, 16'd27638, 16'd11377, 16'd9733, 16'd20707, 16'd20806, 16'd49088, 16'd37340, 16'd41402, 16'd5191, 16'd59112, 16'd57388, 16'd49712, 16'd48287, 16'd50854, 16'd38877, 16'd7379});
	test_expansion(128'h5889af8bb3204d353e78d6af71ab51cb, {16'd53288, 16'd21061, 16'd29591, 16'd11992, 16'd58791, 16'd8397, 16'd51763, 16'd64225, 16'd38230, 16'd19276, 16'd13099, 16'd27994, 16'd999, 16'd44343, 16'd25992, 16'd32672, 16'd35964, 16'd12400, 16'd15518, 16'd55106, 16'd16186, 16'd35781, 16'd32876, 16'd19245, 16'd43684, 16'd14088});
	test_expansion(128'haeda181aafbbdfaa941ed942150efe3a, {16'd14121, 16'd48175, 16'd8236, 16'd42150, 16'd28909, 16'd51992, 16'd38917, 16'd24283, 16'd21077, 16'd11000, 16'd25348, 16'd56450, 16'd26750, 16'd36498, 16'd64175, 16'd15431, 16'd17814, 16'd4797, 16'd19683, 16'd53783, 16'd11693, 16'd9266, 16'd26156, 16'd29390, 16'd32214, 16'd61396});
	test_expansion(128'h6808617c0ea3e19e9329014db5d6fb29, {16'd35800, 16'd41215, 16'd12037, 16'd59920, 16'd60976, 16'd59793, 16'd48195, 16'd53271, 16'd2953, 16'd15263, 16'd31578, 16'd34598, 16'd24245, 16'd55527, 16'd38214, 16'd19770, 16'd45233, 16'd61043, 16'd9750, 16'd6727, 16'd98, 16'd25865, 16'd2554, 16'd63305, 16'd10783, 16'd44418});
	test_expansion(128'h7d4b0e73e0f655940885c962a7ec706e, {16'd7508, 16'd27813, 16'd27183, 16'd52842, 16'd43443, 16'd39568, 16'd14233, 16'd41871, 16'd64248, 16'd51205, 16'd2483, 16'd62184, 16'd21070, 16'd22853, 16'd37741, 16'd54172, 16'd47910, 16'd24234, 16'd12853, 16'd65101, 16'd21312, 16'd53578, 16'd39406, 16'd17971, 16'd50921, 16'd43619});
	test_expansion(128'hdf6959c6cc07ec065aa7413482a6b066, {16'd13798, 16'd56968, 16'd48688, 16'd17081, 16'd42323, 16'd37886, 16'd29509, 16'd62129, 16'd46695, 16'd58497, 16'd57290, 16'd44398, 16'd26789, 16'd61741, 16'd35226, 16'd49671, 16'd58441, 16'd53407, 16'd10698, 16'd51546, 16'd25814, 16'd31947, 16'd44303, 16'd51002, 16'd29148, 16'd64711});
	test_expansion(128'h7f978d59dac3471c32773b187d78cf1e, {16'd55906, 16'd822, 16'd14734, 16'd19055, 16'd64963, 16'd36455, 16'd54625, 16'd10070, 16'd38309, 16'd60284, 16'd59689, 16'd23320, 16'd32441, 16'd10375, 16'd367, 16'd46683, 16'd37405, 16'd56066, 16'd17374, 16'd16180, 16'd11850, 16'd45451, 16'd17027, 16'd33307, 16'd10993, 16'd3426});
	test_expansion(128'hd2a78bbc1bb35f77873c189ef7049402, {16'd4676, 16'd44465, 16'd18823, 16'd52650, 16'd33441, 16'd63445, 16'd25925, 16'd15210, 16'd36968, 16'd16052, 16'd54069, 16'd34752, 16'd24623, 16'd43441, 16'd39963, 16'd27789, 16'd3433, 16'd65198, 16'd26439, 16'd5029, 16'd49106, 16'd52306, 16'd44443, 16'd42752, 16'd19737, 16'd21754});
	test_expansion(128'hbd83477d1f7e608017669aee21d61674, {16'd55349, 16'd5463, 16'd41683, 16'd7058, 16'd3043, 16'd13588, 16'd27282, 16'd18523, 16'd335, 16'd60942, 16'd7719, 16'd26417, 16'd63156, 16'd55023, 16'd141, 16'd6619, 16'd14364, 16'd30888, 16'd36892, 16'd45409, 16'd34570, 16'd3292, 16'd51525, 16'd47355, 16'd45101, 16'd46115});
	test_expansion(128'h5e5881d40cdbd6cc28bf99f2f4f8644e, {16'd42763, 16'd39303, 16'd54492, 16'd526, 16'd31912, 16'd15327, 16'd3239, 16'd60937, 16'd42970, 16'd33955, 16'd64176, 16'd4760, 16'd865, 16'd43306, 16'd65431, 16'd46998, 16'd2890, 16'd21858, 16'd31236, 16'd3542, 16'd32604, 16'd21998, 16'd28164, 16'd22956, 16'd53472, 16'd35738});
	test_expansion(128'h6a6fefd1514ea49c64cc58430ffbbeb1, {16'd58844, 16'd240, 16'd45131, 16'd10876, 16'd42654, 16'd59713, 16'd14409, 16'd32130, 16'd42730, 16'd25623, 16'd6297, 16'd46316, 16'd50686, 16'd16399, 16'd22177, 16'd22486, 16'd33155, 16'd1066, 16'd49906, 16'd32014, 16'd40374, 16'd36192, 16'd48051, 16'd13178, 16'd59598, 16'd5780});
	test_expansion(128'hbd168a3b9d2ebca78caedcfb7eaa3176, {16'd49844, 16'd65456, 16'd7219, 16'd43920, 16'd10608, 16'd57929, 16'd10921, 16'd37635, 16'd23144, 16'd25933, 16'd24968, 16'd34119, 16'd22298, 16'd17261, 16'd29253, 16'd31068, 16'd22028, 16'd65474, 16'd25984, 16'd60311, 16'd13341, 16'd21092, 16'd51013, 16'd48947, 16'd63991, 16'd43794});
	test_expansion(128'h4ab6ff29663e67e5a7638860eba6e020, {16'd64849, 16'd7518, 16'd22146, 16'd37026, 16'd16687, 16'd48073, 16'd25925, 16'd32050, 16'd30120, 16'd58077, 16'd39057, 16'd7757, 16'd5091, 16'd14681, 16'd20366, 16'd24158, 16'd35545, 16'd8613, 16'd4900, 16'd21005, 16'd44463, 16'd28644, 16'd11780, 16'd7079, 16'd47170, 16'd64219});
	test_expansion(128'hcbb8672236c7934e2fb3db47b266dc43, {16'd39149, 16'd16087, 16'd4145, 16'd52932, 16'd40802, 16'd38593, 16'd45787, 16'd22920, 16'd38813, 16'd25055, 16'd34000, 16'd57448, 16'd33511, 16'd43784, 16'd60748, 16'd45651, 16'd27184, 16'd42663, 16'd50422, 16'd24722, 16'd4071, 16'd32585, 16'd27392, 16'd3682, 16'd52741, 16'd27021});
	test_expansion(128'hfe918a79ab0ae06225321d4e34b2a3e4, {16'd62859, 16'd59733, 16'd23775, 16'd30900, 16'd17494, 16'd55999, 16'd7775, 16'd5890, 16'd7409, 16'd13876, 16'd46903, 16'd22568, 16'd64269, 16'd54154, 16'd7902, 16'd54859, 16'd48259, 16'd11406, 16'd36956, 16'd56758, 16'd22647, 16'd22001, 16'd36901, 16'd53852, 16'd55222, 16'd60634});
	test_expansion(128'hd555992bbe980eda7d2bd6c29c919659, {16'd52926, 16'd59077, 16'd34885, 16'd11099, 16'd29189, 16'd56495, 16'd15997, 16'd520, 16'd35524, 16'd32655, 16'd15332, 16'd46713, 16'd30222, 16'd7318, 16'd33298, 16'd45087, 16'd47436, 16'd15998, 16'd6745, 16'd20435, 16'd59392, 16'd9770, 16'd15003, 16'd29849, 16'd3411, 16'd65056});
	test_expansion(128'hc4292a78714d1216ffd7e2fa21c4d8e9, {16'd18667, 16'd41426, 16'd35062, 16'd33880, 16'd46395, 16'd58971, 16'd44832, 16'd33961, 16'd33788, 16'd31014, 16'd42734, 16'd18528, 16'd6532, 16'd65049, 16'd7890, 16'd9072, 16'd7785, 16'd8631, 16'd38636, 16'd37628, 16'd4178, 16'd1223, 16'd64688, 16'd42637, 16'd25641, 16'd6504});
	test_expansion(128'h42b85e35e5b81cd44b138ab2e367da39, {16'd24091, 16'd358, 16'd16839, 16'd27294, 16'd27315, 16'd14175, 16'd53664, 16'd8194, 16'd32802, 16'd34547, 16'd63438, 16'd48080, 16'd57311, 16'd43403, 16'd62167, 16'd20832, 16'd3415, 16'd59911, 16'd43812, 16'd18684, 16'd64835, 16'd38915, 16'd38328, 16'd16825, 16'd7120, 16'd3661});
	test_expansion(128'h2b1e8349fbfdc0308ccd2eaf48c5db29, {16'd46928, 16'd9632, 16'd8495, 16'd63048, 16'd42755, 16'd13892, 16'd64661, 16'd41550, 16'd51763, 16'd59156, 16'd3130, 16'd54331, 16'd11195, 16'd61217, 16'd16913, 16'd54069, 16'd10990, 16'd63105, 16'd41084, 16'd21510, 16'd10028, 16'd23724, 16'd34800, 16'd31146, 16'd33558, 16'd21923});
	test_expansion(128'h5c32a42e579797a44748bb58c34c2eeb, {16'd12861, 16'd35050, 16'd17150, 16'd12130, 16'd59899, 16'd45270, 16'd59651, 16'd59497, 16'd63372, 16'd54554, 16'd40412, 16'd7853, 16'd46342, 16'd50727, 16'd21434, 16'd59604, 16'd8863, 16'd23472, 16'd23259, 16'd31820, 16'd39725, 16'd29129, 16'd21812, 16'd54866, 16'd26437, 16'd30945});
	test_expansion(128'hb0b18b0f07921111ea730650ff4b95e9, {16'd10275, 16'd110, 16'd4232, 16'd36446, 16'd8796, 16'd2640, 16'd44838, 16'd4228, 16'd56559, 16'd11270, 16'd39637, 16'd41807, 16'd31110, 16'd17396, 16'd31431, 16'd31052, 16'd58489, 16'd61065, 16'd58128, 16'd23252, 16'd45344, 16'd63443, 16'd5141, 16'd46537, 16'd23586, 16'd2730});
	test_expansion(128'h71641b9c7a4751897c04e97c8bfb1e0b, {16'd61915, 16'd15039, 16'd12771, 16'd6852, 16'd60584, 16'd52072, 16'd32094, 16'd2914, 16'd12552, 16'd64410, 16'd36088, 16'd38233, 16'd50496, 16'd15506, 16'd10371, 16'd58671, 16'd65509, 16'd53022, 16'd62353, 16'd25811, 16'd6008, 16'd56355, 16'd35124, 16'd40102, 16'd17611, 16'd56516});
	test_expansion(128'hcbc25b0ac976a3a9cbff1435fe499be2, {16'd36464, 16'd43269, 16'd2244, 16'd35358, 16'd35910, 16'd22068, 16'd63220, 16'd22945, 16'd10324, 16'd62906, 16'd42250, 16'd64484, 16'd17521, 16'd18010, 16'd55431, 16'd20464, 16'd7283, 16'd3745, 16'd47183, 16'd2295, 16'd17239, 16'd1966, 16'd1583, 16'd43040, 16'd3025, 16'd50745});
	test_expansion(128'h8b12744775fa1509a2543757edae3c65, {16'd5246, 16'd15694, 16'd5353, 16'd12929, 16'd40407, 16'd220, 16'd41526, 16'd28382, 16'd51985, 16'd33041, 16'd3216, 16'd29841, 16'd6652, 16'd42711, 16'd41611, 16'd16864, 16'd43511, 16'd44769, 16'd30247, 16'd10167, 16'd47277, 16'd37609, 16'd39843, 16'd2118, 16'd24007, 16'd61319});
	test_expansion(128'h27908d5b1323f26082c521d5e4edf12c, {16'd18383, 16'd3237, 16'd3181, 16'd10042, 16'd12503, 16'd47959, 16'd6941, 16'd6232, 16'd3902, 16'd20103, 16'd4836, 16'd19540, 16'd16506, 16'd42315, 16'd48870, 16'd2600, 16'd54574, 16'd39932, 16'd58792, 16'd33067, 16'd60272, 16'd2550, 16'd58139, 16'd11688, 16'd15405, 16'd37122});
	test_expansion(128'hb9b484080bf1be6e079b29a98c981d2f, {16'd22368, 16'd7704, 16'd5197, 16'd38771, 16'd58081, 16'd50733, 16'd61524, 16'd19811, 16'd34382, 16'd13092, 16'd21490, 16'd41386, 16'd8353, 16'd15680, 16'd7226, 16'd45632, 16'd25047, 16'd14009, 16'd38550, 16'd49790, 16'd2088, 16'd51670, 16'd60292, 16'd43182, 16'd3200, 16'd32488});
	test_expansion(128'h5f43bf003504b3ae3fc004b42ed03448, {16'd7917, 16'd58085, 16'd29827, 16'd29002, 16'd47976, 16'd63506, 16'd28167, 16'd50737, 16'd13523, 16'd45615, 16'd22887, 16'd64010, 16'd3362, 16'd6742, 16'd25176, 16'd31886, 16'd41455, 16'd14262, 16'd45721, 16'd49214, 16'd64156, 16'd54963, 16'd44142, 16'd48822, 16'd31855, 16'd42550});
	test_expansion(128'h526f0195961cfd2f08b62476021f0d6e, {16'd4615, 16'd3034, 16'd26297, 16'd13128, 16'd1092, 16'd11580, 16'd14290, 16'd62188, 16'd63347, 16'd14248, 16'd14915, 16'd62289, 16'd35502, 16'd27911, 16'd15526, 16'd3489, 16'd4931, 16'd9305, 16'd19454, 16'd5676, 16'd46316, 16'd34433, 16'd4204, 16'd8578, 16'd57946, 16'd42421});
	test_expansion(128'h38e83658e2861665c0e32abb1d7aa421, {16'd36710, 16'd62803, 16'd63089, 16'd55365, 16'd1385, 16'd53523, 16'd51396, 16'd33101, 16'd24967, 16'd57376, 16'd40565, 16'd35348, 16'd52745, 16'd18649, 16'd39503, 16'd41038, 16'd53251, 16'd34466, 16'd12467, 16'd5346, 16'd35241, 16'd47415, 16'd6199, 16'd10846, 16'd35691, 16'd58939});
	test_expansion(128'hf33e5bcfc0d1e395f3d893b866eebe25, {16'd11112, 16'd46651, 16'd16538, 16'd5003, 16'd7660, 16'd45517, 16'd4811, 16'd62885, 16'd60942, 16'd43212, 16'd53800, 16'd26112, 16'd50242, 16'd47399, 16'd12436, 16'd25074, 16'd16409, 16'd16706, 16'd51570, 16'd45983, 16'd34398, 16'd2617, 16'd57136, 16'd30833, 16'd38690, 16'd52683});
	test_expansion(128'h62d50660fdd3bc9fa15b8a656896a23e, {16'd36781, 16'd25333, 16'd42562, 16'd60189, 16'd27616, 16'd30891, 16'd46501, 16'd23041, 16'd50528, 16'd31318, 16'd25674, 16'd22121, 16'd58540, 16'd17030, 16'd16063, 16'd24215, 16'd44990, 16'd50349, 16'd13915, 16'd19214, 16'd11574, 16'd27149, 16'd49596, 16'd50655, 16'd11452, 16'd28109});
	test_expansion(128'h41451325081115673ec25ef0c3087bda, {16'd2503, 16'd14251, 16'd64261, 16'd34015, 16'd62550, 16'd44616, 16'd25553, 16'd27077, 16'd38821, 16'd1259, 16'd12282, 16'd18090, 16'd27682, 16'd44771, 16'd37172, 16'd60603, 16'd16798, 16'd12879, 16'd46036, 16'd44499, 16'd64706, 16'd19535, 16'd42897, 16'd2239, 16'd63777, 16'd38060});
	test_expansion(128'h6f836df7d97950eb1a69ec200ecb49ab, {16'd64240, 16'd55583, 16'd60313, 16'd39355, 16'd26153, 16'd61300, 16'd19732, 16'd9923, 16'd27428, 16'd12021, 16'd58492, 16'd64509, 16'd40575, 16'd37983, 16'd919, 16'd39086, 16'd25417, 16'd8788, 16'd57138, 16'd52838, 16'd9310, 16'd23867, 16'd14443, 16'd36295, 16'd31293, 16'd19022});
	test_expansion(128'h24f22ad456ac1759577a3575317b86af, {16'd35169, 16'd15315, 16'd16360, 16'd51118, 16'd65, 16'd56583, 16'd37124, 16'd26336, 16'd3621, 16'd36745, 16'd22090, 16'd40055, 16'd63703, 16'd58375, 16'd13654, 16'd33344, 16'd46699, 16'd30340, 16'd29680, 16'd41059, 16'd57038, 16'd18540, 16'd3220, 16'd29401, 16'd39307, 16'd64686});
	test_expansion(128'hc2d17b8c53d3645d0b4c0551f320f091, {16'd55501, 16'd34067, 16'd38458, 16'd50674, 16'd45823, 16'd63673, 16'd58542, 16'd40706, 16'd23487, 16'd26241, 16'd4265, 16'd58345, 16'd1766, 16'd48138, 16'd15619, 16'd43713, 16'd26436, 16'd34489, 16'd44647, 16'd22732, 16'd51587, 16'd45076, 16'd8590, 16'd24457, 16'd44418, 16'd24606});
	test_expansion(128'h0a63aa3423f6d475093c8d231bc8b3b4, {16'd8817, 16'd36487, 16'd33640, 16'd51310, 16'd17730, 16'd41092, 16'd13444, 16'd54132, 16'd15542, 16'd32914, 16'd39722, 16'd54183, 16'd61918, 16'd1532, 16'd53350, 16'd11611, 16'd23679, 16'd53511, 16'd53153, 16'd48785, 16'd54794, 16'd36531, 16'd38955, 16'd10547, 16'd55266, 16'd32123});
	test_expansion(128'hcb3ef72033fad1d9141fbe67628484d1, {16'd51270, 16'd48588, 16'd11706, 16'd19286, 16'd13051, 16'd56602, 16'd25577, 16'd32935, 16'd58407, 16'd31942, 16'd61128, 16'd6972, 16'd38792, 16'd26077, 16'd30794, 16'd47344, 16'd5122, 16'd3522, 16'd3855, 16'd10563, 16'd61263, 16'd6884, 16'd56069, 16'd1613, 16'd2905, 16'd46552});
	test_expansion(128'hf3f7f271264e9e4e1541d34eee20fbbe, {16'd26444, 16'd40607, 16'd33923, 16'd24763, 16'd12112, 16'd20602, 16'd12211, 16'd63186, 16'd59474, 16'd52232, 16'd42121, 16'd61908, 16'd45807, 16'd50885, 16'd34876, 16'd15316, 16'd4583, 16'd49977, 16'd19678, 16'd45875, 16'd38628, 16'd45534, 16'd43660, 16'd47806, 16'd16430, 16'd32117});
	test_expansion(128'h76da3e9bfaf3885a9862e204dc3b0498, {16'd14064, 16'd45207, 16'd49811, 16'd3484, 16'd52317, 16'd18486, 16'd39191, 16'd58264, 16'd54934, 16'd27833, 16'd863, 16'd3344, 16'd15049, 16'd37488, 16'd2216, 16'd17721, 16'd37894, 16'd41291, 16'd40350, 16'd5075, 16'd6636, 16'd2935, 16'd15761, 16'd39793, 16'd30926, 16'd7532});
	test_expansion(128'h4bf754576496e14a50ae2ef2c1319205, {16'd43742, 16'd22835, 16'd44578, 16'd18289, 16'd52409, 16'd30924, 16'd12775, 16'd40082, 16'd41296, 16'd8159, 16'd24079, 16'd3001, 16'd38216, 16'd13730, 16'd42607, 16'd9059, 16'd47684, 16'd42798, 16'd38997, 16'd31669, 16'd62502, 16'd30908, 16'd28624, 16'd61571, 16'd11795, 16'd40983});
	test_expansion(128'h10035574e86e1f87fbf8c36df482f8a8, {16'd19924, 16'd28655, 16'd47824, 16'd57474, 16'd26226, 16'd10188, 16'd46863, 16'd30349, 16'd9363, 16'd2050, 16'd4994, 16'd36253, 16'd33937, 16'd2759, 16'd10971, 16'd30572, 16'd31250, 16'd22614, 16'd30117, 16'd64413, 16'd10840, 16'd4659, 16'd37416, 16'd59716, 16'd51443, 16'd16472});
	test_expansion(128'h358325f2bf538f5b6cfe6eccdd48ebd8, {16'd47060, 16'd53461, 16'd30625, 16'd53363, 16'd61628, 16'd11650, 16'd31587, 16'd56441, 16'd57834, 16'd64285, 16'd12096, 16'd14701, 16'd17216, 16'd60040, 16'd14274, 16'd41023, 16'd34488, 16'd64817, 16'd57774, 16'd7024, 16'd22524, 16'd8879, 16'd28701, 16'd7105, 16'd1945, 16'd11021});
	test_expansion(128'h91982e479aaef9bbe3c07b97170f4d75, {16'd17025, 16'd23999, 16'd3154, 16'd19054, 16'd36056, 16'd43869, 16'd59739, 16'd43040, 16'd64543, 16'd19201, 16'd9769, 16'd29923, 16'd57773, 16'd6199, 16'd15404, 16'd34783, 16'd53567, 16'd2415, 16'd31117, 16'd34006, 16'd438, 16'd34285, 16'd5373, 16'd39898, 16'd2552, 16'd64527});
	test_expansion(128'h915848ac1208589daf1b67180528b41e, {16'd21960, 16'd20571, 16'd44539, 16'd37158, 16'd23477, 16'd63077, 16'd265, 16'd57581, 16'd10412, 16'd64672, 16'd1893, 16'd50009, 16'd10092, 16'd30085, 16'd4319, 16'd6063, 16'd18789, 16'd58384, 16'd60838, 16'd45566, 16'd50301, 16'd36334, 16'd16772, 16'd26104, 16'd6426, 16'd14305});
	test_expansion(128'hc3d8df17c5eb5948fa3cc728d614dc02, {16'd27281, 16'd28746, 16'd43754, 16'd21869, 16'd7600, 16'd41186, 16'd60140, 16'd43018, 16'd8500, 16'd12698, 16'd21247, 16'd54422, 16'd14064, 16'd35439, 16'd38811, 16'd43774, 16'd11676, 16'd7625, 16'd14053, 16'd27892, 16'd29578, 16'd1308, 16'd54693, 16'd60711, 16'd15945, 16'd64078});
	test_expansion(128'h254342ae46fe7815cbb7897865fbb28e, {16'd18398, 16'd27049, 16'd49720, 16'd28715, 16'd50504, 16'd37456, 16'd56232, 16'd13385, 16'd41743, 16'd36809, 16'd51266, 16'd61590, 16'd39107, 16'd61553, 16'd17862, 16'd258, 16'd29986, 16'd14127, 16'd35217, 16'd8449, 16'd6877, 16'd29001, 16'd21846, 16'd61530, 16'd11763, 16'd61953});
	test_expansion(128'h9127904fece5a9e73486e69481fe95e2, {16'd7938, 16'd36132, 16'd19285, 16'd17653, 16'd62725, 16'd5351, 16'd54499, 16'd26733, 16'd43574, 16'd38700, 16'd65141, 16'd12622, 16'd35407, 16'd42564, 16'd43220, 16'd5751, 16'd28530, 16'd24732, 16'd65258, 16'd53288, 16'd51939, 16'd38675, 16'd23709, 16'd31878, 16'd2840, 16'd8825});
	test_expansion(128'h22113eb2686542ab61b58bdd1ec62350, {16'd58256, 16'd40735, 16'd6550, 16'd37751, 16'd5415, 16'd35315, 16'd59340, 16'd36259, 16'd9388, 16'd14286, 16'd43407, 16'd46663, 16'd54830, 16'd3322, 16'd37212, 16'd16892, 16'd11277, 16'd24519, 16'd29389, 16'd62056, 16'd32616, 16'd58103, 16'd61175, 16'd32867, 16'd1692, 16'd39970});
	test_expansion(128'h2fcdb04979ef1210a932dbd7ca6b391c, {16'd14600, 16'd15864, 16'd35963, 16'd14904, 16'd47306, 16'd44263, 16'd21409, 16'd32094, 16'd12406, 16'd24593, 16'd36304, 16'd57638, 16'd27945, 16'd5612, 16'd13495, 16'd39945, 16'd22343, 16'd58339, 16'd56887, 16'd39518, 16'd43288, 16'd40210, 16'd48280, 16'd23997, 16'd27641, 16'd13192});
	test_expansion(128'haa09d3fec7f2f74489219022dd8ba5c9, {16'd32186, 16'd8966, 16'd58607, 16'd6703, 16'd24354, 16'd39016, 16'd64184, 16'd58994, 16'd31777, 16'd29667, 16'd15770, 16'd20590, 16'd63489, 16'd41292, 16'd24012, 16'd22073, 16'd63274, 16'd59326, 16'd6722, 16'd30490, 16'd22380, 16'd6963, 16'd30323, 16'd39562, 16'd20798, 16'd14583});
	test_expansion(128'hdb6503b0cad37c08e733b5e260e255d5, {16'd58807, 16'd54841, 16'd37571, 16'd22939, 16'd52567, 16'd299, 16'd27423, 16'd18488, 16'd40645, 16'd49495, 16'd9822, 16'd32385, 16'd53064, 16'd55778, 16'd32141, 16'd64376, 16'd38546, 16'd12113, 16'd15509, 16'd58545, 16'd40737, 16'd24377, 16'd55095, 16'd28411, 16'd59492, 16'd2864});
	test_expansion(128'h1bb12b67163513bef8c9bed5de6ca31f, {16'd16170, 16'd44680, 16'd46939, 16'd6051, 16'd942, 16'd36752, 16'd12344, 16'd2433, 16'd39503, 16'd12170, 16'd59505, 16'd3599, 16'd10431, 16'd37659, 16'd22713, 16'd23769, 16'd18799, 16'd40378, 16'd18034, 16'd47582, 16'd34202, 16'd25779, 16'd47767, 16'd2301, 16'd32044, 16'd19614});
	test_expansion(128'h2f7a490034fc2bd3fa40c14f22804c20, {16'd43271, 16'd63525, 16'd35831, 16'd61887, 16'd57005, 16'd30893, 16'd48654, 16'd3951, 16'd51542, 16'd15697, 16'd47001, 16'd9686, 16'd147, 16'd56619, 16'd55728, 16'd27957, 16'd30548, 16'd38322, 16'd29257, 16'd13359, 16'd33490, 16'd25280, 16'd63036, 16'd39661, 16'd12810, 16'd4921});
	test_expansion(128'he9b22faf470b3318ef0490eaa8e7b7ad, {16'd39153, 16'd5191, 16'd3342, 16'd28396, 16'd30046, 16'd30303, 16'd8777, 16'd12380, 16'd65244, 16'd41454, 16'd34315, 16'd43585, 16'd55170, 16'd36243, 16'd4508, 16'd61258, 16'd3212, 16'd36723, 16'd48364, 16'd43938, 16'd19421, 16'd1339, 16'd11231, 16'd21522, 16'd8721, 16'd40417});
	test_expansion(128'hdeafeb0a8eef546cab65bbb5db1a0654, {16'd14464, 16'd63083, 16'd6857, 16'd16150, 16'd65190, 16'd50106, 16'd32744, 16'd24285, 16'd38432, 16'd48234, 16'd47449, 16'd51313, 16'd39856, 16'd18101, 16'd46928, 16'd61851, 16'd41458, 16'd20332, 16'd19186, 16'd62604, 16'd37999, 16'd27393, 16'd25442, 16'd16566, 16'd55095, 16'd32611});
	test_expansion(128'h2138b4b4b871ff94b39a93b0ea5fbab8, {16'd11397, 16'd26402, 16'd33915, 16'd43355, 16'd44075, 16'd48656, 16'd33170, 16'd34441, 16'd43525, 16'd17437, 16'd24945, 16'd55183, 16'd13642, 16'd38789, 16'd52846, 16'd18011, 16'd46651, 16'd38617, 16'd31620, 16'd45312, 16'd29565, 16'd43542, 16'd23228, 16'd32162, 16'd13872, 16'd4926});
	test_expansion(128'hba56df0450eed98129f3087d921c4a18, {16'd40038, 16'd22301, 16'd48083, 16'd4003, 16'd58107, 16'd40345, 16'd29566, 16'd15828, 16'd12499, 16'd47951, 16'd14020, 16'd33978, 16'd40080, 16'd34435, 16'd60730, 16'd61697, 16'd44990, 16'd39405, 16'd45315, 16'd25790, 16'd7131, 16'd39502, 16'd34838, 16'd23036, 16'd48291, 16'd35392});
	test_expansion(128'h3ac5048996a1f2d88343a2d16c935fa3, {16'd28435, 16'd29806, 16'd29860, 16'd39176, 16'd5995, 16'd29057, 16'd64915, 16'd20894, 16'd55946, 16'd15319, 16'd57730, 16'd42988, 16'd42339, 16'd54745, 16'd34266, 16'd28046, 16'd61788, 16'd2758, 16'd54697, 16'd64957, 16'd31477, 16'd33438, 16'd26734, 16'd24946, 16'd54057, 16'd52995});
	test_expansion(128'hedca0c70a593429ed898d4bda5356745, {16'd36590, 16'd23675, 16'd21089, 16'd13061, 16'd20713, 16'd47425, 16'd33001, 16'd7819, 16'd1098, 16'd28721, 16'd25414, 16'd14035, 16'd31103, 16'd60410, 16'd34362, 16'd61734, 16'd28597, 16'd29226, 16'd65129, 16'd917, 16'd21190, 16'd47044, 16'd14696, 16'd63274, 16'd27774, 16'd42448});
	test_expansion(128'ha4156fec75f12450b2a9080873e390b4, {16'd6131, 16'd44841, 16'd43066, 16'd43642, 16'd38590, 16'd47275, 16'd1847, 16'd29290, 16'd32443, 16'd11785, 16'd56066, 16'd34345, 16'd33398, 16'd7484, 16'd14718, 16'd16356, 16'd27544, 16'd50052, 16'd46300, 16'd43662, 16'd41210, 16'd24244, 16'd60081, 16'd33468, 16'd17062, 16'd38562});
	test_expansion(128'hcc24fa0a6ecc85e5158420092d68e2bd, {16'd8176, 16'd63556, 16'd56224, 16'd61575, 16'd36642, 16'd39984, 16'd18693, 16'd6906, 16'd87, 16'd57596, 16'd20558, 16'd20365, 16'd49731, 16'd49588, 16'd31447, 16'd5084, 16'd31229, 16'd63839, 16'd55225, 16'd9161, 16'd39623, 16'd37215, 16'd64526, 16'd61601, 16'd32899, 16'd19760});
	test_expansion(128'haa3f0b13e5a2dc9ba56b4948b245964e, {16'd60951, 16'd10864, 16'd36914, 16'd18043, 16'd50920, 16'd44379, 16'd45771, 16'd46884, 16'd49204, 16'd45319, 16'd10672, 16'd27791, 16'd13529, 16'd44742, 16'd51438, 16'd36695, 16'd10462, 16'd17385, 16'd13319, 16'd1202, 16'd14873, 16'd11608, 16'd998, 16'd64148, 16'd62229, 16'd25295});
	test_expansion(128'h4d1f641f79bcdad44d9305bb02c7edb3, {16'd16849, 16'd23138, 16'd27467, 16'd56197, 16'd55028, 16'd20999, 16'd33072, 16'd11184, 16'd12096, 16'd45405, 16'd41825, 16'd61345, 16'd12412, 16'd56752, 16'd58518, 16'd35946, 16'd14281, 16'd51221, 16'd61967, 16'd47642, 16'd59322, 16'd4915, 16'd16643, 16'd26831, 16'd39721, 16'd22652});
	test_expansion(128'h5b7a4afc7aeffc75ac245c3860e9c35e, {16'd7264, 16'd56381, 16'd15582, 16'd45978, 16'd35678, 16'd21378, 16'd28944, 16'd58922, 16'd29454, 16'd56889, 16'd6039, 16'd30459, 16'd41663, 16'd20202, 16'd16542, 16'd8183, 16'd63399, 16'd47597, 16'd32662, 16'd34956, 16'd5377, 16'd43145, 16'd57898, 16'd3687, 16'd9177, 16'd63948});
	test_expansion(128'h1ab40e755ca4ebb01180cb5a6efe5728, {16'd39732, 16'd48274, 16'd44572, 16'd36714, 16'd61431, 16'd53088, 16'd27142, 16'd7827, 16'd34721, 16'd51997, 16'd14843, 16'd16425, 16'd14798, 16'd13460, 16'd35236, 16'd47147, 16'd49059, 16'd37339, 16'd40464, 16'd27034, 16'd11718, 16'd45144, 16'd59966, 16'd11343, 16'd12451, 16'd57464});
	test_expansion(128'h3b1a5a6b5f9f873ca66fcb82cab919c0, {16'd57295, 16'd12569, 16'd43781, 16'd61743, 16'd9953, 16'd53458, 16'd33585, 16'd26666, 16'd55370, 16'd9081, 16'd42771, 16'd23582, 16'd2687, 16'd18099, 16'd21630, 16'd52208, 16'd24252, 16'd52083, 16'd18313, 16'd53863, 16'd49906, 16'd52312, 16'd45342, 16'd38196, 16'd65169, 16'd45421});
	test_expansion(128'habea005700df31c61b03019a71a30085, {16'd38252, 16'd7340, 16'd50224, 16'd23700, 16'd23568, 16'd59333, 16'd28904, 16'd62016, 16'd10172, 16'd24377, 16'd20868, 16'd30823, 16'd65142, 16'd57992, 16'd36019, 16'd42145, 16'd50683, 16'd40679, 16'd59185, 16'd28426, 16'd50905, 16'd8775, 16'd35691, 16'd36860, 16'd23306, 16'd21451});
	test_expansion(128'h165a413d57ed24236d7829d0e5347f0d, {16'd22204, 16'd5786, 16'd11103, 16'd36964, 16'd4072, 16'd17615, 16'd53359, 16'd7643, 16'd24627, 16'd21123, 16'd59005, 16'd13734, 16'd37475, 16'd52427, 16'd37933, 16'd52851, 16'd24176, 16'd7606, 16'd53284, 16'd26895, 16'd20550, 16'd62093, 16'd15524, 16'd19723, 16'd52669, 16'd47461});
	test_expansion(128'h37252a8401cc7e6135fb8b0d340f9a78, {16'd21406, 16'd14231, 16'd10300, 16'd31947, 16'd6281, 16'd6290, 16'd1635, 16'd7791, 16'd33576, 16'd27170, 16'd23423, 16'd15849, 16'd42466, 16'd57920, 16'd31484, 16'd895, 16'd38305, 16'd33637, 16'd27671, 16'd16877, 16'd61003, 16'd12227, 16'd42671, 16'd59937, 16'd11358, 16'd48625});
	test_expansion(128'hfbc20b9f8f60da8294e08ad21936b280, {16'd412, 16'd59628, 16'd36177, 16'd19652, 16'd27206, 16'd39557, 16'd13037, 16'd29740, 16'd37707, 16'd54819, 16'd19074, 16'd39523, 16'd28046, 16'd42069, 16'd59542, 16'd25777, 16'd53133, 16'd49893, 16'd47356, 16'd20897, 16'd9544, 16'd31145, 16'd53817, 16'd13912, 16'd20287, 16'd53686});
	test_expansion(128'h476c55f4c80d8b1807bd6d08ea0bd1bc, {16'd61158, 16'd52229, 16'd59437, 16'd37267, 16'd45808, 16'd36184, 16'd23814, 16'd28895, 16'd25913, 16'd31911, 16'd44367, 16'd10030, 16'd28998, 16'd26588, 16'd861, 16'd64853, 16'd5104, 16'd29938, 16'd37257, 16'd52990, 16'd50685, 16'd50416, 16'd35505, 16'd29016, 16'd25865, 16'd42561});
	test_expansion(128'h03821ed8b1d84724a3bcb6c08fbaa2d5, {16'd1536, 16'd31433, 16'd41045, 16'd9206, 16'd15762, 16'd15521, 16'd34421, 16'd57450, 16'd11454, 16'd40451, 16'd58478, 16'd26596, 16'd63895, 16'd34948, 16'd1925, 16'd14078, 16'd50512, 16'd25508, 16'd38575, 16'd569, 16'd38291, 16'd34250, 16'd3931, 16'd28177, 16'd37147, 16'd24947});
	test_expansion(128'h7849aa9cb7cf7778d8c74a3a5ab73eef, {16'd54808, 16'd17357, 16'd35927, 16'd58342, 16'd9129, 16'd16832, 16'd33801, 16'd16611, 16'd35429, 16'd6637, 16'd10917, 16'd54991, 16'd41077, 16'd3647, 16'd22845, 16'd13315, 16'd24888, 16'd61631, 16'd48341, 16'd64131, 16'd38210, 16'd64461, 16'd59283, 16'd21606, 16'd25759, 16'd6649});
	test_expansion(128'he0a3e3187b219680304e7954bcfcac20, {16'd6976, 16'd47196, 16'd13122, 16'd7978, 16'd20056, 16'd44759, 16'd60376, 16'd16140, 16'd35790, 16'd38395, 16'd57023, 16'd23039, 16'd59735, 16'd54813, 16'd29476, 16'd16910, 16'd1074, 16'd20479, 16'd31072, 16'd28368, 16'd1615, 16'd49218, 16'd27302, 16'd110, 16'd14322, 16'd60267});
	test_expansion(128'hb8df10ce191f0c1c6e02385ae66704fa, {16'd61384, 16'd36032, 16'd35421, 16'd36193, 16'd56867, 16'd46975, 16'd27870, 16'd41857, 16'd23760, 16'd64785, 16'd40172, 16'd59555, 16'd55093, 16'd57480, 16'd50520, 16'd37712, 16'd38639, 16'd37348, 16'd28703, 16'd24186, 16'd14641, 16'd226, 16'd60880, 16'd11884, 16'd21445, 16'd62422});
	test_expansion(128'hccac5e4ab68a72cf0e024c04571aa949, {16'd52632, 16'd18631, 16'd29398, 16'd20997, 16'd63546, 16'd20865, 16'd38945, 16'd52353, 16'd62, 16'd23423, 16'd34259, 16'd28831, 16'd31172, 16'd37635, 16'd51796, 16'd41858, 16'd14809, 16'd54764, 16'd1416, 16'd29381, 16'd7410, 16'd33795, 16'd39533, 16'd6644, 16'd11058, 16'd12517});
	test_expansion(128'hce83a54408e0d1edccfc6b4ed47074f0, {16'd31670, 16'd14405, 16'd29626, 16'd37588, 16'd61766, 16'd33962, 16'd16184, 16'd49708, 16'd18115, 16'd28438, 16'd27397, 16'd56102, 16'd39282, 16'd33855, 16'd18970, 16'd47993, 16'd33945, 16'd48394, 16'd63969, 16'd51975, 16'd14972, 16'd5297, 16'd56360, 16'd12704, 16'd59583, 16'd26823});
	test_expansion(128'h012c5c6c200c31631b898c5ed1d5636c, {16'd53628, 16'd15746, 16'd62670, 16'd56054, 16'd42389, 16'd50803, 16'd52505, 16'd38856, 16'd12278, 16'd41614, 16'd6144, 16'd29127, 16'd46371, 16'd38410, 16'd27326, 16'd36012, 16'd2427, 16'd63156, 16'd58853, 16'd50830, 16'd53869, 16'd8344, 16'd48038, 16'd65454, 16'd16632, 16'd20237});
	test_expansion(128'h1be2472d9f241de20abbcd2291ebbbca, {16'd12607, 16'd55789, 16'd39000, 16'd42208, 16'd65043, 16'd11824, 16'd62267, 16'd58453, 16'd57220, 16'd48178, 16'd18069, 16'd42907, 16'd50057, 16'd4630, 16'd21435, 16'd12822, 16'd29360, 16'd12966, 16'd33449, 16'd19545, 16'd1377, 16'd12889, 16'd60400, 16'd29833, 16'd29030, 16'd62956});
	test_expansion(128'h3da2a2809f1969e4978adf1c6e02ea60, {16'd54087, 16'd39615, 16'd3819, 16'd45290, 16'd31255, 16'd26201, 16'd28485, 16'd4402, 16'd30690, 16'd13765, 16'd17387, 16'd34649, 16'd28676, 16'd11781, 16'd29645, 16'd23415, 16'd15063, 16'd22974, 16'd8100, 16'd50149, 16'd35420, 16'd92, 16'd14100, 16'd62062, 16'd7755, 16'd64398});
	test_expansion(128'h6108365f4ebb03608d6c09ef774b84dc, {16'd49131, 16'd12238, 16'd445, 16'd45999, 16'd24845, 16'd4448, 16'd42092, 16'd34844, 16'd55156, 16'd27657, 16'd15817, 16'd21750, 16'd10850, 16'd47326, 16'd48990, 16'd200, 16'd11809, 16'd15690, 16'd63786, 16'd28806, 16'd3430, 16'd65030, 16'd44920, 16'd44090, 16'd46236, 16'd30100});
	test_expansion(128'h3a0fd58655654c8a00e06b926489c5f4, {16'd13338, 16'd25612, 16'd22946, 16'd1697, 16'd59895, 16'd49716, 16'd374, 16'd10443, 16'd52319, 16'd27302, 16'd31954, 16'd37342, 16'd3282, 16'd9723, 16'd60527, 16'd43836, 16'd23978, 16'd36706, 16'd8302, 16'd7324, 16'd44345, 16'd13060, 16'd26953, 16'd50665, 16'd34940, 16'd41146});
	test_expansion(128'hb30c4f03379d2131e92a3b5436e80bfa, {16'd63585, 16'd65172, 16'd50952, 16'd56263, 16'd50448, 16'd27602, 16'd23859, 16'd4997, 16'd23124, 16'd28168, 16'd35155, 16'd56077, 16'd53933, 16'd31972, 16'd55838, 16'd53625, 16'd58323, 16'd15815, 16'd60705, 16'd42973, 16'd29589, 16'd50900, 16'd23147, 16'd37486, 16'd17381, 16'd6859});
	test_expansion(128'h716ff6c4200b9c82baf67fd55a63a624, {16'd4755, 16'd47694, 16'd63932, 16'd12112, 16'd35908, 16'd61921, 16'd61981, 16'd29651, 16'd60896, 16'd21450, 16'd3927, 16'd53324, 16'd3277, 16'd32159, 16'd51302, 16'd30414, 16'd48196, 16'd182, 16'd30786, 16'd47635, 16'd48759, 16'd25533, 16'd1833, 16'd29951, 16'd48310, 16'd28308});
	test_expansion(128'h72eb76decfe568ea026a04e94c0d2a1f, {16'd48919, 16'd37556, 16'd50741, 16'd340, 16'd36718, 16'd10043, 16'd34176, 16'd19970, 16'd13183, 16'd37721, 16'd2442, 16'd15748, 16'd15864, 16'd31464, 16'd47649, 16'd46960, 16'd49585, 16'd25264, 16'd21715, 16'd54175, 16'd23700, 16'd36490, 16'd40682, 16'd45667, 16'd10531, 16'd24061});
	test_expansion(128'ha86f6f9563c586612e7c3aba4954ddb4, {16'd45781, 16'd46232, 16'd60610, 16'd55435, 16'd28908, 16'd8344, 16'd44807, 16'd29608, 16'd8309, 16'd21234, 16'd4303, 16'd43636, 16'd9560, 16'd9839, 16'd25622, 16'd40757, 16'd30274, 16'd35010, 16'd22389, 16'd12734, 16'd17760, 16'd18552, 16'd40339, 16'd31946, 16'd5712, 16'd5396});
	test_expansion(128'h47de237d393f3ed8194f3d0df7b98a40, {16'd3954, 16'd64881, 16'd47262, 16'd50310, 16'd14263, 16'd11501, 16'd1310, 16'd16791, 16'd1320, 16'd9871, 16'd12013, 16'd17110, 16'd3860, 16'd12019, 16'd17055, 16'd24171, 16'd53768, 16'd19845, 16'd13054, 16'd39694, 16'd35688, 16'd27378, 16'd27101, 16'd60015, 16'd7513, 16'd6861});
	test_expansion(128'hd8b29b847d18d108be70d870af361311, {16'd40342, 16'd10940, 16'd46708, 16'd48106, 16'd53154, 16'd46228, 16'd64412, 16'd57024, 16'd52768, 16'd65322, 16'd54861, 16'd59225, 16'd56433, 16'd40864, 16'd49018, 16'd63642, 16'd24909, 16'd23737, 16'd27854, 16'd56519, 16'd9487, 16'd58267, 16'd45503, 16'd8133, 16'd48683, 16'd56121});
	test_expansion(128'h966bb54eb56935367c9beba2ab7ee88e, {16'd16780, 16'd8195, 16'd24229, 16'd60572, 16'd41707, 16'd24393, 16'd57220, 16'd49532, 16'd62322, 16'd36865, 16'd15289, 16'd37045, 16'd44258, 16'd288, 16'd22140, 16'd39296, 16'd32400, 16'd13557, 16'd25088, 16'd63622, 16'd60331, 16'd65325, 16'd12676, 16'd29785, 16'd49604, 16'd51145});
	test_expansion(128'h201a91102ec5e794170842e5b7737b9c, {16'd62040, 16'd64625, 16'd23822, 16'd60478, 16'd51228, 16'd11186, 16'd8373, 16'd55192, 16'd5581, 16'd21627, 16'd5328, 16'd11814, 16'd11837, 16'd11651, 16'd59637, 16'd57518, 16'd33279, 16'd33638, 16'd39785, 16'd6327, 16'd47790, 16'd11538, 16'd26713, 16'd57916, 16'd411, 16'd42966});
	test_expansion(128'h0876fa9c431c121642ee2f6704750f0f, {16'd28443, 16'd34378, 16'd17057, 16'd21572, 16'd2076, 16'd33993, 16'd25931, 16'd36001, 16'd47840, 16'd29538, 16'd17969, 16'd47351, 16'd54437, 16'd22668, 16'd42146, 16'd26572, 16'd23460, 16'd9423, 16'd63251, 16'd59165, 16'd42071, 16'd53610, 16'd10872, 16'd28562, 16'd23781, 16'd8159});
	test_expansion(128'h9994e9a5dbfeda91c50abfb3d29a914a, {16'd22949, 16'd29577, 16'd63213, 16'd7896, 16'd6162, 16'd53150, 16'd25478, 16'd12629, 16'd34089, 16'd54747, 16'd43506, 16'd55327, 16'd6872, 16'd4805, 16'd35642, 16'd290, 16'd5, 16'd64163, 16'd30609, 16'd58487, 16'd52364, 16'd35213, 16'd60404, 16'd46991, 16'd24424, 16'd12446});
	test_expansion(128'h23e52b023299b96d10fb7a06b039b219, {16'd38619, 16'd58190, 16'd13751, 16'd22305, 16'd14270, 16'd45599, 16'd1267, 16'd41414, 16'd62358, 16'd29004, 16'd15888, 16'd55817, 16'd12240, 16'd25463, 16'd57138, 16'd9302, 16'd37740, 16'd24403, 16'd58251, 16'd9758, 16'd19170, 16'd8624, 16'd39181, 16'd27611, 16'd45512, 16'd10573});
	test_expansion(128'h2e64ce42cc52c09cf04e82f9e90d9475, {16'd55271, 16'd1426, 16'd33496, 16'd41843, 16'd5654, 16'd48970, 16'd5699, 16'd20253, 16'd33847, 16'd37264, 16'd61388, 16'd32778, 16'd34404, 16'd27655, 16'd13258, 16'd30165, 16'd65431, 16'd31810, 16'd17202, 16'd44717, 16'd28045, 16'd6734, 16'd5398, 16'd65442, 16'd35378, 16'd63882});
	test_expansion(128'h00409d50ccf8bd73f0746b5d1cbf4ae6, {16'd9642, 16'd13420, 16'd63917, 16'd14707, 16'd60632, 16'd63423, 16'd31035, 16'd54932, 16'd1402, 16'd24139, 16'd28488, 16'd31098, 16'd48273, 16'd7651, 16'd44036, 16'd52721, 16'd57887, 16'd51246, 16'd59371, 16'd57638, 16'd31794, 16'd34631, 16'd1960, 16'd46793, 16'd52367, 16'd53679});
	test_expansion(128'hffccaed94cf1cabacc7e85af723fbf59, {16'd62922, 16'd32217, 16'd14616, 16'd20641, 16'd24376, 16'd1823, 16'd59125, 16'd4712, 16'd42221, 16'd12708, 16'd25897, 16'd20168, 16'd44854, 16'd5989, 16'd13257, 16'd37578, 16'd41757, 16'd13760, 16'd32925, 16'd35509, 16'd7162, 16'd5154, 16'd20021, 16'd34667, 16'd18558, 16'd15165});
	test_expansion(128'h58190c783d104b2a33dccd6d1752282e, {16'd61276, 16'd54037, 16'd26469, 16'd35168, 16'd39315, 16'd8879, 16'd35495, 16'd18013, 16'd63356, 16'd29887, 16'd25645, 16'd59386, 16'd1970, 16'd45211, 16'd62405, 16'd16902, 16'd2938, 16'd6826, 16'd37557, 16'd48652, 16'd36206, 16'd39125, 16'd27483, 16'd56893, 16'd33302, 16'd58048});
	test_expansion(128'ha321d1d5102a5a594d1fd261d586aeb8, {16'd3421, 16'd45859, 16'd36279, 16'd27233, 16'd11083, 16'd20188, 16'd51578, 16'd38479, 16'd56969, 16'd21801, 16'd5725, 16'd44977, 16'd47264, 16'd10320, 16'd3264, 16'd35527, 16'd1375, 16'd46029, 16'd2003, 16'd54570, 16'd25621, 16'd7996, 16'd5980, 16'd9583, 16'd56661, 16'd43165});
	test_expansion(128'h513487af998d1e75a04a1b92e7f69b0f, {16'd51912, 16'd25611, 16'd2421, 16'd7491, 16'd48017, 16'd30212, 16'd53091, 16'd17861, 16'd44307, 16'd19870, 16'd64741, 16'd43484, 16'd48380, 16'd21644, 16'd36211, 16'd2339, 16'd11150, 16'd42104, 16'd34012, 16'd3163, 16'd39467, 16'd59373, 16'd12255, 16'd28732, 16'd17671, 16'd63528});
	test_expansion(128'h6c5fc31bc6424028bef01bbea7feef4b, {16'd3251, 16'd49615, 16'd8841, 16'd34452, 16'd3974, 16'd18612, 16'd29550, 16'd4637, 16'd1930, 16'd22523, 16'd36496, 16'd38804, 16'd29381, 16'd59021, 16'd24617, 16'd14297, 16'd40617, 16'd18326, 16'd8410, 16'd43653, 16'd32986, 16'd22915, 16'd54963, 16'd10825, 16'd25898, 16'd15901});
	test_expansion(128'hdc0e63f1db0ad2408baf26de7e3900d6, {16'd2713, 16'd11506, 16'd14117, 16'd61478, 16'd61359, 16'd41452, 16'd36998, 16'd65413, 16'd60448, 16'd28845, 16'd63364, 16'd63875, 16'd44901, 16'd38034, 16'd17568, 16'd61458, 16'd32746, 16'd62164, 16'd18998, 16'd63082, 16'd57217, 16'd25013, 16'd4440, 16'd28157, 16'd32839, 16'd33250});
	test_expansion(128'hd15f5cf3d44f3f6f3409267772cab0e2, {16'd46326, 16'd27563, 16'd31649, 16'd59137, 16'd60478, 16'd29904, 16'd30563, 16'd9996, 16'd49283, 16'd6685, 16'd10376, 16'd41226, 16'd13890, 16'd53896, 16'd62622, 16'd17974, 16'd28104, 16'd36090, 16'd48461, 16'd16206, 16'd32011, 16'd44733, 16'd9592, 16'd33357, 16'd16311, 16'd9177});
	test_expansion(128'h53dad7d241f76892a45f721dbd861950, {16'd44965, 16'd9623, 16'd53781, 16'd2283, 16'd14300, 16'd5636, 16'd60521, 16'd43809, 16'd65369, 16'd26002, 16'd13167, 16'd38495, 16'd50837, 16'd57135, 16'd44310, 16'd8398, 16'd45117, 16'd35858, 16'd3253, 16'd15015, 16'd26724, 16'd55014, 16'd26088, 16'd14093, 16'd54121, 16'd61371});
	test_expansion(128'hbf875c03a14d6d77c409b7777945dae1, {16'd54610, 16'd59526, 16'd59515, 16'd52249, 16'd50648, 16'd19697, 16'd45264, 16'd54271, 16'd385, 16'd44041, 16'd21321, 16'd56116, 16'd41490, 16'd28015, 16'd12213, 16'd8350, 16'd31615, 16'd14985, 16'd49914, 16'd31237, 16'd3861, 16'd50657, 16'd21608, 16'd10932, 16'd23261, 16'd29296});
	test_expansion(128'h62f3e969da090d9eba6bcdc622352f74, {16'd19839, 16'd55308, 16'd40781, 16'd58067, 16'd11109, 16'd542, 16'd5888, 16'd50198, 16'd7303, 16'd37723, 16'd61383, 16'd1622, 16'd54596, 16'd7658, 16'd37735, 16'd27191, 16'd10109, 16'd19623, 16'd42343, 16'd19965, 16'd32037, 16'd57838, 16'd20687, 16'd37893, 16'd46968, 16'd43178});
	test_expansion(128'h4113d67555e629a363cb296074fdc652, {16'd35757, 16'd13792, 16'd12942, 16'd41656, 16'd26610, 16'd18451, 16'd3379, 16'd38317, 16'd19946, 16'd36737, 16'd52080, 16'd44299, 16'd15686, 16'd23855, 16'd47460, 16'd23198, 16'd62703, 16'd9772, 16'd4419, 16'd33486, 16'd23352, 16'd13662, 16'd2, 16'd33142, 16'd3588, 16'd24809});
	test_expansion(128'hb8d998401d2ad3f239be7572ee492735, {16'd31582, 16'd29659, 16'd7750, 16'd28552, 16'd5569, 16'd61357, 16'd22899, 16'd16186, 16'd12018, 16'd21385, 16'd36988, 16'd28093, 16'd59330, 16'd51610, 16'd7427, 16'd669, 16'd36005, 16'd15853, 16'd12617, 16'd12393, 16'd53727, 16'd52902, 16'd47892, 16'd24574, 16'd21039, 16'd63556});
	test_expansion(128'h5351b11c59def87bd7a81f5f3756343e, {16'd41018, 16'd6464, 16'd464, 16'd5023, 16'd52028, 16'd35758, 16'd27246, 16'd30026, 16'd51226, 16'd55717, 16'd17414, 16'd3097, 16'd1111, 16'd12917, 16'd29094, 16'd26651, 16'd55842, 16'd53518, 16'd43607, 16'd64693, 16'd17044, 16'd6238, 16'd22860, 16'd61661, 16'd50572, 16'd34606});
	test_expansion(128'h1b98d047cfb344d15ff1bf109032ce11, {16'd63035, 16'd53397, 16'd50270, 16'd43840, 16'd10808, 16'd36733, 16'd51962, 16'd24241, 16'd56608, 16'd36389, 16'd1433, 16'd53647, 16'd20209, 16'd53585, 16'd64032, 16'd47033, 16'd55016, 16'd30255, 16'd62466, 16'd52156, 16'd44324, 16'd3051, 16'd20185, 16'd16091, 16'd26712, 16'd48076});
	test_expansion(128'h5ed686268e95441a58ef67c46e9bf353, {16'd38973, 16'd58131, 16'd54479, 16'd47048, 16'd37200, 16'd7427, 16'd12362, 16'd19187, 16'd65231, 16'd16769, 16'd8393, 16'd938, 16'd58988, 16'd28093, 16'd48408, 16'd57208, 16'd42127, 16'd60802, 16'd14979, 16'd25740, 16'd41896, 16'd41465, 16'd24826, 16'd23072, 16'd58949, 16'd24180});
	test_expansion(128'h5527a47925714d434aea225842875b8a, {16'd54492, 16'd64943, 16'd34396, 16'd12675, 16'd5989, 16'd46925, 16'd48033, 16'd64987, 16'd13971, 16'd25645, 16'd29200, 16'd20918, 16'd17941, 16'd58944, 16'd4981, 16'd26369, 16'd56153, 16'd45237, 16'd8245, 16'd16673, 16'd22966, 16'd10422, 16'd8317, 16'd55298, 16'd8116, 16'd53734});
	test_expansion(128'haedf421fc4eb271b9541d07ba37f93e2, {16'd58384, 16'd39561, 16'd61840, 16'd10119, 16'd53275, 16'd15868, 16'd16377, 16'd24955, 16'd13699, 16'd9971, 16'd3343, 16'd3226, 16'd16851, 16'd5598, 16'd25350, 16'd25707, 16'd32526, 16'd30524, 16'd7039, 16'd409, 16'd45325, 16'd21859, 16'd58371, 16'd12641, 16'd48184, 16'd25040});
	test_expansion(128'h38a1bb0ce94a6d64ba1462dcc5528351, {16'd18402, 16'd26863, 16'd47630, 16'd61040, 16'd18579, 16'd1966, 16'd20169, 16'd45566, 16'd12065, 16'd45411, 16'd58646, 16'd56082, 16'd33128, 16'd57549, 16'd57187, 16'd49207, 16'd45600, 16'd7597, 16'd5539, 16'd28269, 16'd20209, 16'd1779, 16'd49312, 16'd35967, 16'd51375, 16'd31794});
	test_expansion(128'h79d8e0b0e85727d27c10c659b3c80492, {16'd25231, 16'd53823, 16'd2169, 16'd50340, 16'd26139, 16'd9235, 16'd51552, 16'd36809, 16'd44202, 16'd36701, 16'd60844, 16'd62470, 16'd11768, 16'd60432, 16'd29601, 16'd54871, 16'd7314, 16'd62423, 16'd19649, 16'd33949, 16'd10508, 16'd61523, 16'd25775, 16'd47674, 16'd14225, 16'd33916});
	test_expansion(128'h7a61d1ef78f8ed173bf470d62a7f4cdc, {16'd4843, 16'd3454, 16'd17244, 16'd26486, 16'd63812, 16'd15444, 16'd10489, 16'd5156, 16'd8275, 16'd38253, 16'd7549, 16'd43292, 16'd43163, 16'd54367, 16'd8529, 16'd28276, 16'd39278, 16'd41674, 16'd60597, 16'd50413, 16'd8070, 16'd27396, 16'd24237, 16'd57139, 16'd63609, 16'd7400});
	test_expansion(128'h9ba2b15203d57d7cb68951448feb75dc, {16'd58767, 16'd42368, 16'd47105, 16'd10944, 16'd40034, 16'd24193, 16'd27461, 16'd50092, 16'd48242, 16'd17480, 16'd1454, 16'd45876, 16'd21686, 16'd56769, 16'd6520, 16'd62438, 16'd18263, 16'd23962, 16'd10911, 16'd21164, 16'd37055, 16'd58005, 16'd54796, 16'd24036, 16'd46517, 16'd4281});
	test_expansion(128'h226e1282d67b30d4806613d4b12337e0, {16'd31561, 16'd18046, 16'd7065, 16'd33547, 16'd49548, 16'd12489, 16'd13837, 16'd46758, 16'd3002, 16'd64471, 16'd20393, 16'd492, 16'd46793, 16'd17953, 16'd44127, 16'd34596, 16'd30486, 16'd40946, 16'd52378, 16'd24282, 16'd426, 16'd38642, 16'd39746, 16'd62229, 16'd52716, 16'd55460});
	test_expansion(128'h41a57cc5fa8ac67f654a2f048d34db17, {16'd14679, 16'd15790, 16'd44900, 16'd53189, 16'd58731, 16'd32329, 16'd13678, 16'd8917, 16'd29834, 16'd12817, 16'd62184, 16'd2486, 16'd23484, 16'd1466, 16'd25580, 16'd32101, 16'd37125, 16'd52452, 16'd34695, 16'd3314, 16'd59606, 16'd31465, 16'd40613, 16'd56273, 16'd6904, 16'd54791});
	test_expansion(128'hd521367565c0d43b81e9bcd5650a8f22, {16'd11089, 16'd24655, 16'd32148, 16'd35127, 16'd56609, 16'd28916, 16'd30651, 16'd34395, 16'd35502, 16'd48737, 16'd39595, 16'd16606, 16'd24191, 16'd13129, 16'd30561, 16'd17312, 16'd57829, 16'd10207, 16'd44697, 16'd50046, 16'd2119, 16'd18911, 16'd46701, 16'd39951, 16'd15020, 16'd50569});
	test_expansion(128'hf288f6b0a8bb7872a8174ba965fbb4f6, {16'd28610, 16'd28905, 16'd57776, 16'd55344, 16'd54422, 16'd18178, 16'd57692, 16'd54542, 16'd7540, 16'd32981, 16'd39142, 16'd39813, 16'd9133, 16'd46249, 16'd8808, 16'd50511, 16'd48092, 16'd29673, 16'd25035, 16'd59083, 16'd8418, 16'd24187, 16'd18839, 16'd60102, 16'd9056, 16'd42274});
	test_expansion(128'h6de2f4f4d33be53083b9a83ee753f6f3, {16'd51556, 16'd6208, 16'd52403, 16'd42615, 16'd6351, 16'd16449, 16'd34507, 16'd19541, 16'd2437, 16'd60625, 16'd57186, 16'd57193, 16'd46341, 16'd57812, 16'd23604, 16'd54983, 16'd14781, 16'd897, 16'd119, 16'd60782, 16'd35024, 16'd35570, 16'd40653, 16'd43298, 16'd13052, 16'd7879});
	test_expansion(128'hff8a68c2abbc03702c0c42faec6c8c90, {16'd33939, 16'd7214, 16'd6567, 16'd26093, 16'd811, 16'd2478, 16'd37943, 16'd35592, 16'd38551, 16'd4226, 16'd26796, 16'd18518, 16'd14427, 16'd28355, 16'd35814, 16'd45145, 16'd15582, 16'd36708, 16'd9469, 16'd1553, 16'd21442, 16'd46885, 16'd58201, 16'd51263, 16'd565, 16'd536});
	test_expansion(128'h50d0b79baaaa47a82119df3069d0d26a, {16'd30615, 16'd17394, 16'd4817, 16'd26431, 16'd56465, 16'd39054, 16'd7545, 16'd26, 16'd62127, 16'd21706, 16'd17518, 16'd7523, 16'd27661, 16'd42341, 16'd24882, 16'd9882, 16'd16832, 16'd56010, 16'd36642, 16'd53306, 16'd61757, 16'd12084, 16'd31612, 16'd49920, 16'd11865, 16'd58940});
	test_expansion(128'he5286e7539f279a8de5ce5139f63046f, {16'd38924, 16'd55827, 16'd9336, 16'd23979, 16'd54730, 16'd30578, 16'd43557, 16'd19865, 16'd32317, 16'd46045, 16'd64008, 16'd50387, 16'd58170, 16'd23125, 16'd4640, 16'd61859, 16'd18639, 16'd27749, 16'd64914, 16'd717, 16'd20108, 16'd52632, 16'd12322, 16'd34007, 16'd51338, 16'd46740});
	test_expansion(128'h5faf342acc71205314335fadf713c6af, {16'd3129, 16'd6506, 16'd25842, 16'd27985, 16'd35957, 16'd35398, 16'd41765, 16'd37462, 16'd23726, 16'd42732, 16'd24876, 16'd34973, 16'd30409, 16'd53765, 16'd60201, 16'd49339, 16'd59827, 16'd8268, 16'd42483, 16'd37495, 16'd40898, 16'd63383, 16'd17492, 16'd19737, 16'd20911, 16'd54506});
	test_expansion(128'hbec64178c8633b1da5e1f6e037fc6dd2, {16'd5573, 16'd9673, 16'd58962, 16'd13110, 16'd27912, 16'd60114, 16'd14157, 16'd12131, 16'd10709, 16'd60465, 16'd63308, 16'd8445, 16'd2043, 16'd29771, 16'd42609, 16'd34629, 16'd15678, 16'd46696, 16'd49109, 16'd28161, 16'd33867, 16'd53051, 16'd25770, 16'd24573, 16'd8078, 16'd52313});
	test_expansion(128'h7ad9b3164b3be90d01b646b6661808af, {16'd54707, 16'd25449, 16'd95, 16'd33622, 16'd62612, 16'd65239, 16'd47794, 16'd13374, 16'd42714, 16'd10745, 16'd40744, 16'd27515, 16'd35893, 16'd56201, 16'd1694, 16'd27859, 16'd61086, 16'd43461, 16'd47024, 16'd47209, 16'd29687, 16'd58852, 16'd29928, 16'd5230, 16'd36692, 16'd44818});
	test_expansion(128'h95f81ed4c8e1e6a25cf74424e80c486b, {16'd26931, 16'd37191, 16'd26459, 16'd707, 16'd22118, 16'd44510, 16'd46017, 16'd59472, 16'd65123, 16'd17926, 16'd62414, 16'd34886, 16'd49946, 16'd17780, 16'd53319, 16'd24721, 16'd9028, 16'd17311, 16'd35571, 16'd41783, 16'd34320, 16'd37954, 16'd61338, 16'd54172, 16'd55141, 16'd61979});
	test_expansion(128'hfe8d1a1b9bbfb1d474a48af7486505d1, {16'd55510, 16'd15041, 16'd46360, 16'd29434, 16'd7523, 16'd8407, 16'd52575, 16'd7553, 16'd57508, 16'd53543, 16'd64993, 16'd39586, 16'd45933, 16'd27099, 16'd5328, 16'd27791, 16'd17683, 16'd10791, 16'd60393, 16'd61803, 16'd2232, 16'd44064, 16'd24274, 16'd42918, 16'd61762, 16'd17483});
	test_expansion(128'h6dfe9b1afeda91193378a1e420501b72, {16'd7010, 16'd34613, 16'd20441, 16'd22466, 16'd48518, 16'd9434, 16'd4328, 16'd17408, 16'd38286, 16'd49987, 16'd18950, 16'd11713, 16'd36628, 16'd53438, 16'd17565, 16'd21455, 16'd12705, 16'd33905, 16'd8018, 16'd44121, 16'd33578, 16'd62649, 16'd53854, 16'd13053, 16'd51055, 16'd36208});
	test_expansion(128'h32ef04e1d6c770e41fe9dd52563cf76e, {16'd47641, 16'd26711, 16'd27580, 16'd3000, 16'd49130, 16'd57417, 16'd23840, 16'd1323, 16'd22391, 16'd37179, 16'd45211, 16'd56546, 16'd34493, 16'd58671, 16'd38995, 16'd26562, 16'd34196, 16'd9597, 16'd49521, 16'd52327, 16'd31786, 16'd60053, 16'd56588, 16'd19663, 16'd30296, 16'd10126});
	test_expansion(128'h4533b5e5fe40770f69ab3f46a15c57d5, {16'd9397, 16'd10728, 16'd92, 16'd64329, 16'd45272, 16'd44873, 16'd54010, 16'd46630, 16'd15638, 16'd404, 16'd62470, 16'd63725, 16'd19918, 16'd41309, 16'd17621, 16'd42064, 16'd24202, 16'd17206, 16'd32490, 16'd50850, 16'd17008, 16'd9116, 16'd3527, 16'd36315, 16'd10787, 16'd28828});
	test_expansion(128'hbd7dcc40dc49c897a0c24877600d503e, {16'd34462, 16'd60779, 16'd57030, 16'd57010, 16'd46454, 16'd30029, 16'd28758, 16'd4990, 16'd26746, 16'd26312, 16'd41463, 16'd1585, 16'd63794, 16'd14630, 16'd13417, 16'd31267, 16'd47533, 16'd51957, 16'd48843, 16'd34567, 16'd11394, 16'd55455, 16'd4055, 16'd39519, 16'd41905, 16'd7692});
	test_expansion(128'h83a0560cd246f707e369c6819ac4a217, {16'd22152, 16'd35770, 16'd23979, 16'd65400, 16'd50862, 16'd22938, 16'd37309, 16'd14639, 16'd59171, 16'd61620, 16'd64657, 16'd14087, 16'd61140, 16'd11327, 16'd29402, 16'd52052, 16'd144, 16'd53983, 16'd41406, 16'd268, 16'd45777, 16'd3478, 16'd19155, 16'd59314, 16'd11658, 16'd27210});
	test_expansion(128'h8487913a382eebbe2cbbf01a5d85649d, {16'd25326, 16'd64840, 16'd47204, 16'd8389, 16'd22893, 16'd57576, 16'd36587, 16'd3171, 16'd2789, 16'd16501, 16'd40371, 16'd35791, 16'd55827, 16'd33335, 16'd2471, 16'd4030, 16'd43212, 16'd48638, 16'd7414, 16'd63432, 16'd59078, 16'd20552, 16'd37714, 16'd51672, 16'd15666, 16'd53957});
	test_expansion(128'hc5d57a2548fcfa5a671330f4454477c7, {16'd28172, 16'd18690, 16'd38922, 16'd44315, 16'd43456, 16'd3377, 16'd22850, 16'd50865, 16'd5222, 16'd41741, 16'd61258, 16'd47058, 16'd33157, 16'd36642, 16'd27214, 16'd981, 16'd7388, 16'd60686, 16'd9002, 16'd50870, 16'd16574, 16'd33910, 16'd62461, 16'd10448, 16'd51916, 16'd19659});
	test_expansion(128'h657f0e724a340f0a65f2061cac01f84a, {16'd59258, 16'd19776, 16'd935, 16'd31917, 16'd28431, 16'd26693, 16'd41373, 16'd1350, 16'd50800, 16'd11401, 16'd6542, 16'd34200, 16'd61592, 16'd4819, 16'd57727, 16'd1289, 16'd46426, 16'd55497, 16'd50323, 16'd64952, 16'd31784, 16'd47611, 16'd60253, 16'd39220, 16'd26067, 16'd19102});
	test_expansion(128'h2ce4592613bb33782abdd88d739951c2, {16'd19003, 16'd35466, 16'd25814, 16'd42785, 16'd10878, 16'd47669, 16'd24912, 16'd42976, 16'd64172, 16'd18710, 16'd2549, 16'd16432, 16'd12974, 16'd24262, 16'd45417, 16'd24846, 16'd59751, 16'd63599, 16'd48998, 16'd54364, 16'd17305, 16'd61864, 16'd56832, 16'd4540, 16'd57795, 16'd26587});
	test_expansion(128'h2a6cfbc4bf2979872a00af74ad438eb8, {16'd56050, 16'd11853, 16'd38926, 16'd24825, 16'd13930, 16'd61998, 16'd62342, 16'd23842, 16'd63894, 16'd800, 16'd38872, 16'd33780, 16'd5940, 16'd10904, 16'd21168, 16'd44464, 16'd54418, 16'd63744, 16'd32069, 16'd41075, 16'd29918, 16'd20360, 16'd17760, 16'd47966, 16'd52100, 16'd33636});
	test_expansion(128'h798c734fd439eb629d6f12ce3ac8cd07, {16'd16722, 16'd31613, 16'd29338, 16'd52958, 16'd43626, 16'd31475, 16'd19777, 16'd58943, 16'd64773, 16'd35246, 16'd48630, 16'd33574, 16'd19612, 16'd48193, 16'd40473, 16'd50165, 16'd17348, 16'd13367, 16'd54814, 16'd57221, 16'd53372, 16'd55758, 16'd22228, 16'd63326, 16'd58615, 16'd35172});
	test_expansion(128'h6cbc4bd639b6fb6d1434d08e3a74858b, {16'd14978, 16'd6631, 16'd1975, 16'd50261, 16'd20258, 16'd13625, 16'd2308, 16'd54148, 16'd851, 16'd33097, 16'd39377, 16'd53284, 16'd49333, 16'd44659, 16'd46222, 16'd17614, 16'd60921, 16'd43689, 16'd2760, 16'd27042, 16'd58972, 16'd14280, 16'd50742, 16'd6171, 16'd47589, 16'd43749});
	test_expansion(128'h291c7d1e30673cbae96ff9aa986f59e2, {16'd11207, 16'd24893, 16'd13656, 16'd4549, 16'd16748, 16'd44802, 16'd21952, 16'd49089, 16'd65039, 16'd7800, 16'd54569, 16'd3590, 16'd25397, 16'd12341, 16'd62350, 16'd29229, 16'd61026, 16'd51582, 16'd18361, 16'd19885, 16'd21810, 16'd57506, 16'd10111, 16'd38770, 16'd27799, 16'd30489});
	test_expansion(128'h8005dbf6db67a72edec0990a811a1f6f, {16'd19655, 16'd3472, 16'd2853, 16'd29205, 16'd20853, 16'd41001, 16'd19109, 16'd64603, 16'd13631, 16'd24002, 16'd39753, 16'd49441, 16'd53197, 16'd35352, 16'd61224, 16'd6372, 16'd8234, 16'd14264, 16'd36159, 16'd31886, 16'd40253, 16'd47482, 16'd9418, 16'd2796, 16'd25605, 16'd43987});
	test_expansion(128'h35997ef589340c66f9a075760c539ff3, {16'd56482, 16'd3111, 16'd54285, 16'd64399, 16'd38137, 16'd25558, 16'd8331, 16'd33129, 16'd1690, 16'd33397, 16'd51225, 16'd42591, 16'd2637, 16'd51788, 16'd37065, 16'd7764, 16'd24975, 16'd25571, 16'd21056, 16'd37854, 16'd7711, 16'd32090, 16'd52702, 16'd5352, 16'd32510, 16'd46522});
	test_expansion(128'hafc074fdac25bb2d271c6bc36ab2d27c, {16'd63372, 16'd4174, 16'd25940, 16'd44547, 16'd63793, 16'd16568, 16'd26373, 16'd21319, 16'd64963, 16'd22482, 16'd41262, 16'd59583, 16'd3869, 16'd29191, 16'd16242, 16'd15673, 16'd55224, 16'd65379, 16'd50178, 16'd42968, 16'd40523, 16'd63076, 16'd5439, 16'd60194, 16'd35211, 16'd16179});
	test_expansion(128'haeeef6ad330e3b046718e9e89932a86a, {16'd28939, 16'd13543, 16'd48117, 16'd59624, 16'd12121, 16'd48296, 16'd25476, 16'd6861, 16'd59433, 16'd40630, 16'd20748, 16'd11383, 16'd16917, 16'd11129, 16'd21640, 16'd62265, 16'd43937, 16'd6026, 16'd50850, 16'd51981, 16'd55527, 16'd4130, 16'd4607, 16'd1933, 16'd24881, 16'd13337});
	test_expansion(128'hdf14bb2d97963fc94eed056a59c9ec34, {16'd44432, 16'd40043, 16'd13265, 16'd29446, 16'd64350, 16'd58879, 16'd51170, 16'd29306, 16'd26671, 16'd11098, 16'd54051, 16'd47270, 16'd33732, 16'd2213, 16'd19965, 16'd24825, 16'd62890, 16'd21130, 16'd4814, 16'd13587, 16'd20887, 16'd42038, 16'd38179, 16'd16698, 16'd4519, 16'd50644});
	test_expansion(128'h6619ac82a7521fd938aba2bdfdabd364, {16'd24095, 16'd11927, 16'd24926, 16'd16301, 16'd35430, 16'd38647, 16'd18484, 16'd15876, 16'd64514, 16'd9650, 16'd41330, 16'd8145, 16'd46114, 16'd42258, 16'd2079, 16'd24830, 16'd24614, 16'd26577, 16'd8441, 16'd54422, 16'd49746, 16'd23770, 16'd47096, 16'd16868, 16'd20367, 16'd8667});
	test_expansion(128'hf083f112857ae703e870ec2d0a465fe4, {16'd52622, 16'd30014, 16'd59002, 16'd1281, 16'd50563, 16'd33707, 16'd32457, 16'd18494, 16'd7645, 16'd30929, 16'd41504, 16'd34423, 16'd5670, 16'd51689, 16'd55304, 16'd1812, 16'd8524, 16'd34571, 16'd45634, 16'd10884, 16'd31317, 16'd25773, 16'd51963, 16'd33831, 16'd38199, 16'd10147});
	test_expansion(128'hd5b298c2c56c2a36fe9113b6f47d8485, {16'd42739, 16'd6927, 16'd61139, 16'd38856, 16'd48544, 16'd40646, 16'd4022, 16'd13508, 16'd57007, 16'd45640, 16'd22186, 16'd33753, 16'd61818, 16'd34269, 16'd43982, 16'd50069, 16'd128, 16'd53362, 16'd30011, 16'd780, 16'd52156, 16'd53410, 16'd18659, 16'd4976, 16'd18363, 16'd51678});
	test_expansion(128'h4749248c590e595eed4fdea3dcc1e0da, {16'd32505, 16'd51379, 16'd58764, 16'd19094, 16'd48870, 16'd53648, 16'd42790, 16'd20230, 16'd6092, 16'd22182, 16'd56147, 16'd64095, 16'd12025, 16'd29472, 16'd24876, 16'd59965, 16'd3250, 16'd56270, 16'd20218, 16'd15396, 16'd9559, 16'd64738, 16'd7867, 16'd50195, 16'd7043, 16'd19870});
	test_expansion(128'hba5b5fe7c9cadbc10458786b9f1a8bdd, {16'd19969, 16'd29808, 16'd9156, 16'd61157, 16'd39998, 16'd27380, 16'd55969, 16'd44725, 16'd61343, 16'd62863, 16'd28796, 16'd52081, 16'd15302, 16'd54456, 16'd57717, 16'd14250, 16'd50451, 16'd54861, 16'd2385, 16'd46676, 16'd46453, 16'd47444, 16'd56384, 16'd56330, 16'd30879, 16'd39876});
	test_expansion(128'h0a5ac991ea0562e4711430472a4de0e0, {16'd6301, 16'd39264, 16'd4251, 16'd48301, 16'd34608, 16'd53627, 16'd45489, 16'd16045, 16'd866, 16'd19558, 16'd52701, 16'd29388, 16'd36631, 16'd63345, 16'd59780, 16'd43231, 16'd58408, 16'd30258, 16'd26826, 16'd36910, 16'd1410, 16'd5380, 16'd53821, 16'd40862, 16'd33696, 16'd14237});
	test_expansion(128'h3eed239178327caaeec1cd13276d985e, {16'd11025, 16'd12855, 16'd58958, 16'd17032, 16'd44131, 16'd26976, 16'd35758, 16'd9397, 16'd33035, 16'd35397, 16'd36238, 16'd43843, 16'd2752, 16'd32696, 16'd16520, 16'd36083, 16'd33528, 16'd16800, 16'd8075, 16'd59060, 16'd33568, 16'd55276, 16'd50875, 16'd230, 16'd50451, 16'd16363});
	test_expansion(128'hda7d5833f320260a55bd597d56eacd9c, {16'd39810, 16'd24320, 16'd20037, 16'd27305, 16'd45715, 16'd21832, 16'd44443, 16'd33315, 16'd3554, 16'd34605, 16'd6944, 16'd53252, 16'd45157, 16'd888, 16'd43000, 16'd17468, 16'd25550, 16'd45304, 16'd51642, 16'd15196, 16'd15661, 16'd40428, 16'd43869, 16'd32882, 16'd16932, 16'd34290});
	test_expansion(128'h7134a35420e256d7d1d02e97c222fbd1, {16'd52181, 16'd39869, 16'd19280, 16'd50498, 16'd52063, 16'd1424, 16'd46421, 16'd25814, 16'd63017, 16'd58530, 16'd35902, 16'd41191, 16'd49616, 16'd32406, 16'd14328, 16'd61702, 16'd64764, 16'd31195, 16'd13816, 16'd60418, 16'd55655, 16'd2629, 16'd29014, 16'd16433, 16'd45218, 16'd18333});
	test_expansion(128'h51a8ad6b5339566ef8ea5798d571f103, {16'd19051, 16'd29849, 16'd11196, 16'd35524, 16'd46183, 16'd9383, 16'd3370, 16'd18356, 16'd40057, 16'd43164, 16'd36941, 16'd63022, 16'd64961, 16'd35521, 16'd4787, 16'd37270, 16'd12829, 16'd35971, 16'd11388, 16'd7261, 16'd7932, 16'd4543, 16'd36024, 16'd62902, 16'd33803, 16'd6095});
	test_expansion(128'h103b5139d0d496550dca418ef9f312cc, {16'd13248, 16'd7357, 16'd54125, 16'd1049, 16'd42550, 16'd3395, 16'd20580, 16'd16198, 16'd9988, 16'd63137, 16'd15550, 16'd24707, 16'd47511, 16'd51217, 16'd48314, 16'd35657, 16'd7992, 16'd55694, 16'd2737, 16'd46163, 16'd12896, 16'd16405, 16'd15427, 16'd6983, 16'd21344, 16'd65491});
	test_expansion(128'h30b4e46fedfaafe6b0a97af24490f860, {16'd23031, 16'd14603, 16'd5102, 16'd32815, 16'd2427, 16'd21459, 16'd18202, 16'd35016, 16'd32950, 16'd945, 16'd3363, 16'd44311, 16'd43331, 16'd17709, 16'd10314, 16'd11455, 16'd59659, 16'd32608, 16'd6214, 16'd1056, 16'd28925, 16'd15334, 16'd19810, 16'd52788, 16'd33375, 16'd50329});
	test_expansion(128'hf9251e6f33d73362898c374139600304, {16'd43514, 16'd10573, 16'd20514, 16'd3044, 16'd2470, 16'd32421, 16'd27014, 16'd13530, 16'd36009, 16'd31809, 16'd39552, 16'd61149, 16'd50606, 16'd41751, 16'd51339, 16'd8737, 16'd60984, 16'd17973, 16'd30481, 16'd48923, 16'd50811, 16'd18718, 16'd50852, 16'd48857, 16'd35951, 16'd6099});
	test_expansion(128'h58ec6fb25879cf6376bcac6726f9f139, {16'd32050, 16'd31786, 16'd8714, 16'd22245, 16'd8181, 16'd6487, 16'd45225, 16'd327, 16'd31658, 16'd14802, 16'd13660, 16'd50904, 16'd3275, 16'd579, 16'd46871, 16'd2347, 16'd34587, 16'd24623, 16'd13156, 16'd39551, 16'd24632, 16'd14057, 16'd10195, 16'd11382, 16'd4887, 16'd30704});
	test_expansion(128'h760e10975f43cf2cffc9160dc68062e5, {16'd24740, 16'd11650, 16'd16158, 16'd23451, 16'd32879, 16'd18474, 16'd5762, 16'd33874, 16'd41891, 16'd4128, 16'd41583, 16'd49083, 16'd19781, 16'd17704, 16'd44783, 16'd13044, 16'd39803, 16'd61610, 16'd5232, 16'd23335, 16'd20916, 16'd60752, 16'd30427, 16'd9342, 16'd48698, 16'd57291});
	test_expansion(128'h8df09088c0f64a9f677699541dad5c82, {16'd13883, 16'd23615, 16'd12762, 16'd1795, 16'd19007, 16'd20058, 16'd5305, 16'd53387, 16'd18773, 16'd52105, 16'd34011, 16'd11640, 16'd41820, 16'd1666, 16'd57813, 16'd59109, 16'd57238, 16'd2183, 16'd46196, 16'd61667, 16'd44527, 16'd43421, 16'd11664, 16'd33603, 16'd56312, 16'd9051});
	test_expansion(128'h5f33779493956b715d00f7899f2ba639, {16'd31808, 16'd35137, 16'd49138, 16'd42630, 16'd39185, 16'd54535, 16'd56377, 16'd53057, 16'd34710, 16'd41533, 16'd48137, 16'd36050, 16'd16240, 16'd33257, 16'd61016, 16'd58257, 16'd3843, 16'd56421, 16'd35742, 16'd60842, 16'd41366, 16'd1700, 16'd3304, 16'd5920, 16'd40182, 16'd10449});
	test_expansion(128'hfcb6cad86d195b587d23fd758a5e47e1, {16'd23294, 16'd63866, 16'd40262, 16'd31366, 16'd46024, 16'd56100, 16'd45149, 16'd18745, 16'd19741, 16'd6746, 16'd20784, 16'd23829, 16'd5076, 16'd34705, 16'd40619, 16'd60725, 16'd58566, 16'd58133, 16'd51252, 16'd47671, 16'd9325, 16'd32819, 16'd18379, 16'd40969, 16'd22700, 16'd31859});
	test_expansion(128'h1ff91edb03bfa0387ccb700a1322c40b, {16'd53042, 16'd37116, 16'd53434, 16'd64171, 16'd32618, 16'd58400, 16'd60426, 16'd53711, 16'd39460, 16'd8198, 16'd27446, 16'd12946, 16'd37793, 16'd53169, 16'd51924, 16'd4648, 16'd24295, 16'd10889, 16'd21971, 16'd11703, 16'd2009, 16'd52958, 16'd23464, 16'd46307, 16'd39891, 16'd36735});
	test_expansion(128'hc95f4ba7d484dbb858eed67f4315698c, {16'd50419, 16'd55843, 16'd25443, 16'd6152, 16'd35492, 16'd3122, 16'd16906, 16'd55133, 16'd46159, 16'd33471, 16'd23953, 16'd14258, 16'd52845, 16'd17845, 16'd52304, 16'd60320, 16'd50346, 16'd11066, 16'd774, 16'd50371, 16'd17497, 16'd39882, 16'd54667, 16'd11867, 16'd43609, 16'd23950});
	test_expansion(128'h41f89381199a2f83ede1207c90d3200e, {16'd61137, 16'd14511, 16'd52508, 16'd42297, 16'd58137, 16'd38338, 16'd58332, 16'd25587, 16'd64065, 16'd38025, 16'd30140, 16'd41813, 16'd53648, 16'd5486, 16'd41133, 16'd20792, 16'd4481, 16'd64788, 16'd41495, 16'd11663, 16'd65029, 16'd34291, 16'd59651, 16'd58416, 16'd31093, 16'd58636});
	test_expansion(128'h613fb45cf07dd8dabd62027f2e441bb9, {16'd25846, 16'd35293, 16'd5728, 16'd55963, 16'd43501, 16'd26375, 16'd54125, 16'd59310, 16'd62959, 16'd34375, 16'd1102, 16'd54212, 16'd10371, 16'd56043, 16'd34569, 16'd29965, 16'd18799, 16'd27188, 16'd56116, 16'd57861, 16'd1816, 16'd35582, 16'd3322, 16'd7516, 16'd37605, 16'd22893});
	test_expansion(128'h82b286ebb80418dbf4a829b37cbebbda, {16'd42458, 16'd51396, 16'd46447, 16'd29762, 16'd53619, 16'd13748, 16'd22598, 16'd44627, 16'd19006, 16'd48975, 16'd22719, 16'd9351, 16'd1072, 16'd1196, 16'd15492, 16'd63834, 16'd23437, 16'd18669, 16'd64432, 16'd38993, 16'd50405, 16'd37286, 16'd58261, 16'd5714, 16'd47060, 16'd41638});
	test_expansion(128'h87ad36513596b9181648b8a216d70e66, {16'd6330, 16'd14109, 16'd5822, 16'd3096, 16'd47731, 16'd59251, 16'd23921, 16'd29044, 16'd55235, 16'd40399, 16'd22394, 16'd53946, 16'd11307, 16'd33711, 16'd18030, 16'd64423, 16'd2634, 16'd30291, 16'd30870, 16'd53902, 16'd4597, 16'd64343, 16'd21679, 16'd4905, 16'd60551, 16'd55224});
	test_expansion(128'hb9243bf17189ca5723be425b04f6151f, {16'd50494, 16'd60964, 16'd15135, 16'd44213, 16'd5133, 16'd33820, 16'd30101, 16'd45276, 16'd52780, 16'd12973, 16'd59022, 16'd58954, 16'd23778, 16'd3592, 16'd50260, 16'd10140, 16'd28322, 16'd5205, 16'd51280, 16'd14396, 16'd64168, 16'd33991, 16'd25699, 16'd58545, 16'd2098, 16'd37207});
	test_expansion(128'h5fedcd3316576093ee8bcd654599204b, {16'd45087, 16'd27791, 16'd54246, 16'd2081, 16'd39457, 16'd41840, 16'd17611, 16'd56388, 16'd935, 16'd27702, 16'd32348, 16'd58491, 16'd44620, 16'd6775, 16'd8785, 16'd56236, 16'd54171, 16'd38705, 16'd5647, 16'd29001, 16'd31650, 16'd58799, 16'd22602, 16'd64412, 16'd48400, 16'd8118});
	test_expansion(128'h0ed840d03105471e759a1dff3248ba01, {16'd33345, 16'd33689, 16'd5280, 16'd51420, 16'd32304, 16'd10702, 16'd18332, 16'd40244, 16'd13273, 16'd34348, 16'd7368, 16'd38954, 16'd60754, 16'd5431, 16'd1154, 16'd56479, 16'd42225, 16'd19617, 16'd8380, 16'd43265, 16'd35988, 16'd42401, 16'd2061, 16'd1086, 16'd44929, 16'd41950});
	test_expansion(128'h4475585c596cc3ce2852b2a5980388b7, {16'd7533, 16'd23258, 16'd46361, 16'd46704, 16'd45895, 16'd15766, 16'd60644, 16'd47679, 16'd4322, 16'd36407, 16'd34486, 16'd51500, 16'd59482, 16'd40185, 16'd36591, 16'd14846, 16'd14654, 16'd19787, 16'd18493, 16'd53503, 16'd746, 16'd26938, 16'd36175, 16'd19217, 16'd24457, 16'd49525});
	test_expansion(128'h745608bbc2a5b3095c8ae92cc189f845, {16'd63139, 16'd584, 16'd20094, 16'd25282, 16'd52841, 16'd32663, 16'd32023, 16'd6910, 16'd48016, 16'd25692, 16'd46460, 16'd12713, 16'd1916, 16'd17574, 16'd32365, 16'd57910, 16'd41399, 16'd42147, 16'd29073, 16'd26728, 16'd3695, 16'd16891, 16'd20362, 16'd33099, 16'd54451, 16'd10091});
	test_expansion(128'h28bc0ebc204257804f3b9329aa408e83, {16'd42773, 16'd6023, 16'd18979, 16'd39122, 16'd38149, 16'd35594, 16'd6923, 16'd12406, 16'd2569, 16'd49235, 16'd54031, 16'd21435, 16'd32921, 16'd58202, 16'd15240, 16'd19859, 16'd15356, 16'd605, 16'd4050, 16'd14433, 16'd43628, 16'd11033, 16'd64142, 16'd29192, 16'd60288, 16'd6657});
	test_expansion(128'h40dbbe4109a17728ffe9ac6ee2adc17e, {16'd46720, 16'd8594, 16'd22520, 16'd31656, 16'd444, 16'd8705, 16'd10219, 16'd60314, 16'd57101, 16'd41704, 16'd11789, 16'd37638, 16'd13102, 16'd34699, 16'd35066, 16'd32183, 16'd2129, 16'd25740, 16'd33317, 16'd43162, 16'd56573, 16'd37381, 16'd60375, 16'd57288, 16'd57791, 16'd26501});
	test_expansion(128'h483763af6497c71d7ed89cad19bbdd7e, {16'd20587, 16'd45663, 16'd51041, 16'd57685, 16'd36965, 16'd17964, 16'd43556, 16'd51406, 16'd32837, 16'd13396, 16'd40178, 16'd36720, 16'd35957, 16'd54838, 16'd10934, 16'd56069, 16'd32279, 16'd64434, 16'd18668, 16'd13124, 16'd48339, 16'd64549, 16'd56223, 16'd17556, 16'd56794, 16'd22721});
	test_expansion(128'hf958bfb39f9588ee91d5a0943f608274, {16'd2440, 16'd64315, 16'd12053, 16'd24380, 16'd10656, 16'd3107, 16'd37395, 16'd27329, 16'd18995, 16'd26554, 16'd58635, 16'd25271, 16'd14899, 16'd41218, 16'd7953, 16'd18678, 16'd20315, 16'd28561, 16'd55533, 16'd59657, 16'd21550, 16'd27766, 16'd40128, 16'd41012, 16'd43454, 16'd47310});
	test_expansion(128'h9ce058ad99e1a9b6071594535c0b03d9, {16'd30036, 16'd11792, 16'd59829, 16'd7315, 16'd18174, 16'd45739, 16'd1766, 16'd12328, 16'd1208, 16'd62723, 16'd25773, 16'd46937, 16'd5027, 16'd759, 16'd61726, 16'd22011, 16'd35511, 16'd14842, 16'd51726, 16'd7535, 16'd37241, 16'd2821, 16'd54890, 16'd9584, 16'd11154, 16'd1065});
	test_expansion(128'h2e1c666c2632a1082bb441712dc52d7d, {16'd33493, 16'd19125, 16'd5048, 16'd33161, 16'd25157, 16'd61944, 16'd48778, 16'd57878, 16'd51863, 16'd33128, 16'd26865, 16'd29736, 16'd5580, 16'd22187, 16'd46781, 16'd15224, 16'd41357, 16'd64394, 16'd661, 16'd52020, 16'd16717, 16'd64895, 16'd24512, 16'd65418, 16'd48888, 16'd41783});
	test_expansion(128'h531f3b0800ff77d54a0aab61917e18f6, {16'd4277, 16'd54652, 16'd4531, 16'd52148, 16'd64264, 16'd22888, 16'd9848, 16'd61112, 16'd8715, 16'd51212, 16'd52542, 16'd38844, 16'd28545, 16'd39733, 16'd28050, 16'd63933, 16'd32423, 16'd23261, 16'd35490, 16'd34694, 16'd35234, 16'd31354, 16'd40995, 16'd46609, 16'd24204, 16'd27977});
	test_expansion(128'h837d0f5eaf0c621b06534d1f442327a7, {16'd7192, 16'd52509, 16'd26552, 16'd34925, 16'd8822, 16'd6567, 16'd46003, 16'd13573, 16'd25227, 16'd18169, 16'd28747, 16'd21073, 16'd37653, 16'd6665, 16'd56908, 16'd7273, 16'd23071, 16'd21594, 16'd3575, 16'd55530, 16'd5248, 16'd52219, 16'd13189, 16'd48688, 16'd21042, 16'd43200});
	test_expansion(128'h8ce17f8f50dc7cd4a7d76a7a9e397d5c, {16'd33759, 16'd44832, 16'd35049, 16'd17048, 16'd40842, 16'd55826, 16'd33114, 16'd39940, 16'd30322, 16'd19691, 16'd27742, 16'd4633, 16'd36645, 16'd3887, 16'd51156, 16'd17311, 16'd28830, 16'd16411, 16'd23328, 16'd25908, 16'd40750, 16'd32429, 16'd13753, 16'd37706, 16'd46357, 16'd31248});
	test_expansion(128'h3baeb25c2d48db2ca55d5e4185cdc6cd, {16'd21230, 16'd54398, 16'd20925, 16'd55, 16'd4351, 16'd54607, 16'd12546, 16'd40673, 16'd50157, 16'd59533, 16'd23028, 16'd21773, 16'd6157, 16'd28964, 16'd58889, 16'd60389, 16'd58623, 16'd11110, 16'd37523, 16'd60274, 16'd7108, 16'd6588, 16'd25997, 16'd18660, 16'd58582, 16'd32813});
	test_expansion(128'h4375c4fcfdfdef18346a17804a4e18ce, {16'd38175, 16'd39786, 16'd30790, 16'd14948, 16'd22320, 16'd21068, 16'd56191, 16'd7921, 16'd26314, 16'd35823, 16'd18701, 16'd25936, 16'd55641, 16'd36475, 16'd2709, 16'd46930, 16'd16011, 16'd12155, 16'd48987, 16'd40200, 16'd33709, 16'd41435, 16'd7048, 16'd41639, 16'd24358, 16'd42084});
	test_expansion(128'hcc23ee1c7f4cbfa7cbc1565dd538ad30, {16'd10546, 16'd40891, 16'd15039, 16'd29779, 16'd15203, 16'd22903, 16'd10294, 16'd27477, 16'd35809, 16'd6625, 16'd11902, 16'd47603, 16'd580, 16'd61563, 16'd36352, 16'd13071, 16'd16008, 16'd46084, 16'd33729, 16'd23137, 16'd57009, 16'd40926, 16'd60435, 16'd54736, 16'd12990, 16'd46252});
	test_expansion(128'hd445355ebc565100640f17deea9d4a52, {16'd58150, 16'd22800, 16'd14689, 16'd58298, 16'd27506, 16'd59794, 16'd4605, 16'd45729, 16'd5992, 16'd1568, 16'd60837, 16'd22778, 16'd41621, 16'd55172, 16'd21770, 16'd40446, 16'd32584, 16'd968, 16'd40241, 16'd64352, 16'd55188, 16'd7857, 16'd57438, 16'd28590, 16'd54456, 16'd30709});
	test_expansion(128'h53bf07d5e6277438f620f7dfc6e9d3b0, {16'd3425, 16'd34325, 16'd40310, 16'd65344, 16'd3611, 16'd20587, 16'd12010, 16'd39481, 16'd38136, 16'd18699, 16'd58468, 16'd8463, 16'd33968, 16'd60101, 16'd2593, 16'd44813, 16'd29439, 16'd47059, 16'd49469, 16'd2121, 16'd47036, 16'd37207, 16'd53729, 16'd43098, 16'd46889, 16'd44424});
	test_expansion(128'h382b4335dbdad87587d1d3f1380a9d89, {16'd40732, 16'd53002, 16'd44765, 16'd3037, 16'd22092, 16'd904, 16'd23091, 16'd130, 16'd12881, 16'd27190, 16'd9086, 16'd25731, 16'd17687, 16'd58992, 16'd28003, 16'd50911, 16'd59260, 16'd51375, 16'd55528, 16'd12133, 16'd31957, 16'd29639, 16'd40045, 16'd23209, 16'd36469, 16'd37436});
	test_expansion(128'ha5fd0583279a128f193ea55304295b7a, {16'd65107, 16'd15474, 16'd18224, 16'd32190, 16'd892, 16'd13529, 16'd60697, 16'd62579, 16'd32170, 16'd24553, 16'd33281, 16'd42681, 16'd55987, 16'd10091, 16'd44931, 16'd57587, 16'd18470, 16'd51049, 16'd39270, 16'd9057, 16'd46722, 16'd48661, 16'd54379, 16'd44182, 16'd47709, 16'd14774});
	test_expansion(128'h2981f0755d0089bd4e0c87f1db7fd2a0, {16'd8522, 16'd55062, 16'd56723, 16'd41469, 16'd29221, 16'd34964, 16'd6902, 16'd287, 16'd58344, 16'd32430, 16'd53167, 16'd13467, 16'd37292, 16'd1609, 16'd19153, 16'd60596, 16'd26912, 16'd56459, 16'd16844, 16'd64063, 16'd38668, 16'd55935, 16'd31049, 16'd39961, 16'd34164, 16'd58166});
	test_expansion(128'he81f018642abb8dec2e1912ab20a29db, {16'd30439, 16'd56738, 16'd56933, 16'd30996, 16'd32844, 16'd36984, 16'd49981, 16'd33350, 16'd53059, 16'd5056, 16'd40018, 16'd41288, 16'd4468, 16'd29913, 16'd59093, 16'd47601, 16'd17147, 16'd54960, 16'd27466, 16'd10752, 16'd21644, 16'd65492, 16'd45135, 16'd4919, 16'd53641, 16'd20649});
	test_expansion(128'h336b56b4b43756219e60bf5a0743fb33, {16'd7039, 16'd22422, 16'd32921, 16'd60326, 16'd48629, 16'd50376, 16'd19622, 16'd25282, 16'd30727, 16'd37238, 16'd20143, 16'd3552, 16'd30949, 16'd32900, 16'd31583, 16'd43214, 16'd18373, 16'd40453, 16'd13553, 16'd28235, 16'd39674, 16'd20448, 16'd22256, 16'd21870, 16'd63965, 16'd10241});
	test_expansion(128'h8febd4255e0ddc967077d9ec83b81616, {16'd31370, 16'd57864, 16'd53392, 16'd64174, 16'd47443, 16'd17239, 16'd12159, 16'd1949, 16'd17029, 16'd27475, 16'd61555, 16'd16549, 16'd11366, 16'd58110, 16'd3918, 16'd48461, 16'd65410, 16'd24978, 16'd3033, 16'd4147, 16'd42599, 16'd50915, 16'd43975, 16'd27152, 16'd49063, 16'd14108});
	test_expansion(128'he4f7dccd80754f459b4c40a434214258, {16'd48328, 16'd32662, 16'd3295, 16'd34902, 16'd16321, 16'd41047, 16'd42175, 16'd41851, 16'd62838, 16'd63240, 16'd45388, 16'd10264, 16'd61126, 16'd52376, 16'd51542, 16'd32558, 16'd30243, 16'd1273, 16'd49464, 16'd7773, 16'd14699, 16'd10378, 16'd21251, 16'd25879, 16'd4384, 16'd17282});
	test_expansion(128'ha218fb5b28ae4c83af14694c4ad92daf, {16'd23459, 16'd27060, 16'd51539, 16'd2726, 16'd53523, 16'd42414, 16'd2162, 16'd50830, 16'd8059, 16'd35180, 16'd54763, 16'd46920, 16'd62853, 16'd18042, 16'd20156, 16'd28613, 16'd54465, 16'd8700, 16'd5960, 16'd36767, 16'd31940, 16'd18057, 16'd39764, 16'd11789, 16'd23496, 16'd33975});
	test_expansion(128'ha42e6d8b85e6e27f29869939591a9fbc, {16'd40920, 16'd9285, 16'd10551, 16'd9849, 16'd27992, 16'd38658, 16'd18161, 16'd50474, 16'd45388, 16'd60413, 16'd5899, 16'd29038, 16'd50889, 16'd32193, 16'd41862, 16'd63514, 16'd12148, 16'd11240, 16'd36608, 16'd51687, 16'd37982, 16'd10338, 16'd18919, 16'd60522, 16'd62227, 16'd50762});
	test_expansion(128'he3935790ca42d325aee7066301b41a1f, {16'd33585, 16'd7968, 16'd44169, 16'd64472, 16'd26880, 16'd7752, 16'd33127, 16'd43714, 16'd43952, 16'd10934, 16'd65119, 16'd33208, 16'd2209, 16'd36955, 16'd31305, 16'd32569, 16'd48395, 16'd61542, 16'd39461, 16'd21656, 16'd53875, 16'd51439, 16'd60847, 16'd45093, 16'd13805, 16'd53711});
	test_expansion(128'h884997cc0392396b0c11717cbaa47ec1, {16'd28518, 16'd50438, 16'd49616, 16'd63057, 16'd25677, 16'd55232, 16'd2032, 16'd7417, 16'd58037, 16'd46465, 16'd14594, 16'd29557, 16'd45750, 16'd2586, 16'd47452, 16'd34592, 16'd37736, 16'd5583, 16'd43263, 16'd38012, 16'd27014, 16'd32508, 16'd2876, 16'd65012, 16'd7270, 16'd10358});
	test_expansion(128'h4add224945511b2d80c77139931b0b95, {16'd65226, 16'd59117, 16'd1002, 16'd60254, 16'd35601, 16'd27098, 16'd56199, 16'd45269, 16'd34640, 16'd18761, 16'd51539, 16'd39409, 16'd38580, 16'd52077, 16'd53799, 16'd10055, 16'd40746, 16'd58249, 16'd3413, 16'd7523, 16'd59413, 16'd38999, 16'd23251, 16'd64408, 16'd7880, 16'd21334});
	test_expansion(128'h118f0f3424cddd7c14fe6d470ced00dd, {16'd23511, 16'd11965, 16'd41241, 16'd4665, 16'd8823, 16'd52347, 16'd29965, 16'd8179, 16'd48258, 16'd41869, 16'd30082, 16'd64904, 16'd18904, 16'd17242, 16'd30639, 16'd11595, 16'd7987, 16'd30125, 16'd54683, 16'd45296, 16'd32624, 16'd1461, 16'd63215, 16'd35088, 16'd47011, 16'd65415});
	test_expansion(128'h790aef047c92d36003df3b998e41aa9c, {16'd46056, 16'd63274, 16'd42167, 16'd5968, 16'd15625, 16'd33801, 16'd37520, 16'd57438, 16'd49119, 16'd36920, 16'd41852, 16'd18548, 16'd40541, 16'd37505, 16'd25586, 16'd49036, 16'd62139, 16'd4564, 16'd31973, 16'd61160, 16'd59011, 16'd4480, 16'd9560, 16'd13346, 16'd6096, 16'd23540});
	test_expansion(128'hf1af869d9956c04f9688a094d5be84ed, {16'd62811, 16'd840, 16'd34172, 16'd10292, 16'd63375, 16'd12154, 16'd64061, 16'd52868, 16'd13962, 16'd64643, 16'd61664, 16'd38173, 16'd8302, 16'd19593, 16'd33416, 16'd12225, 16'd5000, 16'd28038, 16'd4414, 16'd37116, 16'd1225, 16'd1047, 16'd20890, 16'd37091, 16'd43547, 16'd57437});
	test_expansion(128'h6f9c5d9f3445e21c0f2ef69d26136638, {16'd10459, 16'd30149, 16'd26794, 16'd61907, 16'd23658, 16'd40268, 16'd34725, 16'd28635, 16'd63807, 16'd6756, 16'd65086, 16'd13625, 16'd52292, 16'd14929, 16'd60439, 16'd13820, 16'd21613, 16'd3766, 16'd48113, 16'd64029, 16'd940, 16'd34847, 16'd31763, 16'd61136, 16'd13809, 16'd7449});
	test_expansion(128'hb1acc9a244720cb28dd557046d05dc24, {16'd28313, 16'd29129, 16'd24531, 16'd4039, 16'd53581, 16'd8015, 16'd37595, 16'd43640, 16'd55357, 16'd36013, 16'd60518, 16'd26155, 16'd15340, 16'd59748, 16'd49785, 16'd32111, 16'd47287, 16'd27764, 16'd7956, 16'd10592, 16'd5236, 16'd47689, 16'd22985, 16'd44008, 16'd28223, 16'd29758});
	test_expansion(128'h56a7d16cb408104c06fbfcfe784be2b2, {16'd20282, 16'd24630, 16'd16494, 16'd17993, 16'd1068, 16'd58123, 16'd19982, 16'd40704, 16'd62027, 16'd64759, 16'd28630, 16'd29062, 16'd3840, 16'd63283, 16'd22051, 16'd53460, 16'd12820, 16'd60728, 16'd48993, 16'd44330, 16'd12556, 16'd32082, 16'd35730, 16'd34803, 16'd57300, 16'd38214});
	test_expansion(128'h50266e0193cfc3fd1b2cc617393f5f68, {16'd31648, 16'd41819, 16'd43879, 16'd58165, 16'd47208, 16'd51578, 16'd49638, 16'd43001, 16'd12968, 16'd3874, 16'd23750, 16'd38788, 16'd10353, 16'd28239, 16'd40786, 16'd8177, 16'd63347, 16'd58154, 16'd4674, 16'd43524, 16'd4782, 16'd28222, 16'd13601, 16'd2496, 16'd56034, 16'd59590});
	test_expansion(128'h57040d23a1aaf23536ba5bcf5727ccd6, {16'd16340, 16'd23931, 16'd35167, 16'd51455, 16'd40600, 16'd60895, 16'd11688, 16'd39879, 16'd61813, 16'd6, 16'd53120, 16'd49672, 16'd13941, 16'd1091, 16'd34406, 16'd29779, 16'd14230, 16'd8702, 16'd51827, 16'd14418, 16'd64090, 16'd4898, 16'd64139, 16'd16312, 16'd53279, 16'd47481});
	test_expansion(128'ha9325c8f60a858ec9b3241cf647a9a5a, {16'd47129, 16'd21541, 16'd3460, 16'd39412, 16'd35639, 16'd40876, 16'd27764, 16'd38291, 16'd40588, 16'd1087, 16'd8406, 16'd1928, 16'd7890, 16'd17488, 16'd61224, 16'd9143, 16'd42997, 16'd44846, 16'd5302, 16'd48366, 16'd12974, 16'd21844, 16'd7575, 16'd62645, 16'd38568, 16'd36922});
	test_expansion(128'ha8a8f1873df8404725d5e82baff3128a, {16'd26541, 16'd9480, 16'd38315, 16'd48055, 16'd59356, 16'd31438, 16'd43666, 16'd32625, 16'd45858, 16'd4817, 16'd28616, 16'd41975, 16'd19324, 16'd38566, 16'd29822, 16'd48836, 16'd38577, 16'd13069, 16'd13792, 16'd17676, 16'd8892, 16'd54367, 16'd45739, 16'd40646, 16'd49433, 16'd57734});
	test_expansion(128'hddc53aee66f22a729eab76267f286fd5, {16'd53571, 16'd62523, 16'd10466, 16'd37996, 16'd58091, 16'd4401, 16'd36536, 16'd13538, 16'd56498, 16'd19369, 16'd39035, 16'd6478, 16'd40734, 16'd35308, 16'd56476, 16'd41685, 16'd58690, 16'd20330, 16'd21115, 16'd42630, 16'd41003, 16'd11710, 16'd31304, 16'd15175, 16'd4208, 16'd8786});
	test_expansion(128'h1f2d25a2006d44f01d0c85fa272ce5ce, {16'd18683, 16'd48979, 16'd13266, 16'd25580, 16'd43637, 16'd5963, 16'd61241, 16'd12251, 16'd32723, 16'd41723, 16'd33956, 16'd47879, 16'd27865, 16'd63896, 16'd41289, 16'd31167, 16'd45096, 16'd6997, 16'd29458, 16'd222, 16'd8673, 16'd43114, 16'd15412, 16'd16838, 16'd44684, 16'd55847});
	test_expansion(128'h770fe00dd7ed7e2dfba8a4735b45db27, {16'd14780, 16'd1102, 16'd41885, 16'd42052, 16'd13309, 16'd28522, 16'd63056, 16'd33630, 16'd49624, 16'd25998, 16'd30384, 16'd44429, 16'd29079, 16'd3979, 16'd35334, 16'd5855, 16'd27995, 16'd62440, 16'd4467, 16'd39043, 16'd40511, 16'd50836, 16'd62613, 16'd4466, 16'd14762, 16'd21440});
	test_expansion(128'he92e1238bb94088998923fafa120a696, {16'd62449, 16'd19883, 16'd18405, 16'd52808, 16'd36445, 16'd16702, 16'd31361, 16'd1491, 16'd37963, 16'd55047, 16'd25057, 16'd21674, 16'd35355, 16'd39401, 16'd33004, 16'd45297, 16'd55008, 16'd16213, 16'd21198, 16'd1400, 16'd21985, 16'd30803, 16'd44285, 16'd5920, 16'd17388, 16'd19179});
	test_expansion(128'h3b189f7919274e6b11aa61e4f05dfea9, {16'd30473, 16'd49041, 16'd24203, 16'd44574, 16'd59651, 16'd41161, 16'd6673, 16'd6317, 16'd40399, 16'd9532, 16'd32878, 16'd18888, 16'd32398, 16'd5614, 16'd24519, 16'd43473, 16'd6957, 16'd608, 16'd38023, 16'd23900, 16'd50928, 16'd52996, 16'd54543, 16'd13092, 16'd15023, 16'd27408});
	test_expansion(128'hdc23e5c76375f2245f8b05432d2b2acd, {16'd1546, 16'd4146, 16'd14548, 16'd22667, 16'd26245, 16'd62418, 16'd4525, 16'd45498, 16'd20557, 16'd60046, 16'd21842, 16'd21554, 16'd30710, 16'd34782, 16'd10303, 16'd23778, 16'd13064, 16'd59142, 16'd43916, 16'd59068, 16'd6159, 16'd43743, 16'd46681, 16'd65070, 16'd41841, 16'd46230});
	test_expansion(128'ha7f4e10f070c9ea8d4977312977321ec, {16'd32898, 16'd30283, 16'd43450, 16'd14084, 16'd665, 16'd15253, 16'd22731, 16'd23411, 16'd58329, 16'd13921, 16'd20876, 16'd38091, 16'd59042, 16'd14929, 16'd28402, 16'd48519, 16'd30121, 16'd28893, 16'd31552, 16'd62804, 16'd51060, 16'd61802, 16'd34493, 16'd53377, 16'd5144, 16'd3139});
	test_expansion(128'h4cdf22cd24910aea9281891244989885, {16'd5252, 16'd16153, 16'd53328, 16'd50036, 16'd2961, 16'd63418, 16'd20819, 16'd31317, 16'd38253, 16'd52245, 16'd18594, 16'd65268, 16'd64367, 16'd5981, 16'd23107, 16'd2688, 16'd43475, 16'd24645, 16'd8476, 16'd37995, 16'd64100, 16'd47316, 16'd35798, 16'd27440, 16'd13373, 16'd861});
	test_expansion(128'h0ec6adfc96a5cbdb4c4a9a98f761f69a, {16'd60649, 16'd7009, 16'd14132, 16'd10694, 16'd52398, 16'd61263, 16'd65195, 16'd40558, 16'd17451, 16'd17709, 16'd59157, 16'd54126, 16'd11358, 16'd43903, 16'd41293, 16'd5156, 16'd56985, 16'd32198, 16'd62275, 16'd57807, 16'd48335, 16'd45962, 16'd9797, 16'd5522, 16'd9427, 16'd43107});
	test_expansion(128'h151e912fb846a865f15e81a6eca60625, {16'd20735, 16'd4262, 16'd16693, 16'd17805, 16'd4257, 16'd21823, 16'd4592, 16'd50722, 16'd52009, 16'd38925, 16'd24611, 16'd19606, 16'd4436, 16'd42052, 16'd18672, 16'd51577, 16'd64132, 16'd14092, 16'd11417, 16'd43149, 16'd7588, 16'd36366, 16'd47344, 16'd31883, 16'd4831, 16'd59831});
	test_expansion(128'he4f30442f4ad1ba04354402dd5a7f8fd, {16'd41944, 16'd1071, 16'd49476, 16'd1196, 16'd4936, 16'd99, 16'd14710, 16'd49136, 16'd24277, 16'd61040, 16'd28784, 16'd39569, 16'd16696, 16'd19755, 16'd17231, 16'd16044, 16'd39576, 16'd28134, 16'd19589, 16'd11074, 16'd21554, 16'd62940, 16'd7087, 16'd19538, 16'd3036, 16'd36939});
	test_expansion(128'hea38c72f42a5cac5b6b46d64def2e53f, {16'd10709, 16'd30879, 16'd37468, 16'd27234, 16'd52471, 16'd34991, 16'd20962, 16'd33303, 16'd62393, 16'd43136, 16'd19764, 16'd46829, 16'd59934, 16'd30052, 16'd15008, 16'd52688, 16'd14085, 16'd38425, 16'd44263, 16'd64331, 16'd28880, 16'd52903, 16'd13654, 16'd58319, 16'd57612, 16'd18136});
	test_expansion(128'h2db6e580f293b77b2263ceabfb8009df, {16'd58296, 16'd12004, 16'd18931, 16'd34364, 16'd8205, 16'd5195, 16'd31357, 16'd39057, 16'd46100, 16'd48732, 16'd60557, 16'd34883, 16'd24683, 16'd43711, 16'd63501, 16'd48269, 16'd11262, 16'd31853, 16'd15446, 16'd20593, 16'd15876, 16'd65125, 16'd29185, 16'd41878, 16'd3480, 16'd11586});
	test_expansion(128'h89fc30763fdfdd7d2832677e66707b00, {16'd26523, 16'd6356, 16'd43596, 16'd14694, 16'd19176, 16'd2716, 16'd32944, 16'd33358, 16'd33201, 16'd51817, 16'd8464, 16'd63759, 16'd7418, 16'd7821, 16'd9605, 16'd7784, 16'd29319, 16'd31976, 16'd52510, 16'd19557, 16'd3754, 16'd10774, 16'd6329, 16'd57689, 16'd15215, 16'd50265});
	test_expansion(128'h78f9ba43fcbe379a3b00887c959d2182, {16'd27390, 16'd56335, 16'd18318, 16'd47933, 16'd4671, 16'd17049, 16'd45218, 16'd23715, 16'd20678, 16'd59559, 16'd36967, 16'd59390, 16'd15773, 16'd12604, 16'd14114, 16'd38198, 16'd17949, 16'd32447, 16'd45107, 16'd18461, 16'd50130, 16'd25376, 16'd38312, 16'd41146, 16'd15904, 16'd54421});
	test_expansion(128'heea72b4ddbcba389c8ba5f5291204784, {16'd21415, 16'd18250, 16'd62443, 16'd19183, 16'd40316, 16'd45538, 16'd42918, 16'd44084, 16'd22683, 16'd53281, 16'd30555, 16'd42817, 16'd10076, 16'd24245, 16'd36650, 16'd63629, 16'd64659, 16'd33356, 16'd56384, 16'd46851, 16'd21534, 16'd11648, 16'd64395, 16'd35474, 16'd15372, 16'd61524});
	test_expansion(128'h67c2aba67c6dd5d18c1e832d198f649e, {16'd5830, 16'd55407, 16'd47311, 16'd9370, 16'd12092, 16'd39818, 16'd22899, 16'd57529, 16'd29192, 16'd22957, 16'd53441, 16'd62847, 16'd9272, 16'd33412, 16'd62275, 16'd1839, 16'd60397, 16'd15789, 16'd24361, 16'd31784, 16'd2580, 16'd64274, 16'd39323, 16'd32632, 16'd28042, 16'd14234});
	test_expansion(128'h6da8da086d487bfbdb390af8295aebf4, {16'd1397, 16'd25042, 16'd61739, 16'd3039, 16'd35061, 16'd6062, 16'd59828, 16'd29015, 16'd37828, 16'd23249, 16'd33093, 16'd34014, 16'd53074, 16'd28204, 16'd14294, 16'd51643, 16'd40450, 16'd57650, 16'd4041, 16'd59831, 16'd20422, 16'd65377, 16'd60055, 16'd39424, 16'd64222, 16'd65452});
	test_expansion(128'h5b93285274dc4e40cf2f3b456409271b, {16'd42305, 16'd817, 16'd38428, 16'd26569, 16'd4153, 16'd31147, 16'd36855, 16'd24770, 16'd58749, 16'd46617, 16'd25580, 16'd46827, 16'd12532, 16'd4301, 16'd27004, 16'd29846, 16'd56336, 16'd25020, 16'd43249, 16'd27251, 16'd39398, 16'd63745, 16'd64834, 16'd38264, 16'd48371, 16'd2187});
	test_expansion(128'hef50fefb9190ebccd46f6345f8ff9b3e, {16'd64392, 16'd5331, 16'd57756, 16'd26275, 16'd9281, 16'd43868, 16'd38046, 16'd55385, 16'd13527, 16'd44567, 16'd566, 16'd19808, 16'd40438, 16'd57998, 16'd19096, 16'd43195, 16'd29828, 16'd26066, 16'd48620, 16'd10523, 16'd52631, 16'd63826, 16'd27268, 16'd62861, 16'd1214, 16'd54850});
	test_expansion(128'h4c219337fa80b1e1cc4975734f87dc19, {16'd18237, 16'd9695, 16'd24489, 16'd50605, 16'd8772, 16'd65072, 16'd54612, 16'd28004, 16'd29752, 16'd34581, 16'd55781, 16'd14917, 16'd42444, 16'd13106, 16'd36814, 16'd40878, 16'd43152, 16'd64797, 16'd45236, 16'd849, 16'd15730, 16'd64062, 16'd15706, 16'd9178, 16'd4441, 16'd56511});
	test_expansion(128'hb99f39d5f31cfac45dcf6d8c9967ee45, {16'd53932, 16'd43914, 16'd37766, 16'd37545, 16'd1069, 16'd38618, 16'd29765, 16'd5981, 16'd8546, 16'd61962, 16'd49289, 16'd23382, 16'd5210, 16'd30043, 16'd46387, 16'd46652, 16'd26085, 16'd63230, 16'd836, 16'd16214, 16'd4928, 16'd49092, 16'd26434, 16'd17369, 16'd41018, 16'd39165});
	test_expansion(128'h07b74af81ece445f9c6c82c9d2d61c6e, {16'd62345, 16'd37510, 16'd21874, 16'd43944, 16'd37326, 16'd49643, 16'd2458, 16'd48780, 16'd15800, 16'd30045, 16'd13257, 16'd37887, 16'd1105, 16'd63622, 16'd12184, 16'd58082, 16'd46646, 16'd18037, 16'd47818, 16'd5142, 16'd16593, 16'd61646, 16'd33934, 16'd8102, 16'd50514, 16'd65167});
	test_expansion(128'h486c5432f3a744f382cad9e700669da7, {16'd30764, 16'd23264, 16'd16495, 16'd12358, 16'd42126, 16'd36886, 16'd11425, 16'd10807, 16'd31983, 16'd34075, 16'd8010, 16'd26185, 16'd39204, 16'd35678, 16'd23886, 16'd20059, 16'd31545, 16'd37859, 16'd50228, 16'd5827, 16'd41545, 16'd13663, 16'd61728, 16'd43709, 16'd47364, 16'd57343});
	test_expansion(128'hedded1c2b3173c03111e61efd3dd7824, {16'd47236, 16'd57205, 16'd64997, 16'd35334, 16'd29930, 16'd13491, 16'd30745, 16'd6283, 16'd4987, 16'd41482, 16'd51562, 16'd48752, 16'd10336, 16'd2274, 16'd20352, 16'd5110, 16'd52986, 16'd57574, 16'd2781, 16'd40406, 16'd60646, 16'd54438, 16'd51719, 16'd6289, 16'd10743, 16'd12249});
	test_expansion(128'h0d8c3029e19cc0880ef3219a0b671eac, {16'd8794, 16'd1139, 16'd4422, 16'd45924, 16'd26749, 16'd26901, 16'd33711, 16'd9178, 16'd55419, 16'd44990, 16'd13028, 16'd40575, 16'd47313, 16'd22565, 16'd22634, 16'd18102, 16'd26966, 16'd57066, 16'd33123, 16'd39044, 16'd63632, 16'd53708, 16'd58046, 16'd11764, 16'd60771, 16'd60726});
	test_expansion(128'hd88c386d95c47d5e421c14ff2a494181, {16'd9475, 16'd62635, 16'd64629, 16'd462, 16'd18303, 16'd24383, 16'd19321, 16'd14401, 16'd55155, 16'd13999, 16'd51834, 16'd55111, 16'd5462, 16'd35142, 16'd4255, 16'd41654, 16'd60807, 16'd37839, 16'd31996, 16'd8107, 16'd31990, 16'd1383, 16'd27220, 16'd3941, 16'd57619, 16'd57562});
	test_expansion(128'h23754b70393894befdd4728fd94dd032, {16'd2838, 16'd52129, 16'd4676, 16'd6938, 16'd1050, 16'd26468, 16'd23330, 16'd7448, 16'd6773, 16'd1852, 16'd52701, 16'd2976, 16'd13421, 16'd9372, 16'd14240, 16'd49961, 16'd30834, 16'd4017, 16'd55580, 16'd2067, 16'd42979, 16'd47724, 16'd50315, 16'd40387, 16'd52516, 16'd57009});
	test_expansion(128'heda1ca84d6904a4523abae2c16c8ec4a, {16'd30329, 16'd53200, 16'd36739, 16'd37459, 16'd41782, 16'd62779, 16'd35790, 16'd41267, 16'd2274, 16'd27800, 16'd13127, 16'd18984, 16'd22948, 16'd38988, 16'd37719, 16'd8605, 16'd2662, 16'd14354, 16'd8352, 16'd35375, 16'd57969, 16'd40502, 16'd27014, 16'd33335, 16'd48025, 16'd51942});
	test_expansion(128'ha8938b299fde93aa9c6dac42447f36e4, {16'd11175, 16'd44113, 16'd28849, 16'd39965, 16'd44974, 16'd47056, 16'd43040, 16'd1184, 16'd45305, 16'd57990, 16'd7515, 16'd34331, 16'd33311, 16'd55483, 16'd58432, 16'd51987, 16'd57391, 16'd46850, 16'd62699, 16'd23119, 16'd1210, 16'd45952, 16'd36269, 16'd53983, 16'd19089, 16'd50901});
	test_expansion(128'h111107a719578d859bd81b0e4dbd44b6, {16'd12396, 16'd11813, 16'd36853, 16'd17447, 16'd51448, 16'd52660, 16'd64537, 16'd9886, 16'd40836, 16'd31683, 16'd44135, 16'd3442, 16'd35139, 16'd51129, 16'd10686, 16'd49866, 16'd20851, 16'd9386, 16'd16833, 16'd32551, 16'd47915, 16'd9530, 16'd56247, 16'd61590, 16'd16561, 16'd46913});
	test_expansion(128'h8897a7aea07b2d5fa1d088feea796d13, {16'd52057, 16'd18387, 16'd46802, 16'd33238, 16'd21273, 16'd15023, 16'd57843, 16'd41756, 16'd8736, 16'd8508, 16'd19339, 16'd13928, 16'd18145, 16'd7247, 16'd57480, 16'd60533, 16'd43628, 16'd6053, 16'd23641, 16'd62654, 16'd3409, 16'd20270, 16'd21640, 16'd57475, 16'd11453, 16'd48099});
	test_expansion(128'hb037cbfe10cd9bae625869e4d70ef18e, {16'd51572, 16'd34413, 16'd3050, 16'd62410, 16'd47666, 16'd54606, 16'd60435, 16'd47409, 16'd898, 16'd49154, 16'd47539, 16'd567, 16'd59467, 16'd58294, 16'd29066, 16'd34114, 16'd14247, 16'd58959, 16'd58345, 16'd1416, 16'd36671, 16'd36104, 16'd48032, 16'd49781, 16'd59690, 16'd22723});
	test_expansion(128'h32a3085cefd81499fea9d7e2cfd83f00, {16'd63894, 16'd19557, 16'd21963, 16'd55457, 16'd43528, 16'd34707, 16'd38561, 16'd33942, 16'd34312, 16'd31108, 16'd18341, 16'd23813, 16'd13038, 16'd36206, 16'd36291, 16'd8138, 16'd13952, 16'd57158, 16'd63373, 16'd8379, 16'd3410, 16'd15943, 16'd26088, 16'd52648, 16'd4919, 16'd23404});
	test_expansion(128'hcceba836e04e660362cd2822336318b9, {16'd24116, 16'd37999, 16'd8208, 16'd59514, 16'd3723, 16'd39490, 16'd31206, 16'd37854, 16'd32029, 16'd37070, 16'd63375, 16'd57811, 16'd41312, 16'd52246, 16'd19040, 16'd25454, 16'd41357, 16'd52383, 16'd973, 16'd51542, 16'd25072, 16'd13557, 16'd63632, 16'd2542, 16'd7057, 16'd23890});
	test_expansion(128'h20a37f1c2edec273370fa4c2c42ec602, {16'd11294, 16'd34677, 16'd37772, 16'd43908, 16'd21585, 16'd60959, 16'd22910, 16'd43394, 16'd29334, 16'd60207, 16'd65465, 16'd64759, 16'd37435, 16'd54299, 16'd1504, 16'd25116, 16'd65500, 16'd65182, 16'd35075, 16'd31048, 16'd60158, 16'd7178, 16'd47814, 16'd31262, 16'd43034, 16'd39736});
	test_expansion(128'h279764624e8e6e1fa4476f28cb1923dd, {16'd53366, 16'd10902, 16'd55405, 16'd33470, 16'd31049, 16'd8824, 16'd34440, 16'd60949, 16'd53907, 16'd12347, 16'd9259, 16'd6273, 16'd19840, 16'd30428, 16'd19067, 16'd60808, 16'd39007, 16'd54830, 16'd14859, 16'd26568, 16'd63426, 16'd30944, 16'd46304, 16'd37911, 16'd29629, 16'd63353});
	test_expansion(128'h472a16cbd9efcb8a2aafa0a372631b98, {16'd62802, 16'd15170, 16'd2763, 16'd34461, 16'd7948, 16'd40025, 16'd55966, 16'd51482, 16'd63299, 16'd47549, 16'd64130, 16'd61493, 16'd51235, 16'd12842, 16'd56332, 16'd1684, 16'd32375, 16'd136, 16'd59352, 16'd7278, 16'd39883, 16'd14971, 16'd42672, 16'd26114, 16'd63959, 16'd24151});
	test_expansion(128'h0300e2f268907b4d80a823a7ccf1518e, {16'd56818, 16'd28670, 16'd35936, 16'd12687, 16'd43856, 16'd26025, 16'd14246, 16'd34863, 16'd50561, 16'd48855, 16'd8442, 16'd20095, 16'd24269, 16'd25601, 16'd21345, 16'd12480, 16'd47816, 16'd54602, 16'd56311, 16'd45932, 16'd16721, 16'd26205, 16'd36427, 16'd51930, 16'd26342, 16'd993});
	test_expansion(128'h69283b5d9f3d2ba2f10474a86b4f9153, {16'd24325, 16'd30723, 16'd31250, 16'd14735, 16'd1124, 16'd46408, 16'd46593, 16'd51186, 16'd30951, 16'd3839, 16'd7867, 16'd34161, 16'd28583, 16'd39748, 16'd64490, 16'd30297, 16'd1224, 16'd13070, 16'd29062, 16'd38819, 16'd51558, 16'd48516, 16'd33702, 16'd16678, 16'd47784, 16'd2758});
	test_expansion(128'h7adbe3b6cd59a734c6f7798cfe0bf728, {16'd50419, 16'd15294, 16'd48004, 16'd47501, 16'd33181, 16'd34643, 16'd5501, 16'd51410, 16'd50221, 16'd28775, 16'd45759, 16'd32985, 16'd59963, 16'd988, 16'd55206, 16'd19728, 16'd57283, 16'd56986, 16'd41937, 16'd25203, 16'd4743, 16'd17384, 16'd2826, 16'd51004, 16'd34329, 16'd22359});
	test_expansion(128'hf4e7716cc2544d3d486dad474753e660, {16'd21555, 16'd46018, 16'd40072, 16'd33035, 16'd3764, 16'd30610, 16'd27336, 16'd39196, 16'd51569, 16'd45831, 16'd42488, 16'd20463, 16'd24392, 16'd15333, 16'd34536, 16'd38977, 16'd57312, 16'd177, 16'd55868, 16'd35245, 16'd15105, 16'd29401, 16'd16358, 16'd43234, 16'd64482, 16'd58141});
	test_expansion(128'h10581d30abdf9750e7becf588439c30f, {16'd5237, 16'd31106, 16'd52003, 16'd26063, 16'd41232, 16'd19892, 16'd44567, 16'd14804, 16'd57842, 16'd33971, 16'd64687, 16'd33931, 16'd25501, 16'd16573, 16'd45606, 16'd63611, 16'd30841, 16'd28860, 16'd31986, 16'd35199, 16'd60503, 16'd3421, 16'd62399, 16'd39783, 16'd47012, 16'd47562});
	test_expansion(128'hc42051bc1446a77e2645b98cedc6a517, {16'd49563, 16'd33897, 16'd19500, 16'd38537, 16'd12138, 16'd4190, 16'd54234, 16'd8716, 16'd28785, 16'd8597, 16'd28490, 16'd48299, 16'd15227, 16'd8851, 16'd27398, 16'd43602, 16'd55303, 16'd63646, 16'd49239, 16'd8004, 16'd4254, 16'd31017, 16'd44865, 16'd16215, 16'd31571, 16'd39229});
	test_expansion(128'hf4f4afa15224c878b865bd74e230c1ed, {16'd10029, 16'd20343, 16'd3746, 16'd65033, 16'd48287, 16'd34179, 16'd63065, 16'd25601, 16'd47065, 16'd60090, 16'd19764, 16'd20494, 16'd56536, 16'd4633, 16'd35849, 16'd47215, 16'd13604, 16'd23171, 16'd41162, 16'd962, 16'd61287, 16'd60382, 16'd65374, 16'd11716, 16'd56289, 16'd5517});
	test_expansion(128'h13fdbb564dd638df13b7f57965722cca, {16'd59711, 16'd7607, 16'd57128, 16'd29291, 16'd59346, 16'd16780, 16'd63025, 16'd3897, 16'd9673, 16'd9259, 16'd25297, 16'd32516, 16'd56390, 16'd6631, 16'd60195, 16'd63995, 16'd44063, 16'd9715, 16'd52272, 16'd34558, 16'd26842, 16'd45209, 16'd18509, 16'd871, 16'd23271, 16'd27259});
	test_expansion(128'hfe95d322738aae08870073c9d9eb6f2d, {16'd391, 16'd61130, 16'd43609, 16'd47008, 16'd52937, 16'd20503, 16'd25973, 16'd38568, 16'd48519, 16'd2514, 16'd37990, 16'd43227, 16'd64160, 16'd5281, 16'd35553, 16'd42091, 16'd62318, 16'd40134, 16'd10557, 16'd12502, 16'd54151, 16'd643, 16'd31623, 16'd25702, 16'd63154, 16'd31123});
	test_expansion(128'hfb8cf505eeaf4b3f7379b236e438d728, {16'd5034, 16'd65017, 16'd37142, 16'd55344, 16'd24300, 16'd51942, 16'd13897, 16'd31551, 16'd47883, 16'd46237, 16'd17109, 16'd43288, 16'd55812, 16'd9443, 16'd36114, 16'd55188, 16'd59991, 16'd21722, 16'd26375, 16'd64229, 16'd12982, 16'd30560, 16'd36569, 16'd55417, 16'd35820, 16'd21800});
	test_expansion(128'h8a8ae9d2bac4e6aa660b4dbfa01cdf88, {16'd54745, 16'd14946, 16'd52345, 16'd31118, 16'd26702, 16'd4246, 16'd6542, 16'd61805, 16'd37481, 16'd62409, 16'd1800, 16'd37469, 16'd8073, 16'd2819, 16'd22680, 16'd15304, 16'd45125, 16'd37188, 16'd46435, 16'd31618, 16'd48133, 16'd45323, 16'd14592, 16'd5860, 16'd169, 16'd62634});
	test_expansion(128'h928696b6d505cd74a84b354f3d35bf17, {16'd6003, 16'd8259, 16'd55191, 16'd62707, 16'd11731, 16'd56172, 16'd58670, 16'd40285, 16'd41124, 16'd4435, 16'd58675, 16'd1558, 16'd9246, 16'd38464, 16'd26392, 16'd23695, 16'd44570, 16'd9174, 16'd39320, 16'd6108, 16'd15248, 16'd63007, 16'd27031, 16'd58684, 16'd12418, 16'd33562});
	test_expansion(128'hbe13e61cb7fb539a0c71c278321c76d0, {16'd53343, 16'd11329, 16'd54948, 16'd61966, 16'd29819, 16'd59792, 16'd47270, 16'd6394, 16'd6574, 16'd52939, 16'd31621, 16'd29308, 16'd58722, 16'd19795, 16'd60901, 16'd58891, 16'd59224, 16'd55472, 16'd20268, 16'd16761, 16'd45787, 16'd13965, 16'd16734, 16'd61838, 16'd6118, 16'd20710});
	test_expansion(128'hd9947e6480a6eb7ece2be1907d3ed307, {16'd40058, 16'd23877, 16'd21915, 16'd59452, 16'd16556, 16'd57852, 16'd47060, 16'd57503, 16'd23522, 16'd29142, 16'd21987, 16'd11347, 16'd45501, 16'd17339, 16'd8055, 16'd1992, 16'd28736, 16'd3339, 16'd17153, 16'd45965, 16'd62116, 16'd57981, 16'd38919, 16'd65288, 16'd14135, 16'd56875});
	test_expansion(128'h01eff10a73cb5b6806ae73fc31d4729a, {16'd50597, 16'd30805, 16'd49632, 16'd50136, 16'd62793, 16'd10839, 16'd35605, 16'd39720, 16'd56753, 16'd15479, 16'd60170, 16'd29247, 16'd48955, 16'd31329, 16'd51790, 16'd62481, 16'd52036, 16'd42684, 16'd45354, 16'd41353, 16'd12080, 16'd12601, 16'd50035, 16'd23568, 16'd20173, 16'd2162});
	test_expansion(128'h72a409da3d7528933468d2e307a81343, {16'd30095, 16'd38088, 16'd63049, 16'd3806, 16'd11716, 16'd17815, 16'd30565, 16'd21605, 16'd36061, 16'd47707, 16'd42624, 16'd55012, 16'd55597, 16'd18478, 16'd59927, 16'd26059, 16'd15006, 16'd28772, 16'd53451, 16'd44259, 16'd21658, 16'd47614, 16'd33889, 16'd45438, 16'd47915, 16'd41580});
	test_expansion(128'hd64477b6fcf515ad9033defcc85b02ff, {16'd60513, 16'd47252, 16'd40710, 16'd10337, 16'd9116, 16'd4459, 16'd42720, 16'd43028, 16'd64389, 16'd54721, 16'd18011, 16'd15983, 16'd53622, 16'd51878, 16'd4506, 16'd48581, 16'd10927, 16'd32250, 16'd9006, 16'd23652, 16'd30657, 16'd23217, 16'd11375, 16'd53307, 16'd31717, 16'd5835});
	test_expansion(128'hec32464a0bf61fbf949721d2aa2326fc, {16'd42522, 16'd32541, 16'd16583, 16'd4074, 16'd44128, 16'd47389, 16'd55482, 16'd3133, 16'd27819, 16'd41229, 16'd6729, 16'd62107, 16'd8751, 16'd58483, 16'd46007, 16'd1137, 16'd15265, 16'd37929, 16'd62702, 16'd8941, 16'd65213, 16'd57370, 16'd39554, 16'd50252, 16'd29617, 16'd37631});
	test_expansion(128'h75de0fa6a73ca2374c888322408f9912, {16'd3731, 16'd26895, 16'd27886, 16'd53659, 16'd60965, 16'd2747, 16'd32322, 16'd36831, 16'd31484, 16'd52138, 16'd59351, 16'd34942, 16'd11241, 16'd22072, 16'd33159, 16'd2025, 16'd49121, 16'd3959, 16'd11628, 16'd12220, 16'd19680, 16'd4357, 16'd44176, 16'd48350, 16'd58726, 16'd3071});
	test_expansion(128'h8bb5c6958d0e8d3bc33a1ad98810ebad, {16'd7337, 16'd3944, 16'd49044, 16'd26188, 16'd20028, 16'd42986, 16'd23677, 16'd54558, 16'd26192, 16'd57552, 16'd26075, 16'd6007, 16'd62335, 16'd12095, 16'd59915, 16'd64588, 16'd52669, 16'd41485, 16'd42956, 16'd52969, 16'd647, 16'd47970, 16'd52690, 16'd609, 16'd63170, 16'd40032});
	test_expansion(128'h9211d53547d057e4e078ce706d8195fd, {16'd15120, 16'd53800, 16'd46854, 16'd58613, 16'd48711, 16'd8869, 16'd33473, 16'd43490, 16'd58682, 16'd10041, 16'd15973, 16'd27137, 16'd63429, 16'd46067, 16'd53487, 16'd60430, 16'd39322, 16'd36758, 16'd17290, 16'd55778, 16'd55540, 16'd37755, 16'd35850, 16'd60841, 16'd28559, 16'd53406});
	test_expansion(128'h85339802c9b5b3cc91d8707171915a23, {16'd58220, 16'd5030, 16'd30785, 16'd15546, 16'd39998, 16'd19549, 16'd48098, 16'd29717, 16'd13326, 16'd29677, 16'd18429, 16'd39938, 16'd49756, 16'd27276, 16'd38207, 16'd40946, 16'd32924, 16'd56110, 16'd40855, 16'd44959, 16'd29739, 16'd3935, 16'd34845, 16'd27818, 16'd44361, 16'd29268});
	test_expansion(128'h40dc2ddf9f8f41b93ffe761bd930f220, {16'd60703, 16'd49530, 16'd13038, 16'd8461, 16'd44233, 16'd63255, 16'd30107, 16'd46823, 16'd36348, 16'd28537, 16'd42870, 16'd25792, 16'd12363, 16'd23303, 16'd25942, 16'd10110, 16'd16733, 16'd63469, 16'd20891, 16'd52178, 16'd61010, 16'd34972, 16'd57761, 16'd24494, 16'd62915, 16'd58337});
	test_expansion(128'hd9617436bb115fc24b86f7040dcb58a4, {16'd47806, 16'd62021, 16'd32302, 16'd18162, 16'd26940, 16'd43980, 16'd33305, 16'd14792, 16'd60364, 16'd36044, 16'd16852, 16'd47652, 16'd55760, 16'd50208, 16'd28589, 16'd58411, 16'd40630, 16'd27522, 16'd22011, 16'd23081, 16'd52370, 16'd37383, 16'd40138, 16'd29881, 16'd21211, 16'd17228});
	test_expansion(128'h411cdfaa02c4340d2e76efda727fed2c, {16'd45830, 16'd40785, 16'd6971, 16'd4021, 16'd16424, 16'd2276, 16'd22008, 16'd42461, 16'd20686, 16'd65133, 16'd54051, 16'd43306, 16'd61715, 16'd64400, 16'd35307, 16'd18540, 16'd41207, 16'd11063, 16'd32128, 16'd27808, 16'd17036, 16'd30806, 16'd40864, 16'd35592, 16'd4965, 16'd17996});
	test_expansion(128'hed98fcd39dfedd2c07178a48d7670255, {16'd26473, 16'd55796, 16'd7370, 16'd15337, 16'd41519, 16'd50495, 16'd63750, 16'd21901, 16'd63630, 16'd51642, 16'd64269, 16'd58581, 16'd48639, 16'd63920, 16'd39464, 16'd54507, 16'd27548, 16'd53034, 16'd47232, 16'd22087, 16'd7176, 16'd5311, 16'd2839, 16'd3390, 16'd12508, 16'd53529});
	test_expansion(128'h9a839f8e03b4f26350ac68db12b00076, {16'd46389, 16'd24996, 16'd47045, 16'd15707, 16'd18638, 16'd27837, 16'd60416, 16'd2859, 16'd50766, 16'd10656, 16'd15428, 16'd60437, 16'd24608, 16'd24136, 16'd52601, 16'd24410, 16'd32097, 16'd20253, 16'd47025, 16'd39209, 16'd3623, 16'd18657, 16'd1326, 16'd783, 16'd2622, 16'd12658});
	test_expansion(128'hb1405a9de64f4bed19c6f78967ac2d67, {16'd51538, 16'd51623, 16'd8162, 16'd32278, 16'd4176, 16'd33141, 16'd15656, 16'd12624, 16'd2126, 16'd18618, 16'd54725, 16'd16207, 16'd20547, 16'd41712, 16'd30549, 16'd47730, 16'd7192, 16'd59886, 16'd21533, 16'd62931, 16'd6063, 16'd2929, 16'd27057, 16'd12133, 16'd59483, 16'd40116});
	test_expansion(128'h66f3c970b85a6a7be635a443aec3797b, {16'd50538, 16'd32752, 16'd374, 16'd40917, 16'd49313, 16'd2820, 16'd7925, 16'd27967, 16'd57547, 16'd58884, 16'd29521, 16'd7744, 16'd44327, 16'd52206, 16'd16286, 16'd30458, 16'd14032, 16'd62325, 16'd51207, 16'd44750, 16'd41570, 16'd5263, 16'd40559, 16'd56007, 16'd29739, 16'd50156});
	test_expansion(128'h6717f92c3b2629ea39cd0e444b7450bc, {16'd12672, 16'd42192, 16'd56359, 16'd18491, 16'd56748, 16'd21497, 16'd13125, 16'd23549, 16'd3088, 16'd39225, 16'd47613, 16'd14094, 16'd34904, 16'd40325, 16'd44077, 16'd27069, 16'd35364, 16'd57454, 16'd22887, 16'd18349, 16'd48596, 16'd26125, 16'd21148, 16'd19167, 16'd25, 16'd5037});
	test_expansion(128'hddecf07348546c9b6cc2ed0ff2e9da35, {16'd15277, 16'd33374, 16'd45066, 16'd47631, 16'd40593, 16'd22724, 16'd39350, 16'd28330, 16'd63929, 16'd513, 16'd5089, 16'd34463, 16'd42657, 16'd6567, 16'd48117, 16'd22124, 16'd9018, 16'd60855, 16'd10089, 16'd48735, 16'd8750, 16'd3758, 16'd34712, 16'd38720, 16'd61153, 16'd61271});
	test_expansion(128'h6368b526248d7f14727198ca00b53c0b, {16'd14741, 16'd33708, 16'd61366, 16'd34279, 16'd44284, 16'd11472, 16'd36583, 16'd48176, 16'd14637, 16'd5681, 16'd51988, 16'd1829, 16'd59668, 16'd33899, 16'd53320, 16'd10216, 16'd6198, 16'd64508, 16'd35223, 16'd33870, 16'd34773, 16'd36101, 16'd36019, 16'd45652, 16'd40536, 16'd43391});
	test_expansion(128'he4b3cd72b63b449c7c1b3bcc2d5d63ae, {16'd38794, 16'd60412, 16'd41171, 16'd31029, 16'd34646, 16'd48920, 16'd33323, 16'd34254, 16'd42440, 16'd28367, 16'd53993, 16'd20895, 16'd48475, 16'd50713, 16'd34017, 16'd1959, 16'd58127, 16'd37535, 16'd9886, 16'd37122, 16'd47977, 16'd21077, 16'd46871, 16'd51784, 16'd21443, 16'd2337});
	test_expansion(128'h3b22009a64e2361140d6c8c4765d0348, {16'd51222, 16'd33463, 16'd23899, 16'd39583, 16'd15491, 16'd4889, 16'd15330, 16'd49184, 16'd51415, 16'd40705, 16'd41835, 16'd13149, 16'd54338, 16'd35173, 16'd59946, 16'd21010, 16'd63421, 16'd35798, 16'd44187, 16'd49914, 16'd60935, 16'd60935, 16'd16593, 16'd47648, 16'd4987, 16'd42854});
	test_expansion(128'haa91abe7220c61ea3b81be9c5f9f2d4b, {16'd32168, 16'd48901, 16'd50868, 16'd32045, 16'd39449, 16'd20492, 16'd17157, 16'd2777, 16'd22299, 16'd8849, 16'd54063, 16'd5082, 16'd42036, 16'd1612, 16'd758, 16'd58789, 16'd40887, 16'd31742, 16'd48196, 16'd21076, 16'd36287, 16'd61170, 16'd7617, 16'd21226, 16'd6993, 16'd6169});
	test_expansion(128'hd6d2a0750f62e0e531654d0f46f836e6, {16'd6453, 16'd42304, 16'd52478, 16'd63776, 16'd20587, 16'd31440, 16'd64672, 16'd39851, 16'd43926, 16'd13817, 16'd59584, 16'd41874, 16'd19074, 16'd29069, 16'd17132, 16'd24408, 16'd29336, 16'd32585, 16'd41604, 16'd63129, 16'd31953, 16'd50437, 16'd51051, 16'd25506, 16'd56577, 16'd41556});
	test_expansion(128'h8b54af4a1e4f377401183390345df77a, {16'd43786, 16'd31047, 16'd33252, 16'd55513, 16'd59293, 16'd18567, 16'd41243, 16'd45244, 16'd25841, 16'd26803, 16'd3457, 16'd58670, 16'd26566, 16'd9964, 16'd31426, 16'd35656, 16'd27311, 16'd39877, 16'd41252, 16'd6174, 16'd27708, 16'd6833, 16'd9393, 16'd47913, 16'd14022, 16'd6164});
	test_expansion(128'h795367cb5f324cb249c7926a846d2769, {16'd65438, 16'd12521, 16'd54522, 16'd47757, 16'd52778, 16'd19130, 16'd31307, 16'd35404, 16'd34398, 16'd51825, 16'd45594, 16'd33389, 16'd876, 16'd6902, 16'd56430, 16'd224, 16'd28593, 16'd25478, 16'd47118, 16'd50229, 16'd32989, 16'd19669, 16'd21644, 16'd51949, 16'd13715, 16'd13633});
	test_expansion(128'h23b69ebb33fcc755ee7ffb697818d862, {16'd3461, 16'd40255, 16'd28759, 16'd58174, 16'd1278, 16'd8777, 16'd59080, 16'd24498, 16'd41013, 16'd61078, 16'd7305, 16'd21737, 16'd7560, 16'd11248, 16'd4538, 16'd50780, 16'd34955, 16'd40278, 16'd11740, 16'd18054, 16'd57926, 16'd28411, 16'd21239, 16'd1872, 16'd42610, 16'd36667});
	test_expansion(128'h8fd74b7a6b439c4a91f0e11a0e284f75, {16'd60512, 16'd57771, 16'd27797, 16'd15556, 16'd9084, 16'd25664, 16'd3122, 16'd39621, 16'd52438, 16'd30384, 16'd35142, 16'd21607, 16'd20368, 16'd8405, 16'd61859, 16'd45347, 16'd57890, 16'd19185, 16'd33667, 16'd705, 16'd4199, 16'd40628, 16'd881, 16'd47062, 16'd29286, 16'd60822});
	test_expansion(128'h2f248a50d81043657664802cbba7274a, {16'd51688, 16'd3600, 16'd30352, 16'd36113, 16'd18985, 16'd9987, 16'd14872, 16'd40149, 16'd31947, 16'd15127, 16'd65204, 16'd57597, 16'd4827, 16'd21100, 16'd12347, 16'd3730, 16'd56769, 16'd38943, 16'd58759, 16'd5115, 16'd25075, 16'd41308, 16'd51620, 16'd30457, 16'd54087, 16'd25464});
	test_expansion(128'h7ba1fc98ad12c9c958253bfdf5da059b, {16'd32219, 16'd10604, 16'd8216, 16'd12693, 16'd36696, 16'd47721, 16'd55610, 16'd32309, 16'd42352, 16'd34121, 16'd27400, 16'd17360, 16'd64151, 16'd31787, 16'd3316, 16'd11062, 16'd52063, 16'd42884, 16'd61788, 16'd16608, 16'd12323, 16'd52038, 16'd38501, 16'd50731, 16'd28385, 16'd1707});
	test_expansion(128'hf7ab347e5ae15386446f1b62e7be0a8f, {16'd1077, 16'd31792, 16'd52655, 16'd13034, 16'd45326, 16'd51626, 16'd24960, 16'd44965, 16'd52035, 16'd50421, 16'd25119, 16'd51767, 16'd28862, 16'd997, 16'd25905, 16'd45253, 16'd30489, 16'd58882, 16'd60841, 16'd48336, 16'd63793, 16'd32070, 16'd12922, 16'd41751, 16'd59947, 16'd49236});
	test_expansion(128'hc9dfa03b04cced7932815f05cbc40114, {16'd32631, 16'd64169, 16'd33816, 16'd55130, 16'd44006, 16'd53139, 16'd54855, 16'd20103, 16'd3875, 16'd30941, 16'd6921, 16'd35204, 16'd33734, 16'd842, 16'd12475, 16'd17116, 16'd51267, 16'd42002, 16'd29436, 16'd14745, 16'd18649, 16'd55207, 16'd36115, 16'd24353, 16'd35081, 16'd6068});
	test_expansion(128'h3a404e02d4a1e7ed1e7abe624e1230d7, {16'd10479, 16'd16814, 16'd1988, 16'd35525, 16'd60443, 16'd11686, 16'd51428, 16'd55852, 16'd44558, 16'd56480, 16'd46659, 16'd52095, 16'd18848, 16'd59455, 16'd54344, 16'd684, 16'd11440, 16'd63266, 16'd62702, 16'd25501, 16'd28364, 16'd63042, 16'd63474, 16'd61206, 16'd25598, 16'd37146});
	test_expansion(128'h83f62a964f7e72183c1e7478539e5b52, {16'd42712, 16'd14486, 16'd58267, 16'd9506, 16'd35892, 16'd39283, 16'd420, 16'd32903, 16'd6158, 16'd62396, 16'd20710, 16'd30910, 16'd37180, 16'd61573, 16'd39151, 16'd34550, 16'd56698, 16'd53834, 16'd64916, 16'd51695, 16'd15627, 16'd1963, 16'd7203, 16'd42959, 16'd16149, 16'd59459});
	test_expansion(128'hb324f0050f0aaedce59137421c6dd8d4, {16'd56725, 16'd13888, 16'd41776, 16'd20114, 16'd58106, 16'd18159, 16'd30329, 16'd53786, 16'd27638, 16'd26920, 16'd28053, 16'd15402, 16'd8136, 16'd64722, 16'd15520, 16'd55397, 16'd23371, 16'd11186, 16'd51831, 16'd50120, 16'd36097, 16'd57513, 16'd61880, 16'd16364, 16'd23979, 16'd5027});
	test_expansion(128'h9a2ef616dd49ee5bb7855fb370170909, {16'd58401, 16'd31173, 16'd50627, 16'd37692, 16'd17634, 16'd59772, 16'd30977, 16'd41421, 16'd38404, 16'd20404, 16'd56376, 16'd46659, 16'd16822, 16'd21558, 16'd1730, 16'd5722, 16'd50761, 16'd13875, 16'd30815, 16'd11184, 16'd31483, 16'd62502, 16'd30655, 16'd7866, 16'd13482, 16'd23550});
	test_expansion(128'hc83acdb0b56ada6155c6d107d4f3827d, {16'd421, 16'd31540, 16'd57747, 16'd13303, 16'd30299, 16'd6842, 16'd17288, 16'd43420, 16'd32575, 16'd20391, 16'd54589, 16'd60119, 16'd35768, 16'd18518, 16'd53614, 16'd14023, 16'd14430, 16'd24859, 16'd24572, 16'd51437, 16'd65051, 16'd16774, 16'd49909, 16'd28857, 16'd40896, 16'd15700});
	test_expansion(128'h8d12203f87641d4c2ba1a6fdc9bb4803, {16'd22698, 16'd55118, 16'd28074, 16'd13109, 16'd49667, 16'd51567, 16'd52359, 16'd11311, 16'd12921, 16'd23611, 16'd46335, 16'd4212, 16'd24063, 16'd26047, 16'd2364, 16'd55875, 16'd42659, 16'd31785, 16'd30603, 16'd59113, 16'd3655, 16'd43571, 16'd8781, 16'd59041, 16'd18222, 16'd43792});
	test_expansion(128'hf5886b86a0617b133f0c0a6639c639cb, {16'd45617, 16'd65391, 16'd64797, 16'd1271, 16'd1837, 16'd11822, 16'd65354, 16'd5191, 16'd10503, 16'd39180, 16'd6012, 16'd40433, 16'd18614, 16'd50527, 16'd17805, 16'd52563, 16'd27196, 16'd45696, 16'd38856, 16'd50062, 16'd28006, 16'd18945, 16'd1832, 16'd31006, 16'd37117, 16'd38989});
	test_expansion(128'h8c00e27f3119b40700b7e504d57210f5, {16'd10576, 16'd19973, 16'd3313, 16'd41935, 16'd31796, 16'd59372, 16'd20053, 16'd28033, 16'd58234, 16'd49650, 16'd31399, 16'd23333, 16'd5602, 16'd28248, 16'd37562, 16'd46159, 16'd15459, 16'd33991, 16'd14098, 16'd51247, 16'd41682, 16'd23985, 16'd10481, 16'd10139, 16'd31595, 16'd39586});
	test_expansion(128'he6599a77e251b55bbcd9cfb48dd32e85, {16'd60975, 16'd19723, 16'd2489, 16'd40748, 16'd10082, 16'd38584, 16'd32386, 16'd3673, 16'd48634, 16'd64817, 16'd27445, 16'd41414, 16'd3485, 16'd48499, 16'd25810, 16'd50224, 16'd4736, 16'd12352, 16'd33741, 16'd1132, 16'd23173, 16'd23711, 16'd61641, 16'd45438, 16'd43177, 16'd53770});
	test_expansion(128'ha878f018bab005c8af7200fe390dc186, {16'd7493, 16'd5457, 16'd35178, 16'd7322, 16'd18334, 16'd25501, 16'd52435, 16'd18599, 16'd24099, 16'd36245, 16'd9786, 16'd31373, 16'd46595, 16'd10822, 16'd44220, 16'd11654, 16'd906, 16'd23089, 16'd35017, 16'd48551, 16'd55314, 16'd32695, 16'd20225, 16'd29442, 16'd4770, 16'd29838});
	test_expansion(128'hb474f4667911e4350b4fe395d4cf75fc, {16'd54013, 16'd2471, 16'd3244, 16'd13854, 16'd38035, 16'd10101, 16'd38763, 16'd42171, 16'd7934, 16'd19707, 16'd11973, 16'd59231, 16'd32742, 16'd2928, 16'd25805, 16'd30590, 16'd28792, 16'd50063, 16'd4703, 16'd42195, 16'd39428, 16'd63892, 16'd51616, 16'd34485, 16'd36644, 16'd13592});
	test_expansion(128'h7aaae45258684f8f2b8e6ad46a39e1a6, {16'd64320, 16'd5119, 16'd30798, 16'd12765, 16'd54032, 16'd17626, 16'd56749, 16'd2160, 16'd586, 16'd5830, 16'd22222, 16'd42767, 16'd2550, 16'd27122, 16'd3618, 16'd47794, 16'd45862, 16'd30306, 16'd49913, 16'd15256, 16'd26419, 16'd25859, 16'd34035, 16'd54585, 16'd33375, 16'd46603});
	test_expansion(128'he3cb929fa3ff106de2bc823b9ee38727, {16'd26473, 16'd40173, 16'd38924, 16'd58639, 16'd53869, 16'd385, 16'd12843, 16'd30260, 16'd62910, 16'd10302, 16'd43572, 16'd25379, 16'd24660, 16'd11, 16'd62419, 16'd33827, 16'd58247, 16'd39661, 16'd48693, 16'd14829, 16'd61705, 16'd21864, 16'd719, 16'd16236, 16'd63433, 16'd64533});
	test_expansion(128'ha82c96b36813cb80cedeaaa2c1fa303c, {16'd15470, 16'd15655, 16'd59687, 16'd3559, 16'd25197, 16'd7860, 16'd51702, 16'd183, 16'd38958, 16'd58789, 16'd16994, 16'd28692, 16'd22394, 16'd1864, 16'd57172, 16'd26598, 16'd48785, 16'd29643, 16'd48127, 16'd13932, 16'd37469, 16'd29372, 16'd58155, 16'd28064, 16'd27699, 16'd5589});
	test_expansion(128'h0e6e9d59df6731b8a35f69eb16eadfea, {16'd28104, 16'd14111, 16'd58511, 16'd56987, 16'd18287, 16'd41170, 16'd20000, 16'd43573, 16'd29958, 16'd10057, 16'd10403, 16'd11920, 16'd42880, 16'd18124, 16'd16213, 16'd25553, 16'd5255, 16'd40747, 16'd29813, 16'd17166, 16'd4880, 16'd17801, 16'd4937, 16'd23462, 16'd34897, 16'd58726});
	test_expansion(128'h753c634fdd7eebd90a40c295155690fe, {16'd24798, 16'd37419, 16'd58931, 16'd20796, 16'd1950, 16'd33585, 16'd3511, 16'd56478, 16'd10105, 16'd22145, 16'd7868, 16'd7615, 16'd9215, 16'd40625, 16'd5997, 16'd61674, 16'd45096, 16'd46614, 16'd26207, 16'd2506, 16'd62743, 16'd50578, 16'd19116, 16'd63749, 16'd43257, 16'd5966});
	test_expansion(128'hf2e1e2310cd09066f2199614bd4e610d, {16'd47189, 16'd40593, 16'd22293, 16'd21543, 16'd3178, 16'd2161, 16'd32628, 16'd61206, 16'd61331, 16'd26139, 16'd60467, 16'd45584, 16'd57199, 16'd62848, 16'd42763, 16'd15102, 16'd4898, 16'd8185, 16'd11701, 16'd38164, 16'd54613, 16'd23666, 16'd54674, 16'd46733, 16'd7155, 16'd20002});
	test_expansion(128'hdef9a5f61d93bb3e0890d3be80215cce, {16'd42423, 16'd25316, 16'd53217, 16'd9645, 16'd13469, 16'd57709, 16'd54290, 16'd53159, 16'd7729, 16'd64728, 16'd4116, 16'd42305, 16'd56273, 16'd38283, 16'd58603, 16'd30298, 16'd34738, 16'd4492, 16'd10024, 16'd45189, 16'd20521, 16'd62028, 16'd51880, 16'd19226, 16'd27794, 16'd63234});
	test_expansion(128'h43db9197377d216ad2cba4db15ad1de8, {16'd1082, 16'd15689, 16'd33062, 16'd16853, 16'd11434, 16'd4017, 16'd50219, 16'd17897, 16'd53848, 16'd30534, 16'd28564, 16'd17884, 16'd29197, 16'd1885, 16'd58992, 16'd51465, 16'd11040, 16'd47620, 16'd15648, 16'd35078, 16'd31782, 16'd16669, 16'd50280, 16'd53555, 16'd42689, 16'd59384});
	test_expansion(128'hca6845fa876ef058f42e8a3886579a5e, {16'd59984, 16'd14530, 16'd20721, 16'd15715, 16'd64620, 16'd22166, 16'd38134, 16'd60575, 16'd3211, 16'd56475, 16'd7148, 16'd7781, 16'd59711, 16'd2438, 16'd20482, 16'd53037, 16'd47695, 16'd20229, 16'd34586, 16'd43682, 16'd13893, 16'd54988, 16'd4504, 16'd13119, 16'd28425, 16'd29355});
	test_expansion(128'h93f87c5ac67a99479196b94a6f185571, {16'd6057, 16'd49542, 16'd34025, 16'd15130, 16'd29297, 16'd6902, 16'd58289, 16'd12293, 16'd27859, 16'd23535, 16'd54358, 16'd25590, 16'd42552, 16'd11151, 16'd60376, 16'd49997, 16'd24285, 16'd14758, 16'd54012, 16'd60553, 16'd16524, 16'd44642, 16'd9042, 16'd11509, 16'd13899, 16'd2432});
	test_expansion(128'h4c37043f1534faf4c37011fee8ec9c24, {16'd22597, 16'd40915, 16'd18028, 16'd28515, 16'd41029, 16'd46651, 16'd63043, 16'd58004, 16'd4714, 16'd21873, 16'd2226, 16'd32830, 16'd52174, 16'd37619, 16'd50370, 16'd31255, 16'd19788, 16'd6814, 16'd35007, 16'd44838, 16'd5360, 16'd37535, 16'd65436, 16'd17558, 16'd17805, 16'd55414});
	test_expansion(128'h68dff0e99f9ab6c9446a984a14b7c88e, {16'd27506, 16'd43208, 16'd10788, 16'd19534, 16'd48012, 16'd14868, 16'd5963, 16'd61855, 16'd6157, 16'd39498, 16'd35214, 16'd18698, 16'd45506, 16'd7650, 16'd5676, 16'd58515, 16'd31871, 16'd44513, 16'd25210, 16'd1186, 16'd38346, 16'd51621, 16'd22707, 16'd59793, 16'd5395, 16'd5338});
	test_expansion(128'hfa9cd7293ac22bcdf63364db1f4a26e4, {16'd7041, 16'd6639, 16'd31757, 16'd34662, 16'd50407, 16'd13249, 16'd9365, 16'd135, 16'd49950, 16'd60291, 16'd17413, 16'd47609, 16'd65335, 16'd12989, 16'd3258, 16'd28707, 16'd58471, 16'd42221, 16'd31369, 16'd22257, 16'd39415, 16'd31961, 16'd20171, 16'd6342, 16'd11782, 16'd24638});
	test_expansion(128'h566cb83b86062499ea3c5b8430c271b4, {16'd38833, 16'd2139, 16'd11163, 16'd54784, 16'd59831, 16'd32919, 16'd12194, 16'd1226, 16'd8274, 16'd7085, 16'd17687, 16'd47127, 16'd29825, 16'd65179, 16'd14227, 16'd35959, 16'd48387, 16'd12692, 16'd58912, 16'd47928, 16'd3254, 16'd36000, 16'd45802, 16'd16973, 16'd10755, 16'd57099});
	test_expansion(128'hb982d6306e018939e2e8e9f80449114f, {16'd33178, 16'd8279, 16'd58279, 16'd54972, 16'd52974, 16'd25766, 16'd31545, 16'd42924, 16'd8819, 16'd10457, 16'd34002, 16'd26652, 16'd61310, 16'd64039, 16'd4874, 16'd14406, 16'd11117, 16'd30472, 16'd25547, 16'd29208, 16'd24245, 16'd47096, 16'd61420, 16'd36253, 16'd54420, 16'd62670});
	test_expansion(128'h291334628ccaafbb36b2a36324db9a94, {16'd44942, 16'd45414, 16'd7033, 16'd45111, 16'd25970, 16'd43183, 16'd53075, 16'd31900, 16'd39553, 16'd17666, 16'd37165, 16'd40777, 16'd46020, 16'd46671, 16'd47298, 16'd2791, 16'd24, 16'd55970, 16'd43988, 16'd46172, 16'd47341, 16'd44127, 16'd53326, 16'd5137, 16'd38060, 16'd61467});
	test_expansion(128'hce1c8f3668a7a8eae084b88cd95175da, {16'd41005, 16'd58848, 16'd61070, 16'd25156, 16'd24870, 16'd14351, 16'd62076, 16'd20309, 16'd29489, 16'd43231, 16'd29993, 16'd17670, 16'd57137, 16'd30183, 16'd18466, 16'd43036, 16'd17909, 16'd6470, 16'd34678, 16'd43115, 16'd31961, 16'd49939, 16'd25890, 16'd34647, 16'd1010, 16'd64042});
	test_expansion(128'h9917dfe19cc195faf36447bbfefa20eb, {16'd56068, 16'd4658, 16'd15512, 16'd56003, 16'd61, 16'd10307, 16'd9556, 16'd29857, 16'd58467, 16'd3519, 16'd22604, 16'd8117, 16'd29020, 16'd11746, 16'd36111, 16'd57681, 16'd58266, 16'd3813, 16'd63977, 16'd14780, 16'd612, 16'd1702, 16'd34154, 16'd24590, 16'd51377, 16'd52546});
	test_expansion(128'h0e0a0e232bc85b2f4ad23fe6a655129a, {16'd45762, 16'd24225, 16'd29015, 16'd61370, 16'd59183, 16'd2978, 16'd4567, 16'd22440, 16'd19754, 16'd2247, 16'd22618, 16'd63962, 16'd25801, 16'd12985, 16'd27743, 16'd41867, 16'd65436, 16'd38136, 16'd21724, 16'd680, 16'd39875, 16'd49185, 16'd15443, 16'd6277, 16'd23426, 16'd4583});
	test_expansion(128'hd6c081b17319b68cae000c1db48ea9c3, {16'd39719, 16'd42313, 16'd37673, 16'd9747, 16'd10987, 16'd43522, 16'd63576, 16'd60979, 16'd20494, 16'd7683, 16'd14021, 16'd20741, 16'd46600, 16'd22093, 16'd40174, 16'd65322, 16'd47881, 16'd54926, 16'd19705, 16'd20445, 16'd26410, 16'd14042, 16'd4330, 16'd47, 16'd27506, 16'd37694});
	test_expansion(128'h17b1ee5b02c422f306aa63cdda2c8480, {16'd5431, 16'd50623, 16'd56432, 16'd45183, 16'd22736, 16'd63651, 16'd33972, 16'd58580, 16'd17859, 16'd37787, 16'd42730, 16'd44965, 16'd24701, 16'd25308, 16'd48614, 16'd23982, 16'd32092, 16'd59515, 16'd21447, 16'd40752, 16'd45738, 16'd4157, 16'd52584, 16'd48906, 16'd42836, 16'd24753});
	test_expansion(128'hae31c4b2c303b61480136210c96df48b, {16'd59005, 16'd31372, 16'd59038, 16'd21920, 16'd54265, 16'd59143, 16'd16194, 16'd38953, 16'd57976, 16'd48026, 16'd51682, 16'd25427, 16'd29144, 16'd57374, 16'd52079, 16'd61416, 16'd28331, 16'd3527, 16'd23050, 16'd443, 16'd35419, 16'd33131, 16'd49494, 16'd49847, 16'd3344, 16'd14039});
	test_expansion(128'h593b66aea2ae4e3e9ce3bd88a49a1b63, {16'd32993, 16'd28220, 16'd9703, 16'd36892, 16'd59931, 16'd17992, 16'd18050, 16'd21078, 16'd40486, 16'd46987, 16'd62946, 16'd31710, 16'd50241, 16'd34399, 16'd29166, 16'd34369, 16'd21949, 16'd55312, 16'd61765, 16'd64904, 16'd58495, 16'd10527, 16'd57304, 16'd47811, 16'd29552, 16'd59301});
	test_expansion(128'h45e469b8fff8d48c010ccec48cc5754b, {16'd56562, 16'd32760, 16'd44985, 16'd53681, 16'd1775, 16'd42729, 16'd53382, 16'd59803, 16'd35833, 16'd36567, 16'd22517, 16'd14221, 16'd2151, 16'd12575, 16'd44338, 16'd44179, 16'd40856, 16'd355, 16'd26271, 16'd42421, 16'd39793, 16'd27394, 16'd16171, 16'd46064, 16'd18344, 16'd15889});
	test_expansion(128'h690e16c48b799c880baa237a5f085c60, {16'd10532, 16'd35650, 16'd53253, 16'd61525, 16'd53025, 16'd3057, 16'd56465, 16'd27816, 16'd34441, 16'd65269, 16'd3311, 16'd40661, 16'd31167, 16'd23962, 16'd60579, 16'd39675, 16'd9366, 16'd1129, 16'd50613, 16'd35576, 16'd15485, 16'd21956, 16'd31944, 16'd61321, 16'd65355, 16'd47022});
	test_expansion(128'h19cfe5cf73e245e861c66c464eb3c981, {16'd40286, 16'd26930, 16'd45609, 16'd2364, 16'd34095, 16'd7872, 16'd37005, 16'd56515, 16'd63821, 16'd23577, 16'd49609, 16'd6347, 16'd44200, 16'd23178, 16'd8215, 16'd20964, 16'd50040, 16'd44588, 16'd3740, 16'd7143, 16'd59654, 16'd48111, 16'd15786, 16'd3737, 16'd56602, 16'd21740});
	test_expansion(128'h734edb10b30270e084293fed594bf4b1, {16'd48496, 16'd17201, 16'd48136, 16'd62158, 16'd53146, 16'd42125, 16'd14629, 16'd58255, 16'd56413, 16'd63738, 16'd46990, 16'd62125, 16'd46364, 16'd7530, 16'd55853, 16'd49739, 16'd31048, 16'd19030, 16'd50004, 16'd50673, 16'd5041, 16'd52881, 16'd2733, 16'd18117, 16'd21124, 16'd6106});
	test_expansion(128'h3f496e859ec65be07fc71f4879345ca3, {16'd54748, 16'd28185, 16'd48198, 16'd10412, 16'd21257, 16'd63019, 16'd22593, 16'd54011, 16'd33378, 16'd24082, 16'd61796, 16'd39401, 16'd26859, 16'd43844, 16'd49973, 16'd54621, 16'd13906, 16'd45126, 16'd63375, 16'd12163, 16'd62488, 16'd46714, 16'd20701, 16'd33735, 16'd48497, 16'd48788});
	test_expansion(128'haea6dc3b695b14af7704338631f3d85b, {16'd30183, 16'd36912, 16'd65404, 16'd49516, 16'd5918, 16'd37839, 16'd56380, 16'd52455, 16'd50995, 16'd36674, 16'd40569, 16'd31231, 16'd3719, 16'd47669, 16'd3218, 16'd14170, 16'd42219, 16'd31994, 16'd11479, 16'd47843, 16'd9270, 16'd718, 16'd9951, 16'd43024, 16'd59554, 16'd54874});
	test_expansion(128'h8d4b0abce7344eb6edbf6d7082057f23, {16'd54685, 16'd19564, 16'd30025, 16'd30388, 16'd17173, 16'd14188, 16'd65196, 16'd12922, 16'd2915, 16'd40691, 16'd46340, 16'd53356, 16'd65138, 16'd38468, 16'd37513, 16'd16867, 16'd62325, 16'd45166, 16'd8563, 16'd30009, 16'd24843, 16'd24039, 16'd3882, 16'd65467, 16'd33391, 16'd8916});
	test_expansion(128'h1b88b21066edaca3329a8421246ee8dc, {16'd56663, 16'd7059, 16'd30602, 16'd61751, 16'd33790, 16'd19288, 16'd61494, 16'd26194, 16'd52471, 16'd11710, 16'd47586, 16'd61080, 16'd12553, 16'd7145, 16'd10660, 16'd42903, 16'd28240, 16'd50717, 16'd47634, 16'd36532, 16'd56286, 16'd33371, 16'd11470, 16'd52376, 16'd47302, 16'd44264});
	test_expansion(128'hb8ee2edce4cb44abd45f1afcb6928f62, {16'd2766, 16'd44702, 16'd17538, 16'd51317, 16'd61569, 16'd18078, 16'd53469, 16'd45668, 16'd51202, 16'd8354, 16'd34913, 16'd3298, 16'd54734, 16'd1603, 16'd9254, 16'd41483, 16'd54823, 16'd56356, 16'd20027, 16'd13884, 16'd55079, 16'd44379, 16'd32207, 16'd2265, 16'd34744, 16'd63628});
	test_expansion(128'hfdc99e82bcf9df05d052da8e2697da3f, {16'd35717, 16'd630, 16'd7920, 16'd39744, 16'd51428, 16'd14613, 16'd42874, 16'd47147, 16'd43849, 16'd46054, 16'd1950, 16'd12912, 16'd1118, 16'd64143, 16'd63582, 16'd48890, 16'd31653, 16'd58992, 16'd23615, 16'd49523, 16'd27221, 16'd2763, 16'd46996, 16'd53183, 16'd7053, 16'd62864});
	test_expansion(128'hf43611b0cd9b25b7f45d37e07772585e, {16'd19026, 16'd5071, 16'd62382, 16'd13710, 16'd12021, 16'd49837, 16'd60146, 16'd36402, 16'd34366, 16'd32360, 16'd18918, 16'd56526, 16'd20770, 16'd4042, 16'd48995, 16'd12486, 16'd14600, 16'd59932, 16'd27083, 16'd32302, 16'd43534, 16'd44605, 16'd16483, 16'd34393, 16'd10629, 16'd41737});
	test_expansion(128'hbca0441c256cd7cb9d7a2042a2d2e572, {16'd9618, 16'd48051, 16'd51836, 16'd38256, 16'd16071, 16'd33829, 16'd55857, 16'd16602, 16'd20758, 16'd52265, 16'd428, 16'd15278, 16'd23467, 16'd7360, 16'd9231, 16'd42033, 16'd31378, 16'd63914, 16'd29828, 16'd40851, 16'd30211, 16'd55182, 16'd50864, 16'd29555, 16'd17181, 16'd59708});
	test_expansion(128'hccdbdc3a0043f7b4cbf3945b46aa9064, {16'd9992, 16'd52494, 16'd17687, 16'd45812, 16'd34544, 16'd35668, 16'd31888, 16'd13085, 16'd60914, 16'd40790, 16'd39644, 16'd50622, 16'd31869, 16'd56330, 16'd51658, 16'd45199, 16'd28494, 16'd56362, 16'd36270, 16'd47313, 16'd27877, 16'd30182, 16'd65453, 16'd65172, 16'd9470, 16'd60748});
	test_expansion(128'h4fe8b2cd28cf985394c272b5ff203470, {16'd51853, 16'd36450, 16'd10576, 16'd14401, 16'd30916, 16'd31774, 16'd55245, 16'd47165, 16'd39905, 16'd10867, 16'd1951, 16'd62506, 16'd43601, 16'd55633, 16'd31114, 16'd6372, 16'd31031, 16'd64037, 16'd2834, 16'd58215, 16'd11467, 16'd389, 16'd34199, 16'd31124, 16'd15920, 16'd7748});
	test_expansion(128'hc2036453432691278d36d12848855b9c, {16'd55148, 16'd21935, 16'd35446, 16'd36102, 16'd48576, 16'd39554, 16'd17103, 16'd17861, 16'd32706, 16'd32176, 16'd9114, 16'd30871, 16'd43539, 16'd22304, 16'd27943, 16'd8979, 16'd11657, 16'd45423, 16'd53982, 16'd51408, 16'd5281, 16'd43911, 16'd17432, 16'd60724, 16'd29776, 16'd42153});
	test_expansion(128'h757966532e21f3db3b3cdaa1f18858e8, {16'd53053, 16'd18965, 16'd64237, 16'd38337, 16'd4075, 16'd46523, 16'd57346, 16'd34681, 16'd31165, 16'd29313, 16'd51757, 16'd15051, 16'd57355, 16'd10045, 16'd51346, 16'd638, 16'd38760, 16'd17415, 16'd187, 16'd60492, 16'd47222, 16'd8906, 16'd49246, 16'd1292, 16'd8534, 16'd53427});
	test_expansion(128'h960e354c3e55192d747c4e8991ac2a8f, {16'd63190, 16'd11817, 16'd20345, 16'd60181, 16'd32178, 16'd58673, 16'd18970, 16'd7032, 16'd63879, 16'd50175, 16'd30067, 16'd17189, 16'd30726, 16'd64725, 16'd2489, 16'd38784, 16'd44283, 16'd61215, 16'd18840, 16'd51361, 16'd19740, 16'd57405, 16'd13064, 16'd32363, 16'd43343, 16'd14590});
	test_expansion(128'had15a7c2c7a04dd16024dc025e636198, {16'd5532, 16'd62140, 16'd41716, 16'd15097, 16'd2585, 16'd11538, 16'd25811, 16'd14793, 16'd56161, 16'd53418, 16'd4852, 16'd51754, 16'd51664, 16'd991, 16'd49451, 16'd28159, 16'd225, 16'd64790, 16'd29160, 16'd50548, 16'd55981, 16'd16969, 16'd415, 16'd22503, 16'd51179, 16'd58780});
	test_expansion(128'h1a97c04cd55f1dbe7dc260e5f78a2971, {16'd59187, 16'd36656, 16'd16877, 16'd49856, 16'd21368, 16'd23166, 16'd31699, 16'd26630, 16'd7158, 16'd35442, 16'd55068, 16'd52467, 16'd28377, 16'd6701, 16'd26484, 16'd1026, 16'd41, 16'd64382, 16'd63468, 16'd11085, 16'd24301, 16'd458, 16'd17010, 16'd28540, 16'd40005, 16'd31330});
	test_expansion(128'h9b7124737833f36dfa5201d026a2717f, {16'd48455, 16'd20324, 16'd51747, 16'd60823, 16'd13868, 16'd39880, 16'd17370, 16'd25509, 16'd37196, 16'd3863, 16'd47720, 16'd23404, 16'd1261, 16'd18943, 16'd52717, 16'd27744, 16'd60112, 16'd26840, 16'd58234, 16'd51764, 16'd48460, 16'd31214, 16'd32099, 16'd38097, 16'd11609, 16'd35050});
	test_expansion(128'h0b05af6dc02d1b93ccd50ab2fe92fe68, {16'd50070, 16'd31763, 16'd5428, 16'd35332, 16'd34019, 16'd23037, 16'd330, 16'd5577, 16'd56337, 16'd28135, 16'd10964, 16'd64021, 16'd32935, 16'd2977, 16'd5219, 16'd24343, 16'd54025, 16'd47857, 16'd43588, 16'd5835, 16'd23338, 16'd18533, 16'd3619, 16'd47884, 16'd18429, 16'd55434});
	test_expansion(128'hdf4d8226d543aa5a23c588b03ea08648, {16'd37313, 16'd46414, 16'd22622, 16'd3709, 16'd60866, 16'd49920, 16'd34026, 16'd22853, 16'd58158, 16'd18307, 16'd64304, 16'd5906, 16'd15639, 16'd37256, 16'd2021, 16'd36892, 16'd8270, 16'd213, 16'd13553, 16'd13843, 16'd23930, 16'd24609, 16'd10707, 16'd43616, 16'd27063, 16'd53652});
	test_expansion(128'h8024ef9f4a5f7b253431fff9a1c443ca, {16'd30831, 16'd33919, 16'd64105, 16'd5016, 16'd4819, 16'd50986, 16'd19963, 16'd64367, 16'd31098, 16'd46386, 16'd41285, 16'd44651, 16'd15727, 16'd13555, 16'd6731, 16'd5074, 16'd53844, 16'd29942, 16'd6655, 16'd52851, 16'd64524, 16'd32405, 16'd10725, 16'd24048, 16'd10498, 16'd39118});
	test_expansion(128'hf94818d28fa5000c22326b70cac117ab, {16'd1732, 16'd60023, 16'd38409, 16'd52602, 16'd4516, 16'd29541, 16'd534, 16'd63385, 16'd40076, 16'd57347, 16'd40891, 16'd43098, 16'd58695, 16'd61135, 16'd41065, 16'd1875, 16'd59984, 16'd13642, 16'd19838, 16'd40371, 16'd55830, 16'd60455, 16'd63677, 16'd45266, 16'd59973, 16'd28244});
	test_expansion(128'h2cf4a2c9ad1bff534fe1e199ddd5a43c, {16'd27165, 16'd18697, 16'd14344, 16'd7778, 16'd5356, 16'd38105, 16'd59257, 16'd34924, 16'd15771, 16'd38543, 16'd60405, 16'd57034, 16'd5017, 16'd39748, 16'd41343, 16'd33711, 16'd26161, 16'd57195, 16'd62367, 16'd39003, 16'd65365, 16'd18350, 16'd978, 16'd53583, 16'd60845, 16'd34153});
	test_expansion(128'ha28eab1f4aedb454dbea9a9b91a9ceac, {16'd54306, 16'd53476, 16'd22061, 16'd17207, 16'd47320, 16'd12321, 16'd40290, 16'd28294, 16'd6089, 16'd3718, 16'd47659, 16'd11581, 16'd6280, 16'd17393, 16'd15145, 16'd48327, 16'd16812, 16'd59721, 16'd44174, 16'd47080, 16'd51192, 16'd15634, 16'd12657, 16'd32233, 16'd15613, 16'd24667});
	test_expansion(128'h27f0339d8f56660d93a1e7001b857175, {16'd44981, 16'd46596, 16'd3496, 16'd13790, 16'd6374, 16'd28537, 16'd8736, 16'd40501, 16'd22559, 16'd63146, 16'd27808, 16'd7752, 16'd47308, 16'd39308, 16'd36682, 16'd50455, 16'd32039, 16'd11707, 16'd3539, 16'd12267, 16'd28944, 16'd54535, 16'd53249, 16'd8405, 16'd53764, 16'd25127});
	test_expansion(128'h42441503cd1cfa6a0ef4e75f51183d32, {16'd11103, 16'd2418, 16'd58656, 16'd23710, 16'd36175, 16'd30754, 16'd7989, 16'd33670, 16'd44464, 16'd10497, 16'd19931, 16'd20792, 16'd13448, 16'd30732, 16'd49658, 16'd3440, 16'd21297, 16'd44903, 16'd46895, 16'd27490, 16'd39449, 16'd3138, 16'd61207, 16'd262, 16'd61370, 16'd21296});
	test_expansion(128'h80add6e08b3c58df6bdc6547bc34f6c5, {16'd59589, 16'd43519, 16'd42048, 16'd30727, 16'd62846, 16'd33851, 16'd31162, 16'd21718, 16'd30908, 16'd3280, 16'd23525, 16'd24754, 16'd11571, 16'd62664, 16'd61400, 16'd60455, 16'd18587, 16'd16849, 16'd37355, 16'd53955, 16'd35201, 16'd18399, 16'd60701, 16'd57431, 16'd33748, 16'd47144});
	test_expansion(128'hd57f9b67fc49ec330ebf0ece976099e6, {16'd38761, 16'd21362, 16'd9760, 16'd36671, 16'd429, 16'd43093, 16'd63790, 16'd59097, 16'd21469, 16'd3243, 16'd61099, 16'd43372, 16'd63106, 16'd60123, 16'd28004, 16'd57556, 16'd24742, 16'd17307, 16'd4055, 16'd20165, 16'd22197, 16'd17911, 16'd835, 16'd20601, 16'd14795, 16'd45065});
	test_expansion(128'h5ca06e38687f37b57eb3b6d7ac26f842, {16'd48814, 16'd34412, 16'd36224, 16'd62578, 16'd14025, 16'd64981, 16'd2373, 16'd65257, 16'd49711, 16'd13319, 16'd4037, 16'd41510, 16'd23972, 16'd22179, 16'd39246, 16'd26399, 16'd30648, 16'd16779, 16'd17699, 16'd36593, 16'd9000, 16'd57973, 16'd48963, 16'd33409, 16'd52019, 16'd39547});
	test_expansion(128'h119df087cc924eb2a71c58b2b0be47bf, {16'd48143, 16'd22036, 16'd51150, 16'd27947, 16'd19578, 16'd18714, 16'd54075, 16'd6023, 16'd27430, 16'd45079, 16'd28895, 16'd46851, 16'd7175, 16'd45279, 16'd50219, 16'd16371, 16'd39788, 16'd51858, 16'd11365, 16'd47142, 16'd18326, 16'd47953, 16'd33112, 16'd50571, 16'd40882, 16'd48905});
	test_expansion(128'h14f5e7c78b8e1893d714b85e346eec8e, {16'd2189, 16'd57830, 16'd27806, 16'd18615, 16'd55470, 16'd1158, 16'd46265, 16'd63687, 16'd24846, 16'd3734, 16'd5279, 16'd6351, 16'd52953, 16'd12070, 16'd50905, 16'd228, 16'd49734, 16'd20672, 16'd24840, 16'd62038, 16'd10559, 16'd31857, 16'd56605, 16'd13862, 16'd2301, 16'd22725});
	test_expansion(128'hcadd49fa765ad943997127220915fa28, {16'd54606, 16'd13990, 16'd22798, 16'd55400, 16'd50337, 16'd53869, 16'd38528, 16'd40796, 16'd27009, 16'd2340, 16'd9035, 16'd50847, 16'd64437, 16'd53413, 16'd38780, 16'd12726, 16'd11606, 16'd28946, 16'd60590, 16'd19746, 16'd5420, 16'd16167, 16'd49962, 16'd5882, 16'd50648, 16'd30099});
	test_expansion(128'h43634218b15fba478a615fa3b9c06f46, {16'd22515, 16'd32683, 16'd58955, 16'd6152, 16'd3437, 16'd38553, 16'd27924, 16'd61919, 16'd5551, 16'd42093, 16'd37091, 16'd56147, 16'd42894, 16'd24363, 16'd3685, 16'd37264, 16'd13144, 16'd54669, 16'd36449, 16'd16706, 16'd15423, 16'd62115, 16'd35650, 16'd34989, 16'd5381, 16'd26500});
	test_expansion(128'h537de4b086f887aff1f98765cb7c1d37, {16'd40687, 16'd42026, 16'd64277, 16'd21688, 16'd16642, 16'd23382, 16'd31337, 16'd10276, 16'd51163, 16'd31348, 16'd35891, 16'd18496, 16'd45619, 16'd62737, 16'd4205, 16'd49608, 16'd49277, 16'd16266, 16'd49435, 16'd62428, 16'd41319, 16'd16770, 16'd18894, 16'd27786, 16'd32787, 16'd34902});
	test_expansion(128'h1b8608f12b15a17a516296174563a572, {16'd14249, 16'd61135, 16'd63899, 16'd24108, 16'd20448, 16'd48850, 16'd17638, 16'd46652, 16'd55462, 16'd40649, 16'd52106, 16'd55352, 16'd41468, 16'd30849, 16'd40204, 16'd3416, 16'd9501, 16'd2027, 16'd20397, 16'd58727, 16'd61753, 16'd26896, 16'd3002, 16'd35004, 16'd31057, 16'd20575});
	test_expansion(128'ha797c428dbb90ebe3f90f6f3c764a545, {16'd47691, 16'd12824, 16'd48960, 16'd64904, 16'd4523, 16'd45670, 16'd56316, 16'd24888, 16'd56863, 16'd62367, 16'd49929, 16'd45521, 16'd58849, 16'd13369, 16'd20536, 16'd10835, 16'd2575, 16'd22181, 16'd39571, 16'd54146, 16'd1687, 16'd58421, 16'd9702, 16'd23537, 16'd39926, 16'd49183});
	test_expansion(128'h377143ed8a9eab8a95118e3b6bd41ae6, {16'd9396, 16'd29997, 16'd29645, 16'd53634, 16'd24557, 16'd53018, 16'd50955, 16'd15571, 16'd54464, 16'd33530, 16'd64135, 16'd21256, 16'd47580, 16'd35948, 16'd4122, 16'd3950, 16'd5124, 16'd49351, 16'd12502, 16'd25528, 16'd28640, 16'd14864, 16'd44857, 16'd47708, 16'd47320, 16'd26391});
	test_expansion(128'h16b105bcbde295e5e9b76ae5335fc811, {16'd30004, 16'd46309, 16'd39994, 16'd34795, 16'd43342, 16'd30221, 16'd47878, 16'd41723, 16'd12448, 16'd4916, 16'd59270, 16'd21031, 16'd41106, 16'd36286, 16'd44226, 16'd26852, 16'd47132, 16'd10752, 16'd16227, 16'd17292, 16'd54509, 16'd51485, 16'd25850, 16'd49608, 16'd49559, 16'd50579});
	test_expansion(128'h38fa5ce96db5b2c65f6484578adc473d, {16'd30472, 16'd16288, 16'd12475, 16'd24687, 16'd55194, 16'd10382, 16'd4588, 16'd39072, 16'd19794, 16'd5898, 16'd40518, 16'd2068, 16'd45039, 16'd38510, 16'd28760, 16'd11611, 16'd6416, 16'd5814, 16'd64086, 16'd4246, 16'd211, 16'd49735, 16'd2272, 16'd47731, 16'd19985, 16'd60328});
	test_expansion(128'h18ee2b588a997ad61e556b2946001e28, {16'd51106, 16'd1299, 16'd37721, 16'd29001, 16'd301, 16'd16877, 16'd26135, 16'd44442, 16'd61395, 16'd32408, 16'd6360, 16'd65289, 16'd28090, 16'd26819, 16'd37720, 16'd42041, 16'd59526, 16'd11950, 16'd61797, 16'd60323, 16'd42613, 16'd43669, 16'd39891, 16'd53582, 16'd50705, 16'd49750});
	test_expansion(128'hbb415c4bee39e9a4f03a2d0225442d3d, {16'd40994, 16'd46989, 16'd18480, 16'd44527, 16'd21280, 16'd43025, 16'd58141, 16'd65484, 16'd51549, 16'd57418, 16'd20829, 16'd46331, 16'd26676, 16'd61670, 16'd36267, 16'd13894, 16'd28131, 16'd33056, 16'd23504, 16'd24039, 16'd50195, 16'd6554, 16'd45120, 16'd10096, 16'd17786, 16'd42965});
	test_expansion(128'h6b067808a6b8b8dc37cc904362e0e9fa, {16'd40184, 16'd5181, 16'd57215, 16'd13580, 16'd3582, 16'd59926, 16'd1689, 16'd14718, 16'd4755, 16'd53192, 16'd55606, 16'd59082, 16'd36404, 16'd4163, 16'd50392, 16'd64659, 16'd36387, 16'd47872, 16'd12929, 16'd4604, 16'd8488, 16'd14382, 16'd40067, 16'd8455, 16'd22502, 16'd58130});
	test_expansion(128'h0bae38c1683a6683d0542a9492583558, {16'd57497, 16'd44844, 16'd55719, 16'd35688, 16'd56052, 16'd58249, 16'd53357, 16'd55353, 16'd54262, 16'd23928, 16'd32332, 16'd36824, 16'd43599, 16'd58894, 16'd21334, 16'd15824, 16'd60853, 16'd6222, 16'd65321, 16'd58082, 16'd57001, 16'd26715, 16'd48527, 16'd20518, 16'd892, 16'd39274});
	test_expansion(128'ha60f34836d4448d3002064403ad6f903, {16'd24400, 16'd253, 16'd63744, 16'd54071, 16'd57579, 16'd28048, 16'd63156, 16'd45297, 16'd45357, 16'd4841, 16'd32849, 16'd48097, 16'd65311, 16'd49952, 16'd19040, 16'd41440, 16'd20364, 16'd707, 16'd53958, 16'd12779, 16'd29030, 16'd13586, 16'd51797, 16'd59328, 16'd26411, 16'd9873});
	test_expansion(128'hf42b12ab50b659071e10c079ddcbb02d, {16'd14417, 16'd34304, 16'd18711, 16'd14222, 16'd17656, 16'd45854, 16'd24656, 16'd51820, 16'd18206, 16'd9705, 16'd42574, 16'd43826, 16'd63608, 16'd35000, 16'd62622, 16'd37288, 16'd51148, 16'd27572, 16'd17407, 16'd62665, 16'd13862, 16'd51618, 16'd63812, 16'd29760, 16'd833, 16'd3553});
	test_expansion(128'hbae27518bad15407533e435705ca5f8c, {16'd11207, 16'd33682, 16'd30448, 16'd34994, 16'd35213, 16'd30533, 16'd54034, 16'd44971, 16'd55309, 16'd54678, 16'd35566, 16'd38217, 16'd45940, 16'd31685, 16'd30123, 16'd16771, 16'd62464, 16'd29554, 16'd62790, 16'd2252, 16'd19059, 16'd27196, 16'd46734, 16'd15769, 16'd24474, 16'd43927});
	test_expansion(128'h2c9802df2c80d2daf66e1c87621139cd, {16'd44154, 16'd19814, 16'd30373, 16'd43551, 16'd37669, 16'd38837, 16'd8117, 16'd34995, 16'd57896, 16'd19588, 16'd10147, 16'd62091, 16'd57842, 16'd31419, 16'd57093, 16'd64680, 16'd15569, 16'd7909, 16'd34566, 16'd64430, 16'd58562, 16'd44082, 16'd24616, 16'd1809, 16'd30560, 16'd35859});
	test_expansion(128'h48794a88694089221a477503d96e355b, {16'd15311, 16'd32418, 16'd28244, 16'd25531, 16'd11598, 16'd46591, 16'd15942, 16'd18356, 16'd56705, 16'd28072, 16'd15819, 16'd41840, 16'd46512, 16'd36189, 16'd22989, 16'd57028, 16'd36806, 16'd33042, 16'd50492, 16'd28955, 16'd55748, 16'd2391, 16'd34810, 16'd11580, 16'd42960, 16'd49073});
	test_expansion(128'hfebfe7b0f9115ef68f3217de71323bbf, {16'd28084, 16'd54998, 16'd52303, 16'd26639, 16'd40373, 16'd33763, 16'd45084, 16'd49059, 16'd20250, 16'd12658, 16'd5145, 16'd50663, 16'd25945, 16'd64, 16'd64491, 16'd12937, 16'd2452, 16'd29176, 16'd52886, 16'd31407, 16'd10530, 16'd25815, 16'd132, 16'd53483, 16'd35749, 16'd12663});
	test_expansion(128'h81d7a09b43d2d3d5af21ea18bc9ed74d, {16'd43967, 16'd52442, 16'd63146, 16'd60001, 16'd63203, 16'd23006, 16'd16453, 16'd14249, 16'd49284, 16'd39783, 16'd50708, 16'd9443, 16'd31875, 16'd55555, 16'd57185, 16'd8215, 16'd52446, 16'd31858, 16'd62263, 16'd16540, 16'd19347, 16'd29747, 16'd14346, 16'd24769, 16'd36869, 16'd62204});
	test_expansion(128'h17390e1f2e2fde2ce246f9f0615107ab, {16'd36515, 16'd57781, 16'd46510, 16'd53655, 16'd37096, 16'd710, 16'd10593, 16'd49803, 16'd25674, 16'd48999, 16'd46683, 16'd19154, 16'd30042, 16'd59550, 16'd50523, 16'd34506, 16'd50202, 16'd32556, 16'd62660, 16'd294, 16'd13318, 16'd37383, 16'd60771, 16'd8056, 16'd28210, 16'd32046});
	test_expansion(128'h8b879228c8c981e4ebebbaee4957ee97, {16'd36201, 16'd49214, 16'd32066, 16'd47136, 16'd2185, 16'd30253, 16'd49699, 16'd23500, 16'd53097, 16'd12442, 16'd10100, 16'd49109, 16'd41878, 16'd51140, 16'd8454, 16'd49225, 16'd18627, 16'd33430, 16'd56216, 16'd5401, 16'd61211, 16'd21265, 16'd40445, 16'd30882, 16'd14861, 16'd32022});
	test_expansion(128'hfb297e5e74b0988deeff8df1517d2011, {16'd55045, 16'd24887, 16'd28796, 16'd30097, 16'd62957, 16'd49984, 16'd59054, 16'd44874, 16'd4139, 16'd39808, 16'd10031, 16'd23189, 16'd43706, 16'd19902, 16'd29868, 16'd64821, 16'd56696, 16'd56670, 16'd50628, 16'd26810, 16'd46476, 16'd64172, 16'd47692, 16'd65489, 16'd63324, 16'd38931});
	test_expansion(128'hf95a83f61ef7c6cc943ed4254bb3b77f, {16'd19792, 16'd31614, 16'd8889, 16'd14958, 16'd27898, 16'd2476, 16'd18004, 16'd50955, 16'd12649, 16'd54436, 16'd29853, 16'd45478, 16'd31458, 16'd29111, 16'd962, 16'd32204, 16'd60331, 16'd56442, 16'd53951, 16'd12264, 16'd14985, 16'd43320, 16'd36430, 16'd44221, 16'd13798, 16'd48152});
	test_expansion(128'hf837af0b416e1053d3e2dd8c70f79072, {16'd38270, 16'd22752, 16'd20563, 16'd62990, 16'd59550, 16'd50867, 16'd3049, 16'd20708, 16'd58331, 16'd21108, 16'd64768, 16'd17567, 16'd22987, 16'd43898, 16'd15765, 16'd61610, 16'd56434, 16'd29663, 16'd37648, 16'd40772, 16'd22007, 16'd13624, 16'd64530, 16'd38247, 16'd51496, 16'd43608});
	test_expansion(128'hd34092468810941e58d9ef14297d4f1d, {16'd18571, 16'd58309, 16'd13180, 16'd4532, 16'd20748, 16'd18785, 16'd31267, 16'd62233, 16'd56375, 16'd31152, 16'd38426, 16'd2712, 16'd49104, 16'd16965, 16'd53692, 16'd39580, 16'd26460, 16'd65483, 16'd21398, 16'd59708, 16'd58908, 16'd59750, 16'd62215, 16'd60647, 16'd64038, 16'd45592});
	test_expansion(128'h2b60fa8e651c18c5de2b9488352e9d22, {16'd26725, 16'd22003, 16'd43051, 16'd24317, 16'd5815, 16'd59791, 16'd33524, 16'd38379, 16'd46095, 16'd47764, 16'd5879, 16'd5562, 16'd43720, 16'd44394, 16'd48176, 16'd41078, 16'd42620, 16'd49916, 16'd10637, 16'd21360, 16'd15396, 16'd65412, 16'd62178, 16'd3388, 16'd58936, 16'd37632});
	test_expansion(128'hfcdd7f5f85fe31f5096f1ca4ad3a0fc5, {16'd45302, 16'd40108, 16'd481, 16'd8890, 16'd36389, 16'd41853, 16'd42740, 16'd34236, 16'd46939, 16'd10692, 16'd34024, 16'd13185, 16'd2015, 16'd42997, 16'd59546, 16'd44717, 16'd23454, 16'd6053, 16'd1698, 16'd45089, 16'd6634, 16'd20635, 16'd19397, 16'd16584, 16'd13492, 16'd42958});
	test_expansion(128'h214ed0dc54fccd548322d2a0584cce4c, {16'd46976, 16'd20386, 16'd31691, 16'd21827, 16'd17730, 16'd2796, 16'd64, 16'd14500, 16'd1839, 16'd27884, 16'd12373, 16'd43462, 16'd50090, 16'd42013, 16'd6951, 16'd21081, 16'd65359, 16'd13193, 16'd12611, 16'd42546, 16'd20061, 16'd47776, 16'd51959, 16'd64194, 16'd40132, 16'd48954});
	test_expansion(128'h08e594b3d5e92c62fcd424d75c967122, {16'd54461, 16'd38194, 16'd29823, 16'd44915, 16'd21647, 16'd8037, 16'd60213, 16'd10562, 16'd35979, 16'd29613, 16'd17687, 16'd40069, 16'd33996, 16'd31216, 16'd61581, 16'd28949, 16'd9625, 16'd13427, 16'd43995, 16'd40813, 16'd21214, 16'd8458, 16'd11432, 16'd41008, 16'd31959, 16'd41379});
	test_expansion(128'hf631b78a3fe1e68d334b9aa7386c0b55, {16'd64915, 16'd44723, 16'd36165, 16'd17041, 16'd28241, 16'd34641, 16'd54718, 16'd2953, 16'd39054, 16'd23663, 16'd21392, 16'd4388, 16'd10419, 16'd32945, 16'd8360, 16'd8371, 16'd64626, 16'd39309, 16'd16791, 16'd16531, 16'd61264, 16'd52082, 16'd60139, 16'd2284, 16'd54931, 16'd3204});
	test_expansion(128'h034307e75c45b0aaaff0a34f776e5bb2, {16'd17420, 16'd2522, 16'd36443, 16'd23547, 16'd60632, 16'd59144, 16'd14406, 16'd23043, 16'd30701, 16'd64923, 16'd12357, 16'd55817, 16'd29648, 16'd51531, 16'd60821, 16'd2434, 16'd41468, 16'd7991, 16'd59511, 16'd63940, 16'd51628, 16'd35957, 16'd41339, 16'd56178, 16'd18007, 16'd56684});
	test_expansion(128'hc04961f4d3e3097c3b3c492edc38af9a, {16'd16381, 16'd60872, 16'd30193, 16'd9121, 16'd37413, 16'd45490, 16'd60248, 16'd29687, 16'd14618, 16'd7152, 16'd56944, 16'd59903, 16'd54188, 16'd13808, 16'd17898, 16'd57778, 16'd38946, 16'd21579, 16'd13419, 16'd48365, 16'd38249, 16'd39895, 16'd26389, 16'd52535, 16'd36574, 16'd30191});
	test_expansion(128'hdc1d245f9c6ed613e45650398f27e252, {16'd25746, 16'd8659, 16'd50787, 16'd16012, 16'd60809, 16'd26021, 16'd7653, 16'd58419, 16'd34628, 16'd35293, 16'd41290, 16'd53791, 16'd8856, 16'd46616, 16'd25025, 16'd20250, 16'd30549, 16'd32517, 16'd25270, 16'd19789, 16'd64705, 16'd23821, 16'd44350, 16'd49392, 16'd28392, 16'd34781});
	test_expansion(128'h0eb8cc4fad19c56b73fd34318678bf4a, {16'd57628, 16'd47200, 16'd12221, 16'd54016, 16'd11411, 16'd19453, 16'd24100, 16'd49087, 16'd36198, 16'd14403, 16'd25345, 16'd9336, 16'd38250, 16'd54928, 16'd18584, 16'd19294, 16'd58720, 16'd35018, 16'd42207, 16'd61558, 16'd34560, 16'd11587, 16'd25315, 16'd15449, 16'd15592, 16'd57170});
	test_expansion(128'h800e721bde3698238f0dfa9ae228924e, {16'd28006, 16'd63279, 16'd37122, 16'd25570, 16'd40392, 16'd12511, 16'd24596, 16'd61033, 16'd4067, 16'd56689, 16'd25348, 16'd61473, 16'd34839, 16'd40779, 16'd47237, 16'd41447, 16'd7919, 16'd61563, 16'd20588, 16'd41740, 16'd50557, 16'd11133, 16'd33446, 16'd9465, 16'd20439, 16'd53568});
	test_expansion(128'h14d2db181d7d07bc89eb5dac5fdf299c, {16'd24773, 16'd47502, 16'd64130, 16'd32007, 16'd59319, 16'd65351, 16'd9857, 16'd2341, 16'd64854, 16'd23806, 16'd25941, 16'd4035, 16'd52122, 16'd32783, 16'd6314, 16'd26308, 16'd29525, 16'd45091, 16'd57030, 16'd181, 16'd8654, 16'd40172, 16'd41750, 16'd11899, 16'd19923, 16'd12617});
	test_expansion(128'ha74d5091444047e8eafbb575dea41b65, {16'd25242, 16'd1991, 16'd63918, 16'd7832, 16'd13242, 16'd14267, 16'd19210, 16'd5266, 16'd6268, 16'd43256, 16'd415, 16'd13906, 16'd16253, 16'd9169, 16'd20875, 16'd31812, 16'd57874, 16'd56684, 16'd52625, 16'd17978, 16'd22337, 16'd37804, 16'd35901, 16'd34738, 16'd24202, 16'd53428});
	test_expansion(128'h42ca3d852c03a5a39a458159c9e286b6, {16'd36345, 16'd7973, 16'd56499, 16'd10255, 16'd38497, 16'd7439, 16'd36710, 16'd43673, 16'd22896, 16'd2186, 16'd32193, 16'd38387, 16'd62345, 16'd23767, 16'd30742, 16'd8386, 16'd5308, 16'd6631, 16'd24440, 16'd64759, 16'd14388, 16'd55590, 16'd36509, 16'd10347, 16'd11253, 16'd17149});
	test_expansion(128'h0feee44ceec34a73ff761355de3d9848, {16'd15535, 16'd44444, 16'd23332, 16'd35335, 16'd13061, 16'd17356, 16'd49732, 16'd49309, 16'd38156, 16'd25253, 16'd61291, 16'd9962, 16'd55430, 16'd36561, 16'd21447, 16'd13130, 16'd16708, 16'd39717, 16'd35487, 16'd26216, 16'd23720, 16'd62077, 16'd43931, 16'd15267, 16'd15, 16'd42238});
	test_expansion(128'h069ffb707aa8fcf34cbaca772d9dee99, {16'd14259, 16'd53012, 16'd3686, 16'd46086, 16'd56502, 16'd59796, 16'd65225, 16'd31827, 16'd58341, 16'd38831, 16'd20807, 16'd31548, 16'd26001, 16'd3207, 16'd64837, 16'd8303, 16'd41910, 16'd25384, 16'd44220, 16'd34011, 16'd57727, 16'd21563, 16'd53744, 16'd57084, 16'd9551, 16'd21189});
	test_expansion(128'h6dcc8ead508332223a9d205baa1e7a92, {16'd58657, 16'd48515, 16'd15163, 16'd58640, 16'd34186, 16'd11921, 16'd22763, 16'd39715, 16'd49555, 16'd31263, 16'd41439, 16'd64341, 16'd41520, 16'd61287, 16'd59104, 16'd58883, 16'd15297, 16'd2087, 16'd33701, 16'd6857, 16'd56083, 16'd54007, 16'd42189, 16'd20907, 16'd47018, 16'd44970});
	test_expansion(128'h7385e7be2ef4a35cc60a398c432c0371, {16'd15633, 16'd8697, 16'd55034, 16'd44518, 16'd64339, 16'd26383, 16'd17308, 16'd61390, 16'd4482, 16'd54553, 16'd36936, 16'd7040, 16'd47702, 16'd29662, 16'd36170, 16'd43673, 16'd27652, 16'd37138, 16'd15114, 16'd19575, 16'd22846, 16'd30711, 16'd32267, 16'd60094, 16'd29474, 16'd31707});
	test_expansion(128'h08626a27b761ddc4451a0056d1eadaa0, {16'd59945, 16'd52365, 16'd47855, 16'd61442, 16'd14903, 16'd16886, 16'd43526, 16'd47782, 16'd32776, 16'd4634, 16'd44544, 16'd33381, 16'd43712, 16'd43966, 16'd44230, 16'd35314, 16'd49847, 16'd51323, 16'd783, 16'd65134, 16'd57775, 16'd29248, 16'd12210, 16'd2056, 16'd52783, 16'd50776});
	test_expansion(128'h5a9272b1b7ee7c6b5d618d833d7abf7d, {16'd13918, 16'd5560, 16'd6560, 16'd2962, 16'd58347, 16'd65214, 16'd14058, 16'd52234, 16'd20947, 16'd18452, 16'd25730, 16'd29588, 16'd61651, 16'd13875, 16'd21793, 16'd62633, 16'd60996, 16'd48253, 16'd29141, 16'd11223, 16'd59652, 16'd29186, 16'd4037, 16'd34979, 16'd21793, 16'd1672});
	test_expansion(128'h68682ff186fcd100e2f49996ea8e4c07, {16'd64675, 16'd64910, 16'd12595, 16'd33304, 16'd46148, 16'd9673, 16'd1313, 16'd57750, 16'd52542, 16'd18459, 16'd4623, 16'd36838, 16'd64323, 16'd9980, 16'd37268, 16'd57141, 16'd53409, 16'd55836, 16'd53268, 16'd22203, 16'd8782, 16'd19744, 16'd50385, 16'd40999, 16'd32521, 16'd18558});
	test_expansion(128'hba18214868707b96916bccbb364e0df8, {16'd43358, 16'd11101, 16'd48340, 16'd34279, 16'd16060, 16'd37712, 16'd53014, 16'd39305, 16'd8775, 16'd19863, 16'd4994, 16'd31066, 16'd17395, 16'd23286, 16'd98, 16'd46914, 16'd31410, 16'd45003, 16'd31969, 16'd27982, 16'd36430, 16'd23395, 16'd51442, 16'd10595, 16'd63722, 16'd39947});
	test_expansion(128'hbf03f5a14bdf6958908884f78de7e9f9, {16'd56241, 16'd25586, 16'd10504, 16'd5951, 16'd33270, 16'd53225, 16'd32516, 16'd33309, 16'd35565, 16'd2171, 16'd52686, 16'd33588, 16'd27986, 16'd47685, 16'd49693, 16'd32403, 16'd35351, 16'd9080, 16'd34151, 16'd39558, 16'd926, 16'd37049, 16'd10563, 16'd34710, 16'd29832, 16'd41784});
	test_expansion(128'hc0621650a25ec7feec710c3c693ea90a, {16'd15134, 16'd11102, 16'd59404, 16'd650, 16'd41235, 16'd34475, 16'd23968, 16'd36136, 16'd60687, 16'd2630, 16'd59384, 16'd8337, 16'd30079, 16'd4242, 16'd60415, 16'd52346, 16'd27501, 16'd49843, 16'd53472, 16'd46736, 16'd26413, 16'd18242, 16'd53352, 16'd4372, 16'd55650, 16'd4703});
	test_expansion(128'h9e03d01a5610d34b4b8fef0534113285, {16'd48611, 16'd48911, 16'd50785, 16'd5734, 16'd4359, 16'd8865, 16'd56322, 16'd36041, 16'd59544, 16'd34162, 16'd49818, 16'd44515, 16'd39360, 16'd55062, 16'd61042, 16'd63194, 16'd42081, 16'd14039, 16'd20799, 16'd58482, 16'd63454, 16'd36840, 16'd32231, 16'd54275, 16'd2133, 16'd10578});
	test_expansion(128'h47c7ddb8337926f73735f47d29097d7b, {16'd8862, 16'd33484, 16'd58931, 16'd41995, 16'd10661, 16'd40795, 16'd61252, 16'd11162, 16'd5866, 16'd29094, 16'd45583, 16'd6738, 16'd4185, 16'd32279, 16'd45926, 16'd26842, 16'd44391, 16'd19057, 16'd50403, 16'd23964, 16'd37857, 16'd28985, 16'd21778, 16'd48995, 16'd9847, 16'd34871});
	test_expansion(128'h4a1e681f56f83a65d21a7af46896891d, {16'd24613, 16'd4728, 16'd21387, 16'd44277, 16'd7088, 16'd23744, 16'd16114, 16'd37487, 16'd31752, 16'd31356, 16'd26042, 16'd33844, 16'd39980, 16'd34095, 16'd7065, 16'd6035, 16'd63223, 16'd57286, 16'd28288, 16'd15654, 16'd22326, 16'd16857, 16'd61402, 16'd39232, 16'd1285, 16'd15847});
	test_expansion(128'h7287ec1cdf76f2581a8a40bc070c3099, {16'd10016, 16'd54036, 16'd2607, 16'd2957, 16'd18392, 16'd47427, 16'd30968, 16'd61723, 16'd17491, 16'd1810, 16'd14619, 16'd16812, 16'd58272, 16'd1441, 16'd844, 16'd31554, 16'd22839, 16'd53982, 16'd50894, 16'd29353, 16'd21009, 16'd37515, 16'd18422, 16'd54322, 16'd52214, 16'd636});
	test_expansion(128'he6a64a6f69899213546266e283f11d6e, {16'd6264, 16'd26150, 16'd53837, 16'd26562, 16'd5459, 16'd16554, 16'd932, 16'd35928, 16'd26851, 16'd42166, 16'd31003, 16'd21372, 16'd8535, 16'd3580, 16'd29586, 16'd1726, 16'd918, 16'd34003, 16'd18829, 16'd28799, 16'd45304, 16'd20901, 16'd55893, 16'd61673, 16'd16339, 16'd44619});
	test_expansion(128'h4a941b176b3d1971149dd0d501dba63e, {16'd22576, 16'd36629, 16'd6599, 16'd49378, 16'd47522, 16'd55679, 16'd2072, 16'd27192, 16'd61705, 16'd45427, 16'd3231, 16'd56869, 16'd40055, 16'd40298, 16'd54102, 16'd20657, 16'd49626, 16'd18147, 16'd38421, 16'd12887, 16'd28114, 16'd25257, 16'd51072, 16'd42174, 16'd56122, 16'd16015});
	test_expansion(128'hb13c2ccb5f49679c0cad8f820f441e07, {16'd1361, 16'd29786, 16'd60933, 16'd51257, 16'd4667, 16'd53500, 16'd671, 16'd39618, 16'd12894, 16'd18917, 16'd6909, 16'd59981, 16'd45428, 16'd15763, 16'd62945, 16'd7173, 16'd60138, 16'd61233, 16'd23744, 16'd31294, 16'd36790, 16'd294, 16'd18984, 16'd40442, 16'd13511, 16'd39876});
	test_expansion(128'h643b719f6061d53ff13a2ba9395a56d7, {16'd19884, 16'd61333, 16'd61518, 16'd16623, 16'd63499, 16'd33618, 16'd46661, 16'd20716, 16'd25968, 16'd45537, 16'd52793, 16'd33966, 16'd30536, 16'd56252, 16'd29137, 16'd9884, 16'd1721, 16'd64961, 16'd33781, 16'd49263, 16'd25777, 16'd29690, 16'd18353, 16'd48911, 16'd64698, 16'd7249});
	test_expansion(128'hbfa726bb65057559127843e369963fbd, {16'd48028, 16'd64253, 16'd39480, 16'd57856, 16'd14651, 16'd47205, 16'd15101, 16'd25257, 16'd11514, 16'd37455, 16'd43605, 16'd58220, 16'd17593, 16'd2310, 16'd45902, 16'd30978, 16'd28014, 16'd476, 16'd64295, 16'd58035, 16'd19412, 16'd2627, 16'd13159, 16'd3847, 16'd42436, 16'd64748});
	test_expansion(128'h03e5135e1af7ff246fd9790464f9d25e, {16'd3073, 16'd24522, 16'd12340, 16'd6809, 16'd35841, 16'd42221, 16'd39514, 16'd29910, 16'd34750, 16'd39973, 16'd15607, 16'd36301, 16'd1861, 16'd27461, 16'd39808, 16'd36854, 16'd50063, 16'd30754, 16'd42207, 16'd3284, 16'd4181, 16'd25938, 16'd30166, 16'd3110, 16'd39952, 16'd7103});
	test_expansion(128'ha50cc64232da80d2daed9dcdce3536b7, {16'd43437, 16'd57359, 16'd56887, 16'd64198, 16'd44165, 16'd50994, 16'd37658, 16'd9454, 16'd18747, 16'd40277, 16'd20633, 16'd1134, 16'd36519, 16'd1143, 16'd22444, 16'd44280, 16'd52698, 16'd450, 16'd6298, 16'd58880, 16'd57339, 16'd49878, 16'd1195, 16'd37232, 16'd30112, 16'd47758});
	test_expansion(128'h9d6fd8e976f9b7660a484b421ac4c3ce, {16'd11521, 16'd9145, 16'd39363, 16'd39197, 16'd12336, 16'd40895, 16'd2636, 16'd32108, 16'd60850, 16'd58420, 16'd59642, 16'd15675, 16'd41324, 16'd18807, 16'd16754, 16'd24925, 16'd44254, 16'd12807, 16'd34069, 16'd55177, 16'd42901, 16'd54139, 16'd714, 16'd33439, 16'd64294, 16'd49541});
	test_expansion(128'h16d2bb5e24d6c170a69675b53f2f49f1, {16'd11799, 16'd10785, 16'd24638, 16'd46856, 16'd2839, 16'd58393, 16'd51052, 16'd20053, 16'd49763, 16'd9339, 16'd62009, 16'd32826, 16'd17602, 16'd31913, 16'd43456, 16'd7534, 16'd11677, 16'd48956, 16'd42626, 16'd25363, 16'd23640, 16'd37849, 16'd25839, 16'd27967, 16'd40877, 16'd19681});
	test_expansion(128'h3dd30772943a3334cfc6ed944fa7c13a, {16'd22134, 16'd30333, 16'd62092, 16'd49365, 16'd7429, 16'd32064, 16'd38143, 16'd51645, 16'd26770, 16'd62136, 16'd40580, 16'd25255, 16'd1121, 16'd52416, 16'd8949, 16'd1763, 16'd56252, 16'd15812, 16'd54591, 16'd52656, 16'd12470, 16'd14600, 16'd51907, 16'd19081, 16'd59728, 16'd57872});
	test_expansion(128'h75bddf8ec64dbc4ae495b1e897413a31, {16'd15920, 16'd30269, 16'd56282, 16'd46963, 16'd1113, 16'd3406, 16'd35953, 16'd12060, 16'd55390, 16'd43371, 16'd46287, 16'd828, 16'd52972, 16'd11749, 16'd51817, 16'd3153, 16'd29893, 16'd28211, 16'd13430, 16'd46334, 16'd22565, 16'd44592, 16'd11704, 16'd51078, 16'd3304, 16'd2528});
	test_expansion(128'hda8e48d6d9691a51a4f2a032ddb6e8b2, {16'd26259, 16'd31629, 16'd47443, 16'd35791, 16'd19847, 16'd12279, 16'd55467, 16'd22210, 16'd34090, 16'd16253, 16'd14725, 16'd33326, 16'd33467, 16'd20900, 16'd22565, 16'd20152, 16'd17863, 16'd22114, 16'd28299, 16'd9202, 16'd36643, 16'd59340, 16'd33951, 16'd58481, 16'd49515, 16'd6436});
	test_expansion(128'h0420faef92244ae246962854560ec404, {16'd41867, 16'd17944, 16'd22923, 16'd47722, 16'd58193, 16'd31842, 16'd37640, 16'd31849, 16'd44931, 16'd29229, 16'd1711, 16'd65192, 16'd27455, 16'd7822, 16'd26239, 16'd1976, 16'd7287, 16'd20127, 16'd16713, 16'd55407, 16'd61908, 16'd1106, 16'd7957, 16'd55627, 16'd54266, 16'd63292});
	test_expansion(128'h14e59d82ded41e22327bb57d78582020, {16'd63607, 16'd233, 16'd36341, 16'd2109, 16'd25725, 16'd3155, 16'd39198, 16'd36499, 16'd704, 16'd20563, 16'd4433, 16'd57171, 16'd39862, 16'd38193, 16'd37447, 16'd39644, 16'd58683, 16'd6717, 16'd39125, 16'd45013, 16'd2784, 16'd52989, 16'd49055, 16'd10278, 16'd37223, 16'd15221});
	test_expansion(128'hae568bbd7f56f00a9525e765d886638b, {16'd32356, 16'd16917, 16'd19758, 16'd49598, 16'd53495, 16'd5569, 16'd49803, 16'd45348, 16'd18068, 16'd40136, 16'd52588, 16'd13019, 16'd16945, 16'd4992, 16'd24761, 16'd56293, 16'd49052, 16'd52915, 16'd7021, 16'd43676, 16'd58327, 16'd47807, 16'd21697, 16'd41463, 16'd22099, 16'd42721});
	test_expansion(128'h14784d9e349ecd78820cbc0250ad254a, {16'd32572, 16'd45281, 16'd47853, 16'd8540, 16'd34345, 16'd60298, 16'd56996, 16'd54412, 16'd25265, 16'd31603, 16'd57814, 16'd44596, 16'd7902, 16'd37525, 16'd58085, 16'd34182, 16'd6, 16'd3621, 16'd42268, 16'd17072, 16'd40624, 16'd61097, 16'd35642, 16'd43359, 16'd26344, 16'd27278});
	test_expansion(128'h7dc53cc2e0f301e302e89237fe0598f8, {16'd58765, 16'd33645, 16'd19087, 16'd39015, 16'd36498, 16'd60163, 16'd25036, 16'd37229, 16'd43599, 16'd36005, 16'd10717, 16'd40948, 16'd49813, 16'd61250, 16'd21941, 16'd55824, 16'd17757, 16'd21679, 16'd15824, 16'd37207, 16'd52976, 16'd10688, 16'd27369, 16'd1656, 16'd36747, 16'd27570});
	test_expansion(128'hcda6c11fbf88b21742525a7e6bc40fcc, {16'd2357, 16'd34402, 16'd46447, 16'd31635, 16'd28182, 16'd29799, 16'd17892, 16'd50530, 16'd30685, 16'd57508, 16'd20225, 16'd62010, 16'd22190, 16'd47163, 16'd33263, 16'd5375, 16'd20172, 16'd11301, 16'd34602, 16'd54825, 16'd55601, 16'd54433, 16'd34201, 16'd16750, 16'd48506, 16'd12550});
	test_expansion(128'h2ffe4a760a0c82a77da8d4beef1bfbd6, {16'd1784, 16'd45958, 16'd60176, 16'd60106, 16'd65493, 16'd63606, 16'd58276, 16'd8997, 16'd14827, 16'd38847, 16'd49432, 16'd40002, 16'd23887, 16'd24284, 16'd36936, 16'd1762, 16'd16926, 16'd19540, 16'd46656, 16'd37497, 16'd17648, 16'd51726, 16'd52804, 16'd27620, 16'd56844, 16'd28095});
	test_expansion(128'hf5a6472817a89231bac385f3a6a12ca5, {16'd23236, 16'd57262, 16'd64912, 16'd33019, 16'd31446, 16'd34702, 16'd6644, 16'd863, 16'd35346, 16'd61257, 16'd53656, 16'd2683, 16'd48547, 16'd54964, 16'd28420, 16'd62205, 16'd33787, 16'd35975, 16'd31100, 16'd42052, 16'd255, 16'd46827, 16'd7057, 16'd14725, 16'd15724, 16'd42434});
	test_expansion(128'h488195f2f50760e75ed50080c4add3da, {16'd3723, 16'd51173, 16'd41691, 16'd46148, 16'd56317, 16'd2999, 16'd53639, 16'd33231, 16'd54170, 16'd24590, 16'd54551, 16'd32230, 16'd25687, 16'd19737, 16'd39587, 16'd23581, 16'd7239, 16'd45688, 16'd47990, 16'd62062, 16'd60278, 16'd15587, 16'd7610, 16'd25484, 16'd46645, 16'd42026});
	test_expansion(128'h4fa36d58cae992d09d8827773ae7943a, {16'd6982, 16'd38188, 16'd3250, 16'd53340, 16'd11971, 16'd13699, 16'd1850, 16'd4778, 16'd38631, 16'd33067, 16'd38602, 16'd23782, 16'd28887, 16'd51458, 16'd17313, 16'd29876, 16'd7695, 16'd15978, 16'd57068, 16'd64626, 16'd1657, 16'd24141, 16'd38987, 16'd38385, 16'd34571, 16'd8354});
	test_expansion(128'hc843d5d6c71b08e59f0ce7793eeeafe8, {16'd15168, 16'd41502, 16'd60153, 16'd39478, 16'd35903, 16'd45858, 16'd35423, 16'd30980, 16'd13682, 16'd47453, 16'd3198, 16'd40425, 16'd34655, 16'd58980, 16'd50897, 16'd60138, 16'd26997, 16'd35943, 16'd42273, 16'd46902, 16'd40177, 16'd8041, 16'd60806, 16'd2727, 16'd43280, 16'd34908});
	test_expansion(128'h94187d0bc39924c98a54b7f38bb9fb93, {16'd1979, 16'd16036, 16'd54199, 16'd59116, 16'd40827, 16'd56222, 16'd6540, 16'd1112, 16'd22543, 16'd33184, 16'd18648, 16'd4837, 16'd1469, 16'd30435, 16'd21207, 16'd20204, 16'd3356, 16'd22354, 16'd19161, 16'd35361, 16'd51211, 16'd60590, 16'd7032, 16'd35486, 16'd60909, 16'd52710});
	test_expansion(128'h9ede1eea7971e58be50af177c132b787, {16'd42032, 16'd16865, 16'd1551, 16'd48460, 16'd16393, 16'd2669, 16'd29694, 16'd55153, 16'd51088, 16'd12601, 16'd23937, 16'd36082, 16'd559, 16'd47614, 16'd21784, 16'd36970, 16'd44197, 16'd1204, 16'd46510, 16'd37639, 16'd3215, 16'd43634, 16'd26286, 16'd1277, 16'd38633, 16'd31260});
	test_expansion(128'h38814db08df6ed8b9c7477da5dd5e578, {16'd2289, 16'd45776, 16'd24790, 16'd4869, 16'd57786, 16'd2932, 16'd54749, 16'd43648, 16'd30098, 16'd14149, 16'd26409, 16'd11322, 16'd54986, 16'd6518, 16'd15107, 16'd41545, 16'd18141, 16'd36928, 16'd14062, 16'd11476, 16'd64361, 16'd3772, 16'd27344, 16'd34456, 16'd33397, 16'd45006});
	test_expansion(128'h2e07a0bab66ca1adceafc09e5c4081d4, {16'd36754, 16'd47886, 16'd55067, 16'd31052, 16'd63330, 16'd19453, 16'd44418, 16'd28290, 16'd14922, 16'd21642, 16'd1824, 16'd29317, 16'd56417, 16'd56156, 16'd55531, 16'd63283, 16'd28981, 16'd24439, 16'd1375, 16'd26444, 16'd19371, 16'd8565, 16'd17877, 16'd20583, 16'd34449, 16'd32121});
	test_expansion(128'h21b75fb50945a76afa8091d27bdb5d2b, {16'd48137, 16'd2334, 16'd22005, 16'd43018, 16'd36786, 16'd14130, 16'd61654, 16'd26478, 16'd13657, 16'd56210, 16'd22054, 16'd17669, 16'd21763, 16'd28282, 16'd65100, 16'd16594, 16'd42191, 16'd17541, 16'd46466, 16'd25722, 16'd1948, 16'd9011, 16'd5675, 16'd20283, 16'd52796, 16'd11608});
	test_expansion(128'h98d8d226172b7f8bc16f4a9b62873a62, {16'd39556, 16'd56164, 16'd65328, 16'd42624, 16'd40818, 16'd50575, 16'd7559, 16'd37036, 16'd27793, 16'd40505, 16'd53465, 16'd34498, 16'd46644, 16'd53653, 16'd11917, 16'd3816, 16'd57677, 16'd2330, 16'd291, 16'd56536, 16'd37455, 16'd15304, 16'd14850, 16'd5221, 16'd11656, 16'd53409});
	test_expansion(128'h093c0271009785b3872a84cc3a66f9ea, {16'd32452, 16'd14359, 16'd16862, 16'd15073, 16'd46662, 16'd54900, 16'd37351, 16'd18768, 16'd35500, 16'd37349, 16'd30994, 16'd60400, 16'd7451, 16'd21665, 16'd46943, 16'd57967, 16'd24451, 16'd42305, 16'd23719, 16'd11464, 16'd18336, 16'd9193, 16'd47133, 16'd829, 16'd11511, 16'd13752});
	test_expansion(128'h123ab0e625463217d403315e53db799a, {16'd41655, 16'd14863, 16'd11442, 16'd58056, 16'd23951, 16'd43230, 16'd33659, 16'd27406, 16'd31803, 16'd54816, 16'd49057, 16'd41399, 16'd50806, 16'd57173, 16'd4743, 16'd14545, 16'd16172, 16'd23723, 16'd51676, 16'd23095, 16'd28004, 16'd22957, 16'd49357, 16'd49312, 16'd14157, 16'd3231});
	test_expansion(128'h73c82ae69382fcef9759d71e49038f7d, {16'd34347, 16'd33031, 16'd14383, 16'd34093, 16'd2057, 16'd53326, 16'd64774, 16'd45923, 16'd27216, 16'd34020, 16'd51503, 16'd35138, 16'd6317, 16'd61663, 16'd34178, 16'd39359, 16'd15639, 16'd9274, 16'd30270, 16'd6714, 16'd15907, 16'd29616, 16'd34300, 16'd47319, 16'd10245, 16'd54934});
	test_expansion(128'hcbf7fa08aa54ea9864551bb1c83aa094, {16'd9493, 16'd19865, 16'd57179, 16'd20784, 16'd51398, 16'd10686, 16'd5823, 16'd51165, 16'd50530, 16'd21309, 16'd13703, 16'd15530, 16'd49208, 16'd63303, 16'd58190, 16'd16806, 16'd62320, 16'd15660, 16'd2750, 16'd34780, 16'd54733, 16'd5675, 16'd48006, 16'd21653, 16'd8350, 16'd60470});
	test_expansion(128'h28031e978113fe24ca46f89fedc00221, {16'd22783, 16'd32173, 16'd15460, 16'd28859, 16'd12668, 16'd47729, 16'd18783, 16'd55870, 16'd11689, 16'd36992, 16'd51105, 16'd61340, 16'd41941, 16'd37825, 16'd33546, 16'd39650, 16'd42999, 16'd50643, 16'd27087, 16'd12525, 16'd55871, 16'd18912, 16'd18895, 16'd22396, 16'd52986, 16'd35019});
	test_expansion(128'h48d703ec2f4290dcf23fae6b362b804d, {16'd33695, 16'd63726, 16'd18517, 16'd31156, 16'd4471, 16'd38212, 16'd64216, 16'd13870, 16'd50397, 16'd44176, 16'd21876, 16'd60619, 16'd38388, 16'd18801, 16'd27674, 16'd24643, 16'd41879, 16'd41194, 16'd20380, 16'd33182, 16'd49524, 16'd48373, 16'd54116, 16'd5906, 16'd61215, 16'd50934});
	test_expansion(128'hbc675b87af2da6fe451d551df552d35d, {16'd37459, 16'd46115, 16'd30710, 16'd18343, 16'd25946, 16'd33902, 16'd32065, 16'd11727, 16'd4302, 16'd17840, 16'd41954, 16'd4733, 16'd48612, 16'd2784, 16'd5074, 16'd57718, 16'd7979, 16'd55503, 16'd31905, 16'd35703, 16'd16541, 16'd9144, 16'd7571, 16'd42957, 16'd24227, 16'd666});
	test_expansion(128'hef2dac040acf822ed33bff2d8f23690a, {16'd11764, 16'd62415, 16'd59665, 16'd62466, 16'd35092, 16'd62917, 16'd10839, 16'd53344, 16'd4949, 16'd34022, 16'd12825, 16'd59537, 16'd3871, 16'd24982, 16'd41310, 16'd17598, 16'd41910, 16'd11673, 16'd12762, 16'd45860, 16'd55226, 16'd48934, 16'd28057, 16'd38199, 16'd32181, 16'd14039});
	test_expansion(128'h9f4e222340327b0d7e07cc4e07162cde, {16'd64991, 16'd64189, 16'd43002, 16'd44999, 16'd11259, 16'd42346, 16'd5224, 16'd24296, 16'd44672, 16'd36886, 16'd25017, 16'd34069, 16'd51170, 16'd42096, 16'd18653, 16'd61109, 16'd23315, 16'd48138, 16'd29500, 16'd29637, 16'd12378, 16'd4081, 16'd25063, 16'd40813, 16'd40439, 16'd15926});
	test_expansion(128'hef5a341e73b869d1f4097eca635b402d, {16'd56590, 16'd30373, 16'd11033, 16'd15760, 16'd28937, 16'd59325, 16'd52683, 16'd29451, 16'd21834, 16'd16027, 16'd47957, 16'd55400, 16'd54104, 16'd63833, 16'd2589, 16'd29313, 16'd30576, 16'd45112, 16'd27515, 16'd55577, 16'd48870, 16'd2783, 16'd23829, 16'd57593, 16'd37398, 16'd49390});
	test_expansion(128'hfeb0070d2fd82a18973ef4976a37137b, {16'd17731, 16'd59246, 16'd63010, 16'd29296, 16'd50916, 16'd9526, 16'd55989, 16'd12326, 16'd5897, 16'd62870, 16'd59979, 16'd30664, 16'd26692, 16'd48186, 16'd52867, 16'd52736, 16'd3090, 16'd45913, 16'd11755, 16'd44542, 16'd12269, 16'd59279, 16'd35931, 16'd43936, 16'd30332, 16'd17761});
	test_expansion(128'h3badb9a1f04efb4074484fa8d8fc5d95, {16'd3126, 16'd8669, 16'd39948, 16'd1762, 16'd6966, 16'd5013, 16'd18797, 16'd33741, 16'd18045, 16'd46082, 16'd60820, 16'd34205, 16'd8609, 16'd64907, 16'd5329, 16'd26155, 16'd44517, 16'd1250, 16'd48703, 16'd33111, 16'd13509, 16'd33313, 16'd11339, 16'd34646, 16'd42482, 16'd12808});
	test_expansion(128'he0dc8ec9fabd05aa6e77fe14a03e7df3, {16'd54163, 16'd8330, 16'd56895, 16'd18670, 16'd34272, 16'd3330, 16'd42234, 16'd39596, 16'd54599, 16'd54311, 16'd48568, 16'd47003, 16'd28138, 16'd40704, 16'd59913, 16'd1802, 16'd29650, 16'd6271, 16'd4436, 16'd15939, 16'd2870, 16'd35244, 16'd40050, 16'd15704, 16'd51993, 16'd50069});
	test_expansion(128'h832561e52f6a637dd48c7333423feb18, {16'd4860, 16'd63618, 16'd17525, 16'd51107, 16'd8465, 16'd1921, 16'd52986, 16'd1830, 16'd61546, 16'd61041, 16'd1093, 16'd54089, 16'd26294, 16'd64187, 16'd44090, 16'd51881, 16'd44634, 16'd19930, 16'd38023, 16'd14141, 16'd10358, 16'd9620, 16'd55992, 16'd5679, 16'd26491, 16'd22871});
	test_expansion(128'h2e3e9ab4a90eebc0795d0be6d99cccd0, {16'd27198, 16'd47984, 16'd50417, 16'd20229, 16'd11867, 16'd1948, 16'd61075, 16'd31742, 16'd17167, 16'd53134, 16'd8997, 16'd28676, 16'd33420, 16'd31551, 16'd61065, 16'd34330, 16'd27033, 16'd49857, 16'd45891, 16'd24993, 16'd3479, 16'd23083, 16'd29887, 16'd63430, 16'd55860, 16'd28800});
	test_expansion(128'h97b9a085a780a4183de83bbd3f9eeee0, {16'd46487, 16'd3136, 16'd28643, 16'd65093, 16'd50352, 16'd39226, 16'd31828, 16'd16308, 16'd38424, 16'd41260, 16'd24912, 16'd7736, 16'd65114, 16'd19552, 16'd52151, 16'd53421, 16'd29833, 16'd53872, 16'd53287, 16'd26695, 16'd35654, 16'd34275, 16'd15616, 16'd17813, 16'd19952, 16'd9658});
	test_expansion(128'hd71b30009cc583deece9efbc0eb49521, {16'd62578, 16'd337, 16'd20622, 16'd42780, 16'd43468, 16'd62111, 16'd42573, 16'd53997, 16'd12453, 16'd14364, 16'd51291, 16'd12612, 16'd64124, 16'd21138, 16'd17614, 16'd36032, 16'd2179, 16'd58499, 16'd20238, 16'd50576, 16'd43883, 16'd39854, 16'd11201, 16'd25481, 16'd51448, 16'd14353});
	test_expansion(128'h9424619283cc5ac2c69f3da310143702, {16'd17278, 16'd25662, 16'd40787, 16'd20125, 16'd15922, 16'd26310, 16'd42941, 16'd23703, 16'd65188, 16'd19507, 16'd21575, 16'd30074, 16'd4831, 16'd4422, 16'd405, 16'd35161, 16'd33576, 16'd54208, 16'd64027, 16'd9047, 16'd20354, 16'd44130, 16'd31767, 16'd64777, 16'd7656, 16'd50348});
	test_expansion(128'h77481b335cace897d287806490a6cb54, {16'd41417, 16'd18531, 16'd38262, 16'd25019, 16'd27450, 16'd40921, 16'd39772, 16'd13341, 16'd19070, 16'd52573, 16'd29522, 16'd39398, 16'd38378, 16'd51300, 16'd37210, 16'd13196, 16'd6061, 16'd27554, 16'd28703, 16'd39354, 16'd47695, 16'd57929, 16'd46457, 16'd629, 16'd36941, 16'd7459});
	test_expansion(128'h48b3b6087e2f1fd74effb214645a569f, {16'd47501, 16'd40957, 16'd10469, 16'd42825, 16'd39091, 16'd16899, 16'd39216, 16'd59652, 16'd40649, 16'd50418, 16'd52467, 16'd31618, 16'd15219, 16'd27226, 16'd22949, 16'd21088, 16'd34137, 16'd8465, 16'd40624, 16'd33078, 16'd30363, 16'd63983, 16'd30194, 16'd46653, 16'd52420, 16'd19373});
	test_expansion(128'haf454d1a691677dcbcd16794fec55cd8, {16'd51975, 16'd849, 16'd54979, 16'd6979, 16'd54367, 16'd43079, 16'd64914, 16'd24715, 16'd57994, 16'd60969, 16'd51037, 16'd40443, 16'd34201, 16'd50284, 16'd36515, 16'd19520, 16'd50947, 16'd38257, 16'd43074, 16'd55872, 16'd3201, 16'd13410, 16'd26752, 16'd43201, 16'd53589, 16'd35198});
	test_expansion(128'hcd8c828d460fa63906f6304a868218d0, {16'd20554, 16'd28936, 16'd44078, 16'd49434, 16'd33092, 16'd41330, 16'd55130, 16'd28384, 16'd29602, 16'd24009, 16'd11917, 16'd39983, 16'd58697, 16'd35000, 16'd53743, 16'd25418, 16'd13427, 16'd31720, 16'd28324, 16'd29556, 16'd19480, 16'd26654, 16'd20516, 16'd64027, 16'd37912, 16'd59471});
	test_expansion(128'h0d0b8abd2abc9045ccb7cc2ca6ad9b9b, {16'd48925, 16'd12203, 16'd33801, 16'd54633, 16'd26843, 16'd31062, 16'd59964, 16'd27886, 16'd52924, 16'd31062, 16'd62025, 16'd58934, 16'd44499, 16'd59281, 16'd22534, 16'd54180, 16'd62534, 16'd7608, 16'd44881, 16'd29145, 16'd3454, 16'd42003, 16'd415, 16'd35402, 16'd27999, 16'd63136});
	test_expansion(128'hffae7036047283c27d8c070b061c3a60, {16'd15858, 16'd58804, 16'd64640, 16'd23850, 16'd46317, 16'd50421, 16'd27513, 16'd31922, 16'd9116, 16'd45761, 16'd64534, 16'd57665, 16'd26749, 16'd58762, 16'd31849, 16'd11026, 16'd60934, 16'd7991, 16'd47547, 16'd55324, 16'd10963, 16'd48628, 16'd44133, 16'd62931, 16'd13136, 16'd60581});
	test_expansion(128'hd15da52603a2a0e517e555177e408a86, {16'd64676, 16'd472, 16'd57532, 16'd2951, 16'd32015, 16'd5529, 16'd6219, 16'd9955, 16'd3291, 16'd62609, 16'd18196, 16'd43989, 16'd34013, 16'd12141, 16'd37655, 16'd19589, 16'd3434, 16'd20995, 16'd15816, 16'd12756, 16'd57495, 16'd24981, 16'd13544, 16'd22646, 16'd23206, 16'd63241});
	test_expansion(128'hcabb2c82b5b7fd01f6342b735a4a2a6d, {16'd41366, 16'd32124, 16'd18898, 16'd7225, 16'd15389, 16'd33483, 16'd57699, 16'd11461, 16'd45960, 16'd32067, 16'd44081, 16'd59598, 16'd47366, 16'd40246, 16'd28996, 16'd31447, 16'd26634, 16'd14254, 16'd64167, 16'd23137, 16'd40972, 16'd24863, 16'd63451, 16'd20413, 16'd4538, 16'd3927});
	test_expansion(128'he509bb518eacf01e2f16fd812595864e, {16'd59574, 16'd19366, 16'd10232, 16'd62385, 16'd47403, 16'd35633, 16'd55543, 16'd54416, 16'd49960, 16'd35512, 16'd39983, 16'd46814, 16'd16457, 16'd20236, 16'd36049, 16'd27540, 16'd64165, 16'd46493, 16'd329, 16'd45535, 16'd63671, 16'd49042, 16'd8958, 16'd29101, 16'd29247, 16'd64401});
	test_expansion(128'hcc356c2621b79f0e86d31cbf6a6e605d, {16'd62266, 16'd52859, 16'd50301, 16'd39859, 16'd16707, 16'd43875, 16'd37256, 16'd18422, 16'd1846, 16'd34263, 16'd34445, 16'd60138, 16'd58096, 16'd11413, 16'd18838, 16'd63152, 16'd5201, 16'd19137, 16'd34649, 16'd46295, 16'd64929, 16'd63473, 16'd20075, 16'd33269, 16'd6829, 16'd7829});
	test_expansion(128'hb19c76e2551caa2cb8947fd5908d2eb9, {16'd21631, 16'd9812, 16'd18651, 16'd5701, 16'd10083, 16'd35628, 16'd19232, 16'd42635, 16'd14672, 16'd34673, 16'd36404, 16'd7382, 16'd17869, 16'd24217, 16'd48655, 16'd3607, 16'd62498, 16'd13074, 16'd15984, 16'd3408, 16'd52452, 16'd51907, 16'd6879, 16'd55178, 16'd16444, 16'd29322});
	test_expansion(128'hd4768abc77abe6f44c6ba69cef8a7f45, {16'd64124, 16'd65436, 16'd7415, 16'd45875, 16'd41846, 16'd45047, 16'd24776, 16'd13124, 16'd59123, 16'd7662, 16'd8224, 16'd7658, 16'd2791, 16'd44224, 16'd46231, 16'd45537, 16'd62960, 16'd41982, 16'd28791, 16'd15220, 16'd6494, 16'd31230, 16'd26114, 16'd29993, 16'd34177, 16'd34885});
	test_expansion(128'h7c61a50ffa4c6ed3a37c3a98becdeed2, {16'd59772, 16'd11339, 16'd58662, 16'd41114, 16'd44356, 16'd48020, 16'd11272, 16'd11615, 16'd43231, 16'd48726, 16'd59231, 16'd27993, 16'd18342, 16'd38986, 16'd35281, 16'd20213, 16'd46654, 16'd49960, 16'd55709, 16'd56435, 16'd8101, 16'd58408, 16'd55365, 16'd40966, 16'd55218, 16'd3230});
	test_expansion(128'hbd0cfc350c1028c0d1ebbcaed5a7d960, {16'd37558, 16'd18910, 16'd24057, 16'd4839, 16'd44944, 16'd40062, 16'd5099, 16'd44503, 16'd25051, 16'd33565, 16'd19572, 16'd27362, 16'd52024, 16'd5336, 16'd53554, 16'd9525, 16'd33407, 16'd24855, 16'd9842, 16'd33901, 16'd47030, 16'd60163, 16'd36656, 16'd52908, 16'd43013, 16'd40895});
	test_expansion(128'h12acf09108bd60e4528c0171b32dcbd9, {16'd23585, 16'd50208, 16'd16873, 16'd52664, 16'd46657, 16'd47963, 16'd12067, 16'd45811, 16'd54931, 16'd28953, 16'd57478, 16'd7819, 16'd56495, 16'd39931, 16'd41307, 16'd61383, 16'd3917, 16'd52033, 16'd21096, 16'd2844, 16'd3694, 16'd45517, 16'd41057, 16'd59121, 16'd7950, 16'd38963});
	test_expansion(128'hc71d659258c8753d953106b44d4e2bf4, {16'd17621, 16'd11853, 16'd9460, 16'd39979, 16'd56444, 16'd13528, 16'd15157, 16'd40209, 16'd62488, 16'd37220, 16'd21885, 16'd45623, 16'd14032, 16'd11139, 16'd53885, 16'd50262, 16'd37362, 16'd52807, 16'd33998, 16'd58447, 16'd12872, 16'd23300, 16'd59984, 16'd64427, 16'd13526, 16'd15559});
	test_expansion(128'he635834fa87024dcfe2c41aa37091b5a, {16'd14912, 16'd50002, 16'd37385, 16'd34982, 16'd35582, 16'd61293, 16'd29975, 16'd64670, 16'd31509, 16'd11412, 16'd7712, 16'd41248, 16'd16511, 16'd1098, 16'd25770, 16'd17257, 16'd30693, 16'd32193, 16'd57298, 16'd49153, 16'd60097, 16'd54639, 16'd25227, 16'd41829, 16'd34875, 16'd59455});
	test_expansion(128'h2675194e0347633ac9d73dfb2b1a7d6d, {16'd38303, 16'd48625, 16'd56664, 16'd51058, 16'd11349, 16'd12657, 16'd56127, 16'd11629, 16'd43461, 16'd50718, 16'd32180, 16'd14482, 16'd48040, 16'd40754, 16'd62570, 16'd24498, 16'd10737, 16'd20863, 16'd23267, 16'd42705, 16'd62649, 16'd63203, 16'd11775, 16'd26963, 16'd37900, 16'd17715});
	test_expansion(128'ha812e334740443b4bbacd7ef7e957343, {16'd34449, 16'd23521, 16'd47152, 16'd51753, 16'd40938, 16'd27252, 16'd32069, 16'd62028, 16'd45389, 16'd59352, 16'd50, 16'd31924, 16'd52306, 16'd19740, 16'd46868, 16'd6285, 16'd16407, 16'd53520, 16'd61325, 16'd23535, 16'd28058, 16'd49444, 16'd36961, 16'd56391, 16'd47659, 16'd56263});
	test_expansion(128'ha6875e13d61374423752c5cfbfa915b2, {16'd53611, 16'd37723, 16'd25202, 16'd48889, 16'd12054, 16'd37934, 16'd34419, 16'd33610, 16'd18802, 16'd1705, 16'd7174, 16'd45190, 16'd29069, 16'd13587, 16'd19002, 16'd60125, 16'd15619, 16'd19866, 16'd28212, 16'd21065, 16'd58706, 16'd49187, 16'd2964, 16'd17159, 16'd12928, 16'd6277});
	test_expansion(128'hb8b5c1a137f478ddfc1deb0f7144304f, {16'd26425, 16'd37965, 16'd63341, 16'd51908, 16'd4873, 16'd26940, 16'd43208, 16'd55022, 16'd19035, 16'd52861, 16'd4272, 16'd33982, 16'd55622, 16'd54888, 16'd58111, 16'd18543, 16'd18510, 16'd46655, 16'd20140, 16'd6755, 16'd21157, 16'd15171, 16'd63888, 16'd32575, 16'd12859, 16'd4841});
	test_expansion(128'h3cafc189bc6caf8a9894cd372a021d03, {16'd30737, 16'd64771, 16'd20652, 16'd41654, 16'd9577, 16'd17908, 16'd40560, 16'd29576, 16'd64158, 16'd38767, 16'd58913, 16'd10594, 16'd29237, 16'd23866, 16'd45740, 16'd50716, 16'd10177, 16'd41399, 16'd34480, 16'd1069, 16'd44569, 16'd26964, 16'd56246, 16'd9961, 16'd54787, 16'd9138});
	test_expansion(128'h8212301ec3b6a6c4a64ef424fe40029b, {16'd43620, 16'd31498, 16'd14910, 16'd54432, 16'd20937, 16'd10430, 16'd27256, 16'd39525, 16'd7225, 16'd30143, 16'd59131, 16'd23613, 16'd23662, 16'd26576, 16'd36508, 16'd2211, 16'd54362, 16'd46734, 16'd8025, 16'd14158, 16'd60243, 16'd27395, 16'd59223, 16'd21534, 16'd34641, 16'd43449});
	test_expansion(128'h2b696a07fa77ea1e76c095b70f5d2799, {16'd21654, 16'd43479, 16'd19076, 16'd6851, 16'd6646, 16'd19829, 16'd17015, 16'd40066, 16'd51043, 16'd43622, 16'd60178, 16'd4150, 16'd14507, 16'd52789, 16'd31853, 16'd30327, 16'd24652, 16'd1163, 16'd7985, 16'd4493, 16'd50177, 16'd31531, 16'd37723, 16'd17989, 16'd47550, 16'd45085});
	test_expansion(128'h91faba430fb27396195ff8208ef01c44, {16'd1289, 16'd21038, 16'd39122, 16'd55432, 16'd63396, 16'd40620, 16'd36043, 16'd31212, 16'd9839, 16'd5753, 16'd56422, 16'd18818, 16'd1630, 16'd22923, 16'd21389, 16'd16530, 16'd46768, 16'd44748, 16'd64643, 16'd49658, 16'd17668, 16'd7799, 16'd4857, 16'd49868, 16'd13733, 16'd51473});
	test_expansion(128'hb8af3256fa2b3633c8387a99ee02ec25, {16'd52387, 16'd46760, 16'd28251, 16'd4630, 16'd58723, 16'd64923, 16'd22883, 16'd64886, 16'd10094, 16'd39063, 16'd25996, 16'd47651, 16'd44581, 16'd62403, 16'd38829, 16'd65401, 16'd14173, 16'd28709, 16'd19369, 16'd34041, 16'd57477, 16'd54104, 16'd61922, 16'd24805, 16'd57025, 16'd54944});
	test_expansion(128'h2a12ca45b805f589476fe9969c8a5912, {16'd48248, 16'd60862, 16'd17941, 16'd1977, 16'd53215, 16'd11830, 16'd25296, 16'd12287, 16'd41210, 16'd14705, 16'd55544, 16'd35271, 16'd36558, 16'd42733, 16'd46958, 16'd29119, 16'd9484, 16'd46162, 16'd20096, 16'd28226, 16'd457, 16'd62026, 16'd14677, 16'd2385, 16'd48958, 16'd17157});
	test_expansion(128'h52a9462c9939e6f51d6d7eee0b0e33dd, {16'd24658, 16'd30075, 16'd21532, 16'd40129, 16'd31579, 16'd33452, 16'd28015, 16'd16579, 16'd59072, 16'd761, 16'd5598, 16'd17014, 16'd34575, 16'd28718, 16'd9674, 16'd9926, 16'd58031, 16'd15649, 16'd54039, 16'd28458, 16'd62982, 16'd26639, 16'd62609, 16'd41833, 16'd55024, 16'd47732});
	test_expansion(128'he5fb7a8da52b5f0dc0c93b5b935da6fb, {16'd799, 16'd9171, 16'd19250, 16'd12096, 16'd51751, 16'd64023, 16'd40934, 16'd13212, 16'd28141, 16'd13017, 16'd58896, 16'd41212, 16'd13369, 16'd7609, 16'd22492, 16'd33299, 16'd25498, 16'd55716, 16'd13521, 16'd23487, 16'd6129, 16'd41770, 16'd9282, 16'd3212, 16'd55859, 16'd3021});
	test_expansion(128'hb884bf591737dae18e22a109acc70f99, {16'd40145, 16'd56002, 16'd62956, 16'd22145, 16'd49181, 16'd21409, 16'd37843, 16'd25854, 16'd27586, 16'd55938, 16'd15802, 16'd57792, 16'd4327, 16'd56158, 16'd17759, 16'd46895, 16'd8457, 16'd48006, 16'd425, 16'd25293, 16'd4690, 16'd62407, 16'd48143, 16'd36511, 16'd11280, 16'd63292});
	test_expansion(128'h0fbd1e77ac13081d846d0fe9cf08fe89, {16'd31060, 16'd59739, 16'd60304, 16'd18245, 16'd22357, 16'd12065, 16'd26830, 16'd2170, 16'd61460, 16'd26679, 16'd14953, 16'd32424, 16'd8150, 16'd51983, 16'd50188, 16'd6985, 16'd36568, 16'd47249, 16'd57752, 16'd28251, 16'd37112, 16'd55615, 16'd42621, 16'd41682, 16'd36730, 16'd16818});
	test_expansion(128'h8a0c50c427d63417652da872996494e5, {16'd53582, 16'd4310, 16'd873, 16'd36749, 16'd49797, 16'd24426, 16'd65308, 16'd5468, 16'd55761, 16'd64733, 16'd58680, 16'd7272, 16'd3610, 16'd10635, 16'd20519, 16'd35317, 16'd53349, 16'd50848, 16'd40990, 16'd10042, 16'd22531, 16'd36977, 16'd8657, 16'd12267, 16'd7857, 16'd27864});
	test_expansion(128'heafeca2bf1fdabf09ff3656f2a084f03, {16'd63146, 16'd46790, 16'd43776, 16'd22596, 16'd61132, 16'd42171, 16'd31442, 16'd52695, 16'd8590, 16'd60674, 16'd4702, 16'd5207, 16'd17538, 16'd50108, 16'd2064, 16'd48414, 16'd34110, 16'd11939, 16'd3640, 16'd21766, 16'd44129, 16'd9028, 16'd6463, 16'd13093, 16'd63018, 16'd42792});
	test_expansion(128'h49a063eacfd9d8989b33d52feca44939, {16'd14650, 16'd19255, 16'd2715, 16'd25262, 16'd14148, 16'd40760, 16'd56613, 16'd27221, 16'd3230, 16'd51338, 16'd44047, 16'd47373, 16'd814, 16'd30098, 16'd27235, 16'd42105, 16'd33834, 16'd25654, 16'd43903, 16'd20695, 16'd44256, 16'd2683, 16'd14577, 16'd28553, 16'd50663, 16'd50308});
	test_expansion(128'hceab6618693f33606605065eba24fc04, {16'd11894, 16'd42251, 16'd8783, 16'd18797, 16'd50537, 16'd20561, 16'd55639, 16'd48527, 16'd59513, 16'd58833, 16'd28351, 16'd61871, 16'd29242, 16'd26158, 16'd44278, 16'd3306, 16'd32332, 16'd36209, 16'd18137, 16'd59802, 16'd37675, 16'd25021, 16'd43948, 16'd63954, 16'd32871, 16'd16082});
	test_expansion(128'h1cb20210e2e249739e5e778408464da4, {16'd27098, 16'd48044, 16'd43437, 16'd41683, 16'd24902, 16'd34430, 16'd33126, 16'd40281, 16'd60600, 16'd40366, 16'd28116, 16'd23398, 16'd54893, 16'd6123, 16'd16984, 16'd16919, 16'd49231, 16'd56659, 16'd53713, 16'd54331, 16'd30903, 16'd40760, 16'd7916, 16'd4816, 16'd7667, 16'd63467});
	test_expansion(128'h1b54c490dd300f87f569c3834f561468, {16'd61750, 16'd37402, 16'd15284, 16'd34190, 16'd391, 16'd27814, 16'd45623, 16'd25756, 16'd43586, 16'd21503, 16'd5387, 16'd59302, 16'd64882, 16'd37895, 16'd58365, 16'd48980, 16'd45882, 16'd7624, 16'd41, 16'd614, 16'd53435, 16'd22125, 16'd40551, 16'd49209, 16'd33838, 16'd32083});
	test_expansion(128'hb5f4c851789565fad336fc209615b670, {16'd61348, 16'd23067, 16'd41250, 16'd33890, 16'd1656, 16'd23208, 16'd33701, 16'd24695, 16'd35620, 16'd31771, 16'd58444, 16'd37225, 16'd53190, 16'd39801, 16'd50070, 16'd18884, 16'd12243, 16'd7776, 16'd39835, 16'd22291, 16'd15514, 16'd36910, 16'd64981, 16'd2651, 16'd51961, 16'd61931});
	test_expansion(128'hade74a682d02bf36aab2eb7d746a8f93, {16'd18970, 16'd20026, 16'd50308, 16'd2634, 16'd46778, 16'd34051, 16'd50146, 16'd21693, 16'd17685, 16'd48949, 16'd35165, 16'd65082, 16'd58552, 16'd19963, 16'd19789, 16'd2395, 16'd56472, 16'd26055, 16'd12905, 16'd39790, 16'd60527, 16'd5886, 16'd22393, 16'd27142, 16'd27300, 16'd7563});
	test_expansion(128'h48e1fa0afc536f2844cc91bc222a4032, {16'd8230, 16'd60450, 16'd40332, 16'd13037, 16'd40978, 16'd29021, 16'd42263, 16'd13428, 16'd53265, 16'd32907, 16'd41737, 16'd63434, 16'd65061, 16'd8212, 16'd54664, 16'd50555, 16'd11286, 16'd24646, 16'd30878, 16'd45150, 16'd57171, 16'd33579, 16'd62413, 16'd23981, 16'd6868, 16'd25092});
	test_expansion(128'h581a4666479936463f268558a45abfbc, {16'd50786, 16'd55848, 16'd2020, 16'd43658, 16'd49171, 16'd30973, 16'd51234, 16'd38007, 16'd43344, 16'd38328, 16'd17908, 16'd2557, 16'd33110, 16'd35608, 16'd61697, 16'd23479, 16'd64684, 16'd61113, 16'd56343, 16'd31396, 16'd34021, 16'd50486, 16'd48879, 16'd10576, 16'd6219, 16'd33352});
	test_expansion(128'h69980d78b7d6b6ae9b56fcec709678fe, {16'd43054, 16'd15488, 16'd14910, 16'd15092, 16'd28545, 16'd37219, 16'd16060, 16'd27942, 16'd39992, 16'd12158, 16'd16970, 16'd21506, 16'd40444, 16'd33652, 16'd18511, 16'd48471, 16'd4927, 16'd11159, 16'd47911, 16'd41429, 16'd9911, 16'd31944, 16'd32414, 16'd37610, 16'd35544, 16'd45576});
	test_expansion(128'h6d5961db8f203d54690d10b88d039104, {16'd43871, 16'd57306, 16'd41729, 16'd33165, 16'd42966, 16'd41291, 16'd54290, 16'd61184, 16'd43269, 16'd11804, 16'd31351, 16'd22104, 16'd61586, 16'd55270, 16'd35412, 16'd28604, 16'd7333, 16'd57005, 16'd4803, 16'd93, 16'd50544, 16'd12813, 16'd38945, 16'd59135, 16'd38958, 16'd43694});
	test_expansion(128'hede7c4d059b6f8688976d676edb2f377, {16'd19346, 16'd17553, 16'd14434, 16'd23153, 16'd42213, 16'd13016, 16'd49151, 16'd15153, 16'd58066, 16'd51084, 16'd49580, 16'd16230, 16'd30650, 16'd17309, 16'd8584, 16'd43093, 16'd6994, 16'd23080, 16'd23166, 16'd47439, 16'd2406, 16'd10823, 16'd32335, 16'd24325, 16'd45554, 16'd45519});
	test_expansion(128'h5695a423c6215c990a139faabe9af18a, {16'd15701, 16'd43770, 16'd10938, 16'd41229, 16'd37974, 16'd17479, 16'd32527, 16'd53239, 16'd31838, 16'd23732, 16'd52890, 16'd15358, 16'd30181, 16'd62372, 16'd2196, 16'd2269, 16'd9040, 16'd15798, 16'd45473, 16'd58734, 16'd65289, 16'd61610, 16'd5902, 16'd103, 16'd45047, 16'd4216});
	test_expansion(128'hbc10cbf32f525487470ede75c870b684, {16'd35704, 16'd27653, 16'd15310, 16'd49971, 16'd22624, 16'd37083, 16'd4624, 16'd43286, 16'd64264, 16'd8515, 16'd26009, 16'd36362, 16'd32083, 16'd42349, 16'd63758, 16'd59649, 16'd42639, 16'd64944, 16'd35860, 16'd47487, 16'd54478, 16'd37262, 16'd32098, 16'd22274, 16'd11444, 16'd59759});
	test_expansion(128'h0f36b6ae48b0a8d135950d97d07a3ff1, {16'd16290, 16'd47040, 16'd34941, 16'd49538, 16'd58834, 16'd58095, 16'd11398, 16'd36735, 16'd11522, 16'd25110, 16'd47380, 16'd35999, 16'd50087, 16'd65220, 16'd46943, 16'd32185, 16'd29741, 16'd35650, 16'd29640, 16'd52111, 16'd50895, 16'd30645, 16'd65113, 16'd49989, 16'd27428, 16'd17635});
	test_expansion(128'h0f681212d4fb3392fc2a5b6309f622e6, {16'd60837, 16'd35235, 16'd16698, 16'd31932, 16'd5929, 16'd53439, 16'd54095, 16'd32081, 16'd18442, 16'd43776, 16'd52153, 16'd41097, 16'd7641, 16'd30650, 16'd29104, 16'd26593, 16'd30337, 16'd31195, 16'd18307, 16'd36886, 16'd52013, 16'd9717, 16'd35022, 16'd14089, 16'd52113, 16'd55504});
	test_expansion(128'h8035357668bbba4abe614b9151794e48, {16'd46546, 16'd29562, 16'd9299, 16'd1039, 16'd43951, 16'd20973, 16'd9193, 16'd62132, 16'd33147, 16'd45027, 16'd43032, 16'd33588, 16'd15571, 16'd60730, 16'd45474, 16'd52854, 16'd10718, 16'd41543, 16'd192, 16'd62810, 16'd48441, 16'd16109, 16'd64349, 16'd35022, 16'd11261, 16'd63337});
	test_expansion(128'h94bb1a58fe0ea46d6020af64e1c3b79e, {16'd40569, 16'd8087, 16'd46287, 16'd60429, 16'd46906, 16'd1263, 16'd11840, 16'd146, 16'd16188, 16'd61427, 16'd15445, 16'd57125, 16'd63745, 16'd1094, 16'd53458, 16'd25040, 16'd44996, 16'd17250, 16'd28242, 16'd9844, 16'd34382, 16'd40049, 16'd2789, 16'd39632, 16'd7240, 16'd58249});
	test_expansion(128'h302ac8af9a053d919e2276e96e21de71, {16'd5744, 16'd31447, 16'd26016, 16'd27009, 16'd21651, 16'd47679, 16'd43143, 16'd27035, 16'd16918, 16'd2595, 16'd446, 16'd30530, 16'd31293, 16'd61461, 16'd5070, 16'd19825, 16'd62854, 16'd14423, 16'd60199, 16'd20123, 16'd16575, 16'd40553, 16'd61086, 16'd44215, 16'd8379, 16'd60270});
	test_expansion(128'hd882984de1ea123ba5d552a5ba6e4ebd, {16'd54358, 16'd46850, 16'd48403, 16'd26688, 16'd11638, 16'd37715, 16'd15654, 16'd56157, 16'd33650, 16'd27143, 16'd10052, 16'd36113, 16'd2578, 16'd10473, 16'd18637, 16'd4830, 16'd30217, 16'd8227, 16'd35673, 16'd33365, 16'd60661, 16'd26126, 16'd41310, 16'd17587, 16'd38232, 16'd47609});
	test_expansion(128'h8f6a2c11e2bd74e70e3184f15082befb, {16'd41914, 16'd41753, 16'd34957, 16'd13443, 16'd53164, 16'd22584, 16'd58700, 16'd7143, 16'd32724, 16'd25284, 16'd51818, 16'd4705, 16'd52953, 16'd775, 16'd49661, 16'd18702, 16'd32009, 16'd40769, 16'd48722, 16'd42538, 16'd45026, 16'd11195, 16'd22888, 16'd18990, 16'd14201, 16'd23671});
	test_expansion(128'h6fdcd79e3a2d77ea315972c0602d3eb5, {16'd52716, 16'd41760, 16'd39204, 16'd64915, 16'd35065, 16'd35973, 16'd46558, 16'd36342, 16'd57104, 16'd22342, 16'd26139, 16'd7359, 16'd23975, 16'd45311, 16'd19125, 16'd13250, 16'd58398, 16'd60770, 16'd2645, 16'd44052, 16'd13817, 16'd52880, 16'd4524, 16'd13140, 16'd38346, 16'd1782});
	test_expansion(128'h2cc140e54a9c9e0668de870963dc8de1, {16'd38501, 16'd51886, 16'd33247, 16'd3801, 16'd37206, 16'd2345, 16'd37373, 16'd32280, 16'd2457, 16'd10674, 16'd7810, 16'd4706, 16'd41925, 16'd6436, 16'd11507, 16'd57450, 16'd45715, 16'd40315, 16'd63313, 16'd40467, 16'd43582, 16'd5277, 16'd47318, 16'd31102, 16'd19107, 16'd27850});
	test_expansion(128'h9fdc40966fa71deb74bdf26319c66c5e, {16'd50657, 16'd35254, 16'd60473, 16'd3551, 16'd17494, 16'd37185, 16'd42948, 16'd6975, 16'd48282, 16'd8481, 16'd54704, 16'd29881, 16'd58263, 16'd12063, 16'd3966, 16'd5015, 16'd11426, 16'd6078, 16'd1374, 16'd60383, 16'd20970, 16'd58532, 16'd43356, 16'd33896, 16'd4133, 16'd14140});
	test_expansion(128'h027d619d8fc95f0b96c28f0d7a3e4976, {16'd14727, 16'd27167, 16'd8794, 16'd61376, 16'd44137, 16'd31230, 16'd16016, 16'd62229, 16'd4185, 16'd28373, 16'd51075, 16'd10189, 16'd43867, 16'd3291, 16'd34754, 16'd7085, 16'd46450, 16'd58154, 16'd13374, 16'd12719, 16'd39139, 16'd6490, 16'd37913, 16'd1902, 16'd28132, 16'd58223});
	test_expansion(128'h7d176516b2504ab4a1364667a8e97609, {16'd13129, 16'd39818, 16'd65171, 16'd19435, 16'd36180, 16'd40969, 16'd33239, 16'd44047, 16'd49140, 16'd52884, 16'd4426, 16'd41189, 16'd32672, 16'd10710, 16'd12773, 16'd64136, 16'd33288, 16'd12307, 16'd19482, 16'd62992, 16'd63141, 16'd56177, 16'd38725, 16'd226, 16'd16757, 16'd48412});
	test_expansion(128'hbe00d6acf00007deb4c7cba9968a4dfc, {16'd33472, 16'd9848, 16'd40774, 16'd15025, 16'd37496, 16'd34302, 16'd27523, 16'd38267, 16'd57989, 16'd39739, 16'd22985, 16'd28998, 16'd36067, 16'd41735, 16'd33008, 16'd46759, 16'd52903, 16'd36156, 16'd6654, 16'd2562, 16'd57056, 16'd13595, 16'd6754, 16'd60368, 16'd61977, 16'd33804});
	test_expansion(128'h5a6b10a904da6fe86be21051957bd37a, {16'd42557, 16'd33803, 16'd39588, 16'd11109, 16'd3744, 16'd16045, 16'd21111, 16'd63294, 16'd22675, 16'd27926, 16'd5927, 16'd52373, 16'd8934, 16'd44191, 16'd21413, 16'd65073, 16'd32867, 16'd11463, 16'd29210, 16'd29567, 16'd44113, 16'd20362, 16'd7571, 16'd14349, 16'd61306, 16'd20895});
	test_expansion(128'he3d699d7fb15f14982b11b7a24c72bf6, {16'd3807, 16'd26407, 16'd10095, 16'd46816, 16'd9978, 16'd47356, 16'd61714, 16'd24737, 16'd24224, 16'd47184, 16'd62344, 16'd1815, 16'd33826, 16'd16150, 16'd40197, 16'd47031, 16'd41182, 16'd60103, 16'd1041, 16'd19597, 16'd38723, 16'd9744, 16'd51391, 16'd17932, 16'd26801, 16'd63202});
	test_expansion(128'hcdd5dc6779d949351f85132cd06bf9c4, {16'd47872, 16'd21408, 16'd27551, 16'd47845, 16'd56236, 16'd57536, 16'd28166, 16'd23952, 16'd54158, 16'd47701, 16'd37598, 16'd55706, 16'd34456, 16'd50643, 16'd21066, 16'd35027, 16'd1719, 16'd36434, 16'd13156, 16'd61860, 16'd17922, 16'd18034, 16'd44606, 16'd9514, 16'd23396, 16'd8629});
	test_expansion(128'h1526ebebcf2356a665e5a8affd91ffc9, {16'd17050, 16'd24492, 16'd11541, 16'd3292, 16'd34825, 16'd47760, 16'd18154, 16'd59819, 16'd16783, 16'd12358, 16'd61332, 16'd59456, 16'd33978, 16'd38839, 16'd15341, 16'd49482, 16'd11123, 16'd48897, 16'd38448, 16'd8656, 16'd28984, 16'd61728, 16'd58027, 16'd24319, 16'd60050, 16'd55112});
	test_expansion(128'h951a6c7b6ff8480618f5effcf636072e, {16'd10512, 16'd9895, 16'd47605, 16'd25483, 16'd11710, 16'd28902, 16'd28614, 16'd15112, 16'd33572, 16'd20559, 16'd35441, 16'd48660, 16'd27249, 16'd20758, 16'd12722, 16'd50755, 16'd8707, 16'd59605, 16'd19297, 16'd51332, 16'd55864, 16'd25736, 16'd19092, 16'd43884, 16'd33692, 16'd62926});
	test_expansion(128'h564470ee3d03919f2acdbde8b79ef844, {16'd60160, 16'd53177, 16'd54876, 16'd60808, 16'd10978, 16'd55883, 16'd45259, 16'd40033, 16'd64717, 16'd38596, 16'd38214, 16'd21678, 16'd45538, 16'd39149, 16'd37238, 16'd64722, 16'd42283, 16'd43528, 16'd8739, 16'd45619, 16'd38399, 16'd23200, 16'd18341, 16'd4134, 16'd32407, 16'd50384});
	test_expansion(128'hd00834d623817d21ad9ce652684558f7, {16'd45019, 16'd55227, 16'd8934, 16'd41404, 16'd61711, 16'd1313, 16'd33415, 16'd64811, 16'd7993, 16'd29826, 16'd24752, 16'd12343, 16'd3812, 16'd4454, 16'd5410, 16'd49172, 16'd55002, 16'd38751, 16'd52767, 16'd36315, 16'd43765, 16'd13401, 16'd9148, 16'd33, 16'd58817, 16'd32639});
	test_expansion(128'h22a1177dc2d96328ccece8abc55b725f, {16'd25568, 16'd54798, 16'd52148, 16'd52720, 16'd52207, 16'd14602, 16'd35494, 16'd13152, 16'd10721, 16'd38553, 16'd9477, 16'd27652, 16'd38557, 16'd16300, 16'd43316, 16'd63930, 16'd18959, 16'd14465, 16'd60795, 16'd27494, 16'd1205, 16'd44503, 16'd6350, 16'd19485, 16'd30784, 16'd39679});
	test_expansion(128'h7c710c12d299aa24944a519062c03e81, {16'd33015, 16'd27680, 16'd9048, 16'd10701, 16'd32772, 16'd10368, 16'd58219, 16'd29628, 16'd55488, 16'd28389, 16'd27200, 16'd57152, 16'd61591, 16'd38144, 16'd36982, 16'd49829, 16'd62426, 16'd53517, 16'd24971, 16'd32213, 16'd41056, 16'd26608, 16'd62704, 16'd65366, 16'd28609, 16'd42515});
	test_expansion(128'h812ac95ddcb8739ad2aee7d31386b54c, {16'd36218, 16'd9224, 16'd61793, 16'd10573, 16'd50399, 16'd38575, 16'd13319, 16'd36851, 16'd31280, 16'd36563, 16'd60501, 16'd31674, 16'd16666, 16'd6614, 16'd60577, 16'd53914, 16'd9265, 16'd52572, 16'd21630, 16'd8117, 16'd51752, 16'd61546, 16'd60909, 16'd38554, 16'd2896, 16'd12792});
	test_expansion(128'h10a7a953f40ebb7af76f4532740a11a1, {16'd16142, 16'd40183, 16'd7238, 16'd36581, 16'd25957, 16'd50069, 16'd22807, 16'd19589, 16'd11577, 16'd64532, 16'd57743, 16'd19920, 16'd40018, 16'd31452, 16'd63747, 16'd24479, 16'd28995, 16'd53520, 16'd49170, 16'd3226, 16'd56916, 16'd55772, 16'd36264, 16'd26190, 16'd17768, 16'd34093});
	test_expansion(128'h5a0ca98eb1fe31bb8d8becfd46df5847, {16'd25473, 16'd6576, 16'd25999, 16'd1768, 16'd41698, 16'd48125, 16'd2636, 16'd15013, 16'd30327, 16'd36673, 16'd20157, 16'd44451, 16'd58059, 16'd61580, 16'd2621, 16'd32569, 16'd33864, 16'd12314, 16'd26421, 16'd5967, 16'd54730, 16'd18499, 16'd17226, 16'd13514, 16'd6251, 16'd36294});
	test_expansion(128'h22ed0135dafe132da9ded3cd4fd6cf4d, {16'd8310, 16'd26148, 16'd60618, 16'd16802, 16'd29045, 16'd59377, 16'd53695, 16'd28000, 16'd44828, 16'd13974, 16'd38236, 16'd38048, 16'd38516, 16'd594, 16'd50434, 16'd7266, 16'd17349, 16'd6548, 16'd48723, 16'd14495, 16'd11949, 16'd12315, 16'd17177, 16'd30415, 16'd39299, 16'd52404});
	test_expansion(128'hfc618bb8b2b8ebe1543ab7e3fcf0102d, {16'd24444, 16'd25834, 16'd27272, 16'd17596, 16'd63064, 16'd40869, 16'd37061, 16'd46397, 16'd17403, 16'd54899, 16'd41648, 16'd21973, 16'd60335, 16'd8952, 16'd36897, 16'd41272, 16'd8584, 16'd46572, 16'd27604, 16'd64310, 16'd24763, 16'd58933, 16'd50071, 16'd7436, 16'd31725, 16'd6122});
	test_expansion(128'h25045efd97ac84b266066d9300234c16, {16'd8787, 16'd2737, 16'd57371, 16'd25509, 16'd2966, 16'd24792, 16'd36095, 16'd21020, 16'd28795, 16'd58236, 16'd4611, 16'd46431, 16'd47686, 16'd40989, 16'd47856, 16'd5949, 16'd45574, 16'd19002, 16'd65153, 16'd51636, 16'd17624, 16'd7864, 16'd36211, 16'd17966, 16'd29940, 16'd7347});
	test_expansion(128'h85f95a5ceeaa890fe9a9574798ff857f, {16'd39722, 16'd6429, 16'd18682, 16'd4332, 16'd64864, 16'd28745, 16'd49864, 16'd43558, 16'd1466, 16'd6211, 16'd431, 16'd13214, 16'd18228, 16'd29649, 16'd14544, 16'd33179, 16'd44348, 16'd10509, 16'd28375, 16'd35879, 16'd24747, 16'd27447, 16'd22742, 16'd18412, 16'd65512, 16'd6778});
	test_expansion(128'hd56d2cc94e573c2570b25ec358dce8cc, {16'd17062, 16'd23826, 16'd7610, 16'd58904, 16'd23898, 16'd57297, 16'd737, 16'd32006, 16'd12346, 16'd30442, 16'd37810, 16'd17483, 16'd54389, 16'd12522, 16'd62647, 16'd60088, 16'd48988, 16'd18261, 16'd8009, 16'd53948, 16'd62649, 16'd39597, 16'd20101, 16'd2905, 16'd26079, 16'd22936});
	test_expansion(128'hecd9cdb57914b8bc2203f390226d6cd8, {16'd42597, 16'd21184, 16'd34425, 16'd26311, 16'd48275, 16'd13541, 16'd34757, 16'd11783, 16'd62568, 16'd10419, 16'd39902, 16'd38101, 16'd25915, 16'd31878, 16'd54911, 16'd34624, 16'd5013, 16'd41585, 16'd17320, 16'd51986, 16'd65328, 16'd4619, 16'd38138, 16'd40806, 16'd52503, 16'd45224});
	test_expansion(128'h4f0bc389ed73a6451960937131b446fc, {16'd1811, 16'd38684, 16'd18837, 16'd5269, 16'd52688, 16'd8504, 16'd24807, 16'd60500, 16'd49327, 16'd26334, 16'd10, 16'd60281, 16'd18917, 16'd26332, 16'd22516, 16'd20115, 16'd18802, 16'd58291, 16'd8266, 16'd2503, 16'd6364, 16'd16127, 16'd13032, 16'd63065, 16'd57843, 16'd13323});
	test_expansion(128'hd166f87c6077d11ba879e157f4770437, {16'd35421, 16'd31175, 16'd50477, 16'd21794, 16'd4020, 16'd25396, 16'd7647, 16'd3365, 16'd37421, 16'd64779, 16'd38278, 16'd55138, 16'd61764, 16'd6772, 16'd32919, 16'd55229, 16'd44749, 16'd37943, 16'd48787, 16'd55131, 16'd52257, 16'd64441, 16'd56615, 16'd42743, 16'd18539, 16'd47939});
	test_expansion(128'hfd2fc81f15906be80db994b80687c03d, {16'd62320, 16'd52988, 16'd36873, 16'd28191, 16'd53906, 16'd8034, 16'd38601, 16'd48531, 16'd58123, 16'd1726, 16'd24791, 16'd63783, 16'd7457, 16'd37817, 16'd60454, 16'd5455, 16'd37864, 16'd19126, 16'd32608, 16'd14919, 16'd61938, 16'd29717, 16'd25212, 16'd50350, 16'd65202, 16'd22330});
	test_expansion(128'hcea470f625f1fbe3ff5bd8d4f9bdd8ec, {16'd5410, 16'd3620, 16'd54974, 16'd63365, 16'd54112, 16'd29315, 16'd31165, 16'd11579, 16'd31359, 16'd21651, 16'd60841, 16'd37833, 16'd54393, 16'd25533, 16'd9750, 16'd61518, 16'd13956, 16'd50600, 16'd16514, 16'd26347, 16'd38021, 16'd41010, 16'd38194, 16'd9634, 16'd8976, 16'd60060});
	test_expansion(128'hc8ec0f96472de888055e7631a8bd26fa, {16'd22182, 16'd8342, 16'd57128, 16'd44703, 16'd40038, 16'd50186, 16'd17568, 16'd41551, 16'd31557, 16'd34426, 16'd3859, 16'd2598, 16'd25464, 16'd27585, 16'd48466, 16'd950, 16'd15534, 16'd32377, 16'd63805, 16'd1437, 16'd37305, 16'd27877, 16'd63242, 16'd33372, 16'd23635, 16'd13790});
	test_expansion(128'h2e49d7dc0d5a9408c069d257e6ee5beb, {16'd63896, 16'd8472, 16'd29342, 16'd49468, 16'd20876, 16'd32510, 16'd64295, 16'd1755, 16'd3071, 16'd61306, 16'd10459, 16'd64970, 16'd157, 16'd3860, 16'd51398, 16'd25857, 16'd35492, 16'd34750, 16'd34607, 16'd29129, 16'd5085, 16'd21805, 16'd25639, 16'd7657, 16'd400, 16'd28202});
	test_expansion(128'hea9b293239d7c593c01994ed6962daa6, {16'd36918, 16'd15792, 16'd22070, 16'd36062, 16'd49302, 16'd38011, 16'd53902, 16'd35540, 16'd25380, 16'd59172, 16'd8473, 16'd29735, 16'd21027, 16'd11832, 16'd51052, 16'd21063, 16'd40894, 16'd53527, 16'd58383, 16'd51900, 16'd21638, 16'd39672, 16'd48222, 16'd60091, 16'd33860, 16'd59235});
	test_expansion(128'h8206055d4dd1cac7ee30a0a68b90eaad, {16'd7038, 16'd29012, 16'd28040, 16'd28927, 16'd40515, 16'd50057, 16'd24141, 16'd64232, 16'd39124, 16'd5451, 16'd3458, 16'd46978, 16'd44593, 16'd32426, 16'd62546, 16'd31743, 16'd661, 16'd45781, 16'd19786, 16'd48227, 16'd23230, 16'd6373, 16'd107, 16'd38492, 16'd599, 16'd48276});
	test_expansion(128'hd38352b54b31cf96c5388f6d6076d70e, {16'd39491, 16'd22709, 16'd26915, 16'd10205, 16'd5107, 16'd16322, 16'd8506, 16'd7273, 16'd46177, 16'd39143, 16'd63559, 16'd31990, 16'd45092, 16'd26533, 16'd27357, 16'd952, 16'd35207, 16'd2107, 16'd29168, 16'd33761, 16'd56882, 16'd32436, 16'd43173, 16'd43261, 16'd12435, 16'd5572});
	test_expansion(128'hacd383768ebcfcf7fcc0c81938fd200f, {16'd6942, 16'd23549, 16'd46864, 16'd1751, 16'd43797, 16'd38374, 16'd10291, 16'd35217, 16'd50478, 16'd20146, 16'd39080, 16'd31800, 16'd21911, 16'd2187, 16'd40592, 16'd10510, 16'd64982, 16'd65132, 16'd40164, 16'd52729, 16'd12091, 16'd21265, 16'd9978, 16'd11622, 16'd26451, 16'd12134});
	test_expansion(128'h75ef083cf24ff09e22542c7ff4d6c4d2, {16'd60087, 16'd47708, 16'd3068, 16'd12255, 16'd33845, 16'd13664, 16'd21072, 16'd53314, 16'd58800, 16'd46882, 16'd8410, 16'd46152, 16'd29541, 16'd41775, 16'd6510, 16'd42827, 16'd854, 16'd23280, 16'd4753, 16'd10777, 16'd15806, 16'd27523, 16'd15113, 16'd59111, 16'd39544, 16'd9521});
	test_expansion(128'h615f895c437e3f05e19db619067b97c4, {16'd53024, 16'd5698, 16'd38555, 16'd27479, 16'd40755, 16'd21264, 16'd11750, 16'd13132, 16'd11783, 16'd52405, 16'd1182, 16'd36413, 16'd17852, 16'd62635, 16'd61294, 16'd25885, 16'd54947, 16'd14689, 16'd10281, 16'd54949, 16'd63351, 16'd36055, 16'd18061, 16'd60750, 16'd40706, 16'd14610});
	test_expansion(128'h3ad53b62a94c626245bde8b62af7edc0, {16'd32936, 16'd64382, 16'd22766, 16'd8344, 16'd39721, 16'd38460, 16'd46720, 16'd64155, 16'd1698, 16'd63164, 16'd61900, 16'd19961, 16'd5264, 16'd15481, 16'd46422, 16'd14732, 16'd36594, 16'd668, 16'd61217, 16'd61532, 16'd40253, 16'd56244, 16'd28067, 16'd10301, 16'd38795, 16'd10290});
	test_expansion(128'h598c30859927f426a1854dd254adf356, {16'd24413, 16'd59523, 16'd50623, 16'd15521, 16'd26206, 16'd22813, 16'd31197, 16'd45464, 16'd59407, 16'd51303, 16'd28510, 16'd50941, 16'd32913, 16'd54002, 16'd63479, 16'd49969, 16'd25316, 16'd50227, 16'd2062, 16'd29452, 16'd2165, 16'd43857, 16'd39612, 16'd13515, 16'd57579, 16'd16711});
	test_expansion(128'hfcb0ea119cca4279686503d3a71cfc17, {16'd16559, 16'd53745, 16'd53579, 16'd15099, 16'd57636, 16'd25706, 16'd37083, 16'd30767, 16'd8685, 16'd20687, 16'd36629, 16'd33562, 16'd17631, 16'd10682, 16'd31546, 16'd42124, 16'd5332, 16'd42396, 16'd18902, 16'd28992, 16'd13724, 16'd58849, 16'd42727, 16'd43706, 16'd2945, 16'd9971});
	test_expansion(128'hbf0d1f8a732523bf1f5e21f53d1f0518, {16'd58587, 16'd32799, 16'd40462, 16'd64826, 16'd5517, 16'd1848, 16'd53709, 16'd4770, 16'd52345, 16'd45880, 16'd32838, 16'd2927, 16'd8502, 16'd59696, 16'd15206, 16'd64205, 16'd35660, 16'd2011, 16'd1167, 16'd39017, 16'd40275, 16'd7697, 16'd28471, 16'd42976, 16'd24021, 16'd20867});
	test_expansion(128'h7cee7cdaec9e2e0c3aff3ca03a8a90aa, {16'd27244, 16'd33942, 16'd52207, 16'd14778, 16'd32571, 16'd30760, 16'd10991, 16'd55124, 16'd45589, 16'd39368, 16'd28325, 16'd10304, 16'd27505, 16'd32932, 16'd27551, 16'd25352, 16'd23763, 16'd8643, 16'd35671, 16'd50589, 16'd15728, 16'd33549, 16'd46614, 16'd12270, 16'd60994, 16'd23985});
	test_expansion(128'h63ff68b28cfa7143317956b77d49d05b, {16'd1269, 16'd17442, 16'd52858, 16'd9902, 16'd25390, 16'd6301, 16'd40492, 16'd6632, 16'd60104, 16'd9124, 16'd64118, 16'd65367, 16'd44396, 16'd26160, 16'd19003, 16'd58276, 16'd48787, 16'd1809, 16'd57392, 16'd48982, 16'd28778, 16'd47160, 16'd14446, 16'd49779, 16'd40344, 16'd20818});
	test_expansion(128'h55fcbf1546bb053865aeac3386c0c781, {16'd323, 16'd11355, 16'd43960, 16'd47522, 16'd46391, 16'd49043, 16'd45052, 16'd45863, 16'd18309, 16'd49522, 16'd17939, 16'd32439, 16'd16552, 16'd15332, 16'd57630, 16'd7620, 16'd63920, 16'd36716, 16'd33050, 16'd14587, 16'd4649, 16'd35368, 16'd57195, 16'd63545, 16'd65085, 16'd52684});
	test_expansion(128'h398e42a343b29a20039af2e8773d07ef, {16'd49697, 16'd64101, 16'd49390, 16'd53665, 16'd19231, 16'd47195, 16'd8294, 16'd11101, 16'd46814, 16'd26913, 16'd30714, 16'd40090, 16'd26471, 16'd17831, 16'd41063, 16'd51129, 16'd43889, 16'd16734, 16'd40970, 16'd58451, 16'd28372, 16'd52376, 16'd15305, 16'd63363, 16'd25607, 16'd46569});
	test_expansion(128'h29167cd38001cd98b54245b1e8a1e29e, {16'd9391, 16'd22364, 16'd27564, 16'd63120, 16'd32351, 16'd4009, 16'd39859, 16'd679, 16'd54097, 16'd4126, 16'd46691, 16'd46662, 16'd21375, 16'd56771, 16'd54766, 16'd56244, 16'd52748, 16'd34825, 16'd28276, 16'd62893, 16'd19083, 16'd14965, 16'd39796, 16'd62036, 16'd59460, 16'd43484});
	test_expansion(128'h65b32ad14aa0e8eca46be16e687dbdb8, {16'd35251, 16'd39846, 16'd48301, 16'd16982, 16'd6598, 16'd58434, 16'd4049, 16'd20533, 16'd29911, 16'd39024, 16'd5292, 16'd61373, 16'd7158, 16'd4827, 16'd3863, 16'd64245, 16'd21542, 16'd30201, 16'd38041, 16'd3555, 16'd11432, 16'd26733, 16'd44885, 16'd2764, 16'd30128, 16'd63204});
	test_expansion(128'h1d93494b78a0d3450753518bd5d82e79, {16'd6260, 16'd54805, 16'd8907, 16'd30774, 16'd55249, 16'd12529, 16'd48004, 16'd12139, 16'd41794, 16'd60166, 16'd45240, 16'd65453, 16'd818, 16'd26847, 16'd13672, 16'd41312, 16'd12369, 16'd14307, 16'd44065, 16'd18231, 16'd51412, 16'd9741, 16'd18413, 16'd4691, 16'd31985, 16'd37112});
	test_expansion(128'ha6623a68deabd57d9b372467e546d769, {16'd15015, 16'd5205, 16'd46788, 16'd1738, 16'd19540, 16'd37220, 16'd7428, 16'd39409, 16'd64302, 16'd12470, 16'd32627, 16'd10232, 16'd49994, 16'd35452, 16'd21567, 16'd16034, 16'd57903, 16'd55215, 16'd52535, 16'd25196, 16'd24733, 16'd51774, 16'd22340, 16'd15726, 16'd28338, 16'd47687});
	test_expansion(128'h68d93e9489e5652277724108b2a126f8, {16'd22414, 16'd34586, 16'd60855, 16'd2601, 16'd23163, 16'd60903, 16'd44318, 16'd7949, 16'd37526, 16'd27279, 16'd12929, 16'd45264, 16'd36336, 16'd5046, 16'd49271, 16'd41439, 16'd57067, 16'd7018, 16'd5196, 16'd30832, 16'd28402, 16'd57015, 16'd45364, 16'd10875, 16'd46316, 16'd6294});
	test_expansion(128'he4549043b05dc9e8bc490e878f3310b3, {16'd33291, 16'd59703, 16'd26040, 16'd32345, 16'd16245, 16'd64164, 16'd64722, 16'd16889, 16'd12993, 16'd55707, 16'd40069, 16'd19984, 16'd56601, 16'd47909, 16'd12368, 16'd9243, 16'd53132, 16'd22548, 16'd43485, 16'd37879, 16'd16294, 16'd38227, 16'd44384, 16'd59641, 16'd45773, 16'd37428});
	test_expansion(128'ha7090055438e648215b7e70ae4c4f330, {16'd8146, 16'd45857, 16'd60307, 16'd42176, 16'd16053, 16'd44642, 16'd57807, 16'd29401, 16'd60102, 16'd32024, 16'd26534, 16'd27124, 16'd22046, 16'd7763, 16'd49846, 16'd42046, 16'd35930, 16'd20286, 16'd43978, 16'd64060, 16'd42789, 16'd40521, 16'd50081, 16'd18583, 16'd33132, 16'd40520});
	test_expansion(128'h32421489df1051ca867ab1413d875a98, {16'd4888, 16'd51247, 16'd47229, 16'd10133, 16'd40506, 16'd29817, 16'd32807, 16'd49949, 16'd47685, 16'd24278, 16'd52311, 16'd5481, 16'd31368, 16'd26656, 16'd24059, 16'd10490, 16'd19779, 16'd20060, 16'd12191, 16'd38255, 16'd30445, 16'd19319, 16'd22775, 16'd25485, 16'd52121, 16'd61125});
	test_expansion(128'h68cefba54fe44d647d5924de68930679, {16'd14566, 16'd53996, 16'd59740, 16'd27459, 16'd20828, 16'd415, 16'd32495, 16'd12193, 16'd16739, 16'd9396, 16'd9544, 16'd54165, 16'd4753, 16'd257, 16'd43400, 16'd65439, 16'd33674, 16'd19493, 16'd37875, 16'd48593, 16'd42399, 16'd40724, 16'd44704, 16'd24572, 16'd14473, 16'd23454});
	test_expansion(128'h8430608554f8d07674702d8de098833d, {16'd29031, 16'd8870, 16'd65342, 16'd25519, 16'd13369, 16'd58728, 16'd64520, 16'd48118, 16'd39546, 16'd9, 16'd49896, 16'd32532, 16'd26142, 16'd16964, 16'd63062, 16'd2616, 16'd29677, 16'd47245, 16'd32885, 16'd6636, 16'd20131, 16'd62586, 16'd45367, 16'd58196, 16'd1624, 16'd26330});
	test_expansion(128'h26718791caa4fb84b625aa62be3f9d8e, {16'd52471, 16'd38583, 16'd29350, 16'd57870, 16'd59533, 16'd57910, 16'd59005, 16'd57419, 16'd64555, 16'd3922, 16'd38697, 16'd52577, 16'd11491, 16'd40039, 16'd44788, 16'd47068, 16'd33900, 16'd9920, 16'd19397, 16'd63341, 16'd43483, 16'd38366, 16'd58419, 16'd45644, 16'd8319, 16'd28337});
	test_expansion(128'h6774773cfe13df8b4518898bb74b21c8, {16'd22297, 16'd33552, 16'd52139, 16'd53558, 16'd38116, 16'd7760, 16'd62915, 16'd52869, 16'd10022, 16'd63586, 16'd36398, 16'd12132, 16'd62904, 16'd56911, 16'd62991, 16'd40272, 16'd21190, 16'd38212, 16'd13949, 16'd18128, 16'd18511, 16'd12877, 16'd53673, 16'd24619, 16'd3743, 16'd41971});
	test_expansion(128'h9e056d6684d3048e807fbb4aed7876f6, {16'd59159, 16'd48164, 16'd46198, 16'd45185, 16'd17043, 16'd15132, 16'd38105, 16'd26486, 16'd50802, 16'd50364, 16'd25502, 16'd30862, 16'd643, 16'd1847, 16'd38169, 16'd16400, 16'd36894, 16'd63156, 16'd14543, 16'd64778, 16'd53330, 16'd19689, 16'd36635, 16'd2486, 16'd7030, 16'd39015});
	test_expansion(128'hf7298fe170ba1e313d7007989ef7fa58, {16'd4247, 16'd58719, 16'd46920, 16'd31698, 16'd19634, 16'd59106, 16'd28532, 16'd13205, 16'd22514, 16'd14419, 16'd55166, 16'd35900, 16'd17287, 16'd14371, 16'd57740, 16'd36809, 16'd22144, 16'd61278, 16'd44068, 16'd36594, 16'd10380, 16'd22663, 16'd44412, 16'd14603, 16'd63984, 16'd54425});
	test_expansion(128'h378ee93b8f0fd1916ded1a557b8c3731, {16'd57525, 16'd7278, 16'd39685, 16'd61738, 16'd59249, 16'd8187, 16'd60407, 16'd33932, 16'd22510, 16'd3384, 16'd9973, 16'd28091, 16'd22557, 16'd3178, 16'd50114, 16'd7226, 16'd46571, 16'd56615, 16'd10852, 16'd24561, 16'd29348, 16'd3314, 16'd49014, 16'd46987, 16'd9166, 16'd20223});
	test_expansion(128'hbfa2a7c5956da8e5fd2fd381dadd5d52, {16'd31894, 16'd49246, 16'd43858, 16'd26023, 16'd16767, 16'd14162, 16'd41357, 16'd56575, 16'd2339, 16'd60224, 16'd21002, 16'd5352, 16'd60335, 16'd14258, 16'd64657, 16'd879, 16'd31676, 16'd44982, 16'd29657, 16'd4560, 16'd9709, 16'd389, 16'd37315, 16'd39382, 16'd20425, 16'd19958});
	test_expansion(128'h50acdfb62245ab3a20985946d70e91c8, {16'd46566, 16'd29143, 16'd50991, 16'd26994, 16'd52659, 16'd39866, 16'd60619, 16'd16260, 16'd10199, 16'd44129, 16'd19243, 16'd42710, 16'd32974, 16'd2219, 16'd32528, 16'd4349, 16'd19168, 16'd42617, 16'd57819, 16'd11214, 16'd49454, 16'd38253, 16'd30610, 16'd30377, 16'd57058, 16'd2256});
	test_expansion(128'hfce92b68491cce38a262f88d579b4123, {16'd12152, 16'd13299, 16'd23257, 16'd28957, 16'd37048, 16'd5267, 16'd53138, 16'd46106, 16'd19693, 16'd37588, 16'd2244, 16'd51564, 16'd45577, 16'd407, 16'd45868, 16'd42118, 16'd53544, 16'd41709, 16'd40020, 16'd36288, 16'd1831, 16'd12555, 16'd47414, 16'd48709, 16'd32199, 16'd55860});
	test_expansion(128'h8f2e3f21a51c135a7e4770936d92b05c, {16'd39582, 16'd58218, 16'd52754, 16'd1004, 16'd64839, 16'd2172, 16'd32196, 16'd30399, 16'd28071, 16'd18048, 16'd58868, 16'd45199, 16'd46514, 16'd15737, 16'd64882, 16'd61467, 16'd5505, 16'd24489, 16'd28027, 16'd42407, 16'd48298, 16'd7146, 16'd11067, 16'd45945, 16'd58765, 16'd32159});
	test_expansion(128'h14fa88211727c3176ec72eadd8cf629e, {16'd58985, 16'd27478, 16'd36422, 16'd22681, 16'd9239, 16'd16469, 16'd5231, 16'd9897, 16'd63803, 16'd12728, 16'd64980, 16'd22494, 16'd35131, 16'd53064, 16'd13482, 16'd50262, 16'd36883, 16'd53925, 16'd18322, 16'd41033, 16'd47227, 16'd9721, 16'd65276, 16'd10411, 16'd48662, 16'd11474});
	test_expansion(128'hfeaee51220d36bd9e962fc62151c1074, {16'd59505, 16'd35928, 16'd37420, 16'd6558, 16'd28080, 16'd36180, 16'd2167, 16'd30191, 16'd41530, 16'd35441, 16'd16924, 16'd9977, 16'd58259, 16'd45354, 16'd50663, 16'd58068, 16'd621, 16'd27898, 16'd29420, 16'd43672, 16'd21884, 16'd18387, 16'd31844, 16'd56185, 16'd21627, 16'd45561});
	test_expansion(128'h4e56c30a94644d2501ff9e2f5361a8fe, {16'd37131, 16'd38145, 16'd61228, 16'd52600, 16'd52599, 16'd16232, 16'd46952, 16'd25082, 16'd34133, 16'd57450, 16'd20901, 16'd58441, 16'd5588, 16'd254, 16'd36855, 16'd4940, 16'd23761, 16'd58356, 16'd8448, 16'd61967, 16'd10420, 16'd9929, 16'd46329, 16'd16886, 16'd34334, 16'd2519});
	test_expansion(128'ha472dc12834465e2f3e6515b4d682107, {16'd14255, 16'd4484, 16'd33460, 16'd36197, 16'd42772, 16'd3427, 16'd18324, 16'd5116, 16'd29778, 16'd44552, 16'd30429, 16'd13991, 16'd14635, 16'd14803, 16'd27251, 16'd19012, 16'd15741, 16'd28956, 16'd41001, 16'd39816, 16'd30208, 16'd21061, 16'd6128, 16'd8389, 16'd35394, 16'd26736});
	test_expansion(128'h83b89e5103bb752df6af250bbe630e48, {16'd27928, 16'd11091, 16'd52890, 16'd57696, 16'd44829, 16'd16419, 16'd17248, 16'd57877, 16'd42446, 16'd10616, 16'd56997, 16'd14697, 16'd18106, 16'd64840, 16'd61019, 16'd61975, 16'd29222, 16'd12824, 16'd8122, 16'd2528, 16'd31544, 16'd474, 16'd29627, 16'd34382, 16'd8851, 16'd36741});
	test_expansion(128'h5552fa2a1abbe4b522629fdc71e609c4, {16'd53006, 16'd61995, 16'd14606, 16'd27113, 16'd22449, 16'd17254, 16'd41821, 16'd42504, 16'd58650, 16'd33349, 16'd11505, 16'd7385, 16'd47327, 16'd55769, 16'd18500, 16'd33013, 16'd59187, 16'd13771, 16'd51999, 16'd31958, 16'd8036, 16'd45532, 16'd26420, 16'd54792, 16'd15526, 16'd60113});
	test_expansion(128'hd8a7a77e2ade57d99cfca73d6d490005, {16'd32309, 16'd13736, 16'd31581, 16'd59620, 16'd13533, 16'd17616, 16'd63758, 16'd61132, 16'd58776, 16'd49638, 16'd58676, 16'd57370, 16'd3060, 16'd954, 16'd65232, 16'd35204, 16'd51063, 16'd54008, 16'd47852, 16'd61430, 16'd5976, 16'd35196, 16'd25809, 16'd8548, 16'd28410, 16'd51128});
	test_expansion(128'h3054c75f9e66f50ec14cc122dec5b2d3, {16'd51803, 16'd59637, 16'd8274, 16'd27946, 16'd62166, 16'd22575, 16'd49377, 16'd51108, 16'd513, 16'd12350, 16'd18098, 16'd27365, 16'd41767, 16'd43716, 16'd13764, 16'd53901, 16'd51785, 16'd34457, 16'd1980, 16'd47348, 16'd38010, 16'd19308, 16'd512, 16'd32762, 16'd52153, 16'd48801});
	test_expansion(128'hb366affe65f5e08b5e8720cc25840e60, {16'd11984, 16'd11565, 16'd48163, 16'd37647, 16'd4482, 16'd4773, 16'd45960, 16'd57644, 16'd15515, 16'd28447, 16'd62395, 16'd62809, 16'd36139, 16'd23706, 16'd27673, 16'd34209, 16'd7713, 16'd13703, 16'd17771, 16'd55168, 16'd37959, 16'd300, 16'd36022, 16'd41648, 16'd2861, 16'd34542});
	test_expansion(128'h77cf562c12e196d116d3eaaf832a23ae, {16'd17897, 16'd16472, 16'd12535, 16'd37170, 16'd62608, 16'd61683, 16'd30097, 16'd62005, 16'd62320, 16'd39989, 16'd56922, 16'd15108, 16'd4251, 16'd40780, 16'd43784, 16'd49575, 16'd9389, 16'd61165, 16'd33874, 16'd27140, 16'd23204, 16'd34028, 16'd53288, 16'd61264, 16'd4368, 16'd40184});
	test_expansion(128'h9fa2e657b81e396519879690714758af, {16'd13548, 16'd44035, 16'd13004, 16'd52576, 16'd24481, 16'd27820, 16'd15918, 16'd3179, 16'd47701, 16'd43626, 16'd17588, 16'd42518, 16'd57872, 16'd51258, 16'd58579, 16'd63256, 16'd18610, 16'd44654, 16'd9274, 16'd59986, 16'd15013, 16'd56978, 16'd37191, 16'd44610, 16'd11890, 16'd52811});
	test_expansion(128'hc4c91ecddaf8597cb9ada752d17efe30, {16'd6045, 16'd10172, 16'd47922, 16'd5841, 16'd12494, 16'd25105, 16'd42870, 16'd57533, 16'd20416, 16'd40894, 16'd54060, 16'd40623, 16'd17491, 16'd40542, 16'd48502, 16'd45644, 16'd25416, 16'd4715, 16'd1593, 16'd29435, 16'd6652, 16'd25559, 16'd6276, 16'd63631, 16'd32024, 16'd57850});
	test_expansion(128'h6d34a4ef70c35e109d2d55821818e63d, {16'd51688, 16'd20340, 16'd45100, 16'd27035, 16'd54085, 16'd59524, 16'd36564, 16'd24536, 16'd6525, 16'd55732, 16'd35073, 16'd26634, 16'd6216, 16'd51937, 16'd20979, 16'd59346, 16'd50636, 16'd61103, 16'd5032, 16'd9783, 16'd62678, 16'd37258, 16'd57305, 16'd11171, 16'd44541, 16'd49773});
	test_expansion(128'h73a6b1ed6d10170aa3d9333e4297490c, {16'd24366, 16'd13742, 16'd19542, 16'd53732, 16'd35327, 16'd45011, 16'd9760, 16'd59430, 16'd38349, 16'd4859, 16'd54148, 16'd25252, 16'd16968, 16'd16756, 16'd44040, 16'd59772, 16'd29959, 16'd55745, 16'd55875, 16'd30241, 16'd2615, 16'd46247, 16'd22106, 16'd11844, 16'd33650, 16'd48426});
	test_expansion(128'h996443c0f9187a590ff686b503809616, {16'd37500, 16'd50542, 16'd27356, 16'd62967, 16'd65381, 16'd5780, 16'd22873, 16'd21223, 16'd13185, 16'd47602, 16'd46412, 16'd64350, 16'd62816, 16'd11389, 16'd34515, 16'd63875, 16'd9310, 16'd50390, 16'd6482, 16'd23788, 16'd16597, 16'd63037, 16'd49717, 16'd9332, 16'd32503, 16'd61751});
	test_expansion(128'h9a38abb82501ed0a73d46ff955e65985, {16'd45721, 16'd39248, 16'd14937, 16'd8222, 16'd60384, 16'd52528, 16'd65294, 16'd21389, 16'd49361, 16'd58266, 16'd30090, 16'd22405, 16'd36656, 16'd42530, 16'd15859, 16'd7291, 16'd30469, 16'd58086, 16'd30585, 16'd34535, 16'd5791, 16'd29402, 16'd58846, 16'd24830, 16'd42494, 16'd45661});
	test_expansion(128'h42e466ba67f9cb273c8efb55909b80ad, {16'd35798, 16'd28667, 16'd24856, 16'd13234, 16'd54064, 16'd8462, 16'd49876, 16'd58135, 16'd7482, 16'd48687, 16'd14363, 16'd9687, 16'd23607, 16'd5983, 16'd35473, 16'd57435, 16'd34495, 16'd40797, 16'd27204, 16'd34515, 16'd35779, 16'd49592, 16'd46351, 16'd24089, 16'd12561, 16'd26239});
	test_expansion(128'hc475062486e619bf5a6a2605ffda855d, {16'd41085, 16'd21192, 16'd44578, 16'd52180, 16'd15837, 16'd22972, 16'd56227, 16'd3193, 16'd41152, 16'd10138, 16'd19843, 16'd5679, 16'd56685, 16'd60339, 16'd61500, 16'd63302, 16'd12615, 16'd36057, 16'd28811, 16'd22067, 16'd62116, 16'd1804, 16'd3748, 16'd45673, 16'd56563, 16'd45716});
	test_expansion(128'h70f2525f7e6201e1fb269ef97f9c8c15, {16'd7269, 16'd37935, 16'd2574, 16'd18947, 16'd44558, 16'd57007, 16'd17889, 16'd1544, 16'd27019, 16'd26753, 16'd24631, 16'd36352, 16'd50303, 16'd140, 16'd42093, 16'd15242, 16'd8954, 16'd59513, 16'd23800, 16'd33048, 16'd39037, 16'd52272, 16'd9910, 16'd18278, 16'd18075, 16'd862});
	test_expansion(128'h36adb328fa18c17c5a29691cb29cc077, {16'd4650, 16'd21539, 16'd45200, 16'd10715, 16'd6637, 16'd41356, 16'd17690, 16'd52507, 16'd8185, 16'd46882, 16'd25747, 16'd5084, 16'd11564, 16'd30472, 16'd12730, 16'd59596, 16'd17672, 16'd57070, 16'd12970, 16'd10625, 16'd31508, 16'd51654, 16'd30998, 16'd20669, 16'd63261, 16'd4855});
	test_expansion(128'h6483d189d35677af53aa96910b72d575, {16'd43826, 16'd42899, 16'd48961, 16'd6276, 16'd49824, 16'd5775, 16'd13114, 16'd28596, 16'd7641, 16'd20972, 16'd46736, 16'd40750, 16'd54480, 16'd49018, 16'd40567, 16'd60737, 16'd31299, 16'd24217, 16'd53623, 16'd45322, 16'd4895, 16'd9491, 16'd9147, 16'd32531, 16'd28089, 16'd59876});
	test_expansion(128'h78a04df836b698163a67bdf55e699a9e, {16'd35291, 16'd31694, 16'd26699, 16'd34301, 16'd43323, 16'd10279, 16'd62558, 16'd366, 16'd14063, 16'd24623, 16'd51327, 16'd51926, 16'd50864, 16'd17877, 16'd43675, 16'd54354, 16'd30845, 16'd38242, 16'd8404, 16'd36696, 16'd26239, 16'd5767, 16'd65465, 16'd57724, 16'd14300, 16'd50548});
	test_expansion(128'h641ce9528ff489ff011adf079f2839a5, {16'd34766, 16'd13587, 16'd27400, 16'd55471, 16'd51152, 16'd7012, 16'd7786, 16'd9216, 16'd26061, 16'd32854, 16'd10011, 16'd22805, 16'd55252, 16'd46905, 16'd38717, 16'd16515, 16'd36403, 16'd59604, 16'd27284, 16'd11463, 16'd707, 16'd44681, 16'd41670, 16'd20562, 16'd38505, 16'd18907});
	test_expansion(128'h03f30deb8fb74526f2c33423f0b6ec87, {16'd26076, 16'd23252, 16'd23476, 16'd58665, 16'd47119, 16'd31287, 16'd5613, 16'd33831, 16'd45206, 16'd58428, 16'd42522, 16'd26044, 16'd19006, 16'd59703, 16'd10227, 16'd58012, 16'd58471, 16'd56510, 16'd1492, 16'd10963, 16'd30673, 16'd42752, 16'd5353, 16'd53690, 16'd45965, 16'd26126});
	test_expansion(128'h540990b68570c8703d2c0826bea7ff31, {16'd61017, 16'd27787, 16'd63603, 16'd28224, 16'd43580, 16'd47170, 16'd15319, 16'd25569, 16'd9817, 16'd17155, 16'd14996, 16'd47344, 16'd55423, 16'd17856, 16'd52586, 16'd28461, 16'd50435, 16'd14752, 16'd25717, 16'd41441, 16'd17516, 16'd13600, 16'd45332, 16'd51009, 16'd52645, 16'd36631});
	test_expansion(128'h83bac56dd438823fdaa8ccccaf2e696d, {16'd31693, 16'd53955, 16'd25792, 16'd23694, 16'd47409, 16'd6882, 16'd33828, 16'd44583, 16'd64157, 16'd42229, 16'd53906, 16'd42507, 16'd31597, 16'd57627, 16'd43970, 16'd18013, 16'd19255, 16'd2904, 16'd42311, 16'd40986, 16'd7819, 16'd57464, 16'd7963, 16'd24038, 16'd18856, 16'd42746});
	test_expansion(128'hcbb0fa200df6c73692b4470f57584b96, {16'd20166, 16'd21501, 16'd26901, 16'd14657, 16'd46549, 16'd60628, 16'd13770, 16'd52493, 16'd17994, 16'd3937, 16'd33960, 16'd23703, 16'd27609, 16'd32404, 16'd31779, 16'd53161, 16'd1894, 16'd10268, 16'd13600, 16'd53652, 16'd15803, 16'd749, 16'd10009, 16'd9039, 16'd14151, 16'd8969});
	test_expansion(128'h7e13ed1fbda00635492597e8f11d2503, {16'd59672, 16'd48367, 16'd57053, 16'd64362, 16'd33387, 16'd30954, 16'd7416, 16'd63911, 16'd35989, 16'd52130, 16'd43055, 16'd20322, 16'd32996, 16'd57590, 16'd2838, 16'd4785, 16'd19768, 16'd27039, 16'd38079, 16'd22149, 16'd52060, 16'd48014, 16'd11459, 16'd41163, 16'd6119, 16'd9663});
	test_expansion(128'haed03c79ecf545aeab5e345ad295a2e8, {16'd35061, 16'd17144, 16'd63150, 16'd21777, 16'd40618, 16'd14713, 16'd59076, 16'd52203, 16'd65074, 16'd40093, 16'd47041, 16'd237, 16'd31190, 16'd8925, 16'd20313, 16'd16607, 16'd42936, 16'd56714, 16'd7033, 16'd53166, 16'd18754, 16'd23983, 16'd56419, 16'd27736, 16'd23138, 16'd49868});
	test_expansion(128'hfee715a0d9ceb6ef6765e1f754566083, {16'd5629, 16'd40790, 16'd7942, 16'd54401, 16'd31972, 16'd16934, 16'd15634, 16'd27645, 16'd4378, 16'd40368, 16'd54536, 16'd53566, 16'd25296, 16'd63633, 16'd44471, 16'd48087, 16'd2172, 16'd64435, 16'd5044, 16'd46578, 16'd32320, 16'd10036, 16'd36833, 16'd30173, 16'd65531, 16'd33695});
	test_expansion(128'hb5a1d0eb0144615bbcfdd42a1aab2e24, {16'd30991, 16'd29070, 16'd56122, 16'd24235, 16'd4601, 16'd6895, 16'd37900, 16'd18163, 16'd63735, 16'd20, 16'd63490, 16'd55818, 16'd55279, 16'd19742, 16'd43399, 16'd24532, 16'd40070, 16'd17577, 16'd45191, 16'd6041, 16'd3137, 16'd5805, 16'd24340, 16'd59928, 16'd32972, 16'd48896});
	test_expansion(128'h7a4a9f5ea00c778ea3174be572461c6d, {16'd40707, 16'd31288, 16'd52495, 16'd25230, 16'd11644, 16'd62435, 16'd8132, 16'd10824, 16'd42298, 16'd57227, 16'd27336, 16'd32470, 16'd38448, 16'd4273, 16'd61632, 16'd28483, 16'd48229, 16'd49288, 16'd55704, 16'd9797, 16'd21656, 16'd40993, 16'd43599, 16'd39995, 16'd53152, 16'd58370});
	test_expansion(128'h7c5af760dd1292b280cde00292faa499, {16'd39629, 16'd53289, 16'd31454, 16'd46648, 16'd26838, 16'd57626, 16'd29568, 16'd59554, 16'd35024, 16'd42787, 16'd50458, 16'd53425, 16'd15477, 16'd51780, 16'd14075, 16'd15269, 16'd12690, 16'd40619, 16'd43683, 16'd9409, 16'd60659, 16'd37261, 16'd53938, 16'd12713, 16'd57403, 16'd16247});
	test_expansion(128'hcb426dceab5edba4ebfdf5981f14bfdf, {16'd14063, 16'd54004, 16'd473, 16'd51390, 16'd41622, 16'd59401, 16'd2741, 16'd43290, 16'd65165, 16'd19621, 16'd61406, 16'd19978, 16'd18974, 16'd8084, 16'd2199, 16'd44478, 16'd52604, 16'd59128, 16'd43788, 16'd8150, 16'd59894, 16'd23137, 16'd16377, 16'd23528, 16'd32793, 16'd25085});
	test_expansion(128'h0d3eaee6852f3035e7d370c3939fc09a, {16'd60870, 16'd37889, 16'd43785, 16'd36849, 16'd62796, 16'd33015, 16'd58553, 16'd43847, 16'd47463, 16'd19517, 16'd11813, 16'd10598, 16'd32359, 16'd8446, 16'd22791, 16'd7023, 16'd30282, 16'd47930, 16'd14105, 16'd22402, 16'd18375, 16'd34433, 16'd35305, 16'd52793, 16'd24368, 16'd27948});
	test_expansion(128'hcc19e2473d2b5d0ff0215c0b1cf4e3b3, {16'd60119, 16'd149, 16'd28483, 16'd56360, 16'd18787, 16'd38580, 16'd19650, 16'd49535, 16'd21702, 16'd39893, 16'd11821, 16'd55751, 16'd5034, 16'd43473, 16'd53939, 16'd58154, 16'd41815, 16'd45757, 16'd51990, 16'd9245, 16'd21062, 16'd30209, 16'd53823, 16'd55198, 16'd11813, 16'd44401});
	test_expansion(128'hd96eb27ec63eee49a6f8039a5d7261fa, {16'd30714, 16'd20083, 16'd30715, 16'd47767, 16'd33256, 16'd31059, 16'd63445, 16'd60025, 16'd53299, 16'd30659, 16'd34570, 16'd43448, 16'd12932, 16'd1403, 16'd56907, 16'd47121, 16'd49608, 16'd46304, 16'd53500, 16'd11877, 16'd54391, 16'd19319, 16'd26590, 16'd64040, 16'd32962, 16'd5500});
	test_expansion(128'h44d685b5c913196c8980ec17bc779cfe, {16'd54606, 16'd12087, 16'd63815, 16'd52765, 16'd25021, 16'd52197, 16'd57844, 16'd40943, 16'd16652, 16'd41997, 16'd53790, 16'd49585, 16'd15997, 16'd22287, 16'd50980, 16'd14824, 16'd38532, 16'd27924, 16'd46311, 16'd17543, 16'd26419, 16'd28542, 16'd10037, 16'd32650, 16'd10948, 16'd43526});
	test_expansion(128'had72cdefd8af4d3b97b9c9c0b5abed44, {16'd14611, 16'd17675, 16'd30314, 16'd48460, 16'd29167, 16'd15946, 16'd24447, 16'd19936, 16'd1105, 16'd9840, 16'd46033, 16'd44267, 16'd16917, 16'd12772, 16'd30512, 16'd22512, 16'd16897, 16'd6928, 16'd3685, 16'd3215, 16'd33063, 16'd10015, 16'd10869, 16'd15245, 16'd43598, 16'd41210});
	test_expansion(128'h2058efd5263b303f7c0ba3bd1ae9a7ab, {16'd60826, 16'd29675, 16'd52606, 16'd30170, 16'd30887, 16'd50503, 16'd48842, 16'd28944, 16'd29689, 16'd19746, 16'd24954, 16'd1043, 16'd61573, 16'd21972, 16'd15894, 16'd47168, 16'd24931, 16'd5352, 16'd65410, 16'd35953, 16'd47472, 16'd8108, 16'd26641, 16'd2261, 16'd10768, 16'd11705});
	test_expansion(128'he4c311d1761739602416c57e2fd5cc04, {16'd55585, 16'd57155, 16'd29762, 16'd15476, 16'd61204, 16'd37660, 16'd48063, 16'd60227, 16'd50383, 16'd37583, 16'd33099, 16'd39199, 16'd49260, 16'd4225, 16'd14655, 16'd16084, 16'd49595, 16'd26041, 16'd15922, 16'd23913, 16'd15871, 16'd9200, 16'd4590, 16'd44146, 16'd30088, 16'd1245});
	test_expansion(128'hf268dd4a4784a999b02f2a2fc72927e4, {16'd12074, 16'd41369, 16'd18570, 16'd34211, 16'd33729, 16'd16395, 16'd22607, 16'd51390, 16'd36358, 16'd53057, 16'd1915, 16'd46899, 16'd52397, 16'd40152, 16'd47557, 16'd341, 16'd11271, 16'd36261, 16'd40955, 16'd14119, 16'd33537, 16'd6630, 16'd49497, 16'd46027, 16'd65500, 16'd48705});
	test_expansion(128'h69656e7cdd2be9e7c4143cfafac1f134, {16'd25832, 16'd33781, 16'd44739, 16'd27565, 16'd3640, 16'd15172, 16'd41895, 16'd35959, 16'd61627, 16'd45870, 16'd48443, 16'd61488, 16'd41904, 16'd42160, 16'd18004, 16'd62858, 16'd30356, 16'd39294, 16'd31058, 16'd62422, 16'd61593, 16'd15470, 16'd47150, 16'd48754, 16'd591, 16'd12525});
	test_expansion(128'ha1d218d53edb2a5adb9f14d4acb5e819, {16'd34343, 16'd5282, 16'd32280, 16'd64460, 16'd34599, 16'd37975, 16'd46114, 16'd12396, 16'd26744, 16'd38931, 16'd40524, 16'd58443, 16'd54803, 16'd17025, 16'd2258, 16'd58270, 16'd5963, 16'd29897, 16'd7384, 16'd41075, 16'd16796, 16'd14505, 16'd17635, 16'd57209, 16'd39278, 16'd16273});
	test_expansion(128'hf2bb3c82ff3bf0ce87f3d9a986c8dbdd, {16'd2013, 16'd57039, 16'd60503, 16'd61390, 16'd6889, 16'd34995, 16'd7566, 16'd51256, 16'd48738, 16'd22499, 16'd55230, 16'd3685, 16'd2966, 16'd31599, 16'd23096, 16'd31536, 16'd49625, 16'd65238, 16'd57728, 16'd19768, 16'd51735, 16'd50319, 16'd62460, 16'd8639, 16'd52577, 16'd41715});
	test_expansion(128'h2ffe88dcd0c31e1692161254febc5f8d, {16'd42663, 16'd55531, 16'd36000, 16'd32648, 16'd48349, 16'd65449, 16'd2785, 16'd40750, 16'd2128, 16'd58015, 16'd39062, 16'd52825, 16'd51745, 16'd50245, 16'd52231, 16'd34700, 16'd23216, 16'd56315, 16'd21935, 16'd32110, 16'd56180, 16'd36250, 16'd56396, 16'd6813, 16'd27775, 16'd49219});
	test_expansion(128'h382fa4e8789540fd703c6892ff398cf3, {16'd2916, 16'd27668, 16'd6441, 16'd34635, 16'd35275, 16'd10791, 16'd18999, 16'd64440, 16'd7058, 16'd61863, 16'd813, 16'd37580, 16'd5922, 16'd39119, 16'd47934, 16'd28364, 16'd42934, 16'd42163, 16'd13168, 16'd49873, 16'd35163, 16'd4323, 16'd30015, 16'd62825, 16'd63920, 16'd24527});
	test_expansion(128'h6b9fd2d8ab463fd09a810db5d41dcf2f, {16'd44916, 16'd33439, 16'd36974, 16'd61820, 16'd2365, 16'd40896, 16'd64301, 16'd64095, 16'd18246, 16'd29285, 16'd3572, 16'd65107, 16'd23248, 16'd10981, 16'd59921, 16'd64297, 16'd55675, 16'd15928, 16'd22357, 16'd28714, 16'd34115, 16'd41073, 16'd6987, 16'd15757, 16'd24015, 16'd64180});
	test_expansion(128'h96ba096c4e627527eb274ae662b0173a, {16'd52069, 16'd65292, 16'd18810, 16'd8486, 16'd26858, 16'd12850, 16'd27135, 16'd41794, 16'd56694, 16'd2383, 16'd10969, 16'd60163, 16'd14516, 16'd11302, 16'd12821, 16'd51098, 16'd39060, 16'd26119, 16'd30877, 16'd52954, 16'd7929, 16'd1669, 16'd58905, 16'd46855, 16'd21350, 16'd38465});
	test_expansion(128'hf0ee92e26d2f5721be3b1e323a3b801c, {16'd21461, 16'd1929, 16'd14717, 16'd55220, 16'd9768, 16'd16565, 16'd32305, 16'd36465, 16'd37661, 16'd12295, 16'd55864, 16'd13783, 16'd61129, 16'd56672, 16'd41036, 16'd13316, 16'd44720, 16'd33470, 16'd32917, 16'd2357, 16'd36154, 16'd30814, 16'd61950, 16'd34639, 16'd3612, 16'd22288});
	test_expansion(128'h4c38dd8749154f0eaf791e8168c24a92, {16'd50237, 16'd22055, 16'd5328, 16'd45008, 16'd15928, 16'd42038, 16'd55290, 16'd24751, 16'd33623, 16'd54400, 16'd5652, 16'd410, 16'd57300, 16'd55221, 16'd60700, 16'd34142, 16'd50850, 16'd7500, 16'd24743, 16'd38322, 16'd25565, 16'd56588, 16'd45853, 16'd15092, 16'd57900, 16'd64593});
	test_expansion(128'habfe697ae428746b04bde5dcc9f39842, {16'd31573, 16'd57110, 16'd44240, 16'd33614, 16'd36586, 16'd34494, 16'd27690, 16'd13749, 16'd21294, 16'd61800, 16'd12358, 16'd30833, 16'd63261, 16'd50709, 16'd2506, 16'd64139, 16'd65118, 16'd24451, 16'd64080, 16'd8713, 16'd47094, 16'd31385, 16'd36282, 16'd47536, 16'd3890, 16'd60150});
	test_expansion(128'h227a45356f85ec7cf068115e5a212994, {16'd65512, 16'd2436, 16'd34952, 16'd43831, 16'd24601, 16'd30998, 16'd21386, 16'd6013, 16'd12272, 16'd36347, 16'd23939, 16'd51815, 16'd65377, 16'd26385, 16'd56988, 16'd17708, 16'd38693, 16'd63685, 16'd63200, 16'd57102, 16'd1232, 16'd54815, 16'd63220, 16'd8452, 16'd8239, 16'd57258});
	test_expansion(128'hb117d56513d3b3ee82915b18b0bb1c77, {16'd49681, 16'd56807, 16'd36756, 16'd45078, 16'd48696, 16'd59722, 16'd39837, 16'd41443, 16'd20657, 16'd54491, 16'd20238, 16'd39720, 16'd25067, 16'd46119, 16'd63164, 16'd64188, 16'd7602, 16'd25860, 16'd4843, 16'd23648, 16'd21096, 16'd15690, 16'd63598, 16'd56575, 16'd25618, 16'd27456});
	test_expansion(128'hd330294c13a57a986fb4a20ea128c288, {16'd56710, 16'd5253, 16'd45202, 16'd14948, 16'd13985, 16'd6190, 16'd3158, 16'd14440, 16'd34919, 16'd33193, 16'd57059, 16'd51759, 16'd59263, 16'd28039, 16'd20856, 16'd51970, 16'd26575, 16'd51529, 16'd43483, 16'd46401, 16'd21751, 16'd19885, 16'd47290, 16'd39802, 16'd63040, 16'd18194});
	test_expansion(128'h3e938b9795ce76c649cf2d7c2e6c3de5, {16'd20441, 16'd62825, 16'd41706, 16'd30620, 16'd9730, 16'd28686, 16'd9523, 16'd46282, 16'd47960, 16'd28445, 16'd9531, 16'd38542, 16'd8411, 16'd43984, 16'd3513, 16'd44167, 16'd10853, 16'd50134, 16'd11869, 16'd49115, 16'd62483, 16'd1832, 16'd39714, 16'd64292, 16'd35479, 16'd64479});
	test_expansion(128'h30870b8b6d1205e5c6c55c5de695dd1e, {16'd49348, 16'd57093, 16'd20158, 16'd40631, 16'd1620, 16'd60763, 16'd37418, 16'd13534, 16'd36158, 16'd1116, 16'd52881, 16'd63393, 16'd1975, 16'd38965, 16'd58751, 16'd26320, 16'd2479, 16'd46775, 16'd14996, 16'd57733, 16'd31725, 16'd50268, 16'd56697, 16'd58004, 16'd26838, 16'd37613});
	test_expansion(128'h8a3d6546c8367feac86fd072560989cf, {16'd26821, 16'd38973, 16'd31830, 16'd54130, 16'd40256, 16'd62327, 16'd35125, 16'd32743, 16'd11535, 16'd41669, 16'd12573, 16'd46742, 16'd61033, 16'd51505, 16'd54862, 16'd17076, 16'd53096, 16'd52017, 16'd33568, 16'd46004, 16'd8205, 16'd40905, 16'd465, 16'd20674, 16'd50581, 16'd65239});
	test_expansion(128'h2f7029bb493ec16cebe3aafd7a5baa8d, {16'd27568, 16'd555, 16'd46145, 16'd11579, 16'd1808, 16'd7759, 16'd64345, 16'd6866, 16'd21609, 16'd14214, 16'd2844, 16'd38310, 16'd35287, 16'd58526, 16'd40129, 16'd43291, 16'd47210, 16'd29784, 16'd57038, 16'd54962, 16'd31888, 16'd37756, 16'd18951, 16'd12110, 16'd20041, 16'd26322});
	test_expansion(128'h06fab94a192586834e1cf4db813d23f1, {16'd8078, 16'd1254, 16'd20504, 16'd10145, 16'd28875, 16'd42352, 16'd50785, 16'd12258, 16'd25966, 16'd64079, 16'd39764, 16'd52242, 16'd40664, 16'd16216, 16'd21629, 16'd25271, 16'd53376, 16'd56739, 16'd29984, 16'd14613, 16'd45391, 16'd30786, 16'd43054, 16'd22244, 16'd50104, 16'd24755});
	test_expansion(128'hbec5ce93b22992e92340769fbbd97ded, {16'd13721, 16'd50093, 16'd47549, 16'd21519, 16'd31524, 16'd10767, 16'd44902, 16'd20118, 16'd9316, 16'd30852, 16'd57930, 16'd61005, 16'd24426, 16'd62894, 16'd17200, 16'd45271, 16'd11874, 16'd49620, 16'd11778, 16'd15219, 16'd51195, 16'd26510, 16'd34587, 16'd64715, 16'd47949, 16'd10708});
	test_expansion(128'h27c9ae1ab17183cdc9b64e4731fcb225, {16'd48872, 16'd2806, 16'd16079, 16'd53791, 16'd4097, 16'd14445, 16'd46750, 16'd22292, 16'd2713, 16'd3031, 16'd25725, 16'd28176, 16'd41290, 16'd8894, 16'd46952, 16'd25853, 16'd15248, 16'd6682, 16'd25846, 16'd39418, 16'd10671, 16'd58424, 16'd9022, 16'd35403, 16'd52992, 16'd20981});
	test_expansion(128'h25fbd12523065ef8ae51590192fd9a5c, {16'd37991, 16'd12095, 16'd56510, 16'd37912, 16'd1303, 16'd34464, 16'd63137, 16'd457, 16'd56754, 16'd38881, 16'd59021, 16'd10769, 16'd58403, 16'd57232, 16'd32028, 16'd50583, 16'd1326, 16'd22779, 16'd30702, 16'd8861, 16'd32103, 16'd33059, 16'd17143, 16'd30108, 16'd18564, 16'd24656});
	test_expansion(128'h065006ff452f74aaa74f8509860508e2, {16'd60162, 16'd15637, 16'd10788, 16'd5177, 16'd20827, 16'd13201, 16'd55743, 16'd60883, 16'd8289, 16'd10831, 16'd61622, 16'd17404, 16'd6600, 16'd36068, 16'd23341, 16'd13997, 16'd59783, 16'd61247, 16'd4889, 16'd34983, 16'd22949, 16'd24630, 16'd32111, 16'd6533, 16'd2507, 16'd17232});
	test_expansion(128'h39b13d1e8a9698d0df84923b11f06c3f, {16'd5907, 16'd38654, 16'd45783, 16'd18158, 16'd27424, 16'd46414, 16'd58693, 16'd58081, 16'd41011, 16'd6706, 16'd30457, 16'd40367, 16'd43835, 16'd46439, 16'd29052, 16'd5450, 16'd32181, 16'd14675, 16'd36128, 16'd57842, 16'd28769, 16'd31108, 16'd32193, 16'd58590, 16'd15311, 16'd44419});
	test_expansion(128'h138b19fb17109735a8879f7ae77a2776, {16'd62070, 16'd48648, 16'd19245, 16'd3806, 16'd65277, 16'd62330, 16'd53412, 16'd20205, 16'd25728, 16'd35257, 16'd16757, 16'd17176, 16'd1254, 16'd8484, 16'd58229, 16'd29519, 16'd44854, 16'd53116, 16'd62350, 16'd21322, 16'd12754, 16'd55342, 16'd44874, 16'd25412, 16'd18345, 16'd52557});
	test_expansion(128'h50ed0ad7c3fa7d83ca8f8853dd38e5ac, {16'd43072, 16'd12682, 16'd33682, 16'd49883, 16'd47646, 16'd38995, 16'd43703, 16'd25227, 16'd44330, 16'd49211, 16'd20144, 16'd30646, 16'd56170, 16'd16156, 16'd31794, 16'd37198, 16'd20217, 16'd25010, 16'd51166, 16'd42553, 16'd3192, 16'd43862, 16'd61875, 16'd56875, 16'd35345, 16'd12797});
	test_expansion(128'h17a9ce8550d34a4eeea479e150cd4429, {16'd40119, 16'd28165, 16'd40312, 16'd35160, 16'd20366, 16'd63602, 16'd48787, 16'd50794, 16'd27208, 16'd18888, 16'd39324, 16'd14018, 16'd9873, 16'd2104, 16'd55147, 16'd65005, 16'd50437, 16'd12436, 16'd36558, 16'd28616, 16'd7957, 16'd23124, 16'd44664, 16'd1453, 16'd35101, 16'd64205});
	test_expansion(128'h3d5ea7f2a909d0457eb221d52bda4749, {16'd17567, 16'd54690, 16'd24958, 16'd37878, 16'd29008, 16'd55979, 16'd58389, 16'd64454, 16'd54442, 16'd29444, 16'd20184, 16'd15862, 16'd2278, 16'd1300, 16'd22638, 16'd37831, 16'd45154, 16'd21522, 16'd4228, 16'd28656, 16'd5608, 16'd7213, 16'd50476, 16'd51496, 16'd24553, 16'd26371});
	test_expansion(128'hcd5c369c4fd3e8bb97190f875ea9c3b5, {16'd42842, 16'd22430, 16'd13558, 16'd4113, 16'd47467, 16'd35328, 16'd18151, 16'd28651, 16'd35550, 16'd41634, 16'd2561, 16'd61263, 16'd14985, 16'd23013, 16'd9172, 16'd40874, 16'd23092, 16'd43482, 16'd23870, 16'd21040, 16'd59239, 16'd39869, 16'd4449, 16'd27566, 16'd30278, 16'd2143});
	test_expansion(128'h5db1fe62cc0f1a58cfeab343ddc1b359, {16'd30615, 16'd42181, 16'd53974, 16'd43378, 16'd56025, 16'd9568, 16'd41466, 16'd64534, 16'd27390, 16'd48731, 16'd62741, 16'd60724, 16'd63690, 16'd46442, 16'd16793, 16'd49391, 16'd42850, 16'd55488, 16'd39821, 16'd9373, 16'd59630, 16'd9063, 16'd11153, 16'd64513, 16'd34302, 16'd24003});
	test_expansion(128'h904882d8a2a9603d0d8b455ca8f07fcb, {16'd41350, 16'd61853, 16'd62733, 16'd484, 16'd28788, 16'd2899, 16'd39550, 16'd19785, 16'd17587, 16'd58, 16'd51127, 16'd34794, 16'd60391, 16'd31804, 16'd19428, 16'd45569, 16'd49198, 16'd34401, 16'd13318, 16'd28797, 16'd26764, 16'd2756, 16'd46393, 16'd56817, 16'd25510, 16'd62529});
	test_expansion(128'h98750ec53820566efb2f04d3334f5775, {16'd22726, 16'd25685, 16'd19298, 16'd7472, 16'd45764, 16'd44925, 16'd11489, 16'd37798, 16'd48335, 16'd56792, 16'd7756, 16'd6809, 16'd48385, 16'd37752, 16'd45834, 16'd1677, 16'd782, 16'd11859, 16'd21192, 16'd41631, 16'd34630, 16'd32589, 16'd26184, 16'd5559, 16'd5394, 16'd57917});
	test_expansion(128'h84652d445b10872cb6cd7c810342cc51, {16'd22706, 16'd59191, 16'd53229, 16'd215, 16'd25801, 16'd26575, 16'd49329, 16'd27574, 16'd49575, 16'd12300, 16'd25585, 16'd1529, 16'd58734, 16'd49754, 16'd42381, 16'd58639, 16'd32090, 16'd41122, 16'd36782, 16'd58416, 16'd19504, 16'd2090, 16'd59061, 16'd28148, 16'd17909, 16'd18073});
	test_expansion(128'h8b7469789cd8696bc383c52c198c4321, {16'd11856, 16'd29901, 16'd45092, 16'd24194, 16'd2428, 16'd44277, 16'd302, 16'd42514, 16'd15676, 16'd57543, 16'd119, 16'd49251, 16'd59062, 16'd3147, 16'd10673, 16'd39659, 16'd17714, 16'd54524, 16'd52529, 16'd8480, 16'd230, 16'd33544, 16'd26262, 16'd33453, 16'd18806, 16'd45367});
	test_expansion(128'ha61cccabb03f351c988e39c2b01cf463, {16'd50763, 16'd7241, 16'd28287, 16'd52182, 16'd41822, 16'd61681, 16'd20164, 16'd4162, 16'd1196, 16'd37569, 16'd18632, 16'd63056, 16'd47594, 16'd51342, 16'd15213, 16'd53077, 16'd55300, 16'd64950, 16'd50426, 16'd8597, 16'd64958, 16'd61179, 16'd20046, 16'd51531, 16'd17827, 16'd64573});
	test_expansion(128'h82d06520006ca3bbfa5d959b9f29a973, {16'd35794, 16'd28311, 16'd10605, 16'd27085, 16'd29717, 16'd38149, 16'd25190, 16'd8348, 16'd15794, 16'd64918, 16'd49364, 16'd11171, 16'd42465, 16'd22885, 16'd28080, 16'd50889, 16'd8942, 16'd55846, 16'd48718, 16'd51649, 16'd28886, 16'd32965, 16'd45807, 16'd56192, 16'd57751, 16'd2966});
	test_expansion(128'h578af914d463f0e4032b5c0cd3d5d713, {16'd32033, 16'd64356, 16'd57877, 16'd38062, 16'd26139, 16'd39087, 16'd57516, 16'd3103, 16'd61373, 16'd26740, 16'd16497, 16'd57148, 16'd19268, 16'd43707, 16'd55483, 16'd48051, 16'd42846, 16'd9351, 16'd19664, 16'd60709, 16'd14128, 16'd5671, 16'd9650, 16'd31492, 16'd51208, 16'd43010});
	test_expansion(128'hf6ebd7c608d80686e6cfb33263a0a3dc, {16'd24132, 16'd53458, 16'd35634, 16'd54076, 16'd44839, 16'd60909, 16'd62332, 16'd54938, 16'd11409, 16'd40540, 16'd19150, 16'd61472, 16'd39084, 16'd49642, 16'd15763, 16'd52205, 16'd55433, 16'd26848, 16'd50490, 16'd32873, 16'd36183, 16'd40674, 16'd57222, 16'd47014, 16'd38430, 16'd36907});
	test_expansion(128'h2f5bee0919c58a81cc0f14b7ef7273d5, {16'd47877, 16'd29226, 16'd40246, 16'd39395, 16'd3247, 16'd21854, 16'd26896, 16'd52549, 16'd26904, 16'd9003, 16'd26666, 16'd30468, 16'd16852, 16'd58090, 16'd24614, 16'd50008, 16'd39504, 16'd57389, 16'd57695, 16'd60836, 16'd60701, 16'd14614, 16'd31772, 16'd61190, 16'd18974, 16'd36439});
	test_expansion(128'h3bee19e9e58d99f09d26cb803fdd5450, {16'd27314, 16'd14416, 16'd13826, 16'd38777, 16'd7266, 16'd62867, 16'd53542, 16'd25637, 16'd19750, 16'd8636, 16'd9472, 16'd18548, 16'd20601, 16'd27385, 16'd31851, 16'd46257, 16'd12275, 16'd33903, 16'd17795, 16'd24652, 16'd65323, 16'd15420, 16'd18725, 16'd63988, 16'd51960, 16'd64492});
	test_expansion(128'hf15a4d5f3582429241ac2bdadf50acec, {16'd23641, 16'd32374, 16'd40404, 16'd63998, 16'd43901, 16'd23478, 16'd581, 16'd59885, 16'd39425, 16'd30582, 16'd50300, 16'd16702, 16'd15529, 16'd2267, 16'd33557, 16'd56101, 16'd3024, 16'd12114, 16'd39123, 16'd4189, 16'd58716, 16'd21249, 16'd5418, 16'd47981, 16'd56800, 16'd24546});
	test_expansion(128'hdf9fe6a96c434287dd4f54f1e0077991, {16'd33225, 16'd58801, 16'd38162, 16'd53143, 16'd63988, 16'd38787, 16'd4536, 16'd17516, 16'd56930, 16'd26169, 16'd21550, 16'd12057, 16'd16354, 16'd43042, 16'd14796, 16'd31833, 16'd21645, 16'd25660, 16'd53261, 16'd20338, 16'd26937, 16'd62485, 16'd61630, 16'd54423, 16'd19022, 16'd917});
	test_expansion(128'h548d52138eb779166863d3ae9c1026b8, {16'd25560, 16'd11639, 16'd38476, 16'd33227, 16'd34372, 16'd64224, 16'd25139, 16'd5070, 16'd48977, 16'd42548, 16'd38718, 16'd38485, 16'd29594, 16'd51340, 16'd5425, 16'd29925, 16'd59428, 16'd52666, 16'd4485, 16'd62578, 16'd35470, 16'd58823, 16'd14984, 16'd63003, 16'd27788, 16'd19938});
	test_expansion(128'h7d13dc227164d4eeddb6159d37920cb9, {16'd35231, 16'd28858, 16'd54350, 16'd16652, 16'd31250, 16'd17814, 16'd18579, 16'd54820, 16'd2105, 16'd26115, 16'd36558, 16'd26450, 16'd52378, 16'd21423, 16'd20464, 16'd943, 16'd32860, 16'd41932, 16'd50561, 16'd23421, 16'd53172, 16'd4281, 16'd31785, 16'd64703, 16'd29247, 16'd38417});
	test_expansion(128'h2a2ad8893df7c567f97ab75ebe4f1063, {16'd2740, 16'd14544, 16'd53881, 16'd6352, 16'd64661, 16'd12683, 16'd52765, 16'd52365, 16'd61628, 16'd35350, 16'd58542, 16'd62949, 16'd15651, 16'd17406, 16'd25026, 16'd52813, 16'd34493, 16'd58744, 16'd62171, 16'd9065, 16'd24895, 16'd44977, 16'd21229, 16'd27820, 16'd50332, 16'd20729});
	test_expansion(128'hb03f26e57cdfc158134448032eba99c0, {16'd49338, 16'd5705, 16'd15135, 16'd34281, 16'd51284, 16'd7476, 16'd29797, 16'd6828, 16'd10381, 16'd240, 16'd19453, 16'd2104, 16'd33456, 16'd56575, 16'd26243, 16'd22166, 16'd37386, 16'd36446, 16'd57708, 16'd28588, 16'd56273, 16'd47096, 16'd16334, 16'd14985, 16'd31101, 16'd17170});
	test_expansion(128'h7ebcac180d159ad86a27a69c483aed6f, {16'd53039, 16'd56108, 16'd52308, 16'd6712, 16'd3631, 16'd40203, 16'd46921, 16'd62013, 16'd37229, 16'd36827, 16'd59667, 16'd40255, 16'd18617, 16'd15891, 16'd38219, 16'd38067, 16'd39129, 16'd19334, 16'd17036, 16'd27584, 16'd11364, 16'd55273, 16'd7254, 16'd54552, 16'd12164, 16'd27534});
	test_expansion(128'h14e586037776c038286ce4065a363b03, {16'd63312, 16'd21366, 16'd29375, 16'd44477, 16'd44223, 16'd19352, 16'd7114, 16'd62968, 16'd4802, 16'd11249, 16'd21377, 16'd13646, 16'd18352, 16'd54063, 16'd32623, 16'd208, 16'd48150, 16'd368, 16'd45252, 16'd57289, 16'd269, 16'd26502, 16'd2222, 16'd52071, 16'd26959, 16'd12630});
	test_expansion(128'hb974754ea52802cc7f018a3a3f51d7c2, {16'd18080, 16'd45646, 16'd50870, 16'd31728, 16'd57976, 16'd63568, 16'd321, 16'd62923, 16'd44522, 16'd39832, 16'd31586, 16'd29134, 16'd31657, 16'd62547, 16'd54480, 16'd49811, 16'd10632, 16'd49948, 16'd58498, 16'd17515, 16'd27363, 16'd6101, 16'd48841, 16'd34998, 16'd39099, 16'd60725});
	test_expansion(128'hc0dd7660b06fdf48836439babfeb2de7, {16'd23842, 16'd5292, 16'd13154, 16'd34051, 16'd21898, 16'd54991, 16'd22430, 16'd37042, 16'd54000, 16'd60996, 16'd52073, 16'd61975, 16'd46236, 16'd11210, 16'd37375, 16'd64233, 16'd18615, 16'd54523, 16'd2476, 16'd20468, 16'd56026, 16'd44793, 16'd14189, 16'd16193, 16'd28088, 16'd49463});
	test_expansion(128'he461088ffb443ef9c7f0eacac2db6f3e, {16'd10829, 16'd49617, 16'd57798, 16'd31057, 16'd2740, 16'd55528, 16'd38857, 16'd6490, 16'd62727, 16'd12858, 16'd23304, 16'd52159, 16'd48526, 16'd1680, 16'd47402, 16'd61594, 16'd55485, 16'd50803, 16'd26122, 16'd46277, 16'd48723, 16'd4053, 16'd63482, 16'd2027, 16'd40049, 16'd26085});
	test_expansion(128'h956536aa1503e2427435250616682776, {16'd1598, 16'd32602, 16'd39289, 16'd56382, 16'd60889, 16'd21936, 16'd31321, 16'd22264, 16'd319, 16'd30692, 16'd19493, 16'd62573, 16'd44166, 16'd19894, 16'd56403, 16'd26180, 16'd28845, 16'd19583, 16'd40466, 16'd37362, 16'd13668, 16'd256, 16'd57335, 16'd41242, 16'd48552, 16'd16396});
	test_expansion(128'hdf16a0b4772ff36008ac37baee48d587, {16'd6982, 16'd26181, 16'd46566, 16'd40580, 16'd45895, 16'd47977, 16'd58024, 16'd54738, 16'd5664, 16'd47742, 16'd55571, 16'd51877, 16'd56233, 16'd35407, 16'd16568, 16'd65174, 16'd2676, 16'd46930, 16'd21239, 16'd14589, 16'd49542, 16'd198, 16'd11136, 16'd50191, 16'd44386, 16'd56102});
	test_expansion(128'he57813991f51fe09765041bb0c30685f, {16'd38141, 16'd29706, 16'd24616, 16'd54116, 16'd24257, 16'd53631, 16'd30469, 16'd42316, 16'd57701, 16'd60593, 16'd33180, 16'd46947, 16'd41362, 16'd54976, 16'd17797, 16'd31459, 16'd243, 16'd42656, 16'd5047, 16'd16954, 16'd959, 16'd41342, 16'd32520, 16'd41384, 16'd34217, 16'd41900});
	test_expansion(128'hcaae20a2106a867dab96e02b8ef119c3, {16'd17571, 16'd17027, 16'd19489, 16'd32126, 16'd23810, 16'd10756, 16'd52368, 16'd24255, 16'd22628, 16'd35374, 16'd41562, 16'd6750, 16'd54601, 16'd39507, 16'd50335, 16'd283, 16'd22624, 16'd39606, 16'd46269, 16'd55405, 16'd43623, 16'd25200, 16'd12420, 16'd59602, 16'd36749, 16'd21605});
	test_expansion(128'hfd3b0f3a450108b668cba2363786b197, {16'd33259, 16'd29454, 16'd6914, 16'd54691, 16'd26812, 16'd2137, 16'd5651, 16'd43478, 16'd27437, 16'd9724, 16'd5108, 16'd45261, 16'd29822, 16'd41559, 16'd57183, 16'd57531, 16'd6274, 16'd6784, 16'd33693, 16'd26173, 16'd9649, 16'd30295, 16'd33665, 16'd49027, 16'd9035, 16'd47682});
	test_expansion(128'hf3721b3d089b7587757662c52c784176, {16'd53630, 16'd15246, 16'd48343, 16'd10871, 16'd43987, 16'd49651, 16'd9471, 16'd25613, 16'd26851, 16'd28687, 16'd48178, 16'd6871, 16'd7400, 16'd2816, 16'd15338, 16'd15325, 16'd24847, 16'd6751, 16'd3453, 16'd28707, 16'd37764, 16'd30997, 16'd23186, 16'd25288, 16'd39739, 16'd10690});
	test_expansion(128'hb581786c4354d6277a366c864c4b1640, {16'd30703, 16'd44666, 16'd15370, 16'd52328, 16'd8241, 16'd38750, 16'd2638, 16'd11936, 16'd1003, 16'd22617, 16'd27709, 16'd47956, 16'd25591, 16'd45341, 16'd58296, 16'd34388, 16'd8862, 16'd6678, 16'd35323, 16'd25056, 16'd46932, 16'd17930, 16'd60919, 16'd58859, 16'd56257, 16'd1741});
	test_expansion(128'hc135c70cba3b6bbfa624d217b30c5559, {16'd49326, 16'd17905, 16'd26744, 16'd33192, 16'd2156, 16'd52094, 16'd26804, 16'd27937, 16'd38198, 16'd32030, 16'd14957, 16'd12645, 16'd33107, 16'd13414, 16'd32195, 16'd1461, 16'd43522, 16'd55123, 16'd24335, 16'd47711, 16'd62744, 16'd38208, 16'd21928, 16'd50951, 16'd4062, 16'd14268});
	test_expansion(128'hc84c49673ee2ca5b55b6705678f5cadc, {16'd13651, 16'd17384, 16'd25538, 16'd21503, 16'd7166, 16'd53115, 16'd51406, 16'd50073, 16'd8356, 16'd16213, 16'd61299, 16'd49950, 16'd20348, 16'd11097, 16'd50784, 16'd8284, 16'd65004, 16'd17595, 16'd32737, 16'd4110, 16'd22514, 16'd9991, 16'd19348, 16'd9143, 16'd287, 16'd46156});
	test_expansion(128'he94af4e71503a3fcebb327dd7f82a7bc, {16'd55657, 16'd26727, 16'd20613, 16'd15756, 16'd14052, 16'd25529, 16'd3222, 16'd22964, 16'd11599, 16'd59238, 16'd49519, 16'd58255, 16'd28780, 16'd38998, 16'd24760, 16'd8457, 16'd37703, 16'd47432, 16'd54579, 16'd12229, 16'd45202, 16'd65257, 16'd39711, 16'd5638, 16'd12448, 16'd57141});
	test_expansion(128'hb1a33c63e1a8a31d6ce36d1b530f2c1d, {16'd46353, 16'd26261, 16'd63823, 16'd19867, 16'd44171, 16'd2764, 16'd33434, 16'd32261, 16'd57382, 16'd14184, 16'd52637, 16'd50195, 16'd20261, 16'd25324, 16'd57249, 16'd19736, 16'd26017, 16'd28125, 16'd46367, 16'd59275, 16'd30140, 16'd51605, 16'd30478, 16'd50229, 16'd40457, 16'd38618});
	test_expansion(128'hb771eb233ea0bd0e90a00e9aea6886f9, {16'd1293, 16'd12681, 16'd63268, 16'd39578, 16'd57760, 16'd51699, 16'd18531, 16'd42074, 16'd38513, 16'd18849, 16'd29953, 16'd16702, 16'd21769, 16'd8916, 16'd27240, 16'd31940, 16'd6379, 16'd14393, 16'd14515, 16'd22701, 16'd13956, 16'd18708, 16'd30290, 16'd1338, 16'd55394, 16'd1912});
	test_expansion(128'hcd681f67cdb0df4a93f846446b5e8ca5, {16'd1100, 16'd13094, 16'd52492, 16'd16189, 16'd28771, 16'd35824, 16'd7157, 16'd15187, 16'd16394, 16'd17735, 16'd47236, 16'd20778, 16'd30038, 16'd57055, 16'd44802, 16'd49739, 16'd1314, 16'd55329, 16'd16303, 16'd26728, 16'd45251, 16'd22856, 16'd27019, 16'd63564, 16'd16734, 16'd52456});
	test_expansion(128'h44a9ee29f3f95255c9f0f283ba252d99, {16'd24692, 16'd1852, 16'd31231, 16'd41570, 16'd10287, 16'd43255, 16'd56457, 16'd62245, 16'd56783, 16'd21532, 16'd2018, 16'd47975, 16'd7479, 16'd25865, 16'd17010, 16'd6309, 16'd24717, 16'd57223, 16'd25574, 16'd49764, 16'd14372, 16'd39753, 16'd64997, 16'd18664, 16'd22074, 16'd38426});
	test_expansion(128'h766cd4ede6d9d1278bbc2ce7fced7613, {16'd11604, 16'd32278, 16'd52162, 16'd4893, 16'd34465, 16'd8429, 16'd49857, 16'd49396, 16'd1966, 16'd43605, 16'd26659, 16'd41900, 16'd54316, 16'd7543, 16'd55600, 16'd43319, 16'd54920, 16'd45280, 16'd3511, 16'd10956, 16'd63294, 16'd37726, 16'd57507, 16'd28151, 16'd55288, 16'd55589});
	test_expansion(128'hf1f73bc92811cd03d5d1603bee825cce, {16'd204, 16'd21893, 16'd9539, 16'd33001, 16'd27246, 16'd57294, 16'd35246, 16'd7415, 16'd63613, 16'd2413, 16'd47102, 16'd39503, 16'd23121, 16'd19211, 16'd6524, 16'd41117, 16'd63510, 16'd28560, 16'd39207, 16'd21983, 16'd57566, 16'd59229, 16'd39506, 16'd29451, 16'd61296, 16'd55900});
	test_expansion(128'h8c8f97b605c654fd00ffbbec49e3a59d, {16'd2686, 16'd36874, 16'd56540, 16'd4512, 16'd27302, 16'd39159, 16'd58635, 16'd64372, 16'd13814, 16'd64927, 16'd56923, 16'd13051, 16'd22808, 16'd50728, 16'd20087, 16'd22547, 16'd43188, 16'd4577, 16'd57159, 16'd1941, 16'd48466, 16'd63237, 16'd34225, 16'd28467, 16'd56911, 16'd17261});
	test_expansion(128'hcf5499ea341909f1c9fc4234e62f8e75, {16'd62459, 16'd1550, 16'd58380, 16'd4265, 16'd62719, 16'd64007, 16'd16599, 16'd58008, 16'd11482, 16'd53775, 16'd27980, 16'd57530, 16'd42203, 16'd10842, 16'd63992, 16'd61403, 16'd1096, 16'd34145, 16'd60234, 16'd3487, 16'd37789, 16'd38692, 16'd18347, 16'd5809, 16'd30108, 16'd50978});
	test_expansion(128'h09f2ac6f427b16f4eac0321a0c3b9253, {16'd28673, 16'd30511, 16'd47514, 16'd24278, 16'd5450, 16'd62084, 16'd62114, 16'd36491, 16'd31845, 16'd609, 16'd44997, 16'd37627, 16'd41929, 16'd65049, 16'd9627, 16'd5424, 16'd17171, 16'd52220, 16'd62629, 16'd37291, 16'd60868, 16'd36643, 16'd49907, 16'd54041, 16'd9595, 16'd26755});
	test_expansion(128'h7eeff45d1952b1e6caefb3cf89b9756d, {16'd13003, 16'd31551, 16'd38566, 16'd20829, 16'd26214, 16'd42696, 16'd64760, 16'd54824, 16'd52427, 16'd57573, 16'd52437, 16'd63456, 16'd6909, 16'd7167, 16'd10034, 16'd17771, 16'd48053, 16'd3243, 16'd24865, 16'd22874, 16'd10267, 16'd1102, 16'd20928, 16'd33965, 16'd11940, 16'd30614});
	test_expansion(128'hc1f46a137d10a2384dec90dad8b97b4c, {16'd62627, 16'd17889, 16'd18632, 16'd21071, 16'd42120, 16'd47882, 16'd51057, 16'd16108, 16'd34102, 16'd27269, 16'd36030, 16'd29384, 16'd46826, 16'd52871, 16'd19856, 16'd21835, 16'd9305, 16'd5981, 16'd61143, 16'd22122, 16'd26628, 16'd722, 16'd199, 16'd14520, 16'd52117, 16'd23839});
	test_expansion(128'hb2e3f96e6f6e5a214dd12e5c99520933, {16'd56232, 16'd56596, 16'd37020, 16'd46139, 16'd42322, 16'd31621, 16'd49654, 16'd49475, 16'd44038, 16'd64458, 16'd35030, 16'd2815, 16'd8331, 16'd63567, 16'd47320, 16'd63319, 16'd35291, 16'd62899, 16'd18692, 16'd38226, 16'd43547, 16'd16521, 16'd19960, 16'd33943, 16'd61124, 16'd52716});
	test_expansion(128'h60298460b43fc6987f20dbf83bbaef11, {16'd794, 16'd27919, 16'd3544, 16'd60794, 16'd802, 16'd30011, 16'd33700, 16'd20897, 16'd62130, 16'd58463, 16'd31800, 16'd53078, 16'd40676, 16'd60826, 16'd8808, 16'd45766, 16'd34908, 16'd10003, 16'd31784, 16'd63677, 16'd5247, 16'd33378, 16'd60344, 16'd13615, 16'd60180, 16'd5153});
	test_expansion(128'h14a3762fd78bfd9df1fff25703d84855, {16'd38862, 16'd21510, 16'd4381, 16'd44839, 16'd3643, 16'd40658, 16'd25158, 16'd11443, 16'd48050, 16'd39967, 16'd34285, 16'd63252, 16'd12984, 16'd5810, 16'd29080, 16'd40190, 16'd13837, 16'd16142, 16'd2488, 16'd1580, 16'd46769, 16'd36058, 16'd33728, 16'd52578, 16'd46123, 16'd51583});
	test_expansion(128'h97ff0b523ea2e9c87a736d2c4bef2072, {16'd54792, 16'd11374, 16'd33699, 16'd30641, 16'd23571, 16'd33066, 16'd11652, 16'd63254, 16'd19175, 16'd20150, 16'd3145, 16'd64941, 16'd53223, 16'd4371, 16'd24078, 16'd43539, 16'd33120, 16'd23046, 16'd35565, 16'd46634, 16'd437, 16'd11576, 16'd8750, 16'd46213, 16'd28912, 16'd25720});
	test_expansion(128'h2297b22c88ee4418cbc4202e4c1cecfd, {16'd52663, 16'd63324, 16'd60091, 16'd27951, 16'd28034, 16'd37829, 16'd25653, 16'd10641, 16'd42139, 16'd669, 16'd62632, 16'd8542, 16'd16340, 16'd21967, 16'd50741, 16'd18608, 16'd42179, 16'd31623, 16'd32566, 16'd9886, 16'd3224, 16'd64649, 16'd46349, 16'd35478, 16'd49612, 16'd52006});
	test_expansion(128'h6de87b9eefb2bdd7dbbcc5f158bd0a77, {16'd2119, 16'd42720, 16'd20582, 16'd44500, 16'd31492, 16'd50963, 16'd31376, 16'd54118, 16'd45205, 16'd23660, 16'd52693, 16'd56272, 16'd58428, 16'd30460, 16'd6509, 16'd51642, 16'd49699, 16'd9206, 16'd59256, 16'd48914, 16'd43647, 16'd15867, 16'd38860, 16'd745, 16'd8285, 16'd15388});
	test_expansion(128'h1d167e716a72019a7a3da7f1d5c5bed2, {16'd58656, 16'd63055, 16'd10528, 16'd28132, 16'd16303, 16'd38216, 16'd7186, 16'd24020, 16'd42041, 16'd20720, 16'd8076, 16'd49608, 16'd32824, 16'd14812, 16'd8482, 16'd47127, 16'd52615, 16'd38878, 16'd53936, 16'd32211, 16'd27810, 16'd43188, 16'd7845, 16'd12684, 16'd17340, 16'd41514});
	test_expansion(128'h0c06865120447a8bafc46db87ed33123, {16'd16537, 16'd44378, 16'd49547, 16'd62609, 16'd10242, 16'd55315, 16'd27380, 16'd20140, 16'd56895, 16'd65043, 16'd62805, 16'd40967, 16'd21054, 16'd48281, 16'd58408, 16'd49069, 16'd22774, 16'd52958, 16'd38290, 16'd27823, 16'd48533, 16'd13469, 16'd10922, 16'd7946, 16'd45543, 16'd56413});
	test_expansion(128'h699f9e3ee9d61a6e32f8cd68c2732079, {16'd60466, 16'd29734, 16'd20937, 16'd910, 16'd8288, 16'd23278, 16'd36782, 16'd9498, 16'd42605, 16'd1325, 16'd8489, 16'd19983, 16'd63657, 16'd4550, 16'd2866, 16'd33656, 16'd2980, 16'd60683, 16'd44670, 16'd15267, 16'd53432, 16'd11305, 16'd28544, 16'd58040, 16'd51473, 16'd17038});
	test_expansion(128'hdb08d701116e21d615e97871a585ddf3, {16'd9378, 16'd51695, 16'd30625, 16'd48717, 16'd22327, 16'd20442, 16'd9669, 16'd60930, 16'd56307, 16'd32384, 16'd52435, 16'd5958, 16'd33454, 16'd10351, 16'd25900, 16'd30534, 16'd23861, 16'd44185, 16'd36341, 16'd35453, 16'd2848, 16'd64917, 16'd43063, 16'd2570, 16'd49713, 16'd44898});
	test_expansion(128'hd17b79a7dd38baf1de6eaf9b236ba331, {16'd18746, 16'd39888, 16'd58307, 16'd4105, 16'd24680, 16'd37393, 16'd46058, 16'd64227, 16'd10086, 16'd49521, 16'd37641, 16'd40333, 16'd46694, 16'd18890, 16'd51172, 16'd42649, 16'd59272, 16'd38433, 16'd48321, 16'd6101, 16'd48488, 16'd54674, 16'd16759, 16'd45139, 16'd60924, 16'd55896});
	test_expansion(128'h9d6d7b31b91bbcb986dce83dd85d3648, {16'd11571, 16'd50706, 16'd44809, 16'd22287, 16'd34746, 16'd64284, 16'd41665, 16'd14489, 16'd40556, 16'd37490, 16'd46861, 16'd18663, 16'd2859, 16'd34910, 16'd32972, 16'd17967, 16'd1841, 16'd5775, 16'd31288, 16'd6457, 16'd55794, 16'd9730, 16'd28867, 16'd56928, 16'd8066, 16'd27008});
	test_expansion(128'h7f9cec73b57d14a8823b9697e0d494fb, {16'd5020, 16'd14675, 16'd45961, 16'd32899, 16'd9782, 16'd41215, 16'd15212, 16'd44194, 16'd54958, 16'd57199, 16'd58309, 16'd14085, 16'd3959, 16'd62635, 16'd28691, 16'd39818, 16'd28891, 16'd62954, 16'd42, 16'd24852, 16'd32206, 16'd28107, 16'd15683, 16'd56400, 16'd42291, 16'd44883});
	test_expansion(128'h47d44b60d3ad6a03bb4e921eafe3a521, {16'd12299, 16'd40866, 16'd58261, 16'd30125, 16'd49216, 16'd159, 16'd45156, 16'd54906, 16'd11250, 16'd51550, 16'd33853, 16'd24720, 16'd65004, 16'd18620, 16'd54870, 16'd32618, 16'd22169, 16'd33099, 16'd27974, 16'd40557, 16'd27859, 16'd13457, 16'd17181, 16'd18253, 16'd29173, 16'd50007});
	test_expansion(128'h487bf685402ea391e30c13e4668baac9, {16'd59250, 16'd14578, 16'd13070, 16'd43861, 16'd27697, 16'd55181, 16'd10864, 16'd63532, 16'd26936, 16'd55245, 16'd17561, 16'd57746, 16'd23439, 16'd60049, 16'd43083, 16'd39405, 16'd13025, 16'd21541, 16'd45515, 16'd20648, 16'd56022, 16'd34236, 16'd15587, 16'd35311, 16'd51951, 16'd20423});
	test_expansion(128'ha5a8060a1a64aee5d678b4731b1e5210, {16'd40604, 16'd548, 16'd49742, 16'd13401, 16'd43217, 16'd20703, 16'd62638, 16'd4687, 16'd17679, 16'd36723, 16'd31607, 16'd2104, 16'd61687, 16'd64798, 16'd18165, 16'd5720, 16'd19499, 16'd26247, 16'd51024, 16'd17055, 16'd28652, 16'd21527, 16'd23138, 16'd33307, 16'd25130, 16'd1145});
	test_expansion(128'hfabb0367e66aa1853f4ac31945cfa586, {16'd37582, 16'd18813, 16'd43873, 16'd53760, 16'd5838, 16'd41997, 16'd50506, 16'd17839, 16'd56660, 16'd26891, 16'd5388, 16'd11563, 16'd51957, 16'd35988, 16'd7379, 16'd5536, 16'd58708, 16'd42293, 16'd6117, 16'd22201, 16'd10804, 16'd30249, 16'd8457, 16'd3850, 16'd25654, 16'd28071});
	test_expansion(128'h78ee23de1288fa25ddcf827d25da243b, {16'd65209, 16'd8420, 16'd43381, 16'd34177, 16'd6299, 16'd3954, 16'd43441, 16'd40008, 16'd56657, 16'd49973, 16'd26158, 16'd30482, 16'd7950, 16'd31054, 16'd11097, 16'd49797, 16'd18734, 16'd56991, 16'd47730, 16'd44592, 16'd50427, 16'd487, 16'd39509, 16'd53836, 16'd60150, 16'd40024});
	test_expansion(128'h78e7eb592372c2e13e6baae31a63cce9, {16'd11168, 16'd14089, 16'd60776, 16'd11063, 16'd42756, 16'd28479, 16'd39949, 16'd28669, 16'd54397, 16'd41029, 16'd226, 16'd49580, 16'd42382, 16'd60850, 16'd50653, 16'd37652, 16'd33884, 16'd13282, 16'd53917, 16'd21641, 16'd49240, 16'd12926, 16'd53733, 16'd11507, 16'd11052, 16'd52847});
	test_expansion(128'h844f5ad513cc4fba7e8e967e6967876f, {16'd1611, 16'd46577, 16'd33892, 16'd21509, 16'd41734, 16'd59381, 16'd26841, 16'd36820, 16'd59839, 16'd3034, 16'd32576, 16'd62494, 16'd49333, 16'd49763, 16'd23491, 16'd36421, 16'd4991, 16'd62097, 16'd55122, 16'd10614, 16'd41309, 16'd25549, 16'd63266, 16'd36010, 16'd65410, 16'd5323});
	test_expansion(128'hfbb171e8807bd8518bf448fc59cf70c2, {16'd46945, 16'd27457, 16'd39678, 16'd39599, 16'd3958, 16'd26012, 16'd44312, 16'd11380, 16'd49671, 16'd48973, 16'd15653, 16'd12928, 16'd35188, 16'd33172, 16'd20097, 16'd1328, 16'd53788, 16'd35886, 16'd36392, 16'd46825, 16'd42406, 16'd42059, 16'd36000, 16'd14319, 16'd57307, 16'd30435});
	test_expansion(128'h135a14716075424137cddbaba1f9a209, {16'd58129, 16'd63214, 16'd62807, 16'd48932, 16'd42386, 16'd49121, 16'd5984, 16'd44722, 16'd37909, 16'd37165, 16'd21891, 16'd65372, 16'd59368, 16'd37125, 16'd22751, 16'd31645, 16'd31560, 16'd10996, 16'd59105, 16'd31287, 16'd14159, 16'd7268, 16'd9783, 16'd50159, 16'd42944, 16'd10364});
	test_expansion(128'h847517dd9f8d446ec098a2f80a477223, {16'd59278, 16'd42810, 16'd14691, 16'd62886, 16'd1168, 16'd56503, 16'd35832, 16'd14660, 16'd23205, 16'd51400, 16'd58824, 16'd30899, 16'd16942, 16'd51287, 16'd48568, 16'd51522, 16'd39557, 16'd45470, 16'd57349, 16'd48915, 16'd13648, 16'd20992, 16'd25363, 16'd36237, 16'd5225, 16'd45514});
	test_expansion(128'h2bebfb1f6d96ed2fab2a563ea529f0f7, {16'd12495, 16'd11283, 16'd2921, 16'd44902, 16'd37885, 16'd37495, 16'd50991, 16'd30694, 16'd33080, 16'd51327, 16'd6106, 16'd43908, 16'd26655, 16'd20760, 16'd17346, 16'd61987, 16'd3528, 16'd22731, 16'd64710, 16'd35555, 16'd6544, 16'd39179, 16'd8630, 16'd33909, 16'd53055, 16'd15707});
	test_expansion(128'hd2fc6db6df91c71643059c0903c7c951, {16'd34810, 16'd17221, 16'd14148, 16'd27017, 16'd24377, 16'd56947, 16'd36061, 16'd12921, 16'd5832, 16'd52107, 16'd18957, 16'd32143, 16'd38689, 16'd12180, 16'd57164, 16'd16288, 16'd2554, 16'd24248, 16'd48792, 16'd55647, 16'd31438, 16'd14077, 16'd19655, 16'd64795, 16'd25535, 16'd55474});
	test_expansion(128'hce759a2709ab6ed217f06335296ab7e4, {16'd37982, 16'd27184, 16'd3167, 16'd65509, 16'd59928, 16'd9953, 16'd19896, 16'd17180, 16'd14724, 16'd60540, 16'd11774, 16'd51249, 16'd51904, 16'd33310, 16'd16144, 16'd61288, 16'd41437, 16'd57132, 16'd61065, 16'd52605, 16'd58483, 16'd59787, 16'd48599, 16'd30546, 16'd44480, 16'd49750});
	test_expansion(128'he0b0ca936087268ec016d7aad106cd8c, {16'd54311, 16'd32813, 16'd7938, 16'd21091, 16'd39435, 16'd23711, 16'd16554, 16'd37691, 16'd40585, 16'd41997, 16'd9531, 16'd50812, 16'd3289, 16'd23221, 16'd7791, 16'd50342, 16'd3857, 16'd37377, 16'd16301, 16'd39009, 16'd8558, 16'd64788, 16'd32177, 16'd37481, 16'd37109, 16'd11152});
	test_expansion(128'h21f0d1a8da598e4b9a43652f3cc443b7, {16'd25622, 16'd12796, 16'd59682, 16'd15351, 16'd59149, 16'd54447, 16'd20394, 16'd53765, 16'd17240, 16'd4232, 16'd23699, 16'd9189, 16'd40775, 16'd47434, 16'd27481, 16'd9658, 16'd37015, 16'd42228, 16'd14926, 16'd13650, 16'd34875, 16'd21294, 16'd37550, 16'd8260, 16'd54086, 16'd12120});
	test_expansion(128'hbba07d0feee9faf8523750f42933d67d, {16'd9003, 16'd32817, 16'd55935, 16'd56165, 16'd47209, 16'd38751, 16'd8352, 16'd58780, 16'd19800, 16'd61353, 16'd47127, 16'd7548, 16'd43543, 16'd18573, 16'd2620, 16'd58161, 16'd37112, 16'd26382, 16'd56050, 16'd54370, 16'd29122, 16'd62131, 16'd31693, 16'd1608, 16'd19983, 16'd23276});
	test_expansion(128'h568f4d6db535c410049906022a82e9e0, {16'd41028, 16'd39886, 16'd27354, 16'd37775, 16'd56964, 16'd48841, 16'd58728, 16'd56893, 16'd3369, 16'd7155, 16'd36350, 16'd43236, 16'd53700, 16'd46450, 16'd21526, 16'd54132, 16'd39845, 16'd60309, 16'd50222, 16'd14102, 16'd34438, 16'd36310, 16'd49786, 16'd54033, 16'd54374, 16'd27628});
	test_expansion(128'hfe9f435f780842530faa87f917357bd8, {16'd11465, 16'd35045, 16'd20652, 16'd8590, 16'd64872, 16'd8473, 16'd37860, 16'd13943, 16'd37475, 16'd63030, 16'd17889, 16'd60356, 16'd26331, 16'd10582, 16'd25369, 16'd35534, 16'd16921, 16'd3248, 16'd45882, 16'd5971, 16'd15343, 16'd64764, 16'd64123, 16'd35304, 16'd36020, 16'd23742});
	test_expansion(128'ha1145d41e81586f382f48cc6138b8602, {16'd46298, 16'd1606, 16'd28310, 16'd961, 16'd64131, 16'd51890, 16'd35272, 16'd17565, 16'd49, 16'd5991, 16'd31521, 16'd7309, 16'd32889, 16'd43347, 16'd38263, 16'd34686, 16'd59920, 16'd543, 16'd58392, 16'd45677, 16'd11108, 16'd37446, 16'd9354, 16'd26000, 16'd785, 16'd10799});
	test_expansion(128'h2418d224d0652bdfc223e06520a7a85d, {16'd59651, 16'd52474, 16'd63226, 16'd47420, 16'd56408, 16'd7875, 16'd65125, 16'd36270, 16'd34575, 16'd25115, 16'd50996, 16'd62102, 16'd31126, 16'd61106, 16'd7664, 16'd27319, 16'd65046, 16'd43326, 16'd50278, 16'd51835, 16'd6851, 16'd18696, 16'd51389, 16'd12367, 16'd10393, 16'd6728});
	test_expansion(128'hb56b4f9637c84bf9ca76dfed342b343a, {16'd8923, 16'd12386, 16'd3123, 16'd15259, 16'd41108, 16'd54340, 16'd12786, 16'd19547, 16'd25666, 16'd37873, 16'd60262, 16'd53387, 16'd58033, 16'd63917, 16'd32996, 16'd24751, 16'd60746, 16'd41785, 16'd30243, 16'd50113, 16'd4284, 16'd44382, 16'd18739, 16'd21355, 16'd62020, 16'd39667});
	test_expansion(128'h1ae44f0d201ef4d875347e9964fbc36c, {16'd11032, 16'd38367, 16'd17092, 16'd24709, 16'd42267, 16'd23342, 16'd29553, 16'd62677, 16'd42256, 16'd43997, 16'd42361, 16'd38874, 16'd35436, 16'd20741, 16'd27784, 16'd16417, 16'd33207, 16'd20991, 16'd28271, 16'd42025, 16'd32168, 16'd58290, 16'd31062, 16'd3590, 16'd44676, 16'd39368});
	test_expansion(128'h250764011734fbd3ca1ad514a37992f7, {16'd2859, 16'd13126, 16'd58750, 16'd1742, 16'd13760, 16'd61338, 16'd40976, 16'd28257, 16'd15249, 16'd5529, 16'd38963, 16'd25671, 16'd22076, 16'd23185, 16'd13221, 16'd18567, 16'd174, 16'd1734, 16'd53174, 16'd55028, 16'd52985, 16'd3999, 16'd61027, 16'd20692, 16'd9767, 16'd17158});
	test_expansion(128'hebe798ebcbd336123009294a02974274, {16'd1051, 16'd6362, 16'd22352, 16'd29883, 16'd17383, 16'd14083, 16'd32040, 16'd57351, 16'd44885, 16'd7155, 16'd16983, 16'd50562, 16'd20396, 16'd28765, 16'd2150, 16'd10152, 16'd5251, 16'd44702, 16'd6873, 16'd7504, 16'd787, 16'd56822, 16'd58223, 16'd60228, 16'd8016, 16'd15724});
	test_expansion(128'h4a9d29b5fb43d112ee47f8bd85b061aa, {16'd41206, 16'd41507, 16'd11497, 16'd36416, 16'd36123, 16'd48612, 16'd3799, 16'd4504, 16'd9944, 16'd8406, 16'd43393, 16'd41221, 16'd21741, 16'd26162, 16'd36152, 16'd20884, 16'd51788, 16'd51389, 16'd6924, 16'd33269, 16'd7405, 16'd59280, 16'd40791, 16'd38739, 16'd22691, 16'd16953});
	test_expansion(128'hc1bf5fe67b481f4cf35df8640516accc, {16'd54058, 16'd41094, 16'd14876, 16'd29561, 16'd20575, 16'd37904, 16'd12762, 16'd50003, 16'd9432, 16'd5563, 16'd22759, 16'd21324, 16'd41622, 16'd4999, 16'd46591, 16'd10898, 16'd28386, 16'd18217, 16'd48361, 16'd40689, 16'd44505, 16'd56185, 16'd55160, 16'd9903, 16'd11583, 16'd6183});
	test_expansion(128'hd17033c3cfffd6301e0302c76606b296, {16'd26447, 16'd14061, 16'd19326, 16'd49922, 16'd40247, 16'd3355, 16'd40264, 16'd13170, 16'd65385, 16'd8386, 16'd29055, 16'd51834, 16'd61850, 16'd64754, 16'd39193, 16'd56817, 16'd43911, 16'd47025, 16'd7802, 16'd15235, 16'd18718, 16'd62920, 16'd28255, 16'd40331, 16'd13982, 16'd45097});
	test_expansion(128'h10a9de9774a297584195d6c9c50ca084, {16'd1960, 16'd54217, 16'd65289, 16'd33391, 16'd16102, 16'd51846, 16'd22643, 16'd51477, 16'd39817, 16'd8637, 16'd43518, 16'd62729, 16'd19415, 16'd6388, 16'd26375, 16'd11429, 16'd41265, 16'd11004, 16'd54821, 16'd49095, 16'd9957, 16'd11218, 16'd29341, 16'd20468, 16'd48125, 16'd47985});
	test_expansion(128'h2b344e3e91c377dd4981e94878b599c6, {16'd41050, 16'd57412, 16'd31860, 16'd12611, 16'd60245, 16'd34431, 16'd58506, 16'd38502, 16'd38811, 16'd8162, 16'd62759, 16'd3415, 16'd48533, 16'd55145, 16'd25440, 16'd15298, 16'd54386, 16'd53793, 16'd35198, 16'd57518, 16'd36384, 16'd12770, 16'd17519, 16'd63210, 16'd42654, 16'd56936});
	test_expansion(128'h5ed234af912daa44357c153fbd3b4647, {16'd50627, 16'd2081, 16'd3651, 16'd27124, 16'd335, 16'd18693, 16'd6551, 16'd36978, 16'd55828, 16'd14000, 16'd4389, 16'd28130, 16'd4612, 16'd41459, 16'd61607, 16'd16346, 16'd20296, 16'd51416, 16'd48245, 16'd9321, 16'd50499, 16'd14995, 16'd62303, 16'd64064, 16'd28653, 16'd53699});
	test_expansion(128'h933132c43e5711379dfc0e83fbeb9838, {16'd9852, 16'd22532, 16'd3933, 16'd57517, 16'd61592, 16'd4658, 16'd347, 16'd29109, 16'd13699, 16'd30661, 16'd40629, 16'd10524, 16'd16404, 16'd23066, 16'd24686, 16'd17607, 16'd25816, 16'd11336, 16'd19706, 16'd39346, 16'd36968, 16'd21961, 16'd54586, 16'd60949, 16'd59522, 16'd61371});
	test_expansion(128'hee0007753c817e0cef338a2f0e4e6f33, {16'd27171, 16'd39586, 16'd11578, 16'd12286, 16'd47974, 16'd18554, 16'd32561, 16'd5835, 16'd35071, 16'd1133, 16'd52792, 16'd31306, 16'd5079, 16'd14374, 16'd60843, 16'd18534, 16'd62434, 16'd7361, 16'd13593, 16'd26512, 16'd31236, 16'd29856, 16'd60642, 16'd57870, 16'd45089, 16'd30953});
	test_expansion(128'hee34836895a8dbfe28048d0838d225c3, {16'd31679, 16'd32921, 16'd63489, 16'd26468, 16'd49558, 16'd48384, 16'd10133, 16'd17285, 16'd62891, 16'd16200, 16'd15910, 16'd39396, 16'd37199, 16'd1514, 16'd23038, 16'd49687, 16'd61672, 16'd973, 16'd24482, 16'd11028, 16'd52492, 16'd37454, 16'd33206, 16'd31268, 16'd1370, 16'd46440});
	test_expansion(128'h70faf814c853a1498b17cb8a9b08592b, {16'd28404, 16'd6866, 16'd61702, 16'd12828, 16'd13772, 16'd13799, 16'd45602, 16'd3026, 16'd3931, 16'd36378, 16'd18303, 16'd51588, 16'd40926, 16'd25200, 16'd3659, 16'd39183, 16'd43676, 16'd62992, 16'd33324, 16'd13587, 16'd54853, 16'd1546, 16'd19767, 16'd2643, 16'd5710, 16'd24179});
	test_expansion(128'he20f2f605bccd669f41cb0a5d45284d6, {16'd43477, 16'd45417, 16'd8626, 16'd9696, 16'd55355, 16'd33913, 16'd32030, 16'd6482, 16'd15126, 16'd7540, 16'd48984, 16'd30697, 16'd54787, 16'd42064, 16'd61793, 16'd47851, 16'd59477, 16'd2264, 16'd59810, 16'd55065, 16'd12086, 16'd58008, 16'd33239, 16'd22110, 16'd25198, 16'd15570});
	test_expansion(128'h15160d900b51b4d117adcd85de905490, {16'd12797, 16'd43298, 16'd18943, 16'd4875, 16'd14295, 16'd43324, 16'd11867, 16'd25843, 16'd36766, 16'd38328, 16'd8736, 16'd26569, 16'd63614, 16'd3688, 16'd6913, 16'd25572, 16'd48870, 16'd2222, 16'd29192, 16'd2937, 16'd39407, 16'd37043, 16'd54080, 16'd56055, 16'd39025, 16'd44834});
	test_expansion(128'h3b9e75a7a94be4c00addf840bc8e4985, {16'd63455, 16'd15125, 16'd58229, 16'd24248, 16'd54217, 16'd40190, 16'd6669, 16'd17077, 16'd36120, 16'd59220, 16'd18344, 16'd6334, 16'd34323, 16'd24640, 16'd43316, 16'd7375, 16'd19813, 16'd33658, 16'd34222, 16'd42865, 16'd48213, 16'd46311, 16'd64874, 16'd46080, 16'd52950, 16'd62978});
	test_expansion(128'h0a23ab984b94ec87dcf5778134a2c10b, {16'd28449, 16'd10301, 16'd51518, 16'd62443, 16'd40439, 16'd49786, 16'd65423, 16'd15983, 16'd19526, 16'd7862, 16'd33372, 16'd47329, 16'd53811, 16'd18015, 16'd15882, 16'd3823, 16'd44697, 16'd52440, 16'd47199, 16'd31230, 16'd25795, 16'd39759, 16'd10755, 16'd10521, 16'd18599, 16'd60011});
	test_expansion(128'h1da9eba193387204f8d73bab210ef670, {16'd61083, 16'd38935, 16'd15903, 16'd23444, 16'd5715, 16'd34895, 16'd25256, 16'd45983, 16'd1824, 16'd8944, 16'd5462, 16'd27673, 16'd57248, 16'd34778, 16'd40977, 16'd7129, 16'd37665, 16'd7457, 16'd24193, 16'd38085, 16'd55436, 16'd54625, 16'd19892, 16'd56973, 16'd50968, 16'd6540});
	test_expansion(128'hbbb3b7f17bf9fca877ed2e27964700eb, {16'd5888, 16'd4159, 16'd41321, 16'd1280, 16'd15198, 16'd19666, 16'd57530, 16'd27791, 16'd64240, 16'd14987, 16'd1398, 16'd59799, 16'd32433, 16'd7618, 16'd12967, 16'd48790, 16'd51379, 16'd63857, 16'd8044, 16'd21637, 16'd26712, 16'd38324, 16'd42423, 16'd39404, 16'd37915, 16'd50276});
	test_expansion(128'hf83354d7b65cb34cfb120a35ae512238, {16'd37225, 16'd11931, 16'd34227, 16'd6157, 16'd47878, 16'd51447, 16'd57720, 16'd60315, 16'd30111, 16'd59752, 16'd51807, 16'd19310, 16'd17537, 16'd47087, 16'd43359, 16'd1450, 16'd49807, 16'd24265, 16'd56108, 16'd50546, 16'd42585, 16'd8818, 16'd19998, 16'd15697, 16'd31678, 16'd27300});
	test_expansion(128'hb08502d70be4bb6181896fd67984adf4, {16'd53401, 16'd53230, 16'd61620, 16'd10524, 16'd34911, 16'd59048, 16'd6242, 16'd35683, 16'd56283, 16'd25185, 16'd5245, 16'd28633, 16'd2657, 16'd4847, 16'd10940, 16'd22729, 16'd24906, 16'd2703, 16'd24905, 16'd50586, 16'd35625, 16'd16444, 16'd14057, 16'd36782, 16'd23251, 16'd28945});
	test_expansion(128'h08925d274e6b5434f4be11d462130331, {16'd36332, 16'd22224, 16'd41787, 16'd8622, 16'd4531, 16'd48207, 16'd44646, 16'd8784, 16'd55686, 16'd14921, 16'd62758, 16'd51534, 16'd2603, 16'd1753, 16'd21107, 16'd7915, 16'd54852, 16'd57259, 16'd21729, 16'd36090, 16'd17170, 16'd62859, 16'd56401, 16'd64036, 16'd13920, 16'd40345});
	test_expansion(128'h9c8d3989eb134cbc7c8d1bd2ed3402ea, {16'd49669, 16'd34004, 16'd5022, 16'd29565, 16'd36409, 16'd48401, 16'd33878, 16'd56413, 16'd45880, 16'd61086, 16'd43455, 16'd42368, 16'd20430, 16'd45744, 16'd63034, 16'd43625, 16'd56220, 16'd63248, 16'd41688, 16'd2020, 16'd40663, 16'd5603, 16'd10527, 16'd37326, 16'd63398, 16'd3245});
	test_expansion(128'hdbf5b12e7ff7eee8f164e0a5c9ddf68a, {16'd28958, 16'd10522, 16'd62590, 16'd57590, 16'd33456, 16'd45774, 16'd11378, 16'd2084, 16'd3297, 16'd56124, 16'd45824, 16'd50175, 16'd4313, 16'd56483, 16'd13812, 16'd55990, 16'd18330, 16'd27261, 16'd37135, 16'd22063, 16'd63737, 16'd33309, 16'd30737, 16'd19279, 16'd13868, 16'd37914});
	test_expansion(128'h3bcec4a451c61370794c77185f48d582, {16'd58362, 16'd9170, 16'd4384, 16'd57384, 16'd45347, 16'd7388, 16'd29395, 16'd49861, 16'd11288, 16'd6766, 16'd17576, 16'd24550, 16'd20, 16'd2282, 16'd57254, 16'd47989, 16'd52769, 16'd27297, 16'd24745, 16'd63405, 16'd44934, 16'd21993, 16'd63570, 16'd16274, 16'd50297, 16'd31480});
	test_expansion(128'h88d24254baaed34c0b6679d5dec81556, {16'd31083, 16'd61225, 16'd31911, 16'd57447, 16'd62528, 16'd7001, 16'd16948, 16'd54073, 16'd54409, 16'd37949, 16'd53586, 16'd36551, 16'd35976, 16'd24367, 16'd42269, 16'd32380, 16'd39990, 16'd41899, 16'd17174, 16'd35586, 16'd65204, 16'd51415, 16'd8853, 16'd10850, 16'd45523, 16'd15881});
	test_expansion(128'h3181b2baeca2895f809efb70a34a79d7, {16'd52889, 16'd55049, 16'd45344, 16'd20993, 16'd47992, 16'd36930, 16'd33251, 16'd36778, 16'd43542, 16'd336, 16'd53757, 16'd47427, 16'd22699, 16'd52622, 16'd4952, 16'd34126, 16'd60122, 16'd54006, 16'd15467, 16'd8958, 16'd64872, 16'd5433, 16'd56913, 16'd24107, 16'd4231, 16'd3962});
	test_expansion(128'hec38f7ad3778ce9ae2b54718f13e1cc0, {16'd17876, 16'd6749, 16'd12906, 16'd45083, 16'd58286, 16'd11728, 16'd54959, 16'd36127, 16'd16472, 16'd24556, 16'd4277, 16'd50498, 16'd52912, 16'd19156, 16'd506, 16'd23759, 16'd43016, 16'd24791, 16'd3430, 16'd15322, 16'd49323, 16'd21908, 16'd35897, 16'd48828, 16'd65218, 16'd52917});
	test_expansion(128'hefe6bab71f5afa23cf78f92150918824, {16'd36365, 16'd46768, 16'd32668, 16'd60291, 16'd10972, 16'd28623, 16'd56748, 16'd42481, 16'd58279, 16'd28706, 16'd9554, 16'd1700, 16'd8698, 16'd63973, 16'd30363, 16'd24439, 16'd19960, 16'd20630, 16'd47071, 16'd11519, 16'd57122, 16'd15641, 16'd30578, 16'd8610, 16'd57234, 16'd52507});
	test_expansion(128'h60167608f03e0099281c4dd0f9a475f5, {16'd27448, 16'd56252, 16'd61506, 16'd32146, 16'd29361, 16'd63799, 16'd2698, 16'd52076, 16'd19395, 16'd21502, 16'd7380, 16'd62836, 16'd34010, 16'd25729, 16'd4316, 16'd18228, 16'd30598, 16'd15483, 16'd1411, 16'd10522, 16'd62951, 16'd31724, 16'd46128, 16'd3843, 16'd20660, 16'd25015});
	test_expansion(128'h028caff7498dca07034e192468d9a9dd, {16'd14895, 16'd57023, 16'd42379, 16'd735, 16'd6126, 16'd8343, 16'd59714, 16'd1521, 16'd26382, 16'd25422, 16'd10955, 16'd22566, 16'd19951, 16'd59407, 16'd47705, 16'd15878, 16'd37472, 16'd60528, 16'd5375, 16'd22016, 16'd29777, 16'd47822, 16'd19874, 16'd10118, 16'd11444, 16'd37493});
	test_expansion(128'hd9c0776f725158831e5aff10325d61a1, {16'd26898, 16'd62038, 16'd25402, 16'd57258, 16'd41438, 16'd21609, 16'd8404, 16'd52263, 16'd8827, 16'd64409, 16'd32932, 16'd60986, 16'd20223, 16'd17092, 16'd56937, 16'd47908, 16'd23301, 16'd5109, 16'd48772, 16'd16420, 16'd44593, 16'd10324, 16'd17443, 16'd21099, 16'd20246, 16'd25500});
	test_expansion(128'hdaa981ae48597c099fd03ea822d032a5, {16'd45040, 16'd58194, 16'd5667, 16'd54818, 16'd20528, 16'd10022, 16'd60341, 16'd12484, 16'd17356, 16'd57586, 16'd59739, 16'd47341, 16'd54425, 16'd36731, 16'd60847, 16'd11390, 16'd40486, 16'd21989, 16'd52038, 16'd17286, 16'd17021, 16'd7372, 16'd50498, 16'd60813, 16'd49310, 16'd6545});
	test_expansion(128'h70dd355f2e114aa275f25824643418fd, {16'd14192, 16'd4519, 16'd5191, 16'd3731, 16'd41337, 16'd15467, 16'd56034, 16'd60993, 16'd57214, 16'd28916, 16'd49343, 16'd23152, 16'd34533, 16'd49997, 16'd8622, 16'd36222, 16'd9363, 16'd18889, 16'd47253, 16'd61499, 16'd12302, 16'd13341, 16'd38928, 16'd10214, 16'd32514, 16'd41538});
	test_expansion(128'h9f7fffcd243ac4363ec59e2fe82cb2d6, {16'd11690, 16'd17082, 16'd62080, 16'd57455, 16'd55899, 16'd8104, 16'd2109, 16'd24123, 16'd12063, 16'd48997, 16'd409, 16'd17351, 16'd55335, 16'd32424, 16'd5028, 16'd4229, 16'd16748, 16'd50533, 16'd22027, 16'd59408, 16'd8129, 16'd30487, 16'd51789, 16'd14327, 16'd29508, 16'd8462});
	test_expansion(128'h431e3a8dfd4c5fa54e0d62890cff2a21, {16'd20676, 16'd22801, 16'd63807, 16'd13699, 16'd28857, 16'd41766, 16'd139, 16'd7900, 16'd59918, 16'd14222, 16'd15358, 16'd55945, 16'd30516, 16'd65169, 16'd63465, 16'd10058, 16'd49772, 16'd19841, 16'd13946, 16'd38170, 16'd7825, 16'd57638, 16'd59716, 16'd41089, 16'd61606, 16'd23435});
	test_expansion(128'heb130802f750c946f2fcf2f572fe3b97, {16'd55827, 16'd46221, 16'd44310, 16'd56580, 16'd8182, 16'd27520, 16'd54770, 16'd31553, 16'd55694, 16'd22157, 16'd17344, 16'd23170, 16'd518, 16'd25761, 16'd55616, 16'd37625, 16'd7910, 16'd48234, 16'd22464, 16'd23230, 16'd45189, 16'd61931, 16'd21983, 16'd20286, 16'd32288, 16'd27910});
	test_expansion(128'h7c706059d325d74ed95d5f4b297fe709, {16'd15701, 16'd12449, 16'd12433, 16'd41618, 16'd11083, 16'd23507, 16'd2552, 16'd3955, 16'd40282, 16'd4206, 16'd31526, 16'd58742, 16'd64153, 16'd45375, 16'd9303, 16'd7301, 16'd40194, 16'd55069, 16'd13320, 16'd8658, 16'd14718, 16'd26506, 16'd61117, 16'd22890, 16'd49437, 16'd62774});
	test_expansion(128'h16df2063a81029ba01f4ea5f3602a782, {16'd50941, 16'd50443, 16'd5305, 16'd9604, 16'd38137, 16'd7107, 16'd49057, 16'd41529, 16'd35112, 16'd17732, 16'd3, 16'd48254, 16'd8259, 16'd11106, 16'd42994, 16'd4965, 16'd4270, 16'd33972, 16'd39865, 16'd4197, 16'd29647, 16'd9851, 16'd64259, 16'd29930, 16'd2248, 16'd21465});
	test_expansion(128'h3b43e961942aef00121f97b962e26839, {16'd42833, 16'd10615, 16'd52224, 16'd25438, 16'd41271, 16'd43842, 16'd33902, 16'd31890, 16'd40547, 16'd49390, 16'd8448, 16'd56550, 16'd9697, 16'd8265, 16'd58690, 16'd36167, 16'd42891, 16'd52154, 16'd41160, 16'd37880, 16'd27683, 16'd7066, 16'd19886, 16'd22424, 16'd7716, 16'd37873});
	test_expansion(128'hc73c80f4a938dd896b0f968db2686594, {16'd46039, 16'd64567, 16'd33522, 16'd38816, 16'd51961, 16'd32732, 16'd24511, 16'd193, 16'd44201, 16'd20830, 16'd24517, 16'd35893, 16'd29801, 16'd24648, 16'd3240, 16'd59074, 16'd48542, 16'd54839, 16'd47072, 16'd40185, 16'd57213, 16'd31158, 16'd27923, 16'd2866, 16'd19913, 16'd62616});
	test_expansion(128'h20ec957e5641384e290a47bfbfc7906e, {16'd43941, 16'd28764, 16'd10287, 16'd4662, 16'd44857, 16'd47081, 16'd15091, 16'd36614, 16'd2601, 16'd7139, 16'd17273, 16'd19314, 16'd43162, 16'd54956, 16'd21283, 16'd34400, 16'd3709, 16'd31178, 16'd23747, 16'd1124, 16'd42813, 16'd40929, 16'd7309, 16'd36712, 16'd57309, 16'd2102});
	test_expansion(128'hfee7ed4ddb26379d0b88cdf4e2fcfa20, {16'd51179, 16'd8807, 16'd30347, 16'd31732, 16'd14053, 16'd46061, 16'd35967, 16'd40687, 16'd39042, 16'd35628, 16'd52383, 16'd8969, 16'd59079, 16'd63211, 16'd407, 16'd43707, 16'd26530, 16'd55120, 16'd58058, 16'd7095, 16'd49973, 16'd56991, 16'd9027, 16'd49270, 16'd37071, 16'd13002});
	test_expansion(128'h6d9e8fa50f8a8ddda2c54317f290140c, {16'd10588, 16'd31247, 16'd33523, 16'd1038, 16'd21194, 16'd20294, 16'd4168, 16'd39575, 16'd34818, 16'd55687, 16'd41763, 16'd3609, 16'd25071, 16'd10121, 16'd37128, 16'd4703, 16'd1107, 16'd46069, 16'd28713, 16'd36756, 16'd56678, 16'd20203, 16'd15762, 16'd3590, 16'd10899, 16'd39964});
	test_expansion(128'h63e6f751bb8096ed3893c26c354460ce, {16'd57139, 16'd60719, 16'd60824, 16'd34657, 16'd19634, 16'd65124, 16'd8745, 16'd60519, 16'd12288, 16'd54445, 16'd52844, 16'd27416, 16'd22687, 16'd63242, 16'd4243, 16'd43916, 16'd36506, 16'd53047, 16'd40544, 16'd4650, 16'd10937, 16'd8649, 16'd41814, 16'd28085, 16'd61929, 16'd37793});
	test_expansion(128'h35826eab5338c10a9797188ea3067e68, {16'd20442, 16'd23170, 16'd26612, 16'd31629, 16'd57196, 16'd37043, 16'd37181, 16'd55053, 16'd60012, 16'd26351, 16'd29662, 16'd58423, 16'd55648, 16'd26943, 16'd50376, 16'd3161, 16'd39443, 16'd20330, 16'd46178, 16'd10757, 16'd23042, 16'd50510, 16'd61202, 16'd17840, 16'd63714, 16'd45610});
	test_expansion(128'h563e2c173ddbc83d1e1a93046ffabffb, {16'd31996, 16'd61939, 16'd60363, 16'd55131, 16'd3977, 16'd46674, 16'd7045, 16'd14582, 16'd17265, 16'd27876, 16'd10363, 16'd32133, 16'd41278, 16'd7740, 16'd13639, 16'd31945, 16'd9446, 16'd2850, 16'd29491, 16'd22738, 16'd3942, 16'd10261, 16'd29143, 16'd11937, 16'd58084, 16'd52424});
	test_expansion(128'hdc4043dd7bfe884bd252112b001cce0f, {16'd14540, 16'd42741, 16'd12112, 16'd58065, 16'd39371, 16'd43586, 16'd627, 16'd20457, 16'd41620, 16'd18846, 16'd5595, 16'd29620, 16'd21605, 16'd44032, 16'd49553, 16'd34565, 16'd10850, 16'd44542, 16'd45164, 16'd52651, 16'd48492, 16'd44418, 16'd64345, 16'd1702, 16'd44262, 16'd44639});
	test_expansion(128'ha66cb10954aa38c335baf6496a9f9299, {16'd34977, 16'd3556, 16'd47301, 16'd38493, 16'd28512, 16'd57793, 16'd41730, 16'd29906, 16'd46658, 16'd33456, 16'd39548, 16'd12249, 16'd7188, 16'd896, 16'd61173, 16'd59306, 16'd59504, 16'd61304, 16'd35249, 16'd34023, 16'd56453, 16'd59128, 16'd59716, 16'd61402, 16'd53868, 16'd61186});
	test_expansion(128'h56a3536430d5090cfff808157f1248b7, {16'd61996, 16'd32903, 16'd14445, 16'd14330, 16'd61397, 16'd40058, 16'd58575, 16'd5557, 16'd61336, 16'd25855, 16'd30404, 16'd31943, 16'd6057, 16'd49874, 16'd23165, 16'd38496, 16'd5921, 16'd17243, 16'd61533, 16'd63883, 16'd44360, 16'd24484, 16'd33579, 16'd34464, 16'd9383, 16'd58614});
	test_expansion(128'h532c554febc0a2e35d6a53ed6d76b0d3, {16'd22325, 16'd8663, 16'd20917, 16'd65219, 16'd46209, 16'd3307, 16'd1680, 16'd2881, 16'd27980, 16'd7243, 16'd26234, 16'd52252, 16'd57804, 16'd39648, 16'd24296, 16'd12794, 16'd53679, 16'd37336, 16'd18565, 16'd23152, 16'd44315, 16'd15626, 16'd38505, 16'd50559, 16'd7948, 16'd45575});
	test_expansion(128'h4c8b5ba9e56304586d019760db4ecf9c, {16'd10475, 16'd65013, 16'd28024, 16'd28922, 16'd21272, 16'd17219, 16'd43274, 16'd58225, 16'd16870, 16'd48795, 16'd31643, 16'd25241, 16'd65059, 16'd55538, 16'd40463, 16'd52288, 16'd31452, 16'd12664, 16'd28683, 16'd23393, 16'd39280, 16'd51118, 16'd7162, 16'd22501, 16'd30477, 16'd26967});
	test_expansion(128'h4d82cd020e9df3f69c90a006f46434aa, {16'd39947, 16'd10154, 16'd28707, 16'd48486, 16'd11440, 16'd21098, 16'd55036, 16'd5344, 16'd1648, 16'd62303, 16'd5301, 16'd9122, 16'd16175, 16'd23473, 16'd27804, 16'd7295, 16'd54157, 16'd60487, 16'd51540, 16'd31068, 16'd32737, 16'd56620, 16'd4926, 16'd51154, 16'd23757, 16'd6770});
	test_expansion(128'h7525eab2e1a6dfb320070e93bd82ac3e, {16'd1287, 16'd7768, 16'd3676, 16'd34974, 16'd13911, 16'd1672, 16'd29500, 16'd51947, 16'd12832, 16'd55785, 16'd18787, 16'd9221, 16'd65286, 16'd57224, 16'd64990, 16'd2374, 16'd29397, 16'd782, 16'd4665, 16'd16636, 16'd2914, 16'd26376, 16'd44944, 16'd2073, 16'd8714, 16'd60054});
	test_expansion(128'h9afeecc42279e2f6381b98b6b5c96dcf, {16'd36418, 16'd37722, 16'd27347, 16'd4748, 16'd27918, 16'd5089, 16'd12817, 16'd11668, 16'd5931, 16'd31596, 16'd59626, 16'd20091, 16'd190, 16'd9963, 16'd54884, 16'd34079, 16'd38665, 16'd1966, 16'd23321, 16'd30277, 16'd7441, 16'd8139, 16'd47708, 16'd51200, 16'd28800, 16'd39668});
	test_expansion(128'h23998030d21fb4f1c10dc13c810f555e, {16'd10038, 16'd5298, 16'd22252, 16'd17132, 16'd1045, 16'd43018, 16'd27932, 16'd2605, 16'd50610, 16'd1714, 16'd1002, 16'd43393, 16'd13810, 16'd11894, 16'd46044, 16'd9565, 16'd5411, 16'd7135, 16'd51501, 16'd24175, 16'd16502, 16'd28957, 16'd39679, 16'd51543, 16'd42726, 16'd45500});
	test_expansion(128'hc3976601c1e796798b86325cceb72584, {16'd60340, 16'd25122, 16'd65135, 16'd17531, 16'd58748, 16'd54698, 16'd35671, 16'd48835, 16'd46025, 16'd28690, 16'd28163, 16'd9578, 16'd17470, 16'd37364, 16'd63882, 16'd63056, 16'd55235, 16'd2674, 16'd17275, 16'd58330, 16'd10881, 16'd15786, 16'd63606, 16'd42685, 16'd59331, 16'd49259});
	test_expansion(128'hae2f8b09d91bf54c21821ff5e4bb0875, {16'd24600, 16'd12471, 16'd64762, 16'd39038, 16'd11293, 16'd27857, 16'd32551, 16'd36753, 16'd41076, 16'd57787, 16'd2822, 16'd21304, 16'd45344, 16'd48544, 16'd16022, 16'd17966, 16'd39542, 16'd32754, 16'd48490, 16'd28228, 16'd3277, 16'd8092, 16'd49604, 16'd59482, 16'd60671, 16'd57684});
	test_expansion(128'h392658b91e85a87eda54dcbace5e1385, {16'd64189, 16'd31597, 16'd60793, 16'd33889, 16'd61283, 16'd45277, 16'd29673, 16'd4704, 16'd23564, 16'd63522, 16'd2419, 16'd8213, 16'd24120, 16'd15179, 16'd53976, 16'd64152, 16'd33262, 16'd43205, 16'd60919, 16'd24715, 16'd50035, 16'd57759, 16'd20122, 16'd29979, 16'd4819, 16'd48654});
	test_expansion(128'h0ae4791a0803c329416db0a1b4ac0570, {16'd48006, 16'd8243, 16'd35736, 16'd36625, 16'd20125, 16'd12287, 16'd20515, 16'd38991, 16'd7001, 16'd7562, 16'd41206, 16'd9543, 16'd49463, 16'd12719, 16'd30565, 16'd1621, 16'd53023, 16'd13198, 16'd55969, 16'd11314, 16'd43658, 16'd41694, 16'd57915, 16'd24391, 16'd25126, 16'd17859});
	test_expansion(128'h941cf29fb46baba42e5e2187120c15e1, {16'd37326, 16'd24331, 16'd46409, 16'd25753, 16'd51615, 16'd60566, 16'd57935, 16'd6824, 16'd30809, 16'd9961, 16'd7208, 16'd12578, 16'd38092, 16'd1973, 16'd11024, 16'd41213, 16'd39089, 16'd63683, 16'd40051, 16'd5546, 16'd46161, 16'd26406, 16'd51804, 16'd29763, 16'd1502, 16'd63933});
	test_expansion(128'h1d655296adbd415d0fa99fc1b72609e0, {16'd16676, 16'd26593, 16'd14201, 16'd14942, 16'd62176, 16'd4636, 16'd24492, 16'd41560, 16'd61493, 16'd63834, 16'd53190, 16'd49221, 16'd60980, 16'd63141, 16'd59632, 16'd7272, 16'd52308, 16'd34695, 16'd18342, 16'd25122, 16'd4710, 16'd29458, 16'd45347, 16'd39276, 16'd28890, 16'd29653});
	test_expansion(128'h4e712c3d03a70a99a7507be4e9c22550, {16'd7888, 16'd45871, 16'd29313, 16'd18071, 16'd7934, 16'd45217, 16'd58796, 16'd18678, 16'd23059, 16'd3130, 16'd14162, 16'd11583, 16'd37033, 16'd63215, 16'd53052, 16'd61203, 16'd3511, 16'd23560, 16'd49111, 16'd7251, 16'd11916, 16'd27782, 16'd1793, 16'd56689, 16'd36150, 16'd10285});
	test_expansion(128'h3b8dd4d86ca8ecc6636e9bc649d5e95a, {16'd7836, 16'd5291, 16'd4065, 16'd29653, 16'd8602, 16'd33752, 16'd55782, 16'd12010, 16'd6896, 16'd15359, 16'd57825, 16'd51411, 16'd5842, 16'd35998, 16'd52883, 16'd63717, 16'd60868, 16'd22137, 16'd14964, 16'd21095, 16'd22230, 16'd13477, 16'd19666, 16'd630, 16'd35196, 16'd28840});
	test_expansion(128'h400296b18d639809f7fa6325dad238db, {16'd58027, 16'd22015, 16'd7134, 16'd26253, 16'd38909, 16'd5303, 16'd10042, 16'd2224, 16'd12635, 16'd12686, 16'd26444, 16'd27394, 16'd61102, 16'd47003, 16'd37120, 16'd408, 16'd13521, 16'd21363, 16'd34236, 16'd31397, 16'd32507, 16'd12985, 16'd38158, 16'd31570, 16'd39429, 16'd25367});
	test_expansion(128'h05d53547815cf0946031b5f29d0d6615, {16'd18641, 16'd46867, 16'd56468, 16'd52648, 16'd1097, 16'd20303, 16'd48850, 16'd22486, 16'd14711, 16'd9196, 16'd45431, 16'd23519, 16'd30617, 16'd48040, 16'd16104, 16'd10974, 16'd53763, 16'd29929, 16'd53921, 16'd57040, 16'd35776, 16'd54260, 16'd26333, 16'd10661, 16'd48687, 16'd36350});
	test_expansion(128'h80bbbd204936a3fa49a94b35f726572b, {16'd29484, 16'd52658, 16'd2457, 16'd61660, 16'd16241, 16'd63210, 16'd7514, 16'd53697, 16'd14319, 16'd65128, 16'd29706, 16'd32112, 16'd16105, 16'd32045, 16'd41418, 16'd24514, 16'd11943, 16'd16243, 16'd16444, 16'd54613, 16'd49751, 16'd3546, 16'd56119, 16'd59872, 16'd49176, 16'd18043});
	test_expansion(128'h8dc654bd8b9c44e44d99d5542fd1a313, {16'd47851, 16'd9170, 16'd28088, 16'd61658, 16'd57752, 16'd38546, 16'd27132, 16'd40715, 16'd50121, 16'd65171, 16'd23747, 16'd34768, 16'd931, 16'd14038, 16'd1092, 16'd1513, 16'd40233, 16'd40802, 16'd27743, 16'd61215, 16'd5064, 16'd8885, 16'd64387, 16'd35621, 16'd10013, 16'd26694});
	test_expansion(128'h9300ed4a773186f5d8afbd2f71ca45a9, {16'd28122, 16'd50747, 16'd29175, 16'd7035, 16'd1316, 16'd4105, 16'd26946, 16'd4704, 16'd29199, 16'd38390, 16'd37317, 16'd18978, 16'd7599, 16'd7742, 16'd32538, 16'd11516, 16'd58741, 16'd61948, 16'd37662, 16'd40806, 16'd62539, 16'd53170, 16'd56371, 16'd45624, 16'd25784, 16'd34742});
	test_expansion(128'h545af67d1e3b81076a9085e3cb733460, {16'd64997, 16'd8249, 16'd50521, 16'd20660, 16'd19706, 16'd45370, 16'd2152, 16'd504, 16'd1144, 16'd34855, 16'd27938, 16'd24972, 16'd3313, 16'd46865, 16'd15739, 16'd33339, 16'd42791, 16'd16973, 16'd11779, 16'd46811, 16'd35015, 16'd30778, 16'd41957, 16'd23611, 16'd22452, 16'd43157});
	test_expansion(128'h4a6c19edee9ccd79924458367c473249, {16'd31909, 16'd2806, 16'd19388, 16'd47566, 16'd5436, 16'd55917, 16'd63692, 16'd14409, 16'd49612, 16'd7559, 16'd2315, 16'd6219, 16'd41995, 16'd39409, 16'd19289, 16'd31103, 16'd18658, 16'd51624, 16'd43192, 16'd45103, 16'd65283, 16'd48403, 16'd12007, 16'd17735, 16'd10951, 16'd20976});
	test_expansion(128'hf33d8a84ebb2fce8ae40a1bc6ed9e9b0, {16'd4038, 16'd39841, 16'd45397, 16'd21981, 16'd28199, 16'd31078, 16'd30042, 16'd32150, 16'd38420, 16'd64875, 16'd25876, 16'd23346, 16'd38895, 16'd45386, 16'd18859, 16'd6827, 16'd26603, 16'd24984, 16'd50866, 16'd62141, 16'd19158, 16'd62642, 16'd50317, 16'd4995, 16'd10462, 16'd7935});
	test_expansion(128'hb052b5945a2a06b4306717622f0c6a76, {16'd42198, 16'd44122, 16'd58900, 16'd36021, 16'd36492, 16'd38396, 16'd59738, 16'd26060, 16'd4763, 16'd28560, 16'd25294, 16'd42070, 16'd53942, 16'd58672, 16'd8206, 16'd23567, 16'd48392, 16'd36039, 16'd57508, 16'd10986, 16'd25964, 16'd49175, 16'd46654, 16'd64319, 16'd61887, 16'd4194});
	test_expansion(128'hfd6d51e6667f390e281db6c3a7a29285, {16'd35881, 16'd625, 16'd20406, 16'd12054, 16'd17197, 16'd50426, 16'd16312, 16'd54145, 16'd57955, 16'd1327, 16'd23106, 16'd44898, 16'd14304, 16'd41745, 16'd51797, 16'd13581, 16'd10431, 16'd20998, 16'd21916, 16'd27987, 16'd60947, 16'd33807, 16'd61862, 16'd9881, 16'd5487, 16'd56165});
	test_expansion(128'h1fd886b777e02df2a231d03695b844ea, {16'd27847, 16'd56279, 16'd15095, 16'd15352, 16'd64996, 16'd57794, 16'd23855, 16'd58641, 16'd25969, 16'd12179, 16'd44609, 16'd17007, 16'd13195, 16'd42699, 16'd17837, 16'd18390, 16'd47545, 16'd29633, 16'd41247, 16'd51415, 16'd4596, 16'd33977, 16'd59975, 16'd53099, 16'd45710, 16'd27874});
	test_expansion(128'hcdafac03b591383e6219744bc32da71d, {16'd27590, 16'd63922, 16'd59868, 16'd12717, 16'd33481, 16'd54255, 16'd40828, 16'd10926, 16'd28671, 16'd39070, 16'd31932, 16'd11694, 16'd32206, 16'd9094, 16'd38500, 16'd43098, 16'd56246, 16'd44202, 16'd10407, 16'd22457, 16'd7981, 16'd39595, 16'd61191, 16'd38346, 16'd15223, 16'd31918});
	test_expansion(128'he14fcb2b73ae66179a01f76a8a4f96b5, {16'd19234, 16'd52337, 16'd18794, 16'd48588, 16'd63956, 16'd24450, 16'd44202, 16'd65194, 16'd57147, 16'd33660, 16'd34219, 16'd47397, 16'd2674, 16'd17406, 16'd3639, 16'd23779, 16'd9439, 16'd48697, 16'd19223, 16'd63607, 16'd42048, 16'd26704, 16'd49169, 16'd47977, 16'd28857, 16'd37493});
	test_expansion(128'ha1574015bb65026cbffce3729d5c7419, {16'd20699, 16'd26614, 16'd47584, 16'd62288, 16'd13304, 16'd14901, 16'd34738, 16'd36754, 16'd8503, 16'd56633, 16'd58191, 16'd9358, 16'd29799, 16'd49686, 16'd31205, 16'd25986, 16'd34619, 16'd35345, 16'd63920, 16'd19534, 16'd26273, 16'd44389, 16'd35891, 16'd3541, 16'd62076, 16'd2871});
	test_expansion(128'had2331c2770a56c4ab70db9642fbfe57, {16'd52873, 16'd5820, 16'd8031, 16'd6295, 16'd19891, 16'd22884, 16'd46256, 16'd49884, 16'd50217, 16'd20796, 16'd28986, 16'd13927, 16'd44479, 16'd54484, 16'd46234, 16'd32970, 16'd25352, 16'd60846, 16'd45047, 16'd13172, 16'd14291, 16'd38691, 16'd24771, 16'd44983, 16'd48845, 16'd46784});
	test_expansion(128'h78ccaa54112536dc768016880042cbe7, {16'd49619, 16'd21553, 16'd26755, 16'd35182, 16'd2860, 16'd12736, 16'd55798, 16'd1200, 16'd29748, 16'd20092, 16'd32735, 16'd6043, 16'd57148, 16'd12425, 16'd61301, 16'd5373, 16'd11695, 16'd61110, 16'd5920, 16'd6755, 16'd56959, 16'd56336, 16'd30744, 16'd46582, 16'd17557, 16'd8928});
	test_expansion(128'h89af408dd4dd16f7f03e2fadf5d7079a, {16'd54681, 16'd43983, 16'd57942, 16'd7529, 16'd31819, 16'd50515, 16'd61213, 16'd7518, 16'd2106, 16'd60671, 16'd62439, 16'd32554, 16'd20753, 16'd21743, 16'd9418, 16'd22341, 16'd53760, 16'd25202, 16'd23213, 16'd50933, 16'd25597, 16'd35998, 16'd30357, 16'd205, 16'd29456, 16'd4088});
	test_expansion(128'hce31035f2418bda8a950f89cfb50a56d, {16'd5597, 16'd60044, 16'd36660, 16'd53247, 16'd62572, 16'd57936, 16'd30910, 16'd2228, 16'd5508, 16'd10881, 16'd20801, 16'd1021, 16'd25350, 16'd37224, 16'd52174, 16'd35242, 16'd2552, 16'd36239, 16'd35838, 16'd42880, 16'd64283, 16'd28441, 16'd5635, 16'd53505, 16'd16744, 16'd16934});
	test_expansion(128'h414fdca62750f2cb94c6fd5755ddc36a, {16'd62256, 16'd37780, 16'd39458, 16'd1634, 16'd27775, 16'd4373, 16'd55519, 16'd35869, 16'd60401, 16'd51649, 16'd39361, 16'd65295, 16'd60327, 16'd27978, 16'd16655, 16'd13036, 16'd8505, 16'd8594, 16'd39698, 16'd64328, 16'd34773, 16'd16260, 16'd52303, 16'd13414, 16'd55255, 16'd7390});
	test_expansion(128'hf5d47f0371a055b9a8f114a685f4da52, {16'd63480, 16'd21314, 16'd47755, 16'd25452, 16'd26269, 16'd40436, 16'd27862, 16'd24816, 16'd10715, 16'd25236, 16'd10029, 16'd22507, 16'd12681, 16'd26920, 16'd2440, 16'd53279, 16'd20840, 16'd7960, 16'd63744, 16'd10610, 16'd15114, 16'd28153, 16'd23440, 16'd4621, 16'd6012, 16'd9669});
	test_expansion(128'hb0f6b3caa8d0f56267422fca5bc503a0, {16'd64517, 16'd33586, 16'd50746, 16'd29129, 16'd14556, 16'd61508, 16'd29792, 16'd23848, 16'd55730, 16'd4606, 16'd22821, 16'd52601, 16'd25788, 16'd8611, 16'd29226, 16'd28510, 16'd52244, 16'd48536, 16'd62092, 16'd54476, 16'd23285, 16'd6060, 16'd22674, 16'd39374, 16'd61341, 16'd53755});
	test_expansion(128'h1fb6939799b5b6c7329b44a1681c37ad, {16'd38109, 16'd44897, 16'd49398, 16'd44662, 16'd38099, 16'd61973, 16'd28231, 16'd52807, 16'd24317, 16'd65216, 16'd45511, 16'd64536, 16'd1709, 16'd44874, 16'd28703, 16'd533, 16'd62602, 16'd6312, 16'd29071, 16'd55715, 16'd524, 16'd29590, 16'd61103, 16'd39747, 16'd5057, 16'd1208});
	test_expansion(128'h93b8017152d03954a5b0c1bd77030e19, {16'd46197, 16'd4394, 16'd51039, 16'd20957, 16'd63077, 16'd42356, 16'd5908, 16'd26166, 16'd36431, 16'd35066, 16'd4349, 16'd38814, 16'd6274, 16'd54610, 16'd440, 16'd63449, 16'd65245, 16'd64286, 16'd38599, 16'd29933, 16'd17944, 16'd51638, 16'd42010, 16'd21644, 16'd46927, 16'd44924});
	test_expansion(128'h38f9381e725252fd85dc95bfc524a1c6, {16'd53262, 16'd9978, 16'd45635, 16'd11208, 16'd43886, 16'd48446, 16'd60769, 16'd12860, 16'd6299, 16'd10295, 16'd35112, 16'd10822, 16'd30448, 16'd28963, 16'd2098, 16'd65081, 16'd16250, 16'd59636, 16'd26192, 16'd34692, 16'd51636, 16'd9857, 16'd63643, 16'd1985, 16'd30611, 16'd32834});
	test_expansion(128'hc3938b41527e5d8e842b8bcb67d42366, {16'd54266, 16'd17879, 16'd1275, 16'd53491, 16'd19298, 16'd14662, 16'd56620, 16'd15923, 16'd21702, 16'd73, 16'd59571, 16'd58768, 16'd20679, 16'd27980, 16'd1754, 16'd11975, 16'd14502, 16'd28947, 16'd38869, 16'd21555, 16'd47644, 16'd38619, 16'd24388, 16'd32881, 16'd5985, 16'd48002});
	test_expansion(128'hdb5abe2e1b1afe25c6b570d682bc7225, {16'd57816, 16'd50642, 16'd23527, 16'd3798, 16'd49091, 16'd16256, 16'd36548, 16'd38433, 16'd23400, 16'd47657, 16'd464, 16'd58966, 16'd65056, 16'd45352, 16'd36140, 16'd20014, 16'd34259, 16'd41911, 16'd7398, 16'd15474, 16'd31745, 16'd14372, 16'd64336, 16'd54487, 16'd48796, 16'd17265});
	test_expansion(128'h2da67a9dbe977271051018ed2f43fe85, {16'd23073, 16'd42858, 16'd7649, 16'd12032, 16'd56091, 16'd63052, 16'd49466, 16'd50370, 16'd52825, 16'd15496, 16'd44020, 16'd51103, 16'd12266, 16'd28479, 16'd59174, 16'd4278, 16'd4266, 16'd5639, 16'd5238, 16'd56104, 16'd15015, 16'd57053, 16'd47191, 16'd38115, 16'd26832, 16'd56883});
	test_expansion(128'h552f90d2dd93828589821b4ae0c45c17, {16'd27371, 16'd42533, 16'd36579, 16'd23706, 16'd2237, 16'd35250, 16'd21024, 16'd45563, 16'd27503, 16'd55635, 16'd4312, 16'd54295, 16'd42220, 16'd60926, 16'd60446, 16'd18216, 16'd52805, 16'd5686, 16'd21283, 16'd28582, 16'd21781, 16'd45785, 16'd4901, 16'd21558, 16'd12595, 16'd64012});
	test_expansion(128'hfafa1c8381a0fe50d906128c4060285c, {16'd58988, 16'd43178, 16'd59992, 16'd27015, 16'd38297, 16'd53086, 16'd29941, 16'd37462, 16'd20695, 16'd23205, 16'd35886, 16'd55966, 16'd54442, 16'd40735, 16'd57841, 16'd22650, 16'd33772, 16'd16781, 16'd58448, 16'd15767, 16'd53465, 16'd51115, 16'd64380, 16'd49068, 16'd32222, 16'd21132});
	test_expansion(128'heb9312750a47113b9e0653fd846df6af, {16'd45210, 16'd4857, 16'd41256, 16'd22007, 16'd18484, 16'd22322, 16'd26554, 16'd5382, 16'd32007, 16'd42162, 16'd31853, 16'd42055, 16'd63602, 16'd16386, 16'd38550, 16'd1771, 16'd14933, 16'd21249, 16'd10940, 16'd62243, 16'd64792, 16'd63240, 16'd36833, 16'd63650, 16'd40557, 16'd14630});
	test_expansion(128'hbcfae5cdab7e533ed693bad9c306a23a, {16'd13149, 16'd18601, 16'd35337, 16'd36774, 16'd44814, 16'd14965, 16'd52534, 16'd22117, 16'd1839, 16'd13299, 16'd14751, 16'd33596, 16'd39481, 16'd31398, 16'd32339, 16'd22502, 16'd25131, 16'd39471, 16'd33227, 16'd31930, 16'd56558, 16'd14166, 16'd65038, 16'd4448, 16'd64776, 16'd6650});
	test_expansion(128'h2a47298a8068b2d132f0f447d8294722, {16'd30945, 16'd63185, 16'd38783, 16'd6461, 16'd4085, 16'd30965, 16'd18860, 16'd9078, 16'd10908, 16'd3068, 16'd5997, 16'd46588, 16'd49406, 16'd9659, 16'd49663, 16'd861, 16'd30945, 16'd31860, 16'd64716, 16'd11328, 16'd54548, 16'd63476, 16'd62216, 16'd54486, 16'd23559, 16'd51850});
	test_expansion(128'h1560f311e4b0c43abec861146bb38215, {16'd33183, 16'd7513, 16'd52311, 16'd25226, 16'd61661, 16'd63758, 16'd42746, 16'd41085, 16'd2821, 16'd23921, 16'd45218, 16'd64730, 16'd16384, 16'd45958, 16'd20497, 16'd55087, 16'd60892, 16'd32689, 16'd28315, 16'd56132, 16'd29554, 16'd1753, 16'd52838, 16'd6116, 16'd50925, 16'd28419});
	test_expansion(128'hd557b269414960c3aeeeede1593eb6e3, {16'd6317, 16'd10660, 16'd26030, 16'd9637, 16'd29531, 16'd15524, 16'd37377, 16'd48518, 16'd18228, 16'd38718, 16'd44666, 16'd57335, 16'd51930, 16'd51207, 16'd39695, 16'd15948, 16'd53707, 16'd9488, 16'd4714, 16'd42932, 16'd45127, 16'd21925, 16'd46352, 16'd45512, 16'd52833, 16'd2387});
	test_expansion(128'hc7fe36e16781106b8af4087db1519bb0, {16'd62568, 16'd55124, 16'd18046, 16'd30521, 16'd63573, 16'd54575, 16'd63052, 16'd36875, 16'd280, 16'd59214, 16'd62747, 16'd8874, 16'd25602, 16'd28385, 16'd8112, 16'd7257, 16'd25179, 16'd30514, 16'd18706, 16'd19186, 16'd179, 16'd20204, 16'd35743, 16'd59707, 16'd250, 16'd51343});
	test_expansion(128'hc1c77863bf1de63b036be3fc5204dd40, {16'd3320, 16'd64050, 16'd46907, 16'd4346, 16'd8915, 16'd19876, 16'd59294, 16'd59033, 16'd45060, 16'd7229, 16'd47784, 16'd26855, 16'd39702, 16'd27462, 16'd4664, 16'd48263, 16'd6358, 16'd43963, 16'd4960, 16'd15994, 16'd45901, 16'd29051, 16'd32510, 16'd12364, 16'd36058, 16'd33000});
	test_expansion(128'hc85013350a88d1f893bf5f0a51b543fa, {16'd31627, 16'd56107, 16'd3566, 16'd57666, 16'd6143, 16'd15401, 16'd43857, 16'd34278, 16'd29290, 16'd6301, 16'd45152, 16'd58359, 16'd25558, 16'd29184, 16'd9661, 16'd25029, 16'd51403, 16'd12673, 16'd47257, 16'd15736, 16'd32351, 16'd8115, 16'd229, 16'd890, 16'd17730, 16'd20858});
	test_expansion(128'he2ae4899bc1161824017997296e2e8a8, {16'd6988, 16'd30353, 16'd58838, 16'd20171, 16'd52005, 16'd40319, 16'd21887, 16'd16575, 16'd55214, 16'd17962, 16'd30775, 16'd25097, 16'd39745, 16'd31606, 16'd37669, 16'd50640, 16'd35791, 16'd25684, 16'd45128, 16'd48767, 16'd5380, 16'd26559, 16'd2531, 16'd44857, 16'd62041, 16'd24815});
	test_expansion(128'h804a81b675f5c28f4968bf402aa9ce96, {16'd43295, 16'd24197, 16'd6734, 16'd39215, 16'd40592, 16'd29662, 16'd37399, 16'd15724, 16'd8571, 16'd49982, 16'd13081, 16'd23006, 16'd15866, 16'd30765, 16'd4052, 16'd49071, 16'd57301, 16'd2983, 16'd7733, 16'd55171, 16'd10402, 16'd52826, 16'd22926, 16'd61707, 16'd47250, 16'd35479});
	test_expansion(128'h5f41345d19f760a4885d32b6fa5fcde9, {16'd59462, 16'd3282, 16'd55938, 16'd44152, 16'd25464, 16'd18961, 16'd19033, 16'd5708, 16'd12581, 16'd57369, 16'd42817, 16'd44954, 16'd38088, 16'd20833, 16'd25655, 16'd2000, 16'd61688, 16'd2161, 16'd34725, 16'd35411, 16'd64258, 16'd35691, 16'd30001, 16'd36714, 16'd53902, 16'd42073});
	test_expansion(128'h15c31fba9aba7825fdee66fa809e016b, {16'd46369, 16'd49048, 16'd47446, 16'd40153, 16'd61266, 16'd10831, 16'd21834, 16'd20176, 16'd39100, 16'd13878, 16'd32121, 16'd40383, 16'd10558, 16'd64195, 16'd2890, 16'd65363, 16'd42103, 16'd10955, 16'd24615, 16'd61139, 16'd20039, 16'd45488, 16'd8221, 16'd43318, 16'd35999, 16'd2397});
	test_expansion(128'hbfe0657d490a11236bdb892768dd027b, {16'd33142, 16'd44001, 16'd63166, 16'd38493, 16'd64336, 16'd60841, 16'd53490, 16'd37215, 16'd16361, 16'd1889, 16'd57562, 16'd28368, 16'd46779, 16'd48455, 16'd25321, 16'd49292, 16'd19767, 16'd49552, 16'd23875, 16'd27995, 16'd24175, 16'd22749, 16'd18463, 16'd12785, 16'd43082, 16'd57586});
	test_expansion(128'h0b17c3b85065ad2867f1b466205d9923, {16'd23652, 16'd51476, 16'd51256, 16'd53927, 16'd18597, 16'd35760, 16'd11251, 16'd15788, 16'd12820, 16'd34857, 16'd33852, 16'd60483, 16'd47988, 16'd5404, 16'd16131, 16'd16710, 16'd42517, 16'd46427, 16'd5333, 16'd36965, 16'd10112, 16'd43206, 16'd36932, 16'd10263, 16'd10479, 16'd39715});
	test_expansion(128'hd3085050dbe4d5f3b66cc7493357b304, {16'd3474, 16'd48117, 16'd59401, 16'd48251, 16'd47953, 16'd49204, 16'd7729, 16'd42290, 16'd10221, 16'd43375, 16'd57279, 16'd13524, 16'd44278, 16'd35180, 16'd62186, 16'd44591, 16'd17652, 16'd39649, 16'd38809, 16'd59865, 16'd5756, 16'd18621, 16'd46936, 16'd37408, 16'd22291, 16'd30039});
	test_expansion(128'hb6129a1d35289a415dc37e2b8f34bca2, {16'd30154, 16'd12630, 16'd52989, 16'd25856, 16'd22310, 16'd7588, 16'd12266, 16'd43194, 16'd13722, 16'd36659, 16'd23784, 16'd10396, 16'd52335, 16'd23692, 16'd49061, 16'd21413, 16'd20940, 16'd30639, 16'd4142, 16'd47374, 16'd45349, 16'd9982, 16'd35055, 16'd33733, 16'd14743, 16'd13646});
	test_expansion(128'hb6c809ddbc0744b7c1a1e02128cbd671, {16'd48517, 16'd56926, 16'd39586, 16'd43328, 16'd885, 16'd49115, 16'd52989, 16'd13998, 16'd37500, 16'd14484, 16'd59888, 16'd15678, 16'd65436, 16'd17751, 16'd54587, 16'd30029, 16'd30114, 16'd32878, 16'd11411, 16'd61108, 16'd29478, 16'd31272, 16'd64340, 16'd48624, 16'd36556, 16'd55656});
	test_expansion(128'h934381d5f0e9e6a93ee6e0b7acbca980, {16'd64642, 16'd52881, 16'd38718, 16'd61903, 16'd60552, 16'd18422, 16'd2744, 16'd38108, 16'd47605, 16'd28344, 16'd8622, 16'd3546, 16'd56474, 16'd7928, 16'd59822, 16'd28776, 16'd30089, 16'd15070, 16'd32111, 16'd52660, 16'd53465, 16'd13032, 16'd623, 16'd22949, 16'd65070, 16'd34683});
	test_expansion(128'h4b5d332d709a1843c6b04fdcd94ca49d, {16'd6810, 16'd56217, 16'd17833, 16'd6362, 16'd21148, 16'd57736, 16'd9881, 16'd51603, 16'd29273, 16'd50894, 16'd20974, 16'd5843, 16'd10354, 16'd35860, 16'd37027, 16'd24871, 16'd46054, 16'd9481, 16'd38043, 16'd17096, 16'd35237, 16'd33320, 16'd59645, 16'd26013, 16'd3125, 16'd48444});
	test_expansion(128'h729a985d78f152aa2ebff0a9be30a2ab, {16'd1516, 16'd36405, 16'd12416, 16'd16486, 16'd18117, 16'd32551, 16'd7837, 16'd46878, 16'd49254, 16'd35411, 16'd20810, 16'd62844, 16'd10448, 16'd21793, 16'd54090, 16'd7262, 16'd55382, 16'd24019, 16'd9593, 16'd19744, 16'd51506, 16'd3514, 16'd64344, 16'd22415, 16'd41665, 16'd12506});
	test_expansion(128'h3ecf0866202fb44c0e8d838d8be062cb, {16'd5810, 16'd1699, 16'd15046, 16'd416, 16'd61237, 16'd64720, 16'd25761, 16'd30617, 16'd11649, 16'd46594, 16'd44199, 16'd23785, 16'd64985, 16'd28925, 16'd62148, 16'd54389, 16'd43546, 16'd59008, 16'd33665, 16'd45547, 16'd9704, 16'd1112, 16'd31016, 16'd36371, 16'd53863, 16'd60734});
	test_expansion(128'h40b612924fc9143ebd8d82e1ee5eba85, {16'd17816, 16'd62683, 16'd56274, 16'd59358, 16'd62336, 16'd33967, 16'd65168, 16'd5768, 16'd981, 16'd30347, 16'd36582, 16'd58295, 16'd60954, 16'd22765, 16'd47512, 16'd6047, 16'd45252, 16'd11203, 16'd50941, 16'd12989, 16'd5397, 16'd25482, 16'd63142, 16'd52072, 16'd42636, 16'd4442});
	test_expansion(128'hdecf209930e4b2585220807025552e79, {16'd27823, 16'd26624, 16'd38657, 16'd52685, 16'd65501, 16'd10719, 16'd38087, 16'd45571, 16'd15411, 16'd11223, 16'd3055, 16'd25703, 16'd32991, 16'd40962, 16'd321, 16'd48531, 16'd55102, 16'd48099, 16'd3637, 16'd21696, 16'd34398, 16'd65225, 16'd6683, 16'd6907, 16'd13488, 16'd39742});
	test_expansion(128'h3e4d2f34355f6136cabba95e2735a608, {16'd50464, 16'd11475, 16'd61034, 16'd164, 16'd23681, 16'd36207, 16'd24568, 16'd34214, 16'd33146, 16'd65495, 16'd24198, 16'd16229, 16'd40758, 16'd8813, 16'd62633, 16'd56601, 16'd34783, 16'd60358, 16'd36468, 16'd3769, 16'd787, 16'd17161, 16'd60520, 16'd62684, 16'd10495, 16'd17260});
	test_expansion(128'hc4f2b30fb2fd25d9e03341eaca3c7c50, {16'd53494, 16'd7829, 16'd24154, 16'd42377, 16'd37706, 16'd12881, 16'd28259, 16'd34372, 16'd55721, 16'd18054, 16'd8024, 16'd20370, 16'd24270, 16'd18321, 16'd25831, 16'd57391, 16'd7791, 16'd9959, 16'd15891, 16'd40905, 16'd19076, 16'd42730, 16'd33781, 16'd14716, 16'd54806, 16'd11140});
	test_expansion(128'h62258d1b866f190d9d65c20d0c154f57, {16'd43022, 16'd3743, 16'd21329, 16'd23879, 16'd55019, 16'd18884, 16'd34902, 16'd52324, 16'd5403, 16'd38614, 16'd24035, 16'd58890, 16'd62820, 16'd580, 16'd303, 16'd34989, 16'd51945, 16'd54723, 16'd51894, 16'd63133, 16'd40823, 16'd15518, 16'd7208, 16'd20290, 16'd35304, 16'd24733});
	test_expansion(128'hd48df5748c9675d16a3221b303349070, {16'd25845, 16'd50577, 16'd41477, 16'd15038, 16'd61577, 16'd44631, 16'd22039, 16'd48878, 16'd52760, 16'd40008, 16'd56836, 16'd11140, 16'd18242, 16'd10119, 16'd42954, 16'd9963, 16'd52715, 16'd6983, 16'd1984, 16'd57225, 16'd3939, 16'd53007, 16'd28173, 16'd1015, 16'd27850, 16'd45951});
	test_expansion(128'hc2a2e09f0610f7fbda4da089da89f9f6, {16'd7837, 16'd64715, 16'd13907, 16'd63513, 16'd14306, 16'd16261, 16'd2823, 16'd47375, 16'd58679, 16'd60349, 16'd3648, 16'd61041, 16'd14197, 16'd3315, 16'd11576, 16'd61074, 16'd4952, 16'd49205, 16'd53686, 16'd1420, 16'd23484, 16'd22719, 16'd58178, 16'd29683, 16'd39178, 16'd16091});
	test_expansion(128'h049e401c833154fc56100b167fb0d088, {16'd2933, 16'd21243, 16'd36425, 16'd57476, 16'd59208, 16'd11954, 16'd39443, 16'd6420, 16'd32396, 16'd35587, 16'd51056, 16'd14390, 16'd58251, 16'd12710, 16'd12266, 16'd51118, 16'd14862, 16'd64284, 16'd54050, 16'd51645, 16'd21646, 16'd59067, 16'd23397, 16'd58838, 16'd42617, 16'd20618});
	test_expansion(128'hade7a2b7b47bcb3b3f1d0fdb4080c0df, {16'd22963, 16'd44442, 16'd39228, 16'd39677, 16'd54841, 16'd51582, 16'd59400, 16'd54490, 16'd16531, 16'd14935, 16'd54224, 16'd37005, 16'd30022, 16'd61176, 16'd29168, 16'd30271, 16'd49426, 16'd13691, 16'd64193, 16'd56822, 16'd39951, 16'd10283, 16'd7918, 16'd14731, 16'd24130, 16'd20180});
	test_expansion(128'he334663376698b00bab4f343cc107be9, {16'd33156, 16'd41028, 16'd61554, 16'd47045, 16'd39161, 16'd30566, 16'd56306, 16'd50133, 16'd63412, 16'd52729, 16'd15770, 16'd43035, 16'd60070, 16'd10783, 16'd27882, 16'd12514, 16'd58627, 16'd7272, 16'd13934, 16'd9914, 16'd61393, 16'd12376, 16'd28487, 16'd2685, 16'd56471, 16'd47996});
	test_expansion(128'had6fb1c06a34e0ae77126c25ea571e34, {16'd30375, 16'd6419, 16'd39880, 16'd43228, 16'd32636, 16'd282, 16'd22096, 16'd59315, 16'd5057, 16'd64434, 16'd35856, 16'd37918, 16'd9495, 16'd47264, 16'd63289, 16'd34396, 16'd21933, 16'd46540, 16'd58192, 16'd41539, 16'd47388, 16'd50077, 16'd6254, 16'd39295, 16'd59222, 16'd6852});
	test_expansion(128'h8ddcf5341b77a2da84d16f14c50bf86e, {16'd13792, 16'd47435, 16'd16571, 16'd61353, 16'd62248, 16'd11433, 16'd31168, 16'd59253, 16'd17653, 16'd49197, 16'd26984, 16'd27924, 16'd63594, 16'd17296, 16'd49106, 16'd58149, 16'd50652, 16'd35794, 16'd21625, 16'd61809, 16'd24873, 16'd102, 16'd28395, 16'd17497, 16'd51371, 16'd54293});
	test_expansion(128'h1f94b6139c709c96e376b705e3180747, {16'd47294, 16'd48529, 16'd14005, 16'd24660, 16'd45033, 16'd30278, 16'd21565, 16'd45164, 16'd7005, 16'd22118, 16'd5550, 16'd55277, 16'd39546, 16'd15656, 16'd48450, 16'd20330, 16'd228, 16'd34154, 16'd12240, 16'd62668, 16'd40613, 16'd52093, 16'd22219, 16'd4996, 16'd38656, 16'd7263});
	test_expansion(128'h690b0948ddc0be86bf2858df0cc04c9d, {16'd32472, 16'd12513, 16'd35320, 16'd4429, 16'd31389, 16'd27564, 16'd17122, 16'd6019, 16'd20331, 16'd35184, 16'd43507, 16'd42566, 16'd31055, 16'd29646, 16'd32667, 16'd1923, 16'd18382, 16'd51152, 16'd36110, 16'd9215, 16'd43272, 16'd19093, 16'd19253, 16'd43667, 16'd42085, 16'd4761});
	test_expansion(128'ha37d72607b84205c9af7aceaad9c912e, {16'd33542, 16'd28039, 16'd3852, 16'd23178, 16'd64344, 16'd58823, 16'd56458, 16'd8762, 16'd321, 16'd9782, 16'd46407, 16'd18946, 16'd12801, 16'd47865, 16'd63008, 16'd55106, 16'd47435, 16'd28502, 16'd33216, 16'd32, 16'd19936, 16'd44096, 16'd31111, 16'd37174, 16'd12867, 16'd13239});
	test_expansion(128'h34233242d4794cadb19376cf65e9bc6a, {16'd52325, 16'd7782, 16'd62188, 16'd31710, 16'd65267, 16'd31149, 16'd18281, 16'd42252, 16'd35854, 16'd36701, 16'd17707, 16'd36697, 16'd59257, 16'd17313, 16'd24218, 16'd50562, 16'd33824, 16'd31592, 16'd26574, 16'd64868, 16'd17321, 16'd29909, 16'd6330, 16'd27072, 16'd29073, 16'd40202});
	test_expansion(128'hfd3f8b82ecdd9040c6c3437ce4d100f7, {16'd27152, 16'd22473, 16'd25838, 16'd272, 16'd10209, 16'd56988, 16'd19551, 16'd9021, 16'd7272, 16'd48178, 16'd64945, 16'd65484, 16'd13740, 16'd2077, 16'd40807, 16'd26380, 16'd47483, 16'd6236, 16'd48600, 16'd27245, 16'd2606, 16'd60992, 16'd44975, 16'd59745, 16'd52079, 16'd34195});
	test_expansion(128'hbb18e280f6e9ed141e813501278394ee, {16'd10450, 16'd36092, 16'd25319, 16'd19089, 16'd26904, 16'd38516, 16'd7511, 16'd5151, 16'd38011, 16'd38135, 16'd17284, 16'd33514, 16'd40381, 16'd11245, 16'd54880, 16'd52001, 16'd45375, 16'd50051, 16'd23597, 16'd9634, 16'd59099, 16'd45754, 16'd35721, 16'd48477, 16'd22309, 16'd25478});
	test_expansion(128'h6018af9f20f7bf1857b48d703954305d, {16'd37942, 16'd15049, 16'd2997, 16'd31119, 16'd28714, 16'd39656, 16'd32914, 16'd24484, 16'd39053, 16'd27335, 16'd31583, 16'd60273, 16'd38904, 16'd7890, 16'd56348, 16'd18378, 16'd58568, 16'd20349, 16'd63190, 16'd8617, 16'd11175, 16'd35608, 16'd1978, 16'd53918, 16'd47222, 16'd51450});
	test_expansion(128'h8e47ebbe07aea440e57b5090a26e71e0, {16'd5097, 16'd42974, 16'd20532, 16'd59256, 16'd12129, 16'd61142, 16'd46068, 16'd44458, 16'd47516, 16'd67, 16'd5643, 16'd18833, 16'd15023, 16'd25844, 16'd33361, 16'd2030, 16'd61881, 16'd14966, 16'd28137, 16'd39687, 16'd56068, 16'd62048, 16'd31411, 16'd20037, 16'd25840, 16'd13966});
	test_expansion(128'ha92dcadddf8e8c14d44d2926fe7d0233, {16'd7734, 16'd5072, 16'd22054, 16'd25682, 16'd52295, 16'd55538, 16'd61737, 16'd35385, 16'd49052, 16'd10525, 16'd29312, 16'd19597, 16'd53690, 16'd44124, 16'd4166, 16'd60435, 16'd41787, 16'd24910, 16'd16864, 16'd15127, 16'd39307, 16'd15714, 16'd8345, 16'd35196, 16'd3491, 16'd9696});
	test_expansion(128'h0886b019c7473a520fb163fff204e9b3, {16'd43029, 16'd51519, 16'd45228, 16'd29038, 16'd8568, 16'd12573, 16'd2738, 16'd3008, 16'd11359, 16'd39319, 16'd59689, 16'd61148, 16'd38652, 16'd22120, 16'd30729, 16'd27865, 16'd17992, 16'd10593, 16'd3202, 16'd36671, 16'd2496, 16'd44985, 16'd15133, 16'd43976, 16'd10203, 16'd42302});
	test_expansion(128'h80a679edf9f3cf12333053ce01bd623f, {16'd48499, 16'd43891, 16'd915, 16'd59492, 16'd32183, 16'd33821, 16'd44355, 16'd44179, 16'd56564, 16'd63941, 16'd51823, 16'd30657, 16'd15152, 16'd54101, 16'd53471, 16'd37618, 16'd436, 16'd44689, 16'd30578, 16'd62837, 16'd32921, 16'd49784, 16'd62179, 16'd62864, 16'd65274, 16'd24787});
	test_expansion(128'hd105bff17407d77b1bb910ab8b2b2542, {16'd10317, 16'd6207, 16'd6528, 16'd14799, 16'd10805, 16'd62836, 16'd13098, 16'd41880, 16'd37432, 16'd33156, 16'd5146, 16'd37236, 16'd61381, 16'd10660, 16'd56534, 16'd40984, 16'd24129, 16'd32528, 16'd41256, 16'd52653, 16'd2719, 16'd10872, 16'd44721, 16'd6863, 16'd45619, 16'd38321});
	test_expansion(128'h652ac0a376767876d376c2473f11b4f8, {16'd61471, 16'd24977, 16'd24064, 16'd10433, 16'd31133, 16'd62651, 16'd23749, 16'd37129, 16'd31312, 16'd31480, 16'd30633, 16'd64276, 16'd33243, 16'd37887, 16'd62377, 16'd10931, 16'd59060, 16'd50387, 16'd33443, 16'd12154, 16'd58977, 16'd33884, 16'd64577, 16'd10559, 16'd56273, 16'd61780});
	test_expansion(128'haaf1764f38a38b02b44100b0dd730517, {16'd44602, 16'd41335, 16'd19037, 16'd19668, 16'd16595, 16'd19329, 16'd35420, 16'd37097, 16'd21764, 16'd39366, 16'd41796, 16'd13382, 16'd45290, 16'd10827, 16'd6387, 16'd12845, 16'd22042, 16'd49161, 16'd46904, 16'd17858, 16'd42399, 16'd13997, 16'd25596, 16'd40160, 16'd26813, 16'd42517});
	test_expansion(128'ha7a0d6ddbd8567fb9b71fd578e020a27, {16'd16148, 16'd46549, 16'd25527, 16'd11104, 16'd2325, 16'd28438, 16'd62892, 16'd17846, 16'd24805, 16'd59742, 16'd9140, 16'd28577, 16'd31116, 16'd30482, 16'd57056, 16'd41472, 16'd4344, 16'd16451, 16'd20356, 16'd490, 16'd8082, 16'd48577, 16'd34326, 16'd26813, 16'd13565, 16'd4534});
	test_expansion(128'he828645e907d2000ae080af1fd2efd78, {16'd5321, 16'd14304, 16'd39501, 16'd4387, 16'd7317, 16'd49909, 16'd47995, 16'd10445, 16'd60766, 16'd42776, 16'd60981, 16'd5248, 16'd10706, 16'd19582, 16'd33947, 16'd28033, 16'd6297, 16'd34631, 16'd61154, 16'd3256, 16'd34142, 16'd18620, 16'd4420, 16'd6283, 16'd13460, 16'd13468});
	test_expansion(128'hdbc4a0676adb0c6e6eecb60194a03c70, {16'd53085, 16'd1493, 16'd63993, 16'd48176, 16'd45430, 16'd57858, 16'd17835, 16'd44872, 16'd23407, 16'd7323, 16'd2103, 16'd20469, 16'd8935, 16'd6138, 16'd9433, 16'd21698, 16'd15377, 16'd28347, 16'd585, 16'd61498, 16'd23824, 16'd54797, 16'd37808, 16'd48273, 16'd25582, 16'd64164});
	test_expansion(128'h8341b14e85ce6fa418663c8f584b7014, {16'd38380, 16'd37087, 16'd11533, 16'd11202, 16'd52500, 16'd25323, 16'd45202, 16'd13392, 16'd59526, 16'd9843, 16'd3837, 16'd33457, 16'd54045, 16'd15823, 16'd24749, 16'd45687, 16'd5235, 16'd4890, 16'd37758, 16'd35763, 16'd26248, 16'd36237, 16'd52141, 16'd56246, 16'd10013, 16'd19675});
	test_expansion(128'h01fad6fbcde7809a1e3d69201837cd66, {16'd8369, 16'd32454, 16'd17844, 16'd27864, 16'd16877, 16'd21010, 16'd47087, 16'd13520, 16'd52235, 16'd27544, 16'd53196, 16'd42329, 16'd24357, 16'd8403, 16'd33458, 16'd32274, 16'd32276, 16'd17001, 16'd40546, 16'd56914, 16'd10660, 16'd52907, 16'd13071, 16'd18631, 16'd32254, 16'd46008});
	test_expansion(128'ha3b9b700f9be7fdefcaee14655e258da, {16'd56481, 16'd37864, 16'd54795, 16'd26387, 16'd61904, 16'd52986, 16'd5753, 16'd166, 16'd3443, 16'd9594, 16'd63450, 16'd26851, 16'd30971, 16'd34445, 16'd48907, 16'd8268, 16'd529, 16'd32545, 16'd60995, 16'd30379, 16'd17443, 16'd58015, 16'd23786, 16'd54712, 16'd48402, 16'd2213});
	test_expansion(128'hd2aaf07d38e63fea7ee0949bdf5d5f70, {16'd8975, 16'd21211, 16'd3032, 16'd27558, 16'd31222, 16'd14642, 16'd3867, 16'd5828, 16'd35719, 16'd5948, 16'd14075, 16'd38456, 16'd45685, 16'd11222, 16'd37673, 16'd13443, 16'd54691, 16'd11610, 16'd49818, 16'd8035, 16'd14866, 16'd4362, 16'd29374, 16'd16970, 16'd27726, 16'd32741});
	test_expansion(128'he06d65c406bf299fa1a1599234e07dba, {16'd35313, 16'd30486, 16'd34593, 16'd47285, 16'd19571, 16'd63871, 16'd5121, 16'd53187, 16'd62474, 16'd3519, 16'd31734, 16'd55493, 16'd56527, 16'd28254, 16'd59054, 16'd13439, 16'd34136, 16'd58182, 16'd24710, 16'd47271, 16'd30102, 16'd28705, 16'd1186, 16'd16548, 16'd15001, 16'd26529});
	test_expansion(128'h2c3888cd511415894f11498ac9530b8d, {16'd62055, 16'd47736, 16'd39557, 16'd51604, 16'd3389, 16'd8395, 16'd59787, 16'd9207, 16'd29768, 16'd24543, 16'd29308, 16'd20545, 16'd22201, 16'd50122, 16'd12521, 16'd15340, 16'd21283, 16'd12462, 16'd58525, 16'd4180, 16'd1238, 16'd26472, 16'd2375, 16'd9400, 16'd15894, 16'd45905});
	test_expansion(128'hf3a820698c546dd4e0e155c24eea8e41, {16'd63408, 16'd42145, 16'd34666, 16'd62116, 16'd47383, 16'd48226, 16'd34969, 16'd15528, 16'd33047, 16'd14889, 16'd24263, 16'd23682, 16'd29325, 16'd48187, 16'd4757, 16'd20627, 16'd65074, 16'd43633, 16'd65174, 16'd52578, 16'd36765, 16'd14771, 16'd21103, 16'd9457, 16'd39655, 16'd13198});
	test_expansion(128'hcbe4573c26832902d2ea7b34e739220c, {16'd51855, 16'd40133, 16'd52359, 16'd17241, 16'd5109, 16'd34766, 16'd22757, 16'd44155, 16'd19893, 16'd11707, 16'd19101, 16'd13741, 16'd57904, 16'd12579, 16'd36453, 16'd57320, 16'd37282, 16'd25336, 16'd48194, 16'd57886, 16'd15760, 16'd10022, 16'd13798, 16'd18517, 16'd58234, 16'd13236});
	test_expansion(128'h33e01e475a468077e05caba3c30f6150, {16'd26226, 16'd34876, 16'd18442, 16'd55763, 16'd30016, 16'd59888, 16'd17758, 16'd35670, 16'd47290, 16'd14720, 16'd54910, 16'd51849, 16'd41748, 16'd38260, 16'd28447, 16'd44200, 16'd8397, 16'd15937, 16'd13263, 16'd49603, 16'd43507, 16'd55102, 16'd11673, 16'd33846, 16'd21769, 16'd22743});
	test_expansion(128'h00d1e0c7845bda3dd73ae7b2ba9d2ad6, {16'd3971, 16'd24782, 16'd33496, 16'd52740, 16'd62834, 16'd25571, 16'd50752, 16'd33031, 16'd29977, 16'd19679, 16'd13150, 16'd59755, 16'd4934, 16'd42818, 16'd34954, 16'd9809, 16'd43737, 16'd6085, 16'd688, 16'd5915, 16'd17694, 16'd62896, 16'd14667, 16'd51819, 16'd33804, 16'd56421});
	test_expansion(128'haca9ade895a0126f73e77e08cce5a5ee, {16'd14977, 16'd701, 16'd6064, 16'd61825, 16'd46675, 16'd59361, 16'd62442, 16'd12220, 16'd19528, 16'd49180, 16'd47202, 16'd13153, 16'd21827, 16'd64896, 16'd56744, 16'd49628, 16'd8995, 16'd434, 16'd23579, 16'd20, 16'd37143, 16'd28102, 16'd4847, 16'd28848, 16'd7050, 16'd35361});
	test_expansion(128'h8859c62a8bbcdb7df832f6b8a84893b8, {16'd12100, 16'd11903, 16'd56154, 16'd47407, 16'd12827, 16'd46139, 16'd42956, 16'd7167, 16'd49178, 16'd62323, 16'd37957, 16'd57265, 16'd13031, 16'd26265, 16'd29645, 16'd58301, 16'd14046, 16'd4044, 16'd32880, 16'd19153, 16'd47080, 16'd58602, 16'd17488, 16'd54748, 16'd56697, 16'd55060});
	test_expansion(128'hee4e9b888d87a1e057df0dd900e6cf0f, {16'd50795, 16'd59736, 16'd36855, 16'd91, 16'd7459, 16'd35500, 16'd57487, 16'd46834, 16'd52959, 16'd32875, 16'd45944, 16'd29303, 16'd8221, 16'd23937, 16'd37663, 16'd39985, 16'd59275, 16'd33228, 16'd64384, 16'd56764, 16'd53070, 16'd42626, 16'd28865, 16'd14211, 16'd45384, 16'd39497});
	test_expansion(128'h7f4e992d8bd9bf13f6ed80459fc650d1, {16'd47754, 16'd26870, 16'd28056, 16'd17403, 16'd45842, 16'd42984, 16'd5311, 16'd33462, 16'd15049, 16'd53194, 16'd45465, 16'd28182, 16'd53533, 16'd53657, 16'd15052, 16'd22827, 16'd62342, 16'd23447, 16'd12360, 16'd21574, 16'd52669, 16'd16845, 16'd16057, 16'd35044, 16'd28365, 16'd12352});
	test_expansion(128'h0bd723ec76e3e4f5aef7fcd224a2a797, {16'd18927, 16'd4060, 16'd23953, 16'd23232, 16'd3512, 16'd32376, 16'd23640, 16'd14328, 16'd15643, 16'd23371, 16'd63878, 16'd51588, 16'd8090, 16'd34149, 16'd41327, 16'd58038, 16'd30046, 16'd58975, 16'd62809, 16'd35718, 16'd23783, 16'd52822, 16'd14471, 16'd61286, 16'd33788, 16'd64815});
	test_expansion(128'h96484d6be34fdcd7b1b37b04353b8009, {16'd39972, 16'd33885, 16'd18152, 16'd44151, 16'd59065, 16'd47613, 16'd53683, 16'd34333, 16'd61788, 16'd7251, 16'd50702, 16'd62107, 16'd6600, 16'd29293, 16'd36376, 16'd16734, 16'd1152, 16'd35360, 16'd42029, 16'd17664, 16'd20932, 16'd15475, 16'd25610, 16'd22977, 16'd53428, 16'd17830});
	test_expansion(128'hd6399ea45c0c9ad25eb7dfad23d1acec, {16'd47050, 16'd24258, 16'd41283, 16'd38944, 16'd61512, 16'd3343, 16'd56025, 16'd50671, 16'd57787, 16'd34247, 16'd48008, 16'd18340, 16'd64611, 16'd19988, 16'd8978, 16'd65019, 16'd39564, 16'd45230, 16'd32703, 16'd46807, 16'd10329, 16'd6453, 16'd31834, 16'd23908, 16'd59101, 16'd53509});
	test_expansion(128'h469f8fd55cd010a1d3b284b132193bd2, {16'd59777, 16'd35473, 16'd23137, 16'd5934, 16'd29620, 16'd36674, 16'd31109, 16'd27995, 16'd53679, 16'd53371, 16'd555, 16'd48859, 16'd13020, 16'd5523, 16'd62729, 16'd11623, 16'd6205, 16'd7719, 16'd10167, 16'd42308, 16'd45758, 16'd52762, 16'd22978, 16'd57346, 16'd39809, 16'd21474});
	test_expansion(128'h180d1af24ca709f5a2e376a1a314881b, {16'd51389, 16'd184, 16'd17257, 16'd50542, 16'd700, 16'd17999, 16'd27527, 16'd47952, 16'd39254, 16'd10435, 16'd59312, 16'd49508, 16'd42355, 16'd8623, 16'd38936, 16'd4260, 16'd45386, 16'd25601, 16'd22066, 16'd40725, 16'd63048, 16'd25370, 16'd45151, 16'd10515, 16'd2326, 16'd55742});
	test_expansion(128'h1b15dba7365567af8fc008c2f6f6ced3, {16'd26948, 16'd39667, 16'd18161, 16'd7746, 16'd41842, 16'd26943, 16'd24809, 16'd5825, 16'd317, 16'd40867, 16'd63441, 16'd25324, 16'd43065, 16'd59900, 16'd49291, 16'd45626, 16'd61336, 16'd36780, 16'd11058, 16'd36421, 16'd45379, 16'd60494, 16'd9979, 16'd39179, 16'd39084, 16'd150});
	test_expansion(128'hfcb81ca867fd481aa02f36e15af0ddc3, {16'd27858, 16'd51432, 16'd58310, 16'd13802, 16'd58688, 16'd21845, 16'd53453, 16'd18698, 16'd45653, 16'd1398, 16'd58856, 16'd34547, 16'd8585, 16'd26006, 16'd55841, 16'd6894, 16'd13249, 16'd19877, 16'd13189, 16'd2980, 16'd39150, 16'd28806, 16'd40443, 16'd11982, 16'd31206, 16'd54241});
	test_expansion(128'hc092dbf31f6af8e4d16ac167831155a3, {16'd7199, 16'd5531, 16'd38247, 16'd12075, 16'd25634, 16'd54625, 16'd34630, 16'd43761, 16'd8765, 16'd5151, 16'd52382, 16'd48590, 16'd43148, 16'd8581, 16'd18793, 16'd53195, 16'd20, 16'd36055, 16'd19206, 16'd36221, 16'd20244, 16'd64075, 16'd16009, 16'd43604, 16'd48154, 16'd11902});
	test_expansion(128'h398aed7f15f9ead6fcb4369369b6c97b, {16'd30889, 16'd27645, 16'd286, 16'd11263, 16'd6381, 16'd29239, 16'd56535, 16'd27446, 16'd57256, 16'd42082, 16'd20003, 16'd37589, 16'd34726, 16'd32120, 16'd21415, 16'd36354, 16'd34579, 16'd35189, 16'd10019, 16'd3607, 16'd51498, 16'd35878, 16'd47884, 16'd13001, 16'd2196, 16'd57843});
	test_expansion(128'h87f5eaba22f5e30c2a6f6a5c076f04c7, {16'd49058, 16'd5454, 16'd59428, 16'd17525, 16'd24522, 16'd9943, 16'd42312, 16'd31551, 16'd63909, 16'd130, 16'd48977, 16'd35013, 16'd3945, 16'd46985, 16'd46405, 16'd64635, 16'd21018, 16'd22238, 16'd40123, 16'd43292, 16'd57071, 16'd53870, 16'd58161, 16'd46883, 16'd30910, 16'd40596});
	test_expansion(128'hca0eac702e21ff4278545d0e96235f39, {16'd43289, 16'd19041, 16'd61923, 16'd25627, 16'd27715, 16'd11348, 16'd16830, 16'd57038, 16'd23637, 16'd2046, 16'd21342, 16'd21281, 16'd32855, 16'd62040, 16'd49131, 16'd12257, 16'd57582, 16'd35074, 16'd58489, 16'd55800, 16'd59199, 16'd41160, 16'd47247, 16'd21441, 16'd15635, 16'd9315});
	test_expansion(128'hb4ddc4ba5f1022b3cad9ebf87946360a, {16'd28904, 16'd15006, 16'd9429, 16'd50201, 16'd58070, 16'd52511, 16'd18627, 16'd51983, 16'd21993, 16'd33422, 16'd15615, 16'd34465, 16'd12098, 16'd33548, 16'd20191, 16'd24806, 16'd7731, 16'd50022, 16'd48908, 16'd45502, 16'd57803, 16'd17183, 16'd36102, 16'd48998, 16'd64542, 16'd51687});
	test_expansion(128'h955a9a6bd0a5e0dfc53f39854271ce67, {16'd6454, 16'd3390, 16'd48665, 16'd64916, 16'd40663, 16'd54092, 16'd32474, 16'd55110, 16'd20014, 16'd48466, 16'd2079, 16'd22767, 16'd34039, 16'd5141, 16'd22594, 16'd7020, 16'd51564, 16'd37654, 16'd33963, 16'd32922, 16'd27154, 16'd2657, 16'd43568, 16'd14727, 16'd21591, 16'd4401});
	test_expansion(128'h2c8a3692a249d9891649b0b598a3b716, {16'd7776, 16'd10788, 16'd40494, 16'd61955, 16'd3961, 16'd58191, 16'd53109, 16'd26932, 16'd14982, 16'd44364, 16'd30079, 16'd46550, 16'd37880, 16'd48853, 16'd55462, 16'd1873, 16'd44015, 16'd20335, 16'd22724, 16'd8417, 16'd30444, 16'd9704, 16'd21589, 16'd6437, 16'd64736, 16'd50925});
	test_expansion(128'h81431b082bdccf0f0a7b011bb6581b29, {16'd4163, 16'd25616, 16'd4475, 16'd63573, 16'd65368, 16'd17211, 16'd18752, 16'd58354, 16'd42657, 16'd48639, 16'd59973, 16'd37743, 16'd37128, 16'd22379, 16'd43248, 16'd33288, 16'd26006, 16'd13384, 16'd63507, 16'd17906, 16'd19187, 16'd25585, 16'd35164, 16'd25698, 16'd47641, 16'd22902});
	test_expansion(128'haca300584438d9554cf61e4c471db97a, {16'd44951, 16'd52480, 16'd56956, 16'd15512, 16'd29050, 16'd10222, 16'd31215, 16'd25868, 16'd12224, 16'd43483, 16'd14731, 16'd51733, 16'd35169, 16'd13082, 16'd57885, 16'd22169, 16'd26387, 16'd50692, 16'd62747, 16'd20553, 16'd46405, 16'd52657, 16'd29794, 16'd41611, 16'd54189, 16'd17002});
	test_expansion(128'hfc6f7c1163dea22236d7b120820908c2, {16'd65376, 16'd49240, 16'd42567, 16'd30453, 16'd57240, 16'd21181, 16'd55396, 16'd26235, 16'd59828, 16'd14439, 16'd693, 16'd62591, 16'd59542, 16'd35337, 16'd41957, 16'd53542, 16'd62493, 16'd15715, 16'd18108, 16'd58047, 16'd15618, 16'd42221, 16'd62977, 16'd4028, 16'd5514, 16'd41474});
	test_expansion(128'h34b2684e0b112bbfebdbdb8b66c7a321, {16'd21651, 16'd22473, 16'd12553, 16'd62030, 16'd23874, 16'd28489, 16'd33698, 16'd23841, 16'd34258, 16'd2602, 16'd64327, 16'd9613, 16'd44037, 16'd32695, 16'd4620, 16'd7294, 16'd44086, 16'd19685, 16'd36258, 16'd59478, 16'd44123, 16'd33424, 16'd9197, 16'd9599, 16'd28596, 16'd3018});
	test_expansion(128'h84752fcbcd541391a7b324d89d9742f9, {16'd4477, 16'd2307, 16'd3538, 16'd2427, 16'd38302, 16'd55970, 16'd65002, 16'd53044, 16'd42987, 16'd52888, 16'd30861, 16'd7853, 16'd22906, 16'd58565, 16'd40054, 16'd37545, 16'd54515, 16'd24573, 16'd25401, 16'd27959, 16'd29578, 16'd49675, 16'd2620, 16'd4829, 16'd6165, 16'd32399});
	test_expansion(128'h0e8035209e55df97db28bac9406fd3ba, {16'd2829, 16'd40098, 16'd16115, 16'd1965, 16'd48688, 16'd1865, 16'd54635, 16'd64896, 16'd32560, 16'd7009, 16'd35501, 16'd65321, 16'd48699, 16'd6459, 16'd9406, 16'd51097, 16'd6932, 16'd19753, 16'd19565, 16'd37731, 16'd11241, 16'd37110, 16'd12899, 16'd15379, 16'd16420, 16'd8690});
	test_expansion(128'h77d6c678ab7beb2cb64001cfe4b93f64, {16'd4280, 16'd19790, 16'd55596, 16'd51643, 16'd13851, 16'd3791, 16'd44353, 16'd36391, 16'd13703, 16'd56413, 16'd34133, 16'd41645, 16'd59468, 16'd31256, 16'd15441, 16'd64877, 16'd50609, 16'd56813, 16'd18325, 16'd820, 16'd63567, 16'd35452, 16'd54687, 16'd36663, 16'd8274, 16'd24343});
	test_expansion(128'h10028c338ba0fb3c0c3462b920ab453d, {16'd13524, 16'd10796, 16'd64810, 16'd40838, 16'd26212, 16'd27506, 16'd48387, 16'd30239, 16'd10987, 16'd64509, 16'd24310, 16'd33565, 16'd53922, 16'd62058, 16'd54724, 16'd38392, 16'd16120, 16'd56694, 16'd53256, 16'd43529, 16'd31991, 16'd27119, 16'd55691, 16'd65055, 16'd52962, 16'd64733});
	test_expansion(128'he1e5e45e46a83215cb4015189601ab4d, {16'd2631, 16'd7575, 16'd48572, 16'd19625, 16'd53667, 16'd65488, 16'd45995, 16'd39878, 16'd21306, 16'd9165, 16'd58420, 16'd6738, 16'd50144, 16'd512, 16'd54748, 16'd18380, 16'd44386, 16'd46689, 16'd12988, 16'd17996, 16'd58486, 16'd25005, 16'd41499, 16'd52228, 16'd46341, 16'd213});
	test_expansion(128'h6fa6047f75dbcb56b4e37e92d9adbca1, {16'd25337, 16'd34709, 16'd29647, 16'd61782, 16'd55804, 16'd43713, 16'd12438, 16'd53204, 16'd60833, 16'd8365, 16'd2050, 16'd48337, 16'd41054, 16'd15204, 16'd55833, 16'd27132, 16'd4268, 16'd36147, 16'd37422, 16'd27336, 16'd10323, 16'd2704, 16'd38674, 16'd45486, 16'd61451, 16'd14812});
	test_expansion(128'h07655ae49c0a62f3c9caf306e6414ac0, {16'd12333, 16'd716, 16'd26002, 16'd61125, 16'd20395, 16'd19124, 16'd42546, 16'd54868, 16'd19233, 16'd61833, 16'd1176, 16'd12236, 16'd36437, 16'd58798, 16'd25981, 16'd49570, 16'd56267, 16'd14043, 16'd4092, 16'd46637, 16'd42412, 16'd20223, 16'd21302, 16'd35041, 16'd40524, 16'd1375});
	test_expansion(128'h736ea8ccf96c5d45c64913caea078512, {16'd52827, 16'd20919, 16'd28947, 16'd1700, 16'd27830, 16'd25412, 16'd47082, 16'd31044, 16'd45208, 16'd27056, 16'd47064, 16'd7234, 16'd26997, 16'd34111, 16'd45783, 16'd47098, 16'd38979, 16'd30632, 16'd57769, 16'd30146, 16'd29180, 16'd54118, 16'd40011, 16'd4899, 16'd51406, 16'd14243});
	test_expansion(128'h0b66e22790726adcfd4e3cb07b0fd299, {16'd12820, 16'd18018, 16'd44427, 16'd32771, 16'd63708, 16'd10510, 16'd36784, 16'd43298, 16'd27600, 16'd30578, 16'd40013, 16'd53909, 16'd51087, 16'd51878, 16'd24341, 16'd26974, 16'd36520, 16'd25817, 16'd32442, 16'd63418, 16'd21224, 16'd11755, 16'd28808, 16'd41845, 16'd31333, 16'd45039});
	test_expansion(128'h4346a49ab7bd3573ef33de075d49fd7e, {16'd5412, 16'd38383, 16'd31311, 16'd44308, 16'd48835, 16'd51111, 16'd21998, 16'd28056, 16'd48912, 16'd18443, 16'd52897, 16'd45089, 16'd24282, 16'd30462, 16'd50354, 16'd25067, 16'd63493, 16'd43032, 16'd35415, 16'd28456, 16'd795, 16'd54003, 16'd49999, 16'd64648, 16'd42850, 16'd60573});
	test_expansion(128'h1d96a10edf32276c7a98ee994fd15c7d, {16'd53700, 16'd59497, 16'd8843, 16'd43228, 16'd36336, 16'd1257, 16'd15877, 16'd933, 16'd6113, 16'd51609, 16'd1740, 16'd35989, 16'd2656, 16'd19114, 16'd36926, 16'd17463, 16'd11034, 16'd19056, 16'd50809, 16'd9995, 16'd9505, 16'd48629, 16'd60007, 16'd51415, 16'd51834, 16'd29716});
	test_expansion(128'h1e50845dac6fc5fb20832d43d2fd3c4b, {16'd26345, 16'd16902, 16'd15692, 16'd20237, 16'd49780, 16'd38483, 16'd61755, 16'd12463, 16'd45531, 16'd9866, 16'd44657, 16'd58239, 16'd8301, 16'd49242, 16'd53176, 16'd39643, 16'd22281, 16'd55021, 16'd25037, 16'd40655, 16'd39908, 16'd56344, 16'd22031, 16'd21844, 16'd6359, 16'd11405});
	test_expansion(128'hb03e9ceb1e12ceb884ab3693d15a23af, {16'd13508, 16'd40250, 16'd17, 16'd14868, 16'd14670, 16'd23783, 16'd51985, 16'd7396, 16'd22410, 16'd48982, 16'd56203, 16'd4708, 16'd35787, 16'd54479, 16'd2482, 16'd3599, 16'd55704, 16'd36629, 16'd30657, 16'd26045, 16'd1547, 16'd5873, 16'd5693, 16'd8594, 16'd54125, 16'd21862});
	test_expansion(128'h278039b626b03a5654122aea4c5c6dc1, {16'd11876, 16'd16455, 16'd5819, 16'd42509, 16'd39237, 16'd519, 16'd52902, 16'd45745, 16'd37166, 16'd63936, 16'd6952, 16'd656, 16'd31169, 16'd53205, 16'd60702, 16'd8789, 16'd20744, 16'd17385, 16'd29962, 16'd44750, 16'd64098, 16'd12583, 16'd37094, 16'd40283, 16'd28989, 16'd25374});
	test_expansion(128'h1471a66d4af04114be83d4f171737e71, {16'd1777, 16'd14023, 16'd13836, 16'd29457, 16'd18990, 16'd63438, 16'd45779, 16'd15215, 16'd39707, 16'd23369, 16'd60549, 16'd6438, 16'd14596, 16'd34038, 16'd17536, 16'd35, 16'd34979, 16'd64452, 16'd23426, 16'd22495, 16'd51988, 16'd23376, 16'd30138, 16'd41868, 16'd44049, 16'd43415});
	test_expansion(128'hdc6db0a77ef74d21d58f9c314880ec32, {16'd3162, 16'd7849, 16'd16312, 16'd42776, 16'd27344, 16'd44578, 16'd57107, 16'd26891, 16'd14557, 16'd58556, 16'd2993, 16'd16455, 16'd55841, 16'd14355, 16'd12114, 16'd48086, 16'd33987, 16'd46482, 16'd64450, 16'd18606, 16'd40378, 16'd17078, 16'd704, 16'd65023, 16'd33193, 16'd30796});
	test_expansion(128'ha7584f119d4c757a3aafac7b3b45c6b0, {16'd58726, 16'd35733, 16'd27328, 16'd33326, 16'd1471, 16'd51466, 16'd59871, 16'd19016, 16'd24838, 16'd20820, 16'd47655, 16'd9194, 16'd10383, 16'd13085, 16'd59570, 16'd30526, 16'd46143, 16'd24296, 16'd53462, 16'd30059, 16'd34126, 16'd16735, 16'd35323, 16'd245, 16'd23620, 16'd35778});
	test_expansion(128'hb274e4932f639d383a28f1835503c9d2, {16'd62537, 16'd21779, 16'd15717, 16'd62499, 16'd37579, 16'd63218, 16'd23105, 16'd13758, 16'd45680, 16'd2726, 16'd10357, 16'd43343, 16'd43653, 16'd44371, 16'd17075, 16'd53127, 16'd38327, 16'd50419, 16'd34884, 16'd19105, 16'd16085, 16'd7501, 16'd61814, 16'd32692, 16'd55996, 16'd25006});
	test_expansion(128'h37550253845e13f8970a8bb423a11978, {16'd30450, 16'd63979, 16'd32826, 16'd46285, 16'd48013, 16'd19097, 16'd58874, 16'd51675, 16'd27977, 16'd63921, 16'd5101, 16'd41751, 16'd51719, 16'd29679, 16'd63105, 16'd11666, 16'd17700, 16'd50510, 16'd38560, 16'd9689, 16'd52971, 16'd50656, 16'd34063, 16'd30731, 16'd54178, 16'd5715});
	test_expansion(128'h088715065f46dc56209c1a6cc77906a5, {16'd65278, 16'd48893, 16'd15619, 16'd12710, 16'd7701, 16'd19130, 16'd56533, 16'd55212, 16'd18351, 16'd5410, 16'd64472, 16'd32308, 16'd56268, 16'd56413, 16'd34378, 16'd37525, 16'd17683, 16'd47099, 16'd57999, 16'd40613, 16'd48221, 16'd61602, 16'd19629, 16'd3984, 16'd27431, 16'd30359});
	test_expansion(128'h58278db1841f95994ab687cfae4806f2, {16'd24804, 16'd25301, 16'd46324, 16'd49719, 16'd55820, 16'd55716, 16'd24607, 16'd64562, 16'd40902, 16'd44926, 16'd7762, 16'd2993, 16'd11009, 16'd30823, 16'd22964, 16'd36519, 16'd46941, 16'd16939, 16'd11534, 16'd31696, 16'd58449, 16'd16196, 16'd33368, 16'd58551, 16'd30427, 16'd46396});
	test_expansion(128'h9ba85da30e3410900461fa69f1df0093, {16'd14989, 16'd61016, 16'd21068, 16'd61283, 16'd60407, 16'd50228, 16'd33195, 16'd33957, 16'd13968, 16'd50031, 16'd25446, 16'd32992, 16'd20944, 16'd49942, 16'd16951, 16'd57604, 16'd8710, 16'd5030, 16'd21650, 16'd54747, 16'd51931, 16'd42033, 16'd17722, 16'd23950, 16'd44401, 16'd38872});
	test_expansion(128'h6dee3c63a7137743201358dff381ffc1, {16'd65092, 16'd31787, 16'd40407, 16'd33147, 16'd49913, 16'd8516, 16'd64428, 16'd32553, 16'd6267, 16'd12234, 16'd45707, 16'd5777, 16'd9014, 16'd50218, 16'd48138, 16'd33371, 16'd29448, 16'd30598, 16'd45041, 16'd37655, 16'd49445, 16'd54339, 16'd38395, 16'd44266, 16'd11789, 16'd50006});
	test_expansion(128'hb71f1db7c5a3ea8a2e8b66b551bf8cda, {16'd50594, 16'd53337, 16'd11545, 16'd43966, 16'd49223, 16'd17587, 16'd33158, 16'd5992, 16'd26213, 16'd52448, 16'd20485, 16'd8616, 16'd42436, 16'd20414, 16'd49293, 16'd57119, 16'd57002, 16'd18254, 16'd27849, 16'd43504, 16'd37711, 16'd26204, 16'd44320, 16'd62366, 16'd29939, 16'd3654});
	test_expansion(128'hf3142943ffe97706f5a913fb7e299d55, {16'd41334, 16'd12186, 16'd43920, 16'd60537, 16'd45464, 16'd38942, 16'd52262, 16'd60696, 16'd14166, 16'd32514, 16'd31243, 16'd43837, 16'd36924, 16'd57613, 16'd36060, 16'd39376, 16'd32353, 16'd55255, 16'd3706, 16'd15943, 16'd50582, 16'd17071, 16'd48462, 16'd35793, 16'd42068, 16'd37434});
	test_expansion(128'h7c729bf9c50cdb501178723f5e23f025, {16'd41937, 16'd9065, 16'd35711, 16'd63017, 16'd45073, 16'd60920, 16'd4208, 16'd37930, 16'd37663, 16'd56559, 16'd56526, 16'd44818, 16'd22149, 16'd58255, 16'd32075, 16'd32262, 16'd53778, 16'd43636, 16'd14262, 16'd41824, 16'd58572, 16'd3757, 16'd48687, 16'd5990, 16'd47770, 16'd54835});
	test_expansion(128'h80e3c827d4afa99191c797e7df2c63b9, {16'd10683, 16'd386, 16'd15099, 16'd38909, 16'd14772, 16'd8641, 16'd19564, 16'd40538, 16'd38647, 16'd22795, 16'd29849, 16'd11459, 16'd174, 16'd23169, 16'd9284, 16'd32626, 16'd24510, 16'd29800, 16'd28534, 16'd34789, 16'd41981, 16'd9414, 16'd59240, 16'd33835, 16'd25959, 16'd36673});
	test_expansion(128'h7bdc949b5f465e7517b9be2a0b573a3d, {16'd60906, 16'd46381, 16'd46, 16'd28321, 16'd18986, 16'd43196, 16'd5645, 16'd8066, 16'd2021, 16'd34949, 16'd51280, 16'd33793, 16'd10600, 16'd14069, 16'd17163, 16'd32414, 16'd12621, 16'd2043, 16'd558, 16'd36507, 16'd4028, 16'd16079, 16'd11060, 16'd29997, 16'd17931, 16'd25087});
	test_expansion(128'h8e46abe058ab1123745d75f3992a46b5, {16'd62245, 16'd29232, 16'd10400, 16'd34649, 16'd22511, 16'd30174, 16'd2810, 16'd61384, 16'd33331, 16'd52841, 16'd20287, 16'd51403, 16'd43832, 16'd17628, 16'd56991, 16'd7939, 16'd14774, 16'd3532, 16'd27314, 16'd3431, 16'd52028, 16'd12951, 16'd40273, 16'd2490, 16'd59654, 16'd42177});
	test_expansion(128'h21d412f82b58b35a7c0ca2dbc3e6447d, {16'd53758, 16'd37584, 16'd25621, 16'd60698, 16'd30737, 16'd927, 16'd26385, 16'd56567, 16'd2313, 16'd46553, 16'd60704, 16'd22395, 16'd20008, 16'd34495, 16'd33361, 16'd48127, 16'd17175, 16'd50218, 16'd43415, 16'd50750, 16'd16018, 16'd35391, 16'd51894, 16'd44841, 16'd53428, 16'd39608});
	test_expansion(128'h53f1f27f53bc88d50e02fad51b310d89, {16'd64638, 16'd34012, 16'd45744, 16'd47973, 16'd26969, 16'd18887, 16'd32891, 16'd7165, 16'd25766, 16'd56696, 16'd62412, 16'd59015, 16'd43116, 16'd53892, 16'd700, 16'd37336, 16'd4394, 16'd17104, 16'd27618, 16'd63047, 16'd55443, 16'd21327, 16'd43855, 16'd57042, 16'd2499, 16'd52524});
	test_expansion(128'h5ed4878b70abbe93f296f4f25dcb1f2a, {16'd31529, 16'd57307, 16'd11575, 16'd40122, 16'd2579, 16'd63501, 16'd36034, 16'd873, 16'd13941, 16'd56103, 16'd30253, 16'd55072, 16'd55300, 16'd62683, 16'd15399, 16'd9901, 16'd3895, 16'd8595, 16'd39451, 16'd41433, 16'd36807, 16'd63223, 16'd22254, 16'd6597, 16'd14069, 16'd24189});
	test_expansion(128'ha05f5c18ee6c72534360bed6dd342034, {16'd64308, 16'd38421, 16'd1525, 16'd10223, 16'd9327, 16'd23049, 16'd51020, 16'd33252, 16'd50631, 16'd23731, 16'd44126, 16'd23777, 16'd13345, 16'd17179, 16'd48664, 16'd22475, 16'd12200, 16'd37638, 16'd40057, 16'd32539, 16'd372, 16'd11932, 16'd18797, 16'd14371, 16'd45125, 16'd46450});
	test_expansion(128'h024f1abaa04b13c749df6037d88c6b21, {16'd48970, 16'd28079, 16'd13068, 16'd8904, 16'd7014, 16'd52711, 16'd51081, 16'd40358, 16'd49750, 16'd9579, 16'd38779, 16'd36558, 16'd32208, 16'd49668, 16'd53699, 16'd9416, 16'd39113, 16'd22596, 16'd51541, 16'd29931, 16'd16964, 16'd40576, 16'd62606, 16'd53019, 16'd16716, 16'd4256});
	test_expansion(128'h0024f791b7c5d106dde860cf442762a1, {16'd48545, 16'd32245, 16'd34675, 16'd51940, 16'd8346, 16'd48235, 16'd9170, 16'd28651, 16'd63562, 16'd25538, 16'd46952, 16'd50861, 16'd51751, 16'd1433, 16'd4830, 16'd39387, 16'd25991, 16'd37789, 16'd29612, 16'd35986, 16'd29793, 16'd27761, 16'd61147, 16'd16428, 16'd19765, 16'd21346});
	test_expansion(128'hd27562d33124f1e04a7ae60d1fe02464, {16'd57932, 16'd9475, 16'd65428, 16'd45974, 16'd26610, 16'd43766, 16'd53876, 16'd39725, 16'd42458, 16'd62698, 16'd23125, 16'd40668, 16'd56795, 16'd24190, 16'd62607, 16'd40507, 16'd44800, 16'd57509, 16'd8352, 16'd28134, 16'd62455, 16'd1078, 16'd29985, 16'd13267, 16'd37242, 16'd667});
	test_expansion(128'hc46ed103113128978254da6b7583e02c, {16'd27604, 16'd42726, 16'd14463, 16'd6761, 16'd63889, 16'd30132, 16'd36766, 16'd60601, 16'd7481, 16'd29564, 16'd47303, 16'd2236, 16'd8754, 16'd31023, 16'd39732, 16'd33980, 16'd19136, 16'd11185, 16'd6530, 16'd26312, 16'd21240, 16'd40632, 16'd48772, 16'd7030, 16'd31899, 16'd61679});
	test_expansion(128'hbd3364675beea31b285b2143fc076f2a, {16'd53336, 16'd51380, 16'd1724, 16'd9209, 16'd15572, 16'd32374, 16'd7630, 16'd39960, 16'd2076, 16'd45868, 16'd54633, 16'd11184, 16'd55361, 16'd13730, 16'd44717, 16'd86, 16'd59018, 16'd34801, 16'd12377, 16'd49764, 16'd44676, 16'd61721, 16'd2304, 16'd846, 16'd6708, 16'd8525});
	test_expansion(128'he8dd4c3bd148b27736925d4c216c6a18, {16'd47720, 16'd34980, 16'd58681, 16'd11236, 16'd35974, 16'd57946, 16'd1242, 16'd1842, 16'd49583, 16'd14857, 16'd63963, 16'd30619, 16'd24812, 16'd10587, 16'd23830, 16'd62227, 16'd51495, 16'd17685, 16'd14928, 16'd34744, 16'd50890, 16'd32463, 16'd2800, 16'd36989, 16'd28205, 16'd25336});
	test_expansion(128'hf63dd0e1abe3d99d0332e22c88d69a75, {16'd59890, 16'd10393, 16'd32055, 16'd19376, 16'd21461, 16'd59608, 16'd45155, 16'd52244, 16'd47846, 16'd36772, 16'd7293, 16'd11615, 16'd26755, 16'd25562, 16'd6357, 16'd25863, 16'd19738, 16'd39677, 16'd64403, 16'd35943, 16'd13059, 16'd24421, 16'd37267, 16'd20966, 16'd28189, 16'd32625});
	test_expansion(128'hdfca83c469e27fec456f2238f137e467, {16'd35282, 16'd16591, 16'd20538, 16'd52122, 16'd46811, 16'd43360, 16'd45092, 16'd3545, 16'd13782, 16'd16303, 16'd28781, 16'd9675, 16'd46295, 16'd47241, 16'd24033, 16'd58942, 16'd25958, 16'd37717, 16'd25910, 16'd46094, 16'd20723, 16'd32676, 16'd3137, 16'd34670, 16'd40204, 16'd1459});
	test_expansion(128'hbb14b4823419275497a72e97b39e2073, {16'd15143, 16'd12435, 16'd50402, 16'd2368, 16'd22052, 16'd52173, 16'd56725, 16'd17726, 16'd19170, 16'd37948, 16'd26456, 16'd48809, 16'd51558, 16'd35581, 16'd33399, 16'd63189, 16'd20878, 16'd14176, 16'd32227, 16'd685, 16'd49328, 16'd35356, 16'd59315, 16'd19541, 16'd23213, 16'd17028});
	test_expansion(128'h7bc07128829d5e784e1cfff097ca6134, {16'd58080, 16'd53370, 16'd63701, 16'd22795, 16'd50078, 16'd15802, 16'd1684, 16'd32388, 16'd49151, 16'd65030, 16'd24570, 16'd50898, 16'd56219, 16'd15401, 16'd29952, 16'd6738, 16'd10284, 16'd31979, 16'd20052, 16'd38572, 16'd62741, 16'd56952, 16'd31194, 16'd17752, 16'd40204, 16'd29127});
	test_expansion(128'h2ead1d5ecc0b0cf7bd2a38f55f946b2f, {16'd23191, 16'd50023, 16'd33809, 16'd52553, 16'd28861, 16'd36227, 16'd58612, 16'd51843, 16'd12861, 16'd10178, 16'd21010, 16'd59207, 16'd33002, 16'd44936, 16'd29497, 16'd36082, 16'd25466, 16'd17890, 16'd16503, 16'd34283, 16'd40348, 16'd64774, 16'd22182, 16'd12315, 16'd65162, 16'd13232});
	test_expansion(128'hb4254d0aba7613fefa521bb17229c539, {16'd35320, 16'd28452, 16'd22475, 16'd43966, 16'd31375, 16'd34063, 16'd59058, 16'd63547, 16'd48741, 16'd56216, 16'd19111, 16'd7355, 16'd11056, 16'd58413, 16'd28620, 16'd61334, 16'd64725, 16'd10933, 16'd36508, 16'd39016, 16'd14238, 16'd411, 16'd33879, 16'd63025, 16'd11519, 16'd61890});
	test_expansion(128'hb6df815dd4dfd57dcd6da0d909e7ed22, {16'd59867, 16'd43331, 16'd16898, 16'd11170, 16'd16707, 16'd61271, 16'd54516, 16'd30873, 16'd45175, 16'd4267, 16'd32835, 16'd33598, 16'd42345, 16'd24165, 16'd25470, 16'd58358, 16'd31146, 16'd15012, 16'd58831, 16'd7274, 16'd9725, 16'd60878, 16'd54771, 16'd8198, 16'd52156, 16'd16682});
	test_expansion(128'he0e7341597b555cc2b2ab59536dea703, {16'd55824, 16'd53041, 16'd46885, 16'd20326, 16'd11893, 16'd42940, 16'd30589, 16'd31379, 16'd63085, 16'd6874, 16'd1648, 16'd15338, 16'd12045, 16'd8650, 16'd12916, 16'd65033, 16'd27394, 16'd48170, 16'd40956, 16'd29613, 16'd14318, 16'd48571, 16'd57277, 16'd50541, 16'd42773, 16'd50932});
	test_expansion(128'h49ecba68d942c07950822f9fdcc42719, {16'd59021, 16'd54939, 16'd5279, 16'd64744, 16'd16258, 16'd62548, 16'd42880, 16'd64840, 16'd3477, 16'd56590, 16'd11329, 16'd64865, 16'd13880, 16'd15290, 16'd58768, 16'd11014, 16'd30250, 16'd31357, 16'd30766, 16'd11115, 16'd48888, 16'd35913, 16'd13437, 16'd44398, 16'd62965, 16'd45105});
	test_expansion(128'h739cb58440fc26fccb124b9cbeb17f04, {16'd40390, 16'd44483, 16'd6249, 16'd59385, 16'd64389, 16'd47072, 16'd3941, 16'd39512, 16'd11681, 16'd32482, 16'd4601, 16'd62174, 16'd31483, 16'd27401, 16'd52813, 16'd30453, 16'd65483, 16'd57845, 16'd61561, 16'd28603, 16'd65077, 16'd13872, 16'd49479, 16'd31912, 16'd25756, 16'd28804});
	test_expansion(128'h8a586f7f8de54827891bff683da31d9c, {16'd44731, 16'd29584, 16'd35109, 16'd65041, 16'd65221, 16'd1049, 16'd54412, 16'd53535, 16'd63154, 16'd11921, 16'd62562, 16'd49880, 16'd63095, 16'd35191, 16'd32159, 16'd45644, 16'd20381, 16'd65248, 16'd6034, 16'd51320, 16'd35663, 16'd21567, 16'd8390, 16'd62217, 16'd19951, 16'd35489});
	test_expansion(128'h2114f2dae26b40252d1faadb5bfcb6a3, {16'd41699, 16'd29413, 16'd55536, 16'd45373, 16'd26753, 16'd875, 16'd15853, 16'd28644, 16'd22336, 16'd25010, 16'd36196, 16'd34012, 16'd39392, 16'd23873, 16'd15469, 16'd15140, 16'd28158, 16'd14537, 16'd3817, 16'd18395, 16'd45790, 16'd20909, 16'd41430, 16'd39575, 16'd19650, 16'd23220});
	test_expansion(128'h9fba95339ef445e363ef6a919ef4e42b, {16'd55027, 16'd49906, 16'd48930, 16'd32703, 16'd35206, 16'd61840, 16'd25949, 16'd7117, 16'd4661, 16'd43704, 16'd57099, 16'd62413, 16'd38989, 16'd5571, 16'd2671, 16'd18231, 16'd45901, 16'd52758, 16'd29445, 16'd22674, 16'd9981, 16'd34989, 16'd53920, 16'd6529, 16'd17323, 16'd11399});
	test_expansion(128'h166eb7236081dc53626b329e8b0a90d5, {16'd19724, 16'd2028, 16'd12447, 16'd65226, 16'd27178, 16'd35057, 16'd30361, 16'd2249, 16'd53143, 16'd1796, 16'd54815, 16'd45699, 16'd46758, 16'd43702, 16'd43771, 16'd58005, 16'd42018, 16'd13678, 16'd35810, 16'd36064, 16'd9106, 16'd11089, 16'd62920, 16'd60049, 16'd28877, 16'd340});
	test_expansion(128'h6c8dfb2eb2033c2d5a347a67989b9ecb, {16'd62558, 16'd32082, 16'd54667, 16'd18271, 16'd56961, 16'd37051, 16'd58947, 16'd1451, 16'd65436, 16'd41894, 16'd7682, 16'd40165, 16'd6786, 16'd38207, 16'd51588, 16'd16967, 16'd50559, 16'd44935, 16'd45427, 16'd58052, 16'd39381, 16'd48273, 16'd36308, 16'd54469, 16'd39627, 16'd10937});
	test_expansion(128'hf913b12eac1cce0e2ded4514199ec1e1, {16'd14820, 16'd46043, 16'd59652, 16'd26483, 16'd8712, 16'd8993, 16'd2377, 16'd199, 16'd2914, 16'd48703, 16'd26129, 16'd187, 16'd29915, 16'd6279, 16'd16648, 16'd44091, 16'd11973, 16'd40589, 16'd37643, 16'd16510, 16'd25641, 16'd64911, 16'd18684, 16'd61475, 16'd39194, 16'd64209});
	test_expansion(128'ha0c29a89fdcd08c6e30404abbeb20b3c, {16'd12782, 16'd10553, 16'd28216, 16'd44760, 16'd5597, 16'd5526, 16'd28879, 16'd7222, 16'd16694, 16'd35521, 16'd33135, 16'd11032, 16'd55411, 16'd53732, 16'd12275, 16'd45525, 16'd40088, 16'd58016, 16'd42866, 16'd22570, 16'd34676, 16'd40653, 16'd5613, 16'd248, 16'd7842, 16'd31281});
	test_expansion(128'h53eeecf75d8fae67d22d449cf25bbe55, {16'd38697, 16'd18884, 16'd38187, 16'd29221, 16'd63662, 16'd8812, 16'd24948, 16'd41274, 16'd40367, 16'd17127, 16'd51285, 16'd20165, 16'd41011, 16'd12638, 16'd44400, 16'd59865, 16'd32739, 16'd23704, 16'd19920, 16'd22896, 16'd7443, 16'd60673, 16'd1730, 16'd50529, 16'd8344, 16'd51387});
	test_expansion(128'hf69b39f704e69f7545121eab622a8b9a, {16'd23291, 16'd59093, 16'd3109, 16'd57358, 16'd41201, 16'd19565, 16'd50280, 16'd38372, 16'd58491, 16'd63048, 16'd42335, 16'd33739, 16'd28344, 16'd54809, 16'd27476, 16'd65314, 16'd55304, 16'd16379, 16'd30070, 16'd732, 16'd37717, 16'd34714, 16'd6491, 16'd22743, 16'd6541, 16'd993});
	test_expansion(128'hcdeede34af4696ceaa9e62564165874f, {16'd21797, 16'd16746, 16'd24633, 16'd14460, 16'd31173, 16'd31440, 16'd13125, 16'd55954, 16'd7921, 16'd42310, 16'd10915, 16'd24496, 16'd12579, 16'd48793, 16'd37283, 16'd51107, 16'd61796, 16'd51663, 16'd17040, 16'd59839, 16'd42974, 16'd636, 16'd35290, 16'd53020, 16'd36724, 16'd41359});
	test_expansion(128'h4e6de9297cfb64380d31ab63883bef07, {16'd57872, 16'd8609, 16'd45516, 16'd8613, 16'd58705, 16'd22381, 16'd46317, 16'd51650, 16'd38286, 16'd11006, 16'd15350, 16'd5958, 16'd13179, 16'd40442, 16'd33437, 16'd47079, 16'd8532, 16'd38046, 16'd13708, 16'd14535, 16'd29241, 16'd31427, 16'd7684, 16'd40845, 16'd62914, 16'd36638});
	test_expansion(128'h51763474d21eb71433e7343c252f7cf5, {16'd41822, 16'd37110, 16'd3248, 16'd45332, 16'd42957, 16'd23049, 16'd2519, 16'd39738, 16'd42130, 16'd55204, 16'd40428, 16'd23163, 16'd43817, 16'd45098, 16'd33946, 16'd28672, 16'd17440, 16'd60982, 16'd16758, 16'd48499, 16'd13500, 16'd64306, 16'd13430, 16'd46907, 16'd20554, 16'd62311});
	test_expansion(128'h5c47931b18182d4e7ee0a6578a1d8d64, {16'd33442, 16'd43967, 16'd40646, 16'd37999, 16'd38743, 16'd40571, 16'd41526, 16'd55078, 16'd65199, 16'd33479, 16'd41139, 16'd14019, 16'd49068, 16'd32078, 16'd56794, 16'd26503, 16'd13935, 16'd37178, 16'd7012, 16'd28470, 16'd28099, 16'd15143, 16'd49731, 16'd58668, 16'd6987, 16'd29568});
	test_expansion(128'haaadd082c7a355c7005dc3a627c5949c, {16'd40580, 16'd4517, 16'd11840, 16'd15414, 16'd27326, 16'd53237, 16'd59708, 16'd65319, 16'd41309, 16'd33324, 16'd21676, 16'd3587, 16'd43196, 16'd51394, 16'd59648, 16'd13059, 16'd30622, 16'd19555, 16'd19206, 16'd41323, 16'd37932, 16'd63872, 16'd43892, 16'd51110, 16'd36315, 16'd29307});
	test_expansion(128'h2afe320b357365fcc266c6321d0c6e6a, {16'd53632, 16'd42, 16'd34147, 16'd18747, 16'd478, 16'd43651, 16'd1153, 16'd40554, 16'd58112, 16'd29169, 16'd18677, 16'd44109, 16'd20017, 16'd56643, 16'd48271, 16'd10816, 16'd2850, 16'd56359, 16'd23182, 16'd8742, 16'd46211, 16'd1908, 16'd36633, 16'd24675, 16'd18277, 16'd502});
	test_expansion(128'h0860dd824e5d8609a95cb422b9ec4a05, {16'd1591, 16'd61119, 16'd14161, 16'd17142, 16'd4411, 16'd36462, 16'd10291, 16'd45221, 16'd16321, 16'd63383, 16'd21002, 16'd57874, 16'd18374, 16'd51518, 16'd58517, 16'd14988, 16'd64657, 16'd29882, 16'd7217, 16'd33810, 16'd59490, 16'd23668, 16'd3927, 16'd54109, 16'd33670, 16'd62188});
	test_expansion(128'hec28495964d6cbf6a61d1a07c86be09a, {16'd34722, 16'd42688, 16'd15439, 16'd59922, 16'd42682, 16'd54950, 16'd10885, 16'd7318, 16'd27358, 16'd15706, 16'd33954, 16'd63697, 16'd2100, 16'd51108, 16'd61709, 16'd27247, 16'd35572, 16'd27278, 16'd57509, 16'd55292, 16'd49260, 16'd28674, 16'd14445, 16'd36765, 16'd39581, 16'd37760});
	test_expansion(128'h446b1be7e41934775da869bec1783a65, {16'd540, 16'd56741, 16'd51493, 16'd26921, 16'd43801, 16'd21285, 16'd56429, 16'd37610, 16'd31749, 16'd4600, 16'd105, 16'd53264, 16'd28840, 16'd5040, 16'd26340, 16'd10261, 16'd3818, 16'd29391, 16'd17720, 16'd56516, 16'd11326, 16'd5397, 16'd60052, 16'd44073, 16'd237, 16'd8157});
	test_expansion(128'hb845da889978116a4fe2b30f0c483835, {16'd47582, 16'd56987, 16'd46061, 16'd25210, 16'd37681, 16'd33704, 16'd53696, 16'd14190, 16'd45693, 16'd19210, 16'd5913, 16'd64702, 16'd33771, 16'd29944, 16'd54596, 16'd33167, 16'd51942, 16'd15151, 16'd49696, 16'd6284, 16'd26947, 16'd47166, 16'd41950, 16'd53141, 16'd44580, 16'd19587});
	test_expansion(128'h1c1ec9702c35560ba3b74f2d233b3e7a, {16'd57570, 16'd24120, 16'd42503, 16'd41215, 16'd61169, 16'd29222, 16'd33984, 16'd65173, 16'd33826, 16'd13816, 16'd29489, 16'd36820, 16'd59721, 16'd62942, 16'd18103, 16'd24600, 16'd58834, 16'd57216, 16'd54765, 16'd61975, 16'd36136, 16'd58563, 16'd58524, 16'd10494, 16'd64546, 16'd2012});
	test_expansion(128'he0a7cc682a0c7c67cc1a7ceac89786be, {16'd23782, 16'd54448, 16'd36682, 16'd23993, 16'd19152, 16'd37679, 16'd18416, 16'd30935, 16'd11063, 16'd64734, 16'd33253, 16'd14282, 16'd8372, 16'd54223, 16'd47545, 16'd39400, 16'd5447, 16'd31796, 16'd51925, 16'd31566, 16'd9695, 16'd17841, 16'd41441, 16'd1368, 16'd53464, 16'd9708});


	`endif

    $display("SUCCESS :: FINISH CALLED FROM END OF FILE!");
    $finish;

end


endmodule

