
`define W_size 16 // word size (PARAMETER)
`define K_size 128 // Key size (PARAMETER)
`define U 2 // W_size/2
`define T 26 // 2*(number of rounds + 1)
`define B 16 // key size in bytes
`define C 8 // c=b/u=16/2=8
`define P 16'hb7e1
`define Q 16'h9e37

// UNCOMMENT THIS DEFINE FOR ALL 10,000 TEST CASES!!!!
`define FULL

`timescale 1ns / 1ps
module key_tb;

logic start;
logic clk;
logic rst;
logic [128:0] key;
logic [`W_size-1:0] sub [0:`T-1];
logic [4:0] num_rounds;
logic ready;

assign num_rounds = 12;

keygen Keygen(.*);

default clocking ckb @(posedge clk);
    input sub, ready;
    output rst, key, start;
endclocking

always begin
    clk = 1'b0;
    #1;
    clk = 1'b1;
    #1;
end

task reset();
    rst <= 1;
    ##1;
    rst <= 0;
    ##1;
endtask

task test_expansion(logic[`K_size-1:0] test_key, logic [`W_size-1:0] test_subkey [0:`T-1]);
    key <= test_key;

    ##1;

    start <= 1;
    ##1;

    start <= 0;

    while(~ready) begin
        ##1;
    end

    for(int i = 0; i < `T; i++) begin
        assert(test_subkey[i] == sub[i])
            else begin
                $error("Bad Subkey Value: 0x%x at position %0d, should be 0x%x", sub[i], i, test_subkey[i]);
                $finish;
            end
    end
endtask

initial begin
    $fsdbDumpfile("dump.fsdb");
	$fsdbDumpvars(0, "+all");
    key <= 0;
    rst <= 0;
    start <= 0;

    #2;

    reset();

    // Known Test Case
	test_expansion(128'hdeadbeefdeadbeefdeadbeefdeadbeef, {16'd55048, 16'd43744, 16'd48559, 16'd27403, 16'd20374, 16'd33387, 16'd2062, 16'd61013, 16'd49237, 16'd33709, 16'd16278, 16'd65452, 16'd9968, 16'd4572, 16'd34933, 16'd35205, 16'd37470, 16'd42119, 16'd21025, 16'd13567, 16'd19718, 16'd1446, 16'd11664, 16'd40137, 16'd19576, 16'd15720});

    // AUTO GENERATED TEST CASES
	`ifdef FULL

	test_expansion(128'h701d6ca4b5f9cb6eec751243d4fc4117, {16'd53001, 16'd41195, 16'd15524, 16'd53014, 16'd57831, 16'd30487, 16'd21534, 16'd1969, 16'd17535, 16'd35736, 16'd26089, 16'd38976, 16'd9380, 16'd18481, 16'd16318, 16'd62818, 16'd28387, 16'd4160, 16'd20782, 16'd54929, 16'd51509, 16'd59820, 16'd21353, 16'd53083, 16'd31851, 16'd33526});
	test_expansion(128'h0d21f7a29d740da69d94cebae90a73b2, {16'd17926, 16'd52683, 16'd13645, 16'd7564, 16'd58736, 16'd18045, 16'd59198, 16'd25906, 16'd9342, 16'd48639, 16'd36978, 16'd18734, 16'd32236, 16'd54457, 16'd19974, 16'd19623, 16'd59254, 16'd41762, 16'd10718, 16'd916, 16'd38591, 16'd58888, 16'd27719, 16'd39913, 16'd41828, 16'd60178});
	test_expansion(128'h77c0d6190c1c2b373bc0b14535ed89e9, {16'd46994, 16'd22149, 16'd20758, 16'd59893, 16'd51182, 16'd32385, 16'd11793, 16'd59150, 16'd5574, 16'd38406, 16'd17297, 16'd8676, 16'd57008, 16'd34660, 16'd524, 16'd38344, 16'd56945, 16'd5192, 16'd16327, 16'd18444, 16'd10570, 16'd19965, 16'd58431, 16'd39748, 16'd51671, 16'd57769});
	test_expansion(128'h116176d9ce32c83a996a2cc77ec37fb9, {16'd17268, 16'd54786, 16'd37501, 16'd40859, 16'd17280, 16'd27520, 16'd33014, 16'd35596, 16'd43511, 16'd19408, 16'd2029, 16'd25654, 16'd15120, 16'd17139, 16'd47974, 16'd57737, 16'd26941, 16'd24712, 16'd22487, 16'd5394, 16'd59541, 16'd61245, 16'd756, 16'd18141, 16'd41711, 16'd42750});
	test_expansion(128'h9e07c3998c046ca959b5546dd9ce800a, {16'd26544, 16'd6641, 16'd5066, 16'd39243, 16'd17682, 16'd30543, 16'd4705, 16'd43107, 16'd23026, 16'd6917, 16'd31870, 16'd44151, 16'd8619, 16'd20294, 16'd34043, 16'd61960, 16'd45392, 16'd36101, 16'd53113, 16'd40970, 16'd63243, 16'd21806, 16'd24087, 16'd42679, 16'd58683, 16'd28112});
	test_expansion(128'h49cb7022bc6cbedc8033b5820e44fcbb, {16'd50583, 16'd35686, 16'd39522, 16'd4106, 16'd17634, 16'd14875, 16'd20384, 16'd26364, 16'd3464, 16'd4516, 16'd24832, 16'd11372, 16'd29070, 16'd24096, 16'd55526, 16'd13618, 16'd39609, 16'd1567, 16'd18041, 16'd27881, 16'd56325, 16'd19849, 16'd28708, 16'd27638, 16'd700, 16'd28842});
	test_expansion(128'he6ac47a99e4b141fc620d589a028f90e, {16'd35221, 16'd859, 16'd44919, 16'd42679, 16'd45616, 16'd18478, 16'd2440, 16'd7922, 16'd23587, 16'd37796, 16'd34153, 16'd59681, 16'd392, 16'd40091, 16'd17044, 16'd52362, 16'd24483, 16'd57687, 16'd56863, 16'd29629, 16'd5164, 16'd44388, 16'd46699, 16'd36651, 16'd60099, 16'd13407});
	test_expansion(128'hf6922cd155e15d281c7a77ef51ef6958, {16'd43618, 16'd36950, 16'd59638, 16'd22708, 16'd54404, 16'd62250, 16'd29633, 16'd40263, 16'd1321, 16'd60032, 16'd49937, 16'd48755, 16'd54971, 16'd1735, 16'd31463, 16'd4415, 16'd11992, 16'd59379, 16'd31209, 16'd12984, 16'd4535, 16'd62682, 16'd17962, 16'd37900, 16'd41466, 16'd554});
	test_expansion(128'he0b0ff112d3f0df7b52d024f85049142, {16'd14774, 16'd16242, 16'd2379, 16'd22218, 16'd652, 16'd54388, 16'd62260, 16'd31331, 16'd1879, 16'd59418, 16'd60742, 16'd2367, 16'd46433, 16'd14843, 16'd29558, 16'd20773, 16'd41754, 16'd49279, 16'd46535, 16'd43135, 16'd9381, 16'd52961, 16'd1499, 16'd6373, 16'd7544, 16'd7468});
	test_expansion(128'h6372e18787d5b6bc387050a510febc71, {16'd50914, 16'd41712, 16'd61138, 16'd13080, 16'd27120, 16'd19056, 16'd37777, 16'd15715, 16'd15350, 16'd53118, 16'd40408, 16'd4122, 16'd12496, 16'd34096, 16'd59369, 16'd49418, 16'd48066, 16'd2324, 16'd30268, 16'd5359, 16'd34193, 16'd50736, 16'd3126, 16'd4705, 16'd47923, 16'd1847});
	test_expansion(128'h551e354291a1291ce93e23932a80390d, {16'd64187, 16'd48888, 16'd20910, 16'd40587, 16'd2701, 16'd63619, 16'd2459, 16'd46816, 16'd50206, 16'd34683, 16'd60041, 16'd2191, 16'd51985, 16'd37296, 16'd47755, 16'd22185, 16'd64807, 16'd60084, 16'd60141, 16'd14574, 16'd7295, 16'd640, 16'd16612, 16'd15676, 16'd8428, 16'd35652});
	test_expansion(128'hd2cae861da148671fb477d37272d1868, {16'd64125, 16'd2228, 16'd47838, 16'd11569, 16'd25682, 16'd15874, 16'd60980, 16'd9763, 16'd48738, 16'd426, 16'd20591, 16'd32317, 16'd23633, 16'd20275, 16'd20047, 16'd36695, 16'd27328, 16'd22236, 16'd36297, 16'd9969, 16'd11577, 16'd55797, 16'd51447, 16'd56436, 16'd1113, 16'd9358});
	test_expansion(128'h8f64f7f9e454da3939fc19a237d34022, {16'd31052, 16'd51930, 16'd5661, 16'd18521, 16'd63275, 16'd54941, 16'd43933, 16'd22762, 16'd62269, 16'd58929, 16'd59835, 16'd44224, 16'd54752, 16'd65078, 16'd50856, 16'd30701, 16'd47116, 16'd5762, 16'd17583, 16'd33724, 16'd6470, 16'd62473, 16'd44918, 16'd20467, 16'd41067, 16'd35348});
	test_expansion(128'hb46ff9ef8889097496859605438e1ee3, {16'd7300, 16'd16416, 16'd61640, 16'd25897, 16'd34134, 16'd58251, 16'd1031, 16'd6095, 16'd37477, 16'd28617, 16'd47279, 16'd31468, 16'd27930, 16'd32748, 16'd64769, 16'd59480, 16'd8008, 16'd25427, 16'd52627, 16'd37233, 16'd9274, 16'd28369, 16'd28255, 16'd43663, 16'd18659, 16'd16421});
	test_expansion(128'h8bcd68a2327c52b4b0674d289aa43bef, {16'd26933, 16'd51001, 16'd38109, 16'd13152, 16'd23844, 16'd32386, 16'd41646, 16'd30774, 16'd30897, 16'd28696, 16'd26566, 16'd62674, 16'd11155, 16'd38468, 16'd39125, 16'd23956, 16'd14420, 16'd14430, 16'd25425, 16'd59822, 16'd42640, 16'd46484, 16'd6993, 16'd60245, 16'd54208, 16'd37121});
	test_expansion(128'ha5454a0a6be4aaaedbb1c54689da8304, {16'd37291, 16'd62679, 16'd36135, 16'd64927, 16'd20336, 16'd57471, 16'd49561, 16'd44647, 16'd21506, 16'd44984, 16'd25639, 16'd10182, 16'd29677, 16'd24239, 16'd4886, 16'd44632, 16'd65216, 16'd48657, 16'd22964, 16'd50850, 16'd65018, 16'd55002, 16'd8424, 16'd4355, 16'd35009, 16'd6105});
	test_expansion(128'h828f308c0830b66a677de612c7609225, {16'd65304, 16'd20359, 16'd26408, 16'd22271, 16'd24869, 16'd63804, 16'd31442, 16'd35217, 16'd15152, 16'd40789, 16'd17317, 16'd14786, 16'd34487, 16'd10375, 16'd53835, 16'd43148, 16'd29208, 16'd10247, 16'd22222, 16'd36392, 16'd1513, 16'd54676, 16'd59574, 16'd53667, 16'd46928, 16'd53468});
	test_expansion(128'hf02ee46c868532f19dc4605538656768, {16'd6779, 16'd16600, 16'd39394, 16'd61297, 16'd46230, 16'd36696, 16'd19605, 16'd15351, 16'd56757, 16'd55844, 16'd45212, 16'd19549, 16'd56278, 16'd35352, 16'd33325, 16'd52939, 16'd1688, 16'd5897, 16'd45946, 16'd39673, 16'd45287, 16'd3972, 16'd34266, 16'd560, 16'd54886, 16'd14150});
	test_expansion(128'h14e2e85167ecc171ab24a262b9c9d4fb, {16'd19424, 16'd51992, 16'd58138, 16'd58450, 16'd52152, 16'd56447, 16'd55537, 16'd19895, 16'd6290, 16'd33731, 16'd49747, 16'd25616, 16'd65474, 16'd10441, 16'd22106, 16'd20213, 16'd34457, 16'd56006, 16'd44789, 16'd64826, 16'd49910, 16'd6922, 16'd61529, 16'd16337, 16'd49443, 16'd25919});
	test_expansion(128'h3bca7a58d9724da5801e6cf06a8653f7, {16'd34997, 16'd6055, 16'd39067, 16'd14999, 16'd2469, 16'd6046, 16'd14252, 16'd26868, 16'd14483, 16'd33312, 16'd1981, 16'd36869, 16'd45465, 16'd50385, 16'd65400, 16'd1585, 16'd32815, 16'd25135, 16'd64606, 16'd62885, 16'd25775, 16'd59480, 16'd6323, 16'd31692, 16'd25145, 16'd5173});
	test_expansion(128'h8342bd6627f5fd9ffa8b0d8b3058321b, {16'd42911, 16'd56418, 16'd47640, 16'd23601, 16'd1424, 16'd9008, 16'd38636, 16'd31482, 16'd48819, 16'd41195, 16'd2349, 16'd28421, 16'd30418, 16'd1283, 16'd1467, 16'd39189, 16'd36241, 16'd26801, 16'd23232, 16'd2681, 16'd51180, 16'd22019, 16'd15769, 16'd61231, 16'd58472, 16'd39964});
	test_expansion(128'h04cce75c7c059dd2d70bbdc679d6f4c2, {16'd26179, 16'd44209, 16'd50147, 16'd4244, 16'd6929, 16'd21550, 16'd19909, 16'd21281, 16'd62546, 16'd25401, 16'd37324, 16'd30871, 16'd13584, 16'd50880, 16'd22010, 16'd47048, 16'd28415, 16'd11072, 16'd22865, 16'd27107, 16'd8869, 16'd11804, 16'd50322, 16'd47912, 16'd27715, 16'd57401});
	test_expansion(128'hf27eedf1ec3dff3c19ea1370a2ce01c5, {16'd29716, 16'd7578, 16'd12263, 16'd42368, 16'd27194, 16'd62463, 16'd51639, 16'd61908, 16'd40737, 16'd61658, 16'd56988, 16'd15795, 16'd35612, 16'd32356, 16'd8817, 16'd12125, 16'd47008, 16'd10378, 16'd40074, 16'd25821, 16'd43079, 16'd37730, 16'd61029, 16'd37666, 16'd64256, 16'd58074});
	test_expansion(128'haf3c689f2e656c3112b5627e0d397301, {16'd53381, 16'd63442, 16'd32294, 16'd29257, 16'd731, 16'd28456, 16'd1961, 16'd14871, 16'd23287, 16'd15995, 16'd28856, 16'd55392, 16'd38332, 16'd19685, 16'd33105, 16'd16653, 16'd44877, 16'd16841, 16'd42681, 16'd11961, 16'd9221, 16'd52922, 16'd10709, 16'd23102, 16'd39112, 16'd51509});
	test_expansion(128'he9569ef7a60878007564e786ecc72ae3, {16'd8637, 16'd36151, 16'd10946, 16'd47595, 16'd18086, 16'd17968, 16'd5978, 16'd32345, 16'd8548, 16'd3983, 16'd4314, 16'd35837, 16'd41744, 16'd57892, 16'd13935, 16'd35543, 16'd50673, 16'd64563, 16'd56059, 16'd22323, 16'd24539, 16'd3344, 16'd39088, 16'd38827, 16'd23496, 16'd19040});
	test_expansion(128'hd335edb551e21a6ea115024cd833252c, {16'd38123, 16'd52324, 16'd65315, 16'd44918, 16'd21012, 16'd9412, 16'd52775, 16'd48035, 16'd63175, 16'd24763, 16'd34104, 16'd7884, 16'd50304, 16'd48466, 16'd44002, 16'd25, 16'd65201, 16'd21895, 16'd62817, 16'd537, 16'd23071, 16'd38403, 16'd34247, 16'd50330, 16'd56614, 16'd35130});
	test_expansion(128'h3618141da0559b34b6edeb095e6a4b85, {16'd7272, 16'd16602, 16'd3118, 16'd46083, 16'd60718, 16'd43589, 16'd17482, 16'd17712, 16'd11002, 16'd8063, 16'd296, 16'd36028, 16'd53034, 16'd21602, 16'd8972, 16'd36328, 16'd22958, 16'd60280, 16'd51338, 16'd22471, 16'd46869, 16'd32342, 16'd38544, 16'd1479, 16'd51152, 16'd59514});
	test_expansion(128'h9a2b638f1ae7ced17e5ac02739ad0988, {16'd5139, 16'd20524, 16'd61207, 16'd44865, 16'd60516, 16'd42429, 16'd39807, 16'd7962, 16'd18583, 16'd53488, 16'd17476, 16'd15513, 16'd2113, 16'd47980, 16'd41301, 16'd12566, 16'd36816, 16'd58631, 16'd29177, 16'd18269, 16'd36498, 16'd24974, 16'd1166, 16'd21666, 16'd54001, 16'd39117});
	test_expansion(128'hdd9aca7be1a096f7914b16fc7cb765f7, {16'd29047, 16'd48821, 16'd12617, 16'd57466, 16'd53990, 16'd52456, 16'd2475, 16'd55204, 16'd64262, 16'd47691, 16'd8000, 16'd9655, 16'd60321, 16'd64473, 16'd7336, 16'd65389, 16'd35591, 16'd26615, 16'd44494, 16'd14477, 16'd17733, 16'd19824, 16'd46900, 16'd25102, 16'd48759, 16'd65443});
	test_expansion(128'h4b09b0c839eabb77d8161d3ba952f711, {16'd61654, 16'd22836, 16'd58117, 16'd56031, 16'd64600, 16'd16210, 16'd12295, 16'd49449, 16'd48347, 16'd51709, 16'd38630, 16'd19538, 16'd33324, 16'd59674, 16'd50676, 16'd7417, 16'd35781, 16'd58438, 16'd1556, 16'd57266, 16'd42760, 16'd17613, 16'd34835, 16'd56828, 16'd61590, 16'd27703});
	test_expansion(128'h6375aef07a74e4fff22847935b02148b, {16'd21335, 16'd5812, 16'd10292, 16'd23834, 16'd10407, 16'd17062, 16'd56790, 16'd32830, 16'd37502, 16'd57244, 16'd56817, 16'd28216, 16'd50671, 16'd17368, 16'd59128, 16'd51255, 16'd6502, 16'd34556, 16'd39847, 16'd31048, 16'd56556, 16'd38004, 16'd33145, 16'd54341, 16'd50327, 16'd30164});
	test_expansion(128'h1775acd543db1136aa5c6add70bbb564, {16'd60714, 16'd13801, 16'd28124, 16'd17744, 16'd19733, 16'd5051, 16'd382, 16'd50915, 16'd35830, 16'd26426, 16'd32554, 16'd53, 16'd24567, 16'd1359, 16'd61332, 16'd53852, 16'd10521, 16'd64753, 16'd28653, 16'd19661, 16'd48845, 16'd45892, 16'd5356, 16'd22606, 16'd35126, 16'd33866});
	test_expansion(128'h0b6cdf2e028bc9419aa166017b5fe2ca, {16'd49669, 16'd45850, 16'd38960, 16'd39918, 16'd5067, 16'd43006, 16'd16450, 16'd24986, 16'd35036, 16'd32034, 16'd56380, 16'd48727, 16'd12790, 16'd52794, 16'd2597, 16'd1334, 16'd14753, 16'd34988, 16'd44661, 16'd38018, 16'd6691, 16'd45520, 16'd12, 16'd60344, 16'd10688, 16'd23252});
	test_expansion(128'hf13704b272b42498bfbf2b6c76493042, {16'd28825, 16'd29549, 16'd37712, 16'd32001, 16'd20257, 16'd16839, 16'd42458, 16'd12098, 16'd49247, 16'd43242, 16'd52898, 16'd7087, 16'd18570, 16'd33463, 16'd3912, 16'd51769, 16'd1984, 16'd14517, 16'd28528, 16'd42481, 16'd28658, 16'd43755, 16'd11642, 16'd50317, 16'd61925, 16'd22337});
	test_expansion(128'had2e95a6ecc3ea9b3f9d1fcee975dbb9, {16'd17436, 16'd63230, 16'd38722, 16'd3750, 16'd60181, 16'd22834, 16'd53263, 16'd24134, 16'd31591, 16'd36915, 16'd64757, 16'd36835, 16'd29899, 16'd42150, 16'd29977, 16'd163, 16'd44072, 16'd2932, 16'd61908, 16'd57140, 16'd13558, 16'd64821, 16'd42658, 16'd64198, 16'd34770, 16'd42086});
	test_expansion(128'h5d16c228437cd1ec67577f2164e3c964, {16'd25361, 16'd64005, 16'd43420, 16'd40544, 16'd3824, 16'd62356, 16'd38427, 16'd46999, 16'd55247, 16'd1178, 16'd52298, 16'd36226, 16'd39118, 16'd34036, 16'd46283, 16'd9741, 16'd26983, 16'd8058, 16'd44488, 16'd53682, 16'd30251, 16'd30627, 16'd17791, 16'd4143, 16'd8069, 16'd42639});
	test_expansion(128'hb2e7b5bd039e36f8a5dd59b105224147, {16'd47105, 16'd27002, 16'd59624, 16'd2522, 16'd7393, 16'd63574, 16'd20965, 16'd26087, 16'd38335, 16'd28468, 16'd19454, 16'd56852, 16'd47467, 16'd46006, 16'd23266, 16'd53199, 16'd31712, 16'd21767, 16'd8854, 16'd13674, 16'd26328, 16'd46812, 16'd24070, 16'd26379, 16'd59203, 16'd25300});
	test_expansion(128'h8bce3a94da2343574c8b566f5226163a, {16'd11897, 16'd4998, 16'd33012, 16'd6245, 16'd21393, 16'd39592, 16'd11472, 16'd25740, 16'd39904, 16'd58330, 16'd33753, 16'd52961, 16'd39387, 16'd26296, 16'd19853, 16'd6613, 16'd24656, 16'd23057, 16'd11043, 16'd14400, 16'd9255, 16'd40664, 16'd21984, 16'd4289, 16'd61911, 16'd35978});
	test_expansion(128'hb22f67c50fa4c88d99c2f733b9cf68e0, {16'd45756, 16'd44253, 16'd3906, 16'd26430, 16'd28186, 16'd57305, 16'd32988, 16'd23153, 16'd19084, 16'd33575, 16'd5481, 16'd25257, 16'd45569, 16'd41425, 16'd43345, 16'd619, 16'd2987, 16'd39342, 16'd6375, 16'd10900, 16'd43788, 16'd14166, 16'd12237, 16'd9416, 16'd31228, 16'd25949});
	test_expansion(128'he8a008d2100aad75af55837ee4f9f44f, {16'd11638, 16'd10441, 16'd29654, 16'd8045, 16'd45631, 16'd19490, 16'd44344, 16'd57567, 16'd37398, 16'd5718, 16'd39110, 16'd47154, 16'd57693, 16'd32865, 16'd9197, 16'd48012, 16'd10973, 16'd61451, 16'd8611, 16'd30812, 16'd53227, 16'd19503, 16'd26569, 16'd43116, 16'd18709, 16'd44696});
	test_expansion(128'h15acb1ab49a7f3c4e18a3b25a5b2c7fa, {16'd34630, 16'd35081, 16'd48997, 16'd31094, 16'd2039, 16'd50031, 16'd28095, 16'd64993, 16'd53304, 16'd51408, 16'd43609, 16'd19119, 16'd60854, 16'd25931, 16'd19832, 16'd42896, 16'd29553, 16'd64918, 16'd52635, 16'd17344, 16'd14424, 16'd64914, 16'd6798, 16'd43704, 16'd33616, 16'd23230});
	test_expansion(128'h76d85a1eb992ddbe679ea8bee5bb0c25, {16'd7169, 16'd58873, 16'd926, 16'd60290, 16'd58586, 16'd62866, 16'd7437, 16'd21068, 16'd29352, 16'd13697, 16'd46851, 16'd29810, 16'd28139, 16'd60047, 16'd4967, 16'd57744, 16'd56980, 16'd7849, 16'd29039, 16'd40485, 16'd1959, 16'd22981, 16'd15895, 16'd33305, 16'd29473, 16'd31733});
	test_expansion(128'h5cb2943b8a76698ccb6c4b1c2c2d9924, {16'd45087, 16'd24463, 16'd5066, 16'd28854, 16'd54342, 16'd11520, 16'd63934, 16'd7084, 16'd11036, 16'd58788, 16'd42829, 16'd44608, 16'd30267, 16'd18638, 16'd63633, 16'd17578, 16'd44751, 16'd26095, 16'd46761, 16'd249, 16'd63243, 16'd16129, 16'd40898, 16'd33844, 16'd56917, 16'd61828});
	test_expansion(128'h4645c8ba5d44b36c144ca1c7c4d7dbee, {16'd12165, 16'd44585, 16'd34498, 16'd15126, 16'd49745, 16'd53761, 16'd59379, 16'd18602, 16'd61377, 16'd45596, 16'd52913, 16'd56095, 16'd29840, 16'd19984, 16'd18420, 16'd14444, 16'd19486, 16'd6207, 16'd2030, 16'd3292, 16'd43643, 16'd38169, 16'd61493, 16'd38171, 16'd32502, 16'd38050});
	test_expansion(128'h2a10394049c17a98478227f2fde0f845, {16'd11738, 16'd60687, 16'd25468, 16'd53966, 16'd37505, 16'd34681, 16'd5485, 16'd55521, 16'd20478, 16'd24858, 16'd2246, 16'd37381, 16'd21541, 16'd29289, 16'd35549, 16'd35235, 16'd23478, 16'd10274, 16'd27005, 16'd33822, 16'd24685, 16'd6756, 16'd50581, 16'd9250, 16'd62075, 16'd37567});
	test_expansion(128'hc08c87daed4bab5492890a4176181b3a, {16'd61710, 16'd16089, 16'd16100, 16'd34050, 16'd43480, 16'd22523, 16'd17034, 16'd25384, 16'd38701, 16'd48877, 16'd20134, 16'd51190, 16'd56307, 16'd16005, 16'd34369, 16'd21633, 16'd43548, 16'd19418, 16'd45397, 16'd25420, 16'd49102, 16'd56006, 16'd35206, 16'd36166, 16'd25866, 16'd38619});
	test_expansion(128'hb8cdd9391664a591e746d7b5d81c56eb, {16'd8191, 16'd65463, 16'd64237, 16'd8237, 16'd51157, 16'd17266, 16'd51812, 16'd43226, 16'd35713, 16'd20226, 16'd48547, 16'd51366, 16'd26497, 16'd20925, 16'd45721, 16'd13323, 16'd45167, 16'd29211, 16'd30593, 16'd48770, 16'd54473, 16'd5048, 16'd41581, 16'd30562, 16'd43657, 16'd29550});
	test_expansion(128'h0c50ea71476fffb406d10da3d866bc50, {16'd24351, 16'd16421, 16'd46917, 16'd19264, 16'd60688, 16'd63333, 16'd15759, 16'd29939, 16'd50993, 16'd17569, 16'd64699, 16'd9647, 16'd34622, 16'd52096, 16'd2778, 16'd28075, 16'd48130, 16'd52611, 16'd13072, 16'd30349, 16'd8539, 16'd17222, 16'd49708, 16'd48259, 16'd6626, 16'd24679});
	test_expansion(128'h76c51508e7eef84f2e6600bcd59d5461, {16'd18429, 16'd7397, 16'd27538, 16'd42013, 16'd61741, 16'd6573, 16'd63102, 16'd47434, 16'd14360, 16'd4404, 16'd24575, 16'd26272, 16'd59976, 16'd23484, 16'd14822, 16'd11081, 16'd24522, 16'd28494, 16'd31084, 16'd56154, 16'd38938, 16'd48894, 16'd37023, 16'd42496, 16'd37887, 16'd51304});
	test_expansion(128'ha36a1ade3d61d9b25fa4f049bec9f5b4, {16'd61609, 16'd54455, 16'd53920, 16'd1126, 16'd22479, 16'd48766, 16'd12881, 16'd13498, 16'd2061, 16'd52807, 16'd25072, 16'd64252, 16'd58750, 16'd21018, 16'd18225, 16'd58031, 16'd33339, 16'd16387, 16'd40066, 16'd4497, 16'd62634, 16'd61236, 16'd33569, 16'd14229, 16'd6460, 16'd25267});
	test_expansion(128'hbd649706ef18ab35d999473b4bfaaca8, {16'd6767, 16'd25854, 16'd33429, 16'd19698, 16'd20396, 16'd16693, 16'd58046, 16'd34595, 16'd25437, 16'd9327, 16'd25369, 16'd56635, 16'd23523, 16'd50291, 16'd51034, 16'd6184, 16'd46291, 16'd29327, 16'd17432, 16'd18850, 16'd40428, 16'd2604, 16'd15558, 16'd60336, 16'd19705, 16'd46760});
	test_expansion(128'h762c9130306777da89407c04ba21864d, {16'd62121, 16'd13389, 16'd3746, 16'd62982, 16'd57915, 16'd48924, 16'd40531, 16'd27481, 16'd38825, 16'd9667, 16'd29826, 16'd2776, 16'd26394, 16'd37728, 16'd36632, 16'd25990, 16'd49635, 16'd55972, 16'd30895, 16'd5374, 16'd16245, 16'd29187, 16'd53170, 16'd16692, 16'd49811, 16'd46684});
	test_expansion(128'hd9d0b60662d5488d0c082863f6fca18b, {16'd5288, 16'd40866, 16'd30491, 16'd31589, 16'd62808, 16'd11015, 16'd55856, 16'd41012, 16'd10457, 16'd19571, 16'd53479, 16'd27249, 16'd17472, 16'd42198, 16'd54098, 16'd37492, 16'd64989, 16'd45821, 16'd12268, 16'd61104, 16'd57543, 16'd43095, 16'd57242, 16'd62129, 16'd35394, 16'd33594});
	test_expansion(128'hbba535e21a2bef179f1bee9cc2d5e247, {16'd46799, 16'd46056, 16'd38810, 16'd13893, 16'd28317, 16'd55010, 16'd25302, 16'd42552, 16'd46787, 16'd55096, 16'd1086, 16'd33020, 16'd57791, 16'd43844, 16'd62687, 16'd42775, 16'd35876, 16'd33892, 16'd29943, 16'd23634, 16'd63022, 16'd47684, 16'd4647, 16'd30025, 16'd42628, 16'd27777});
	test_expansion(128'hf3b034c809eaa46b27d9743dd007948c, {16'd26600, 16'd17238, 16'd40305, 16'd31806, 16'd63912, 16'd34686, 16'd45690, 16'd89, 16'd26074, 16'd4487, 16'd5435, 16'd63423, 16'd15004, 16'd39088, 16'd35058, 16'd60133, 16'd47030, 16'd52533, 16'd65248, 16'd3542, 16'd41900, 16'd44174, 16'd34230, 16'd63260, 16'd4779, 16'd14755});
	test_expansion(128'h3b6dc79359e6db9d9dc28933e584b8c4, {16'd50010, 16'd44118, 16'd7321, 16'd58274, 16'd50902, 16'd16754, 16'd60109, 16'd58759, 16'd64684, 16'd10354, 16'd44587, 16'd59775, 16'd63186, 16'd2926, 16'd14099, 16'd1173, 16'd23558, 16'd53369, 16'd23836, 16'd62733, 16'd38393, 16'd61814, 16'd8385, 16'd42184, 16'd59915, 16'd8783});
	test_expansion(128'h7e4e32d719e7ab6e599fea1d596393db, {16'd15381, 16'd59514, 16'd42531, 16'd32740, 16'd3477, 16'd14124, 16'd21510, 16'd3412, 16'd27818, 16'd34634, 16'd29316, 16'd55445, 16'd49181, 16'd63866, 16'd43179, 16'd60168, 16'd20331, 16'd34444, 16'd25953, 16'd51362, 16'd64052, 16'd40177, 16'd2144, 16'd367, 16'd38977, 16'd44365});
	test_expansion(128'h61a8c26dc9c7c419e6d61b4efc586608, {16'd12594, 16'd31770, 16'd38267, 16'd19217, 16'd7705, 16'd12453, 16'd45531, 16'd41853, 16'd6134, 16'd18462, 16'd31106, 16'd52000, 16'd35522, 16'd55782, 16'd1886, 16'd31455, 16'd54171, 16'd63625, 16'd7582, 16'd46470, 16'd26364, 16'd38716, 16'd64032, 16'd1033, 16'd29473, 16'd60696});
	test_expansion(128'h3796e8869a877fcb730781875d3b75b9, {16'd38691, 16'd50420, 16'd33768, 16'd39988, 16'd36871, 16'd47685, 16'd38994, 16'd29581, 16'd51607, 16'd10086, 16'd922, 16'd10670, 16'd62983, 16'd49454, 16'd43272, 16'd19953, 16'd42178, 16'd19303, 16'd38257, 16'd47530, 16'd57708, 16'd48987, 16'd52750, 16'd23290, 16'd34496, 16'd52734});
	test_expansion(128'h205b46d2be0dbce0dc3185d9d54410b3, {16'd64072, 16'd7803, 16'd41232, 16'd32423, 16'd45155, 16'd62101, 16'd61315, 16'd45160, 16'd16631, 16'd45682, 16'd7147, 16'd58152, 16'd13632, 16'd57485, 16'd39746, 16'd43804, 16'd29198, 16'd21552, 16'd12916, 16'd48409, 16'd62388, 16'd47039, 16'd21231, 16'd51543, 16'd59710, 16'd45196});
	test_expansion(128'h82b1b1c392793e306edcbb75358acb20, {16'd49980, 16'd11969, 16'd56498, 16'd60873, 16'd31777, 16'd47835, 16'd58055, 16'd18501, 16'd4434, 16'd26024, 16'd37661, 16'd18747, 16'd37532, 16'd26136, 16'd14547, 16'd11593, 16'd30515, 16'd57982, 16'd61239, 16'd39938, 16'd45192, 16'd15939, 16'd50021, 16'd43416, 16'd35895, 16'd14713});
	test_expansion(128'h1da9fec6d9ecf6e603f824f40a682d03, {16'd32041, 16'd50864, 16'd61873, 16'd25200, 16'd22799, 16'd18583, 16'd44364, 16'd19109, 16'd38416, 16'd31826, 16'd32912, 16'd8490, 16'd35870, 16'd60342, 16'd33311, 16'd37315, 16'd55981, 16'd31444, 16'd38600, 16'd63639, 16'd59595, 16'd16674, 16'd41644, 16'd44364, 16'd43849, 16'd47319});
	test_expansion(128'ha2c8665fb762eaf9ee11f62864ea4384, {16'd58377, 16'd13695, 16'd33827, 16'd372, 16'd23495, 16'd41595, 16'd48923, 16'd43133, 16'd5819, 16'd55233, 16'd2064, 16'd28764, 16'd64781, 16'd35621, 16'd13268, 16'd15362, 16'd57088, 16'd48654, 16'd62437, 16'd43302, 16'd23507, 16'd17660, 16'd7047, 16'd3291, 16'd4617, 16'd16308});
	test_expansion(128'h59b8f0144b59050573bf8a040b83fd94, {16'd5104, 16'd1783, 16'd56760, 16'd24548, 16'd47522, 16'd32287, 16'd9829, 16'd32572, 16'd41459, 16'd10411, 16'd50522, 16'd46969, 16'd30130, 16'd2661, 16'd64118, 16'd31038, 16'd16766, 16'd28871, 16'd39370, 16'd57947, 16'd1978, 16'd50695, 16'd44470, 16'd14856, 16'd43391, 16'd14626});
	test_expansion(128'h3c4e0a04dcc42483a05d936a3908f4f6, {16'd583, 16'd49794, 16'd33115, 16'd29631, 16'd38677, 16'd19581, 16'd10936, 16'd60795, 16'd29935, 16'd54602, 16'd15463, 16'd42383, 16'd60457, 16'd39484, 16'd37413, 16'd41007, 16'd19891, 16'd49486, 16'd33045, 16'd31023, 16'd8628, 16'd35368, 16'd22217, 16'd58197, 16'd44950, 16'd54454});
	test_expansion(128'h3bb2bba63373151fae03c1ee732adf6e, {16'd18376, 16'd49281, 16'd26807, 16'd46740, 16'd38397, 16'd49079, 16'd3632, 16'd25921, 16'd23270, 16'd29286, 16'd33384, 16'd23072, 16'd33133, 16'd46570, 16'd12334, 16'd18949, 16'd64156, 16'd41321, 16'd46550, 16'd26175, 16'd44919, 16'd19566, 16'd54722, 16'd60813, 16'd8093, 16'd40627});
	test_expansion(128'h77a8c64c54b221ed1d752998fdd28a84, {16'd20089, 16'd10622, 16'd23374, 16'd9401, 16'd48785, 16'd17693, 16'd55303, 16'd30574, 16'd6218, 16'd10547, 16'd45529, 16'd52156, 16'd7867, 16'd38652, 16'd18665, 16'd42477, 16'd12611, 16'd54779, 16'd60946, 16'd5817, 16'd17280, 16'd31839, 16'd10800, 16'd26432, 16'd9638, 16'd16641});
	test_expansion(128'h998366a96bfa54fb1a58b9fd06ad9be8, {16'd34218, 16'd54750, 16'd34738, 16'd16544, 16'd40101, 16'd39693, 16'd1108, 16'd27242, 16'd20008, 16'd41323, 16'd43758, 16'd42294, 16'd64685, 16'd55422, 16'd54385, 16'd42663, 16'd36160, 16'd34714, 16'd62353, 16'd31190, 16'd65435, 16'd49963, 16'd58613, 16'd25688, 16'd20452, 16'd57433});
	test_expansion(128'ha2b7b1bb1377329073519099fda17129, {16'd11886, 16'd26781, 16'd41704, 16'd48026, 16'd45867, 16'd61932, 16'd65387, 16'd64663, 16'd57462, 16'd29701, 16'd53859, 16'd57459, 16'd51526, 16'd5566, 16'd20117, 16'd50223, 16'd30479, 16'd59793, 16'd49687, 16'd37932, 16'd28846, 16'd58149, 16'd33639, 16'd2650, 16'd35110, 16'd38715});
	test_expansion(128'h9383b44cc2bf6613c1aa617475ceb8a1, {16'd10656, 16'd19105, 16'd61398, 16'd12653, 16'd44035, 16'd46031, 16'd2602, 16'd16377, 16'd20583, 16'd21922, 16'd34895, 16'd24186, 16'd48846, 16'd15140, 16'd10531, 16'd9216, 16'd9686, 16'd4975, 16'd47485, 16'd50361, 16'd11308, 16'd33189, 16'd64559, 16'd30335, 16'd59885, 16'd3602});
	test_expansion(128'hba92fe3017d12f7e21c9c263df8a5f86, {16'd10393, 16'd11052, 16'd16496, 16'd59382, 16'd62519, 16'd58404, 16'd21528, 16'd46228, 16'd39721, 16'd50040, 16'd32114, 16'd3273, 16'd26509, 16'd37367, 16'd33477, 16'd27820, 16'd26802, 16'd7858, 16'd52375, 16'd60944, 16'd30540, 16'd3830, 16'd11607, 16'd25308, 16'd13819, 16'd32644});
	test_expansion(128'h9a3ef4d86a99902d397f276bd53c21c0, {16'd58981, 16'd27884, 16'd47044, 16'd6699, 16'd51054, 16'd33200, 16'd49924, 16'd37537, 16'd14936, 16'd17096, 16'd35200, 16'd48882, 16'd55613, 16'd62559, 16'd38025, 16'd6351, 16'd36287, 16'd31882, 16'd26760, 16'd51817, 16'd3642, 16'd35660, 16'd43240, 16'd12987, 16'd61962, 16'd61560});
	test_expansion(128'h02d7e2f1f797aa8afa7410ec476ae4a0, {16'd54953, 16'd48822, 16'd42725, 16'd54849, 16'd7301, 16'd25558, 16'd53432, 16'd19482, 16'd59401, 16'd63734, 16'd51496, 16'd33986, 16'd9684, 16'd22265, 16'd38020, 16'd35253, 16'd53623, 16'd58691, 16'd52885, 16'd46955, 16'd22074, 16'd25026, 16'd37255, 16'd19426, 16'd63790, 16'd15772});
	test_expansion(128'hb23b8a509a189a2dbf4477ec49987149, {16'd22259, 16'd4538, 16'd62005, 16'd20549, 16'd45916, 16'd15030, 16'd32490, 16'd62997, 16'd47904, 16'd35649, 16'd60003, 16'd24670, 16'd13931, 16'd12945, 16'd14666, 16'd17625, 16'd62695, 16'd14479, 16'd23192, 16'd56496, 16'd12525, 16'd38766, 16'd57674, 16'd63582, 16'd15898, 16'd7415});
	test_expansion(128'ha2c4bd12564ba14ee4ef639339e3c394, {16'd46123, 16'd6407, 16'd59135, 16'd12260, 16'd57681, 16'd61094, 16'd33617, 16'd841, 16'd63190, 16'd49041, 16'd22944, 16'd56644, 16'd45195, 16'd7886, 16'd29232, 16'd8972, 16'd21311, 16'd40784, 16'd6419, 16'd11940, 16'd43727, 16'd48686, 16'd55426, 16'd56900, 16'd3399, 16'd56805});
	test_expansion(128'hca137f1cbc086508460898bc030e5976, {16'd50900, 16'd12596, 16'd28252, 16'd16344, 16'd61598, 16'd31584, 16'd7080, 16'd13400, 16'd61248, 16'd50544, 16'd21095, 16'd55004, 16'd23383, 16'd65198, 16'd46403, 16'd44715, 16'd58745, 16'd8123, 16'd54601, 16'd2713, 16'd10685, 16'd61202, 16'd65150, 16'd49718, 16'd44472, 16'd34584});
	test_expansion(128'h3580cbac2f5d0f7f404756505193407c, {16'd48450, 16'd62430, 16'd17540, 16'd26253, 16'd57919, 16'd23311, 16'd40475, 16'd7580, 16'd30856, 16'd64065, 16'd56434, 16'd40772, 16'd14456, 16'd50455, 16'd42748, 16'd15671, 16'd40226, 16'd29802, 16'd48567, 16'd20564, 16'd282, 16'd41785, 16'd12565, 16'd50099, 16'd14038, 16'd14697});
	test_expansion(128'h56fe867ad33f87a8259a152c6da796a6, {16'd37426, 16'd46336, 16'd47194, 16'd27062, 16'd35425, 16'd1379, 16'd56207, 16'd48909, 16'd20414, 16'd59586, 16'd12977, 16'd40585, 16'd54148, 16'd49294, 16'd45574, 16'd51602, 16'd57080, 16'd53245, 16'd32242, 16'd38878, 16'd40349, 16'd50405, 16'd56601, 16'd36760, 16'd2292, 16'd16436});
	test_expansion(128'h4d30d22d41695f299b677186866ac2e6, {16'd17408, 16'd25751, 16'd47993, 16'd55660, 16'd18300, 16'd28053, 16'd3517, 16'd3216, 16'd33625, 16'd57493, 16'd41197, 16'd31305, 16'd51781, 16'd9929, 16'd43951, 16'd51197, 16'd44056, 16'd8115, 16'd56578, 16'd21851, 16'd42732, 16'd30028, 16'd42268, 16'd7709, 16'd53335, 16'd23253});
	test_expansion(128'ha4db648e1b62573a3962bb997910a768, {16'd43078, 16'd620, 16'd4090, 16'd35149, 16'd55288, 16'd17988, 16'd37151, 16'd17716, 16'd7863, 16'd63017, 16'd65214, 16'd49670, 16'd13024, 16'd3768, 16'd52022, 16'd5682, 16'd37480, 16'd59009, 16'd6476, 16'd28529, 16'd6183, 16'd60751, 16'd9339, 16'd61236, 16'd20708, 16'd47445});
	test_expansion(128'hb4ec8d7825849a140c67bbb67fbcaf1c, {16'd3005, 16'd49010, 16'd60715, 16'd37610, 16'd12699, 16'd53078, 16'd55247, 16'd29500, 16'd3609, 16'd55356, 16'd12736, 16'd62878, 16'd60088, 16'd53728, 16'd1267, 16'd2114, 16'd53391, 16'd52037, 16'd33162, 16'd2042, 16'd5395, 16'd1569, 16'd39254, 16'd32283, 16'd41957, 16'd55602});
	test_expansion(128'h79c1a25afecedc677fdb1f0c359add77, {16'd5846, 16'd1068, 16'd17875, 16'd20107, 16'd51684, 16'd36702, 16'd43454, 16'd43534, 16'd22923, 16'd1532, 16'd56625, 16'd56688, 16'd10889, 16'd64616, 16'd52719, 16'd7242, 16'd16177, 16'd20633, 16'd48385, 16'd50220, 16'd58641, 16'd11424, 16'd45042, 16'd27934, 16'd26999, 16'd3548});
	test_expansion(128'hf0621c9faabd4ac73ec2c2cb4b2445b5, {16'd32293, 16'd384, 16'd61765, 16'd36027, 16'd13812, 16'd10820, 16'd61689, 16'd46381, 16'd40749, 16'd63834, 16'd14298, 16'd4584, 16'd64260, 16'd36476, 16'd30315, 16'd22622, 16'd64285, 16'd18012, 16'd18574, 16'd43683, 16'd5367, 16'd53631, 16'd62265, 16'd53198, 16'd41867, 16'd35837});
	test_expansion(128'h8ebb1c7a7a71ef99a235b7f635d6209b, {16'd13159, 16'd36551, 16'd39145, 16'd27708, 16'd12265, 16'd36237, 16'd36140, 16'd22583, 16'd43472, 16'd47116, 16'd8940, 16'd24054, 16'd14354, 16'd30654, 16'd6394, 16'd65439, 16'd20087, 16'd14023, 16'd47783, 16'd16413, 16'd36873, 16'd47117, 16'd21630, 16'd1160, 16'd52229, 16'd11594});
	test_expansion(128'h27f7668724b2a116e2fb510b8a8fa80f, {16'd15090, 16'd38123, 16'd52896, 16'd56109, 16'd24171, 16'd25981, 16'd45553, 16'd34464, 16'd44434, 16'd4148, 16'd6269, 16'd35427, 16'd38071, 16'd15894, 16'd58965, 16'd19789, 16'd51835, 16'd61575, 16'd39076, 16'd45943, 16'd30488, 16'd36613, 16'd35020, 16'd56749, 16'd1779, 16'd63887});
	test_expansion(128'hd3276ea0505570b53f57c2600da529f6, {16'd13445, 16'd24210, 16'd36830, 16'd47631, 16'd19499, 16'd15355, 16'd39599, 16'd8618, 16'd42413, 16'd5466, 16'd1544, 16'd1159, 16'd25328, 16'd31688, 16'd23306, 16'd397, 16'd63135, 16'd48442, 16'd40909, 16'd48722, 16'd159, 16'd2800, 16'd52647, 16'd50295, 16'd12949, 16'd42790});
	test_expansion(128'hd9ffd2eac3cbd68e80046112d343ef6d, {16'd36793, 16'd54896, 16'd38228, 16'd28953, 16'd5583, 16'd27283, 16'd43245, 16'd8029, 16'd3655, 16'd8791, 16'd40655, 16'd43225, 16'd35949, 16'd12118, 16'd1916, 16'd39725, 16'd57661, 16'd21697, 16'd34619, 16'd40889, 16'd46748, 16'd53499, 16'd18719, 16'd33019, 16'd54598, 16'd32255});
	test_expansion(128'h09d2b1a8915b7d4296e5a0574e0ee2d0, {16'd44505, 16'd23019, 16'd16998, 16'd14269, 16'd46866, 16'd34119, 16'd19877, 16'd44405, 16'd34116, 16'd54959, 16'd43622, 16'd12680, 16'd21201, 16'd16775, 16'd55681, 16'd39993, 16'd54079, 16'd62825, 16'd5690, 16'd63920, 16'd47382, 16'd36703, 16'd34082, 16'd27663, 16'd21687, 16'd8652});
	test_expansion(128'hfa78c37db6b7791afe288140dcac8f40, {16'd3597, 16'd42602, 16'd32030, 16'd35074, 16'd63970, 16'd29111, 16'd56177, 16'd59465, 16'd3193, 16'd45514, 16'd5522, 16'd18334, 16'd8802, 16'd64778, 16'd45155, 16'd30222, 16'd1208, 16'd10517, 16'd18091, 16'd8889, 16'd5173, 16'd34687, 16'd44170, 16'd41777, 16'd24782, 16'd13012});
	test_expansion(128'ha4e3e0a315d57543e943ac2101cdb896, {16'd7690, 16'd15745, 16'd34748, 16'd11802, 16'd35747, 16'd56293, 16'd55872, 16'd35201, 16'd26194, 16'd12008, 16'd5324, 16'd17190, 16'd9681, 16'd41592, 16'd24816, 16'd54077, 16'd28840, 16'd33376, 16'd47931, 16'd13792, 16'd37345, 16'd45728, 16'd2743, 16'd53505, 16'd25381, 16'd43246});
	test_expansion(128'hc1312f7b47032f11b73de931f894ce85, {16'd64341, 16'd56510, 16'd64341, 16'd20918, 16'd45431, 16'd50028, 16'd38211, 16'd10450, 16'd22242, 16'd19650, 16'd63848, 16'd35534, 16'd18882, 16'd11022, 16'd25271, 16'd24492, 16'd45969, 16'd53253, 16'd62900, 16'd40842, 16'd16980, 16'd12132, 16'd48708, 16'd21394, 16'd38988, 16'd56267});
	test_expansion(128'he98220d075eafad0e59170f87db592d6, {16'd17127, 16'd62643, 16'd53584, 16'd37385, 16'd9573, 16'd43957, 16'd59310, 16'd31737, 16'd37197, 16'd32999, 16'd24025, 16'd28743, 16'd64166, 16'd33262, 16'd53772, 16'd5573, 16'd463, 16'd33917, 16'd52378, 16'd15444, 16'd25570, 16'd41924, 16'd62643, 16'd19025, 16'd19585, 16'd31725});
	test_expansion(128'ha88cd32c15242fc837851f1fbf0e3d36, {16'd44275, 16'd34537, 16'd34894, 16'd44269, 16'd54032, 16'd46886, 16'd46568, 16'd64489, 16'd59675, 16'd64152, 16'd7875, 16'd38434, 16'd4660, 16'd40411, 16'd50513, 16'd40820, 16'd37108, 16'd64895, 16'd19765, 16'd23193, 16'd43293, 16'd4074, 16'd8340, 16'd59250, 16'd31713, 16'd15590});
	test_expansion(128'h56a2834d19b6504ba86b0c8f9b03ddde, {16'd58318, 16'd10450, 16'd40945, 16'd41157, 16'd45664, 16'd8444, 16'd37593, 16'd19786, 16'd30356, 16'd24108, 16'd8135, 16'd43697, 16'd20551, 16'd37365, 16'd61309, 16'd11029, 16'd26060, 16'd11871, 16'd15859, 16'd55591, 16'd9696, 16'd8368, 16'd20274, 16'd35176, 16'd36538, 16'd9291});
	test_expansion(128'hd111e0d0faff228d6b9251ee640be90b, {16'd38334, 16'd36397, 16'd16911, 16'd14510, 16'd62010, 16'd17093, 16'd59327, 16'd44524, 16'd26857, 16'd8774, 16'd471, 16'd47464, 16'd23895, 16'd45658, 16'd55387, 16'd65052, 16'd62608, 16'd47267, 16'd54740, 16'd41757, 16'd48945, 16'd18804, 16'd21237, 16'd3844, 16'd14847, 16'd41304});
	test_expansion(128'hc7de93d7c254a0de0968248532bc3584, {16'd15773, 16'd45639, 16'd44933, 16'd18406, 16'd40522, 16'd36120, 16'd45233, 16'd27315, 16'd35575, 16'd27591, 16'd50483, 16'd44255, 16'd55024, 16'd46740, 16'd40089, 16'd10423, 16'd15466, 16'd60346, 16'd52578, 16'd40711, 16'd6661, 16'd41360, 16'd10366, 16'd29724, 16'd53706, 16'd28313});
	test_expansion(128'hf8f26f84b2e9f8f1cabc845b3a077291, {16'd30448, 16'd36262, 16'd38503, 16'd51101, 16'd46953, 16'd20816, 16'd45948, 16'd46904, 16'd9, 16'd17176, 16'd22937, 16'd63226, 16'd23106, 16'd34455, 16'd26528, 16'd12898, 16'd14487, 16'd48934, 16'd8770, 16'd49591, 16'd32632, 16'd54110, 16'd41798, 16'd8577, 16'd24728, 16'd62290});
	test_expansion(128'ha24737b73951d001e14f53c262742440, {16'd1463, 16'd57878, 16'd20995, 16'd31273, 16'd47885, 16'd8963, 16'd16250, 16'd65020, 16'd8865, 16'd13481, 16'd54417, 16'd14517, 16'd16583, 16'd47789, 16'd12871, 16'd1673, 16'd5151, 16'd26234, 16'd10453, 16'd63155, 16'd62682, 16'd20834, 16'd10289, 16'd16092, 16'd43391, 16'd50653});
	test_expansion(128'h5fdde7d5fcf2a80ec0f855c8dd110f07, {16'd43324, 16'd46640, 16'd44891, 16'd43803, 16'd21648, 16'd5995, 16'd16449, 16'd8905, 16'd8337, 16'd38919, 16'd1136, 16'd21332, 16'd56709, 16'd46087, 16'd40617, 16'd51330, 16'd43212, 16'd53831, 16'd35115, 16'd60683, 16'd53653, 16'd15170, 16'd30024, 16'd379, 16'd54221, 16'd814});
	test_expansion(128'hb0fc6ef0024218da37b87ecbb0fd5a09, {16'd63349, 16'd43433, 16'd13460, 16'd3536, 16'd51260, 16'd6191, 16'd53276, 16'd64735, 16'd15482, 16'd42322, 16'd58124, 16'd65258, 16'd12918, 16'd35918, 16'd22338, 16'd8961, 16'd55755, 16'd38988, 16'd16599, 16'd61323, 16'd42336, 16'd41108, 16'd29265, 16'd23043, 16'd40925, 16'd59355});
	test_expansion(128'h71c058302d66ef2ad24fc3569ab70020, {16'd6624, 16'd14709, 16'd39861, 16'd31509, 16'd29378, 16'd33646, 16'd59854, 16'd32428, 16'd57684, 16'd36919, 16'd48269, 16'd30345, 16'd31726, 16'd29943, 16'd51785, 16'd35260, 16'd28905, 16'd20522, 16'd48183, 16'd61719, 16'd36317, 16'd46512, 16'd50724, 16'd152, 16'd30532, 16'd41871});
	test_expansion(128'hbdf7d83e8c9165b01350abe726f6dee2, {16'd19722, 16'd49179, 16'd18537, 16'd33729, 16'd16396, 16'd64732, 16'd16011, 16'd46740, 16'd33358, 16'd6676, 16'd25493, 16'd56062, 16'd7284, 16'd53885, 16'd54548, 16'd16298, 16'd47257, 16'd39048, 16'd6741, 16'd59130, 16'd2054, 16'd9480, 16'd41380, 16'd59982, 16'd60469, 16'd51969});
	test_expansion(128'h33e811a1df389d08e3049698b08f3786, {16'd64540, 16'd921, 16'd61687, 16'd21193, 16'd32457, 16'd30160, 16'd35353, 16'd10811, 16'd15231, 16'd33866, 16'd12807, 16'd11065, 16'd23643, 16'd2331, 16'd42236, 16'd909, 16'd43917, 16'd60199, 16'd31366, 16'd19225, 16'd11316, 16'd60961, 16'd60803, 16'd13496, 16'd44434, 16'd12618});
	test_expansion(128'h554e39038468e8d5f4a32b675fe6d7d5, {16'd5516, 16'd50245, 16'd45307, 16'd52773, 16'd10692, 16'd55274, 16'd19184, 16'd52834, 16'd49156, 16'd27340, 16'd62870, 16'd31208, 16'd61161, 16'd52244, 16'd38512, 16'd21016, 16'd7100, 16'd5618, 16'd51631, 16'd40, 16'd38007, 16'd6540, 16'd57854, 16'd32533, 16'd15472, 16'd11958});
	test_expansion(128'he8ac4c65b3759dd3cdf0974a1004ea34, {16'd25771, 16'd12361, 16'd20232, 16'd33259, 16'd12876, 16'd63225, 16'd45781, 16'd45419, 16'd6401, 16'd54035, 16'd10536, 16'd15479, 16'd65012, 16'd37682, 16'd42942, 16'd38225, 16'd27457, 16'd54116, 16'd47628, 16'd60335, 16'd15401, 16'd51669, 16'd61958, 16'd53903, 16'd50866, 16'd26505});
	test_expansion(128'hdf3462515853e4de7c5d403e541f7566, {16'd39319, 16'd25852, 16'd12815, 16'd29797, 16'd28054, 16'd8340, 16'd38234, 16'd30087, 16'd40066, 16'd26972, 16'd23916, 16'd39149, 16'd27109, 16'd39933, 16'd16306, 16'd34379, 16'd21365, 16'd33048, 16'd41262, 16'd24944, 16'd53347, 16'd62745, 16'd1674, 16'd29097, 16'd637, 16'd25994});
	test_expansion(128'h798aa68e48b2923419e3a6b0c5b594b3, {16'd19139, 16'd10315, 16'd31343, 16'd27574, 16'd32721, 16'd10929, 16'd37133, 16'd24623, 16'd46857, 16'd36744, 16'd64203, 16'd47161, 16'd64250, 16'd26663, 16'd42385, 16'd48316, 16'd35562, 16'd33507, 16'd43843, 16'd26899, 16'd62633, 16'd38961, 16'd5595, 16'd54950, 16'd36045, 16'd60078});
	test_expansion(128'hcb471c012d67de33bc5bcbf43c23dbbd, {16'd39314, 16'd49507, 16'd14295, 16'd42179, 16'd43757, 16'd43745, 16'd21898, 16'd51117, 16'd62940, 16'd44225, 16'd19270, 16'd42480, 16'd36818, 16'd49853, 16'd58624, 16'd59039, 16'd59995, 16'd42704, 16'd45740, 16'd9293, 16'd7542, 16'd5834, 16'd34853, 16'd37426, 16'd4045, 16'd8172});
	test_expansion(128'h6fb725c971377aa77170d1211ac0976b, {16'd17735, 16'd2638, 16'd971, 16'd37526, 16'd40615, 16'd28617, 16'd18517, 16'd22883, 16'd47413, 16'd34711, 16'd2286, 16'd59502, 16'd30691, 16'd47217, 16'd28367, 16'd16528, 16'd37963, 16'd38734, 16'd13830, 16'd7115, 16'd40935, 16'd30920, 16'd59046, 16'd26583, 16'd13035, 16'd53719});
	test_expansion(128'he69dd6c29ef12b28b365a7d265c69074, {16'd38629, 16'd35498, 16'd13863, 16'd7629, 16'd54478, 16'd25493, 16'd28905, 16'd16416, 16'd9209, 16'd65149, 16'd61813, 16'd54830, 16'd16864, 16'd39306, 16'd52325, 16'd30873, 16'd10923, 16'd57123, 16'd60314, 16'd31101, 16'd17186, 16'd53248, 16'd56202, 16'd40268, 16'd23264, 16'd7281});
	test_expansion(128'hd740636e1f8ad31cb805c066f4a1d27f, {16'd27609, 16'd25537, 16'd52826, 16'd30889, 16'd48938, 16'd11906, 16'd46530, 16'd52341, 16'd52897, 16'd23096, 16'd28477, 16'd14267, 16'd39624, 16'd25612, 16'd55192, 16'd12111, 16'd12862, 16'd55569, 16'd10228, 16'd54722, 16'd11899, 16'd40615, 16'd17649, 16'd16656, 16'd29454, 16'd19147});
	test_expansion(128'ha4b157973df18a93b5d408850219e28e, {16'd35578, 16'd40540, 16'd25850, 16'd45687, 16'd27789, 16'd50424, 16'd45185, 16'd5858, 16'd2223, 16'd33229, 16'd11254, 16'd5891, 16'd3645, 16'd56681, 16'd55000, 16'd34014, 16'd20431, 16'd26544, 16'd31407, 16'd4474, 16'd59475, 16'd3501, 16'd25809, 16'd23603, 16'd39273, 16'd43317});
	test_expansion(128'h1d00a6725bd40ef1b53b5698fa336573, {16'd40971, 16'd18236, 16'd4827, 16'd22294, 16'd32000, 16'd37417, 16'd26694, 16'd19765, 16'd16191, 16'd33054, 16'd28872, 16'd31937, 16'd47076, 16'd38358, 16'd44227, 16'd9662, 16'd9985, 16'd43942, 16'd55201, 16'd32985, 16'd56260, 16'd16015, 16'd1084, 16'd55459, 16'd8939, 16'd45118});
	test_expansion(128'h3459a64aee7454cea8f8e239d1b50e90, {16'd1277, 16'd11835, 16'd56278, 16'd65179, 16'd63638, 16'd30210, 16'd29910, 16'd39003, 16'd57067, 16'd63382, 16'd7202, 16'd45076, 16'd57057, 16'd6690, 16'd14791, 16'd38811, 16'd31791, 16'd26403, 16'd61779, 16'd53988, 16'd14589, 16'd25098, 16'd11413, 16'd15426, 16'd3047, 16'd65445});
	test_expansion(128'hc3494d6a0464843ab1991c343ef8e6ff, {16'd39320, 16'd7839, 16'd50202, 16'd45382, 16'd8804, 16'd50800, 16'd46057, 16'd47946, 16'd50189, 16'd12176, 16'd60987, 16'd17415, 16'd40662, 16'd57657, 16'd54268, 16'd46808, 16'd31941, 16'd39159, 16'd23255, 16'd47993, 16'd22605, 16'd40386, 16'd37597, 16'd24609, 16'd62721, 16'd30067});
	test_expansion(128'h64981f213b29ba8bc950ecae6599d242, {16'd44685, 16'd21001, 16'd8980, 16'd14384, 16'd49566, 16'd62776, 16'd34757, 16'd6314, 16'd35077, 16'd62331, 16'd46840, 16'd50457, 16'd20098, 16'd10967, 16'd42121, 16'd25323, 16'd9681, 16'd27541, 16'd65408, 16'd51618, 16'd44295, 16'd53290, 16'd21943, 16'd28141, 16'd59099, 16'd50393});
	test_expansion(128'h050a0454b5d091f44dc5615465c01e78, {16'd24097, 16'd41518, 16'd1370, 16'd4572, 16'd49178, 16'd47343, 16'd35118, 16'd573, 16'd58446, 16'd10576, 16'd24381, 16'd41317, 16'd56118, 16'd37932, 16'd4256, 16'd65274, 16'd4222, 16'd29939, 16'd60930, 16'd8048, 16'd23990, 16'd3442, 16'd23056, 16'd13012, 16'd8050, 16'd8103});
	test_expansion(128'hd68229b7ee6e555ceb31f667acb26f7b, {16'd58002, 16'd20300, 16'd60571, 16'd9897, 16'd33468, 16'd12411, 16'd38338, 16'd5273, 16'd52828, 16'd63244, 16'd33679, 16'd42424, 16'd62740, 16'd48009, 16'd26513, 16'd17620, 16'd53530, 16'd33438, 16'd21275, 16'd62028, 16'd49106, 16'd32489, 16'd43761, 16'd47013, 16'd12477, 16'd39125});
	test_expansion(128'h3964a0a1f30a035e3ecbccc66a17fb84, {16'd14142, 16'd44964, 16'd21691, 16'd28890, 16'd4150, 16'd53646, 16'd39792, 16'd30816, 16'd4041, 16'd65401, 16'd142, 16'd14104, 16'd38231, 16'd33111, 16'd24242, 16'd43646, 16'd1557, 16'd2154, 16'd5152, 16'd21439, 16'd39141, 16'd1919, 16'd38546, 16'd12221, 16'd44335, 16'd36719});
	test_expansion(128'h2ec626269c6b29f69d2f7900817eaf99, {16'd58429, 16'd27446, 16'd38062, 16'd49726, 16'd20137, 16'd28589, 16'd28214, 16'd21242, 16'd2311, 16'd21790, 16'd10405, 16'd40088, 16'd63409, 16'd61051, 16'd40081, 16'd44393, 16'd4270, 16'd55973, 16'd28872, 16'd54148, 16'd13473, 16'd17344, 16'd57540, 16'd54313, 16'd6352, 16'd11406});
	test_expansion(128'heaa4f4cac14b680cec321ed97f56f615, {16'd41592, 16'd38223, 16'd34339, 16'd2176, 16'd56877, 16'd20219, 16'd13923, 16'd58045, 16'd64245, 16'd56875, 16'd24272, 16'd57477, 16'd48846, 16'd42050, 16'd12253, 16'd41908, 16'd50288, 16'd18546, 16'd65238, 16'd18039, 16'd6370, 16'd64939, 16'd40409, 16'd53847, 16'd22055, 16'd23208});
	test_expansion(128'hf52ca823dbc5f2a890614aa944859310, {16'd37621, 16'd37013, 16'd1207, 16'd28933, 16'd4677, 16'd38032, 16'd14502, 16'd34287, 16'd10695, 16'd42685, 16'd50404, 16'd59555, 16'd53031, 16'd27871, 16'd29849, 16'd63271, 16'd41135, 16'd23291, 16'd18750, 16'd45739, 16'd19177, 16'd2128, 16'd56422, 16'd43156, 16'd38424, 16'd37535});
	test_expansion(128'h42668aeb73178791ba25e1f6727c5a23, {16'd26007, 16'd38099, 16'd41144, 16'd8660, 16'd45197, 16'd7316, 16'd35713, 16'd42391, 16'd29431, 16'd13027, 16'd59848, 16'd3035, 16'd54723, 16'd56671, 16'd33220, 16'd34039, 16'd14952, 16'd17378, 16'd10299, 16'd26597, 16'd33613, 16'd24229, 16'd1145, 16'd32227, 16'd39275, 16'd1119});
	test_expansion(128'hdcc818627ebc6f6d7fe1abb669744e02, {16'd3308, 16'd14963, 16'd53080, 16'd13317, 16'd39889, 16'd10250, 16'd24114, 16'd5228, 16'd7793, 16'd55542, 16'd52393, 16'd17520, 16'd7770, 16'd58707, 16'd20004, 16'd7046, 16'd3885, 16'd5708, 16'd12660, 16'd17551, 16'd54188, 16'd58832, 16'd35260, 16'd21604, 16'd56320, 16'd50338});
	test_expansion(128'h02679573abcbd3c9ed5f8cb666c526b6, {16'd8892, 16'd57155, 16'd60428, 16'd184, 16'd1961, 16'd26435, 16'd61810, 16'd12120, 16'd5383, 16'd52290, 16'd2734, 16'd37490, 16'd19791, 16'd18246, 16'd55813, 16'd41827, 16'd22698, 16'd7067, 16'd57468, 16'd53013, 16'd22972, 16'd51968, 16'd58404, 16'd15053, 16'd42702, 16'd61185});
	test_expansion(128'hd8fe063e34a18057a72342fce118025b, {16'd3921, 16'd44751, 16'd21188, 16'd6259, 16'd17584, 16'd2876, 16'd31612, 16'd33354, 16'd12971, 16'd40152, 16'd11625, 16'd60814, 16'd5857, 16'd28294, 16'd33299, 16'd64847, 16'd62383, 16'd56438, 16'd18669, 16'd44362, 16'd47242, 16'd56423, 16'd7830, 16'd24720, 16'd55207, 16'd53793});
	test_expansion(128'h7688743375dea06a2d199ae83a7490d3, {16'd53648, 16'd46831, 16'd38119, 16'd35034, 16'd22725, 16'd52964, 16'd20789, 16'd62178, 16'd9344, 16'd65427, 16'd42881, 16'd51617, 16'd7226, 16'd8567, 16'd54393, 16'd10389, 16'd3494, 16'd48322, 16'd32302, 16'd39206, 16'd9216, 16'd3232, 16'd46791, 16'd45732, 16'd52935, 16'd4343});
	test_expansion(128'h53eb559df9d0f3be48b3de43cc6d1983, {16'd30182, 16'd2649, 16'd13813, 16'd62693, 16'd25485, 16'd12215, 16'd2513, 16'd46497, 16'd49305, 16'd61161, 16'd58125, 16'd44768, 16'd21806, 16'd64693, 16'd58618, 16'd42851, 16'd326, 16'd45595, 16'd52218, 16'd27030, 16'd3401, 16'd48828, 16'd8182, 16'd15540, 16'd39943, 16'd17680});
	test_expansion(128'h5cec329010e4815f98fda22a3f4f4756, {16'd18303, 16'd63064, 16'd31470, 16'd38702, 16'd56939, 16'd686, 16'd25314, 16'd18018, 16'd7407, 16'd61316, 16'd7174, 16'd19004, 16'd17503, 16'd14496, 16'd30852, 16'd16553, 16'd37414, 16'd43149, 16'd4951, 16'd63741, 16'd57383, 16'd35910, 16'd28051, 16'd51876, 16'd30435, 16'd10474});
	test_expansion(128'h066f5858c791718dc7d3eebbf0ff7a56, {16'd20910, 16'd36013, 16'd56771, 16'd25279, 16'd40677, 16'd32667, 16'd421, 16'd55864, 16'd15728, 16'd44021, 16'd32356, 16'd28520, 16'd45499, 16'd46491, 16'd9340, 16'd32779, 16'd50602, 16'd46306, 16'd19391, 16'd55639, 16'd57058, 16'd20617, 16'd30703, 16'd41043, 16'd19471, 16'd5754});
	test_expansion(128'h2e2e1917b65727e61c22dd66fd3f89a2, {16'd64846, 16'd65452, 16'd62818, 16'd50481, 16'd55515, 16'd3067, 16'd31088, 16'd31912, 16'd64741, 16'd21953, 16'd10418, 16'd37238, 16'd39508, 16'd33324, 16'd18438, 16'd56099, 16'd40181, 16'd63298, 16'd29828, 16'd34422, 16'd41645, 16'd50670, 16'd61759, 16'd34995, 16'd35317, 16'd64534});
	test_expansion(128'h607c177995028aa2c109c11ff690ac04, {16'd22483, 16'd22867, 16'd64092, 16'd34323, 16'd30045, 16'd7415, 16'd53760, 16'd7531, 16'd1931, 16'd40655, 16'd8207, 16'd30685, 16'd38467, 16'd14513, 16'd34193, 16'd2279, 16'd61283, 16'd23740, 16'd83, 16'd13696, 16'd52983, 16'd14769, 16'd59684, 16'd6181, 16'd15529, 16'd5146});
	test_expansion(128'h013d3457e858ee6c131105cf67072ef0, {16'd56409, 16'd31839, 16'd40880, 16'd47187, 16'd34073, 16'd19155, 16'd50752, 16'd24298, 16'd3821, 16'd10441, 16'd2752, 16'd17920, 16'd60207, 16'd43501, 16'd37327, 16'd31370, 16'd1367, 16'd33611, 16'd22936, 16'd26857, 16'd40306, 16'd53959, 16'd11145, 16'd36716, 16'd63555, 16'd30226});
	test_expansion(128'hb5914b648aeb8aa7e39696b71030a1da, {16'd17126, 16'd28802, 16'd35302, 16'd6830, 16'd54960, 16'd55812, 16'd53192, 16'd5581, 16'd25639, 16'd48321, 16'd14463, 16'd18923, 16'd11963, 16'd48513, 16'd9383, 16'd11276, 16'd7193, 16'd42319, 16'd40128, 16'd35633, 16'd21156, 16'd29818, 16'd54664, 16'd8250, 16'd6689, 16'd47652});
	test_expansion(128'h07c09ee338170fa056cb8540f06bd315, {16'd24909, 16'd64513, 16'd44592, 16'd15213, 16'd58115, 16'd23653, 16'd58670, 16'd31217, 16'd53895, 16'd48173, 16'd48305, 16'd13434, 16'd14385, 16'd58430, 16'd2787, 16'd763, 16'd49971, 16'd1661, 16'd26481, 16'd46299, 16'd3500, 16'd40079, 16'd1156, 16'd18740, 16'd42323, 16'd5381});
	test_expansion(128'hfbdc116dd337901af870c2c99c091eb2, {16'd64886, 16'd26781, 16'd20880, 16'd54530, 16'd41536, 16'd64705, 16'd53890, 16'd52079, 16'd65, 16'd20674, 16'd46530, 16'd15479, 16'd58664, 16'd52963, 16'd37322, 16'd3706, 16'd12985, 16'd35291, 16'd62911, 16'd43955, 16'd8918, 16'd63208, 16'd6891, 16'd8116, 16'd10391, 16'd39026});
	test_expansion(128'h016a4305f7dea366cf91dd99383797ee, {16'd53048, 16'd1715, 16'd57666, 16'd5358, 16'd5857, 16'd47832, 16'd54423, 16'd27326, 16'd35811, 16'd25827, 16'd28668, 16'd42397, 16'd21497, 16'd452, 16'd52388, 16'd54535, 16'd30918, 16'd60735, 16'd44061, 16'd12782, 16'd10406, 16'd46141, 16'd30640, 16'd20900, 16'd33805, 16'd38510});
	test_expansion(128'h413c605967726207f41b16a90d85e98d, {16'd41137, 16'd21955, 16'd61966, 16'd348, 16'd17306, 16'd10813, 16'd47675, 16'd49153, 16'd34528, 16'd6376, 16'd3553, 16'd52947, 16'd33773, 16'd13777, 16'd31393, 16'd1639, 16'd8406, 16'd45608, 16'd31914, 16'd64253, 16'd37044, 16'd37008, 16'd59188, 16'd793, 16'd26466, 16'd5907});
	test_expansion(128'h67083fe5e1e0fad525f020dc05202d3c, {16'd56572, 16'd62004, 16'd54480, 16'd49138, 16'd39924, 16'd7794, 16'd59328, 16'd37421, 16'd46963, 16'd1176, 16'd37468, 16'd5147, 16'd52577, 16'd3439, 16'd40998, 16'd13943, 16'd38040, 16'd54429, 16'd46464, 16'd55161, 16'd43973, 16'd58415, 16'd9619, 16'd43942, 16'd41133, 16'd11977});
	test_expansion(128'hc8241300e730e29a30e5ad57d53c514a, {16'd32407, 16'd35365, 16'd31976, 16'd4711, 16'd25925, 16'd36444, 16'd22422, 16'd50823, 16'd32703, 16'd44505, 16'd51169, 16'd54347, 16'd57202, 16'd33469, 16'd50520, 16'd11354, 16'd27102, 16'd42367, 16'd12854, 16'd56070, 16'd63052, 16'd234, 16'd45460, 16'd16281, 16'd38152, 16'd60219});
	test_expansion(128'hf958e776bc2bd7a32ae57453bdd8cb79, {16'd34672, 16'd60174, 16'd25537, 16'd29964, 16'd20693, 16'd47460, 16'd47314, 16'd7240, 16'd65053, 16'd61753, 16'd56603, 16'd14381, 16'd30267, 16'd34327, 16'd230, 16'd45765, 16'd16003, 16'd18922, 16'd54785, 16'd58698, 16'd7409, 16'd4071, 16'd47848, 16'd14411, 16'd52932, 16'd52067});
	test_expansion(128'hecce535cb9b58eec85b848755865cf90, {16'd46131, 16'd38560, 16'd62770, 16'd40222, 16'd46126, 16'd46289, 16'd14586, 16'd12428, 16'd27090, 16'd50431, 16'd56446, 16'd39181, 16'd11501, 16'd53843, 16'd50821, 16'd19023, 16'd39799, 16'd14350, 16'd25135, 16'd2647, 16'd3907, 16'd3614, 16'd4640, 16'd29766, 16'd56366, 16'd61331});
	test_expansion(128'hc7ebb7e8af8e70c5125b25ccae3e3f60, {16'd22788, 16'd15045, 16'd14521, 16'd37658, 16'd39162, 16'd52975, 16'd45209, 16'd7, 16'd15945, 16'd2129, 16'd50559, 16'd14640, 16'd49745, 16'd49974, 16'd20987, 16'd40621, 16'd56001, 16'd40986, 16'd40243, 16'd49011, 16'd12621, 16'd35372, 16'd44267, 16'd58413, 16'd4446, 16'd15715});
	test_expansion(128'hbdf11028b2b7a9378e84b509c230b9c9, {16'd24025, 16'd26493, 16'd32196, 16'd12965, 16'd18318, 16'd61221, 16'd1669, 16'd43017, 16'd44808, 16'd22243, 16'd52856, 16'd1738, 16'd55108, 16'd8682, 16'd58707, 16'd7126, 16'd30950, 16'd9149, 16'd48618, 16'd51082, 16'd9376, 16'd49136, 16'd9649, 16'd61955, 16'd63323, 16'd33863});
	test_expansion(128'h0f5c9ac1cf96935dca0cb41ff3965739, {16'd9371, 16'd36896, 16'd23940, 16'd10869, 16'd28094, 16'd48424, 16'd53750, 16'd19270, 16'd15164, 16'd21549, 16'd30552, 16'd94, 16'd43601, 16'd52210, 16'd6236, 16'd1878, 16'd39535, 16'd48481, 16'd51168, 16'd7994, 16'd29690, 16'd47999, 16'd42710, 16'd31737, 16'd28824, 16'd57909});
	test_expansion(128'h05e618f9c75645ca9f01f3a2e883521e, {16'd13378, 16'd197, 16'd50199, 16'd2632, 16'd36558, 16'd46007, 16'd19314, 16'd49097, 16'd25056, 16'd21652, 16'd52623, 16'd58116, 16'd14108, 16'd33790, 16'd37475, 16'd19274, 16'd52672, 16'd13258, 16'd37550, 16'd41843, 16'd55405, 16'd46612, 16'd53707, 16'd2062, 16'd33960, 16'd3598});
	test_expansion(128'h7956d205fade5e7e621abdf6159c5846, {16'd6975, 16'd12131, 16'd17377, 16'd21309, 16'd61598, 16'd45509, 16'd51079, 16'd47065, 16'd14783, 16'd20296, 16'd43519, 16'd21715, 16'd4945, 16'd14054, 16'd46272, 16'd20794, 16'd19382, 16'd56723, 16'd41051, 16'd22116, 16'd11066, 16'd53680, 16'd14713, 16'd34653, 16'd50109, 16'd20512});
	test_expansion(128'hcbf86203967f7b193da72e0025e8abdb, {16'd2024, 16'd34555, 16'd53191, 16'd43747, 16'd17160, 16'd4901, 16'd34896, 16'd53799, 16'd22887, 16'd27633, 16'd14328, 16'd60854, 16'd11075, 16'd22940, 16'd12207, 16'd61639, 16'd8186, 16'd27636, 16'd18714, 16'd48549, 16'd44558, 16'd54911, 16'd34894, 16'd22611, 16'd30322, 16'd34050});
	test_expansion(128'h711b96fd0347a14fe7c7ca9efc2bdc4e, {16'd14720, 16'd26906, 16'd13479, 16'd14484, 16'd38685, 16'd55473, 16'd42324, 16'd21265, 16'd10575, 16'd33600, 16'd13789, 16'd22300, 16'd28470, 16'd44423, 16'd53643, 16'd28821, 16'd49187, 16'd14613, 16'd20, 16'd33879, 16'd43868, 16'd61560, 16'd17640, 16'd9319, 16'd52895, 16'd29591});
	test_expansion(128'hf737d2c09dd608f9fb491f9014173bb4, {16'd15117, 16'd51388, 16'd2867, 16'd58401, 16'd7646, 16'd47881, 16'd9439, 16'd36921, 16'd43033, 16'd51152, 16'd26516, 16'd927, 16'd43761, 16'd14003, 16'd29511, 16'd17665, 16'd19441, 16'd22982, 16'd9301, 16'd54276, 16'd35640, 16'd55505, 16'd55616, 16'd48784, 16'd7461, 16'd172});
	test_expansion(128'hc5a2cc4bb268e53b0a4f8681b5d02580, {16'd37452, 16'd31145, 16'd45536, 16'd61171, 16'd64324, 16'd41288, 16'd2492, 16'd18560, 16'd11958, 16'd1388, 16'd41542, 16'd40252, 16'd14110, 16'd37987, 16'd35771, 16'd24343, 16'd36682, 16'd26041, 16'd56388, 16'd64856, 16'd47497, 16'd11622, 16'd40525, 16'd13395, 16'd3875, 16'd10010});
	test_expansion(128'ha874950ae52377b505529b87f6ddbe93, {16'd16017, 16'd37081, 16'd14423, 16'd37689, 16'd54301, 16'd39357, 16'd15933, 16'd56525, 16'd3654, 16'd44390, 16'd27527, 16'd23786, 16'd26162, 16'd42968, 16'd23747, 16'd62852, 16'd35028, 16'd57352, 16'd33910, 16'd39097, 16'd19538, 16'd53371, 16'd48388, 16'd59765, 16'd43230, 16'd56484});
	test_expansion(128'hb0af9883c9d8383d76f23bb678e5b9db, {16'd46767, 16'd55441, 16'd8368, 16'd13391, 16'd1906, 16'd21701, 16'd47061, 16'd11199, 16'd62614, 16'd13192, 16'd52811, 16'd65340, 16'd18988, 16'd7802, 16'd10909, 16'd29004, 16'd52332, 16'd8741, 16'd61044, 16'd6486, 16'd51956, 16'd27303, 16'd46014, 16'd22573, 16'd18778, 16'd35373});
	test_expansion(128'hb13a24a68dbe3daab10ed42251aeec13, {16'd62528, 16'd15405, 16'd16305, 16'd27062, 16'd46262, 16'd59167, 16'd41410, 16'd7980, 16'd49508, 16'd28783, 16'd3433, 16'd53771, 16'd18923, 16'd57169, 16'd14241, 16'd32679, 16'd21147, 16'd6081, 16'd60454, 16'd42662, 16'd50234, 16'd50897, 16'd17364, 16'd34725, 16'd7091, 16'd54627});
	test_expansion(128'h3a6fd6664e830af1ba4522738e0ad1b9, {16'd23151, 16'd23753, 16'd6900, 16'd37876, 16'd35364, 16'd49514, 16'd51537, 16'd52822, 16'd54287, 16'd48123, 16'd51588, 16'd5726, 16'd28632, 16'd63495, 16'd24028, 16'd9338, 16'd25347, 16'd49884, 16'd21242, 16'd21863, 16'd58611, 16'd12042, 16'd43232, 16'd47318, 16'd63839, 16'd61639});
	test_expansion(128'h35ea6b189a521ebd1a8e831e76237eb2, {16'd35927, 16'd50885, 16'd10332, 16'd52450, 16'd756, 16'd31200, 16'd49353, 16'd6961, 16'd46192, 16'd4108, 16'd54894, 16'd54390, 16'd31856, 16'd47009, 16'd1659, 16'd41259, 16'd15573, 16'd58636, 16'd20792, 16'd33584, 16'd22324, 16'd28972, 16'd1542, 16'd24942, 16'd51859, 16'd64234});
	test_expansion(128'h6ced540196a1f44abb89bb68beebbf33, {16'd28001, 16'd39070, 16'd4359, 16'd55554, 16'd33095, 16'd64602, 16'd19488, 16'd10502, 16'd58157, 16'd7461, 16'd1992, 16'd39846, 16'd7099, 16'd20256, 16'd15125, 16'd57759, 16'd31684, 16'd60141, 16'd39269, 16'd24866, 16'd40668, 16'd31490, 16'd39941, 16'd47180, 16'd40280, 16'd13909});
	test_expansion(128'ha03cd9de238ae7268b892f01e34d9963, {16'd50943, 16'd40966, 16'd45275, 16'd27391, 16'd46014, 16'd48357, 16'd34881, 16'd19595, 16'd10995, 16'd30640, 16'd6470, 16'd12454, 16'd4296, 16'd35505, 16'd64554, 16'd51847, 16'd738, 16'd51953, 16'd42062, 16'd43581, 16'd60422, 16'd42573, 16'd29249, 16'd31860, 16'd60203, 16'd5643});
	test_expansion(128'h1b2b3970553b8e2d719c0b1dfe839129, {16'd58499, 16'd39138, 16'd2851, 16'd54889, 16'd32801, 16'd8633, 16'd24334, 16'd17696, 16'd8515, 16'd31737, 16'd28878, 16'd3491, 16'd19864, 16'd43779, 16'd48887, 16'd21945, 16'd4989, 16'd28448, 16'd9673, 16'd11910, 16'd19591, 16'd33168, 16'd38495, 16'd52800, 16'd1729, 16'd24906});
	test_expansion(128'h6dd06e967b81548c57761bf1c392d23a, {16'd6316, 16'd54520, 16'd51437, 16'd15603, 16'd13159, 16'd49647, 16'd3625, 16'd2693, 16'd64494, 16'd14878, 16'd48255, 16'd13526, 16'd9128, 16'd41277, 16'd50781, 16'd35984, 16'd157, 16'd46970, 16'd121, 16'd8998, 16'd63246, 16'd37069, 16'd31976, 16'd19861, 16'd31944, 16'd39191});
	test_expansion(128'h000b3b31eab88a79625d139566fdb4c8, {16'd23666, 16'd57474, 16'd49549, 16'd29678, 16'd14861, 16'd32192, 16'd20416, 16'd23714, 16'd60918, 16'd5493, 16'd62553, 16'd31372, 16'd38076, 16'd33861, 16'd26552, 16'd1476, 16'd49163, 16'd23566, 16'd58109, 16'd42518, 16'd39591, 16'd8564, 16'd7538, 16'd4681, 16'd36282, 16'd2630});
	test_expansion(128'hca0f11a3f85a7a1eeab0d539ba0abc49, {16'd33537, 16'd11074, 16'd14394, 16'd11631, 16'd27645, 16'd32725, 16'd45840, 16'd34541, 16'd3359, 16'd60874, 16'd9332, 16'd65369, 16'd25905, 16'd4835, 16'd64121, 16'd30661, 16'd62930, 16'd18267, 16'd56322, 16'd6856, 16'd29774, 16'd4884, 16'd51494, 16'd38302, 16'd2421, 16'd10852});
	test_expansion(128'he04950a4aefb8ab60bc44d8caa200d7b, {16'd50202, 16'd26856, 16'd54764, 16'd33131, 16'd59958, 16'd23166, 16'd12014, 16'd25123, 16'd49073, 16'd30541, 16'd49642, 16'd8712, 16'd36287, 16'd15392, 16'd18615, 16'd58491, 16'd57945, 16'd13574, 16'd4363, 16'd60005, 16'd6133, 16'd14257, 16'd63157, 16'd20259, 16'd2524, 16'd52248});
	test_expansion(128'h3998815dc2a786a2b05f4560c0e6bd94, {16'd40217, 16'd54299, 16'd58038, 16'd52859, 16'd56986, 16'd48220, 16'd55963, 16'd50892, 16'd19015, 16'd60605, 16'd8699, 16'd59144, 16'd38760, 16'd616, 16'd58921, 16'd45867, 16'd20966, 16'd32949, 16'd56428, 16'd16920, 16'd22524, 16'd41365, 16'd18377, 16'd11771, 16'd13766, 16'd58338});
	test_expansion(128'h52405b0e40c4560d905e851312f9d5af, {16'd48010, 16'd38114, 16'd19486, 16'd56461, 16'd53421, 16'd42382, 16'd51690, 16'd12487, 16'd53184, 16'd17526, 16'd41445, 16'd19339, 16'd60131, 16'd55694, 16'd57680, 16'd42040, 16'd8608, 16'd37039, 16'd7940, 16'd24336, 16'd21751, 16'd20668, 16'd38130, 16'd30086, 16'd38267, 16'd39007});
	test_expansion(128'h5cce5312dd0f0d820ed8609a106215bf, {16'd48502, 16'd31694, 16'd431, 16'd61472, 16'd21039, 16'd38438, 16'd13638, 16'd12411, 16'd36183, 16'd51018, 16'd7469, 16'd33610, 16'd52484, 16'd7095, 16'd20050, 16'd38596, 16'd41528, 16'd60183, 16'd36866, 16'd12738, 16'd58341, 16'd42395, 16'd28735, 16'd22038, 16'd53346, 16'd55764});
	test_expansion(128'hd40c30bb3d6df09737cdfc1fda178ac6, {16'd50953, 16'd38180, 16'd1765, 16'd50898, 16'd64284, 16'd18287, 16'd48684, 16'd41787, 16'd57136, 16'd51480, 16'd1150, 16'd25339, 16'd8432, 16'd27739, 16'd879, 16'd41212, 16'd51005, 16'd18356, 16'd952, 16'd62710, 16'd42899, 16'd53889, 16'd22754, 16'd65154, 16'd31954, 16'd32991});
	test_expansion(128'h98713dada47d0d61891f1de0711c9306, {16'd15701, 16'd22744, 16'd59711, 16'd43120, 16'd38574, 16'd43513, 16'd4790, 16'd47391, 16'd48071, 16'd42520, 16'd8478, 16'd17598, 16'd7491, 16'd47890, 16'd45048, 16'd12378, 16'd858, 16'd6148, 16'd53555, 16'd275, 16'd52692, 16'd35350, 16'd23308, 16'd19153, 16'd740, 16'd44842});
	test_expansion(128'h765a6a404aa01635163285d6f9963ff0, {16'd57831, 16'd1303, 16'd25228, 16'd53177, 16'd49691, 16'd17548, 16'd19191, 16'd18648, 16'd10531, 16'd51201, 16'd63755, 16'd7668, 16'd48399, 16'd12563, 16'd36845, 16'd61071, 16'd22042, 16'd17825, 16'd5911, 16'd42788, 16'd1073, 16'd16334, 16'd18736, 16'd53761, 16'd62055, 16'd37374});
	test_expansion(128'hff2da026ddb0d5d998265a4eee10bb30, {16'd33316, 16'd44866, 16'd19897, 16'd4230, 16'd33868, 16'd44335, 16'd46526, 16'd16750, 16'd61707, 16'd10686, 16'd53919, 16'd12221, 16'd64449, 16'd62405, 16'd51861, 16'd28304, 16'd43556, 16'd18087, 16'd20947, 16'd6556, 16'd64735, 16'd52318, 16'd63234, 16'd46396, 16'd14256, 16'd35334});
	test_expansion(128'ha7fb2eed32fe6eb3fc4544b98eeea596, {16'd17306, 16'd56927, 16'd26749, 16'd6162, 16'd10360, 16'd6896, 16'd17747, 16'd18894, 16'd50261, 16'd58826, 16'd50446, 16'd58595, 16'd1754, 16'd54417, 16'd18761, 16'd50254, 16'd46, 16'd45265, 16'd6408, 16'd33589, 16'd38811, 16'd20534, 16'd40209, 16'd390, 16'd46358, 16'd47363});
	test_expansion(128'hdf66baab90cb132535ba8b4a20add0ea, {16'd62251, 16'd17975, 16'd10109, 16'd62539, 16'd4076, 16'd6679, 16'd56494, 16'd47189, 16'd55067, 16'd32375, 16'd39329, 16'd27462, 16'd57341, 16'd25783, 16'd16101, 16'd52522, 16'd37383, 16'd23401, 16'd36764, 16'd39811, 16'd58028, 16'd61796, 16'd18457, 16'd23754, 16'd49355, 16'd17258});
	test_expansion(128'hcc0ea52db55d66689ab2ab11cfd1a97f, {16'd12458, 16'd14692, 16'd4908, 16'd12252, 16'd59416, 16'd35585, 16'd7592, 16'd1073, 16'd23213, 16'd28724, 16'd39459, 16'd29162, 16'd12728, 16'd44591, 16'd60790, 16'd45046, 16'd23235, 16'd16070, 16'd23506, 16'd20719, 16'd14477, 16'd9753, 16'd31468, 16'd51028, 16'd25834, 16'd60888});
	test_expansion(128'h18c39b2f3996fa39f0a1010fc8a93a2e, {16'd18974, 16'd44318, 16'd52188, 16'd26342, 16'd62430, 16'd51823, 16'd14866, 16'd19304, 16'd47140, 16'd37873, 16'd3530, 16'd15431, 16'd26622, 16'd26448, 16'd56179, 16'd9002, 16'd12369, 16'd45114, 16'd46863, 16'd60120, 16'd7127, 16'd53712, 16'd26289, 16'd20390, 16'd10959, 16'd60781});
	test_expansion(128'h82d7c7b04e93c323cfa8298716b99005, {16'd16760, 16'd868, 16'd12920, 16'd12165, 16'd41313, 16'd37713, 16'd24039, 16'd40644, 16'd63650, 16'd25611, 16'd2239, 16'd64340, 16'd37972, 16'd41748, 16'd24742, 16'd52959, 16'd30379, 16'd63051, 16'd41714, 16'd37080, 16'd61079, 16'd196, 16'd33177, 16'd28404, 16'd36660, 16'd1959});
	test_expansion(128'h8fbbf194b7cb8897b7293eb2d4fca991, {16'd15060, 16'd57231, 16'd142, 16'd36418, 16'd11091, 16'd31444, 16'd62717, 16'd27136, 16'd8995, 16'd409, 16'd63335, 16'd3999, 16'd45859, 16'd22946, 16'd32264, 16'd45772, 16'd51232, 16'd27258, 16'd53926, 16'd13583, 16'd30369, 16'd32264, 16'd65524, 16'd49050, 16'd7902, 16'd7775});
	test_expansion(128'hed04bdd95fc5a0972a3c32e7dae15251, {16'd43107, 16'd33886, 16'd35016, 16'd53103, 16'd2383, 16'd14455, 16'd7513, 16'd60501, 16'd7402, 16'd45717, 16'd47284, 16'd6130, 16'd20590, 16'd24312, 16'd51566, 16'd32854, 16'd22834, 16'd57202, 16'd52816, 16'd4761, 16'd64247, 16'd65458, 16'd11907, 16'd50520, 16'd36155, 16'd32602});
	test_expansion(128'h46196e54f8facbaa960541a60e1baa27, {16'd7647, 16'd22782, 16'd1337, 16'd58659, 16'd45106, 16'd49438, 16'd16394, 16'd46716, 16'd687, 16'd46209, 16'd15256, 16'd30616, 16'd61073, 16'd29497, 16'd369, 16'd57391, 16'd26773, 16'd47465, 16'd17235, 16'd25926, 16'd27694, 16'd52323, 16'd65411, 16'd45029, 16'd19394, 16'd48947});
	test_expansion(128'habfdca7f68dcf23bb30032d84d254d9b, {16'd26379, 16'd48916, 16'd4691, 16'd26701, 16'd32336, 16'd45494, 16'd63616, 16'd12270, 16'd32301, 16'd30648, 16'd34950, 16'd24078, 16'd50829, 16'd62806, 16'd62899, 16'd6858, 16'd45098, 16'd63414, 16'd49200, 16'd25558, 16'd61271, 16'd17337, 16'd46857, 16'd50417, 16'd61478, 16'd13295});
	test_expansion(128'hee943702fcfd2d3f4ad72f099334a34a, {16'd43496, 16'd4476, 16'd46813, 16'd27822, 16'd34918, 16'd12912, 16'd43303, 16'd51599, 16'd45882, 16'd20348, 16'd65487, 16'd64185, 16'd45517, 16'd34353, 16'd12756, 16'd37614, 16'd46235, 16'd31926, 16'd63231, 16'd31064, 16'd36916, 16'd48181, 16'd50232, 16'd26160, 16'd14735, 16'd19952});
	test_expansion(128'hea282b29d65b636d4f43e5da55d17395, {16'd19987, 16'd23421, 16'd41474, 16'd61151, 16'd3724, 16'd39072, 16'd54429, 16'd15367, 16'd29301, 16'd52864, 16'd56204, 16'd1346, 16'd63554, 16'd57716, 16'd32034, 16'd53189, 16'd37480, 16'd36330, 16'd3576, 16'd2546, 16'd19159, 16'd5823, 16'd13220, 16'd53106, 16'd50876, 16'd29471});
	test_expansion(128'h032bcb1ce55a11cf2833b7c914548286, {16'd14505, 16'd55248, 16'd62275, 16'd9765, 16'd32380, 16'd52794, 16'd27230, 16'd20110, 16'd19418, 16'd4248, 16'd32547, 16'd42562, 16'd53150, 16'd21588, 16'd3083, 16'd23136, 16'd64932, 16'd7036, 16'd33335, 16'd42852, 16'd2413, 16'd44309, 16'd38149, 16'd18152, 16'd21274, 16'd27285});
	test_expansion(128'h3128be62c3c4c44b5755c4f8743cb7a3, {16'd10623, 16'd8449, 16'd29595, 16'd53713, 16'd37503, 16'd14963, 16'd26159, 16'd55281, 16'd18153, 16'd12187, 16'd7591, 16'd35653, 16'd34314, 16'd3921, 16'd14990, 16'd28713, 16'd14156, 16'd52467, 16'd61471, 16'd25976, 16'd51977, 16'd55423, 16'd63652, 16'd19559, 16'd12106, 16'd50966});
	test_expansion(128'hffe3160bb1d60e6fc51e6f1fbe97a34a, {16'd57930, 16'd38826, 16'd53461, 16'd26066, 16'd53092, 16'd59208, 16'd26514, 16'd56137, 16'd21848, 16'd41271, 16'd65332, 16'd19671, 16'd51554, 16'd53843, 16'd38294, 16'd56086, 16'd21693, 16'd49014, 16'd41449, 16'd19390, 16'd9771, 16'd28352, 16'd51669, 16'd28449, 16'd56210, 16'd32192});
	test_expansion(128'h957d7c1f8766380e5215cf2901c907be, {16'd36228, 16'd40406, 16'd26348, 16'd47461, 16'd10345, 16'd62115, 16'd33971, 16'd7461, 16'd327, 16'd47567, 16'd42161, 16'd43394, 16'd11655, 16'd45616, 16'd64401, 16'd47910, 16'd44200, 16'd64877, 16'd6721, 16'd598, 16'd35317, 16'd3782, 16'd60606, 16'd29599, 16'd41597, 16'd29891});
	test_expansion(128'hac4fc51d856408a2e4af1def2ab034bb, {16'd14207, 16'd18907, 16'd35241, 16'd3892, 16'd8584, 16'd37729, 16'd47466, 16'd18463, 16'd46364, 16'd28520, 16'd23211, 16'd13487, 16'd11147, 16'd22201, 16'd25402, 16'd8717, 16'd20814, 16'd12795, 16'd2594, 16'd40340, 16'd4335, 16'd12971, 16'd49206, 16'd8620, 16'd42785, 16'd13961});
	test_expansion(128'h4d7aba5ffbf00211b3ed70ac5d5f7a1b, {16'd20428, 16'd27129, 16'd31685, 16'd50816, 16'd6747, 16'd14431, 16'd32992, 16'd46612, 16'd27214, 16'd54214, 16'd10935, 16'd60710, 16'd50259, 16'd57573, 16'd32169, 16'd10252, 16'd56069, 16'd57217, 16'd26403, 16'd35081, 16'd13591, 16'd59774, 16'd29519, 16'd4433, 16'd53161, 16'd49576});
	test_expansion(128'hcec680e76d70f7f9b2ba16a0aec7b7b6, {16'd49588, 16'd39983, 16'd4932, 16'd30685, 16'd16163, 16'd59155, 16'd5142, 16'd11351, 16'd43444, 16'd30111, 16'd9196, 16'd58307, 16'd27415, 16'd54609, 16'd48383, 16'd5541, 16'd37834, 16'd27293, 16'd35135, 16'd25921, 16'd51118, 16'd30449, 16'd35399, 16'd43766, 16'd37377, 16'd6084});
	test_expansion(128'hdfc0328ef059e40a49d052f40af41231, {16'd4119, 16'd53955, 16'd39829, 16'd40992, 16'd8193, 16'd41408, 16'd42126, 16'd7498, 16'd2989, 16'd62374, 16'd60913, 16'd31394, 16'd33938, 16'd35378, 16'd6410, 16'd55122, 16'd26468, 16'd13831, 16'd51649, 16'd10823, 16'd45976, 16'd49927, 16'd6017, 16'd19323, 16'd21789, 16'd62340});
	test_expansion(128'hce47c258299102d006b8edc34b5aaa52, {16'd13927, 16'd27762, 16'd34529, 16'd46381, 16'd29117, 16'd20006, 16'd9837, 16'd31726, 16'd57764, 16'd10077, 16'd28419, 16'd10187, 16'd8576, 16'd40060, 16'd41617, 16'd1484, 16'd1345, 16'd65157, 16'd10962, 16'd4198, 16'd22247, 16'd22579, 16'd726, 16'd43189, 16'd64997, 16'd25528});
	test_expansion(128'h111889c11bccdff1c58aa9e248c49792, {16'd7664, 16'd62533, 16'd37735, 16'd3454, 16'd834, 16'd18948, 16'd17667, 16'd28484, 16'd33729, 16'd15275, 16'd55529, 16'd32156, 16'd12419, 16'd56014, 16'd8100, 16'd31908, 16'd8181, 16'd58808, 16'd39932, 16'd6536, 16'd55819, 16'd54002, 16'd32254, 16'd36759, 16'd51872, 16'd44123});
	test_expansion(128'hc9d3e77069a4b8604e36c88e11f5a4c4, {16'd39658, 16'd2434, 16'd42746, 16'd47153, 16'd28536, 16'd46929, 16'd28096, 16'd64530, 16'd45599, 16'd53086, 16'd3280, 16'd9491, 16'd7522, 16'd45106, 16'd42981, 16'd59905, 16'd25387, 16'd43100, 16'd22428, 16'd61138, 16'd53216, 16'd10494, 16'd29721, 16'd39553, 16'd34364, 16'd52340});
	test_expansion(128'h0063108466503149f6ffce316cfb7f38, {16'd13277, 16'd10298, 16'd43764, 16'd44020, 16'd64887, 16'd4676, 16'd55144, 16'd42046, 16'd396, 16'd21720, 16'd16642, 16'd22872, 16'd39694, 16'd38467, 16'd22210, 16'd22402, 16'd47061, 16'd3693, 16'd24800, 16'd23053, 16'd64179, 16'd20726, 16'd1918, 16'd53299, 16'd15062, 16'd19945});
	test_expansion(128'he9335bfb8688ae34c13c99a47fb28c17, {16'd19483, 16'd5508, 16'd25184, 16'd32081, 16'd8704, 16'd14622, 16'd10204, 16'd52364, 16'd55402, 16'd7796, 16'd23881, 16'd35569, 16'd48797, 16'd58429, 16'd39959, 16'd48623, 16'd60879, 16'd40467, 16'd40416, 16'd58628, 16'd54738, 16'd10217, 16'd11470, 16'd2708, 16'd61335, 16'd59452});
	test_expansion(128'heb8255afcce2162599f6e65f3d5edced, {16'd6881, 16'd37256, 16'd9996, 16'd11588, 16'd49500, 16'd3813, 16'd7677, 16'd25246, 16'd12379, 16'd12935, 16'd5600, 16'd14263, 16'd56635, 16'd23840, 16'd29636, 16'd36149, 16'd26851, 16'd52454, 16'd52823, 16'd41263, 16'd27749, 16'd6979, 16'd18685, 16'd20165, 16'd62220, 16'd31464});
	test_expansion(128'h9093eaa53d7768a0b5c4020fcd058db3, {16'd4911, 16'd38983, 16'd44264, 16'd24749, 16'd1528, 16'd38034, 16'd56763, 16'd54706, 16'd23739, 16'd35434, 16'd10063, 16'd62906, 16'd1668, 16'd19283, 16'd18469, 16'd29053, 16'd63816, 16'd20208, 16'd9888, 16'd34045, 16'd64496, 16'd46454, 16'd10710, 16'd62339, 16'd48468, 16'd44831});
	test_expansion(128'h849e0959b151aedcfd6343d2c952a925, {16'd49029, 16'd16889, 16'd55299, 16'd14316, 16'd57256, 16'd1696, 16'd13548, 16'd64645, 16'd6958, 16'd8118, 16'd16691, 16'd29642, 16'd16480, 16'd42543, 16'd18728, 16'd61967, 16'd24548, 16'd8089, 16'd64997, 16'd55659, 16'd63465, 16'd12853, 16'd15453, 16'd28637, 16'd33602, 16'd50896});
	test_expansion(128'h7cd02439a0612a2c51660f7b29f1fe14, {16'd37589, 16'd8388, 16'd62319, 16'd24365, 16'd43154, 16'd19474, 16'd47153, 16'd7533, 16'd41163, 16'd55274, 16'd2523, 16'd37341, 16'd38662, 16'd55362, 16'd4330, 16'd25088, 16'd57177, 16'd45346, 16'd5811, 16'd2830, 16'd34897, 16'd28857, 16'd37171, 16'd19623, 16'd62775, 16'd4688});
	test_expansion(128'h9fa413b2bad2cdbac2c6381d62233885, {16'd47395, 16'd60926, 16'd21853, 16'd26066, 16'd30801, 16'd14706, 16'd56929, 16'd46883, 16'd2434, 16'd22249, 16'd47464, 16'd44089, 16'd48112, 16'd35586, 16'd61706, 16'd18939, 16'd53500, 16'd24353, 16'd53045, 16'd25459, 16'd36745, 16'd56702, 16'd42965, 16'd56479, 16'd21846, 16'd20484});
	test_expansion(128'haca595b30d2f98310c762941e33204d3, {16'd21361, 16'd30940, 16'd45999, 16'd55930, 16'd24586, 16'd22652, 16'd20545, 16'd16210, 16'd65111, 16'd45779, 16'd26637, 16'd30893, 16'd33484, 16'd41918, 16'd15943, 16'd12596, 16'd46995, 16'd46991, 16'd16638, 16'd454, 16'd1996, 16'd24614, 16'd46951, 16'd58324, 16'd34436, 16'd14543});
	test_expansion(128'hfe137edbb1a84ed04d2d5c71d69dd5cc, {16'd50010, 16'd42407, 16'd64821, 16'd53253, 16'd1203, 16'd46192, 16'd63144, 16'd44072, 16'd2124, 16'd54548, 16'd62813, 16'd21744, 16'd34090, 16'd38191, 16'd1087, 16'd22483, 16'd14967, 16'd21251, 16'd49787, 16'd25033, 16'd39291, 16'd52300, 16'd55586, 16'd8005, 16'd57599, 16'd20606});
	test_expansion(128'h43d5e35c8fab09c6c7f26e3c8270daf4, {16'd60788, 16'd58768, 16'd49109, 16'd8096, 16'd34206, 16'd28570, 16'd43066, 16'd25342, 16'd33139, 16'd14350, 16'd1063, 16'd46922, 16'd27307, 16'd37737, 16'd11155, 16'd29411, 16'd38137, 16'd63408, 16'd35325, 16'd17337, 16'd1665, 16'd38879, 16'd45578, 16'd53102, 16'd27755, 16'd54220});
	test_expansion(128'h78a8054f1b0b0c98646e4db661e69976, {16'd57764, 16'd42111, 16'd37909, 16'd16502, 16'd16845, 16'd6791, 16'd9809, 16'd34094, 16'd12070, 16'd31097, 16'd6331, 16'd27391, 16'd12639, 16'd6605, 16'd30381, 16'd31713, 16'd32294, 16'd48566, 16'd48836, 16'd31371, 16'd46067, 16'd36376, 16'd10547, 16'd36137, 16'd21350, 16'd33261});
	test_expansion(128'hbf34b612956bb12c3001122ab095156f, {16'd11816, 16'd65047, 16'd22242, 16'd63106, 16'd58265, 16'd56435, 16'd57071, 16'd55280, 16'd42606, 16'd2733, 16'd31398, 16'd2227, 16'd28866, 16'd43633, 16'd22703, 16'd40395, 16'd40025, 16'd59084, 16'd16556, 16'd41871, 16'd22523, 16'd17841, 16'd29769, 16'd58861, 16'd57132, 16'd8242});
	test_expansion(128'hc0fffd88462886cc9357882fef590a47, {16'd3244, 16'd21734, 16'd3728, 16'd29934, 16'd32545, 16'd32002, 16'd37868, 16'd11377, 16'd51712, 16'd33860, 16'd55570, 16'd51382, 16'd81, 16'd33188, 16'd24177, 16'd51937, 16'd56441, 16'd56970, 16'd33931, 16'd41815, 16'd1307, 16'd38520, 16'd57406, 16'd52156, 16'd35555, 16'd45782});
	test_expansion(128'h070373e2aef7b2e2842fbd43df0376dc, {16'd55588, 16'd39557, 16'd32691, 16'd35946, 16'd889, 16'd49106, 16'd23673, 16'd15803, 16'd43548, 16'd3320, 16'd20751, 16'd1826, 16'd29079, 16'd63252, 16'd58662, 16'd32454, 16'd11025, 16'd55518, 16'd47880, 16'd23712, 16'd62815, 16'd55429, 16'd7707, 16'd49204, 16'd48844, 16'd15995});
	test_expansion(128'h72d3621769329f1a0eeed83a8e2c5970, {16'd47583, 16'd65130, 16'd32887, 16'd33123, 16'd50646, 16'd40534, 16'd59971, 16'd64493, 16'd5225, 16'd19474, 16'd41594, 16'd17666, 16'd61539, 16'd60357, 16'd1918, 16'd3577, 16'd45534, 16'd59011, 16'd8272, 16'd51583, 16'd46582, 16'd51303, 16'd58360, 16'd57938, 16'd29639, 16'd43056});
	test_expansion(128'h1939d3c95f3451f7994759b9a449d8ec, {16'd13877, 16'd28822, 16'd42194, 16'd7775, 16'd43785, 16'd16019, 16'd42803, 16'd11225, 16'd64062, 16'd14796, 16'd8792, 16'd7196, 16'd46018, 16'd62117, 16'd13364, 16'd5176, 16'd52015, 16'd52726, 16'd34327, 16'd24289, 16'd31776, 16'd41774, 16'd18435, 16'd22494, 16'd34185, 16'd54463});
	test_expansion(128'hecdd9f0e67cfb854f07818330dd8d071, {16'd54804, 16'd40763, 16'd37219, 16'd46445, 16'd54652, 16'd40098, 16'd16463, 16'd43981, 16'd21583, 16'd40576, 16'd26613, 16'd3451, 16'd47317, 16'd30532, 16'd11048, 16'd60354, 16'd29135, 16'd7140, 16'd61958, 16'd44594, 16'd5447, 16'd2578, 16'd39367, 16'd27327, 16'd3377, 16'd47080});
	test_expansion(128'h60da532ce62da029d626b0d976c6d300, {16'd15950, 16'd35287, 16'd17175, 16'd65380, 16'd9333, 16'd41862, 16'd58278, 16'd42472, 16'd29957, 16'd56455, 16'd13696, 16'd48479, 16'd46145, 16'd16397, 16'd20667, 16'd15417, 16'd53536, 16'd3072, 16'd11116, 16'd47910, 16'd38330, 16'd2357, 16'd49630, 16'd11176, 16'd51948, 16'd13515});
	test_expansion(128'h63e767aa804b343e2b3c46fb1ad65182, {16'd1657, 16'd19848, 16'd64530, 16'd57862, 16'd47946, 16'd64856, 16'd22825, 16'd47568, 16'd6129, 16'd4778, 16'd13254, 16'd32885, 16'd34330, 16'd10444, 16'd50342, 16'd3269, 16'd49721, 16'd64110, 16'd45156, 16'd13749, 16'd42948, 16'd53255, 16'd3851, 16'd24115, 16'd8208, 16'd35165});
	test_expansion(128'h67b9e27a1179434d82a7d243598248b8, {16'd51137, 16'd57746, 16'd42514, 16'd46745, 16'd41106, 16'd32015, 16'd49536, 16'd9703, 16'd6815, 16'd8239, 16'd7081, 16'd18913, 16'd53880, 16'd29170, 16'd672, 16'd26575, 16'd6929, 16'd57625, 16'd19143, 16'd27986, 16'd20972, 16'd35335, 16'd42399, 16'd58341, 16'd51469, 16'd19339});
	test_expansion(128'hb487b630aefa6cb4f2fc2bf01bf240c5, {16'd2868, 16'd64542, 16'd35648, 16'd1258, 16'd48199, 16'd33463, 16'd48518, 16'd47062, 16'd51611, 16'd61295, 16'd45620, 16'd21683, 16'd34291, 16'd3793, 16'd5768, 16'd11471, 16'd33432, 16'd34290, 16'd20459, 16'd48756, 16'd18376, 16'd60244, 16'd41340, 16'd17776, 16'd60745, 16'd45122});
	test_expansion(128'h90e37fad2300d6067d4d7a4a519b5cda, {16'd53549, 16'd56765, 16'd16073, 16'd31316, 16'd61962, 16'd47789, 16'd10910, 16'd65120, 16'd18737, 16'd30678, 16'd38640, 16'd53649, 16'd49875, 16'd20106, 16'd18809, 16'd30124, 16'd35124, 16'd12267, 16'd54598, 16'd8875, 16'd59545, 16'd33838, 16'd53359, 16'd11225, 16'd27556, 16'd58281});
	test_expansion(128'hf85e644456df4ff2f8add239ae61821a, {16'd53347, 16'd48161, 16'd65009, 16'd2078, 16'd44895, 16'd15344, 16'd43403, 16'd42331, 16'd26881, 16'd38851, 16'd52424, 16'd59874, 16'd34575, 16'd40479, 16'd61314, 16'd27518, 16'd64691, 16'd7516, 16'd55919, 16'd46647, 16'd37159, 16'd39085, 16'd3650, 16'd2728, 16'd36773, 16'd21415});
	test_expansion(128'h3a0dfe3bf88214a0654a0a52ba39473f, {16'd38129, 16'd11085, 16'd12688, 16'd14939, 16'd64139, 16'd22905, 16'd23353, 16'd12693, 16'd63542, 16'd43562, 16'd33412, 16'd22693, 16'd50149, 16'd27983, 16'd30216, 16'd1086, 16'd57161, 16'd31327, 16'd935, 16'd17878, 16'd47294, 16'd31331, 16'd20901, 16'd27957, 16'd13308, 16'd2761});
	test_expansion(128'hc4ddf5b741db6536fa1b746557c0ab25, {16'd64972, 16'd48616, 16'd2773, 16'd55541, 16'd48424, 16'd62371, 16'd32835, 16'd56318, 16'd40868, 16'd5714, 16'd12203, 16'd36156, 16'd42001, 16'd46546, 16'd1388, 16'd1271, 16'd62687, 16'd4722, 16'd24142, 16'd57273, 16'd1253, 16'd19866, 16'd12905, 16'd65000, 16'd29492, 16'd44337});
	test_expansion(128'hef379218b2082854aa2d89e79917da45, {16'd30205, 16'd45487, 16'd5094, 16'd8583, 16'd2556, 16'd22238, 16'd34105, 16'd42256, 16'd60409, 16'd51595, 16'd57006, 16'd63694, 16'd58812, 16'd31566, 16'd43758, 16'd24741, 16'd38994, 16'd46864, 16'd29266, 16'd41664, 16'd63119, 16'd17565, 16'd64270, 16'd57322, 16'd24731, 16'd9879});
	test_expansion(128'h00e81bfe902be2ff261fc16f80fbf7b1, {16'd22505, 16'd12308, 16'd8632, 16'd26249, 16'd45096, 16'd52872, 16'd32736, 16'd15275, 16'd46640, 16'd47777, 16'd39347, 16'd50256, 16'd38571, 16'd59993, 16'd20218, 16'd3004, 16'd65490, 16'd12423, 16'd44209, 16'd55468, 16'd44345, 16'd37915, 16'd34990, 16'd31950, 16'd23979, 16'd17794});
	test_expansion(128'h4272ec7700fda0669db28880ae2c5820, {16'd2938, 16'd36914, 16'd22189, 16'd39608, 16'd10696, 16'd10743, 16'd59584, 16'd15672, 16'd26793, 16'd7734, 16'd31644, 16'd56551, 16'd47024, 16'd21709, 16'd45338, 16'd9705, 16'd44279, 16'd46356, 16'd1829, 16'd51282, 16'd16731, 16'd26043, 16'd53708, 16'd46191, 16'd45989, 16'd38542});
	test_expansion(128'h00e61298baacdfdbdf6ac4f77eb56fdf, {16'd28696, 16'd13596, 16'd38795, 16'd25977, 16'd59837, 16'd37328, 16'd50165, 16'd12052, 16'd33107, 16'd19535, 16'd44880, 16'd64725, 16'd27322, 16'd44855, 16'd34876, 16'd34885, 16'd24145, 16'd54649, 16'd48387, 16'd29046, 16'd56484, 16'd22982, 16'd6137, 16'd31278, 16'd16552, 16'd38309});
	test_expansion(128'h08681717415b6491ca67a47b72a1eb5a, {16'd21759, 16'd38262, 16'd41990, 16'd27030, 16'd49031, 16'd13422, 16'd34734, 16'd10683, 16'd8917, 16'd17006, 16'd44922, 16'd25126, 16'd24367, 16'd9291, 16'd50314, 16'd7213, 16'd52964, 16'd49663, 16'd51439, 16'd16212, 16'd4476, 16'd25625, 16'd45584, 16'd57636, 16'd30044, 16'd58738});
	test_expansion(128'h1cae809f8f0ea64be98cfcdc01393f83, {16'd44165, 16'd35287, 16'd64420, 16'd22216, 16'd13938, 16'd11298, 16'd16401, 16'd61494, 16'd11012, 16'd64668, 16'd36778, 16'd23704, 16'd53096, 16'd20102, 16'd7753, 16'd444, 16'd23205, 16'd59440, 16'd9250, 16'd62524, 16'd56772, 16'd12584, 16'd64227, 16'd61650, 16'd31713, 16'd65479});
	test_expansion(128'he4a4968bb7668f69ef1fa75b2efea11e, {16'd324, 16'd4349, 16'd24505, 16'd421, 16'd57374, 16'd13148, 16'd26931, 16'd64590, 16'd61843, 16'd43555, 16'd15400, 16'd50653, 16'd59525, 16'd50081, 16'd15070, 16'd6554, 16'd65276, 16'd37505, 16'd47600, 16'd64220, 16'd51330, 16'd25805, 16'd4455, 16'd29564, 16'd36629, 16'd46461});
	test_expansion(128'ha00f9ec85f7ded3c9ed3a30fd827f03f, {16'd16807, 16'd8897, 16'd47147, 16'd32229, 16'd62187, 16'd62638, 16'd54188, 16'd1450, 16'd22786, 16'd23516, 16'd14554, 16'd13689, 16'd59479, 16'd23266, 16'd59660, 16'd32724, 16'd4271, 16'd59939, 16'd45526, 16'd38613, 16'd18597, 16'd57667, 16'd53164, 16'd4416, 16'd42091, 16'd2365});
	test_expansion(128'hedad5da9d0bb8b20da50817b7e41b9db, {16'd34241, 16'd12159, 16'd46225, 16'd47102, 16'd38850, 16'd51209, 16'd46728, 16'd46949, 16'd17604, 16'd23651, 16'd4201, 16'd52332, 16'd39017, 16'd56300, 16'd25994, 16'd905, 16'd9105, 16'd19264, 16'd3985, 16'd54970, 16'd3429, 16'd32864, 16'd54108, 16'd36937, 16'd64867, 16'd40210});
	test_expansion(128'hb5487b578bd1e341d83af300c0dfd1a7, {16'd22699, 16'd42501, 16'd5815, 16'd54529, 16'd56318, 16'd6466, 16'd42056, 16'd6389, 16'd25536, 16'd14663, 16'd63243, 16'd127, 16'd25953, 16'd52801, 16'd62218, 16'd26898, 16'd3427, 16'd38856, 16'd63172, 16'd35777, 16'd48896, 16'd8983, 16'd51648, 16'd27449, 16'd2871, 16'd22998});
	test_expansion(128'h3e01c3ab3086919de5cad85135ac8c38, {16'd53545, 16'd63163, 16'd15316, 16'd13575, 16'd39551, 16'd34447, 16'd14054, 16'd51770, 16'd22895, 16'd41047, 16'd8373, 16'd38540, 16'd42718, 16'd13109, 16'd33209, 16'd36308, 16'd50031, 16'd39238, 16'd26810, 16'd50138, 16'd6833, 16'd44397, 16'd2809, 16'd59079, 16'd21538, 16'd14604});
	test_expansion(128'hc01bc6dc7819f9781bbc0b98741d6bdd, {16'd10028, 16'd3845, 16'd12920, 16'd58948, 16'd65524, 16'd4221, 16'd45503, 16'd12127, 16'd38435, 16'd37075, 16'd13435, 16'd16180, 16'd55138, 16'd59607, 16'd1421, 16'd2048, 16'd8817, 16'd48603, 16'd61526, 16'd11216, 16'd55914, 16'd61731, 16'd34581, 16'd7948, 16'd26171, 16'd26007});
	test_expansion(128'h0a19fe48fc47c037ad4afae67faa38c5, {16'd21071, 16'd49290, 16'd21884, 16'd8945, 16'd16885, 16'd18204, 16'd19123, 16'd59728, 16'd47881, 16'd60503, 16'd2177, 16'd34708, 16'd21848, 16'd23230, 16'd37397, 16'd6592, 16'd14891, 16'd62926, 16'd33436, 16'd8425, 16'd25721, 16'd11067, 16'd10716, 16'd51908, 16'd58547, 16'd47098});
	test_expansion(128'hc1a2954c3b9991e3801a7a050c51a6f5, {16'd45345, 16'd16430, 16'd31563, 16'd48032, 16'd47665, 16'd34051, 16'd13715, 16'd38094, 16'd27383, 16'd32994, 16'd16528, 16'd18241, 16'd24128, 16'd24678, 16'd52404, 16'd5125, 16'd54329, 16'd15030, 16'd12910, 16'd62249, 16'd14880, 16'd40246, 16'd4190, 16'd37894, 16'd19324, 16'd32984});
	test_expansion(128'head68d9b5c6142cb213790c8c3b662cd, {16'd34348, 16'd28370, 16'd1839, 16'd37785, 16'd8756, 16'd4868, 16'd42618, 16'd59436, 16'd63266, 16'd27354, 16'd7406, 16'd26084, 16'd37560, 16'd18807, 16'd42746, 16'd46095, 16'd43680, 16'd33975, 16'd40372, 16'd25162, 16'd15891, 16'd34259, 16'd44747, 16'd10846, 16'd49387, 16'd3056});
	test_expansion(128'hf038bcc1a93fba0875f8f1e9542cd715, {16'd49094, 16'd26517, 16'd54269, 16'd31736, 16'd58521, 16'd60517, 16'd61148, 16'd4682, 16'd10654, 16'd6781, 16'd29703, 16'd39538, 16'd25547, 16'd31283, 16'd1336, 16'd46823, 16'd19765, 16'd63898, 16'd20661, 16'd58860, 16'd20568, 16'd13008, 16'd14773, 16'd6155, 16'd43023, 16'd11463});
	test_expansion(128'hd7af2a8e179a2acd8c4b71869dbbe807, {16'd41969, 16'd41452, 16'd20689, 16'd18800, 16'd44442, 16'd20678, 16'd15857, 16'd46501, 16'd53904, 16'd11412, 16'd30696, 16'd55417, 16'd35147, 16'd55483, 16'd10041, 16'd62520, 16'd5009, 16'd1359, 16'd19492, 16'd4338, 16'd25445, 16'd29997, 16'd52024, 16'd44243, 16'd37679, 16'd11780});
	test_expansion(128'h398b05f7d309b88ef77a74f6476e3570, {16'd21687, 16'd48756, 16'd2072, 16'd47383, 16'd20188, 16'd24811, 16'd50109, 16'd54601, 16'd42262, 16'd63049, 16'd53284, 16'd55000, 16'd8346, 16'd48704, 16'd5590, 16'd46874, 16'd20963, 16'd6731, 16'd55159, 16'd49907, 16'd3892, 16'd9113, 16'd29987, 16'd45795, 16'd39335, 16'd23249});
	test_expansion(128'hbb3025d2893c0b102a219927b242bb02, {16'd53902, 16'd16484, 16'd19155, 16'd14939, 16'd3664, 16'd41375, 16'd48475, 16'd52145, 16'd15145, 16'd12274, 16'd15823, 16'd18824, 16'd50225, 16'd60074, 16'd13178, 16'd43990, 16'd63713, 16'd36432, 16'd36555, 16'd30970, 16'd60392, 16'd28988, 16'd39955, 16'd8565, 16'd44942, 16'd51754});
	test_expansion(128'h37cbe4b135b4b6f213a4ba966006b34a, {16'd9949, 16'd33203, 16'd42678, 16'd64201, 16'd49247, 16'd28770, 16'd24632, 16'd59517, 16'd55076, 16'd39727, 16'd21612, 16'd37779, 16'd24615, 16'd62783, 16'd57189, 16'd61824, 16'd64979, 16'd24232, 16'd30496, 16'd13312, 16'd43804, 16'd34972, 16'd46100, 16'd48754, 16'd12738, 16'd50887});
	test_expansion(128'hec5e8ab86ab91cf268ad78e8b96b525a, {16'd34792, 16'd39888, 16'd62943, 16'd63206, 16'd59325, 16'd18321, 16'd22801, 16'd19517, 16'd3365, 16'd35610, 16'd10871, 16'd52517, 16'd64179, 16'd20173, 16'd21507, 16'd51410, 16'd55226, 16'd65056, 16'd11897, 16'd21187, 16'd47642, 16'd37726, 16'd8755, 16'd40141, 16'd36099, 16'd35435});
	test_expansion(128'hc7b1da24ff7e6733ec00fd0876591cda, {16'd31415, 16'd63063, 16'd57032, 16'd7044, 16'd15913, 16'd17708, 16'd54294, 16'd12448, 16'd23638, 16'd49616, 16'd51641, 16'd27097, 16'd34324, 16'd3943, 16'd9273, 16'd48365, 16'd49518, 16'd55410, 16'd45200, 16'd21445, 16'd50666, 16'd24982, 16'd7710, 16'd56408, 16'd58352, 16'd57312});
	test_expansion(128'hb716335ca35fc8364a625293d3cc781c, {16'd21555, 16'd14624, 16'd47721, 16'd57033, 16'd49544, 16'd29931, 16'd60904, 16'd41663, 16'd42058, 16'd27996, 16'd62034, 16'd65329, 16'd46322, 16'd4370, 16'd35671, 16'd44590, 16'd32938, 16'd39487, 16'd12916, 16'd58035, 16'd18472, 16'd52601, 16'd3497, 16'd51374, 16'd23107, 16'd7757});
	test_expansion(128'h67a994fa1c22454ed45014fb3c69d0eb, {16'd33903, 16'd16542, 16'd48115, 16'd64222, 16'd40265, 16'd28274, 16'd20619, 16'd14377, 16'd30289, 16'd20143, 16'd44178, 16'd17038, 16'd44601, 16'd14704, 16'd56853, 16'd63120, 16'd29538, 16'd56192, 16'd49964, 16'd46170, 16'd28660, 16'd36179, 16'd29635, 16'd43975, 16'd62098, 16'd42599});
	test_expansion(128'hd0d558730a30c9de1ecb514ecf94b5cb, {16'd40546, 16'd9517, 16'd61714, 16'd33540, 16'd50442, 16'd34123, 16'd33745, 16'd30667, 16'd55114, 16'd46062, 16'd51780, 16'd40209, 16'd22049, 16'd13391, 16'd39819, 16'd44841, 16'd58776, 16'd12555, 16'd48568, 16'd45, 16'd43395, 16'd46401, 16'd52772, 16'd58369, 16'd1336, 16'd4668});
	test_expansion(128'h4f3ff8fb3274f7a210bb8e9b59118972, {16'd56402, 16'd21844, 16'd14257, 16'd32519, 16'd48676, 16'd57442, 16'd56273, 16'd65174, 16'd27271, 16'd56553, 16'd35051, 16'd59238, 16'd3551, 16'd36291, 16'd10293, 16'd43750, 16'd50914, 16'd4456, 16'd12889, 16'd52471, 16'd1539, 16'd23508, 16'd10554, 16'd40061, 16'd32291, 16'd39161});
	test_expansion(128'h462d4b24873e9cd9ba508b69218386ca, {16'd364, 16'd34764, 16'd27082, 16'd11981, 16'd2688, 16'd57443, 16'd24085, 16'd10444, 16'd27934, 16'd55892, 16'd27297, 16'd48211, 16'd58205, 16'd8384, 16'd21821, 16'd31544, 16'd38746, 16'd10663, 16'd35501, 16'd16386, 16'd20032, 16'd36280, 16'd49561, 16'd37831, 16'd16163, 16'd47737});
	test_expansion(128'ha222171a738ffcdc1abe59cd425744df, {16'd1092, 16'd26035, 16'd33757, 16'd23220, 16'd28321, 16'd32807, 16'd59828, 16'd60572, 16'd50730, 16'd59581, 16'd61176, 16'd9275, 16'd51937, 16'd63441, 16'd17574, 16'd21598, 16'd11158, 16'd28696, 16'd14685, 16'd17459, 16'd16774, 16'd30924, 16'd20298, 16'd6025, 16'd49770, 16'd24764});
	test_expansion(128'h111ecc9b3d17caa16e1b39a965ec8965, {16'd7237, 16'd7408, 16'd17049, 16'd38313, 16'd31383, 16'd16546, 16'd39594, 16'd14602, 16'd42467, 16'd49215, 16'd26773, 16'd53138, 16'd34814, 16'd55826, 16'd10444, 16'd2863, 16'd40980, 16'd37278, 16'd44019, 16'd40545, 16'd23812, 16'd32679, 16'd62022, 16'd2988, 16'd21185, 16'd49643});
	test_expansion(128'hae47ecd618ad54e3e3250cdc08f8d148, {16'd17481, 16'd63313, 16'd10230, 16'd44456, 16'd4276, 16'd45388, 16'd37736, 16'd25889, 16'd34102, 16'd21457, 16'd8832, 16'd9910, 16'd8436, 16'd39758, 16'd11578, 16'd55677, 16'd15026, 16'd58955, 16'd60518, 16'd35920, 16'd44877, 16'd2509, 16'd19731, 16'd26906, 16'd1574, 16'd55325});
	test_expansion(128'h2405c08631d033519dc300cbbf094425, {16'd54662, 16'd27426, 16'd29811, 16'd32432, 16'd51445, 16'd50662, 16'd998, 16'd11845, 16'd2447, 16'd34283, 16'd24126, 16'd38649, 16'd42628, 16'd43858, 16'd3953, 16'd50353, 16'd24510, 16'd51316, 16'd58931, 16'd46866, 16'd57398, 16'd25372, 16'd53669, 16'd4395, 16'd41382, 16'd34713});
	test_expansion(128'hd8d65640f0873e4ff064c81ae2473215, {16'd61683, 16'd13485, 16'd50416, 16'd61804, 16'd5042, 16'd14400, 16'd19871, 16'd32487, 16'd30261, 16'd21742, 16'd63606, 16'd16791, 16'd43212, 16'd7120, 16'd52843, 16'd48928, 16'd16025, 16'd6978, 16'd4365, 16'd9404, 16'd30585, 16'd11483, 16'd19701, 16'd511, 16'd29709, 16'd25585});
	test_expansion(128'h31f522301bfef9a06623c13af9d655c0, {16'd55976, 16'd14638, 16'd55999, 16'd6416, 16'd49790, 16'd7514, 16'd2075, 16'd7068, 16'd11104, 16'd33911, 16'd8691, 16'd30283, 16'd8892, 16'd36650, 16'd5008, 16'd49296, 16'd54078, 16'd42798, 16'd20595, 16'd38966, 16'd35371, 16'd53603, 16'd46239, 16'd10336, 16'd22169, 16'd14211});
	test_expansion(128'h009a4c259b8772f5492107571d1a0d4c, {16'd18688, 16'd22529, 16'd1073, 16'd44038, 16'd30028, 16'd55761, 16'd62496, 16'd33213, 16'd803, 16'd33973, 16'd47988, 16'd38441, 16'd36336, 16'd33904, 16'd9150, 16'd63330, 16'd41495, 16'd37008, 16'd31716, 16'd37739, 16'd8934, 16'd32607, 16'd56954, 16'd54511, 16'd21585, 16'd42774});
	test_expansion(128'hd121a2e09156734ecda9ff61e29b7b87, {16'd59489, 16'd8582, 16'd2887, 16'd38707, 16'd16729, 16'd3977, 16'd13144, 16'd2947, 16'd26083, 16'd30214, 16'd6547, 16'd608, 16'd27737, 16'd16840, 16'd13834, 16'd44035, 16'd65203, 16'd17393, 16'd48297, 16'd20233, 16'd36728, 16'd33119, 16'd38246, 16'd14395, 16'd26877, 16'd14672});
	test_expansion(128'he4660f79fe502fdddc652a59cea83f0c, {16'd651, 16'd60062, 16'd16613, 16'd58540, 16'd10095, 16'd23277, 16'd32711, 16'd27327, 16'd64332, 16'd10646, 16'd65130, 16'd51942, 16'd53325, 16'd30250, 16'd23006, 16'd34236, 16'd56197, 16'd3483, 16'd19112, 16'd44035, 16'd54224, 16'd25345, 16'd46486, 16'd26654, 16'd36535, 16'd14890});
	test_expansion(128'h6e7252913b62758b408c63c741d6ef68, {16'd16003, 16'd14970, 16'd14069, 16'd9643, 16'd3609, 16'd33904, 16'd10133, 16'd5674, 16'd12731, 16'd55623, 16'd1787, 16'd15717, 16'd57173, 16'd44974, 16'd4791, 16'd17033, 16'd37326, 16'd2654, 16'd15174, 16'd12579, 16'd46839, 16'd17224, 16'd55710, 16'd22252, 16'd19009, 16'd39008});
	test_expansion(128'h7da270a8b6f6405af05e5555a81a4fac, {16'd20215, 16'd57907, 16'd20025, 16'd2517, 16'd42215, 16'd42626, 16'd60776, 16'd51090, 16'd43412, 16'd62555, 16'd38629, 16'd825, 16'd49784, 16'd39219, 16'd29124, 16'd61926, 16'd17879, 16'd36779, 16'd22627, 16'd25643, 16'd50106, 16'd42004, 16'd11060, 16'd187, 16'd27378, 16'd32927});
	test_expansion(128'hd2cc8359f045e5cb5b5e58833d099734, {16'd32568, 16'd51016, 16'd34978, 16'd61519, 16'd62151, 16'd36867, 16'd25127, 16'd56868, 16'd50906, 16'd28742, 16'd20717, 16'd30005, 16'd33517, 16'd3707, 16'd43445, 16'd34725, 16'd34106, 16'd16363, 16'd63630, 16'd25663, 16'd22447, 16'd18380, 16'd28236, 16'd49740, 16'd65031, 16'd21661});
	test_expansion(128'h87ae49e6d44f7834da88c5f55d6fb082, {16'd11940, 16'd50688, 16'd962, 16'd12371, 16'd18314, 16'd51937, 16'd29897, 16'd4001, 16'd5796, 16'd27805, 16'd28889, 16'd5094, 16'd36229, 16'd10459, 16'd29150, 16'd12699, 16'd62131, 16'd23940, 16'd33298, 16'd6741, 16'd20877, 16'd50397, 16'd63587, 16'd43701, 16'd41676, 16'd56708});
	test_expansion(128'hc1f33c2ee338a2f1443d9127a97cb9a9, {16'd800, 16'd40789, 16'd24644, 16'd3058, 16'd63850, 16'd9844, 16'd2837, 16'd59334, 16'd53607, 16'd9081, 16'd2012, 16'd44484, 16'd31338, 16'd31513, 16'd17398, 16'd7430, 16'd17999, 16'd24621, 16'd665, 16'd50751, 16'd51768, 16'd18422, 16'd14790, 16'd3638, 16'd29519, 16'd24829});
	test_expansion(128'h0de0f6220494a08dd489a9f0e5e86fc3, {16'd44212, 16'd8172, 16'd47736, 16'd5864, 16'd56241, 16'd42807, 16'd40487, 16'd31043, 16'd63520, 16'd57053, 16'd25987, 16'd57781, 16'd7605, 16'd37915, 16'd6512, 16'd3686, 16'd42009, 16'd39573, 16'd33863, 16'd46721, 16'd30118, 16'd23380, 16'd26798, 16'd36868, 16'd14568, 16'd44863});
	test_expansion(128'hb2a1d3e5752a6f3fb8e57b6c0e26effc, {16'd9574, 16'd39446, 16'd56879, 16'd34181, 16'd5664, 16'd3826, 16'd35580, 16'd329, 16'd12137, 16'd58993, 16'd30247, 16'd46019, 16'd7982, 16'd726, 16'd51950, 16'd38001, 16'd53396, 16'd58656, 16'd58962, 16'd27465, 16'd3330, 16'd45205, 16'd25253, 16'd49038, 16'd42525, 16'd11983});
	test_expansion(128'hf898acda8fd0b76bfec55aa77b058a02, {16'd64683, 16'd38804, 16'd16357, 16'd23638, 16'd41683, 16'd49705, 16'd15550, 16'd55681, 16'd13041, 16'd54576, 16'd30198, 16'd44999, 16'd65449, 16'd7398, 16'd39052, 16'd7863, 16'd23659, 16'd49785, 16'd45168, 16'd2227, 16'd51440, 16'd596, 16'd28907, 16'd52258, 16'd52641, 16'd15709});
	test_expansion(128'hd4b144a46db45ac0c008bf903f3ac445, {16'd25974, 16'd55386, 16'd60667, 16'd8887, 16'd2807, 16'd40630, 16'd24001, 16'd35211, 16'd39407, 16'd4058, 16'd13571, 16'd34431, 16'd10087, 16'd41543, 16'd37414, 16'd5625, 16'd3755, 16'd23084, 16'd5087, 16'd28573, 16'd47194, 16'd18287, 16'd47473, 16'd55971, 16'd14947, 16'd54782});
	test_expansion(128'h19af1e2e2518beb13f8456fec3ae16ce, {16'd28564, 16'd28618, 16'd17449, 16'd27364, 16'd53927, 16'd4732, 16'd39760, 16'd14885, 16'd13607, 16'd17494, 16'd8100, 16'd8962, 16'd19081, 16'd47620, 16'd41029, 16'd49946, 16'd28429, 16'd63373, 16'd1736, 16'd40587, 16'd52147, 16'd65479, 16'd27276, 16'd61, 16'd49896, 16'd19771});
	test_expansion(128'he2d3824fa89fb29e2053f121d522c85b, {16'd20035, 16'd31686, 16'd54779, 16'd31244, 16'd33021, 16'd9370, 16'd28018, 16'd39223, 16'd27717, 16'd51736, 16'd65311, 16'd11280, 16'd8377, 16'd64393, 16'd34422, 16'd40053, 16'd44100, 16'd23290, 16'd57762, 16'd15355, 16'd36444, 16'd59104, 16'd21000, 16'd20607, 16'd44218, 16'd24163});
	test_expansion(128'he5d5cc25631f7fd430a5cda07059958d, {16'd10460, 16'd41365, 16'd30071, 16'd44089, 16'd56876, 16'd41841, 16'd43905, 16'd341, 16'd37406, 16'd2739, 16'd34704, 16'd62645, 16'd60242, 16'd21153, 16'd64244, 16'd41901, 16'd28785, 16'd43098, 16'd35237, 16'd12601, 16'd19472, 16'd55514, 16'd12270, 16'd11848, 16'd2629, 16'd25882});
	test_expansion(128'h481796672a3fe4e4627009f41dcb5090, {16'd16740, 16'd3806, 16'd9528, 16'd32619, 16'd26490, 16'd51519, 16'd61128, 16'd58589, 16'd38561, 16'd21380, 16'd50515, 16'd27290, 16'd11108, 16'd40710, 16'd21470, 16'd25565, 16'd19824, 16'd28756, 16'd47051, 16'd20809, 16'd18226, 16'd48165, 16'd46061, 16'd56801, 16'd8495, 16'd52358});
	test_expansion(128'h7fe83425d9a05505cdd968bd2c58de36, {16'd37418, 16'd9344, 16'd39672, 16'd58086, 16'd59244, 16'd34048, 16'd41889, 16'd3509, 16'd20663, 16'd23648, 16'd56471, 16'd8721, 16'd31235, 16'd2354, 16'd64858, 16'd40318, 16'd59486, 16'd17026, 16'd62190, 16'd25537, 16'd54647, 16'd10414, 16'd25396, 16'd20327, 16'd24572, 16'd30399});
	test_expansion(128'ha4378908e19a3e446620af0329b1e515, {16'd16894, 16'd3315, 16'd54118, 16'd18041, 16'd5822, 16'd35391, 16'd46394, 16'd15431, 16'd43314, 16'd37406, 16'd39917, 16'd49184, 16'd43266, 16'd63149, 16'd16761, 16'd4806, 16'd58634, 16'd1097, 16'd32871, 16'd29484, 16'd45079, 16'd21531, 16'd27243, 16'd53190, 16'd6836, 16'd1730});
	test_expansion(128'hf1212ffeb746d5ce1a424ecac690e5e1, {16'd5255, 16'd41508, 16'd19751, 16'd4393, 16'd34610, 16'd39366, 16'd48915, 16'd11774, 16'd47259, 16'd5687, 16'd5156, 16'd15932, 16'd27638, 16'd38192, 16'd3331, 16'd21410, 16'd57613, 16'd7526, 16'd63933, 16'd3280, 16'd58708, 16'd65177, 16'd49813, 16'd10053, 16'd47397, 16'd58857});
	test_expansion(128'h06ab2b0258729bc64eccba719a6b7613, {16'd33950, 16'd29137, 16'd49589, 16'd49146, 16'd28255, 16'd20841, 16'd10752, 16'd60506, 16'd18054, 16'd23496, 16'd43209, 16'd58521, 16'd62404, 16'd63890, 16'd54773, 16'd343, 16'd7438, 16'd22497, 16'd28656, 16'd45068, 16'd56999, 16'd8652, 16'd6616, 16'd50594, 16'd34932, 16'd12541});
	test_expansion(128'h62268dcd9e5074759b595c7fe3935348, {16'd38260, 16'd38253, 16'd42090, 16'd9261, 16'd19436, 16'd157, 16'd23686, 16'd61881, 16'd35228, 16'd59411, 16'd47894, 16'd48628, 16'd2564, 16'd42921, 16'd7428, 16'd24287, 16'd57935, 16'd60902, 16'd13172, 16'd62786, 16'd2558, 16'd32346, 16'd43766, 16'd15392, 16'd7287, 16'd58333});
	test_expansion(128'hddcf6c8c4d990f8dbb4e6047f09288e2, {16'd55481, 16'd14345, 16'd55190, 16'd50898, 16'd40253, 16'd46373, 16'd8460, 16'd5291, 16'd50152, 16'd35888, 16'd9197, 16'd35898, 16'd32627, 16'd2940, 16'd27335, 16'd38285, 16'd54592, 16'd44825, 16'd57737, 16'd15569, 16'd36958, 16'd4523, 16'd4861, 16'd61734, 16'd19898, 16'd41453});
	test_expansion(128'h55bf51546a89b608ed317be1afdf8fdf, {16'd37371, 16'd32929, 16'd58067, 16'd64364, 16'd45280, 16'd21997, 16'd40348, 16'd30639, 16'd10297, 16'd59049, 16'd6707, 16'd41474, 16'd19840, 16'd56260, 16'd22867, 16'd44974, 16'd23305, 16'd16060, 16'd49340, 16'd38867, 16'd65240, 16'd31969, 16'd60437, 16'd56069, 16'd28886, 16'd1222});
	test_expansion(128'h7ee752e3ae03b277f218e4d558e76550, {16'd38779, 16'd54579, 16'd51057, 16'd63064, 16'd46117, 16'd22815, 16'd23688, 16'd7761, 16'd57730, 16'd63201, 16'd9405, 16'd16640, 16'd23248, 16'd61801, 16'd50069, 16'd28608, 16'd15363, 16'd26277, 16'd27639, 16'd55431, 16'd33074, 16'd49698, 16'd5880, 16'd11054, 16'd48450, 16'd11331});
	test_expansion(128'h8b6d488fae126d7c726474d15abf824f, {16'd57834, 16'd64853, 16'd8819, 16'd19140, 16'd12201, 16'd1147, 16'd42213, 16'd37708, 16'd34344, 16'd5790, 16'd33071, 16'd55047, 16'd40491, 16'd59904, 16'd27114, 16'd17021, 16'd51481, 16'd58357, 16'd46944, 16'd10247, 16'd51306, 16'd10648, 16'd48337, 16'd51960, 16'd33551, 16'd42221});
	test_expansion(128'h72221b4d5b0392c7a0c681078348208c, {16'd61483, 16'd6873, 16'd21229, 16'd14168, 16'd44926, 16'd37602, 16'd43202, 16'd55117, 16'd44594, 16'd27305, 16'd23416, 16'd45522, 16'd3293, 16'd6853, 16'd14494, 16'd44530, 16'd13767, 16'd59560, 16'd61253, 16'd60919, 16'd4376, 16'd46944, 16'd25374, 16'd56601, 16'd39054, 16'd4060});
	test_expansion(128'h65b44423e855fdc9f884ab945ae21eb6, {16'd44475, 16'd39321, 16'd20350, 16'd52374, 16'd4894, 16'd43559, 16'd39250, 16'd24353, 16'd18787, 16'd13337, 16'd15312, 16'd30546, 16'd5371, 16'd39001, 16'd27999, 16'd53658, 16'd7763, 16'd64793, 16'd86, 16'd6356, 16'd25456, 16'd40445, 16'd63824, 16'd33086, 16'd10725, 16'd28071});
	test_expansion(128'h3120acf678bb5b13f332d55ede761b41, {16'd44273, 16'd14468, 16'd46071, 16'd23324, 16'd46157, 16'd65496, 16'd53, 16'd62334, 16'd55046, 16'd11912, 16'd23788, 16'd35539, 16'd3399, 16'd27612, 16'd31720, 16'd35269, 16'd7470, 16'd30379, 16'd37236, 16'd31092, 16'd29246, 16'd5173, 16'd53479, 16'd36687, 16'd8091, 16'd6445});
	test_expansion(128'h60e6378fd3ac47818322facce1df0aca, {16'd40355, 16'd23633, 16'd27741, 16'd41446, 16'd53700, 16'd36470, 16'd57776, 16'd54658, 16'd6391, 16'd45151, 16'd42108, 16'd41875, 16'd27536, 16'd125, 16'd42343, 16'd39529, 16'd34554, 16'd41581, 16'd43677, 16'd31770, 16'd27180, 16'd795, 16'd41285, 16'd47155, 16'd53659, 16'd5026});
	test_expansion(128'h0501133288d539a7e8d914980b43963e, {16'd37768, 16'd20084, 16'd57091, 16'd14073, 16'd46124, 16'd796, 16'd48340, 16'd12230, 16'd46939, 16'd61617, 16'd18947, 16'd62064, 16'd1630, 16'd55595, 16'd60639, 16'd15724, 16'd3477, 16'd17780, 16'd26324, 16'd65191, 16'd18619, 16'd39060, 16'd36850, 16'd36274, 16'd10690, 16'd4878});
	test_expansion(128'h83dcdf4c1db657e326d1bbba4586cdf0, {16'd25833, 16'd47270, 16'd12321, 16'd13595, 16'd62126, 16'd36952, 16'd18536, 16'd28027, 16'd17978, 16'd26573, 16'd24387, 16'd54169, 16'd14165, 16'd37701, 16'd12999, 16'd34553, 16'd35262, 16'd32428, 16'd54861, 16'd7669, 16'd11285, 16'd31595, 16'd14956, 16'd28347, 16'd45333, 16'd45804});
	test_expansion(128'hf55da90d4164d2feaf36812b9fbdd87c, {16'd64525, 16'd55248, 16'd62505, 16'd2449, 16'd35185, 16'd29631, 16'd33898, 16'd915, 16'd54362, 16'd53519, 16'd28638, 16'd20086, 16'd35564, 16'd24008, 16'd6190, 16'd44749, 16'd21778, 16'd20731, 16'd55407, 16'd9066, 16'd55277, 16'd8205, 16'd27880, 16'd63535, 16'd30564, 16'd38782});
	test_expansion(128'heca00faa17d0644601622379859b2785, {16'd55737, 16'd7752, 16'd53271, 16'd3620, 16'd19000, 16'd36770, 16'd8355, 16'd23371, 16'd37998, 16'd8439, 16'd62110, 16'd49078, 16'd42826, 16'd18855, 16'd19762, 16'd60474, 16'd51995, 16'd31630, 16'd54088, 16'd14185, 16'd50461, 16'd57157, 16'd26626, 16'd32563, 16'd22806, 16'd61191});
	test_expansion(128'h9597de0701ba899c2e3a645d3b28d348, {16'd7151, 16'd58828, 16'd40649, 16'd50139, 16'd42518, 16'd14975, 16'd54111, 16'd63951, 16'd3850, 16'd22996, 16'd476, 16'd60252, 16'd1884, 16'd34489, 16'd52843, 16'd49507, 16'd31614, 16'd27489, 16'd51357, 16'd34084, 16'd47861, 16'd53874, 16'd33006, 16'd49967, 16'd2632, 16'd5247});
	test_expansion(128'hedee59bea4844a851485e47abd12806e, {16'd22482, 16'd1568, 16'd63498, 16'd60736, 16'd15207, 16'd45540, 16'd42152, 16'd22104, 16'd64857, 16'd2687, 16'd51641, 16'd11908, 16'd3292, 16'd37638, 16'd37852, 16'd39351, 16'd34613, 16'd39077, 16'd52712, 16'd43496, 16'd60630, 16'd19390, 16'd52628, 16'd22312, 16'd46014, 16'd49448});
	test_expansion(128'hc5640ac10a672c95ecf81943b4401ed4, {16'd47734, 16'd45277, 16'd50374, 16'd41201, 16'd15731, 16'd36394, 16'd45488, 16'd55172, 16'd59696, 16'd63665, 16'd22849, 16'd38899, 16'd48889, 16'd35664, 16'd37992, 16'd54966, 16'd7738, 16'd53631, 16'd42259, 16'd11351, 16'd25072, 16'd51842, 16'd55392, 16'd61039, 16'd60192, 16'd37060});
	test_expansion(128'h6c4b34a8c3d585f17441dc5a3ec84681, {16'd31301, 16'd50578, 16'd9661, 16'd39306, 16'd48048, 16'd28940, 16'd7224, 16'd61264, 16'd8752, 16'd20732, 16'd49269, 16'd16621, 16'd53847, 16'd7266, 16'd31228, 16'd51937, 16'd47344, 16'd58907, 16'd5186, 16'd19541, 16'd49729, 16'd6861, 16'd27195, 16'd24840, 16'd10858, 16'd21121});
	test_expansion(128'h422394d39398d45f45e023c2625ee6ef, {16'd35647, 16'd16402, 16'd57811, 16'd10972, 16'd55282, 16'd15719, 16'd9089, 16'd43562, 16'd43195, 16'd47770, 16'd62834, 16'd26723, 16'd40776, 16'd46207, 16'd4053, 16'd25047, 16'd18350, 16'd6331, 16'd64482, 16'd13204, 16'd36718, 16'd62311, 16'd13229, 16'd41184, 16'd6655, 16'd12164});
	test_expansion(128'he36c3f27c16195024cf3878ce855cdda, {16'd18393, 16'd35833, 16'd28968, 16'd33301, 16'd20464, 16'd15667, 16'd33249, 16'd21802, 16'd34611, 16'd34767, 16'd24766, 16'd59261, 16'd44093, 16'd52475, 16'd17467, 16'd40319, 16'd31019, 16'd11501, 16'd16185, 16'd17890, 16'd62287, 16'd51115, 16'd33288, 16'd8635, 16'd46554, 16'd59759});
	test_expansion(128'h608d2bf6cc79a4cf390e1f9af00e7497, {16'd64316, 16'd25903, 16'd44632, 16'd9538, 16'd3474, 16'd54802, 16'd38204, 16'd16935, 16'd55034, 16'd11552, 16'd52347, 16'd63766, 16'd20762, 16'd9236, 16'd16778, 16'd51965, 16'd63868, 16'd13621, 16'd643, 16'd22422, 16'd57228, 16'd44713, 16'd49001, 16'd33891, 16'd6052, 16'd9071});
	test_expansion(128'h52da9b1d142639391e42f597a5f8d2ef, {16'd24343, 16'd5643, 16'd17422, 16'd53502, 16'd1805, 16'd47404, 16'd34688, 16'd10428, 16'd45666, 16'd29885, 16'd51944, 16'd4617, 16'd59868, 16'd28775, 16'd43101, 16'd56241, 16'd17558, 16'd64667, 16'd23961, 16'd5738, 16'd3170, 16'd55605, 16'd8104, 16'd31314, 16'd32464, 16'd41673});
	test_expansion(128'h902184b52d746b7cc2c91b8302cf19ad, {16'd44059, 16'd55998, 16'd38717, 16'd7616, 16'd20334, 16'd46163, 16'd40743, 16'd45088, 16'd20707, 16'd35324, 16'd48046, 16'd34080, 16'd3232, 16'd47137, 16'd36640, 16'd5435, 16'd28014, 16'd59043, 16'd30688, 16'd28831, 16'd40265, 16'd34815, 16'd33511, 16'd54673, 16'd60491, 16'd16879});
	test_expansion(128'h5db0544ec157b1215f1597c63de68055, {16'd62840, 16'd40543, 16'd55101, 16'd55326, 16'd22029, 16'd1416, 16'd32007, 16'd12620, 16'd1001, 16'd25710, 16'd64986, 16'd54062, 16'd20924, 16'd5304, 16'd10328, 16'd27639, 16'd58224, 16'd36252, 16'd27152, 16'd64901, 16'd14432, 16'd38418, 16'd26082, 16'd6607, 16'd35447, 16'd31114});
	test_expansion(128'h3c3fae6feb63c4a183f173b4cff072ef, {16'd10234, 16'd21655, 16'd34777, 16'd64207, 16'd33260, 16'd30065, 16'd284, 16'd56981, 16'd41188, 16'd53029, 16'd32737, 16'd49240, 16'd10545, 16'd21271, 16'd27679, 16'd51210, 16'd31787, 16'd31771, 16'd43104, 16'd972, 16'd62910, 16'd59897, 16'd52965, 16'd60252, 16'd54903, 16'd44838});
	test_expansion(128'hd98fc5512fac2b31dfb91129b4a6e7d1, {16'd59948, 16'd50024, 16'd23807, 16'd46934, 16'd10043, 16'd63664, 16'd33693, 16'd34295, 16'd2794, 16'd43326, 16'd56714, 16'd45753, 16'd7289, 16'd61237, 16'd64541, 16'd29772, 16'd15180, 16'd16418, 16'd30232, 16'd65198, 16'd59043, 16'd26382, 16'd41826, 16'd18537, 16'd6026, 16'd60528});
	test_expansion(128'h05ba3c1c808d0e67077eb219fde30d2f, {16'd22220, 16'd57109, 16'd39952, 16'd46017, 16'd30978, 16'd7587, 16'd32948, 16'd36692, 16'd34849, 16'd39495, 16'd16366, 16'd52703, 16'd13504, 16'd56392, 16'd21135, 16'd4483, 16'd50611, 16'd55426, 16'd20002, 16'd20882, 16'd31831, 16'd43201, 16'd56346, 16'd41905, 16'd917, 16'd13393});
	test_expansion(128'he5b856e916d554a319dcf6baa1369915, {16'd7804, 16'd61688, 16'd31503, 16'd21173, 16'd34787, 16'd9802, 16'd9801, 16'd63391, 16'd42921, 16'd62159, 16'd3894, 16'd4942, 16'd34387, 16'd9236, 16'd46658, 16'd42603, 16'd51029, 16'd14510, 16'd2935, 16'd14131, 16'd43358, 16'd21273, 16'd11737, 16'd3782, 16'd63655, 16'd51594});
	test_expansion(128'h29a3173f0c3eaf52dd79910a1e301c86, {16'd16805, 16'd10091, 16'd15008, 16'd32166, 16'd16257, 16'd41405, 16'd17618, 16'd14657, 16'd39166, 16'd7580, 16'd12286, 16'd11220, 16'd19278, 16'd22209, 16'd63123, 16'd36096, 16'd44784, 16'd46630, 16'd6482, 16'd13017, 16'd56594, 16'd46267, 16'd16338, 16'd26164, 16'd12125, 16'd10019});
	test_expansion(128'h34e2e35e465572b96d7c4483eade6c8d, {16'd45815, 16'd40526, 16'd33916, 16'd61663, 16'd35016, 16'd64315, 16'd40071, 16'd9085, 16'd45849, 16'd28359, 16'd26707, 16'd51670, 16'd1119, 16'd8789, 16'd4514, 16'd8401, 16'd51544, 16'd28349, 16'd17690, 16'd44671, 16'd12318, 16'd29061, 16'd36531, 16'd50621, 16'd62045, 16'd5306});
	test_expansion(128'h88860ab1b340e3b26169dd6769b121d4, {16'd49163, 16'd5241, 16'd5896, 16'd53102, 16'd6282, 16'd41993, 16'd63211, 16'd49582, 16'd26904, 16'd52009, 16'd23791, 16'd60523, 16'd415, 16'd62884, 16'd61633, 16'd52014, 16'd21430, 16'd11976, 16'd16195, 16'd42193, 16'd6773, 16'd37673, 16'd11071, 16'd14399, 16'd49577, 16'd54005});
	test_expansion(128'heaaf62d141bd74e35204b98bce7a0893, {16'd31583, 16'd58697, 16'd50847, 16'd33685, 16'd41094, 16'd29701, 16'd13112, 16'd9692, 16'd64582, 16'd53593, 16'd4499, 16'd3312, 16'd29094, 16'd33465, 16'd14230, 16'd1677, 16'd4676, 16'd17442, 16'd14100, 16'd9049, 16'd17174, 16'd16645, 16'd49492, 16'd40952, 16'd47384, 16'd6468});
	test_expansion(128'h5e7875375d6e491246fb3514c5993b1f, {16'd32630, 16'd62259, 16'd16371, 16'd60286, 16'd35251, 16'd35224, 16'd3433, 16'd57005, 16'd42657, 16'd53885, 16'd46380, 16'd47847, 16'd4828, 16'd6076, 16'd8294, 16'd43007, 16'd62172, 16'd36867, 16'd36257, 16'd26392, 16'd48301, 16'd24861, 16'd46820, 16'd3080, 16'd51351, 16'd12397});
	test_expansion(128'h4c66899e7821aa51a7b36f1fdcc4809d, {16'd63769, 16'd3984, 16'd52109, 16'd18342, 16'd10168, 16'd19585, 16'd58775, 16'd23793, 16'd59999, 16'd61476, 16'd43200, 16'd13437, 16'd57250, 16'd51531, 16'd38682, 16'd42237, 16'd46060, 16'd52000, 16'd46286, 16'd20689, 16'd1499, 16'd60613, 16'd12029, 16'd8141, 16'd29373, 16'd33980});
	test_expansion(128'hd976567b45e71708d52b744c469c2949, {16'd22454, 16'd12503, 16'd33446, 16'd50187, 16'd21106, 16'd52857, 16'd35963, 16'd5207, 16'd39997, 16'd21340, 16'd44769, 16'd48426, 16'd12116, 16'd21750, 16'd11861, 16'd60278, 16'd5586, 16'd39450, 16'd8967, 16'd4801, 16'd18618, 16'd2891, 16'd26140, 16'd17650, 16'd60492, 16'd63113});
	test_expansion(128'h6dc26c7475ad018616e3563db432a97c, {16'd26320, 16'd28709, 16'd43034, 16'd49666, 16'd53294, 16'd44459, 16'd60301, 16'd10455, 16'd22975, 16'd3539, 16'd21760, 16'd53914, 16'd19956, 16'd12417, 16'd47401, 16'd14874, 16'd23793, 16'd21865, 16'd6376, 16'd16651, 16'd62018, 16'd60816, 16'd2942, 16'd16017, 16'd30504, 16'd64841});
	test_expansion(128'h76cd8930b8f9559164547e7c3db2d93f, {16'd5778, 16'd36767, 16'd46606, 16'd20426, 16'd40805, 16'd27677, 16'd62866, 16'd16418, 16'd26042, 16'd21406, 16'd17870, 16'd5380, 16'd47042, 16'd31843, 16'd65229, 16'd28120, 16'd1941, 16'd47144, 16'd31828, 16'd44923, 16'd25216, 16'd63694, 16'd22378, 16'd53563, 16'd28430, 16'd15869});
	test_expansion(128'h5de9e57d210eb3e54870ac62c69a2c6e, {16'd23013, 16'd5326, 16'd7626, 16'd43705, 16'd55788, 16'd65498, 16'd48981, 16'd4935, 16'd52280, 16'd25319, 16'd18899, 16'd45526, 16'd60418, 16'd32884, 16'd61299, 16'd8756, 16'd11502, 16'd8003, 16'd28526, 16'd28106, 16'd52538, 16'd2506, 16'd10038, 16'd23485, 16'd9409, 16'd30457});
	test_expansion(128'hcaaa8667c6eca9560640caa635af08ab, {16'd46359, 16'd51216, 16'd35004, 16'd64618, 16'd45449, 16'd18153, 16'd2843, 16'd35183, 16'd54428, 16'd29312, 16'd45253, 16'd8197, 16'd2007, 16'd45080, 16'd53996, 16'd8634, 16'd40691, 16'd3623, 16'd10471, 16'd55748, 16'd24677, 16'd46255, 16'd8957, 16'd63569, 16'd57450, 16'd20937});
	test_expansion(128'h37c7d5710cee32bbba0a3363279d3b8d, {16'd22862, 16'd24498, 16'd9105, 16'd52571, 16'd64149, 16'd17826, 16'd49928, 16'd8253, 16'd8704, 16'd14696, 16'd20675, 16'd21221, 16'd16971, 16'd51563, 16'd56796, 16'd217, 16'd25253, 16'd49294, 16'd24422, 16'd40709, 16'd5255, 16'd25281, 16'd7444, 16'd37705, 16'd50207, 16'd14737});
	test_expansion(128'h0dd0d1087ec833639864e4440bf6c6e6, {16'd14387, 16'd48514, 16'd64101, 16'd60090, 16'd6748, 16'd64060, 16'd55321, 16'd52130, 16'd2608, 16'd25854, 16'd36864, 16'd31230, 16'd3433, 16'd18058, 16'd46858, 16'd41905, 16'd52181, 16'd50295, 16'd37116, 16'd9111, 16'd22745, 16'd37562, 16'd37676, 16'd63610, 16'd3585, 16'd60944});
	test_expansion(128'h4a20dba1622f5bd9f44bbc141037cd7d, {16'd42843, 16'd47081, 16'd7634, 16'd33740, 16'd12753, 16'd28933, 16'd38868, 16'd48897, 16'd24519, 16'd41312, 16'd37787, 16'd4304, 16'd25982, 16'd52004, 16'd15329, 16'd16067, 16'd38419, 16'd26906, 16'd55463, 16'd56176, 16'd50030, 16'd54077, 16'd44497, 16'd45524, 16'd21706, 16'd12151});
	test_expansion(128'h3f31ea031d8145e35b441766455d5b76, {16'd34639, 16'd14914, 16'd8146, 16'd21268, 16'd38539, 16'd49752, 16'd61964, 16'd47865, 16'd520, 16'd5345, 16'd16162, 16'd60523, 16'd61937, 16'd62394, 16'd6876, 16'd37959, 16'd15818, 16'd55905, 16'd57370, 16'd58439, 16'd7050, 16'd47024, 16'd50336, 16'd13656, 16'd61272, 16'd54743});
	test_expansion(128'h86a9333e2941fd0a43f8a25978ea9b0f, {16'd36975, 16'd48898, 16'd47348, 16'd16734, 16'd58887, 16'd11374, 16'd8960, 16'd13554, 16'd56120, 16'd41487, 16'd64514, 16'd6360, 16'd50846, 16'd14359, 16'd733, 16'd16289, 16'd32255, 16'd49096, 16'd10310, 16'd62280, 16'd43828, 16'd44678, 16'd63282, 16'd59998, 16'd6592, 16'd49664});
	test_expansion(128'hd30339f9e938b6f152bca48c916ccacd, {16'd39097, 16'd10019, 16'd41106, 16'd33894, 16'd33822, 16'd6516, 16'd8320, 16'd51907, 16'd29770, 16'd27041, 16'd34474, 16'd11930, 16'd47753, 16'd62136, 16'd25275, 16'd38170, 16'd49291, 16'd34643, 16'd1262, 16'd20029, 16'd60933, 16'd11855, 16'd5050, 16'd44341, 16'd62487, 16'd9077});
	test_expansion(128'h2350d3dc1cb6cdcc43831fbcced4a191, {16'd4695, 16'd42768, 16'd32077, 16'd45079, 16'd17657, 16'd13493, 16'd15740, 16'd23184, 16'd62675, 16'd57009, 16'd53003, 16'd12633, 16'd64476, 16'd8463, 16'd17257, 16'd24327, 16'd17735, 16'd62267, 16'd23846, 16'd29232, 16'd43244, 16'd39964, 16'd64708, 16'd13290, 16'd36967, 16'd10174});
	test_expansion(128'h3089188c379c3076169293e251e3d746, {16'd28373, 16'd64028, 16'd59366, 16'd29685, 16'd61823, 16'd38893, 16'd50759, 16'd48677, 16'd5262, 16'd18180, 16'd10753, 16'd51838, 16'd40684, 16'd5913, 16'd65085, 16'd43889, 16'd56095, 16'd43679, 16'd61077, 16'd51774, 16'd14357, 16'd32954, 16'd41503, 16'd24167, 16'd21130, 16'd18644});
	test_expansion(128'hc1daee63e6470fea494d6058fd1b13cc, {16'd62070, 16'd47598, 16'd27708, 16'd50469, 16'd47519, 16'd34105, 16'd7882, 16'd37396, 16'd50098, 16'd59838, 16'd30384, 16'd47014, 16'd46962, 16'd45311, 16'd6943, 16'd59004, 16'd54040, 16'd59933, 16'd56766, 16'd51378, 16'd50275, 16'd32420, 16'd61930, 16'd14238, 16'd24401, 16'd1803});
	test_expansion(128'h91aa58ec7d70a88f594f7049aa6354a3, {16'd40224, 16'd9305, 16'd51576, 16'd41937, 16'd26212, 16'd65164, 16'd23070, 16'd60093, 16'd64152, 16'd29833, 16'd8289, 16'd19864, 16'd60314, 16'd38829, 16'd37872, 16'd44966, 16'd12229, 16'd26540, 16'd59566, 16'd23223, 16'd41719, 16'd40395, 16'd39623, 16'd32717, 16'd60871, 16'd11134});
	test_expansion(128'h94e65b543fac9c15012e156ffe36512a, {16'd61169, 16'd63558, 16'd24454, 16'd16321, 16'd52746, 16'd30750, 16'd27081, 16'd10315, 16'd47857, 16'd60524, 16'd33983, 16'd13701, 16'd14246, 16'd9393, 16'd43861, 16'd60736, 16'd13213, 16'd60299, 16'd41488, 16'd60653, 16'd60374, 16'd10577, 16'd26534, 16'd29006, 16'd12017, 16'd23342});
	test_expansion(128'hf54d6b81718d2fbd71741ba53588d10a, {16'd36020, 16'd24150, 16'd38698, 16'd2695, 16'd16265, 16'd31665, 16'd9120, 16'd13842, 16'd57863, 16'd11278, 16'd9159, 16'd9187, 16'd28161, 16'd8357, 16'd44368, 16'd25381, 16'd55118, 16'd36158, 16'd31434, 16'd41170, 16'd25797, 16'd55162, 16'd4874, 16'd303, 16'd50771, 16'd38120});
	test_expansion(128'h443af6e6b3f770408e9c327a5974c2cf, {16'd2466, 16'd21056, 16'd31203, 16'd12425, 16'd24520, 16'd51297, 16'd26047, 16'd12681, 16'd44375, 16'd44762, 16'd42868, 16'd15950, 16'd6947, 16'd60738, 16'd14767, 16'd34822, 16'd1123, 16'd13673, 16'd6089, 16'd56813, 16'd27516, 16'd7523, 16'd64129, 16'd60386, 16'd32880, 16'd33020});
	test_expansion(128'h2ea647d0d31096cab14472b7d61a9c32, {16'd63145, 16'd10546, 16'd29361, 16'd16219, 16'd28478, 16'd62456, 16'd41352, 16'd52266, 16'd16082, 16'd52145, 16'd51275, 16'd58725, 16'd38641, 16'd63338, 16'd46926, 16'd29819, 16'd45710, 16'd41239, 16'd33791, 16'd861, 16'd15219, 16'd15248, 16'd16919, 16'd16315, 16'd41333, 16'd16726});
	test_expansion(128'h6535fe3f576d20a196949ffb55967b5d, {16'd32202, 16'd44926, 16'd350, 16'd39514, 16'd27834, 16'd5507, 16'd20323, 16'd2378, 16'd65484, 16'd3730, 16'd2267, 16'd8605, 16'd14863, 16'd10354, 16'd39574, 16'd16920, 16'd52405, 16'd56084, 16'd22534, 16'd29616, 16'd53798, 16'd13725, 16'd25901, 16'd44950, 16'd34532, 16'd56762});
	test_expansion(128'hed3d6f7ea09419e08d5e04202cb733de, {16'd1457, 16'd48689, 16'd25121, 16'd47412, 16'd26537, 16'd57404, 16'd3106, 16'd34309, 16'd57424, 16'd20441, 16'd22071, 16'd8157, 16'd9583, 16'd47012, 16'd3548, 16'd33865, 16'd16974, 16'd56204, 16'd63109, 16'd41780, 16'd63953, 16'd46949, 16'd26659, 16'd27361, 16'd17479, 16'd47723});
	test_expansion(128'h3f30a5e75f530a40391bbbef9c97e083, {16'd3234, 16'd13580, 16'd58690, 16'd41794, 16'd35798, 16'd25946, 16'd20180, 16'd61193, 16'd11047, 16'd22102, 16'd64628, 16'd47582, 16'd22457, 16'd670, 16'd33707, 16'd4949, 16'd60484, 16'd8010, 16'd57951, 16'd6388, 16'd34958, 16'd52561, 16'd36356, 16'd22684, 16'd27962, 16'd65528});
	test_expansion(128'h31bdfba124cc934d2f689beb86256736, {16'd32000, 16'd17601, 16'd37238, 16'd43856, 16'd4729, 16'd42206, 16'd53759, 16'd6235, 16'd42176, 16'd31525, 16'd977, 16'd47352, 16'd29542, 16'd23024, 16'd58093, 16'd36594, 16'd29386, 16'd24481, 16'd65210, 16'd3351, 16'd37122, 16'd37134, 16'd28835, 16'd1903, 16'd65444, 16'd44378});
	test_expansion(128'h5285740eabde7361628881cf296952e4, {16'd50420, 16'd45069, 16'd53922, 16'd2874, 16'd47123, 16'd1379, 16'd56971, 16'd32183, 16'd19595, 16'd56282, 16'd44056, 16'd31622, 16'd49059, 16'd17098, 16'd11923, 16'd7653, 16'd31799, 16'd28993, 16'd43683, 16'd12642, 16'd35736, 16'd48938, 16'd1838, 16'd12621, 16'd42467, 16'd2279});
	test_expansion(128'h5f280801bdd712fa4693417e0f39ed23, {16'd39847, 16'd7091, 16'd57274, 16'd52682, 16'd47551, 16'd17541, 16'd34012, 16'd56515, 16'd63792, 16'd24811, 16'd53225, 16'd42208, 16'd14405, 16'd63109, 16'd18554, 16'd1528, 16'd54614, 16'd3759, 16'd18344, 16'd26060, 16'd62971, 16'd62010, 16'd46956, 16'd60544, 16'd42635, 16'd13314});
	test_expansion(128'h387c57b31a2ef556256c7921e71f8448, {16'd33295, 16'd41921, 16'd33941, 16'd19513, 16'd29075, 16'd54977, 16'd58114, 16'd58773, 16'd19241, 16'd62764, 16'd52271, 16'd42794, 16'd58444, 16'd38715, 16'd50790, 16'd24924, 16'd43563, 16'd6741, 16'd18221, 16'd42367, 16'd3206, 16'd10231, 16'd23385, 16'd1450, 16'd3543, 16'd46277});
	test_expansion(128'h311f3f719bb15e1562813c115f3466eb, {16'd11377, 16'd28887, 16'd53801, 16'd50264, 16'd21891, 16'd196, 16'd32784, 16'd56836, 16'd38481, 16'd33992, 16'd62551, 16'd32859, 16'd38473, 16'd37559, 16'd11085, 16'd31431, 16'd37093, 16'd61885, 16'd61420, 16'd10456, 16'd58268, 16'd36395, 16'd51559, 16'd24290, 16'd41888, 16'd1686});
	test_expansion(128'h52ff25f1acbf54169030daa7436bb79d, {16'd40331, 16'd2094, 16'd54296, 16'd9659, 16'd55293, 16'd16377, 16'd46162, 16'd53664, 16'd28683, 16'd45097, 16'd790, 16'd30468, 16'd11086, 16'd28599, 16'd5814, 16'd51402, 16'd61615, 16'd2683, 16'd53655, 16'd64099, 16'd21354, 16'd18022, 16'd10183, 16'd37991, 16'd28987, 16'd62233});
	test_expansion(128'h21f6ff42630ef5b6ae3db312d009c03c, {16'd32809, 16'd27793, 16'd6197, 16'd44909, 16'd36106, 16'd8257, 16'd7222, 16'd41216, 16'd11527, 16'd56187, 16'd33937, 16'd16011, 16'd51346, 16'd20225, 16'd48329, 16'd60457, 16'd23558, 16'd1476, 16'd27066, 16'd15760, 16'd61918, 16'd11507, 16'd24291, 16'd23244, 16'd49991, 16'd51036});
	test_expansion(128'haf70edd14f6d32eb1589a1427df61e2c, {16'd930, 16'd39549, 16'd44259, 16'd41735, 16'd4030, 16'd46226, 16'd18598, 16'd7100, 16'd2133, 16'd35251, 16'd48916, 16'd19486, 16'd51081, 16'd4005, 16'd49311, 16'd31831, 16'd38390, 16'd7155, 16'd51946, 16'd8938, 16'd60665, 16'd23532, 16'd14050, 16'd346, 16'd54915, 16'd35210});
	test_expansion(128'h2887e1f5959ba50bbf5bb1f5d1ae71f6, {16'd46107, 16'd31621, 16'd3658, 16'd30592, 16'd53966, 16'd50769, 16'd34339, 16'd55194, 16'd28338, 16'd60522, 16'd29892, 16'd49985, 16'd24177, 16'd3539, 16'd51002, 16'd8709, 16'd8824, 16'd38775, 16'd12051, 16'd17259, 16'd50553, 16'd38727, 16'd39727, 16'd59705, 16'd13526, 16'd38045});
	test_expansion(128'hbc91806c15d0deab181dad1672fd4c6b, {16'd55215, 16'd9690, 16'd55489, 16'd48164, 16'd19995, 16'd4763, 16'd35481, 16'd11408, 16'd8605, 16'd39397, 16'd35877, 16'd2790, 16'd9885, 16'd22224, 16'd6527, 16'd36638, 16'd23091, 16'd55216, 16'd13557, 16'd55153, 16'd6430, 16'd47217, 16'd31222, 16'd53744, 16'd49308, 16'd57128});
	test_expansion(128'hfc0e23ac420df1ac36e37f5bf8710052, {16'd14385, 16'd54311, 16'd50591, 16'd47735, 16'd10804, 16'd21064, 16'd21460, 16'd22898, 16'd24181, 16'd42481, 16'd42294, 16'd4879, 16'd48724, 16'd7532, 16'd35454, 16'd46354, 16'd61066, 16'd21902, 16'd56020, 16'd2097, 16'd8857, 16'd20170, 16'd64016, 16'd18160, 16'd10124, 16'd53696});
	test_expansion(128'hb5274d45b49ab61dce79d3def211d004, {16'd50575, 16'd20173, 16'd29163, 16'd23856, 16'd40431, 16'd3339, 16'd12613, 16'd12416, 16'd15110, 16'd56529, 16'd16896, 16'd28616, 16'd28233, 16'd44644, 16'd60258, 16'd14477, 16'd5696, 16'd37798, 16'd62594, 16'd8958, 16'd17285, 16'd18605, 16'd42924, 16'd13039, 16'd25133, 16'd11000});
	test_expansion(128'h15d02f643a9b6ddfe3263755dae7914b, {16'd32352, 16'd14183, 16'd40406, 16'd46982, 16'd29430, 16'd10840, 16'd63174, 16'd22783, 16'd64489, 16'd15001, 16'd41389, 16'd12817, 16'd36095, 16'd38404, 16'd33997, 16'd64802, 16'd24401, 16'd56559, 16'd5423, 16'd57738, 16'd19232, 16'd52860, 16'd57482, 16'd23146, 16'd29566, 16'd44725});
	test_expansion(128'h5f46c8dcb2e6ccf657d910e759e375a6, {16'd23363, 16'd21236, 16'd27732, 16'd56851, 16'd8715, 16'd29844, 16'd23080, 16'd26732, 16'd53045, 16'd14052, 16'd11748, 16'd16058, 16'd28835, 16'd13031, 16'd63080, 16'd58261, 16'd5770, 16'd227, 16'd41536, 16'd48303, 16'd20215, 16'd7822, 16'd7784, 16'd1402, 16'd53261, 16'd37068});
	test_expansion(128'he9387e32eb4b2ab1628e8e7bb3edde5b, {16'd22353, 16'd53593, 16'd43826, 16'd54073, 16'd47266, 16'd31728, 16'd38138, 16'd7854, 16'd14127, 16'd33163, 16'd63659, 16'd30231, 16'd12619, 16'd60010, 16'd14614, 16'd41727, 16'd23009, 16'd26178, 16'd53383, 16'd48037, 16'd26742, 16'd170, 16'd38760, 16'd13686, 16'd46542, 16'd56108});
	test_expansion(128'hcf02f20d3e492510d4a3c30566b8a905, {16'd28060, 16'd3835, 16'd16308, 16'd26679, 16'd2003, 16'd42727, 16'd31637, 16'd38935, 16'd7879, 16'd18754, 16'd13398, 16'd15207, 16'd9784, 16'd41683, 16'd11787, 16'd5947, 16'd30369, 16'd544, 16'd50052, 16'd22408, 16'd60923, 16'd54190, 16'd51906, 16'd20156, 16'd30998, 16'd5472});
	test_expansion(128'hf2a6434eb2888fd7d3c2c284a23e673d, {16'd2155, 16'd44551, 16'd13198, 16'd25920, 16'd42947, 16'd10990, 16'd64312, 16'd56980, 16'd1192, 16'd49221, 16'd27706, 16'd53730, 16'd1200, 16'd33390, 16'd27442, 16'd12482, 16'd5469, 16'd3675, 16'd62937, 16'd60522, 16'd50397, 16'd5518, 16'd35621, 16'd57416, 16'd60593, 16'd6550});
	test_expansion(128'hc5a24da0835ca0ce108e8785cbde3ceb, {16'd2108, 16'd50291, 16'd11891, 16'd6525, 16'd65366, 16'd24927, 16'd42303, 16'd45649, 16'd7353, 16'd64046, 16'd15695, 16'd53142, 16'd54974, 16'd45022, 16'd5855, 16'd11317, 16'd33247, 16'd19507, 16'd6578, 16'd55253, 16'd35836, 16'd394, 16'd54837, 16'd51909, 16'd46797, 16'd50379});
	test_expansion(128'h30512ea4e040f9cb8957a8c21d06ac04, {16'd62589, 16'd9293, 16'd47496, 16'd39646, 16'd26729, 16'd43594, 16'd32940, 16'd60390, 16'd53395, 16'd41340, 16'd44276, 16'd33893, 16'd4628, 16'd33605, 16'd2346, 16'd329, 16'd45960, 16'd46378, 16'd48045, 16'd30842, 16'd58421, 16'd25527, 16'd17654, 16'd2523, 16'd20990, 16'd23612});
	test_expansion(128'h81ce816374482319de0ffcf4cf22519d, {16'd40723, 16'd60404, 16'd59866, 16'd47123, 16'd43587, 16'd18489, 16'd38018, 16'd12875, 16'd54327, 16'd56748, 16'd16109, 16'd2181, 16'd1520, 16'd8282, 16'd45261, 16'd42664, 16'd23979, 16'd21709, 16'd59321, 16'd49331, 16'd26664, 16'd36176, 16'd60382, 16'd37086, 16'd37868, 16'd52317});
	test_expansion(128'hdb6df96eefa7359ab8e8cc4c2a2678e8, {16'd9691, 16'd32193, 16'd49980, 16'd4453, 16'd41809, 16'd57260, 16'd11416, 16'd18662, 16'd42081, 16'd63063, 16'd39636, 16'd3092, 16'd23729, 16'd10863, 16'd36215, 16'd39565, 16'd33609, 16'd23916, 16'd7856, 16'd50400, 16'd7000, 16'd11450, 16'd54462, 16'd44857, 16'd44915, 16'd49878});
	test_expansion(128'h6fe0b411db96304b4731d570e9b46083, {16'd219, 16'd8284, 16'd46527, 16'd9493, 16'd26544, 16'd30612, 16'd5163, 16'd58902, 16'd43767, 16'd57770, 16'd6666, 16'd52642, 16'd5402, 16'd49846, 16'd63620, 16'd52014, 16'd48131, 16'd48197, 16'd54865, 16'd25711, 16'd47857, 16'd63451, 16'd62217, 16'd39717, 16'd62790, 16'd21464});
	test_expansion(128'h41baa9540061beac79c63b3ec4c5a1a2, {16'd56490, 16'd32841, 16'd28568, 16'd56223, 16'd27071, 16'd13017, 16'd1860, 16'd16375, 16'd8109, 16'd16341, 16'd35756, 16'd46170, 16'd36905, 16'd49948, 16'd23420, 16'd39367, 16'd60745, 16'd55062, 16'd62784, 16'd52181, 16'd32674, 16'd59885, 16'd47340, 16'd41609, 16'd35838, 16'd48098});
	test_expansion(128'hd7353ebc55223782c714ce7bb3a69f55, {16'd19669, 16'd5360, 16'd33961, 16'd45009, 16'd63790, 16'd53059, 16'd21884, 16'd54040, 16'd19973, 16'd32105, 16'd22716, 16'd43531, 16'd41049, 16'd28813, 16'd28605, 16'd18382, 16'd13475, 16'd21125, 16'd47852, 16'd23577, 16'd29645, 16'd28329, 16'd22286, 16'd51081, 16'd11171, 16'd17011});
	test_expansion(128'hc4fb74d8fdc9b5e5c7fce743d2855177, {16'd46341, 16'd25285, 16'd44699, 16'd19580, 16'd21561, 16'd3289, 16'd7144, 16'd19125, 16'd19623, 16'd59257, 16'd61560, 16'd57128, 16'd39916, 16'd59650, 16'd37955, 16'd61322, 16'd10513, 16'd50906, 16'd944, 16'd38154, 16'd20387, 16'd35699, 16'd60976, 16'd41128, 16'd41561, 16'd20437});
	test_expansion(128'h90e5f3b292d010aebd894d6beef2a353, {16'd21948, 16'd45985, 16'd42857, 16'd54282, 16'd34996, 16'd12270, 16'd56923, 16'd18426, 16'd65345, 16'd62945, 16'd35761, 16'd53455, 16'd41982, 16'd60046, 16'd56009, 16'd61271, 16'd29077, 16'd35162, 16'd65117, 16'd36559, 16'd28171, 16'd28267, 16'd32630, 16'd36223, 16'd39931, 16'd27657});
	test_expansion(128'hfbc1a6f8123e585162ced60e7d60653e, {16'd11650, 16'd645, 16'd32835, 16'd3932, 16'd15367, 16'd11205, 16'd3828, 16'd196, 16'd32215, 16'd14084, 16'd25375, 16'd1726, 16'd35782, 16'd51044, 16'd24618, 16'd27856, 16'd38532, 16'd57522, 16'd37383, 16'd24652, 16'd4784, 16'd32288, 16'd33750, 16'd4435, 16'd160, 16'd44369});
	test_expansion(128'he525d6b953071b65563f8a522a5b299d, {16'd12026, 16'd696, 16'd16947, 16'd50492, 16'd14450, 16'd47482, 16'd61903, 16'd11535, 16'd47730, 16'd42262, 16'd59984, 16'd54888, 16'd20971, 16'd32055, 16'd2352, 16'd15718, 16'd1778, 16'd54843, 16'd56481, 16'd12926, 16'd50315, 16'd37467, 16'd56759, 16'd34121, 16'd57606, 16'd21520});
	test_expansion(128'hc39eae35edeb5de8f81d018c068c4820, {16'd9527, 16'd9086, 16'd16371, 16'd21045, 16'd11627, 16'd42743, 16'd27726, 16'd43082, 16'd37613, 16'd40166, 16'd58610, 16'd64794, 16'd50340, 16'd5254, 16'd61984, 16'd56623, 16'd26700, 16'd59069, 16'd55871, 16'd30363, 16'd7881, 16'd27888, 16'd30714, 16'd27730, 16'd27176, 16'd43406});
	test_expansion(128'h8eba6c0860958ee75d65defb4b69e32e, {16'd15990, 16'd37093, 16'd23963, 16'd5957, 16'd34701, 16'd11238, 16'd57731, 16'd42675, 16'd30631, 16'd21774, 16'd63384, 16'd50415, 16'd43173, 16'd6626, 16'd22007, 16'd15962, 16'd25513, 16'd36957, 16'd23215, 16'd27845, 16'd34810, 16'd48584, 16'd19303, 16'd55008, 16'd38142, 16'd57681});
	test_expansion(128'h02020016126338ef438de49c8a1e7bf1, {16'd59071, 16'd37307, 16'd14900, 16'd24804, 16'd3719, 16'd16652, 16'd37120, 16'd20943, 16'd54867, 16'd53942, 16'd50318, 16'd49349, 16'd8365, 16'd409, 16'd62989, 16'd52810, 16'd4538, 16'd54912, 16'd20724, 16'd56075, 16'd51746, 16'd16420, 16'd32639, 16'd48184, 16'd11645, 16'd43140});
	test_expansion(128'h2c29e6a3d0fe4d5ed5e59862d7cb3cbe, {16'd4529, 16'd44945, 16'd28786, 16'd23362, 16'd9201, 16'd35050, 16'd50422, 16'd62141, 16'd25798, 16'd7379, 16'd5530, 16'd44091, 16'd24550, 16'd22478, 16'd46578, 16'd5315, 16'd22006, 16'd35312, 16'd10561, 16'd25211, 16'd23184, 16'd27572, 16'd45109, 16'd19505, 16'd56106, 16'd54952});
	test_expansion(128'hc8799760bdf5116946d9805f4dfb0899, {16'd49969, 16'd6187, 16'd15332, 16'd16382, 16'd61734, 16'd18739, 16'd23566, 16'd13733, 16'd31740, 16'd14457, 16'd424, 16'd7459, 16'd19289, 16'd2307, 16'd55675, 16'd12877, 16'd46867, 16'd48660, 16'd60452, 16'd16788, 16'd24397, 16'd59971, 16'd63815, 16'd7462, 16'd45419, 16'd39032});
	test_expansion(128'hc4ddf6bc600cc78088a4348cb59812a8, {16'd49567, 16'd14677, 16'd40697, 16'd2224, 16'd12300, 16'd61368, 16'd36103, 16'd58490, 16'd15635, 16'd63859, 16'd24483, 16'd2783, 16'd55181, 16'd9541, 16'd12427, 16'd20204, 16'd28691, 16'd32058, 16'd53644, 16'd14602, 16'd25074, 16'd22420, 16'd44691, 16'd61876, 16'd29309, 16'd22207});
	test_expansion(128'hb765f58cf9130c7865449073deba89f0, {16'd28229, 16'd24801, 16'd52556, 16'd4320, 16'd39159, 16'd33782, 16'd42269, 16'd3791, 16'd19686, 16'd738, 16'd40214, 16'd26104, 16'd60036, 16'd9674, 16'd20256, 16'd14092, 16'd63536, 16'd34749, 16'd61639, 16'd61657, 16'd25086, 16'd49078, 16'd7806, 16'd30545, 16'd10821, 16'd48706});
	test_expansion(128'hf2a4852d07bb77a7034194fd0b281a47, {16'd18617, 16'd560, 16'd27604, 16'd55285, 16'd31398, 16'd25362, 16'd59695, 16'd31971, 16'd15217, 16'd20176, 16'd39759, 16'd34787, 16'd23807, 16'd55458, 16'd29391, 16'd60037, 16'd9696, 16'd17742, 16'd49395, 16'd41521, 16'd27552, 16'd1714, 16'd11472, 16'd44779, 16'd55637, 16'd41081});
	test_expansion(128'hb0fc19d41f91c19f07a0e0ca561d76d6, {16'd60411, 16'd28985, 16'd61134, 16'd61065, 16'd50841, 16'd16360, 16'd17220, 16'd43604, 16'd39612, 16'd54017, 16'd58666, 16'd5297, 16'd47623, 16'd38729, 16'd18034, 16'd5, 16'd40895, 16'd44708, 16'd34108, 16'd11194, 16'd16651, 16'd19831, 16'd12030, 16'd61400, 16'd20497, 16'd33373});
	test_expansion(128'h815aa4dd1c90d24e2a9728c731404226, {16'd62546, 16'd25362, 16'd65528, 16'd31431, 16'd47424, 16'd48654, 16'd18829, 16'd39476, 16'd44341, 16'd35210, 16'd47611, 16'd50481, 16'd35066, 16'd32181, 16'd28662, 16'd40464, 16'd9838, 16'd7141, 16'd31003, 16'd25136, 16'd57084, 16'd51252, 16'd23239, 16'd23429, 16'd28478, 16'd64614});
	test_expansion(128'hdba2e107c965a6e958741190d65db78d, {16'd30585, 16'd24184, 16'd12896, 16'd54374, 16'd17650, 16'd13234, 16'd19876, 16'd37697, 16'd64831, 16'd59455, 16'd29964, 16'd13074, 16'd13904, 16'd47345, 16'd52084, 16'd4684, 16'd51296, 16'd12266, 16'd38145, 16'd30132, 16'd41973, 16'd45206, 16'd58545, 16'd7863, 16'd8364, 16'd8996});
	test_expansion(128'h966dceb6379fc97929f3b7489bd45418, {16'd57634, 16'd62405, 16'd22699, 16'd13607, 16'd14360, 16'd42893, 16'd15969, 16'd12907, 16'd15343, 16'd25856, 16'd11555, 16'd4480, 16'd23312, 16'd20022, 16'd10925, 16'd15094, 16'd51998, 16'd19795, 16'd20551, 16'd13593, 16'd33125, 16'd22963, 16'd4915, 16'd22131, 16'd32983, 16'd61971});
	test_expansion(128'h9d6b3d0680c7017c5abd737959aefd9c, {16'd3541, 16'd62440, 16'd64146, 16'd46321, 16'd29365, 16'd16137, 16'd15492, 16'd46518, 16'd64325, 16'd18268, 16'd56247, 16'd8690, 16'd9955, 16'd20615, 16'd58281, 16'd6535, 16'd36346, 16'd11963, 16'd39370, 16'd62105, 16'd59055, 16'd45448, 16'd51407, 16'd37682, 16'd13168, 16'd5486});
	test_expansion(128'h9d4af0a06261e72cc70cff7808d69fd7, {16'd7998, 16'd39764, 16'd41904, 16'd38716, 16'd15410, 16'd52411, 16'd44757, 16'd25110, 16'd18129, 16'd54770, 16'd48945, 16'd59674, 16'd20368, 16'd56133, 16'd10503, 16'd60197, 16'd36588, 16'd1040, 16'd9652, 16'd52556, 16'd5211, 16'd12640, 16'd59377, 16'd55914, 16'd9529, 16'd29430});
	test_expansion(128'h0b151eed56eace1bef26eef4f728490b, {16'd944, 16'd16879, 16'd61549, 16'd60137, 16'd32489, 16'd39007, 16'd63795, 16'd21843, 16'd62840, 16'd24912, 16'd23353, 16'd59970, 16'd31208, 16'd4227, 16'd51616, 16'd43184, 16'd60094, 16'd5496, 16'd45603, 16'd47321, 16'd5906, 16'd5205, 16'd49798, 16'd53310, 16'd44429, 16'd56421});
	test_expansion(128'hedcbf7b1145c04881e6a0b0b2b9ba407, {16'd62228, 16'd51531, 16'd41122, 16'd23795, 16'd59135, 16'd57314, 16'd9747, 16'd17018, 16'd11611, 16'd45453, 16'd31916, 16'd30734, 16'd33107, 16'd43480, 16'd38757, 16'd17816, 16'd18522, 16'd4248, 16'd64303, 16'd30420, 16'd51936, 16'd28076, 16'd1451, 16'd15391, 16'd17901, 16'd51061});
	test_expansion(128'h54897493e88e618d3c0c303b7b4ce49f, {16'd40212, 16'd43340, 16'd57377, 16'd6009, 16'd28742, 16'd18543, 16'd64855, 16'd39219, 16'd63888, 16'd9867, 16'd3822, 16'd48009, 16'd34313, 16'd64794, 16'd6156, 16'd43998, 16'd37415, 16'd13644, 16'd19746, 16'd16160, 16'd56476, 16'd60221, 16'd41272, 16'd15520, 16'd16884, 16'd42144});
	test_expansion(128'h08653c6a1c8206eab5dd0c3197aad005, {16'd36443, 16'd1496, 16'd21766, 16'd45896, 16'd27719, 16'd52029, 16'd15619, 16'd55873, 16'd28408, 16'd2998, 16'd54838, 16'd61011, 16'd8359, 16'd21404, 16'd4989, 16'd9322, 16'd21867, 16'd8298, 16'd58711, 16'd25812, 16'd64363, 16'd58944, 16'd32433, 16'd63185, 16'd52597, 16'd58367});
	test_expansion(128'h28d5585e6bf7d90288ba252622bac74e, {16'd16237, 16'd1280, 16'd31183, 16'd48150, 16'd64314, 16'd62809, 16'd62155, 16'd10850, 16'd48843, 16'd15455, 16'd9584, 16'd57650, 16'd48869, 16'd3645, 16'd58233, 16'd59001, 16'd64947, 16'd35877, 16'd40775, 16'd48961, 16'd51428, 16'd51354, 16'd15220, 16'd23962, 16'd5339, 16'd3718});
	test_expansion(128'h3fe33ee3a8a068becf18ebee796fae68, {16'd13815, 16'd31910, 16'd19495, 16'd46440, 16'd29502, 16'd59602, 16'd56178, 16'd28137, 16'd20392, 16'd44016, 16'd37785, 16'd44140, 16'd19185, 16'd31195, 16'd17063, 16'd36533, 16'd63731, 16'd38668, 16'd48496, 16'd59774, 16'd59804, 16'd61664, 16'd57169, 16'd37189, 16'd15357, 16'd52398});
	test_expansion(128'hcbbc9092e514d88c7789d8917a5215f1, {16'd9113, 16'd4988, 16'd13986, 16'd8714, 16'd41679, 16'd28948, 16'd47306, 16'd41431, 16'd6756, 16'd12828, 16'd31045, 16'd19516, 16'd55293, 16'd26533, 16'd31885, 16'd29991, 16'd27621, 16'd35550, 16'd59260, 16'd63329, 16'd12799, 16'd43182, 16'd62438, 16'd30074, 16'd52708, 16'd12218});
	test_expansion(128'h3bdb7d438e37f73285ba1e09bc28e17a, {16'd11356, 16'd53928, 16'd2354, 16'd57861, 16'd58633, 16'd19022, 16'd44315, 16'd36383, 16'd8600, 16'd57073, 16'd25357, 16'd47625, 16'd46573, 16'd43579, 16'd4757, 16'd13291, 16'd22892, 16'd34117, 16'd6280, 16'd15531, 16'd24343, 16'd62706, 16'd37324, 16'd16625, 16'd8960, 16'd23857});
	test_expansion(128'h3e7b142a3a263038bb77468ebea9e639, {16'd9409, 16'd11818, 16'd46132, 16'd25202, 16'd40843, 16'd35457, 16'd39942, 16'd55327, 16'd17973, 16'd53099, 16'd39379, 16'd28703, 16'd47182, 16'd12797, 16'd28687, 16'd51101, 16'd52572, 16'd35224, 16'd50381, 16'd16460, 16'd703, 16'd4172, 16'd18227, 16'd59446, 16'd54788, 16'd40178});
	test_expansion(128'h1bc70ffed04c6216b6225ab29a93aa09, {16'd2458, 16'd45667, 16'd55733, 16'd54318, 16'd62332, 16'd23777, 16'd21400, 16'd33973, 16'd27522, 16'd7355, 16'd64411, 16'd34234, 16'd7105, 16'd34437, 16'd4496, 16'd25601, 16'd44318, 16'd6245, 16'd61596, 16'd29865, 16'd62767, 16'd47151, 16'd11634, 16'd4834, 16'd31973, 16'd63969});
	test_expansion(128'hd95100913d3bf0f8968acdc5f58a7f21, {16'd46740, 16'd22124, 16'd57763, 16'd11163, 16'd45155, 16'd38814, 16'd43578, 16'd25834, 16'd9769, 16'd21464, 16'd60381, 16'd59342, 16'd29454, 16'd4028, 16'd10149, 16'd11064, 16'd58771, 16'd10268, 16'd1807, 16'd1530, 16'd15369, 16'd23112, 16'd54066, 16'd50944, 16'd23368, 16'd15047});
	test_expansion(128'hc9633a0b043d188b8f5b7f11e8fa6e26, {16'd11796, 16'd46063, 16'd20109, 16'd1121, 16'd35535, 16'd57575, 16'd62931, 16'd52310, 16'd31618, 16'd18715, 16'd27645, 16'd42653, 16'd12317, 16'd26107, 16'd16460, 16'd52642, 16'd53142, 16'd55726, 16'd59186, 16'd47842, 16'd49167, 16'd36373, 16'd40643, 16'd7236, 16'd49451, 16'd2498});
	test_expansion(128'h06083b916d1708f2b06cc2285696525b, {16'd27239, 16'd7283, 16'd62738, 16'd25751, 16'd60746, 16'd55112, 16'd1741, 16'd64220, 16'd62232, 16'd54959, 16'd16263, 16'd52778, 16'd40928, 16'd62805, 16'd5476, 16'd41816, 16'd37799, 16'd49607, 16'd13269, 16'd31930, 16'd45989, 16'd51374, 16'd20217, 16'd32315, 16'd28428, 16'd11726});
	test_expansion(128'hab222ddf7d06ac8bbd8a0e311548aaab, {16'd33512, 16'd27445, 16'd54207, 16'd13312, 16'd15998, 16'd60434, 16'd64084, 16'd39484, 16'd19665, 16'd33646, 16'd57631, 16'd49082, 16'd1326, 16'd29134, 16'd5550, 16'd33511, 16'd7187, 16'd62924, 16'd21086, 16'd1217, 16'd50115, 16'd41170, 16'd40628, 16'd62057, 16'd34548, 16'd29050});
	test_expansion(128'h29703cd06d7b8493eef5a8ec19e19833, {16'd53872, 16'd39530, 16'd61504, 16'd14055, 16'd4268, 16'd38838, 16'd61326, 16'd58369, 16'd22646, 16'd19378, 16'd41619, 16'd16439, 16'd2562, 16'd14125, 16'd6150, 16'd36790, 16'd10582, 16'd16520, 16'd31153, 16'd52901, 16'd18942, 16'd58988, 16'd19961, 16'd27139, 16'd4064, 16'd29568});
	test_expansion(128'ha5127e342867036d310c2f23b33e3aa4, {16'd14993, 16'd44711, 16'd3837, 16'd11620, 16'd49756, 16'd20908, 16'd52244, 16'd2162, 16'd37250, 16'd60085, 16'd14611, 16'd63091, 16'd65531, 16'd58330, 16'd28947, 16'd27144, 16'd49292, 16'd31156, 16'd30853, 16'd33687, 16'd28295, 16'd8330, 16'd58966, 16'd46311, 16'd30307, 16'd23275});
	test_expansion(128'hc4e1940b83122856c700b7c1585a74b2, {16'd31936, 16'd40758, 16'd11380, 16'd65411, 16'd49865, 16'd49165, 16'd52266, 16'd63518, 16'd40919, 16'd57173, 16'd39894, 16'd43668, 16'd11208, 16'd17418, 16'd14162, 16'd13562, 16'd30011, 16'd38801, 16'd2854, 16'd30757, 16'd41060, 16'd14509, 16'd65327, 16'd51401, 16'd57191, 16'd8335});
	test_expansion(128'hb777400d36162e138de26d3e3cfb3508, {16'd46322, 16'd47441, 16'd37259, 16'd48497, 16'd49002, 16'd26192, 16'd49263, 16'd7427, 16'd16253, 16'd15179, 16'd11733, 16'd49907, 16'd58533, 16'd63948, 16'd61890, 16'd25260, 16'd38124, 16'd20843, 16'd20677, 16'd41340, 16'd14340, 16'd57795, 16'd59028, 16'd20940, 16'd55181, 16'd63935});
	test_expansion(128'hec64e326563bcd4c5981f459047207f0, {16'd56781, 16'd41868, 16'd19032, 16'd7032, 16'd8671, 16'd65487, 16'd50104, 16'd11337, 16'd26136, 16'd41256, 16'd25865, 16'd19448, 16'd41332, 16'd49930, 16'd25703, 16'd30151, 16'd60241, 16'd32243, 16'd34600, 16'd48319, 16'd45101, 16'd37721, 16'd52718, 16'd41974, 16'd2008, 16'd33632});
	test_expansion(128'h55e881921c7c04620592626d1a7b680d, {16'd51714, 16'd63982, 16'd57878, 16'd60178, 16'd21263, 16'd25395, 16'd21835, 16'd32065, 16'd5256, 16'd54511, 16'd4388, 16'd40515, 16'd60064, 16'd9915, 16'd48836, 16'd60711, 16'd32067, 16'd5330, 16'd30103, 16'd29614, 16'd46292, 16'd10148, 16'd53509, 16'd35535, 16'd57369, 16'd54124});
	test_expansion(128'h9292eb2cbc1ea71f2a763800ea09ab6d, {16'd44675, 16'd40851, 16'd17320, 16'd44026, 16'd42363, 16'd29584, 16'd53816, 16'd49623, 16'd54402, 16'd62267, 16'd44677, 16'd48845, 16'd963, 16'd31110, 16'd42083, 16'd19965, 16'd54716, 16'd28927, 16'd22204, 16'd64439, 16'd11751, 16'd54768, 16'd18316, 16'd27423, 16'd37010, 16'd8198});
	test_expansion(128'hef68454dafde8d4cb566a2a62d43b8e9, {16'd55511, 16'd40274, 16'd31007, 16'd35753, 16'd15437, 16'd60876, 16'd14355, 16'd48993, 16'd45641, 16'd2676, 16'd23713, 16'd6498, 16'd19687, 16'd32639, 16'd62839, 16'd22291, 16'd35345, 16'd12952, 16'd55520, 16'd55307, 16'd18145, 16'd32298, 16'd57366, 16'd8203, 16'd5963, 16'd59633});
	test_expansion(128'h11dc29c23c1dc4dc27f4a2d2e3e447d1, {16'd22973, 16'd22498, 16'd30326, 16'd30829, 16'd23413, 16'd17610, 16'd32627, 16'd46556, 16'd29520, 16'd18739, 16'd11070, 16'd53710, 16'd46848, 16'd53411, 16'd12949, 16'd65050, 16'd24359, 16'd22816, 16'd30442, 16'd19029, 16'd60236, 16'd47581, 16'd13858, 16'd47730, 16'd8142, 16'd58035});
	test_expansion(128'hb00687ca12825a4e7393f8deb88e7243, {16'd50992, 16'd59804, 16'd62448, 16'd12776, 16'd11244, 16'd64452, 16'd40000, 16'd51489, 16'd6767, 16'd53546, 16'd34915, 16'd1866, 16'd59060, 16'd29150, 16'd61732, 16'd7794, 16'd2232, 16'd20600, 16'd61403, 16'd36169, 16'd5014, 16'd16424, 16'd64715, 16'd61099, 16'd53990, 16'd24132});
	test_expansion(128'h41a29d31a0abb1e2db90773bbcbda665, {16'd14960, 16'd29022, 16'd6670, 16'd20000, 16'd64683, 16'd32048, 16'd61322, 16'd54447, 16'd59101, 16'd64809, 16'd3681, 16'd63153, 16'd2399, 16'd10344, 16'd32942, 16'd41166, 16'd64193, 16'd29612, 16'd13237, 16'd48444, 16'd60240, 16'd25646, 16'd6237, 16'd14731, 16'd38741, 16'd58828});
	test_expansion(128'hb550c3d5ad82bb0122d440d61df9620f, {16'd49248, 16'd10160, 16'd22805, 16'd1638, 16'd12460, 16'd43191, 16'd38037, 16'd56559, 16'd29154, 16'd9240, 16'd24153, 16'd16459, 16'd56069, 16'd15570, 16'd16859, 16'd42794, 16'd7178, 16'd23381, 16'd57441, 16'd40327, 16'd18152, 16'd21096, 16'd21307, 16'd51383, 16'd5309, 16'd24064});
	test_expansion(128'h9010a41232d8df6d9ded6f340a44127d, {16'd10855, 16'd16981, 16'd17835, 16'd63196, 16'd58850, 16'd16576, 16'd9226, 16'd24763, 16'd7359, 16'd36560, 16'd55534, 16'd58269, 16'd41646, 16'd47173, 16'd26340, 16'd25289, 16'd58240, 16'd33500, 16'd48173, 16'd9384, 16'd24628, 16'd7837, 16'd2274, 16'd61482, 16'd37453, 16'd165});
	test_expansion(128'hb7881e6c3fcf3b45b927012ba05ca750, {16'd46430, 16'd49635, 16'd46505, 16'd48487, 16'd47127, 16'd25811, 16'd38552, 16'd64355, 16'd44729, 16'd62666, 16'd41007, 16'd22654, 16'd13385, 16'd53328, 16'd15859, 16'd22674, 16'd3585, 16'd23674, 16'd27680, 16'd22222, 16'd1798, 16'd56824, 16'd49040, 16'd29918, 16'd17086, 16'd40567});
	test_expansion(128'h680bb6ce180003726482c837a4a71965, {16'd30388, 16'd20342, 16'd18431, 16'd29182, 16'd59089, 16'd21264, 16'd9203, 16'd28535, 16'd61436, 16'd48811, 16'd37107, 16'd8615, 16'd57571, 16'd50089, 16'd63295, 16'd1376, 16'd7030, 16'd7334, 16'd54141, 16'd29116, 16'd4546, 16'd3257, 16'd8267, 16'd4427, 16'd41359, 16'd40492});
	test_expansion(128'h0c9b809b99ae22cb9b00134235a809d2, {16'd17766, 16'd54911, 16'd37857, 16'd18489, 16'd37894, 16'd60688, 16'd17888, 16'd28133, 16'd40749, 16'd63670, 16'd42954, 16'd42665, 16'd47114, 16'd58730, 16'd62564, 16'd22935, 16'd43311, 16'd47857, 16'd39159, 16'd24582, 16'd28227, 16'd8838, 16'd25503, 16'd37254, 16'd57820, 16'd7400});
	test_expansion(128'h72d1cae2a444fb38a105af984524e338, {16'd20978, 16'd3498, 16'd5541, 16'd29392, 16'd19119, 16'd10673, 16'd29998, 16'd14936, 16'd2812, 16'd19879, 16'd37569, 16'd24334, 16'd34763, 16'd18973, 16'd20771, 16'd7826, 16'd25895, 16'd30456, 16'd27395, 16'd14783, 16'd53434, 16'd1863, 16'd51345, 16'd24999, 16'd8434, 16'd47651});
	test_expansion(128'h74453b1319e2015100e6d1b246734d91, {16'd55997, 16'd45716, 16'd5370, 16'd30059, 16'd48557, 16'd49798, 16'd38848, 16'd33960, 16'd60316, 16'd43059, 16'd42419, 16'd7526, 16'd33035, 16'd1355, 16'd57488, 16'd61936, 16'd63890, 16'd53423, 16'd130, 16'd28153, 16'd26833, 16'd28085, 16'd25159, 16'd40530, 16'd10128, 16'd19760});
	test_expansion(128'h47f4505c8e9b59ba479742beb2d7e72d, {16'd24492, 16'd3686, 16'd40888, 16'd63972, 16'd9347, 16'd64378, 16'd6557, 16'd35152, 16'd48219, 16'd2388, 16'd39719, 16'd33801, 16'd64770, 16'd9579, 16'd60486, 16'd9939, 16'd3279, 16'd42266, 16'd25128, 16'd28128, 16'd47103, 16'd62775, 16'd57367, 16'd39001, 16'd45308, 16'd26162});
	test_expansion(128'h6fc42957f8ef2ec37b90bca9d2f145da, {16'd34934, 16'd24659, 16'd11747, 16'd19205, 16'd1926, 16'd443, 16'd19094, 16'd54673, 16'd44451, 16'd40938, 16'd64780, 16'd4315, 16'd18435, 16'd1200, 16'd43299, 16'd17005, 16'd27500, 16'd3009, 16'd43447, 16'd17293, 16'd41586, 16'd20244, 16'd26208, 16'd34316, 16'd20564, 16'd3584});
	test_expansion(128'h8c4c62a79ec352be355497fcff7596a9, {16'd31801, 16'd45526, 16'd33446, 16'd23466, 16'd3612, 16'd34446, 16'd61121, 16'd47845, 16'd15560, 16'd56274, 16'd9853, 16'd64079, 16'd25680, 16'd29316, 16'd39574, 16'd8742, 16'd58133, 16'd12714, 16'd62547, 16'd57681, 16'd41409, 16'd54771, 16'd31865, 16'd24288, 16'd30155, 16'd36389});
	test_expansion(128'h8bff3dcd9538b4c13c1c0f4d34890c0e, {16'd8929, 16'd18526, 16'd38586, 16'd26889, 16'd36108, 16'd14170, 16'd13210, 16'd65412, 16'd43393, 16'd62205, 16'd11122, 16'd49189, 16'd51131, 16'd38466, 16'd59876, 16'd24939, 16'd44435, 16'd1112, 16'd61063, 16'd32948, 16'd50605, 16'd7362, 16'd56472, 16'd46616, 16'd24230, 16'd10396});
	test_expansion(128'he8d963af47aeb2ab74f69a064a465af8, {16'd40882, 16'd46031, 16'd35454, 16'd13392, 16'd26227, 16'd61734, 16'd4915, 16'd53935, 16'd62924, 16'd17665, 16'd11906, 16'd18067, 16'd11620, 16'd2435, 16'd36368, 16'd10729, 16'd7135, 16'd36755, 16'd43911, 16'd11756, 16'd16913, 16'd8587, 16'd12927, 16'd48837, 16'd25149, 16'd15653});
	test_expansion(128'h79b9ba24dc73235f77bd93e7685f2816, {16'd37876, 16'd16889, 16'd20666, 16'd56698, 16'd16182, 16'd44417, 16'd9939, 16'd43417, 16'd53231, 16'd30235, 16'd42563, 16'd30706, 16'd25678, 16'd42075, 16'd22040, 16'd58981, 16'd60412, 16'd48254, 16'd30162, 16'd2737, 16'd64611, 16'd39607, 16'd38756, 16'd13719, 16'd19728, 16'd62048});
	test_expansion(128'h90ebb4effdcdb79190ea3cd89821895d, {16'd23558, 16'd9899, 16'd20341, 16'd380, 16'd22809, 16'd24127, 16'd35760, 16'd37810, 16'd38306, 16'd54047, 16'd24260, 16'd59830, 16'd39278, 16'd18247, 16'd20962, 16'd23749, 16'd1938, 16'd35183, 16'd45510, 16'd32280, 16'd15648, 16'd41647, 16'd65166, 16'd15667, 16'd53984, 16'd8687});
	test_expansion(128'h15ab1800851c4662067cb1d3ce54f937, {16'd63984, 16'd24474, 16'd15112, 16'd33077, 16'd14772, 16'd19875, 16'd9028, 16'd40082, 16'd26800, 16'd17054, 16'd47506, 16'd29819, 16'd56772, 16'd61178, 16'd31417, 16'd23117, 16'd60527, 16'd51062, 16'd576, 16'd13944, 16'd35741, 16'd21739, 16'd14650, 16'd17107, 16'd2274, 16'd62505});
	test_expansion(128'h2d60da563b1bbfad9dd37093f0169296, {16'd61521, 16'd750, 16'd29030, 16'd53707, 16'd32830, 16'd40138, 16'd37979, 16'd57215, 16'd27116, 16'd52186, 16'd37341, 16'd21469, 16'd2756, 16'd10789, 16'd42976, 16'd13098, 16'd46747, 16'd21089, 16'd7968, 16'd53962, 16'd45237, 16'd9968, 16'd33147, 16'd34375, 16'd2078, 16'd39214});
	test_expansion(128'h291535eae70dc9c0f8bfa8cfeb7d49b1, {16'd20407, 16'd56166, 16'd8533, 16'd63514, 16'd57511, 16'd40752, 16'd2283, 16'd31708, 16'd24893, 16'd58416, 16'd29276, 16'd61411, 16'd35986, 16'd3379, 16'd33942, 16'd46717, 16'd38937, 16'd64177, 16'd23331, 16'd17202, 16'd24325, 16'd42381, 16'd48789, 16'd44896, 16'd23819, 16'd53782});
	test_expansion(128'h2f1b336e99a153ba61cd75744c03bab7, {16'd7529, 16'd46413, 16'd41893, 16'd46317, 16'd20749, 16'd35111, 16'd36180, 16'd15967, 16'd42910, 16'd61590, 16'd62035, 16'd33374, 16'd40178, 16'd30376, 16'd38070, 16'd28210, 16'd46511, 16'd13637, 16'd43486, 16'd43285, 16'd49971, 16'd12119, 16'd42656, 16'd45805, 16'd42523, 16'd7184});
	test_expansion(128'he1c8463025337566144ba20d284a5f2c, {16'd63661, 16'd22896, 16'd45612, 16'd65465, 16'd15948, 16'd20021, 16'd62792, 16'd52521, 16'd16628, 16'd14155, 16'd51138, 16'd61032, 16'd62152, 16'd56663, 16'd16031, 16'd32905, 16'd2357, 16'd21327, 16'd38581, 16'd8214, 16'd21044, 16'd27501, 16'd42386, 16'd3776, 16'd33340, 16'd12710});
	test_expansion(128'h9199b45a6c56f984e3d8cf721420a299, {16'd16767, 16'd10202, 16'd5373, 16'd11236, 16'd22666, 16'd7971, 16'd30982, 16'd25082, 16'd26338, 16'd9362, 16'd50358, 16'd40534, 16'd19449, 16'd49546, 16'd1540, 16'd9545, 16'd44299, 16'd15829, 16'd14306, 16'd4201, 16'd50499, 16'd23126, 16'd49504, 16'd55128, 16'd12430, 16'd38297});
	test_expansion(128'h4731e093049375408029f2b9054cf250, {16'd46333, 16'd6370, 16'd4039, 16'd38296, 16'd36405, 16'd50206, 16'd23909, 16'd54788, 16'd37105, 16'd32273, 16'd52634, 16'd45624, 16'd37510, 16'd28538, 16'd28349, 16'd49490, 16'd31560, 16'd38388, 16'd4404, 16'd5194, 16'd29307, 16'd138, 16'd20182, 16'd11046, 16'd10503, 16'd43045});
	test_expansion(128'h4cb1b0ac68e950ff178bf17f0c692765, {16'd45314, 16'd57256, 16'd42700, 16'd21469, 16'd63202, 16'd34547, 16'd21419, 16'd3849, 16'd2769, 16'd62081, 16'd52052, 16'd64619, 16'd3906, 16'd40171, 16'd44833, 16'd61853, 16'd22320, 16'd40336, 16'd56924, 16'd37262, 16'd36172, 16'd28590, 16'd13297, 16'd21918, 16'd51331, 16'd44604});
	test_expansion(128'h6027b6b460449160be6a3eaa4eef7737, {16'd6400, 16'd32779, 16'd1662, 16'd56501, 16'd56109, 16'd46299, 16'd24021, 16'd57622, 16'd62061, 16'd24781, 16'd23875, 16'd17156, 16'd51335, 16'd6761, 16'd29505, 16'd56367, 16'd64827, 16'd22494, 16'd9108, 16'd9207, 16'd27671, 16'd55597, 16'd38073, 16'd18644, 16'd1267, 16'd16841});
	test_expansion(128'hc057beedc7632004af33926d9895677b, {16'd7649, 16'd50958, 16'd35230, 16'd45239, 16'd444, 16'd32358, 16'd9455, 16'd20559, 16'd31480, 16'd31620, 16'd9203, 16'd50599, 16'd28635, 16'd57667, 16'd54265, 16'd60887, 16'd4274, 16'd57972, 16'd17754, 16'd48461, 16'd17477, 16'd61555, 16'd52597, 16'd40531, 16'd3673, 16'd684});
	test_expansion(128'hb51ef8502b9aaff40660c39f466fc45d, {16'd62524, 16'd27769, 16'd45250, 16'd1514, 16'd56394, 16'd25156, 16'd21257, 16'd41802, 16'd21667, 16'd3960, 16'd31240, 16'd29018, 16'd48251, 16'd38748, 16'd22383, 16'd36275, 16'd20348, 16'd3002, 16'd21422, 16'd8027, 16'd25343, 16'd18800, 16'd60933, 16'd39652, 16'd29858, 16'd55857});
	test_expansion(128'hc1790be8a36681649e4fcde8cbee13fb, {16'd33484, 16'd65324, 16'd6554, 16'd10317, 16'd20477, 16'd52670, 16'd57072, 16'd63179, 16'd61474, 16'd55463, 16'd12547, 16'd16529, 16'd15951, 16'd16710, 16'd58445, 16'd5896, 16'd62940, 16'd33851, 16'd23944, 16'd39571, 16'd36565, 16'd45676, 16'd14949, 16'd45077, 16'd28819, 16'd29795});
	test_expansion(128'h047009c10bc86074d1d3d102724ee813, {16'd21202, 16'd497, 16'd57357, 16'd46211, 16'd23103, 16'd18758, 16'd63169, 16'd45431, 16'd58489, 16'd29505, 16'd60001, 16'd59254, 16'd38549, 16'd2545, 16'd33134, 16'd25887, 16'd19712, 16'd37763, 16'd17786, 16'd38137, 16'd58357, 16'd34602, 16'd61046, 16'd55821, 16'd4588, 16'd11576});
	test_expansion(128'ha2d42e25f2625110f23e679d6fec71de, {16'd14725, 16'd38058, 16'd37961, 16'd29090, 16'd17603, 16'd18720, 16'd59601, 16'd8256, 16'd41862, 16'd41185, 16'd23662, 16'd41586, 16'd27223, 16'd50371, 16'd9763, 16'd22747, 16'd4283, 16'd29070, 16'd42181, 16'd34140, 16'd46478, 16'd32801, 16'd24477, 16'd44780, 16'd30968, 16'd53113});
	test_expansion(128'he45787e462484cd4c130f6268200e48e, {16'd18194, 16'd34675, 16'd10160, 16'd35592, 16'd30982, 16'd50545, 16'd9400, 16'd32354, 16'd2119, 16'd55133, 16'd46618, 16'd8980, 16'd15583, 16'd59440, 16'd19381, 16'd21286, 16'd22083, 16'd55602, 16'd19072, 16'd1273, 16'd35779, 16'd17529, 16'd4569, 16'd17684, 16'd61046, 16'd18282});
	test_expansion(128'h3a3bbdaad164efd8aa83e381e1089c60, {16'd32064, 16'd29316, 16'd56804, 16'd49759, 16'd8241, 16'd16453, 16'd20015, 16'd22294, 16'd20045, 16'd65241, 16'd26073, 16'd8896, 16'd10449, 16'd4594, 16'd43596, 16'd36496, 16'd3936, 16'd19107, 16'd32612, 16'd16513, 16'd6336, 16'd63135, 16'd44117, 16'd6905, 16'd53658, 16'd50919});
	test_expansion(128'h9a30e0478e60bb284774b26ed57baefd, {16'd37892, 16'd53062, 16'd56875, 16'd26016, 16'd9383, 16'd13886, 16'd24929, 16'd60440, 16'd471, 16'd30938, 16'd26039, 16'd32204, 16'd57246, 16'd25682, 16'd16072, 16'd36336, 16'd41658, 16'd560, 16'd23380, 16'd23771, 16'd34458, 16'd63502, 16'd25176, 16'd63672, 16'd10117, 16'd17517});
	test_expansion(128'h3310ae2ca65c0871336ab0f20c1640c6, {16'd56725, 16'd11958, 16'd476, 16'd55894, 16'd19355, 16'd26782, 16'd31028, 16'd12711, 16'd3047, 16'd25306, 16'd58867, 16'd36494, 16'd3492, 16'd6746, 16'd16371, 16'd7607, 16'd2398, 16'd61731, 16'd19600, 16'd10570, 16'd1523, 16'd64912, 16'd41880, 16'd32952, 16'd49727, 16'd21094});
	test_expansion(128'h49b2543bb643afb1b8338ae028efbcbe, {16'd61029, 16'd17900, 16'd53684, 16'd56419, 16'd63650, 16'd24378, 16'd30099, 16'd38375, 16'd55371, 16'd617, 16'd65117, 16'd47231, 16'd53176, 16'd23280, 16'd26434, 16'd14655, 16'd55303, 16'd10060, 16'd24501, 16'd17883, 16'd39780, 16'd21981, 16'd16317, 16'd62935, 16'd21165, 16'd54950});
	test_expansion(128'hfdbf7f155e38e9537c8f0239c20ae3f8, {16'd37815, 16'd18629, 16'd62560, 16'd49718, 16'd215, 16'd35941, 16'd62806, 16'd32118, 16'd62054, 16'd36803, 16'd49259, 16'd1998, 16'd29771, 16'd63881, 16'd20768, 16'd11170, 16'd47463, 16'd43181, 16'd50729, 16'd13945, 16'd23179, 16'd36026, 16'd49765, 16'd41134, 16'd39120, 16'd41685});
	test_expansion(128'hb28c2cbba6a5820f7a282597e1243bf4, {16'd64419, 16'd28445, 16'd17006, 16'd33339, 16'd48655, 16'd12113, 16'd27658, 16'd25342, 16'd13085, 16'd9313, 16'd18368, 16'd62672, 16'd42107, 16'd4697, 16'd63758, 16'd21097, 16'd31008, 16'd57107, 16'd2022, 16'd2086, 16'd18752, 16'd4102, 16'd22681, 16'd6013, 16'd52144, 16'd6005});
	test_expansion(128'h228277b0063cc391a360e02fd95b1777, {16'd668, 16'd63120, 16'd33662, 16'd39618, 16'd59142, 16'd11597, 16'd8770, 16'd27466, 16'd63148, 16'd19493, 16'd19593, 16'd41174, 16'd42901, 16'd27362, 16'd13071, 16'd58389, 16'd33982, 16'd9668, 16'd12249, 16'd9846, 16'd2410, 16'd29874, 16'd13637, 16'd14135, 16'd4161, 16'd63472});
	test_expansion(128'h41d3f8a202b29c2a013326601e88b128, {16'd28149, 16'd45670, 16'd12103, 16'd31631, 16'd42407, 16'd52897, 16'd31295, 16'd26510, 16'd41893, 16'd8328, 16'd34883, 16'd60724, 16'd14720, 16'd5411, 16'd13575, 16'd16734, 16'd21953, 16'd33652, 16'd12549, 16'd60862, 16'd56598, 16'd49360, 16'd43945, 16'd25797, 16'd2835, 16'd59940});
	test_expansion(128'hbc0f88b649872b83029191adb1e0b9cd, {16'd38472, 16'd54255, 16'd32747, 16'd45638, 16'd31046, 16'd61043, 16'd42222, 16'd2976, 16'd64547, 16'd4455, 16'd50432, 16'd47796, 16'd7923, 16'd55106, 16'd14880, 16'd45432, 16'd7889, 16'd20719, 16'd7637, 16'd14880, 16'd29368, 16'd24320, 16'd46339, 16'd17670, 16'd19371, 16'd31912});
	test_expansion(128'hda0ca43abb89781522c7413e3a6efc0e, {16'd52676, 16'd54195, 16'd22396, 16'd33702, 16'd10600, 16'd24920, 16'd54580, 16'd28126, 16'd37538, 16'd28928, 16'd30348, 16'd42013, 16'd20356, 16'd10982, 16'd61123, 16'd61690, 16'd47088, 16'd29425, 16'd22630, 16'd25892, 16'd42196, 16'd9408, 16'd34312, 16'd36089, 16'd54131, 16'd1005});
	test_expansion(128'hd74fc8d30c8482779a33516fa7329024, {16'd17785, 16'd50205, 16'd7132, 16'd18847, 16'd6935, 16'd20391, 16'd54321, 16'd31244, 16'd44, 16'd5092, 16'd13091, 16'd16809, 16'd358, 16'd33822, 16'd54383, 16'd14974, 16'd42056, 16'd10667, 16'd48406, 16'd9164, 16'd11263, 16'd13657, 16'd37151, 16'd7710, 16'd62259, 16'd51175});
	test_expansion(128'hddff588895a80915f8d3717fa5dbc9f1, {16'd61695, 16'd58086, 16'd57115, 16'd36024, 16'd21846, 16'd58290, 16'd29272, 16'd49328, 16'd54880, 16'd12220, 16'd42746, 16'd11755, 16'd32166, 16'd59185, 16'd10984, 16'd62662, 16'd63169, 16'd56354, 16'd7011, 16'd16005, 16'd21431, 16'd24716, 16'd11995, 16'd12963, 16'd22739, 16'd28132});
	test_expansion(128'hb67eab9c0c122d45d897d2cc255b80a0, {16'd18288, 16'd24616, 16'd26591, 16'd34662, 16'd54893, 16'd56114, 16'd63463, 16'd44332, 16'd3527, 16'd54762, 16'd33177, 16'd29803, 16'd59152, 16'd30662, 16'd42159, 16'd52489, 16'd8735, 16'd57704, 16'd61343, 16'd56886, 16'd18929, 16'd39905, 16'd23772, 16'd29846, 16'd59255, 16'd42467});
	test_expansion(128'hbfc65af1a917bf7361059a1d4e02dd7e, {16'd51112, 16'd33624, 16'd32341, 16'd974, 16'd53767, 16'd12125, 16'd49248, 16'd14067, 16'd49316, 16'd50361, 16'd10944, 16'd16317, 16'd19086, 16'd23712, 16'd34940, 16'd53818, 16'd26354, 16'd21063, 16'd61164, 16'd25743, 16'd13239, 16'd63006, 16'd11183, 16'd21394, 16'd20300, 16'd3521});
	test_expansion(128'h1db1750de2f876d143390bcb2b12f309, {16'd31468, 16'd57439, 16'd21771, 16'd58227, 16'd18719, 16'd42419, 16'd26307, 16'd29489, 16'd3245, 16'd15815, 16'd14707, 16'd2481, 16'd50499, 16'd58985, 16'd33904, 16'd32514, 16'd47838, 16'd36324, 16'd45471, 16'd62749, 16'd46206, 16'd61783, 16'd40828, 16'd11972, 16'd25983, 16'd9575});
	test_expansion(128'h93a214246024f14f0a35936975385035, {16'd41848, 16'd61656, 16'd13074, 16'd38772, 16'd19250, 16'd37221, 16'd27799, 16'd37369, 16'd30905, 16'd1249, 16'd30887, 16'd54491, 16'd55395, 16'd14680, 16'd37109, 16'd6751, 16'd13843, 16'd34813, 16'd42337, 16'd53021, 16'd41896, 16'd21532, 16'd35581, 16'd52258, 16'd25333, 16'd64804});
	test_expansion(128'h10e36404ad0da1ccfe959d58327e1f9f, {16'd13365, 16'd27135, 16'd62536, 16'd43006, 16'd31549, 16'd9770, 16'd59490, 16'd63240, 16'd55993, 16'd38482, 16'd13343, 16'd45956, 16'd8884, 16'd62670, 16'd45067, 16'd22039, 16'd12682, 16'd31300, 16'd27083, 16'd28235, 16'd30486, 16'd45876, 16'd16649, 16'd42929, 16'd48302, 16'd45494});
	test_expansion(128'hea7b2cfb7f164fe5cbbe48616d5bb3c4, {16'd23180, 16'd63150, 16'd19516, 16'd59595, 16'd40620, 16'd14210, 16'd13284, 16'd16666, 16'd44943, 16'd31075, 16'd4788, 16'd46178, 16'd51610, 16'd2248, 16'd39785, 16'd18466, 16'd32286, 16'd44019, 16'd22062, 16'd31645, 16'd6317, 16'd21364, 16'd34220, 16'd43193, 16'd33573, 16'd27783});
	test_expansion(128'h04c9137c19c569350bc350d296d3ff3b, {16'd30608, 16'd2428, 16'd54235, 16'd32482, 16'd13769, 16'd746, 16'd54774, 16'd1756, 16'd56664, 16'd63644, 16'd22796, 16'd16724, 16'd15525, 16'd8163, 16'd46835, 16'd20290, 16'd47636, 16'd49958, 16'd36807, 16'd40969, 16'd41014, 16'd44847, 16'd54259, 16'd39139, 16'd24429, 16'd36970});
	test_expansion(128'h2725832195fd3f95cf47718bc7c08ab3, {16'd1411, 16'd28635, 16'd14182, 16'd13296, 16'd12665, 16'd20121, 16'd1718, 16'd31177, 16'd56240, 16'd37154, 16'd28155, 16'd30243, 16'd43664, 16'd48326, 16'd18980, 16'd6798, 16'd53835, 16'd61988, 16'd36830, 16'd2945, 16'd22052, 16'd46289, 16'd63217, 16'd53153, 16'd33055, 16'd16057});
	test_expansion(128'hc0997e4bed673847346d41ad80d34d83, {16'd10393, 16'd56086, 16'd58493, 16'd65393, 16'd26561, 16'd24005, 16'd24796, 16'd51687, 16'd47994, 16'd7629, 16'd42813, 16'd20165, 16'd1180, 16'd43846, 16'd48554, 16'd22593, 16'd15524, 16'd12148, 16'd2880, 16'd11466, 16'd51876, 16'd61203, 16'd5735, 16'd28108, 16'd23454, 16'd6118});
	test_expansion(128'had4a14e68a45bac994d0878e53dbd073, {16'd20426, 16'd52497, 16'd24078, 16'd4327, 16'd16463, 16'd55025, 16'd13723, 16'd10583, 16'd9415, 16'd31375, 16'd42075, 16'd5565, 16'd32520, 16'd3369, 16'd21833, 16'd27097, 16'd29461, 16'd25509, 16'd12704, 16'd44168, 16'd13894, 16'd4343, 16'd48661, 16'd14467, 16'd52639, 16'd52420});
	test_expansion(128'hef3e4723bb47681622862aa37bc076c7, {16'd34017, 16'd6535, 16'd22779, 16'd4034, 16'd43088, 16'd54781, 16'd38363, 16'd52378, 16'd22680, 16'd10825, 16'd50600, 16'd34172, 16'd1553, 16'd54276, 16'd31072, 16'd50310, 16'd4514, 16'd34220, 16'd49715, 16'd36431, 16'd23513, 16'd62641, 16'd22124, 16'd63501, 16'd23231, 16'd39057});
	test_expansion(128'h13607414afbbc689c3bd226018da6fbf, {16'd28909, 16'd39477, 16'd61748, 16'd31540, 16'd27680, 16'd62528, 16'd29087, 16'd24709, 16'd41519, 16'd26554, 16'd9819, 16'd39406, 16'd35970, 16'd26089, 16'd6433, 16'd46032, 16'd20842, 16'd11194, 16'd50784, 16'd14394, 16'd22624, 16'd18832, 16'd13011, 16'd42474, 16'd22695, 16'd25516});
	test_expansion(128'h3690589b94fbf10d13512509cb9d3aff, {16'd25085, 16'd9442, 16'd12685, 16'd53767, 16'd9591, 16'd799, 16'd47765, 16'd15777, 16'd15234, 16'd61673, 16'd33187, 16'd52673, 16'd46007, 16'd62127, 16'd3487, 16'd10705, 16'd25981, 16'd30180, 16'd36190, 16'd1318, 16'd42171, 16'd51456, 16'd18985, 16'd36702, 16'd14884, 16'd55566});
	test_expansion(128'hb735a93b3230b2e5821d905795d9f68f, {16'd26860, 16'd59440, 16'd59419, 16'd43538, 16'd36134, 16'd45332, 16'd59626, 16'd27792, 16'd10798, 16'd46474, 16'd34105, 16'd19311, 16'd14659, 16'd55151, 16'd49226, 16'd64158, 16'd54177, 16'd7754, 16'd7950, 16'd38041, 16'd9859, 16'd32292, 16'd1190, 16'd65000, 16'd3981, 16'd55630});
	test_expansion(128'hc359ff1f3821607cd92b15ffc65d8321, {16'd50442, 16'd25450, 16'd21211, 16'd23123, 16'd12323, 16'd33023, 16'd62822, 16'd53, 16'd16001, 16'd54688, 16'd29615, 16'd49604, 16'd25733, 16'd38674, 16'd45934, 16'd33778, 16'd34806, 16'd41504, 16'd26147, 16'd27727, 16'd58614, 16'd39786, 16'd52007, 16'd61860, 16'd43135, 16'd59925});
	test_expansion(128'h892b3c8121f2d15d0d77514448212ac6, {16'd8212, 16'd48899, 16'd36301, 16'd3297, 16'd56027, 16'd30147, 16'd26754, 16'd53768, 16'd56115, 16'd49589, 16'd29603, 16'd16596, 16'd38124, 16'd13677, 16'd12756, 16'd46682, 16'd7913, 16'd3037, 16'd14489, 16'd62001, 16'd22144, 16'd30481, 16'd21521, 16'd34254, 16'd45746, 16'd38217});
	test_expansion(128'h4699610d3c2ab6d360713ac48819d579, {16'd7783, 16'd8537, 16'd49366, 16'd9843, 16'd36486, 16'd6048, 16'd64483, 16'd35720, 16'd54246, 16'd47140, 16'd27333, 16'd12665, 16'd33457, 16'd7636, 16'd29129, 16'd30357, 16'd43399, 16'd54669, 16'd34226, 16'd41794, 16'd54733, 16'd4528, 16'd19830, 16'd27880, 16'd63584, 16'd61218});
	test_expansion(128'hf191af0ac18985af1a1e1efb78bea042, {16'd2032, 16'd25452, 16'd55398, 16'd14809, 16'd8413, 16'd8393, 16'd28510, 16'd24539, 16'd43335, 16'd52559, 16'd15635, 16'd58853, 16'd17860, 16'd43717, 16'd7744, 16'd54287, 16'd36355, 16'd37604, 16'd31736, 16'd34321, 16'd32146, 16'd54363, 16'd11574, 16'd50521, 16'd31802, 16'd31717});
	test_expansion(128'h560b3ddb0fca0be56ce9e70c28321c27, {16'd4320, 16'd61810, 16'd31072, 16'd42113, 16'd34427, 16'd27768, 16'd51749, 16'd3155, 16'd51607, 16'd48442, 16'd50499, 16'd4349, 16'd38914, 16'd33142, 16'd38082, 16'd64931, 16'd21167, 16'd11610, 16'd48113, 16'd9327, 16'd49121, 16'd30759, 16'd43390, 16'd13546, 16'd13294, 16'd5915});
	test_expansion(128'h9986d2ab9be7ded993f08bf549c43e3a, {16'd59182, 16'd34400, 16'd27276, 16'd18183, 16'd65444, 16'd10181, 16'd17928, 16'd48497, 16'd35434, 16'd39518, 16'd26899, 16'd9654, 16'd31441, 16'd15958, 16'd27755, 16'd48481, 16'd41307, 16'd1023, 16'd3230, 16'd4672, 16'd52781, 16'd22146, 16'd15012, 16'd63468, 16'd21485, 16'd29469});
	test_expansion(128'h26b2d8421246163f5fbbacbb0b5b18e9, {16'd19361, 16'd29209, 16'd44287, 16'd17653, 16'd36951, 16'd1672, 16'd6703, 16'd28623, 16'd30956, 16'd14345, 16'd30080, 16'd28677, 16'd48210, 16'd61956, 16'd49579, 16'd16115, 16'd18426, 16'd42, 16'd60993, 16'd4173, 16'd1505, 16'd34989, 16'd20542, 16'd27466, 16'd52652, 16'd10164});
	test_expansion(128'h8a8d045b52697f757e104fe8293a41eb, {16'd57735, 16'd58441, 16'd13989, 16'd38061, 16'd8217, 16'd11949, 16'd33610, 16'd13740, 16'd43080, 16'd15765, 16'd21234, 16'd37353, 16'd46359, 16'd45130, 16'd48783, 16'd62043, 16'd2941, 16'd9430, 16'd41600, 16'd58704, 16'd22030, 16'd52384, 16'd63364, 16'd7977, 16'd43874, 16'd61506});
	test_expansion(128'h1bac0f5b498ed8d9133d08dd91e557d5, {16'd63268, 16'd5192, 16'd13019, 16'd1415, 16'd58310, 16'd18660, 16'd62173, 16'd13169, 16'd50561, 16'd44910, 16'd43151, 16'd42714, 16'd47842, 16'd28747, 16'd59100, 16'd16284, 16'd32243, 16'd53944, 16'd41836, 16'd57989, 16'd38183, 16'd60184, 16'd60808, 16'd27806, 16'd54315, 16'd25437});
	test_expansion(128'h05cf18d40197282b4312f4fdf71163e2, {16'd5492, 16'd16553, 16'd24282, 16'd25219, 16'd47031, 16'd33128, 16'd38846, 16'd64195, 16'd9746, 16'd59246, 16'd30305, 16'd3801, 16'd34588, 16'd25722, 16'd16026, 16'd34100, 16'd1152, 16'd15926, 16'd45473, 16'd14222, 16'd21671, 16'd3297, 16'd30237, 16'd54861, 16'd40057, 16'd20756});
	test_expansion(128'h3fa0374e35758295f39ff4240ea0bcc0, {16'd54970, 16'd60402, 16'd44297, 16'd33850, 16'd22187, 16'd35170, 16'd56077, 16'd6798, 16'd35219, 16'd9675, 16'd21919, 16'd38653, 16'd53824, 16'd44712, 16'd59780, 16'd34959, 16'd22227, 16'd27717, 16'd62728, 16'd55946, 16'd52238, 16'd17398, 16'd23675, 16'd16526, 16'd51776, 16'd56817});
	test_expansion(128'hc219dc017edb0a60ee2c9af35b65fddd, {16'd14586, 16'd24146, 16'd40799, 16'd52294, 16'd46664, 16'd17728, 16'd46934, 16'd5459, 16'd5268, 16'd18966, 16'd42549, 16'd14488, 16'd5714, 16'd4080, 16'd51543, 16'd12790, 16'd30522, 16'd9481, 16'd35684, 16'd7482, 16'd56516, 16'd15324, 16'd29076, 16'd1002, 16'd2808, 16'd62401});
	test_expansion(128'h3032c8381cc727c6a716da2dbae8ddc9, {16'd64863, 16'd1853, 16'd64120, 16'd30591, 16'd57093, 16'd49753, 16'd39848, 16'd52091, 16'd304, 16'd40794, 16'd43842, 16'd10290, 16'd41013, 16'd21588, 16'd26175, 16'd46341, 16'd44632, 16'd9284, 16'd52714, 16'd29014, 16'd34369, 16'd34283, 16'd25312, 16'd17989, 16'd31298, 16'd53668});
	test_expansion(128'h0492bc7720db4139fb2aaf6fd9260297, {16'd45789, 16'd58319, 16'd8499, 16'd42283, 16'd31923, 16'd51198, 16'd39198, 16'd26372, 16'd41591, 16'd49171, 16'd23926, 16'd34694, 16'd8352, 16'd28011, 16'd59466, 16'd35845, 16'd32509, 16'd14169, 16'd12588, 16'd39329, 16'd22915, 16'd57401, 16'd7030, 16'd46565, 16'd20755, 16'd30965});
	test_expansion(128'h26786e10b5c4449e1e34a054e0c48022, {16'd16417, 16'd14738, 16'd47293, 16'd1949, 16'd17973, 16'd47407, 16'd42031, 16'd3101, 16'd62905, 16'd34450, 16'd63918, 16'd54028, 16'd1276, 16'd43382, 16'd54341, 16'd35983, 16'd16647, 16'd43480, 16'd33268, 16'd36356, 16'd18114, 16'd50862, 16'd81, 16'd47169, 16'd27621, 16'd46760});
	test_expansion(128'h87efd855c61ead630b0598bc140f9df7, {16'd30177, 16'd15066, 16'd14765, 16'd52570, 16'd57851, 16'd26848, 16'd47735, 16'd46354, 16'd9581, 16'd33937, 16'd24257, 16'd36837, 16'd34971, 16'd24758, 16'd4509, 16'd1117, 16'd53572, 16'd26931, 16'd5003, 16'd58990, 16'd19779, 16'd5540, 16'd53909, 16'd33330, 16'd39438, 16'd18318});
	test_expansion(128'hbe3e40792180eaba2875cecefc12f05a, {16'd21500, 16'd17114, 16'd16569, 16'd59527, 16'd11793, 16'd13973, 16'd58619, 16'd16715, 16'd27681, 16'd20549, 16'd23343, 16'd2758, 16'd28476, 16'd1290, 16'd12409, 16'd731, 16'd15195, 16'd38600, 16'd25465, 16'd25755, 16'd59976, 16'd37043, 16'd12321, 16'd10696, 16'd18875, 16'd48504});
	test_expansion(128'hcee45fb8ce635d3f1fbeac2649793847, {16'd49236, 16'd28246, 16'd48679, 16'd7605, 16'd62338, 16'd22694, 16'd25751, 16'd21312, 16'd3052, 16'd45026, 16'd52045, 16'd50490, 16'd31816, 16'd41214, 16'd4654, 16'd11339, 16'd37787, 16'd38933, 16'd7942, 16'd28126, 16'd14996, 16'd81, 16'd49218, 16'd57317, 16'd45469, 16'd57021});
	test_expansion(128'h347fe4c1a2f114242bbf4f5b5bd982aa, {16'd39561, 16'd9377, 16'd43997, 16'd61447, 16'd59894, 16'd2518, 16'd11474, 16'd45587, 16'd23630, 16'd59709, 16'd21332, 16'd20714, 16'd54250, 16'd55528, 16'd23899, 16'd34130, 16'd6598, 16'd8404, 16'd64841, 16'd3674, 16'd30264, 16'd38766, 16'd19172, 16'd32905, 16'd49573, 16'd39601});
	test_expansion(128'h813e72bb625614befb5b42e8bd1ccf76, {16'd11853, 16'd14352, 16'd26644, 16'd29534, 16'd2665, 16'd56930, 16'd45857, 16'd14360, 16'd4608, 16'd44336, 16'd25459, 16'd44674, 16'd34268, 16'd51299, 16'd13477, 16'd1010, 16'd28842, 16'd53350, 16'd27487, 16'd23702, 16'd3025, 16'd26549, 16'd58539, 16'd21711, 16'd40383, 16'd3522});
	test_expansion(128'h9e60d62e14f570fddec58c38cc0626df, {16'd25173, 16'd9313, 16'd64156, 16'd29711, 16'd25031, 16'd35902, 16'd52767, 16'd31224, 16'd26010, 16'd61423, 16'd46202, 16'd43038, 16'd22554, 16'd42251, 16'd19382, 16'd34103, 16'd52829, 16'd59525, 16'd60758, 16'd36384, 16'd18678, 16'd34541, 16'd33026, 16'd14769, 16'd28900, 16'd57894});
	test_expansion(128'h7b318cd1fd1daca52b5353393bd45c82, {16'd54663, 16'd42826, 16'd56295, 16'd30468, 16'd26567, 16'd43176, 16'd220, 16'd34200, 16'd53903, 16'd30875, 16'd18639, 16'd55575, 16'd52684, 16'd27242, 16'd786, 16'd42004, 16'd23518, 16'd6617, 16'd16334, 16'd33612, 16'd42927, 16'd45797, 16'd49005, 16'd32578, 16'd48373, 16'd31675});
	test_expansion(128'h2d2dabc50a53693a225a99acadc6c552, {16'd49761, 16'd43416, 16'd58179, 16'd14350, 16'd35922, 16'd51594, 16'd43095, 16'd42157, 16'd42110, 16'd34407, 16'd44234, 16'd19779, 16'd55082, 16'd23560, 16'd50737, 16'd50403, 16'd13801, 16'd24016, 16'd1368, 16'd59336, 16'd31290, 16'd35142, 16'd47716, 16'd58832, 16'd31398, 16'd48563});
	test_expansion(128'h1bab8bd7663f54a5c66cfd307a1431f2, {16'd57419, 16'd32597, 16'd18704, 16'd659, 16'd37449, 16'd35335, 16'd11526, 16'd31494, 16'd14839, 16'd631, 16'd7824, 16'd60050, 16'd49558, 16'd15972, 16'd16859, 16'd56263, 16'd50700, 16'd8009, 16'd21633, 16'd39671, 16'd50722, 16'd21649, 16'd35636, 16'd33130, 16'd8798, 16'd40308});
	test_expansion(128'h7255f9608964248f87bc008d60f4f54c, {16'd46906, 16'd38450, 16'd25693, 16'd64382, 16'd28516, 16'd21575, 16'd10113, 16'd63728, 16'd24272, 16'd20893, 16'd15618, 16'd8189, 16'd49110, 16'd39316, 16'd22064, 16'd50497, 16'd9838, 16'd6571, 16'd19151, 16'd55426, 16'd12253, 16'd24002, 16'd26918, 16'd41729, 16'd2587, 16'd20682});
	test_expansion(128'h3dbc871b8660f4018927bf9e9efbe95d, {16'd57365, 16'd9753, 16'd9217, 16'd54613, 16'd24149, 16'd47741, 16'd22801, 16'd56612, 16'd50786, 16'd32011, 16'd9309, 16'd22114, 16'd37767, 16'd61001, 16'd46826, 16'd52161, 16'd46112, 16'd5805, 16'd12000, 16'd17770, 16'd41921, 16'd61161, 16'd29943, 16'd6943, 16'd17056, 16'd36739});
	test_expansion(128'hcaf82409b17605a25405058a20bf20e1, {16'd41519, 16'd51966, 16'd7065, 16'd61658, 16'd18383, 16'd51571, 16'd22002, 16'd64001, 16'd49623, 16'd9462, 16'd11852, 16'd60166, 16'd28394, 16'd33467, 16'd22987, 16'd64790, 16'd63276, 16'd40294, 16'd31325, 16'd48224, 16'd8207, 16'd26022, 16'd64745, 16'd11544, 16'd58245, 16'd33073});
	test_expansion(128'h6fcb009a905a97dd5061b5e824047f65, {16'd3506, 16'd4736, 16'd125, 16'd20722, 16'd39818, 16'd20918, 16'd17833, 16'd55998, 16'd222, 16'd11064, 16'd53903, 16'd28666, 16'd62848, 16'd51871, 16'd20169, 16'd55708, 16'd31047, 16'd57742, 16'd46825, 16'd44511, 16'd49759, 16'd20356, 16'd36406, 16'd47432, 16'd22177, 16'd23639});
	test_expansion(128'h3e21f703dcadb9bc1c373ce7ce77de92, {16'd55165, 16'd42039, 16'd7054, 16'd17661, 16'd65088, 16'd3170, 16'd56052, 16'd54340, 16'd54178, 16'd24838, 16'd29532, 16'd62193, 16'd24056, 16'd53702, 16'd37118, 16'd26268, 16'd35440, 16'd51540, 16'd1694, 16'd54194, 16'd42773, 16'd7900, 16'd5914, 16'd5074, 16'd59977, 16'd37101});
	test_expansion(128'hc316b61d6fa78d010089fd0752933dad, {16'd62220, 16'd30035, 16'd28882, 16'd23687, 16'd16522, 16'd6168, 16'd47079, 16'd26117, 16'd41937, 16'd43005, 16'd38893, 16'd42369, 16'd48010, 16'd46312, 16'd53946, 16'd44902, 16'd15517, 16'd43391, 16'd50752, 16'd5537, 16'd51897, 16'd23226, 16'd43134, 16'd36854, 16'd27090, 16'd21086});
	test_expansion(128'h2b72afc3b70d1b85450a53a7dc2b0651, {16'd24785, 16'd16892, 16'd59622, 16'd7795, 16'd4460, 16'd4303, 16'd53464, 16'd25266, 16'd32004, 16'd12306, 16'd29078, 16'd44908, 16'd16674, 16'd28263, 16'd65089, 16'd58891, 16'd47083, 16'd56408, 16'd40691, 16'd19526, 16'd27337, 16'd12036, 16'd64859, 16'd26518, 16'd44297, 16'd54794});
	test_expansion(128'h280d9a2f6bfc74139c6a5d46de8b195a, {16'd58351, 16'd17740, 16'd6389, 16'd45997, 16'd61358, 16'd48627, 16'd41633, 16'd52435, 16'd6343, 16'd47684, 16'd47113, 16'd57598, 16'd56647, 16'd29479, 16'd7367, 16'd25959, 16'd20136, 16'd19654, 16'd6798, 16'd61655, 16'd22885, 16'd23160, 16'd61693, 16'd30723, 16'd60901, 16'd8071});
	test_expansion(128'h60e4105d5e524cdeab861f256e8f8ea9, {16'd36127, 16'd25406, 16'd41336, 16'd48960, 16'd1584, 16'd39237, 16'd34743, 16'd21342, 16'd19605, 16'd18130, 16'd25930, 16'd6684, 16'd25572, 16'd3532, 16'd61541, 16'd32331, 16'd15755, 16'd9900, 16'd36198, 16'd35545, 16'd16651, 16'd26714, 16'd38175, 16'd47891, 16'd62558, 16'd43504});
	test_expansion(128'h6c98d9247694bab33b14b74c970e3ce8, {16'd42829, 16'd37341, 16'd44668, 16'd54997, 16'd31086, 16'd26779, 16'd10082, 16'd38512, 16'd29390, 16'd22380, 16'd42719, 16'd47665, 16'd63785, 16'd34991, 16'd17465, 16'd37920, 16'd54596, 16'd22446, 16'd15436, 16'd8488, 16'd63836, 16'd47790, 16'd32474, 16'd16450, 16'd12652, 16'd30100});
	test_expansion(128'hd157d63dbf93301518440c8eddaa4b72, {16'd54527, 16'd62768, 16'd58621, 16'd58844, 16'd57231, 16'd55428, 16'd53731, 16'd26066, 16'd290, 16'd60684, 16'd58795, 16'd29419, 16'd2022, 16'd4731, 16'd16002, 16'd1815, 16'd28305, 16'd28594, 16'd17558, 16'd35257, 16'd8520, 16'd63588, 16'd6843, 16'd47785, 16'd44039, 16'd32898});
	test_expansion(128'h46d327dcbaff7b02aa39a71bf4dc9093, {16'd28632, 16'd49167, 16'd63829, 16'd24145, 16'd52479, 16'd16318, 16'd37913, 16'd38167, 16'd49961, 16'd523, 16'd44051, 16'd46228, 16'd17888, 16'd2180, 16'd29857, 16'd45547, 16'd61850, 16'd57494, 16'd54505, 16'd36674, 16'd31901, 16'd28124, 16'd33555, 16'd57745, 16'd17761, 16'd8998});
	test_expansion(128'he57b3c34aaf4c84dc2e688dca8263c74, {16'd11092, 16'd60788, 16'd16159, 16'd52195, 16'd59853, 16'd6378, 16'd51575, 16'd18549, 16'd59317, 16'd16186, 16'd19194, 16'd1754, 16'd47938, 16'd48020, 16'd42978, 16'd28338, 16'd30486, 16'd11815, 16'd43698, 16'd10723, 16'd4713, 16'd14796, 16'd10035, 16'd61212, 16'd19640, 16'd63885});
	test_expansion(128'h3d6ed0fb10049c0464e34992f9b95e60, {16'd7314, 16'd58772, 16'd6840, 16'd63033, 16'd57505, 16'd32508, 16'd44669, 16'd8775, 16'd26962, 16'd58593, 16'd35878, 16'd28912, 16'd11949, 16'd37574, 16'd61322, 16'd44514, 16'd23126, 16'd61713, 16'd47801, 16'd21930, 16'd43855, 16'd16656, 16'd53671, 16'd35110, 16'd40898, 16'd7695});
	test_expansion(128'h0dcb2c325bac274bed78e36f8a048fc3, {16'd52540, 16'd44489, 16'd53206, 16'd55897, 16'd6262, 16'd62710, 16'd57714, 16'd47557, 16'd17448, 16'd21026, 16'd15791, 16'd51519, 16'd57864, 16'd13361, 16'd3415, 16'd38142, 16'd56885, 16'd11299, 16'd47746, 16'd37606, 16'd64056, 16'd56077, 16'd59238, 16'd6471, 16'd57300, 16'd5078});
	test_expansion(128'h16a102ea8ee23db229f39efc63492041, {16'd15337, 16'd18285, 16'd64603, 16'd57180, 16'd11715, 16'd40938, 16'd39365, 16'd56702, 16'd44421, 16'd51373, 16'd39673, 16'd2328, 16'd9571, 16'd45902, 16'd40553, 16'd7368, 16'd20, 16'd41219, 16'd30113, 16'd23869, 16'd21008, 16'd6267, 16'd37715, 16'd8202, 16'd16705, 16'd53455});
	test_expansion(128'he3bfbeb4977bc4e7bfd08fc6d6f86d4e, {16'd46705, 16'd18589, 16'd47861, 16'd54019, 16'd20223, 16'd5965, 16'd13125, 16'd61738, 16'd46936, 16'd49973, 16'd43480, 16'd38996, 16'd8134, 16'd27191, 16'd25426, 16'd58798, 16'd35533, 16'd11271, 16'd44634, 16'd10200, 16'd26055, 16'd31604, 16'd13765, 16'd36097, 16'd62590, 16'd11151});
	test_expansion(128'hd39a38a789c5ae6f00e1a96758831481, {16'd61820, 16'd64783, 16'd32310, 16'd155, 16'd38832, 16'd21363, 16'd43113, 16'd13713, 16'd56509, 16'd44657, 16'd3214, 16'd34271, 16'd64681, 16'd56899, 16'd2979, 16'd58348, 16'd62394, 16'd9111, 16'd59780, 16'd12375, 16'd39860, 16'd26067, 16'd32521, 16'd57306, 16'd62858, 16'd41378});
	test_expansion(128'h278d56d50529312ef28a2809fa8435f2, {16'd61202, 16'd25643, 16'd58798, 16'd24028, 16'd12239, 16'd5296, 16'd43983, 16'd10375, 16'd1565, 16'd62702, 16'd51430, 16'd59096, 16'd33693, 16'd27117, 16'd37489, 16'd25294, 16'd57889, 16'd27044, 16'd53168, 16'd11148, 16'd59861, 16'd10896, 16'd8523, 16'd51288, 16'd47906, 16'd35791});
	test_expansion(128'h801107603d86dc4860d751f151364919, {16'd13718, 16'd60333, 16'd54255, 16'd6590, 16'd59776, 16'd50517, 16'd17232, 16'd42643, 16'd15683, 16'd57577, 16'd30754, 16'd17858, 16'd55169, 16'd58760, 16'd16640, 16'd8755, 16'd4460, 16'd8968, 16'd5547, 16'd18744, 16'd2527, 16'd33950, 16'd47374, 16'd54191, 16'd9884, 16'd12183});
	test_expansion(128'h3b37960d0d85c7df4fe3d13a267b7d1e, {16'd41341, 16'd26639, 16'd12654, 16'd36455, 16'd21493, 16'd44107, 16'd17592, 16'd42171, 16'd62566, 16'd32713, 16'd50247, 16'd48966, 16'd11437, 16'd26175, 16'd29200, 16'd36246, 16'd4534, 16'd8899, 16'd33275, 16'd60412, 16'd11246, 16'd60533, 16'd22106, 16'd9794, 16'd29249, 16'd14236});
	test_expansion(128'h0f9f7d762ce25422736161dbb88d9980, {16'd3022, 16'd34750, 16'd8532, 16'd31715, 16'd8175, 16'd18588, 16'd23040, 16'd54341, 16'd45236, 16'd23791, 16'd33821, 16'd32768, 16'd7742, 16'd60173, 16'd15533, 16'd45092, 16'd58835, 16'd61312, 16'd51743, 16'd55195, 16'd15301, 16'd35495, 16'd53813, 16'd4857, 16'd59292, 16'd13873});
	test_expansion(128'h3f820dbdb453b79a8efcd7298892391d, {16'd14353, 16'd39827, 16'd43071, 16'd52694, 16'd64541, 16'd50765, 16'd14556, 16'd47771, 16'd48207, 16'd14319, 16'd44033, 16'd48973, 16'd1149, 16'd57696, 16'd4615, 16'd8812, 16'd39136, 16'd62962, 16'd9569, 16'd61712, 16'd2616, 16'd27030, 16'd55377, 16'd3886, 16'd59089, 16'd42032});
	test_expansion(128'h296267d88f3b1b0f76e69f412686ac2e, {16'd39997, 16'd51658, 16'd35565, 16'd5137, 16'd29983, 16'd6989, 16'd1914, 16'd60623, 16'd1572, 16'd43085, 16'd57277, 16'd52441, 16'd1692, 16'd33175, 16'd30317, 16'd53452, 16'd53926, 16'd65450, 16'd62862, 16'd39305, 16'd47527, 16'd23434, 16'd59156, 16'd51992, 16'd34746, 16'd22383});
	test_expansion(128'h9015899b58beed69f0009f24185b118a, {16'd29183, 16'd932, 16'd22596, 16'd59501, 16'd10923, 16'd6562, 16'd32832, 16'd2579, 16'd51597, 16'd22627, 16'd10306, 16'd31383, 16'd34999, 16'd34435, 16'd27532, 16'd15874, 16'd58828, 16'd3685, 16'd58459, 16'd26104, 16'd62405, 16'd22607, 16'd44682, 16'd54686, 16'd63258, 16'd24798});
	test_expansion(128'h77603be1a66bccf1b954478dd061da3b, {16'd52812, 16'd18745, 16'd37223, 16'd42673, 16'd22916, 16'd16763, 16'd58919, 16'd7977, 16'd12855, 16'd52846, 16'd479, 16'd49538, 16'd9225, 16'd26423, 16'd2556, 16'd32087, 16'd1451, 16'd17562, 16'd51798, 16'd4172, 16'd18671, 16'd45318, 16'd51744, 16'd43480, 16'd35827, 16'd53044});
	test_expansion(128'h9b26f13c337f806f3e6712943473d654, {16'd64258, 16'd9211, 16'd43631, 16'd13493, 16'd53056, 16'd27867, 16'd63153, 16'd28945, 16'd51004, 16'd32026, 16'd41077, 16'd16077, 16'd50731, 16'd15012, 16'd33147, 16'd20248, 16'd59936, 16'd3604, 16'd34265, 16'd63632, 16'd27669, 16'd20173, 16'd1196, 16'd48459, 16'd53754, 16'd59587});
	test_expansion(128'h981b8126b587df40f146fd0c362704c8, {16'd18469, 16'd42074, 16'd26145, 16'd7537, 16'd44114, 16'd62864, 16'd29967, 16'd19228, 16'd21150, 16'd16722, 16'd18636, 16'd35293, 16'd44991, 16'd4437, 16'd49216, 16'd25179, 16'd53495, 16'd26321, 16'd50787, 16'd7464, 16'd12895, 16'd3453, 16'd23664, 16'd59981, 16'd49422, 16'd9584});
	test_expansion(128'h6bf157933a57cdd30ebd6c4273c33afb, {16'd62040, 16'd34728, 16'd11901, 16'd5473, 16'd33733, 16'd64770, 16'd38523, 16'd34611, 16'd26820, 16'd37794, 16'd40620, 16'd10465, 16'd26697, 16'd36393, 16'd44052, 16'd10925, 16'd32423, 16'd13155, 16'd60135, 16'd23749, 16'd33511, 16'd65015, 16'd5675, 16'd39645, 16'd39960, 16'd26522});
	test_expansion(128'h167a6e02daea737d17dc446cc620cb64, {16'd31632, 16'd51361, 16'd16286, 16'd40324, 16'd25657, 16'd34852, 16'd3863, 16'd55511, 16'd31605, 16'd49795, 16'd35497, 16'd15117, 16'd19274, 16'd11507, 16'd47511, 16'd60718, 16'd62110, 16'd43668, 16'd61310, 16'd4282, 16'd55050, 16'd60488, 16'd41376, 16'd37369, 16'd35329, 16'd27662});
	test_expansion(128'hf9265e9e023888fde9bd09e036a3036d, {16'd32004, 16'd5485, 16'd39428, 16'd40307, 16'd33394, 16'd62736, 16'd55339, 16'd24578, 16'd23681, 16'd65146, 16'd13587, 16'd53152, 16'd43064, 16'd51361, 16'd28202, 16'd33651, 16'd21830, 16'd3554, 16'd53402, 16'd34297, 16'd35213, 16'd61815, 16'd51156, 16'd4031, 16'd42945, 16'd62194});
	test_expansion(128'h000faff44d0e77ee3827f19f14ab8b1d, {16'd32683, 16'd2098, 16'd32406, 16'd31010, 16'd36638, 16'd14534, 16'd28897, 16'd37414, 16'd47470, 16'd5249, 16'd55927, 16'd32618, 16'd25082, 16'd33742, 16'd43376, 16'd6027, 16'd40561, 16'd4410, 16'd11282, 16'd51654, 16'd61945, 16'd51752, 16'd34940, 16'd38446, 16'd15390, 16'd51353});
	test_expansion(128'hb5544ac445fbe36669b4fc2cbce3a8dc, {16'd63854, 16'd59739, 16'd21812, 16'd44037, 16'd60893, 16'd38360, 16'd54738, 16'd14851, 16'd44833, 16'd41468, 16'd34871, 16'd45688, 16'd29859, 16'd50449, 16'd21084, 16'd26699, 16'd4526, 16'd59144, 16'd46073, 16'd64625, 16'd63176, 16'd65252, 16'd33099, 16'd32898, 16'd43706, 16'd50059});
	test_expansion(128'ha57c4c7cb4b6f7f7129d80200433fbc5, {16'd13134, 16'd32159, 16'd35618, 16'd36377, 16'd35600, 16'd44580, 16'd12097, 16'd31734, 16'd17949, 16'd54179, 16'd11407, 16'd62244, 16'd61666, 16'd21544, 16'd31830, 16'd34079, 16'd48862, 16'd46578, 16'd1975, 16'd62094, 16'd62247, 16'd58162, 16'd25563, 16'd18836, 16'd8032, 16'd10286});
	test_expansion(128'ha733cfe8082603a16e6e9c4939410e55, {16'd30277, 16'd1910, 16'd34307, 16'd34358, 16'd9213, 16'd17973, 16'd23606, 16'd52516, 16'd29047, 16'd4482, 16'd17042, 16'd40270, 16'd48027, 16'd23303, 16'd31860, 16'd56445, 16'd40425, 16'd25423, 16'd11306, 16'd2941, 16'd2863, 16'd16726, 16'd36781, 16'd17734, 16'd10580, 16'd24314});
	test_expansion(128'ha5e01c1fefbc368ad653bef1cfa9f022, {16'd4118, 16'd22831, 16'd8249, 16'd30822, 16'd4665, 16'd62779, 16'd41684, 16'd56623, 16'd22778, 16'd31673, 16'd13692, 16'd38741, 16'd64770, 16'd46714, 16'd16642, 16'd6943, 16'd48330, 16'd45339, 16'd57848, 16'd5380, 16'd17, 16'd33926, 16'd19964, 16'd30879, 16'd35984, 16'd40211});
	test_expansion(128'hb9f8b7a7652256c0ceccc28de05a079d, {16'd16456, 16'd44519, 16'd109, 16'd6773, 16'd53748, 16'd45438, 16'd15758, 16'd30217, 16'd60703, 16'd45806, 16'd1570, 16'd1302, 16'd15077, 16'd36025, 16'd63602, 16'd705, 16'd26445, 16'd23024, 16'd59088, 16'd15374, 16'd53494, 16'd17883, 16'd5535, 16'd40558, 16'd30032, 16'd1210});
	test_expansion(128'h39fe269f05b17af52526f968d8dcb5d9, {16'd28010, 16'd40929, 16'd42082, 16'd32970, 16'd22, 16'd34488, 16'd8587, 16'd32042, 16'd40550, 16'd12350, 16'd37166, 16'd5272, 16'd13565, 16'd21232, 16'd49449, 16'd14661, 16'd25511, 16'd50786, 16'd59460, 16'd36161, 16'd29495, 16'd53635, 16'd564, 16'd49463, 16'd22411, 16'd61219});
	test_expansion(128'h6eb7754a246d476fcff7103ce04846aa, {16'd27285, 16'd13740, 16'd23042, 16'd3590, 16'd52459, 16'd7566, 16'd347, 16'd57662, 16'd62263, 16'd12780, 16'd23444, 16'd11506, 16'd48764, 16'd65094, 16'd18355, 16'd45487, 16'd7604, 16'd28107, 16'd39453, 16'd17502, 16'd48688, 16'd50200, 16'd47991, 16'd35753, 16'd19012, 16'd16805});
	test_expansion(128'hbadc07e124bd80898912b5245607c8dd, {16'd14116, 16'd13279, 16'd7679, 16'd20790, 16'd44224, 16'd62119, 16'd59209, 16'd35508, 16'd64424, 16'd35883, 16'd10968, 16'd55384, 16'd24716, 16'd42622, 16'd32548, 16'd60836, 16'd55195, 16'd48095, 16'd44882, 16'd58672, 16'd56498, 16'd58647, 16'd44584, 16'd27745, 16'd1495, 16'd12382});
	test_expansion(128'hdab44987073f01e86aa973db886af952, {16'd23260, 16'd60733, 16'd50282, 16'd54852, 16'd47838, 16'd2549, 16'd2368, 16'd9580, 16'd41217, 16'd16462, 16'd9408, 16'd25200, 16'd26192, 16'd64844, 16'd31270, 16'd7782, 16'd32191, 16'd5189, 16'd62009, 16'd28547, 16'd24024, 16'd7217, 16'd40718, 16'd50462, 16'd56208, 16'd8022});
	test_expansion(128'h9798b8290d8f6b340c6a6a5cbc5c2c6e, {16'd48523, 16'd56704, 16'd2008, 16'd48536, 16'd44703, 16'd31461, 16'd17107, 16'd17023, 16'd55110, 16'd17876, 16'd35303, 16'd12556, 16'd1262, 16'd40409, 16'd56124, 16'd40291, 16'd9205, 16'd34219, 16'd35883, 16'd55700, 16'd58001, 16'd35461, 16'd13013, 16'd40723, 16'd32005, 16'd37126});
	test_expansion(128'h3f0bfbc76cd43436c27ccb462c75d4c6, {16'd4008, 16'd43736, 16'd62284, 16'd31740, 16'd28264, 16'd53892, 16'd51376, 16'd45805, 16'd52403, 16'd41177, 16'd15755, 16'd16315, 16'd34040, 16'd41156, 16'd36713, 16'd8805, 16'd38082, 16'd39556, 16'd10999, 16'd34598, 16'd53853, 16'd46759, 16'd41286, 16'd18842, 16'd45030, 16'd35063});
	test_expansion(128'h739696b1b80cb54d71fd62fb03d4ac9e, {16'd27790, 16'd30279, 16'd3800, 16'd40775, 16'd34261, 16'd61056, 16'd32816, 16'd18093, 16'd34486, 16'd35098, 16'd55509, 16'd43456, 16'd20061, 16'd48034, 16'd42505, 16'd39588, 16'd19057, 16'd48456, 16'd5857, 16'd48607, 16'd16651, 16'd18333, 16'd39741, 16'd50711, 16'd24200, 16'd27547});
	test_expansion(128'h38eaae268513c69145ee42b26d4b1226, {16'd26757, 16'd58610, 16'd48050, 16'd55924, 16'd50082, 16'd42393, 16'd35707, 16'd11278, 16'd24584, 16'd38591, 16'd5750, 16'd111, 16'd32873, 16'd35185, 16'd26875, 16'd63642, 16'd33307, 16'd6854, 16'd53154, 16'd26312, 16'd12168, 16'd30800, 16'd17328, 16'd24331, 16'd17875, 16'd25653});
	test_expansion(128'hcd3843692edfd4b298d3fb864993414d, {16'd32733, 16'd61009, 16'd37713, 16'd52008, 16'd14591, 16'd62434, 16'd1915, 16'd6036, 16'd3882, 16'd17187, 16'd31578, 16'd37708, 16'd13595, 16'd33090, 16'd62709, 16'd27178, 16'd5077, 16'd14626, 16'd53448, 16'd7318, 16'd23800, 16'd30110, 16'd41697, 16'd59273, 16'd808, 16'd63947});
	test_expansion(128'h9b8039077e085c4515381d0c11f120d6, {16'd53022, 16'd44438, 16'd56667, 16'd23129, 16'd63435, 16'd48663, 16'd53040, 16'd36959, 16'd63373, 16'd45580, 16'd38202, 16'd25891, 16'd809, 16'd24183, 16'd51539, 16'd28761, 16'd42621, 16'd30387, 16'd64599, 16'd36837, 16'd6095, 16'd10450, 16'd6908, 16'd30065, 16'd5752, 16'd41555});
	test_expansion(128'hb3f7c8dee7124daa8996d335be0e970b, {16'd49081, 16'd26444, 16'd49515, 16'd29138, 16'd20037, 16'd22465, 16'd17668, 16'd51722, 16'd63107, 16'd62697, 16'd1650, 16'd10763, 16'd37113, 16'd25428, 16'd4115, 16'd56723, 16'd45192, 16'd30385, 16'd23876, 16'd34198, 16'd34606, 16'd37889, 16'd18639, 16'd6650, 16'd16381, 16'd63444});
	test_expansion(128'hc458de191c6d8c9e8e0794651eb6d348, {16'd2828, 16'd43252, 16'd56463, 16'd20585, 16'd45231, 16'd62451, 16'd41203, 16'd26891, 16'd26177, 16'd43271, 16'd59857, 16'd17395, 16'd24336, 16'd39656, 16'd5970, 16'd57455, 16'd11965, 16'd34432, 16'd9060, 16'd51913, 16'd61805, 16'd47335, 16'd4103, 16'd52648, 16'd7268, 16'd2935});
	test_expansion(128'ha8033a171d057f623ea0ec134ec2b482, {16'd33143, 16'd16889, 16'd4956, 16'd31435, 16'd56852, 16'd19456, 16'd15670, 16'd5569, 16'd50040, 16'd30613, 16'd31801, 16'd57616, 16'd57658, 16'd43895, 16'd5854, 16'd13259, 16'd27341, 16'd36854, 16'd63299, 16'd65047, 16'd441, 16'd57444, 16'd40497, 16'd45828, 16'd33045, 16'd11164});
	test_expansion(128'hff112c6a6f22789af9e4da1e599f8556, {16'd63798, 16'd49886, 16'd43265, 16'd58204, 16'd61251, 16'd41691, 16'd6653, 16'd12361, 16'd16957, 16'd56607, 16'd35150, 16'd5349, 16'd65340, 16'd54878, 16'd61672, 16'd45800, 16'd57348, 16'd47304, 16'd50692, 16'd17965, 16'd53638, 16'd20309, 16'd63746, 16'd60867, 16'd18361, 16'd63433});
	test_expansion(128'h2f53a4043e5f78b1c9f1d4f594f0fd07, {16'd104, 16'd2878, 16'd2, 16'd65280, 16'd14784, 16'd7181, 16'd781, 16'd62734, 16'd31207, 16'd24792, 16'd36320, 16'd16032, 16'd531, 16'd57324, 16'd33611, 16'd19702, 16'd58147, 16'd51600, 16'd61460, 16'd53464, 16'd40233, 16'd62428, 16'd38764, 16'd33739, 16'd13415, 16'd26726});
	test_expansion(128'hf2ea7d9dce4f867c98b8bd051c57cd6c, {16'd43606, 16'd13050, 16'd61692, 16'd42529, 16'd19846, 16'd47743, 16'd43486, 16'd58001, 16'd27480, 16'd62306, 16'd11657, 16'd32004, 16'd49490, 16'd42643, 16'd32621, 16'd25499, 16'd54187, 16'd24171, 16'd20887, 16'd56133, 16'd2992, 16'd23990, 16'd57612, 16'd41393, 16'd48611, 16'd54406});
	test_expansion(128'h8f6d886f8a5c4c0519ad28b3054776e7, {16'd17364, 16'd55205, 16'd10901, 16'd42673, 16'd38920, 16'd39659, 16'd55147, 16'd39755, 16'd10366, 16'd21669, 16'd50299, 16'd25462, 16'd3392, 16'd29519, 16'd40312, 16'd19183, 16'd18729, 16'd34151, 16'd50061, 16'd36896, 16'd59791, 16'd64996, 16'd50956, 16'd39760, 16'd6402, 16'd35337});
	test_expansion(128'h0fe31a08f7e2e48bf9013aa097916f99, {16'd16523, 16'd60073, 16'd27418, 16'd25810, 16'd13664, 16'd11798, 16'd36799, 16'd53897, 16'd40458, 16'd12942, 16'd15363, 16'd42505, 16'd33504, 16'd17653, 16'd29403, 16'd56981, 16'd14532, 16'd14223, 16'd18025, 16'd11630, 16'd62769, 16'd47121, 16'd37199, 16'd58760, 16'd61429, 16'd9429});
	test_expansion(128'h7d29331e207b2faf0e7775e3a92ba325, {16'd44438, 16'd21437, 16'd9158, 16'd25097, 16'd41402, 16'd42296, 16'd35609, 16'd17385, 16'd27473, 16'd44783, 16'd46723, 16'd59825, 16'd58663, 16'd17431, 16'd44991, 16'd31551, 16'd425, 16'd28559, 16'd40294, 16'd17417, 16'd17498, 16'd44044, 16'd36685, 16'd45483, 16'd38019, 16'd7721});
	test_expansion(128'he791707eab09fb06157dbdb8ce4a72c2, {16'd58528, 16'd23898, 16'd21386, 16'd6049, 16'd50104, 16'd9470, 16'd64870, 16'd13047, 16'd42351, 16'd47787, 16'd4327, 16'd13302, 16'd37531, 16'd5084, 16'd14630, 16'd31072, 16'd18827, 16'd1767, 16'd24913, 16'd6747, 16'd11099, 16'd38864, 16'd39236, 16'd53018, 16'd4575, 16'd56496});
	test_expansion(128'h7439b855e2e814a198dc0fd75496c99a, {16'd22987, 16'd45256, 16'd24873, 16'd46828, 16'd56200, 16'd4481, 16'd20697, 16'd33697, 16'd1033, 16'd8494, 16'd39365, 16'd42539, 16'd48395, 16'd64558, 16'd42801, 16'd46115, 16'd58071, 16'd13161, 16'd13964, 16'd59171, 16'd29387, 16'd35765, 16'd49960, 16'd34293, 16'd40317, 16'd12359});
	test_expansion(128'h4bf1a1c7044e0b9b26354a45bbb7b525, {16'd31599, 16'd5610, 16'd42220, 16'd53708, 16'd55032, 16'd7633, 16'd58624, 16'd57249, 16'd5343, 16'd25617, 16'd34330, 16'd51202, 16'd49894, 16'd44998, 16'd39274, 16'd64829, 16'd21397, 16'd23497, 16'd16683, 16'd20957, 16'd4308, 16'd37016, 16'd52379, 16'd53394, 16'd46742, 16'd22115});
	test_expansion(128'h638270cce458de9fa5083ab9f948aa5f, {16'd6812, 16'd52288, 16'd6685, 16'd20591, 16'd25779, 16'd11837, 16'd48997, 16'd64698, 16'd37306, 16'd30581, 16'd16656, 16'd54383, 16'd49777, 16'd5687, 16'd4370, 16'd56906, 16'd9885, 16'd63087, 16'd45424, 16'd60130, 16'd27190, 16'd7254, 16'd40693, 16'd46565, 16'd20974, 16'd43205});
	test_expansion(128'h0ac21bf3529d8807a7f5aa953adbe19a, {16'd30516, 16'd26490, 16'd63613, 16'd24950, 16'd55024, 16'd62095, 16'd52590, 16'd4178, 16'd12124, 16'd11680, 16'd63250, 16'd32306, 16'd43800, 16'd63425, 16'd2625, 16'd39960, 16'd54898, 16'd63106, 16'd45862, 16'd13474, 16'd5438, 16'd27043, 16'd5441, 16'd21578, 16'd57156, 16'd55901});
	test_expansion(128'h6434128636896715f3b5bcbb9a464849, {16'd44173, 16'd59738, 16'd63792, 16'd3854, 16'd3699, 16'd18435, 16'd58559, 16'd22133, 16'd65345, 16'd48755, 16'd40397, 16'd3296, 16'd47250, 16'd15836, 16'd14266, 16'd63731, 16'd24290, 16'd46264, 16'd45335, 16'd44101, 16'd56974, 16'd50264, 16'd25456, 16'd59933, 16'd37247, 16'd37898});
	test_expansion(128'h1b57364d87215241326fa0474144ce7c, {16'd31813, 16'd18373, 16'd33166, 16'd57657, 16'd63489, 16'd47134, 16'd29923, 16'd5867, 16'd51001, 16'd20867, 16'd52524, 16'd32291, 16'd11099, 16'd27177, 16'd13130, 16'd48012, 16'd44625, 16'd43780, 16'd53374, 16'd9785, 16'd19692, 16'd22217, 16'd50706, 16'd57292, 16'd46526, 16'd53512});
	test_expansion(128'h3f54fa071ed310c6f81aa3d1d0e53dfc, {16'd527, 16'd62755, 16'd29278, 16'd28433, 16'd60777, 16'd19349, 16'd40620, 16'd31271, 16'd679, 16'd54410, 16'd13978, 16'd41704, 16'd29777, 16'd33534, 16'd43003, 16'd8270, 16'd6234, 16'd53957, 16'd60659, 16'd64876, 16'd20960, 16'd65493, 16'd24320, 16'd65155, 16'd50915, 16'd24259});
	test_expansion(128'h564f53843516369e7620d1dbdb2c7851, {16'd46827, 16'd52707, 16'd4839, 16'd50565, 16'd33555, 16'd27636, 16'd24676, 16'd58558, 16'd59407, 16'd59835, 16'd46939, 16'd19668, 16'd36103, 16'd42912, 16'd44262, 16'd55711, 16'd59337, 16'd17565, 16'd32883, 16'd48966, 16'd48725, 16'd30564, 16'd9383, 16'd64326, 16'd45862, 16'd25332});
	test_expansion(128'h6c237b2f986d33217f169cd81c54277e, {16'd1521, 16'd41437, 16'd51879, 16'd62428, 16'd49411, 16'd64883, 16'd44473, 16'd32216, 16'd19147, 16'd33952, 16'd17792, 16'd61063, 16'd42607, 16'd15976, 16'd15417, 16'd9714, 16'd20832, 16'd39642, 16'd33375, 16'd37186, 16'd50484, 16'd5537, 16'd32210, 16'd37621, 16'd41806, 16'd44113});
	test_expansion(128'h8c37d8f36048cc2b46e28d6391f1e883, {16'd45216, 16'd42161, 16'd45967, 16'd61122, 16'd60209, 16'd12143, 16'd31378, 16'd3961, 16'd3958, 16'd2470, 16'd30402, 16'd63442, 16'd18900, 16'd25785, 16'd13697, 16'd23713, 16'd64916, 16'd30857, 16'd745, 16'd12655, 16'd12824, 16'd17995, 16'd13245, 16'd3534, 16'd18751, 16'd4786});
	test_expansion(128'hbd7e571a856a9189463d7955451d789a, {16'd40867, 16'd8808, 16'd53054, 16'd20914, 16'd17911, 16'd48832, 16'd60395, 16'd28853, 16'd2385, 16'd40153, 16'd25091, 16'd41356, 16'd21498, 16'd25984, 16'd34932, 16'd39864, 16'd6820, 16'd11026, 16'd44162, 16'd13469, 16'd40655, 16'd10472, 16'd56841, 16'd31916, 16'd11350, 16'd9335});
	test_expansion(128'he8d44a241621fcc17d1e6e7ad4f4c438, {16'd63571, 16'd61921, 16'd40968, 16'd32253, 16'd25205, 16'd43355, 16'd59459, 16'd328, 16'd52247, 16'd59973, 16'd35503, 16'd26859, 16'd1785, 16'd43174, 16'd9398, 16'd15840, 16'd53734, 16'd30724, 16'd40153, 16'd51371, 16'd54668, 16'd7381, 16'd2607, 16'd8341, 16'd30597, 16'd26646});
	test_expansion(128'h1bdb6f082b165c9931fc266557cbf2eb, {16'd59290, 16'd36055, 16'd15707, 16'd26552, 16'd15132, 16'd37224, 16'd7897, 16'd11382, 16'd40718, 16'd62561, 16'd2847, 16'd31818, 16'd39222, 16'd27847, 16'd2746, 16'd1321, 16'd41307, 16'd31696, 16'd29295, 16'd26496, 16'd64439, 16'd41213, 16'd41696, 16'd58354, 16'd57277, 16'd48839});
	test_expansion(128'hc707fc73562cb581a6e0e7f461c6ef58, {16'd39945, 16'd47537, 16'd8639, 16'd49089, 16'd27596, 16'd52813, 16'd46140, 16'd49165, 16'd26563, 16'd38036, 16'd16735, 16'd6162, 16'd34355, 16'd11760, 16'd58424, 16'd61097, 16'd43824, 16'd7305, 16'd9754, 16'd63737, 16'd1358, 16'd37146, 16'd26115, 16'd5001, 16'd52805, 16'd13324});
	test_expansion(128'had14339b0b7b5ef4b192623e61313291, {16'd42638, 16'd555, 16'd6643, 16'd35687, 16'd35172, 16'd50979, 16'd8563, 16'd48414, 16'd51544, 16'd8657, 16'd62510, 16'd37678, 16'd31901, 16'd36694, 16'd65087, 16'd23432, 16'd58695, 16'd13220, 16'd8008, 16'd8961, 16'd2849, 16'd8859, 16'd7847, 16'd60065, 16'd62974, 16'd12460});
	test_expansion(128'h5bd1404aee517ecbe23d34814ad06571, {16'd2834, 16'd54787, 16'd35433, 16'd29820, 16'd55940, 16'd52498, 16'd61258, 16'd52651, 16'd13504, 16'd10186, 16'd35257, 16'd7362, 16'd59899, 16'd31655, 16'd26083, 16'd3150, 16'd43534, 16'd61009, 16'd8520, 16'd17222, 16'd4481, 16'd59515, 16'd56739, 16'd47375, 16'd16842, 16'd28230});
	test_expansion(128'h3d887935ced932a1590c3fa03dce5739, {16'd64055, 16'd16804, 16'd1810, 16'd15795, 16'd38314, 16'd51707, 16'd14352, 16'd55295, 16'd65220, 16'd11989, 16'd42920, 16'd60472, 16'd60781, 16'd46319, 16'd24683, 16'd58308, 16'd64593, 16'd9370, 16'd31269, 16'd29112, 16'd16740, 16'd24421, 16'd22037, 16'd6860, 16'd16263, 16'd47955});
	test_expansion(128'h90625c3669eb6faf77931bf027e17180, {16'd19007, 16'd36175, 16'd53923, 16'd57002, 16'd42050, 16'd45728, 16'd63320, 16'd49619, 16'd1048, 16'd30047, 16'd62166, 16'd19454, 16'd54621, 16'd17062, 16'd9762, 16'd2847, 16'd24653, 16'd50138, 16'd24973, 16'd2394, 16'd63719, 16'd27654, 16'd11515, 16'd56123, 16'd42285, 16'd53486});
	test_expansion(128'h67ff4a7c2d092622dff30d2418d3b5f9, {16'd41783, 16'd34052, 16'd29535, 16'd36423, 16'd38621, 16'd52842, 16'd986, 16'd43859, 16'd61100, 16'd49425, 16'd40958, 16'd46669, 16'd61891, 16'd2445, 16'd40184, 16'd58739, 16'd27584, 16'd9318, 16'd42542, 16'd14521, 16'd23971, 16'd47810, 16'd16954, 16'd44378, 16'd55330, 16'd40642});
	test_expansion(128'hed3498b328059e77dadf9e601ecfc490, {16'd51969, 16'd31212, 16'd25364, 16'd32232, 16'd41876, 16'd52413, 16'd42962, 16'd34574, 16'd29129, 16'd22416, 16'd54943, 16'd5916, 16'd54367, 16'd7712, 16'd60784, 16'd12166, 16'd19300, 16'd38270, 16'd3801, 16'd13903, 16'd25973, 16'd21454, 16'd190, 16'd42850, 16'd34029, 16'd63259});
	test_expansion(128'h0635fda57e772ed18a6f8504e3d7248e, {16'd34529, 16'd48759, 16'd45483, 16'd33411, 16'd30785, 16'd14679, 16'd821, 16'd40445, 16'd54797, 16'd48944, 16'd22261, 16'd35990, 16'd38043, 16'd6277, 16'd27792, 16'd12731, 16'd41661, 16'd48047, 16'd51266, 16'd46825, 16'd8753, 16'd59642, 16'd64027, 16'd30963, 16'd33863, 16'd18916});
	test_expansion(128'h2055648e222a93d1bcf8d21df69b4db7, {16'd55004, 16'd38481, 16'd13633, 16'd38916, 16'd9706, 16'd45169, 16'd23626, 16'd20173, 16'd24152, 16'd40126, 16'd63, 16'd21588, 16'd25896, 16'd2931, 16'd11782, 16'd13040, 16'd29684, 16'd22371, 16'd46525, 16'd27579, 16'd32176, 16'd52493, 16'd31963, 16'd16770, 16'd56198, 16'd60196});
	test_expansion(128'he0e1f45ccd83106db34f7bef35dd237b, {16'd65347, 16'd14650, 16'd27842, 16'd43227, 16'd24380, 16'd34686, 16'd41089, 16'd44950, 16'd35656, 16'd36934, 16'd44064, 16'd35221, 16'd37341, 16'd44979, 16'd45859, 16'd51314, 16'd42894, 16'd54728, 16'd30988, 16'd58417, 16'd60616, 16'd9342, 16'd13782, 16'd19776, 16'd14425, 16'd19401});
	test_expansion(128'h4d6484f6e80b36584e6f64a18874c9dd, {16'd32848, 16'd3094, 16'd61496, 16'd45744, 16'd3579, 16'd46942, 16'd64789, 16'd25457, 16'd34903, 16'd6543, 16'd7062, 16'd10624, 16'd15448, 16'd21354, 16'd14371, 16'd42490, 16'd32104, 16'd12586, 16'd31146, 16'd55575, 16'd3479, 16'd51123, 16'd62224, 16'd22784, 16'd14626, 16'd3443});
	test_expansion(128'h1b1c99f25e85a7389816cf44ea35d540, {16'd8921, 16'd15655, 16'd44649, 16'd2539, 16'd12046, 16'd36739, 16'd37661, 16'd8201, 16'd51948, 16'd60159, 16'd1694, 16'd34169, 16'd12960, 16'd636, 16'd3112, 16'd35667, 16'd5874, 16'd30964, 16'd58389, 16'd54966, 16'd22157, 16'd14013, 16'd65128, 16'd27554, 16'd4841, 16'd34095});
	test_expansion(128'h9940aabac2e051f8622912e2c4cbb96f, {16'd37181, 16'd30487, 16'd1951, 16'd36970, 16'd63965, 16'd12234, 16'd5722, 16'd18498, 16'd64419, 16'd19147, 16'd55257, 16'd28560, 16'd56471, 16'd29311, 16'd37451, 16'd40805, 16'd18886, 16'd4738, 16'd53682, 16'd19479, 16'd7629, 16'd2528, 16'd2436, 16'd18806, 16'd53607, 16'd15328});
	test_expansion(128'hdc91a48cb4c82d5da102e15ab76258e3, {16'd29184, 16'd51471, 16'd42604, 16'd34497, 16'd40215, 16'd22094, 16'd20880, 16'd11961, 16'd8557, 16'd2463, 16'd36879, 16'd32771, 16'd61816, 16'd32870, 16'd10284, 16'd48635, 16'd8744, 16'd33224, 16'd16275, 16'd48699, 16'd13743, 16'd53488, 16'd61214, 16'd7807, 16'd17768, 16'd53005});
	test_expansion(128'h8fd4deeb1847ab92461e41a6f3010001, {16'd41070, 16'd35371, 16'd4516, 16'd11917, 16'd12335, 16'd35993, 16'd16292, 16'd27865, 16'd32769, 16'd40757, 16'd12008, 16'd39530, 16'd64862, 16'd9967, 16'd42426, 16'd12114, 16'd52088, 16'd45515, 16'd10269, 16'd15609, 16'd33189, 16'd27074, 16'd45740, 16'd41966, 16'd60519, 16'd59513});
	test_expansion(128'hfb84c4491bc60f52491949654f11b969, {16'd5074, 16'd17037, 16'd56652, 16'd25763, 16'd62261, 16'd20654, 16'd42758, 16'd44801, 16'd12469, 16'd18828, 16'd6484, 16'd15787, 16'd6902, 16'd15943, 16'd21994, 16'd49223, 16'd5779, 16'd22833, 16'd44513, 16'd60694, 16'd63762, 16'd51225, 16'd57066, 16'd52281, 16'd64528, 16'd16934});
	test_expansion(128'h9ebe00790ae2c8b0f131adb7d9d8c05d, {16'd25527, 16'd28914, 16'd14345, 16'd43619, 16'd39006, 16'd56891, 16'd25146, 16'd63557, 16'd50221, 16'd284, 16'd19827, 16'd21323, 16'd15864, 16'd24413, 16'd24156, 16'd11559, 16'd36887, 16'd54196, 16'd39136, 16'd15206, 16'd42949, 16'd21724, 16'd28220, 16'd39741, 16'd3550, 16'd3546});
	test_expansion(128'h0fef1bc14ebd834865aa98632c87b046, {16'd12273, 16'd39976, 16'd51031, 16'd43233, 16'd35157, 16'd28986, 16'd32404, 16'd48954, 16'd35221, 16'd55544, 16'd55381, 16'd57555, 16'd31995, 16'd2588, 16'd47711, 16'd35762, 16'd229, 16'd23676, 16'd62438, 16'd27265, 16'd17216, 16'd34849, 16'd42138, 16'd21754, 16'd19057, 16'd55519});
	test_expansion(128'h464787124b2e6a8b905198f281c747f4, {16'd23910, 16'd58485, 16'd20091, 16'd60878, 16'd55381, 16'd17333, 16'd53958, 16'd46370, 16'd38763, 16'd30626, 16'd28639, 16'd11490, 16'd42924, 16'd4789, 16'd30086, 16'd57797, 16'd2737, 16'd21362, 16'd59030, 16'd51200, 16'd43134, 16'd20777, 16'd25812, 16'd50646, 16'd9911, 16'd24599});
	test_expansion(128'h05020a0b2087833244fab02c4af28a30, {16'd21667, 16'd6778, 16'd12430, 16'd5756, 16'd1675, 16'd4347, 16'd47106, 16'd20408, 16'd45008, 16'd61188, 16'd32793, 16'd36693, 16'd26055, 16'd42814, 16'd31345, 16'd48008, 16'd56771, 16'd41995, 16'd46813, 16'd53301, 16'd35604, 16'd11535, 16'd53754, 16'd21655, 16'd48124, 16'd19255});
	test_expansion(128'hd676932da2a515216e47d1bcc0fd8937, {16'd26997, 16'd63221, 16'd32153, 16'd44484, 16'd7927, 16'd62823, 16'd51683, 16'd21547, 16'd5396, 16'd25252, 16'd34074, 16'd37905, 16'd37099, 16'd61647, 16'd61828, 16'd60310, 16'd4912, 16'd22906, 16'd60960, 16'd15640, 16'd6463, 16'd41376, 16'd47677, 16'd52196, 16'd21130, 16'd19749});
	test_expansion(128'h38334cd4dc410a64bcb3a76bd489fec0, {16'd36479, 16'd18592, 16'd21397, 16'd9711, 16'd36773, 16'd35342, 16'd33925, 16'd33392, 16'd51447, 16'd45328, 16'd28783, 16'd15412, 16'd19620, 16'd28286, 16'd60993, 16'd49279, 16'd11633, 16'd26952, 16'd44095, 16'd16869, 16'd60965, 16'd4142, 16'd21129, 16'd34290, 16'd10758, 16'd47642});
	test_expansion(128'h7bbf940fd04b6ad431f451b49b69b6df, {16'd4559, 16'd56062, 16'd48267, 16'd46967, 16'd51524, 16'd28821, 16'd27063, 16'd17800, 16'd34486, 16'd22808, 16'd20749, 16'd5492, 16'd6230, 16'd40460, 16'd41611, 16'd46635, 16'd18490, 16'd1375, 16'd38375, 16'd15367, 16'd57346, 16'd17492, 16'd8500, 16'd3260, 16'd46862, 16'd30255});
	test_expansion(128'h5b51edb5e103323901cb78cbf25c7a90, {16'd49994, 16'd17230, 16'd62291, 16'd20415, 16'd28279, 16'd37975, 16'd14560, 16'd9051, 16'd44966, 16'd26197, 16'd62728, 16'd49362, 16'd61381, 16'd56812, 16'd44941, 16'd45620, 16'd17497, 16'd50896, 16'd30787, 16'd55604, 16'd48406, 16'd11919, 16'd226, 16'd3437, 16'd27729, 16'd35595});
	test_expansion(128'h1027745b3e9f0cc8be5f493b9a4b713a, {16'd1892, 16'd8401, 16'd38687, 16'd52484, 16'd33806, 16'd38105, 16'd10603, 16'd11150, 16'd55005, 16'd7964, 16'd47854, 16'd11794, 16'd8614, 16'd61117, 16'd60009, 16'd41364, 16'd19023, 16'd64509, 16'd41470, 16'd546, 16'd63380, 16'd41866, 16'd63716, 16'd11040, 16'd17286, 16'd55547});
	test_expansion(128'hf6096142d38f52a7e42f9068a9c21b9f, {16'd43437, 16'd8327, 16'd42514, 16'd53061, 16'd9144, 16'd57424, 16'd20342, 16'd60867, 16'd64354, 16'd29232, 16'd38659, 16'd9247, 16'd13423, 16'd30107, 16'd60715, 16'd49049, 16'd12217, 16'd49151, 16'd39935, 16'd28166, 16'd12837, 16'd6590, 16'd33825, 16'd18269, 16'd46181, 16'd17986});
	test_expansion(128'hf763ce99a270d10cf9350761d14b5731, {16'd50210, 16'd55235, 16'd27261, 16'd58213, 16'd64964, 16'd25425, 16'd39626, 16'd27232, 16'd38260, 16'd1535, 16'd9586, 16'd56273, 16'd39004, 16'd11201, 16'd45088, 16'd26309, 16'd14026, 16'd52888, 16'd64725, 16'd10810, 16'd36375, 16'd58200, 16'd42155, 16'd3141, 16'd30653, 16'd49764});
	test_expansion(128'h563152481117e525555a0f40d4ff7e7a, {16'd60100, 16'd56797, 16'd45071, 16'd34281, 16'd31264, 16'd18364, 16'd48605, 16'd47210, 16'd22530, 16'd62484, 16'd15228, 16'd34731, 16'd51863, 16'd40999, 16'd27877, 16'd30131, 16'd51938, 16'd3094, 16'd21980, 16'd54167, 16'd53988, 16'd11937, 16'd31053, 16'd52321, 16'd23720, 16'd19491});
	test_expansion(128'h5a4275899e9a38a42bc4571e6337582e, {16'd34628, 16'd4253, 16'd36016, 16'd65344, 16'd36045, 16'd29948, 16'd23594, 16'd26177, 16'd54972, 16'd34496, 16'd6089, 16'd36183, 16'd17968, 16'd27734, 16'd4447, 16'd5748, 16'd41850, 16'd63288, 16'd55029, 16'd11646, 16'd63735, 16'd43976, 16'd39551, 16'd1413, 16'd54733, 16'd4544});
	test_expansion(128'ha58153b5fbe93aa4063772d44eeaf1d3, {16'd8334, 16'd7889, 16'd60507, 16'd11082, 16'd43493, 16'd56937, 16'd44057, 16'd11049, 16'd11300, 16'd14460, 16'd48028, 16'd15809, 16'd45720, 16'd17529, 16'd59242, 16'd57717, 16'd33213, 16'd56789, 16'd55578, 16'd33200, 16'd18846, 16'd57376, 16'd27317, 16'd15009, 16'd51050, 16'd55203});
	test_expansion(128'h54af930c3033e7ccafb591009c1bc4c2, {16'd45558, 16'd57880, 16'd22554, 16'd43164, 16'd28105, 16'd25437, 16'd38821, 16'd44993, 16'd12018, 16'd55934, 16'd43607, 16'd55701, 16'd26213, 16'd52072, 16'd54887, 16'd20092, 16'd25003, 16'd24334, 16'd19992, 16'd51531, 16'd23544, 16'd39469, 16'd64116, 16'd863, 16'd40873, 16'd4610});
	test_expansion(128'h989dfb0bb38beb0c1bf7faf6dd168f3e, {16'd28342, 16'd34888, 16'd47783, 16'd16101, 16'd14331, 16'd36218, 16'd39512, 16'd17177, 16'd36333, 16'd15983, 16'd32802, 16'd61004, 16'd3116, 16'd33961, 16'd21932, 16'd63399, 16'd12014, 16'd29088, 16'd51387, 16'd55031, 16'd65527, 16'd45062, 16'd27968, 16'd45374, 16'd21233, 16'd6304});
	test_expansion(128'h312626342f78fb6a09bd2d4488b9fa37, {16'd42508, 16'd30875, 16'd62201, 16'd62642, 16'd25357, 16'd47863, 16'd12235, 16'd557, 16'd61067, 16'd5824, 16'd6841, 16'd16851, 16'd17587, 16'd62694, 16'd34489, 16'd32473, 16'd18210, 16'd9338, 16'd56454, 16'd55191, 16'd62498, 16'd45911, 16'd24467, 16'd34018, 16'd46519, 16'd59899});
	test_expansion(128'hff6bd6664f84c3b7b4c03562ce0e87b4, {16'd34399, 16'd62458, 16'd48994, 16'd34696, 16'd38115, 16'd54694, 16'd38840, 16'd19327, 16'd3511, 16'd54682, 16'd35466, 16'd46406, 16'd52411, 16'd4450, 16'd38475, 16'd16047, 16'd42633, 16'd35283, 16'd8974, 16'd6631, 16'd13546, 16'd24875, 16'd59365, 16'd55441, 16'd16749, 16'd61666});
	test_expansion(128'h57b8eb9506c4dc503b4e252ffba3a371, {16'd33207, 16'd51227, 16'd61982, 16'd55294, 16'd57271, 16'd3545, 16'd46087, 16'd43155, 16'd43826, 16'd38288, 16'd50653, 16'd46735, 16'd39247, 16'd11147, 16'd53529, 16'd48802, 16'd39862, 16'd48661, 16'd43382, 16'd59970, 16'd9107, 16'd43603, 16'd51777, 16'd62728, 16'd14327, 16'd17074});
	test_expansion(128'had5948ba0c15eed2dc512b6da3e7e36d, {16'd61644, 16'd33817, 16'd26638, 16'd53242, 16'd49341, 16'd17752, 16'd65027, 16'd44215, 16'd51360, 16'd10703, 16'd45251, 16'd1914, 16'd13862, 16'd16078, 16'd51654, 16'd45089, 16'd49263, 16'd12870, 16'd38424, 16'd62300, 16'd6434, 16'd64106, 16'd136, 16'd5047, 16'd34752, 16'd8130});
	test_expansion(128'h839cf0801d21cb251896e8f77977004f, {16'd41221, 16'd22207, 16'd64352, 16'd46295, 16'd5534, 16'd21785, 16'd16917, 16'd17590, 16'd34515, 16'd36175, 16'd47033, 16'd56873, 16'd40815, 16'd20206, 16'd33299, 16'd47938, 16'd60351, 16'd24300, 16'd65238, 16'd8254, 16'd53576, 16'd30860, 16'd20443, 16'd30760, 16'd54476, 16'd186});
	test_expansion(128'had24e8fd8b42336f74b0347b557b322d, {16'd49276, 16'd26550, 16'd7509, 16'd18684, 16'd30326, 16'd1561, 16'd29715, 16'd15408, 16'd444, 16'd39553, 16'd10540, 16'd4069, 16'd22095, 16'd23191, 16'd18294, 16'd29040, 16'd58809, 16'd12322, 16'd24357, 16'd54405, 16'd62129, 16'd2721, 16'd58283, 16'd58090, 16'd919, 16'd13165});
	test_expansion(128'hffb0d17f53b88b581b8432a40db91f5d, {16'd61835, 16'd56299, 16'd57999, 16'd4258, 16'd60991, 16'd52982, 16'd52946, 16'd37966, 16'd49206, 16'd45529, 16'd47617, 16'd18955, 16'd22963, 16'd20437, 16'd9877, 16'd28845, 16'd41038, 16'd30538, 16'd42078, 16'd60138, 16'd11276, 16'd64494, 16'd52924, 16'd30680, 16'd43754, 16'd252});
	test_expansion(128'hddab167bca123d8908e3349bda5837d6, {16'd6508, 16'd45156, 16'd14814, 16'd976, 16'd65232, 16'd29441, 16'd6844, 16'd12970, 16'd9517, 16'd64421, 16'd51682, 16'd64245, 16'd32569, 16'd4991, 16'd1845, 16'd57860, 16'd16013, 16'd6734, 16'd63855, 16'd18394, 16'd18330, 16'd3001, 16'd25680, 16'd12384, 16'd15614, 16'd46012});
	test_expansion(128'hd7fbef0a5b09090cff73c8379d3d9629, {16'd12465, 16'd1849, 16'd45751, 16'd55083, 16'd5595, 16'd55241, 16'd25798, 16'd61092, 16'd17219, 16'd48117, 16'd36464, 16'd55704, 16'd44374, 16'd17206, 16'd39503, 16'd55351, 16'd14890, 16'd43562, 16'd27424, 16'd32637, 16'd46446, 16'd8595, 16'd19273, 16'd52195, 16'd56366, 16'd46893});
	test_expansion(128'h97a6f2df246af7e2fab485bdbab2fd3a, {16'd14778, 16'd43216, 16'd64111, 16'd41157, 16'd22848, 16'd48607, 16'd54238, 16'd36591, 16'd7175, 16'd43549, 16'd1841, 16'd42955, 16'd53001, 16'd58610, 16'd6212, 16'd63469, 16'd55223, 16'd53258, 16'd23720, 16'd64390, 16'd4090, 16'd3849, 16'd34071, 16'd8439, 16'd14044, 16'd46388});
	test_expansion(128'hdc3739ed5211495b0cc0772d644e8c71, {16'd43444, 16'd24628, 16'd30455, 16'd17443, 16'd8911, 16'd33541, 16'd10246, 16'd30594, 16'd33183, 16'd46958, 16'd6054, 16'd43119, 16'd64299, 16'd57324, 16'd7872, 16'd27382, 16'd44366, 16'd60865, 16'd4831, 16'd53704, 16'd33563, 16'd3832, 16'd51354, 16'd28399, 16'd45152, 16'd45705});
	test_expansion(128'h6f3647c55a0eed061cf590bfd758d24e, {16'd63815, 16'd4712, 16'd51932, 16'd61447, 16'd33500, 16'd42779, 16'd64443, 16'd55988, 16'd41307, 16'd33955, 16'd46223, 16'd47772, 16'd57980, 16'd56713, 16'd47207, 16'd19661, 16'd18165, 16'd2549, 16'd39795, 16'd43577, 16'd24048, 16'd41226, 16'd52159, 16'd53596, 16'd42625, 16'd56093});
	test_expansion(128'h9ccb40188ca884022d98af84763be1ec, {16'd16215, 16'd5167, 16'd27331, 16'd38282, 16'd20010, 16'd3278, 16'd63921, 16'd4954, 16'd50012, 16'd60475, 16'd45860, 16'd33251, 16'd4993, 16'd36864, 16'd41337, 16'd40391, 16'd48812, 16'd48117, 16'd63165, 16'd34106, 16'd41773, 16'd18451, 16'd48475, 16'd52962, 16'd17937, 16'd43702});
	test_expansion(128'hafc0c04f2eec18c0faf97cbf7878079a, {16'd62894, 16'd18842, 16'd24957, 16'd29096, 16'd21022, 16'd11340, 16'd11105, 16'd51992, 16'd62039, 16'd24702, 16'd29551, 16'd6171, 16'd54349, 16'd15218, 16'd27468, 16'd41271, 16'd18054, 16'd54285, 16'd44959, 16'd49107, 16'd6968, 16'd21955, 16'd17410, 16'd39782, 16'd64437, 16'd56769});
	test_expansion(128'hc14fd7d488f4ee3f0a8fe7d6f8b23432, {16'd46333, 16'd19047, 16'd25568, 16'd27667, 16'd36202, 16'd28705, 16'd35039, 16'd36543, 16'd46652, 16'd60487, 16'd63531, 16'd21275, 16'd3601, 16'd64873, 16'd12184, 16'd54366, 16'd59310, 16'd56647, 16'd56323, 16'd41570, 16'd40929, 16'd59851, 16'd45986, 16'd39357, 16'd32206, 16'd1047});
	test_expansion(128'h7cb49c660a992efc3a45f6b5e9d1e9e1, {16'd64606, 16'd3803, 16'd55352, 16'd22580, 16'd10758, 16'd47394, 16'd60252, 16'd53066, 16'd45547, 16'd22274, 16'd39105, 16'd35333, 16'd28133, 16'd41321, 16'd22218, 16'd20849, 16'd44915, 16'd41479, 16'd46977, 16'd43475, 16'd44725, 16'd15338, 16'd3918, 16'd29718, 16'd46722, 16'd24362});
	test_expansion(128'hce59fbc7d9337a30762636f19788f6a3, {16'd27075, 16'd50642, 16'd38999, 16'd51854, 16'd7266, 16'd27126, 16'd3549, 16'd38427, 16'd27709, 16'd13094, 16'd48721, 16'd57606, 16'd25395, 16'd54216, 16'd48402, 16'd34391, 16'd41594, 16'd36274, 16'd47259, 16'd55360, 16'd47799, 16'd3301, 16'd59516, 16'd40942, 16'd61235, 16'd39377});
	test_expansion(128'h6180ce4fe9253738ff299ddc556602c3, {16'd49249, 16'd50801, 16'd7010, 16'd27212, 16'd40914, 16'd42299, 16'd63267, 16'd53804, 16'd43693, 16'd3949, 16'd43577, 16'd40033, 16'd28546, 16'd14805, 16'd61545, 16'd55089, 16'd49976, 16'd39944, 16'd30124, 16'd62933, 16'd49572, 16'd52591, 16'd1566, 16'd24187, 16'd51994, 16'd4021});
	test_expansion(128'hf55735bb4bbb5da95fbd8a4eb631d5c3, {16'd44244, 16'd34800, 16'd33859, 16'd6916, 16'd47012, 16'd28441, 16'd45714, 16'd12562, 16'd33553, 16'd47637, 16'd51338, 16'd17551, 16'd14970, 16'd59273, 16'd43628, 16'd42555, 16'd25738, 16'd53937, 16'd14240, 16'd31847, 16'd61734, 16'd52272, 16'd59073, 16'd38643, 16'd32422, 16'd35947});
	test_expansion(128'he67146262f43f8f68337e104c2bbc7a9, {16'd23676, 16'd33535, 16'd55862, 16'd37617, 16'd15351, 16'd29944, 16'd49578, 16'd51088, 16'd23168, 16'd64736, 16'd116, 16'd42702, 16'd35533, 16'd61208, 16'd55197, 16'd40218, 16'd21484, 16'd23112, 16'd54861, 16'd60733, 16'd51339, 16'd55117, 16'd21773, 16'd496, 16'd60883, 16'd28304});
	test_expansion(128'h86e759c9e2544328d5dbfa2ecafd711d, {16'd16435, 16'd10366, 16'd1705, 16'd59106, 16'd20829, 16'd23388, 16'd21019, 16'd51836, 16'd15752, 16'd40156, 16'd52513, 16'd43704, 16'd9776, 16'd9161, 16'd4833, 16'd47314, 16'd31402, 16'd13858, 16'd47929, 16'd45566, 16'd17507, 16'd38688, 16'd20816, 16'd55684, 16'd16522, 16'd28048});
	test_expansion(128'h8268b117e221b5cbff870a8fe882e864, {16'd59524, 16'd6428, 16'd27934, 16'd35193, 16'd39841, 16'd6680, 16'd4919, 16'd29438, 16'd34528, 16'd20582, 16'd41010, 16'd56180, 16'd2453, 16'd61190, 16'd22784, 16'd3874, 16'd3770, 16'd6048, 16'd20571, 16'd42416, 16'd58342, 16'd46980, 16'd23586, 16'd61292, 16'd47670, 16'd8711});
	test_expansion(128'h3d2da2fd1a3cf992ea341ed391e5a518, {16'd45622, 16'd2468, 16'd29285, 16'd53796, 16'd57413, 16'd53974, 16'd60494, 16'd60117, 16'd43402, 16'd6629, 16'd21322, 16'd3635, 16'd49045, 16'd65164, 16'd63813, 16'd598, 16'd7451, 16'd62033, 16'd19180, 16'd1226, 16'd19745, 16'd26315, 16'd47688, 16'd32127, 16'd27569, 16'd57146});
	test_expansion(128'h4aa6db83caed5862aa7ff750bdef81fc, {16'd61752, 16'd29533, 16'd9869, 16'd17351, 16'd6224, 16'd6894, 16'd33987, 16'd64888, 16'd8635, 16'd49069, 16'd30971, 16'd56764, 16'd28792, 16'd46921, 16'd61795, 16'd56387, 16'd49534, 16'd20227, 16'd19394, 16'd49700, 16'd54062, 16'd136, 16'd33863, 16'd45153, 16'd47890, 16'd14269});
	test_expansion(128'h383d40eb06aba40b9cdcbcbcdf1f9b66, {16'd41509, 16'd29282, 16'd13850, 16'd10561, 16'd46255, 16'd23049, 16'd61362, 16'd50614, 16'd12183, 16'd17540, 16'd41108, 16'd7369, 16'd28924, 16'd42181, 16'd15287, 16'd14640, 16'd51225, 16'd43552, 16'd4793, 16'd13100, 16'd41540, 16'd56072, 16'd30636, 16'd64697, 16'd3790, 16'd39410});
	test_expansion(128'h2a2a63fdbf59ea5b1ed66da5604a25de, {16'd29631, 16'd4832, 16'd18508, 16'd57891, 16'd65413, 16'd8700, 16'd47355, 16'd8408, 16'd11317, 16'd1425, 16'd12288, 16'd37919, 16'd48757, 16'd14493, 16'd36272, 16'd29421, 16'd10171, 16'd48674, 16'd7721, 16'd27467, 16'd21076, 16'd7951, 16'd45550, 16'd8257, 16'd38273, 16'd8710});
	test_expansion(128'hea7d74788161463363127eca7b98522c, {16'd52992, 16'd21996, 16'd51387, 16'd5731, 16'd11590, 16'd38482, 16'd36600, 16'd2131, 16'd48236, 16'd60378, 16'd37174, 16'd29885, 16'd46084, 16'd11062, 16'd44210, 16'd59381, 16'd63301, 16'd1421, 16'd1589, 16'd19167, 16'd2672, 16'd51647, 16'd6486, 16'd28869, 16'd18547, 16'd8579});
	test_expansion(128'hde0f1efa576ebabef9114f295110959f, {16'd60056, 16'd13040, 16'd18604, 16'd62436, 16'd58209, 16'd57185, 16'd58871, 16'd1964, 16'd40988, 16'd25908, 16'd9834, 16'd20400, 16'd17059, 16'd38462, 16'd56095, 16'd17169, 16'd54431, 16'd19149, 16'd5534, 16'd47594, 16'd40841, 16'd10818, 16'd43184, 16'd31194, 16'd13977, 16'd16538});
	test_expansion(128'h7723c2f7fd63e88af91ba8f8ca0d0f36, {16'd63570, 16'd24625, 16'd53787, 16'd10279, 16'd37619, 16'd7591, 16'd9449, 16'd17773, 16'd42757, 16'd23436, 16'd48411, 16'd32596, 16'd50950, 16'd51229, 16'd8308, 16'd59046, 16'd41718, 16'd20654, 16'd16800, 16'd56768, 16'd12609, 16'd27482, 16'd23544, 16'd33707, 16'd18236, 16'd30689});
	test_expansion(128'h6e3fbdfdfeb747d874e841ee2cc9640c, {16'd17563, 16'd52005, 16'd45785, 16'd17684, 16'd31369, 16'd30311, 16'd2333, 16'd3331, 16'd45420, 16'd33583, 16'd6722, 16'd4916, 16'd41265, 16'd28102, 16'd58549, 16'd62110, 16'd8341, 16'd33217, 16'd39361, 16'd43083, 16'd63216, 16'd45356, 16'd33491, 16'd15587, 16'd11386, 16'd4665});
	test_expansion(128'h98a211ab4529e7292613b45e7b75e7f9, {16'd21854, 16'd5259, 16'd18236, 16'd10104, 16'd25122, 16'd62136, 16'd28612, 16'd54249, 16'd61121, 16'd42192, 16'd11731, 16'd7572, 16'd19263, 16'd26430, 16'd2787, 16'd15575, 16'd43839, 16'd26358, 16'd14766, 16'd23047, 16'd52535, 16'd31321, 16'd12903, 16'd2822, 16'd10492, 16'd22503});
	test_expansion(128'he52d4f24465c7595da09e7792df7a6e9, {16'd19442, 16'd58053, 16'd37885, 16'd27862, 16'd25599, 16'd36320, 16'd28103, 16'd27218, 16'd57847, 16'd41814, 16'd13225, 16'd48095, 16'd40764, 16'd36292, 16'd959, 16'd18099, 16'd5648, 16'd1293, 16'd51977, 16'd5434, 16'd37295, 16'd64787, 16'd53880, 16'd23869, 16'd28768, 16'd22685});
	test_expansion(128'h9026391e890fb9ed790bd6a22e067c10, {16'd13243, 16'd61144, 16'd51248, 16'd31714, 16'd20982, 16'd59756, 16'd49402, 16'd57902, 16'd48396, 16'd40874, 16'd29282, 16'd48806, 16'd1926, 16'd63630, 16'd9361, 16'd52925, 16'd14434, 16'd12165, 16'd17363, 16'd50647, 16'd21903, 16'd17423, 16'd62433, 16'd21246, 16'd61869, 16'd13555});
	test_expansion(128'h89d0ddce2ef2434718e8ecc950c56abd, {16'd12636, 16'd59108, 16'd20253, 16'd41060, 16'd54415, 16'd8862, 16'd44407, 16'd20912, 16'd22857, 16'd62480, 16'd41815, 16'd35137, 16'd58150, 16'd12827, 16'd7501, 16'd57262, 16'd61742, 16'd60189, 16'd36410, 16'd35289, 16'd52055, 16'd56369, 16'd21633, 16'd15691, 16'd17400, 16'd59659});
	test_expansion(128'h0001610464d3cf7d9a66aa33b3ce54d7, {16'd24911, 16'd47612, 16'd25257, 16'd41953, 16'd56979, 16'd3470, 16'd19529, 16'd11149, 16'd117, 16'd56135, 16'd11840, 16'd13504, 16'd59770, 16'd1422, 16'd13775, 16'd32745, 16'd2447, 16'd36820, 16'd52575, 16'd47413, 16'd63372, 16'd48324, 16'd36483, 16'd2464, 16'd1705, 16'd52877});
	test_expansion(128'h026684627267f398263493018c5a7a77, {16'd63330, 16'd21655, 16'd15591, 16'd18714, 16'd14368, 16'd43722, 16'd25382, 16'd38103, 16'd21112, 16'd35470, 16'd20818, 16'd37651, 16'd30224, 16'd39313, 16'd7840, 16'd40433, 16'd6670, 16'd35110, 16'd64587, 16'd6513, 16'd5240, 16'd61462, 16'd25094, 16'd49349, 16'd12301, 16'd39639});
	test_expansion(128'hb908feda9f740210cf3e1e8ef01ae72f, {16'd63181, 16'd16049, 16'd24992, 16'd13277, 16'd23254, 16'd30689, 16'd62321, 16'd43152, 16'd62635, 16'd38179, 16'd58212, 16'd41393, 16'd32114, 16'd15770, 16'd7700, 16'd55407, 16'd8600, 16'd3842, 16'd58327, 16'd24586, 16'd41060, 16'd17269, 16'd24594, 16'd56859, 16'd38626, 16'd22864});
	test_expansion(128'h004b02fe6663546aecf4a2171f733f8d, {16'd39646, 16'd58702, 16'd62849, 16'd64995, 16'd36823, 16'd26091, 16'd29707, 16'd25969, 16'd6772, 16'd44264, 16'd18015, 16'd59200, 16'd18112, 16'd51786, 16'd61958, 16'd40808, 16'd8420, 16'd60387, 16'd57587, 16'd41569, 16'd17968, 16'd37443, 16'd2611, 16'd13712, 16'd51278, 16'd45689});
	test_expansion(128'h25f8cce223c49d0c81daeaa208315c6f, {16'd29227, 16'd54145, 16'd20294, 16'd58233, 16'd50940, 16'd19853, 16'd65434, 16'd62442, 16'd23226, 16'd62033, 16'd15514, 16'd45580, 16'd2250, 16'd59639, 16'd13491, 16'd11554, 16'd19742, 16'd13063, 16'd24512, 16'd30143, 16'd19358, 16'd24570, 16'd7272, 16'd61749, 16'd57799, 16'd21221});
	test_expansion(128'hdec8de29f1d736afb2fcb75a90efec92, {16'd59111, 16'd22964, 16'd22243, 16'd23856, 16'd41039, 16'd11011, 16'd27624, 16'd523, 16'd64934, 16'd14703, 16'd32939, 16'd1734, 16'd64851, 16'd5729, 16'd56423, 16'd52224, 16'd47260, 16'd19762, 16'd5861, 16'd19846, 16'd9355, 16'd142, 16'd28114, 16'd12918, 16'd8879, 16'd13894});
	test_expansion(128'h8e3e86e120c2eb0660b1bc1249d09187, {16'd28308, 16'd9194, 16'd51513, 16'd31459, 16'd33013, 16'd30074, 16'd36460, 16'd25655, 16'd42125, 16'd27056, 16'd35185, 16'd9723, 16'd6668, 16'd49156, 16'd10729, 16'd32226, 16'd36782, 16'd3019, 16'd54963, 16'd19897, 16'd46920, 16'd21184, 16'd56267, 16'd22444, 16'd29835, 16'd51485});
	test_expansion(128'hbf87625fc2fca2a2d6c115145a8f489e, {16'd40333, 16'd58613, 16'd16261, 16'd24553, 16'd20505, 16'd56744, 16'd63955, 16'd48742, 16'd3108, 16'd35144, 16'd65050, 16'd7221, 16'd51284, 16'd41979, 16'd38513, 16'd48477, 16'd58093, 16'd53734, 16'd17476, 16'd48041, 16'd27372, 16'd21654, 16'd59306, 16'd46254, 16'd49697, 16'd43086});
	test_expansion(128'h231e24a520e3cce9c3e76a6fbcbecf01, {16'd45932, 16'd24439, 16'd14167, 16'd14669, 16'd14028, 16'd43023, 16'd53416, 16'd51923, 16'd19726, 16'd4088, 16'd61966, 16'd55374, 16'd48325, 16'd58815, 16'd3980, 16'd2603, 16'd45649, 16'd18594, 16'd46810, 16'd24715, 16'd5128, 16'd65239, 16'd64188, 16'd44204, 16'd63092, 16'd18192});
	test_expansion(128'h6fa2ba345b9469702b35fe4b48f2d761, {16'd9264, 16'd5073, 16'd57072, 16'd59495, 16'd14247, 16'd9771, 16'd6049, 16'd35954, 16'd47446, 16'd16749, 16'd35012, 16'd1092, 16'd40206, 16'd36280, 16'd9230, 16'd20393, 16'd61752, 16'd16356, 16'd53053, 16'd42699, 16'd2554, 16'd28088, 16'd22741, 16'd6041, 16'd17360, 16'd36563});
	test_expansion(128'hccae85be7d495f1ed4d3ec12160ac127, {16'd30441, 16'd21903, 16'd20969, 16'd54673, 16'd769, 16'd276, 16'd29637, 16'd35295, 16'd5685, 16'd7863, 16'd31687, 16'd11077, 16'd7175, 16'd53514, 16'd47724, 16'd39720, 16'd37767, 16'd23227, 16'd34345, 16'd62766, 16'd27265, 16'd41961, 16'd29498, 16'd51576, 16'd47067, 16'd10207});
	test_expansion(128'he9570169bbc42a706eafa4b04b15b941, {16'd614, 16'd22741, 16'd15759, 16'd23678, 16'd46923, 16'd36577, 16'd21904, 16'd4871, 16'd50222, 16'd29750, 16'd65508, 16'd61816, 16'd9731, 16'd56085, 16'd64636, 16'd6485, 16'd23983, 16'd54207, 16'd52221, 16'd15734, 16'd3672, 16'd16010, 16'd53559, 16'd38107, 16'd48195, 16'd63647});
	test_expansion(128'h3967031dee77e6267ca76e6c2590d0e5, {16'd39479, 16'd17497, 16'd2717, 16'd9448, 16'd48020, 16'd33983, 16'd58127, 16'd60661, 16'd22733, 16'd28769, 16'd19207, 16'd41472, 16'd47939, 16'd11787, 16'd9587, 16'd27233, 16'd8247, 16'd24897, 16'd57673, 16'd19741, 16'd27470, 16'd7384, 16'd61110, 16'd60267, 16'd5138, 16'd15416});
	test_expansion(128'h0ddd862b321079027a3c597f4dcd2fd6, {16'd27032, 16'd46065, 16'd63217, 16'd3059, 16'd14266, 16'd1341, 16'd45712, 16'd16177, 16'd47432, 16'd19469, 16'd56073, 16'd14301, 16'd30243, 16'd65229, 16'd4322, 16'd55951, 16'd12771, 16'd55878, 16'd9958, 16'd48982, 16'd22758, 16'd10327, 16'd10052, 16'd50461, 16'd50842, 16'd43783});
	test_expansion(128'h131d6a16466215fcfde4cd81809f8c79, {16'd32536, 16'd55700, 16'd11852, 16'd59504, 16'd57484, 16'd46127, 16'd42673, 16'd20086, 16'd40534, 16'd65293, 16'd56096, 16'd56436, 16'd55538, 16'd20874, 16'd56259, 16'd8021, 16'd31878, 16'd50157, 16'd13596, 16'd64902, 16'd13254, 16'd40884, 16'd4763, 16'd62905, 16'd42557, 16'd4673});
	test_expansion(128'ha921a50a6623c85494e32ec4f90dd473, {16'd25269, 16'd30639, 16'd60206, 16'd23410, 16'd22168, 16'd65209, 16'd54441, 16'd5771, 16'd41203, 16'd3601, 16'd30212, 16'd42080, 16'd17182, 16'd42063, 16'd53661, 16'd60707, 16'd1629, 16'd3933, 16'd51731, 16'd39293, 16'd57504, 16'd47948, 16'd14710, 16'd11456, 16'd28981, 16'd54307});
	test_expansion(128'h417c74f967756fe1a9806f55c6fe95c0, {16'd43479, 16'd10771, 16'd18380, 16'd22906, 16'd43470, 16'd57280, 16'd11016, 16'd52502, 16'd47179, 16'd5825, 16'd48307, 16'd58440, 16'd14077, 16'd10093, 16'd62345, 16'd17811, 16'd29542, 16'd40064, 16'd64665, 16'd57429, 16'd47966, 16'd44124, 16'd2778, 16'd31027, 16'd54087, 16'd45946});
	test_expansion(128'h6199cb831c6dba47b21226964d915327, {16'd8748, 16'd3410, 16'd9045, 16'd29160, 16'd19247, 16'd18479, 16'd26983, 16'd1780, 16'd31437, 16'd63647, 16'd25629, 16'd18861, 16'd60297, 16'd36989, 16'd1222, 16'd53821, 16'd42376, 16'd22241, 16'd5381, 16'd56691, 16'd24554, 16'd12789, 16'd60415, 16'd3109, 16'd28856, 16'd13028});
	test_expansion(128'hecf8338461d8696c8e447e2e5762b395, {16'd48328, 16'd19174, 16'd25739, 16'd37719, 16'd33356, 16'd33148, 16'd49214, 16'd15510, 16'd2363, 16'd50804, 16'd23773, 16'd65059, 16'd13696, 16'd1214, 16'd288, 16'd33491, 16'd46052, 16'd58921, 16'd33861, 16'd4938, 16'd9695, 16'd14606, 16'd37722, 16'd60778, 16'd53917, 16'd2310});
	test_expansion(128'h30db2c01d88d67e84da649b3c746044e, {16'd14228, 16'd39219, 16'd28426, 16'd6124, 16'd2670, 16'd13585, 16'd63765, 16'd53323, 16'd54490, 16'd15453, 16'd3362, 16'd52422, 16'd60066, 16'd27698, 16'd55189, 16'd55716, 16'd60621, 16'd35501, 16'd5446, 16'd64707, 16'd19497, 16'd21150, 16'd28737, 16'd41167, 16'd42200, 16'd44513});
	test_expansion(128'h715db537ae9aca80bd3f818f4a5c30ac, {16'd13997, 16'd28766, 16'd17678, 16'd13082, 16'd48795, 16'd43814, 16'd31877, 16'd11315, 16'd16159, 16'd38846, 16'd57704, 16'd52390, 16'd50762, 16'd60137, 16'd4983, 16'd5181, 16'd63919, 16'd36015, 16'd37279, 16'd37577, 16'd34342, 16'd13865, 16'd42439, 16'd19819, 16'd63910, 16'd4395});
	test_expansion(128'h58a75064f56fd1a21a9e433f298e9ab3, {16'd63650, 16'd64479, 16'd1848, 16'd49825, 16'd8664, 16'd2668, 16'd24933, 16'd34895, 16'd18048, 16'd10699, 16'd19929, 16'd21155, 16'd9156, 16'd54913, 16'd6092, 16'd2267, 16'd1616, 16'd31198, 16'd22316, 16'd15896, 16'd48359, 16'd26009, 16'd21578, 16'd13053, 16'd45313, 16'd5814});
	test_expansion(128'h475e65f1190dc54e081e10855ec28f3e, {16'd9730, 16'd49009, 16'd22838, 16'd46714, 16'd31692, 16'd37742, 16'd41839, 16'd46236, 16'd51325, 16'd48937, 16'd15426, 16'd23253, 16'd19905, 16'd39841, 16'd62221, 16'd31103, 16'd27979, 16'd31567, 16'd4516, 16'd7169, 16'd8506, 16'd2442, 16'd19977, 16'd54668, 16'd21177, 16'd32048});
	test_expansion(128'h1fea940892c55130ca7efdb063163ab6, {16'd50591, 16'd42396, 16'd29734, 16'd52741, 16'd13554, 16'd12726, 16'd23003, 16'd2509, 16'd3943, 16'd1241, 16'd34501, 16'd20956, 16'd52376, 16'd3929, 16'd61272, 16'd8612, 16'd17735, 16'd319, 16'd25321, 16'd25552, 16'd33958, 16'd30494, 16'd36942, 16'd56572, 16'd23805, 16'd10616});
	test_expansion(128'hb028e8819f4a0eabd92d4d10c221aea9, {16'd46325, 16'd1076, 16'd46415, 16'd10956, 16'd49004, 16'd45356, 16'd31472, 16'd27676, 16'd24992, 16'd3669, 16'd27060, 16'd11958, 16'd52046, 16'd16713, 16'd1210, 16'd32258, 16'd623, 16'd6408, 16'd64023, 16'd29016, 16'd61797, 16'd14520, 16'd28347, 16'd50522, 16'd23913, 16'd59255});
	test_expansion(128'h9994d56baed6b3f177d0976c10dc5531, {16'd26437, 16'd17117, 16'd380, 16'd63219, 16'd52115, 16'd36075, 16'd46277, 16'd5313, 16'd12992, 16'd33829, 16'd1109, 16'd16132, 16'd41763, 16'd64005, 16'd23898, 16'd37424, 16'd16909, 16'd26230, 16'd4429, 16'd57718, 16'd13505, 16'd33381, 16'd19157, 16'd30641, 16'd11221, 16'd9501});
	test_expansion(128'h0ce4c450ebbff11243f9f9b634f2efe8, {16'd8002, 16'd29124, 16'd33087, 16'd20080, 16'd43087, 16'd29610, 16'd13266, 16'd38465, 16'd53540, 16'd7850, 16'd16069, 16'd48148, 16'd4292, 16'd46257, 16'd32219, 16'd25541, 16'd14261, 16'd9398, 16'd27052, 16'd64497, 16'd6864, 16'd23878, 16'd32575, 16'd53923, 16'd37334, 16'd26893});
	test_expansion(128'h97b5badadf1c3d27cdfd530a3a08da60, {16'd33852, 16'd52631, 16'd29980, 16'd29904, 16'd17379, 16'd63203, 16'd46388, 16'd24073, 16'd35718, 16'd59372, 16'd62264, 16'd12257, 16'd58062, 16'd14299, 16'd8504, 16'd62163, 16'd43103, 16'd289, 16'd50170, 16'd46567, 16'd13691, 16'd44755, 16'd39253, 16'd57126, 16'd59895, 16'd48919});
	test_expansion(128'hd5fe2d95615147bc462be69f7def8c26, {16'd44697, 16'd65474, 16'd55444, 16'd19360, 16'd3138, 16'd41125, 16'd38428, 16'd54959, 16'd15218, 16'd31811, 16'd63139, 16'd41619, 16'd58287, 16'd5816, 16'd9382, 16'd12661, 16'd57149, 16'd24287, 16'd47097, 16'd11990, 16'd45758, 16'd9879, 16'd51599, 16'd18657, 16'd36226, 16'd2168});
	test_expansion(128'h63b7c9220b6f0255fab5fbf2d1ea51a1, {16'd65070, 16'd51215, 16'd46840, 16'd18258, 16'd18305, 16'd42540, 16'd13702, 16'd29283, 16'd32076, 16'd13471, 16'd58811, 16'd23469, 16'd28996, 16'd34708, 16'd13282, 16'd50747, 16'd61619, 16'd6134, 16'd61507, 16'd34706, 16'd51070, 16'd29727, 16'd63819, 16'd44720, 16'd53905, 16'd17074});
	test_expansion(128'h1010189faa7ff13902921a43bec1971a, {16'd10222, 16'd643, 16'd4740, 16'd35888, 16'd37180, 16'd10321, 16'd60342, 16'd33186, 16'd9592, 16'd48434, 16'd23875, 16'd47690, 16'd52425, 16'd7084, 16'd27422, 16'd47267, 16'd58715, 16'd18245, 16'd24769, 16'd49285, 16'd12845, 16'd47889, 16'd12048, 16'd58603, 16'd14126, 16'd15035});
	test_expansion(128'h0756d578cbb7483fa9d38970411d1139, {16'd26625, 16'd59571, 16'd35975, 16'd52716, 16'd24604, 16'd32019, 16'd49365, 16'd54690, 16'd21109, 16'd35756, 16'd11763, 16'd51804, 16'd39460, 16'd62164, 16'd22987, 16'd62988, 16'd26950, 16'd13631, 16'd15820, 16'd52808, 16'd19392, 16'd51613, 16'd18764, 16'd26538, 16'd61384, 16'd47492});
	test_expansion(128'h990286de511780014b725f4e50204d8b, {16'd4473, 16'd4906, 16'd34849, 16'd27379, 16'd20182, 16'd30516, 16'd58644, 16'd29315, 16'd10161, 16'd34406, 16'd16458, 16'd7780, 16'd27353, 16'd39144, 16'd13475, 16'd39380, 16'd45741, 16'd57051, 16'd59209, 16'd54172, 16'd23794, 16'd65045, 16'd63377, 16'd2296, 16'd2041, 16'd34785});
	test_expansion(128'he2a2f5658ed9a6a6bffd85a16c08593a, {16'd38141, 16'd3837, 16'd9438, 16'd46989, 16'd65243, 16'd954, 16'd4358, 16'd47576, 16'd32121, 16'd19369, 16'd7217, 16'd10826, 16'd31416, 16'd57269, 16'd16051, 16'd59940, 16'd22181, 16'd7958, 16'd19362, 16'd2910, 16'd53704, 16'd53239, 16'd39267, 16'd26278, 16'd62347, 16'd23183});
	test_expansion(128'h53fc96266f9dfcccc847214f549339ac, {16'd44614, 16'd2801, 16'd37326, 16'd1445, 16'd25667, 16'd36314, 16'd19966, 16'd58359, 16'd63995, 16'd24913, 16'd32976, 16'd4433, 16'd2406, 16'd44314, 16'd51995, 16'd39474, 16'd37353, 16'd16107, 16'd63617, 16'd64578, 16'd51816, 16'd3433, 16'd7369, 16'd19785, 16'd20912, 16'd26893});
	test_expansion(128'hc56db69d22a9bd3c419ea17448203f14, {16'd58437, 16'd54166, 16'd1765, 16'd46398, 16'd17478, 16'd60045, 16'd57231, 16'd54416, 16'd32834, 16'd32939, 16'd4140, 16'd54875, 16'd29026, 16'd55219, 16'd64923, 16'd56227, 16'd25766, 16'd23622, 16'd16517, 16'd17719, 16'd61413, 16'd29927, 16'd18403, 16'd34132, 16'd21437, 16'd47040});
	test_expansion(128'h7f8138e858355af848cf942f45ffb50e, {16'd22861, 16'd32262, 16'd45536, 16'd45783, 16'd52105, 16'd3876, 16'd31991, 16'd61905, 16'd24073, 16'd56370, 16'd31760, 16'd46784, 16'd54422, 16'd54471, 16'd8920, 16'd59786, 16'd3948, 16'd7015, 16'd11449, 16'd823, 16'd18331, 16'd38384, 16'd44057, 16'd57962, 16'd47169, 16'd62066});
	test_expansion(128'hcf2060ed42362ad3a7994b02b1921ef7, {16'd46150, 16'd61121, 16'd6193, 16'd9701, 16'd46402, 16'd58797, 16'd6916, 16'd41935, 16'd2716, 16'd7461, 16'd32570, 16'd47820, 16'd48999, 16'd57623, 16'd19462, 16'd39666, 16'd3703, 16'd28277, 16'd33167, 16'd62422, 16'd29130, 16'd62049, 16'd23997, 16'd59982, 16'd19308, 16'd38205});
	test_expansion(128'h8c500254d4a03a5683b2c42a53c272fd, {16'd13657, 16'd22964, 16'd51840, 16'd55530, 16'd50460, 16'd26686, 16'd14711, 16'd34889, 16'd45791, 16'd1385, 16'd22802, 16'd42171, 16'd51215, 16'd59411, 16'd4833, 16'd8205, 16'd34045, 16'd57581, 16'd58460, 16'd29049, 16'd11649, 16'd19547, 16'd16471, 16'd6805, 16'd34614, 16'd8259});
	test_expansion(128'h32c05ea098c000d307858372d4a1f1cd, {16'd57206, 16'd46212, 16'd7267, 16'd53872, 16'd36538, 16'd27843, 16'd11946, 16'd31908, 16'd47587, 16'd30217, 16'd59055, 16'd26897, 16'd36015, 16'd43852, 16'd62512, 16'd8512, 16'd54742, 16'd41575, 16'd20990, 16'd36517, 16'd46753, 16'd45836, 16'd53055, 16'd1852, 16'd4679, 16'd36495});
	test_expansion(128'hcd5b272f5c7fd16c6bace73960ac11bf, {16'd65067, 16'd56662, 16'd4190, 16'd18467, 16'd8506, 16'd16809, 16'd26721, 16'd8214, 16'd59793, 16'd52546, 16'd64676, 16'd20836, 16'd38587, 16'd41492, 16'd21227, 16'd21871, 16'd20567, 16'd38967, 16'd40001, 16'd27384, 16'd31299, 16'd25562, 16'd41127, 16'd47378, 16'd24009, 16'd26847});
	test_expansion(128'hcb391aa72bc3dc7581a710f00713ac76, {16'd26230, 16'd10630, 16'd57012, 16'd27647, 16'd28404, 16'd61681, 16'd15693, 16'd5486, 16'd46669, 16'd57717, 16'd63125, 16'd55490, 16'd48110, 16'd63612, 16'd12278, 16'd37294, 16'd10207, 16'd10495, 16'd63777, 16'd15176, 16'd62019, 16'd35641, 16'd12462, 16'd17291, 16'd48118, 16'd49714});
	test_expansion(128'hcba30a0f808890636f4ad1b9c1770bbf, {16'd35411, 16'd26283, 16'd17275, 16'd62887, 16'd40727, 16'd44531, 16'd40673, 16'd45573, 16'd17529, 16'd14397, 16'd20665, 16'd59426, 16'd54724, 16'd34466, 16'd50565, 16'd63324, 16'd27532, 16'd39447, 16'd26354, 16'd12061, 16'd53918, 16'd33507, 16'd40912, 16'd12388, 16'd25624, 16'd21571});
	test_expansion(128'h7ca88b11006856ece9e9059f8bebf128, {16'd6621, 16'd24676, 16'd60687, 16'd30840, 16'd42033, 16'd41289, 16'd49255, 16'd34295, 16'd60006, 16'd62030, 16'd58308, 16'd21833, 16'd13722, 16'd41101, 16'd15216, 16'd25993, 16'd60755, 16'd4558, 16'd56819, 16'd43152, 16'd29989, 16'd9810, 16'd1704, 16'd61192, 16'd16581, 16'd24931});
	test_expansion(128'ha5b3c657a7db969493572d8743f0385b, {16'd35852, 16'd51408, 16'd6191, 16'd39013, 16'd35443, 16'd18049, 16'd33436, 16'd21775, 16'd43407, 16'd26957, 16'd4796, 16'd36475, 16'd13249, 16'd48687, 16'd17938, 16'd37293, 16'd42139, 16'd49604, 16'd10647, 16'd52963, 16'd48753, 16'd34049, 16'd60353, 16'd26046, 16'd30584, 16'd41545});
	test_expansion(128'hdf14ffa5c69803962cce6cfcaf953b81, {16'd48257, 16'd40380, 16'd22765, 16'd46387, 16'd58300, 16'd17914, 16'd29852, 16'd57152, 16'd3974, 16'd11253, 16'd30722, 16'd37000, 16'd36352, 16'd41229, 16'd6126, 16'd59234, 16'd24314, 16'd12355, 16'd10910, 16'd59485, 16'd20998, 16'd42444, 16'd24892, 16'd53748, 16'd55561, 16'd31900});
	test_expansion(128'hcdcd216a7089ddf636851e28f741f1e1, {16'd10312, 16'd25184, 16'd40270, 16'd11012, 16'd56029, 16'd57424, 16'd36205, 16'd58559, 16'd8961, 16'd8747, 16'd6912, 16'd25738, 16'd17777, 16'd38886, 16'd37822, 16'd49218, 16'd39173, 16'd3007, 16'd31956, 16'd39630, 16'd999, 16'd43544, 16'd35324, 16'd13506, 16'd46107, 16'd39422});
	test_expansion(128'hfc50387560c3b706dd84a2ea5025940a, {16'd14879, 16'd51929, 16'd20178, 16'd35396, 16'd3669, 16'd27874, 16'd626, 16'd24498, 16'd2496, 16'd14586, 16'd24717, 16'd57442, 16'd11590, 16'd21024, 16'd34245, 16'd18092, 16'd30967, 16'd48674, 16'd51109, 16'd18344, 16'd35336, 16'd41361, 16'd36738, 16'd11332, 16'd36444, 16'd17975});
	test_expansion(128'hd3f8aa28a8f89eb970f74ed10a1a794c, {16'd45199, 16'd2688, 16'd37388, 16'd20185, 16'd10370, 16'd29700, 16'd18472, 16'd51979, 16'd62118, 16'd3540, 16'd57315, 16'd28822, 16'd43149, 16'd50351, 16'd13559, 16'd2107, 16'd39141, 16'd33225, 16'd53295, 16'd16110, 16'd25479, 16'd30597, 16'd31526, 16'd53863, 16'd21276, 16'd21731});
	test_expansion(128'hb1f69fbde0b73ed43398fd5c34bf3b99, {16'd47591, 16'd31777, 16'd9600, 16'd64641, 16'd12704, 16'd8213, 16'd58031, 16'd46890, 16'd19248, 16'd46201, 16'd32362, 16'd20038, 16'd64231, 16'd22173, 16'd55614, 16'd55505, 16'd28077, 16'd3398, 16'd16236, 16'd19826, 16'd21261, 16'd49627, 16'd54447, 16'd11456, 16'd41380, 16'd30509});
	test_expansion(128'he2fd9a070f6bc9e15a88e115d0ae0005, {16'd5299, 16'd53830, 16'd19103, 16'd43434, 16'd7785, 16'd3492, 16'd11552, 16'd42804, 16'd16707, 16'd54127, 16'd14450, 16'd25478, 16'd3028, 16'd9306, 16'd19313, 16'd49746, 16'd9253, 16'd16396, 16'd43352, 16'd57447, 16'd16190, 16'd40627, 16'd49302, 16'd48261, 16'd60506, 16'd7559});
	test_expansion(128'habb1784d8aefcaa9f1ef6409753fc93b, {16'd26732, 16'd46734, 16'd20182, 16'd37085, 16'd4536, 16'd18296, 16'd63112, 16'd19342, 16'd38377, 16'd11120, 16'd26098, 16'd55629, 16'd44594, 16'd25411, 16'd43085, 16'd7701, 16'd25275, 16'd12996, 16'd22506, 16'd16392, 16'd47413, 16'd9850, 16'd33105, 16'd2649, 16'd27060, 16'd4444});
	test_expansion(128'h068f6c53bd5e001c17b99ae443142af9, {16'd34250, 16'd7522, 16'd3857, 16'd61909, 16'd43619, 16'd53309, 16'd43887, 16'd31383, 16'd37938, 16'd35436, 16'd48838, 16'd43165, 16'd38561, 16'd61548, 16'd18749, 16'd345, 16'd1743, 16'd61638, 16'd16873, 16'd60653, 16'd62791, 16'd60070, 16'd43003, 16'd6315, 16'd36375, 16'd18595});
	test_expansion(128'h5d9f77fcdcb3a1558c346098729269da, {16'd17183, 16'd25713, 16'd5616, 16'd31937, 16'd11574, 16'd24732, 16'd30655, 16'd63737, 16'd31161, 16'd13548, 16'd47543, 16'd45899, 16'd56041, 16'd61235, 16'd47758, 16'd30479, 16'd33502, 16'd2187, 16'd18237, 16'd43691, 16'd2824, 16'd27426, 16'd28471, 16'd28164, 16'd59342, 16'd1059});
	test_expansion(128'h7a0bf676cac8b2b38e8d06ac893c6f4e, {16'd38839, 16'd20672, 16'd21787, 16'd8376, 16'd6138, 16'd28255, 16'd15272, 16'd57616, 16'd45918, 16'd45696, 16'd26169, 16'd24710, 16'd22200, 16'd32929, 16'd55068, 16'd19293, 16'd25666, 16'd26058, 16'd65505, 16'd31172, 16'd53136, 16'd64962, 16'd6510, 16'd51976, 16'd14439, 16'd20261});
	test_expansion(128'hc0f7e7a2d53c63116fa79d63bfb9b697, {16'd50811, 16'd10433, 16'd47589, 16'd65042, 16'd15181, 16'd49056, 16'd57771, 16'd29834, 16'd46924, 16'd60123, 16'd62937, 16'd41420, 16'd6651, 16'd9533, 16'd54860, 16'd48942, 16'd47737, 16'd55606, 16'd61042, 16'd5626, 16'd6760, 16'd41143, 16'd27354, 16'd64824, 16'd5064, 16'd31349});
	test_expansion(128'hc1aca0ed349fa7b31c1cbf6aa0571a89, {16'd52821, 16'd23211, 16'd37313, 16'd25095, 16'd8384, 16'd9769, 16'd62061, 16'd38108, 16'd27992, 16'd40413, 16'd34480, 16'd64290, 16'd18888, 16'd55836, 16'd63892, 16'd49834, 16'd47573, 16'd32427, 16'd53525, 16'd42748, 16'd24217, 16'd23451, 16'd60538, 16'd17669, 16'd39, 16'd3177});
	test_expansion(128'hf97a182e848cd47a93da65c7a2caa71c, {16'd65245, 16'd20197, 16'd43803, 16'd6703, 16'd14903, 16'd17041, 16'd12906, 16'd53774, 16'd50182, 16'd26081, 16'd63281, 16'd20970, 16'd8894, 16'd14772, 16'd17676, 16'd6881, 16'd24847, 16'd53721, 16'd39655, 16'd10817, 16'd43148, 16'd47703, 16'd25662, 16'd57721, 16'd49903, 16'd43747});
	test_expansion(128'h15f5b3f0d0e379b0b0a8057861217fd4, {16'd9849, 16'd4487, 16'd60484, 16'd31802, 16'd34064, 16'd44592, 16'd65174, 16'd8390, 16'd21751, 16'd54251, 16'd24558, 16'd31799, 16'd658, 16'd16761, 16'd9648, 16'd26263, 16'd13279, 16'd30739, 16'd26810, 16'd10479, 16'd10127, 16'd44435, 16'd38755, 16'd10812, 16'd20098, 16'd13967});
	test_expansion(128'h76a2da31ba23cbeea4e7b7e915863fa5, {16'd18724, 16'd41771, 16'd17938, 16'd58221, 16'd5680, 16'd14627, 16'd39281, 16'd13592, 16'd42246, 16'd231, 16'd19561, 16'd1136, 16'd54029, 16'd49064, 16'd55585, 16'd64354, 16'd39858, 16'd57132, 16'd44157, 16'd38889, 16'd64599, 16'd32308, 16'd64518, 16'd64303, 16'd14133, 16'd34995});
	test_expansion(128'h610d69df6eebd6f8b9f8d67aadf3a03a, {16'd47482, 16'd6611, 16'd34049, 16'd7397, 16'd36397, 16'd15271, 16'd45748, 16'd58945, 16'd17908, 16'd5664, 16'd8508, 16'd45402, 16'd58626, 16'd53309, 16'd57484, 16'd16057, 16'd40199, 16'd58757, 16'd20093, 16'd63829, 16'd40672, 16'd38563, 16'd1862, 16'd63573, 16'd41005, 16'd47926});
	test_expansion(128'hf3d62394b0dcc6c489940befb47e0df1, {16'd60957, 16'd1281, 16'd24314, 16'd63413, 16'd10385, 16'd33838, 16'd4512, 16'd34451, 16'd51758, 16'd36143, 16'd47606, 16'd63102, 16'd38446, 16'd21316, 16'd46445, 16'd42499, 16'd17629, 16'd602, 16'd10479, 16'd20732, 16'd17069, 16'd27738, 16'd55182, 16'd49580, 16'd21699, 16'd35098});
	test_expansion(128'h7b1165fe861e984ab4fd426e5f5480cc, {16'd7500, 16'd19869, 16'd45831, 16'd50714, 16'd11934, 16'd39727, 16'd45950, 16'd43091, 16'd5986, 16'd47923, 16'd769, 16'd20405, 16'd37780, 16'd35380, 16'd10946, 16'd59374, 16'd32573, 16'd21531, 16'd60555, 16'd12741, 16'd55725, 16'd25073, 16'd41897, 16'd45853, 16'd5787, 16'd57476});
	test_expansion(128'hefca248e1c1d0844120c095488568ff6, {16'd57020, 16'd60953, 16'd22387, 16'd38379, 16'd57688, 16'd20052, 16'd35298, 16'd38329, 16'd18676, 16'd62924, 16'd10798, 16'd49519, 16'd20704, 16'd12231, 16'd40754, 16'd54368, 16'd49358, 16'd24819, 16'd41409, 16'd16924, 16'd36246, 16'd25897, 16'd32944, 16'd41788, 16'd45434, 16'd8972});
	test_expansion(128'hfedbe14bd215e98bd9dbbbde84fc0d78, {16'd52109, 16'd42155, 16'd9532, 16'd47652, 16'd2663, 16'd17001, 16'd14678, 16'd50292, 16'd30303, 16'd47230, 16'd48633, 16'd17135, 16'd19649, 16'd65189, 16'd58344, 16'd18839, 16'd40658, 16'd41788, 16'd47312, 16'd6083, 16'd54488, 16'd59116, 16'd37105, 16'd42769, 16'd30483, 16'd51724});
	test_expansion(128'h6092bbf229f8d69e4d223f003323b44b, {16'd13331, 16'd24254, 16'd3144, 16'd23253, 16'd61358, 16'd1439, 16'd7305, 16'd48723, 16'd3445, 16'd62024, 16'd6915, 16'd64742, 16'd15130, 16'd48975, 16'd52072, 16'd51424, 16'd13808, 16'd62418, 16'd62855, 16'd49676, 16'd45172, 16'd3835, 16'd30840, 16'd38062, 16'd22097, 16'd33112});
	test_expansion(128'he9625998df9f7faa9787070a99fdad33, {16'd3843, 16'd51222, 16'd34172, 16'd34475, 16'd13428, 16'd61110, 16'd36726, 16'd17139, 16'd6130, 16'd3527, 16'd3178, 16'd33303, 16'd764, 16'd27484, 16'd8202, 16'd348, 16'd53988, 16'd60593, 16'd14160, 16'd58575, 16'd15214, 16'd32617, 16'd34098, 16'd35707, 16'd60460, 16'd43985});
	test_expansion(128'hff1382b899b45486de084e2a1b45a5dd, {16'd60924, 16'd20383, 16'd60041, 16'd58940, 16'd64287, 16'd56235, 16'd34316, 16'd26936, 16'd7657, 16'd62412, 16'd55830, 16'd10627, 16'd11701, 16'd6549, 16'd28931, 16'd15422, 16'd13533, 16'd30383, 16'd6200, 16'd55622, 16'd47455, 16'd50489, 16'd61260, 16'd24523, 16'd4754, 16'd32679});
	test_expansion(128'h04a86aec647f6adae44e9f3afa03c781, {16'd12127, 16'd41921, 16'd47987, 16'd45797, 16'd39917, 16'd16545, 16'd35926, 16'd25633, 16'd3980, 16'd18207, 16'd39082, 16'd34580, 16'd54525, 16'd41892, 16'd1070, 16'd4831, 16'd49644, 16'd23302, 16'd20777, 16'd27335, 16'd13590, 16'd45854, 16'd9054, 16'd40081, 16'd35396, 16'd6655});
	test_expansion(128'h4f3ed4807e9154658392fc818db9b9ae, {16'd5073, 16'd53221, 16'd54117, 16'd25506, 16'd18915, 16'd56567, 16'd40757, 16'd62339, 16'd12907, 16'd35200, 16'd48864, 16'd42340, 16'd37962, 16'd2460, 16'd62093, 16'd39330, 16'd61491, 16'd46045, 16'd61648, 16'd28442, 16'd45459, 16'd52318, 16'd29226, 16'd14092, 16'd64227, 16'd52331});
	test_expansion(128'h58f53e533850cb203ce97796694f2022, {16'd53651, 16'd64544, 16'd7181, 16'd7532, 16'd27158, 16'd61994, 16'd14656, 16'd53235, 16'd33475, 16'd50825, 16'd10206, 16'd57255, 16'd24597, 16'd38387, 16'd61048, 16'd16513, 16'd38521, 16'd15165, 16'd56864, 16'd52157, 16'd46266, 16'd19722, 16'd63902, 16'd26361, 16'd32064, 16'd19951});
	test_expansion(128'h826cf8e8c3cc9934acf6cb5c4ce6e861, {16'd1136, 16'd13439, 16'd35013, 16'd14549, 16'd50737, 16'd34881, 16'd9873, 16'd15554, 16'd40791, 16'd60376, 16'd26168, 16'd14789, 16'd19691, 16'd58558, 16'd21822, 16'd17992, 16'd2602, 16'd32464, 16'd41638, 16'd35282, 16'd34686, 16'd22353, 16'd50822, 16'd28636, 16'd60510, 16'd36995});
	test_expansion(128'h32211febd0e7060a3b1ef9ef6fad9dcc, {16'd20733, 16'd58618, 16'd48179, 16'd39288, 16'd27802, 16'd32773, 16'd43975, 16'd9684, 16'd44560, 16'd43239, 16'd62707, 16'd24406, 16'd63155, 16'd14102, 16'd36603, 16'd48623, 16'd11352, 16'd25653, 16'd60415, 16'd32718, 16'd64290, 16'd12889, 16'd53599, 16'd21891, 16'd30012, 16'd16331});
	test_expansion(128'h9eee8246f29f097694dc6a23db9d0336, {16'd64856, 16'd48030, 16'd52485, 16'd6243, 16'd30407, 16'd57075, 16'd54724, 16'd24224, 16'd42247, 16'd8265, 16'd30280, 16'd53864, 16'd57186, 16'd42888, 16'd57072, 16'd46480, 16'd214, 16'd33051, 16'd19035, 16'd42547, 16'd26026, 16'd31355, 16'd11337, 16'd12400, 16'd34823, 16'd64526});
	test_expansion(128'h371b4a06a10cbf66989346ffab7dca9d, {16'd44488, 16'd8498, 16'd19660, 16'd63208, 16'd33387, 16'd44276, 16'd65362, 16'd13008, 16'd39709, 16'd20420, 16'd48882, 16'd38779, 16'd10012, 16'd57451, 16'd3531, 16'd50556, 16'd15134, 16'd21166, 16'd32762, 16'd10843, 16'd10570, 16'd48170, 16'd21079, 16'd38219, 16'd63815, 16'd61436});
	test_expansion(128'h59378649b64f3262245696508f71c47e, {16'd55491, 16'd50088, 16'd47512, 16'd54456, 16'd64554, 16'd18591, 16'd17326, 16'd48199, 16'd22059, 16'd57536, 16'd64302, 16'd50614, 16'd61756, 16'd9298, 16'd52195, 16'd2949, 16'd61302, 16'd33206, 16'd9851, 16'd6476, 16'd65533, 16'd1531, 16'd3533, 16'd38736, 16'd24022, 16'd42910});
	test_expansion(128'hceedccfd00595bd013437a1853e6197c, {16'd57951, 16'd8844, 16'd43970, 16'd45345, 16'd23677, 16'd28127, 16'd34969, 16'd28892, 16'd61462, 16'd11345, 16'd32064, 16'd19519, 16'd61567, 16'd15230, 16'd33149, 16'd51514, 16'd53722, 16'd21950, 16'd63984, 16'd61252, 16'd831, 16'd14050, 16'd55273, 16'd5613, 16'd26537, 16'd33842});
	test_expansion(128'h7828ad34b52a432c7bcfde7d1fc2726b, {16'd46197, 16'd6464, 16'd54306, 16'd21162, 16'd48560, 16'd19210, 16'd62504, 16'd708, 16'd20179, 16'd58053, 16'd64208, 16'd10106, 16'd26235, 16'd55865, 16'd19220, 16'd42531, 16'd13639, 16'd16982, 16'd51852, 16'd31677, 16'd25557, 16'd48229, 16'd32315, 16'd34894, 16'd46902, 16'd27436});
	test_expansion(128'h54cf5b89c79ce8aa09fa3121565a43d8, {16'd1733, 16'd5203, 16'd23213, 16'd62632, 16'd25263, 16'd26480, 16'd52307, 16'd26484, 16'd25970, 16'd25935, 16'd40792, 16'd39077, 16'd35296, 16'd24864, 16'd43101, 16'd50296, 16'd5818, 16'd63169, 16'd4119, 16'd28437, 16'd13134, 16'd41751, 16'd25574, 16'd44056, 16'd17365, 16'd23629});
	test_expansion(128'hc71dcfdc76ec8c01a428629550c94668, {16'd61327, 16'd52517, 16'd31383, 16'd22792, 16'd53391, 16'd3888, 16'd25553, 16'd24835, 16'd57685, 16'd54822, 16'd57208, 16'd39867, 16'd17650, 16'd14957, 16'd61529, 16'd12227, 16'd32957, 16'd4895, 16'd27241, 16'd45530, 16'd25183, 16'd58852, 16'd15869, 16'd28634, 16'd38729, 16'd11115});
	test_expansion(128'hed10e661fdabef3aaa6d49fcc62d5b20, {16'd44104, 16'd25462, 16'd11581, 16'd51787, 16'd63070, 16'd32310, 16'd63337, 16'd827, 16'd37929, 16'd38018, 16'd61761, 16'd55073, 16'd23539, 16'd60940, 16'd62104, 16'd44473, 16'd29816, 16'd55198, 16'd50123, 16'd29606, 16'd11971, 16'd14352, 16'd18004, 16'd57140, 16'd33713, 16'd48137});
	test_expansion(128'h1e16c08076eb4b376803a34dc43d5e3a, {16'd36432, 16'd64275, 16'd53225, 16'd8350, 16'd44819, 16'd3359, 16'd9305, 16'd62517, 16'd3390, 16'd64105, 16'd16074, 16'd27495, 16'd2521, 16'd26094, 16'd50974, 16'd24539, 16'd9944, 16'd53033, 16'd31049, 16'd2806, 16'd30228, 16'd271, 16'd28278, 16'd35188, 16'd37704, 16'd63811});
	test_expansion(128'h42ef0051f1bf7de640e0fb8f5295970c, {16'd21244, 16'd22814, 16'd34159, 16'd19101, 16'd17609, 16'd60308, 16'd59788, 16'd32872, 16'd38616, 16'd37115, 16'd19959, 16'd31600, 16'd2830, 16'd17922, 16'd3015, 16'd15076, 16'd57078, 16'd17361, 16'd24877, 16'd38275, 16'd40453, 16'd57381, 16'd45754, 16'd8345, 16'd49502, 16'd60750});
	test_expansion(128'h67c16e87a0dc97da0e462ed787b81cfd, {16'd60559, 16'd64094, 16'd30659, 16'd23859, 16'd33531, 16'd11459, 16'd34842, 16'd63142, 16'd53038, 16'd57663, 16'd30115, 16'd24877, 16'd63072, 16'd30919, 16'd37182, 16'd53539, 16'd54493, 16'd55661, 16'd29831, 16'd47460, 16'd46917, 16'd44067, 16'd30591, 16'd48639, 16'd37417, 16'd55847});
	test_expansion(128'hcdef32acd73c87e0468e17d06321fead, {16'd2387, 16'd12284, 16'd50740, 16'd41457, 16'd64447, 16'd19993, 16'd15514, 16'd38681, 16'd42152, 16'd32045, 16'd8155, 16'd34629, 16'd56159, 16'd36653, 16'd26732, 16'd31265, 16'd21769, 16'd38504, 16'd33813, 16'd42491, 16'd48002, 16'd818, 16'd9168, 16'd7647, 16'd47947, 16'd50181});
	test_expansion(128'h516dd56236509e43b458316d16469a9a, {16'd20155, 16'd31720, 16'd45362, 16'd58518, 16'd9601, 16'd27651, 16'd2687, 16'd44490, 16'd23028, 16'd36943, 16'd53995, 16'd51193, 16'd57995, 16'd21970, 16'd50124, 16'd4598, 16'd40410, 16'd12425, 16'd16141, 16'd46683, 16'd8665, 16'd9, 16'd38596, 16'd11170, 16'd60658, 16'd59313});
	test_expansion(128'h39b03ad047ab82d08157654281f12afa, {16'd33232, 16'd32310, 16'd8940, 16'd65329, 16'd21640, 16'd50047, 16'd31241, 16'd49093, 16'd24338, 16'd16149, 16'd43409, 16'd36905, 16'd59338, 16'd47221, 16'd27858, 16'd26984, 16'd37696, 16'd56432, 16'd55381, 16'd21595, 16'd39655, 16'd36275, 16'd49394, 16'd52604, 16'd56669, 16'd19392});
	test_expansion(128'ha51803ea6e0f8eefd86c7b5536c6a90f, {16'd12454, 16'd49243, 16'd30668, 16'd15031, 16'd44251, 16'd26238, 16'd14857, 16'd39125, 16'd5729, 16'd48725, 16'd30764, 16'd13511, 16'd13233, 16'd51283, 16'd50633, 16'd9457, 16'd64722, 16'd45823, 16'd34892, 16'd30519, 16'd36431, 16'd49400, 16'd1329, 16'd63933, 16'd44693, 16'd38858});
	test_expansion(128'had23104b3e307c6f197ca94cdea8def1, {16'd54462, 16'd64911, 16'd49920, 16'd52336, 16'd23946, 16'd12488, 16'd9942, 16'd11148, 16'd12575, 16'd22399, 16'd7874, 16'd8659, 16'd4829, 16'd23569, 16'd41792, 16'd47481, 16'd53021, 16'd44554, 16'd26586, 16'd36806, 16'd22957, 16'd61667, 16'd46860, 16'd12687, 16'd23701, 16'd56998});
	test_expansion(128'h8a3c36731aa805119c025ea991e8402f, {16'd16822, 16'd26980, 16'd23227, 16'd27178, 16'd64905, 16'd25614, 16'd61378, 16'd39088, 16'd38453, 16'd59873, 16'd41267, 16'd64527, 16'd56663, 16'd4360, 16'd40973, 16'd64011, 16'd30855, 16'd3372, 16'd45157, 16'd38603, 16'd34522, 16'd28789, 16'd53459, 16'd58562, 16'd62318, 16'd19798});
	test_expansion(128'hc1c4544368da5049c8897562228415bc, {16'd56925, 16'd4311, 16'd15825, 16'd23502, 16'd49241, 16'd31328, 16'd11298, 16'd9660, 16'd26415, 16'd44815, 16'd28540, 16'd59193, 16'd14948, 16'd3826, 16'd14823, 16'd27846, 16'd23959, 16'd41932, 16'd9588, 16'd61845, 16'd56393, 16'd16739, 16'd30695, 16'd5790, 16'd5433, 16'd30698});
	test_expansion(128'h541194181f13ad6b19ec3e0124893988, {16'd31426, 16'd41281, 16'd15338, 16'd6773, 16'd5605, 16'd55064, 16'd30156, 16'd43635, 16'd11604, 16'd23696, 16'd20545, 16'd8591, 16'd15729, 16'd57569, 16'd13414, 16'd65446, 16'd31712, 16'd65242, 16'd25952, 16'd54175, 16'd44045, 16'd50644, 16'd60294, 16'd55152, 16'd35228, 16'd63404});
	test_expansion(128'h430eac7115bdfb2dde3dbee0a0991fb2, {16'd13532, 16'd61389, 16'd46145, 16'd20094, 16'd14437, 16'd47292, 16'd3816, 16'd38711, 16'd42616, 16'd64635, 16'd36918, 16'd16980, 16'd56511, 16'd13480, 16'd38224, 16'd2555, 16'd24777, 16'd14690, 16'd29664, 16'd19587, 16'd44199, 16'd48889, 16'd6127, 16'd21243, 16'd53596, 16'd28325});
	test_expansion(128'hfe9299fbed6602a4fceae6bb970038a9, {16'd24157, 16'd31073, 16'd2846, 16'd2888, 16'd55365, 16'd31259, 16'd9424, 16'd53447, 16'd24600, 16'd3737, 16'd65102, 16'd34726, 16'd53759, 16'd18212, 16'd18757, 16'd40043, 16'd8207, 16'd28184, 16'd27461, 16'd16388, 16'd29883, 16'd11885, 16'd7220, 16'd46186, 16'd59791, 16'd38170});
	test_expansion(128'h3b42eccc66479fc918102e5bcbe32bfc, {16'd2107, 16'd20316, 16'd34181, 16'd35578, 16'd40923, 16'd52277, 16'd21549, 16'd9788, 16'd11644, 16'd48509, 16'd14215, 16'd60797, 16'd45195, 16'd18569, 16'd21283, 16'd48506, 16'd22846, 16'd42196, 16'd9822, 16'd12062, 16'd61859, 16'd14659, 16'd27012, 16'd12536, 16'd38874, 16'd44807});
	test_expansion(128'h54be09a1e6cac093138bae8bf95884a9, {16'd3538, 16'd60375, 16'd30086, 16'd1543, 16'd38300, 16'd33044, 16'd18547, 16'd6698, 16'd13272, 16'd17549, 16'd33548, 16'd52244, 16'd56016, 16'd32341, 16'd54548, 16'd34970, 16'd20858, 16'd35560, 16'd62, 16'd51792, 16'd18994, 16'd14910, 16'd47906, 16'd52854, 16'd33039, 16'd57241});
	test_expansion(128'h6130b891673b8b35db3dc55b0e62cf17, {16'd28495, 16'd63956, 16'd61903, 16'd9337, 16'd52840, 16'd45411, 16'd13651, 16'd43479, 16'd17676, 16'd59160, 16'd64139, 16'd47803, 16'd49896, 16'd25424, 16'd30211, 16'd30898, 16'd43771, 16'd25554, 16'd51653, 16'd55936, 16'd59660, 16'd58657, 16'd8606, 16'd15820, 16'd40691, 16'd49175});
	test_expansion(128'hbdf409a2ebf26a4b305b2702defb3e44, {16'd31844, 16'd56807, 16'd42008, 16'd37345, 16'd20756, 16'd33225, 16'd45265, 16'd42361, 16'd38678, 16'd24938, 16'd47849, 16'd54715, 16'd19964, 16'd401, 16'd6177, 16'd24024, 16'd169, 16'd38471, 16'd58344, 16'd17818, 16'd26713, 16'd16426, 16'd54780, 16'd17451, 16'd19295, 16'd60898});
	test_expansion(128'h1723ed1d055516507dd58dbc01b345f6, {16'd24216, 16'd36532, 16'd2368, 16'd56270, 16'd49899, 16'd26418, 16'd50372, 16'd6773, 16'd26886, 16'd26679, 16'd51490, 16'd40823, 16'd17200, 16'd13390, 16'd14415, 16'd63640, 16'd35770, 16'd50466, 16'd18072, 16'd3223, 16'd49521, 16'd61177, 16'd52597, 16'd48855, 16'd5480, 16'd33320});
	test_expansion(128'h090902b37e7655d2d8fd9867d6a2c678, {16'd60839, 16'd41873, 16'd16137, 16'd16281, 16'd33176, 16'd9196, 16'd53184, 16'd21979, 16'd2618, 16'd5215, 16'd15895, 16'd60884, 16'd12937, 16'd12577, 16'd47451, 16'd39161, 16'd15670, 16'd9502, 16'd8992, 16'd4882, 16'd23600, 16'd1795, 16'd3161, 16'd46930, 16'd24291, 16'd42855});
	test_expansion(128'h87fa65927d53ebd6b2d11f498da625ca, {16'd6593, 16'd8484, 16'd1346, 16'd4904, 16'd28869, 16'd23645, 16'd7846, 16'd24788, 16'd54792, 16'd57455, 16'd55199, 16'd55180, 16'd22669, 16'd40926, 16'd4787, 16'd35909, 16'd19884, 16'd30047, 16'd50482, 16'd2691, 16'd20660, 16'd31934, 16'd65281, 16'd42186, 16'd24792, 16'd38427});
	test_expansion(128'ha60c2e1b5812cb4c06729aa06778d0d0, {16'd32084, 16'd21705, 16'd26289, 16'd18734, 16'd3061, 16'd22073, 16'd38058, 16'd37258, 16'd49950, 16'd31030, 16'd19362, 16'd20618, 16'd31214, 16'd18873, 16'd48456, 16'd13978, 16'd42728, 16'd35251, 16'd35253, 16'd9769, 16'd55357, 16'd12525, 16'd56505, 16'd21774, 16'd1543, 16'd35144});
	test_expansion(128'hcd164d5184eb66d14f16d17bf3e574b9, {16'd62656, 16'd26566, 16'd16618, 16'd1770, 16'd64719, 16'd1281, 16'd10149, 16'd31864, 16'd53094, 16'd20438, 16'd64474, 16'd52456, 16'd31647, 16'd51806, 16'd57332, 16'd58356, 16'd29384, 16'd2659, 16'd28844, 16'd5199, 16'd44672, 16'd39427, 16'd10298, 16'd53244, 16'd17862, 16'd44450});
	test_expansion(128'h98c044ca9952dd53d7ffb0cf4a6e9d89, {16'd52407, 16'd8029, 16'd43230, 16'd54258, 16'd33225, 16'd42788, 16'd42847, 16'd45813, 16'd24418, 16'd24558, 16'd60740, 16'd22104, 16'd23144, 16'd43963, 16'd7384, 16'd22160, 16'd34359, 16'd22377, 16'd28713, 16'd53858, 16'd61106, 16'd42405, 16'd19243, 16'd20120, 16'd22000, 16'd12547});
	test_expansion(128'h04d073c1057ed54e27a9be0fa88bcbc8, {16'd1372, 16'd3957, 16'd27210, 16'd27495, 16'd53484, 16'd48029, 16'd2240, 16'd46758, 16'd40307, 16'd25686, 16'd37241, 16'd62426, 16'd48517, 16'd56002, 16'd24510, 16'd63569, 16'd53000, 16'd19619, 16'd58344, 16'd65200, 16'd10716, 16'd12452, 16'd34408, 16'd21924, 16'd9020, 16'd14212});
	test_expansion(128'hb6467907c14b99618a95a4db3d2f7806, {16'd16990, 16'd60882, 16'd33003, 16'd2246, 16'd62272, 16'd62107, 16'd12239, 16'd46198, 16'd53026, 16'd32652, 16'd552, 16'd30905, 16'd22549, 16'd22187, 16'd51641, 16'd62293, 16'd17782, 16'd34331, 16'd27729, 16'd42665, 16'd53314, 16'd17562, 16'd18490, 16'd16706, 16'd45527, 16'd46243});
	test_expansion(128'h83d917ad69d4ae9e3985e0bd74f42dae, {16'd28518, 16'd61803, 16'd1909, 16'd18189, 16'd42467, 16'd22040, 16'd47543, 16'd5366, 16'd45287, 16'd60676, 16'd22658, 16'd64271, 16'd64778, 16'd55309, 16'd44704, 16'd59356, 16'd51464, 16'd16522, 16'd16081, 16'd36370, 16'd45488, 16'd48108, 16'd46011, 16'd40399, 16'd21024, 16'd27820});
	test_expansion(128'h36944a3c3f53607f548e66ade7d0c07b, {16'd53276, 16'd30445, 16'd3196, 16'd51061, 16'd45592, 16'd20452, 16'd56212, 16'd29174, 16'd47613, 16'd25434, 16'd4803, 16'd33376, 16'd48498, 16'd32643, 16'd21138, 16'd48440, 16'd28060, 16'd40985, 16'd33131, 16'd3438, 16'd6296, 16'd55831, 16'd44468, 16'd8817, 16'd18701, 16'd6875});
	test_expansion(128'hfefaee47e17ab891b9b40bacef085b0e, {16'd37533, 16'd52762, 16'd65483, 16'd47461, 16'd15059, 16'd24068, 16'd19281, 16'd37957, 16'd11603, 16'd32400, 16'd39021, 16'd65416, 16'd29689, 16'd7093, 16'd14869, 16'd26864, 16'd280, 16'd49132, 16'd1247, 16'd20628, 16'd1276, 16'd34548, 16'd25273, 16'd50618, 16'd33544, 16'd6389});
	test_expansion(128'h445eeb205f5fec4b60e76873e689befc, {16'd11994, 16'd12465, 16'd42305, 16'd14003, 16'd62694, 16'd34500, 16'd37292, 16'd31540, 16'd43810, 16'd5407, 16'd51136, 16'd11702, 16'd56140, 16'd39624, 16'd1350, 16'd45404, 16'd19390, 16'd51491, 16'd64212, 16'd30660, 16'd14185, 16'd29922, 16'd12046, 16'd44302, 16'd22536, 16'd31706});
	test_expansion(128'h2375e0301d303e301a2a27820c0fa502, {16'd34114, 16'd42942, 16'd55292, 16'd32850, 16'd60314, 16'd56358, 16'd19855, 16'd30949, 16'd30060, 16'd19142, 16'd50304, 16'd43781, 16'd13598, 16'd55308, 16'd41423, 16'd37744, 16'd27074, 16'd28261, 16'd3208, 16'd21086, 16'd45314, 16'd8799, 16'd37770, 16'd2101, 16'd10531, 16'd48193});
	test_expansion(128'hae1d5f0daea210c19da5bc02e067efc3, {16'd28583, 16'd63080, 16'd47672, 16'd25523, 16'd7710, 16'd10365, 16'd27863, 16'd62429, 16'd53728, 16'd29992, 16'd44184, 16'd49191, 16'd41875, 16'd24633, 16'd19810, 16'd55395, 16'd51696, 16'd21519, 16'd22543, 16'd23867, 16'd13901, 16'd467, 16'd18055, 16'd4758, 16'd57911, 16'd7743});
	test_expansion(128'hb5040edfe3d9db5d5dd94caa04ca082e, {16'd48045, 16'd44277, 16'd51353, 16'd15278, 16'd10611, 16'd41524, 16'd52547, 16'd65500, 16'd12382, 16'd5281, 16'd15104, 16'd61052, 16'd14329, 16'd26105, 16'd64935, 16'd52536, 16'd61789, 16'd31879, 16'd43497, 16'd11526, 16'd31005, 16'd17317, 16'd38067, 16'd41118, 16'd57695, 16'd33443});
	test_expansion(128'h78ab7c3a77bf13f405a07ab0dc70adaa, {16'd2663, 16'd62376, 16'd19802, 16'd6484, 16'd61014, 16'd28131, 16'd36563, 16'd4700, 16'd11344, 16'd21109, 16'd37885, 16'd52340, 16'd53024, 16'd58464, 16'd55409, 16'd38045, 16'd28772, 16'd44771, 16'd37770, 16'd7467, 16'd50465, 16'd29474, 16'd61210, 16'd31778, 16'd43234, 16'd46012});
	test_expansion(128'haad1a72945ccdad455a66eafcc9b0644, {16'd29657, 16'd26969, 16'd34120, 16'd7829, 16'd45592, 16'd25321, 16'd54718, 16'd46973, 16'd45820, 16'd18176, 16'd10150, 16'd43601, 16'd61834, 16'd34910, 16'd62641, 16'd4358, 16'd9626, 16'd27572, 16'd2403, 16'd53338, 16'd57716, 16'd40364, 16'd46046, 16'd20401, 16'd37594, 16'd59959});
	test_expansion(128'h8a1dccaf01208d43d00942adb8890e67, {16'd46738, 16'd19820, 16'd49309, 16'd1934, 16'd17772, 16'd15594, 16'd56855, 16'd16352, 16'd21197, 16'd4454, 16'd12950, 16'd7283, 16'd51799, 16'd15639, 16'd18821, 16'd30612, 16'd27594, 16'd18666, 16'd27627, 16'd83, 16'd60624, 16'd30117, 16'd53119, 16'd40319, 16'd50988, 16'd17818});
	test_expansion(128'hcbab7579f498f98728c08b19dd965996, {16'd5818, 16'd65401, 16'd15924, 16'd58054, 16'd23029, 16'd18296, 16'd19275, 16'd43472, 16'd29796, 16'd51263, 16'd19295, 16'd63788, 16'd14511, 16'd39228, 16'd8704, 16'd24634, 16'd57075, 16'd12711, 16'd7283, 16'd36006, 16'd40524, 16'd44875, 16'd5806, 16'd28073, 16'd48841, 16'd48543});
	test_expansion(128'hc220611ea6673414a7af97084a3d174a, {16'd20045, 16'd39033, 16'd22939, 16'd10936, 16'd29089, 16'd993, 16'd5267, 16'd27848, 16'd2780, 16'd2559, 16'd15678, 16'd13512, 16'd37080, 16'd44244, 16'd52924, 16'd18627, 16'd62639, 16'd42795, 16'd9380, 16'd28081, 16'd35237, 16'd45124, 16'd24149, 16'd1208, 16'd14120, 16'd15735});
	test_expansion(128'hb68d01626b698f73e1c57e2c111fc3e2, {16'd52591, 16'd5159, 16'd54658, 16'd20729, 16'd34805, 16'd27974, 16'd3853, 16'd65494, 16'd1348, 16'd437, 16'd4173, 16'd8165, 16'd36354, 16'd49563, 16'd62587, 16'd8053, 16'd64216, 16'd22427, 16'd15606, 16'd2513, 16'd64321, 16'd41188, 16'd20956, 16'd22885, 16'd666, 16'd62782});
	test_expansion(128'hd3c420e41b146f68175017dce16f5ec2, {16'd3051, 16'd30224, 16'd26829, 16'd13099, 16'd31832, 16'd7076, 16'd13713, 16'd45117, 16'd45414, 16'd12154, 16'd25335, 16'd8169, 16'd6420, 16'd37479, 16'd53715, 16'd40594, 16'd31255, 16'd1019, 16'd6164, 16'd17581, 16'd63386, 16'd23174, 16'd3229, 16'd45565, 16'd59117, 16'd21225});
	test_expansion(128'h255cf46788acf17b9450370584de4a2e, {16'd51545, 16'd58673, 16'd61115, 16'd29058, 16'd49356, 16'd52193, 16'd31509, 16'd32817, 16'd21249, 16'd30690, 16'd45688, 16'd15799, 16'd41439, 16'd33199, 16'd3011, 16'd2737, 16'd28712, 16'd41664, 16'd35220, 16'd741, 16'd30239, 16'd39931, 16'd51775, 16'd30789, 16'd43354, 16'd38801});
	test_expansion(128'h4b2796b2088fe19eb2be04722a05da52, {16'd20120, 16'd50651, 16'd44347, 16'd35304, 16'd51550, 16'd7903, 16'd6916, 16'd15746, 16'd7280, 16'd58622, 16'd51391, 16'd48402, 16'd7604, 16'd38338, 16'd25353, 16'd32856, 16'd28046, 16'd14305, 16'd9366, 16'd13890, 16'd46190, 16'd18621, 16'd14396, 16'd24488, 16'd19746, 16'd19698});
	test_expansion(128'h219bb61499a1c2259cb6658a16382c6d, {16'd25905, 16'd23121, 16'd5966, 16'd26436, 16'd28344, 16'd48988, 16'd33367, 16'd58549, 16'd3592, 16'd61255, 16'd54650, 16'd53471, 16'd51425, 16'd8414, 16'd38109, 16'd35377, 16'd23946, 16'd51654, 16'd62400, 16'd62084, 16'd397, 16'd62168, 16'd31397, 16'd5071, 16'd10272, 16'd2443});
	test_expansion(128'hb66849ba0f8d1325545f8fef30429221, {16'd58795, 16'd33959, 16'd372, 16'd39820, 16'd40215, 16'd60682, 16'd25403, 16'd3290, 16'd58296, 16'd25385, 16'd11107, 16'd40879, 16'd54282, 16'd20319, 16'd40746, 16'd23218, 16'd23465, 16'd59639, 16'd60278, 16'd53317, 16'd60209, 16'd10265, 16'd60776, 16'd25644, 16'd56177, 16'd11765});
	test_expansion(128'h05a6ce4282b3beef71416585d8c54ec2, {16'd7642, 16'd22235, 16'd25302, 16'd10100, 16'd45508, 16'd65245, 16'd7187, 16'd7557, 16'd33106, 16'd50878, 16'd48827, 16'd48463, 16'd18582, 16'd34793, 16'd45110, 16'd43688, 16'd30853, 16'd12515, 16'd16779, 16'd14671, 16'd11433, 16'd45610, 16'd23927, 16'd18060, 16'd15876, 16'd31694});
	test_expansion(128'h1e93af2bb6e1fad7d9f46dcbbfd35d16, {16'd64999, 16'd6622, 16'd73, 16'd28719, 16'd45779, 16'd12128, 16'd61455, 16'd14870, 16'd42137, 16'd58804, 16'd12609, 16'd11320, 16'd19447, 16'd50403, 16'd54162, 16'd33195, 16'd4139, 16'd11842, 16'd25103, 16'd65045, 16'd61856, 16'd32916, 16'd36211, 16'd39315, 16'd49228, 16'd39655});
	test_expansion(128'hd0c5514ca93869aab0172dc9fc0830ff, {16'd52612, 16'd32691, 16'd40344, 16'd47660, 16'd6665, 16'd33211, 16'd48164, 16'd24293, 16'd48399, 16'd65003, 16'd16913, 16'd3765, 16'd1980, 16'd64496, 16'd10512, 16'd57321, 16'd11417, 16'd425, 16'd35361, 16'd9851, 16'd37275, 16'd43341, 16'd28581, 16'd38429, 16'd44509, 16'd1594});
	test_expansion(128'hd3b5afd2d7b0a071b177d494da566bc1, {16'd63920, 16'd6217, 16'd20245, 16'd74, 16'd1744, 16'd57215, 16'd37073, 16'd47543, 16'd58204, 16'd52818, 16'd2380, 16'd38502, 16'd59114, 16'd32146, 16'd12370, 16'd48800, 16'd64684, 16'd50625, 16'd6672, 16'd35094, 16'd30488, 16'd17898, 16'd49237, 16'd44694, 16'd63626, 16'd20481});
	test_expansion(128'h627129f45e0c7bede92fbbba136871de, {16'd3706, 16'd34089, 16'd19435, 16'd17808, 16'd35611, 16'd46581, 16'd40699, 16'd8819, 16'd8079, 16'd31675, 16'd46617, 16'd61955, 16'd29089, 16'd21486, 16'd3651, 16'd35160, 16'd44284, 16'd16159, 16'd27719, 16'd47302, 16'd62912, 16'd56865, 16'd40746, 16'd33844, 16'd360, 16'd17279});
	test_expansion(128'hb3a83f509b27f06130d2da1b1352d0ea, {16'd23714, 16'd8230, 16'd21889, 16'd14691, 16'd3941, 16'd56127, 16'd32107, 16'd38421, 16'd34675, 16'd38618, 16'd18923, 16'd4806, 16'd25642, 16'd35116, 16'd54138, 16'd10841, 16'd45645, 16'd49607, 16'd12078, 16'd3270, 16'd37482, 16'd23650, 16'd59352, 16'd16448, 16'd43756, 16'd15369});
	test_expansion(128'h0cd9fd9a21917428ce92f0f62922aca8, {16'd59632, 16'd43665, 16'd21522, 16'd54734, 16'd64902, 16'd45481, 16'd33345, 16'd53029, 16'd46120, 16'd39061, 16'd16122, 16'd61349, 16'd10676, 16'd3508, 16'd18393, 16'd51310, 16'd34410, 16'd12849, 16'd41972, 16'd18313, 16'd26637, 16'd15372, 16'd6814, 16'd49448, 16'd11518, 16'd3894});
	test_expansion(128'h68656a357cb748a6eca9d63a71bf9875, {16'd25190, 16'd19203, 16'd58184, 16'd8659, 16'd63849, 16'd42369, 16'd44136, 16'd17334, 16'd46422, 16'd44740, 16'd58027, 16'd7736, 16'd8502, 16'd20888, 16'd51954, 16'd11575, 16'd53528, 16'd6533, 16'd8431, 16'd50933, 16'd63056, 16'd18689, 16'd18542, 16'd32866, 16'd30258, 16'd56547});
	test_expansion(128'h905d947363cd546adcc7b44ff39b93e5, {16'd13468, 16'd49369, 16'd17446, 16'd10026, 16'd11228, 16'd3995, 16'd27399, 16'd47321, 16'd46531, 16'd16093, 16'd36891, 16'd44521, 16'd43884, 16'd48661, 16'd14983, 16'd3129, 16'd26947, 16'd25411, 16'd58857, 16'd6723, 16'd58317, 16'd42258, 16'd53687, 16'd42915, 16'd59130, 16'd8988});
	test_expansion(128'hb92b07a611eb5375c36752f74dbea183, {16'd4199, 16'd4446, 16'd38698, 16'd39060, 16'd32920, 16'd14489, 16'd9524, 16'd43761, 16'd3427, 16'd49857, 16'd26567, 16'd12490, 16'd11776, 16'd14680, 16'd5443, 16'd55460, 16'd30095, 16'd65532, 16'd19145, 16'd25761, 16'd32135, 16'd37396, 16'd16219, 16'd32310, 16'd26739, 16'd52552});
	test_expansion(128'hfc79129d64f05c911de150a4d09bd603, {16'd58562, 16'd6276, 16'd35548, 16'd53370, 16'd7638, 16'd19387, 16'd37707, 16'd27970, 16'd4472, 16'd955, 16'd8340, 16'd48624, 16'd310, 16'd57522, 16'd56420, 16'd9250, 16'd45970, 16'd49079, 16'd54450, 16'd33366, 16'd24605, 16'd44492, 16'd39426, 16'd19889, 16'd25984, 16'd56342});
	test_expansion(128'h4328a5ab388f536a1d7822e003a24380, {16'd53651, 16'd12277, 16'd52656, 16'd44607, 16'd4064, 16'd34348, 16'd41082, 16'd39422, 16'd26501, 16'd62641, 16'd26315, 16'd30466, 16'd61127, 16'd18675, 16'd2690, 16'd44196, 16'd23671, 16'd53485, 16'd19537, 16'd31860, 16'd32704, 16'd24886, 16'd53798, 16'd21274, 16'd57822, 16'd10659});
	test_expansion(128'h14cc8a268f795a10404194bf4e9f8529, {16'd18438, 16'd10207, 16'd61848, 16'd62125, 16'd41090, 16'd39882, 16'd56318, 16'd58886, 16'd32148, 16'd3188, 16'd33367, 16'd55664, 16'd41669, 16'd58434, 16'd26192, 16'd32284, 16'd21444, 16'd27858, 16'd42125, 16'd20302, 16'd10962, 16'd26278, 16'd59768, 16'd44316, 16'd58498, 16'd53822});
	test_expansion(128'h133c6403b8bdda10688553accc50722a, {16'd11854, 16'd29447, 16'd19977, 16'd27304, 16'd21089, 16'd4194, 16'd33634, 16'd2882, 16'd2816, 16'd52768, 16'd16888, 16'd51683, 16'd57987, 16'd19709, 16'd34653, 16'd32500, 16'd15749, 16'd41603, 16'd26872, 16'd4766, 16'd9058, 16'd625, 16'd36772, 16'd64589, 16'd53316, 16'd42738});
	test_expansion(128'h5a9f76662a0eab10c350f9021cf7392c, {16'd36678, 16'd12733, 16'd38697, 16'd10966, 16'd20687, 16'd52860, 16'd7959, 16'd5107, 16'd55410, 16'd56738, 16'd18493, 16'd2184, 16'd18688, 16'd17589, 16'd22651, 16'd7892, 16'd27142, 16'd47569, 16'd62112, 16'd55057, 16'd20610, 16'd36612, 16'd29346, 16'd34231, 16'd2556, 16'd47696});
	test_expansion(128'ha16f5b61ef37f8eab0f7a885697c1dba, {16'd22390, 16'd12692, 16'd49759, 16'd5110, 16'd14984, 16'd38549, 16'd52050, 16'd10858, 16'd7897, 16'd26178, 16'd27622, 16'd22732, 16'd30182, 16'd16046, 16'd15945, 16'd23406, 16'd50318, 16'd11512, 16'd45332, 16'd1429, 16'd33416, 16'd49831, 16'd32458, 16'd62536, 16'd9852, 16'd20383});
	test_expansion(128'hbf15b641b8d16ca11af4ac2ecfc93124, {16'd9859, 16'd32351, 16'd61018, 16'd63326, 16'd59775, 16'd24690, 16'd24563, 16'd64693, 16'd53698, 16'd56802, 16'd31574, 16'd21265, 16'd12212, 16'd47633, 16'd33229, 16'd63016, 16'd36415, 16'd42874, 16'd17288, 16'd17286, 16'd61120, 16'd31874, 16'd36095, 16'd48439, 16'd34948, 16'd17535});
	test_expansion(128'h110b56f06041aaa81685b4559799c608, {16'd35647, 16'd53100, 16'd10539, 16'd45431, 16'd5101, 16'd64542, 16'd12446, 16'd9970, 16'd1729, 16'd52587, 16'd28527, 16'd2735, 16'd333, 16'd33419, 16'd21252, 16'd38744, 16'd41633, 16'd56647, 16'd49474, 16'd46520, 16'd29417, 16'd21885, 16'd19965, 16'd32566, 16'd30764, 16'd52972});
	test_expansion(128'h5fd395a5d3bd8af28bc8a3baec438a6a, {16'd30046, 16'd37890, 16'd9870, 16'd3982, 16'd13436, 16'd35020, 16'd35535, 16'd5972, 16'd50986, 16'd55312, 16'd62973, 16'd14079, 16'd2196, 16'd6408, 16'd51102, 16'd48437, 16'd19118, 16'd15666, 16'd7466, 16'd1598, 16'd52261, 16'd3191, 16'd7796, 16'd37046, 16'd58732, 16'd26841});
	test_expansion(128'hcff81567740b2212987e63e2e3837ccb, {16'd55682, 16'd8334, 16'd35315, 16'd7691, 16'd37863, 16'd18663, 16'd13406, 16'd20885, 16'd18072, 16'd5040, 16'd25571, 16'd2705, 16'd6683, 16'd60582, 16'd12630, 16'd21924, 16'd37407, 16'd2410, 16'd64210, 16'd14042, 16'd27409, 16'd27412, 16'd35445, 16'd50099, 16'd15793, 16'd9299});
	test_expansion(128'h960d6a05d6048bcac26322637125feb6, {16'd2360, 16'd15284, 16'd50402, 16'd13755, 16'd59435, 16'd49251, 16'd18146, 16'd2045, 16'd51430, 16'd45631, 16'd11714, 16'd10537, 16'd63633, 16'd16464, 16'd14455, 16'd44875, 16'd58105, 16'd63682, 16'd55581, 16'd15592, 16'd43460, 16'd49435, 16'd7263, 16'd51473, 16'd3074, 16'd8096});
	test_expansion(128'h217d768041b6afae8b198ee33bc8abba, {16'd34543, 16'd42012, 16'd50783, 16'd25600, 16'd45247, 16'd46445, 16'd13915, 16'd24634, 16'd37634, 16'd4885, 16'd28171, 16'd34344, 16'd42736, 16'd40613, 16'd5683, 16'd12391, 16'd26800, 16'd29847, 16'd40062, 16'd570, 16'd29938, 16'd51733, 16'd15977, 16'd38596, 16'd18827, 16'd11057});
	test_expansion(128'h651a8d8ffd3a834b3e39aa0b0d7b8e79, {16'd37846, 16'd59716, 16'd34049, 16'd1970, 16'd59265, 16'd18655, 16'd6228, 16'd27388, 16'd46436, 16'd2787, 16'd20185, 16'd21053, 16'd5485, 16'd624, 16'd7419, 16'd9755, 16'd13789, 16'd29809, 16'd9534, 16'd29516, 16'd19051, 16'd39812, 16'd52894, 16'd21110, 16'd29693, 16'd45880});
	test_expansion(128'hfaa6ba0c33e99517014155bb62f24c5d, {16'd35718, 16'd6463, 16'd56688, 16'd18723, 16'd11455, 16'd44817, 16'd31900, 16'd20480, 16'd11031, 16'd43707, 16'd57875, 16'd9275, 16'd16054, 16'd35773, 16'd57117, 16'd47721, 16'd12362, 16'd18813, 16'd26793, 16'd13205, 16'd37103, 16'd42566, 16'd19443, 16'd16359, 16'd11337, 16'd39106});
	test_expansion(128'h3a9f355f506a2a5bf4150c3442304b89, {16'd41339, 16'd5608, 16'd8893, 16'd50061, 16'd22690, 16'd61099, 16'd28814, 16'd45492, 16'd7427, 16'd24861, 16'd5667, 16'd14935, 16'd26355, 16'd25686, 16'd27451, 16'd5608, 16'd62409, 16'd62586, 16'd39527, 16'd55149, 16'd30750, 16'd2954, 16'd5678, 16'd27471, 16'd49604, 16'd47642});
	test_expansion(128'h12ea995253b976a9295f330d2347786f, {16'd55864, 16'd57801, 16'd41400, 16'd5076, 16'd11015, 16'd51159, 16'd56026, 16'd23975, 16'd59803, 16'd55672, 16'd56311, 16'd52181, 16'd30042, 16'd44239, 16'd6507, 16'd33043, 16'd6970, 16'd893, 16'd30536, 16'd32179, 16'd3443, 16'd4664, 16'd28406, 16'd10946, 16'd62871, 16'd19546});
	test_expansion(128'he5d73d59ae246db5a42f735d14fd267e, {16'd61182, 16'd24450, 16'd6996, 16'd33138, 16'd38776, 16'd17167, 16'd11529, 16'd23447, 16'd61617, 16'd42550, 16'd7429, 16'd46988, 16'd56263, 16'd49318, 16'd12241, 16'd40680, 16'd45483, 16'd32570, 16'd49844, 16'd3690, 16'd2848, 16'd15210, 16'd17931, 16'd33793, 16'd2205, 16'd54947});
	test_expansion(128'hd06d2976f3b50b0f93f368848b139da6, {16'd28419, 16'd16927, 16'd39206, 16'd54983, 16'd14303, 16'd27456, 16'd37031, 16'd39369, 16'd11843, 16'd4167, 16'd27277, 16'd44434, 16'd26857, 16'd808, 16'd41553, 16'd29281, 16'd38216, 16'd798, 16'd31320, 16'd55755, 16'd48321, 16'd20384, 16'd40674, 16'd6041, 16'd20679, 16'd45020});
	test_expansion(128'h4a60ab2e2584bc44471d5d95edd1ed36, {16'd26013, 16'd3674, 16'd61742, 16'd52924, 16'd64971, 16'd7220, 16'd36934, 16'd31373, 16'd150, 16'd5452, 16'd64068, 16'd14640, 16'd27853, 16'd34493, 16'd64173, 16'd48473, 16'd46404, 16'd26130, 16'd41160, 16'd36067, 16'd4397, 16'd10487, 16'd14389, 16'd38823, 16'd23110, 16'd4559});
	test_expansion(128'hdfc1563dd988543c7cec1a4ce62eeff9, {16'd26566, 16'd49439, 16'd59319, 16'd30720, 16'd64785, 16'd35198, 16'd52772, 16'd20123, 16'd18230, 16'd9324, 16'd11989, 16'd52632, 16'd39022, 16'd31492, 16'd43650, 16'd44562, 16'd29302, 16'd28642, 16'd46175, 16'd17124, 16'd697, 16'd25037, 16'd4265, 16'd49574, 16'd3944, 16'd47843});
	test_expansion(128'h1cdd85e02a61bb367cb473ac384fb4b1, {16'd21551, 16'd55802, 16'd30071, 16'd52015, 16'd58685, 16'd61609, 16'd35588, 16'd5016, 16'd32171, 16'd30675, 16'd11697, 16'd50322, 16'd29380, 16'd20470, 16'd41919, 16'd48938, 16'd10971, 16'd2750, 16'd35641, 16'd14685, 16'd19165, 16'd23230, 16'd19507, 16'd45390, 16'd46927, 16'd26784});
	test_expansion(128'hd06b7294addd6ae73288934858ea9c87, {16'd39485, 16'd11159, 16'd28203, 16'd62570, 16'd3735, 16'd6463, 16'd24397, 16'd41577, 16'd49160, 16'd7638, 16'd62008, 16'd59891, 16'd36398, 16'd51219, 16'd13276, 16'd53927, 16'd56634, 16'd48833, 16'd47946, 16'd51115, 16'd57354, 16'd28618, 16'd5869, 16'd38957, 16'd22081, 16'd24658});
	test_expansion(128'hbf58da068040af6c80b59c994f15850b, {16'd5853, 16'd50806, 16'd51108, 16'd58396, 16'd58286, 16'd24641, 16'd9774, 16'd30534, 16'd6999, 16'd5365, 16'd61772, 16'd43695, 16'd9680, 16'd1123, 16'd45283, 16'd51405, 16'd15876, 16'd24215, 16'd32423, 16'd36447, 16'd37613, 16'd13736, 16'd13663, 16'd57575, 16'd25283, 16'd45205});
	test_expansion(128'haeaf5cfbfbe7d6d5ea7cbdc2d1a8e926, {16'd5654, 16'd61685, 16'd56052, 16'd15066, 16'd59025, 16'd4678, 16'd43521, 16'd24244, 16'd24679, 16'd30924, 16'd61640, 16'd31323, 16'd29657, 16'd6963, 16'd14476, 16'd52160, 16'd32998, 16'd10016, 16'd29077, 16'd40635, 16'd21176, 16'd52356, 16'd24192, 16'd54267, 16'd58705, 16'd57595});
	test_expansion(128'h102c01cbd816db6c1c7557500254448d, {16'd6565, 16'd40958, 16'd36914, 16'd41815, 16'd25963, 16'd45192, 16'd34778, 16'd22824, 16'd19797, 16'd61576, 16'd44997, 16'd61190, 16'd62230, 16'd19023, 16'd8148, 16'd43802, 16'd22744, 16'd2733, 16'd63685, 16'd62252, 16'd3096, 16'd7177, 16'd19396, 16'd30848, 16'd26002, 16'd54963});
	test_expansion(128'h5896d9b041bd874063396041570678d7, {16'd40444, 16'd62697, 16'd26338, 16'd21772, 16'd27554, 16'd45040, 16'd63006, 16'd9438, 16'd5618, 16'd57664, 16'd12034, 16'd62805, 16'd4123, 16'd22928, 16'd35091, 16'd45816, 16'd59757, 16'd63432, 16'd34938, 16'd17350, 16'd2999, 16'd23750, 16'd13001, 16'd4069, 16'd14615, 16'd24579});
	test_expansion(128'h11f2c1286a1fb1b8206cefa15ad8a26e, {16'd17699, 16'd5984, 16'd57397, 16'd62741, 16'd23589, 16'd7239, 16'd14989, 16'd17809, 16'd54315, 16'd20600, 16'd48501, 16'd11147, 16'd19657, 16'd36546, 16'd24171, 16'd8728, 16'd3564, 16'd986, 16'd62818, 16'd49549, 16'd12772, 16'd38526, 16'd22514, 16'd33494, 16'd8169, 16'd18297});
	test_expansion(128'hb298b040bb63731ecd4733c67327a1e8, {16'd39207, 16'd8528, 16'd11894, 16'd55961, 16'd3189, 16'd47658, 16'd34017, 16'd23737, 16'd3848, 16'd21044, 16'd65239, 16'd63098, 16'd11463, 16'd41589, 16'd63428, 16'd23372, 16'd30401, 16'd13226, 16'd51252, 16'd29565, 16'd59658, 16'd26754, 16'd54047, 16'd16052, 16'd32445, 16'd55923});
	test_expansion(128'h305dab7d61d6afc9be6bc435dd3caa55, {16'd32102, 16'd14725, 16'd16808, 16'd23831, 16'd41975, 16'd51033, 16'd35743, 16'd27077, 16'd30255, 16'd25583, 16'd10120, 16'd39218, 16'd58843, 16'd5918, 16'd2454, 16'd25472, 16'd1672, 16'd52357, 16'd49232, 16'd3445, 16'd133, 16'd31631, 16'd7466, 16'd6480, 16'd19192, 16'd5870});
	test_expansion(128'hce129c4790278f9e70582fe9c792c4d0, {16'd33658, 16'd56730, 16'd50471, 16'd36906, 16'd5291, 16'd30625, 16'd5515, 16'd64335, 16'd50894, 16'd27821, 16'd28507, 16'd33204, 16'd43231, 16'd60225, 16'd17087, 16'd53010, 16'd32030, 16'd12723, 16'd43444, 16'd31865, 16'd51132, 16'd42495, 16'd64225, 16'd13167, 16'd59394, 16'd21349});
	test_expansion(128'h3150431ce1ed5657fe160fa8b55fdfa7, {16'd47877, 16'd61970, 16'd45108, 16'd49954, 16'd31887, 16'd61623, 16'd36919, 16'd31297, 16'd9008, 16'd24717, 16'd28731, 16'd42378, 16'd39021, 16'd57571, 16'd54855, 16'd59317, 16'd50548, 16'd22699, 16'd39596, 16'd13800, 16'd24806, 16'd60423, 16'd47528, 16'd32635, 16'd19429, 16'd59209});
	test_expansion(128'h747afdf1c15b58c6174256980dbad8ff, {16'd22396, 16'd22395, 16'd18496, 16'd20868, 16'd8036, 16'd9510, 16'd40698, 16'd21263, 16'd51470, 16'd35628, 16'd63154, 16'd6859, 16'd5127, 16'd51946, 16'd7454, 16'd16332, 16'd15747, 16'd55573, 16'd27543, 16'd43928, 16'd30485, 16'd5290, 16'd7859, 16'd12124, 16'd19070, 16'd55999});
	test_expansion(128'h35e4ed7861728441eefe8f5ebbc816df, {16'd24794, 16'd4582, 16'd11167, 16'd6231, 16'd54354, 16'd31984, 16'd5593, 16'd26371, 16'd13577, 16'd4983, 16'd19664, 16'd50063, 16'd46116, 16'd6712, 16'd57410, 16'd22159, 16'd42102, 16'd7981, 16'd54365, 16'd5675, 16'd27633, 16'd35188, 16'd38494, 16'd26540, 16'd44119, 16'd43980});
	test_expansion(128'h078b075ea160e31bfe15cc20a6036090, {16'd3854, 16'd45871, 16'd47863, 16'd21873, 16'd9982, 16'd738, 16'd63662, 16'd62840, 16'd968, 16'd43656, 16'd13728, 16'd28557, 16'd30131, 16'd55979, 16'd22891, 16'd63185, 16'd35629, 16'd46045, 16'd16602, 16'd36410, 16'd60917, 16'd25758, 16'd48970, 16'd39191, 16'd35286, 16'd21489});
	test_expansion(128'h466df1d508a5c3a0c77ff0395f2b353d, {16'd22954, 16'd33235, 16'd23029, 16'd33733, 16'd65349, 16'd41126, 16'd54353, 16'd57387, 16'd65404, 16'd58939, 16'd10796, 16'd32051, 16'd53485, 16'd17383, 16'd50021, 16'd25753, 16'd16881, 16'd18605, 16'd45474, 16'd30253, 16'd38769, 16'd4778, 16'd19752, 16'd54005, 16'd4892, 16'd11638});
	test_expansion(128'hff561627bc476209ed17baa0ecd5dcd3, {16'd62258, 16'd62474, 16'd27416, 16'd380, 16'd58651, 16'd61438, 16'd55340, 16'd35568, 16'd56118, 16'd804, 16'd54816, 16'd10293, 16'd5128, 16'd56681, 16'd47878, 16'd31460, 16'd34613, 16'd48886, 16'd58054, 16'd20593, 16'd3760, 16'd61491, 16'd18438, 16'd63615, 16'd37521, 16'd30188});
	test_expansion(128'h0b6ca851f0ef894d89447bd8c5da3743, {16'd35840, 16'd18158, 16'd27010, 16'd30765, 16'd33885, 16'd41780, 16'd36593, 16'd63317, 16'd50306, 16'd40319, 16'd32301, 16'd1859, 16'd59725, 16'd26876, 16'd19045, 16'd18433, 16'd167, 16'd41331, 16'd52196, 16'd17127, 16'd34020, 16'd63662, 16'd22559, 16'd34892, 16'd10022, 16'd22478});
	test_expansion(128'ha957afce60a82db218ff802a25223c3e, {16'd9732, 16'd36791, 16'd13157, 16'd64905, 16'd15180, 16'd176, 16'd2086, 16'd19180, 16'd7210, 16'd17328, 16'd20540, 16'd45622, 16'd62504, 16'd12707, 16'd34681, 16'd25273, 16'd6007, 16'd20547, 16'd64913, 16'd46104, 16'd51289, 16'd59939, 16'd55547, 16'd65380, 16'd27869, 16'd34718});
	test_expansion(128'h945f5f05aabf1c132356b74ff4bbec87, {16'd55147, 16'd53051, 16'd56545, 16'd57775, 16'd40152, 16'd53031, 16'd45731, 16'd5800, 16'd12493, 16'd16758, 16'd30554, 16'd60070, 16'd65093, 16'd22976, 16'd37867, 16'd42638, 16'd47398, 16'd43101, 16'd29792, 16'd12328, 16'd24781, 16'd37442, 16'd37852, 16'd29739, 16'd5307, 16'd6729});
	test_expansion(128'h1aee0e52c3b0eebea9772913f36b0c0c, {16'd63245, 16'd11285, 16'd27876, 16'd62528, 16'd16611, 16'd7531, 16'd15534, 16'd54282, 16'd30705, 16'd6538, 16'd44744, 16'd25609, 16'd62426, 16'd45406, 16'd45693, 16'd38000, 16'd55841, 16'd43141, 16'd23617, 16'd36291, 16'd12177, 16'd18026, 16'd54371, 16'd47480, 16'd61553, 16'd23530});
	test_expansion(128'h1e9ecbdeca320d21bf2859e2fd0dceed, {16'd8153, 16'd64654, 16'd45947, 16'd23398, 16'd30977, 16'd27731, 16'd62127, 16'd41998, 16'd1058, 16'd15586, 16'd21025, 16'd3543, 16'd19846, 16'd17054, 16'd10283, 16'd18524, 16'd33061, 16'd47526, 16'd1807, 16'd8958, 16'd25384, 16'd5955, 16'd23648, 16'd19226, 16'd41668, 16'd12204});
	test_expansion(128'h2f7de7a26c74713b04be8f12d79f561a, {16'd30753, 16'd17890, 16'd62726, 16'd5407, 16'd26251, 16'd23986, 16'd26026, 16'd52939, 16'd13044, 16'd51769, 16'd23797, 16'd39551, 16'd36218, 16'd56943, 16'd26228, 16'd16829, 16'd36954, 16'd19973, 16'd27508, 16'd8748, 16'd48323, 16'd13092, 16'd28071, 16'd21084, 16'd20636, 16'd47624});
	test_expansion(128'hf5b7b1206c50eedaf454fe3e4efd253c, {16'd42404, 16'd9306, 16'd52401, 16'd27988, 16'd6284, 16'd26454, 16'd40575, 16'd6306, 16'd76, 16'd35827, 16'd35002, 16'd14550, 16'd54608, 16'd65001, 16'd3529, 16'd29517, 16'd1910, 16'd1218, 16'd10936, 16'd3204, 16'd4798, 16'd42972, 16'd23792, 16'd56726, 16'd62442, 16'd17489});
	test_expansion(128'h5687a99761465556ef8e4ef2ae9d4f77, {16'd28254, 16'd47909, 16'd7300, 16'd20653, 16'd23013, 16'd10577, 16'd8305, 16'd17672, 16'd12041, 16'd31547, 16'd51920, 16'd35469, 16'd4694, 16'd38701, 16'd46467, 16'd21095, 16'd30870, 16'd39618, 16'd24165, 16'd7922, 16'd37999, 16'd52218, 16'd439, 16'd52257, 16'd58251, 16'd46559});
	test_expansion(128'hbc882fa9e27e39f84ec895bfdb1b379d, {16'd52306, 16'd58361, 16'd4420, 16'd34837, 16'd51874, 16'd60303, 16'd15355, 16'd38160, 16'd27900, 16'd22777, 16'd19263, 16'd38742, 16'd13421, 16'd23911, 16'd56313, 16'd10213, 16'd2824, 16'd11838, 16'd36677, 16'd28635, 16'd52294, 16'd47873, 16'd53176, 16'd32955, 16'd14140, 16'd23367});
	test_expansion(128'ha5b324cca4caff8725979926c194be00, {16'd32843, 16'd23035, 16'd14530, 16'd37543, 16'd13752, 16'd41857, 16'd24118, 16'd3424, 16'd11143, 16'd23706, 16'd8821, 16'd7476, 16'd10788, 16'd24695, 16'd22579, 16'd44496, 16'd63545, 16'd47215, 16'd43214, 16'd15441, 16'd3038, 16'd56594, 16'd31771, 16'd14732, 16'd44797, 16'd16976});
	test_expansion(128'hcb2462a913a6768df9c0dd103e35416d, {16'd8300, 16'd36485, 16'd61147, 16'd3623, 16'd5904, 16'd153, 16'd10724, 16'd36452, 16'd47347, 16'd14836, 16'd50905, 16'd44886, 16'd60582, 16'd12747, 16'd9059, 16'd49426, 16'd55065, 16'd20898, 16'd23435, 16'd42110, 16'd16140, 16'd51502, 16'd36959, 16'd63600, 16'd8748, 16'd1784});
	test_expansion(128'hc7ab65e1060f8970ea1abf158fe6a591, {16'd32114, 16'd36244, 16'd58761, 16'd4667, 16'd35450, 16'd24660, 16'd41786, 16'd13497, 16'd35558, 16'd24017, 16'd18927, 16'd5274, 16'd27733, 16'd61047, 16'd32802, 16'd20123, 16'd5301, 16'd37046, 16'd36371, 16'd16815, 16'd4437, 16'd26625, 16'd3950, 16'd29826, 16'd22371, 16'd46868});
	test_expansion(128'h26fc8372fd8fac60b470063095ba3127, {16'd4069, 16'd23019, 16'd6796, 16'd64322, 16'd63199, 16'd26587, 16'd15809, 16'd6966, 16'd42154, 16'd30306, 16'd61088, 16'd29930, 16'd17954, 16'd16108, 16'd62306, 16'd29380, 16'd51642, 16'd55449, 16'd46407, 16'd48394, 16'd17871, 16'd17440, 16'd56652, 16'd51137, 16'd23162, 16'd50142});
	test_expansion(128'h18412a56ef660f8c50abc0c36b7a6ad6, {16'd37545, 16'd21664, 16'd8505, 16'd25152, 16'd8554, 16'd5515, 16'd18474, 16'd19197, 16'd10145, 16'd6952, 16'd12948, 16'd19875, 16'd52596, 16'd6357, 16'd65439, 16'd15366, 16'd1556, 16'd38660, 16'd13409, 16'd37319, 16'd7384, 16'd53918, 16'd60934, 16'd18387, 16'd44549, 16'd46457});
	test_expansion(128'h0276f9ff215cba078d72b6845b11bfe2, {16'd51060, 16'd36461, 16'd59149, 16'd22433, 16'd56964, 16'd26351, 16'd60427, 16'd48455, 16'd37115, 16'd11605, 16'd40580, 16'd33206, 16'd47315, 16'd52295, 16'd49800, 16'd19954, 16'd56726, 16'd46114, 16'd42662, 16'd28642, 16'd50238, 16'd14939, 16'd12394, 16'd41062, 16'd26283, 16'd42468});
	test_expansion(128'h6be49b824349de7955c09ddf74ec4d0b, {16'd62259, 16'd4261, 16'd54381, 16'd28344, 16'd4210, 16'd22437, 16'd60832, 16'd36861, 16'd55280, 16'd52084, 16'd64869, 16'd41214, 16'd4324, 16'd29715, 16'd15248, 16'd7113, 16'd37600, 16'd3730, 16'd13076, 16'd64281, 16'd25305, 16'd43488, 16'd54067, 16'd39961, 16'd22587, 16'd43787});
	test_expansion(128'ha00b7bb08db857148ecf253cc6f7d690, {16'd39987, 16'd59261, 16'd51992, 16'd28111, 16'd5817, 16'd52652, 16'd58849, 16'd55943, 16'd6635, 16'd49491, 16'd8277, 16'd41272, 16'd16464, 16'd63705, 16'd40505, 16'd38293, 16'd28718, 16'd43348, 16'd31196, 16'd23941, 16'd14485, 16'd40234, 16'd63296, 16'd29232, 16'd17266, 16'd39911});
	test_expansion(128'h8766e7d1406f20f5fca344e7b1701203, {16'd57530, 16'd20526, 16'd26617, 16'd2078, 16'd33193, 16'd52836, 16'd24551, 16'd37718, 16'd46785, 16'd23565, 16'd41215, 16'd16062, 16'd15498, 16'd29734, 16'd32864, 16'd6501, 16'd38867, 16'd63211, 16'd32285, 16'd27303, 16'd44425, 16'd52882, 16'd1376, 16'd27577, 16'd51771, 16'd1903});
	test_expansion(128'h63e381a7bec264a37aeca49d006609ba, {16'd23574, 16'd29420, 16'd38325, 16'd19346, 16'd24667, 16'd63381, 16'd62823, 16'd51127, 16'd52200, 16'd47674, 16'd30600, 16'd12498, 16'd59465, 16'd50030, 16'd28044, 16'd9289, 16'd10294, 16'd59784, 16'd64490, 16'd2325, 16'd28958, 16'd6312, 16'd59284, 16'd21432, 16'd31601, 16'd52650});
	test_expansion(128'h1b5ee6305a6457d493019a40cfa0c4e2, {16'd26746, 16'd63628, 16'd3092, 16'd13392, 16'd33636, 16'd4903, 16'd45726, 16'd4651, 16'd4325, 16'd35891, 16'd26892, 16'd32712, 16'd27050, 16'd26433, 16'd23047, 16'd23613, 16'd39247, 16'd3166, 16'd9894, 16'd42772, 16'd18542, 16'd2068, 16'd4679, 16'd12240, 16'd37392, 16'd2134});
	test_expansion(128'hd86c9f3a14eceac6f292fc346de93647, {16'd35475, 16'd40101, 16'd59553, 16'd58556, 16'd45878, 16'd11686, 16'd60269, 16'd45630, 16'd6603, 16'd7356, 16'd49130, 16'd37480, 16'd31850, 16'd5475, 16'd5909, 16'd9244, 16'd30231, 16'd27755, 16'd22312, 16'd65294, 16'd16525, 16'd22636, 16'd30336, 16'd13994, 16'd5931, 16'd63390});
	test_expansion(128'hb48ac6fa56e029a64eba44365e1a9a09, {16'd33837, 16'd24956, 16'd39201, 16'd11500, 16'd4815, 16'd34391, 16'd35936, 16'd6264, 16'd24847, 16'd14959, 16'd55285, 16'd19825, 16'd12527, 16'd45877, 16'd52858, 16'd35931, 16'd43090, 16'd7261, 16'd42431, 16'd32373, 16'd51594, 16'd2305, 16'd34662, 16'd51210, 16'd5631, 16'd3127});
	test_expansion(128'h9c1bc98e3b8b39ab91115cd6bd5beb5a, {16'd5191, 16'd13387, 16'd28996, 16'd32427, 16'd58110, 16'd19695, 16'd46655, 16'd35335, 16'd64027, 16'd43286, 16'd50874, 16'd65054, 16'd31118, 16'd17691, 16'd29453, 16'd38784, 16'd27874, 16'd49474, 16'd59675, 16'd60234, 16'd56382, 16'd48454, 16'd36598, 16'd10786, 16'd30546, 16'd58651});
	test_expansion(128'h780eab5fbad658afbe5cc25a23df3d71, {16'd59302, 16'd51912, 16'd23910, 16'd64582, 16'd52358, 16'd17743, 16'd4273, 16'd10407, 16'd31208, 16'd51143, 16'd10937, 16'd47688, 16'd9470, 16'd63732, 16'd7401, 16'd22754, 16'd43289, 16'd40178, 16'd49450, 16'd57038, 16'd14483, 16'd63519, 16'd2722, 16'd13501, 16'd58658, 16'd46286});
	test_expansion(128'h37a58538707062a4e72cdd537e9d6d84, {16'd15734, 16'd35666, 16'd7707, 16'd6925, 16'd62426, 16'd12673, 16'd20480, 16'd9009, 16'd51042, 16'd52707, 16'd36659, 16'd31078, 16'd23469, 16'd34236, 16'd11476, 16'd19696, 16'd45959, 16'd65400, 16'd5470, 16'd32816, 16'd64119, 16'd53230, 16'd38346, 16'd52715, 16'd57486, 16'd924});
	test_expansion(128'he5f56d76183424dae9a9740e83ccd912, {16'd46844, 16'd33862, 16'd49692, 16'd5516, 16'd22676, 16'd20142, 16'd34946, 16'd44957, 16'd4286, 16'd41183, 16'd20883, 16'd43592, 16'd50816, 16'd65160, 16'd54362, 16'd1772, 16'd23470, 16'd3245, 16'd26090, 16'd26174, 16'd48411, 16'd42531, 16'd7963, 16'd38106, 16'd5277, 16'd39736});
	test_expansion(128'hff35ec7548c651534abe3b314ad75812, {16'd24428, 16'd41071, 16'd23223, 16'd42035, 16'd11510, 16'd12695, 16'd17115, 16'd48160, 16'd36592, 16'd11264, 16'd12683, 16'd19901, 16'd39068, 16'd17990, 16'd2388, 16'd43075, 16'd25226, 16'd62541, 16'd6133, 16'd5340, 16'd10611, 16'd57104, 16'd12143, 16'd18932, 16'd1291, 16'd64771});
	test_expansion(128'h7fc644da19ebc08f3de2bae1dc93e2d9, {16'd63113, 16'd24830, 16'd44106, 16'd62910, 16'd32126, 16'd18113, 16'd27170, 16'd9106, 16'd16504, 16'd32762, 16'd18782, 16'd28063, 16'd22443, 16'd52184, 16'd4264, 16'd34582, 16'd48360, 16'd54974, 16'd13565, 16'd51235, 16'd17711, 16'd55228, 16'd4239, 16'd34247, 16'd35040, 16'd63678});
	test_expansion(128'h628652b20368ebdfe9a65462618994a8, {16'd10134, 16'd20218, 16'd64885, 16'd12017, 16'd5847, 16'd43341, 16'd34734, 16'd21354, 16'd52434, 16'd31293, 16'd51040, 16'd14703, 16'd18137, 16'd61441, 16'd47513, 16'd535, 16'd34810, 16'd35372, 16'd32951, 16'd4768, 16'd55524, 16'd2678, 16'd24330, 16'd49220, 16'd36098, 16'd55568});
	test_expansion(128'h77fd6166d02430df89ecdd260958e8f8, {16'd4115, 16'd58106, 16'd53537, 16'd52025, 16'd15211, 16'd48825, 16'd3790, 16'd62383, 16'd23462, 16'd36389, 16'd7788, 16'd17927, 16'd129, 16'd56278, 16'd13287, 16'd42856, 16'd38927, 16'd63428, 16'd51328, 16'd55229, 16'd4844, 16'd37831, 16'd19639, 16'd504, 16'd60339, 16'd35892});
	test_expansion(128'h2102a7b4721f1c368b60766a92940a6a, {16'd29042, 16'd51678, 16'd62439, 16'd9346, 16'd51337, 16'd665, 16'd59941, 16'd33413, 16'd32290, 16'd39674, 16'd59474, 16'd5668, 16'd61983, 16'd44497, 16'd31095, 16'd36018, 16'd52308, 16'd14718, 16'd22434, 16'd29082, 16'd12671, 16'd14009, 16'd53322, 16'd30949, 16'd36378, 16'd6186});
	test_expansion(128'hfb250f8ef1b6644b5689963f7ef642f1, {16'd49956, 16'd21085, 16'd60338, 16'd33617, 16'd29126, 16'd27343, 16'd445, 16'd10452, 16'd41897, 16'd12273, 16'd17463, 16'd43629, 16'd2683, 16'd14734, 16'd2200, 16'd14308, 16'd21508, 16'd45751, 16'd16712, 16'd25579, 16'd13263, 16'd15885, 16'd601, 16'd33611, 16'd15845, 16'd5515});
	test_expansion(128'h1cfefec4c14d00f64fee88cc864a218e, {16'd42071, 16'd57946, 16'd53029, 16'd13790, 16'd12800, 16'd59227, 16'd38753, 16'd59403, 16'd27381, 16'd28784, 16'd63314, 16'd21451, 16'd21849, 16'd45934, 16'd11164, 16'd11107, 16'd38353, 16'd15710, 16'd61628, 16'd10055, 16'd7606, 16'd31511, 16'd13328, 16'd49797, 16'd59513, 16'd43230});
	test_expansion(128'hf5ad125b287bfedde2d48aced0b2689d, {16'd35259, 16'd47874, 16'd10175, 16'd58549, 16'd36626, 16'd57773, 16'd55501, 16'd23925, 16'd21748, 16'd26905, 16'd56758, 16'd1116, 16'd10829, 16'd39087, 16'd57412, 16'd19199, 16'd8674, 16'd52935, 16'd61343, 16'd19984, 16'd60396, 16'd33972, 16'd39231, 16'd22546, 16'd38795, 16'd45060});
	test_expansion(128'h3dba9661a219469bb44b6b917ba4aec7, {16'd42342, 16'd1894, 16'd39579, 16'd27903, 16'd32511, 16'd3080, 16'd22604, 16'd25850, 16'd34234, 16'd10857, 16'd60233, 16'd19408, 16'd42553, 16'd37297, 16'd46642, 16'd64928, 16'd28886, 16'd7151, 16'd5910, 16'd53168, 16'd29010, 16'd47001, 16'd9462, 16'd48690, 16'd36310, 16'd48303});
	test_expansion(128'h12a6e39cd851a87b0278faa916ba776f, {16'd51396, 16'd11349, 16'd20135, 16'd15416, 16'd30588, 16'd20241, 16'd53631, 16'd13205, 16'd4709, 16'd33267, 16'd36136, 16'd27609, 16'd15004, 16'd54248, 16'd51953, 16'd11150, 16'd23476, 16'd64124, 16'd26936, 16'd44105, 16'd40381, 16'd53266, 16'd55239, 16'd10025, 16'd2710, 16'd57785});
	test_expansion(128'h765845bf5e3d36fb49ec87cb1aa23188, {16'd62281, 16'd43160, 16'd17595, 16'd51438, 16'd62878, 16'd23077, 16'd15203, 16'd57920, 16'd59801, 16'd535, 16'd56346, 16'd934, 16'd57177, 16'd48132, 16'd56454, 16'd30301, 16'd25443, 16'd45848, 16'd5238, 16'd31397, 16'd59970, 16'd57041, 16'd10563, 16'd34649, 16'd7766, 16'd9311});
	test_expansion(128'he77cc19af9a77df446bbb5f1bdd175ee, {16'd20015, 16'd29376, 16'd3319, 16'd23129, 16'd4531, 16'd59604, 16'd1569, 16'd2638, 16'd59669, 16'd64058, 16'd36973, 16'd14455, 16'd630, 16'd7529, 16'd46951, 16'd42741, 16'd63195, 16'd48544, 16'd12507, 16'd40465, 16'd21735, 16'd28873, 16'd26017, 16'd18633, 16'd33592, 16'd58939});
	test_expansion(128'h66c83ca1cf2e986dddec0221bac60d34, {16'd7010, 16'd59944, 16'd55561, 16'd17696, 16'd18202, 16'd64652, 16'd34940, 16'd48535, 16'd55414, 16'd46901, 16'd33279, 16'd4373, 16'd53946, 16'd35733, 16'd64240, 16'd44874, 16'd30841, 16'd52402, 16'd13956, 16'd9620, 16'd21793, 16'd4605, 16'd57058, 16'd50840, 16'd15478, 16'd21338});
	test_expansion(128'h7d370f48bc2a737d309ac440bdba5515, {16'd37250, 16'd17637, 16'd8072, 16'd23915, 16'd17937, 16'd2663, 16'd3223, 16'd16717, 16'd39616, 16'd45323, 16'd56063, 16'd37830, 16'd556, 16'd24348, 16'd33721, 16'd55189, 16'd33030, 16'd18800, 16'd41582, 16'd16977, 16'd33132, 16'd55676, 16'd65018, 16'd29762, 16'd34690, 16'd18958});
	test_expansion(128'h16bd47f04706946025161a3a7d0cbbe0, {16'd14206, 16'd41205, 16'd40976, 16'd60009, 16'd44555, 16'd3281, 16'd40360, 16'd10759, 16'd24762, 16'd64511, 16'd43561, 16'd63497, 16'd64242, 16'd56591, 16'd59019, 16'd27449, 16'd7534, 16'd808, 16'd14356, 16'd9681, 16'd4543, 16'd3469, 16'd37378, 16'd41756, 16'd29362, 16'd35247});
	test_expansion(128'h3e6549f0fab1785426f03e403b2f8528, {16'd51054, 16'd18451, 16'd38483, 16'd13913, 16'd4804, 16'd13820, 16'd24818, 16'd62173, 16'd28854, 16'd38844, 16'd33698, 16'd28815, 16'd4176, 16'd59229, 16'd48586, 16'd4342, 16'd59699, 16'd14251, 16'd40585, 16'd40110, 16'd25192, 16'd24107, 16'd47823, 16'd50071, 16'd708, 16'd9190});
	test_expansion(128'ha22c50c348991283ac1d96999e046732, {16'd14496, 16'd10258, 16'd4072, 16'd46615, 16'd47324, 16'd31963, 16'd56999, 16'd54765, 16'd19868, 16'd23599, 16'd32570, 16'd12, 16'd40211, 16'd38622, 16'd15012, 16'd58506, 16'd31278, 16'd48173, 16'd4413, 16'd38998, 16'd39519, 16'd29161, 16'd45868, 16'd10237, 16'd62789, 16'd39675});
	test_expansion(128'hbb1ee335dc2735b6f7dace4abebf7117, {16'd34605, 16'd9897, 16'd24309, 16'd51873, 16'd28168, 16'd40577, 16'd21908, 16'd39427, 16'd52694, 16'd44340, 16'd29944, 16'd42640, 16'd28272, 16'd18617, 16'd51644, 16'd56771, 16'd58158, 16'd49484, 16'd25639, 16'd47025, 16'd7327, 16'd12563, 16'd5421, 16'd15812, 16'd8116, 16'd8432});
	test_expansion(128'h369101a1122bc0d8a4466db3f3490d9b, {16'd51336, 16'd21411, 16'd39881, 16'd10017, 16'd57854, 16'd8450, 16'd59226, 16'd3937, 16'd58844, 16'd20696, 16'd27424, 16'd60227, 16'd10940, 16'd62593, 16'd42391, 16'd31300, 16'd34083, 16'd31260, 16'd29480, 16'd36350, 16'd10875, 16'd48304, 16'd16899, 16'd64633, 16'd9172, 16'd57961});
	test_expansion(128'hb4a9acf684a650d611e0a9a89eeffc90, {16'd47792, 16'd61188, 16'd27751, 16'd11291, 16'd40926, 16'd6797, 16'd55429, 16'd18438, 16'd62520, 16'd55707, 16'd52220, 16'd2220, 16'd29913, 16'd58041, 16'd36767, 16'd6067, 16'd56204, 16'd50704, 16'd41140, 16'd30860, 16'd59330, 16'd20326, 16'd64811, 16'd55500, 16'd14923, 16'd28265});
	test_expansion(128'h8b4d1413996f957778619601ef501031, {16'd23508, 16'd39195, 16'd32311, 16'd30043, 16'd48269, 16'd33830, 16'd18198, 16'd4507, 16'd60886, 16'd31589, 16'd12724, 16'd53042, 16'd6541, 16'd26697, 16'd47872, 16'd21685, 16'd40610, 16'd36602, 16'd1386, 16'd38381, 16'd20652, 16'd9120, 16'd16112, 16'd42855, 16'd36614, 16'd37019});
	test_expansion(128'ha460b0252b273c8d1e962e7a90fb9cf1, {16'd14654, 16'd27063, 16'd13249, 16'd64327, 16'd29340, 16'd49250, 16'd13845, 16'd45942, 16'd48772, 16'd3019, 16'd32707, 16'd65528, 16'd39572, 16'd57500, 16'd29102, 16'd33506, 16'd22067, 16'd8894, 16'd58365, 16'd6630, 16'd20070, 16'd160, 16'd55502, 16'd53287, 16'd63645, 16'd55277});
	test_expansion(128'ha99ec6ab285c329d8c6b7428ab1bdf25, {16'd57162, 16'd41628, 16'd42578, 16'd18053, 16'd61005, 16'd36430, 16'd47222, 16'd2782, 16'd62898, 16'd46965, 16'd13066, 16'd51154, 16'd24482, 16'd33993, 16'd23297, 16'd27876, 16'd18883, 16'd43257, 16'd13721, 16'd5664, 16'd6094, 16'd3278, 16'd14396, 16'd47632, 16'd14867, 16'd36485});
	test_expansion(128'hd0761fcc7fdf577c9081459c9fce85cd, {16'd35693, 16'd40855, 16'd14941, 16'd58733, 16'd50043, 16'd3193, 16'd51228, 16'd11280, 16'd27637, 16'd57957, 16'd10468, 16'd45818, 16'd25653, 16'd59116, 16'd63108, 16'd59269, 16'd53609, 16'd45997, 16'd49140, 16'd18950, 16'd64071, 16'd59103, 16'd58885, 16'd56207, 16'd57822, 16'd43975});
	test_expansion(128'h2ea5e357fbccf04fc89c9ac0a547d182, {16'd654, 16'd56362, 16'd31670, 16'd40020, 16'd41018, 16'd33629, 16'd43420, 16'd10465, 16'd39494, 16'd63268, 16'd43476, 16'd59371, 16'd13581, 16'd4658, 16'd5977, 16'd20919, 16'd32015, 16'd29181, 16'd60920, 16'd59513, 16'd30084, 16'd36508, 16'd5736, 16'd12699, 16'd13689, 16'd18633});
	test_expansion(128'hd8ba80b22153e8825cc8332a75e26bf6, {16'd49760, 16'd49229, 16'd11533, 16'd45373, 16'd32881, 16'd12599, 16'd54587, 16'd14956, 16'd12566, 16'd28336, 16'd44219, 16'd11297, 16'd55010, 16'd28316, 16'd13226, 16'd44625, 16'd38196, 16'd42889, 16'd9874, 16'd15024, 16'd27765, 16'd18373, 16'd62463, 16'd31883, 16'd12448, 16'd49340});
	test_expansion(128'hd37b554827a49e8959d17d89e1811629, {16'd55854, 16'd52827, 16'd50764, 16'd28073, 16'd6055, 16'd29255, 16'd6810, 16'd52752, 16'd18609, 16'd21161, 16'd26946, 16'd6682, 16'd62953, 16'd32378, 16'd64592, 16'd52646, 16'd63443, 16'd7578, 16'd29687, 16'd45936, 16'd33713, 16'd46551, 16'd18648, 16'd27712, 16'd3536, 16'd33695});
	test_expansion(128'hd71961a3bcd275c1bb146cf06a78be2b, {16'd53507, 16'd9503, 16'd41854, 16'd19146, 16'd3367, 16'd60752, 16'd264, 16'd64343, 16'd23557, 16'd40643, 16'd19872, 16'd19953, 16'd1876, 16'd10922, 16'd44687, 16'd1889, 16'd34671, 16'd11854, 16'd63867, 16'd47682, 16'd62152, 16'd56631, 16'd30026, 16'd16437, 16'd23864, 16'd23392});
	test_expansion(128'h3f422360dbcbc61b619bee99effd373e, {16'd56598, 16'd21590, 16'd8684, 16'd50715, 16'd41082, 16'd22672, 16'd5504, 16'd12497, 16'd14063, 16'd25035, 16'd10796, 16'd46116, 16'd41631, 16'd57540, 16'd60784, 16'd17693, 16'd47575, 16'd5730, 16'd57789, 16'd3389, 16'd29699, 16'd49994, 16'd7225, 16'd20279, 16'd50534, 16'd27373});
	test_expansion(128'h6a30215879b390d1926fab5511468ee4, {16'd43763, 16'd63387, 16'd13981, 16'd1650, 16'd14430, 16'd49670, 16'd24060, 16'd4859, 16'd29356, 16'd60118, 16'd1063, 16'd1918, 16'd8209, 16'd57762, 16'd27668, 16'd65150, 16'd43692, 16'd23402, 16'd42315, 16'd55022, 16'd62436, 16'd40179, 16'd57972, 16'd20547, 16'd48111, 16'd35217});
	test_expansion(128'h0f089b63375715d6f568fb0601a227ec, {16'd10035, 16'd14008, 16'd61874, 16'd26643, 16'd25416, 16'd61581, 16'd13497, 16'd1702, 16'd49278, 16'd14995, 16'd6917, 16'd40811, 16'd18537, 16'd7405, 16'd22743, 16'd35219, 16'd44406, 16'd59567, 16'd36184, 16'd63915, 16'd25140, 16'd54941, 16'd64012, 16'd15750, 16'd51062, 16'd46284});
	test_expansion(128'h617514e75cba7472db43e96b30ce0650, {16'd55595, 16'd17016, 16'd49606, 16'd30201, 16'd25795, 16'd24666, 16'd33505, 16'd32951, 16'd32637, 16'd10053, 16'd9031, 16'd5588, 16'd30321, 16'd28007, 16'd64482, 16'd55543, 16'd49555, 16'd50795, 16'd51175, 16'd7104, 16'd37707, 16'd11228, 16'd15919, 16'd45540, 16'd14461, 16'd44097});
	test_expansion(128'hbd560e84aa781b15d260b9a58322aef3, {16'd9339, 16'd12392, 16'd29530, 16'd8910, 16'd14443, 16'd51471, 16'd8613, 16'd21104, 16'd52323, 16'd30309, 16'd52917, 16'd60139, 16'd3379, 16'd42338, 16'd26098, 16'd47973, 16'd39761, 16'd65319, 16'd24771, 16'd10874, 16'd15187, 16'd38310, 16'd63226, 16'd47347, 16'd48154, 16'd53739});
	test_expansion(128'h24e509052b79d2a73c8865588ee636f0, {16'd52986, 16'd22480, 16'd14793, 16'd3718, 16'd59656, 16'd10254, 16'd21923, 16'd7136, 16'd27824, 16'd2903, 16'd60918, 16'd27892, 16'd44252, 16'd6726, 16'd7475, 16'd20795, 16'd53439, 16'd63173, 16'd36960, 16'd4108, 16'd64936, 16'd44262, 16'd35798, 16'd64503, 16'd40384, 16'd51368});
	test_expansion(128'h0ac2bc9d4ce193812c0ff3f59a67f727, {16'd23687, 16'd31807, 16'd1766, 16'd29695, 16'd50739, 16'd61233, 16'd9823, 16'd29335, 16'd42738, 16'd25669, 16'd13497, 16'd19966, 16'd15932, 16'd56958, 16'd40181, 16'd9569, 16'd38912, 16'd31038, 16'd44475, 16'd32723, 16'd58117, 16'd38269, 16'd57851, 16'd26623, 16'd30345, 16'd26281});
	test_expansion(128'h32a1ac379959566e13862318d5fc35c2, {16'd5103, 16'd49451, 16'd33975, 16'd62231, 16'd55212, 16'd2945, 16'd24099, 16'd29366, 16'd11863, 16'd11973, 16'd40086, 16'd23060, 16'd34557, 16'd64165, 16'd31884, 16'd24492, 16'd4753, 16'd3911, 16'd36442, 16'd18029, 16'd6686, 16'd59552, 16'd1355, 16'd58190, 16'd13284, 16'd60252});
	test_expansion(128'ha9426d8ad06889703a8c01667bc97626, {16'd6528, 16'd10052, 16'd31801, 16'd41715, 16'd33388, 16'd27, 16'd3928, 16'd15545, 16'd38052, 16'd24916, 16'd34756, 16'd26205, 16'd24132, 16'd22441, 16'd28448, 16'd65333, 16'd62451, 16'd23660, 16'd54755, 16'd54267, 16'd24547, 16'd65429, 16'd40022, 16'd18351, 16'd30378, 16'd53344});
	test_expansion(128'h6d1aa36352872a7f62296b16ddfa5c2b, {16'd32772, 16'd4191, 16'd50889, 16'd8844, 16'd13931, 16'd62984, 16'd16666, 16'd34830, 16'd27808, 16'd53946, 16'd29847, 16'd58319, 16'd33403, 16'd58975, 16'd61453, 16'd43790, 16'd61322, 16'd22171, 16'd2467, 16'd24586, 16'd52793, 16'd44926, 16'd29410, 16'd829, 16'd20051, 16'd17440});
	test_expansion(128'hcb94ea622d9493f4b4dadc642cfcbf71, {16'd24271, 16'd39937, 16'd61280, 16'd57870, 16'd27606, 16'd35912, 16'd52979, 16'd30566, 16'd34314, 16'd2702, 16'd3795, 16'd57491, 16'd59196, 16'd31083, 16'd59231, 16'd7097, 16'd36586, 16'd39434, 16'd8759, 16'd30034, 16'd60626, 16'd51956, 16'd27114, 16'd48874, 16'd161, 16'd56376});
	test_expansion(128'h4d20a3bd41b1b330e2cf830a31fd29c1, {16'd56608, 16'd37753, 16'd16327, 16'd45004, 16'd59390, 16'd9666, 16'd36242, 16'd64252, 16'd20367, 16'd45077, 16'd7016, 16'd34870, 16'd55690, 16'd60249, 16'd44031, 16'd613, 16'd7969, 16'd9785, 16'd31544, 16'd62172, 16'd8957, 16'd34613, 16'd51184, 16'd24779, 16'd19707, 16'd21564});
	test_expansion(128'h9c5a73a65fd8252d4543644faa009785, {16'd15634, 16'd42750, 16'd2278, 16'd59409, 16'd5678, 16'd40041, 16'd47028, 16'd42437, 16'd10423, 16'd43132, 16'd62573, 16'd31796, 16'd54358, 16'd13477, 16'd55996, 16'd26693, 16'd19685, 16'd29542, 16'd28345, 16'd46152, 16'd29167, 16'd37843, 16'd3119, 16'd18930, 16'd9487, 16'd44921});
	test_expansion(128'h861542b87f56d7f1a1fb8863656502dd, {16'd62039, 16'd60713, 16'd28541, 16'd18406, 16'd2494, 16'd15123, 16'd57831, 16'd42624, 16'd64456, 16'd41607, 16'd61735, 16'd44776, 16'd50844, 16'd51364, 16'd63022, 16'd33728, 16'd4449, 16'd65115, 16'd31412, 16'd18545, 16'd26276, 16'd56723, 16'd24544, 16'd41146, 16'd1826, 16'd2778});
	test_expansion(128'h5e8ad30cd54923951938240da3ffd4c6, {16'd46609, 16'd22698, 16'd43446, 16'd41447, 16'd39949, 16'd37693, 16'd27264, 16'd23911, 16'd4691, 16'd26079, 16'd39196, 16'd95, 16'd30856, 16'd23146, 16'd38600, 16'd33968, 16'd13510, 16'd42508, 16'd52169, 16'd8313, 16'd26335, 16'd52879, 16'd1085, 16'd40988, 16'd60942, 16'd63317});
	test_expansion(128'h827a789e9d0708acf0959d012f2ed0d5, {16'd13499, 16'd32753, 16'd55766, 16'd29268, 16'd1235, 16'd1600, 16'd29016, 16'd29390, 16'd17045, 16'd44597, 16'd44410, 16'd56289, 16'd53415, 16'd20373, 16'd21607, 16'd1734, 16'd47395, 16'd41515, 16'd63563, 16'd7164, 16'd18409, 16'd31826, 16'd64775, 16'd3417, 16'd65275, 16'd26883});
	test_expansion(128'h06e5cdb7bb17c5ac109730b65e90dee7, {16'd2430, 16'd55992, 16'd7056, 16'd64681, 16'd45764, 16'd45024, 16'd34666, 16'd32877, 16'd53046, 16'd27961, 16'd17180, 16'd12980, 16'd56837, 16'd38502, 16'd52080, 16'd20027, 16'd3671, 16'd41638, 16'd43847, 16'd39194, 16'd30570, 16'd58937, 16'd64835, 16'd3198, 16'd21451, 16'd43478});
	test_expansion(128'h0b6662dfc592e8c8e779c4414ecd3ebe, {16'd31964, 16'd27579, 16'd52397, 16'd6373, 16'd19542, 16'd31019, 16'd9853, 16'd41801, 16'd58065, 16'd41283, 16'd45556, 16'd55489, 16'd41261, 16'd37145, 16'd5250, 16'd18813, 16'd44340, 16'd46972, 16'd47917, 16'd32722, 16'd55720, 16'd17915, 16'd35079, 16'd58639, 16'd45718, 16'd29187});
	test_expansion(128'hd2303a9ffb86c20ac58e3a29c0ee1c85, {16'd31217, 16'd45488, 16'd5227, 16'd45341, 16'd46877, 16'd15303, 16'd38232, 16'd31792, 16'd50825, 16'd13199, 16'd15996, 16'd56810, 16'd49396, 16'd13735, 16'd35334, 16'd11436, 16'd20920, 16'd22598, 16'd891, 16'd31466, 16'd2158, 16'd46848, 16'd4204, 16'd6053, 16'd32950, 16'd36151});
	test_expansion(128'h13524c0c64b7fae22d970a3f49056bd4, {16'd16804, 16'd47788, 16'd11341, 16'd24023, 16'd40026, 16'd62448, 16'd31766, 16'd45366, 16'd9366, 16'd37835, 16'd2572, 16'd26340, 16'd48986, 16'd11302, 16'd41260, 16'd11125, 16'd62019, 16'd53722, 16'd1943, 16'd50240, 16'd52283, 16'd46926, 16'd520, 16'd22395, 16'd34754, 16'd27811});
	test_expansion(128'h2cd737125f2e2d94611c81a46a9338f4, {16'd36838, 16'd25924, 16'd29111, 16'd60465, 16'd16979, 16'd42820, 16'd2149, 16'd19879, 16'd60873, 16'd18235, 16'd23218, 16'd65392, 16'd43766, 16'd24767, 16'd13972, 16'd16760, 16'd50652, 16'd35714, 16'd58970, 16'd63049, 16'd6845, 16'd16171, 16'd24528, 16'd17664, 16'd17640, 16'd28193});
	test_expansion(128'h18ac6a42e911df625d0a8fc20fe93295, {16'd7943, 16'd52872, 16'd50133, 16'd15472, 16'd53584, 16'd37783, 16'd21475, 16'd27514, 16'd23074, 16'd42986, 16'd55890, 16'd43577, 16'd16577, 16'd15132, 16'd2596, 16'd61634, 16'd2305, 16'd57978, 16'd59661, 16'd52595, 16'd58517, 16'd41815, 16'd27064, 16'd48327, 16'd6688, 16'd61888});
	test_expansion(128'h0890d1b6f649786f2fadc57f2a2c48a2, {16'd9228, 16'd64952, 16'd15812, 16'd933, 16'd56305, 16'd31779, 16'd33166, 16'd15875, 16'd30847, 16'd33461, 16'd40376, 16'd23769, 16'd2463, 16'd46800, 16'd24260, 16'd5003, 16'd54106, 16'd50011, 16'd58585, 16'd26268, 16'd27550, 16'd61462, 16'd54533, 16'd56642, 16'd60420, 16'd37760});
	test_expansion(128'hfbee42a1d166dc33cd25b2a01a67abf4, {16'd37827, 16'd49204, 16'd42260, 16'd42396, 16'd63927, 16'd31636, 16'd62726, 16'd58663, 16'd44874, 16'd62464, 16'd28090, 16'd27362, 16'd12851, 16'd4973, 16'd30544, 16'd36664, 16'd38709, 16'd5414, 16'd3821, 16'd484, 16'd45469, 16'd64581, 16'd57194, 16'd10573, 16'd53682, 16'd6389});
	test_expansion(128'h9b7821b52d8ea269ed13e6d2e6d4a6a0, {16'd46179, 16'd60481, 16'd1283, 16'd49817, 16'd26672, 16'd17311, 16'd19381, 16'd13373, 16'd22746, 16'd56819, 16'd20151, 16'd13033, 16'd19213, 16'd61596, 16'd46020, 16'd6804, 16'd28726, 16'd22411, 16'd24468, 16'd59647, 16'd45700, 16'd62984, 16'd52739, 16'd28194, 16'd6667, 16'd45086});
	test_expansion(128'h53c938159eda560f93f920bda8356210, {16'd63720, 16'd6029, 16'd44047, 16'd65428, 16'd35072, 16'd32997, 16'd7576, 16'd684, 16'd53778, 16'd4139, 16'd36763, 16'd44768, 16'd60257, 16'd42547, 16'd23396, 16'd37791, 16'd2679, 16'd9111, 16'd16498, 16'd49953, 16'd33795, 16'd57959, 16'd31786, 16'd33538, 16'd32785, 16'd48875});
	test_expansion(128'hff27fa89876643e19f7c068ad6f5a408, {16'd21034, 16'd24251, 16'd61287, 16'd24656, 16'd8657, 16'd10198, 16'd8807, 16'd28653, 16'd16956, 16'd42501, 16'd29108, 16'd33844, 16'd32316, 16'd35155, 16'd34191, 16'd5645, 16'd63178, 16'd24061, 16'd11848, 16'd30556, 16'd36548, 16'd60207, 16'd20592, 16'd7341, 16'd34228, 16'd58246});
	test_expansion(128'h4fe6625ad3d62ecc76b5d6a0cb56eeaf, {16'd7163, 16'd29557, 16'd35899, 16'd56639, 16'd34850, 16'd26088, 16'd44913, 16'd30647, 16'd56028, 16'd9893, 16'd6876, 16'd30742, 16'd42101, 16'd40975, 16'd64933, 16'd39334, 16'd52264, 16'd12985, 16'd8047, 16'd49450, 16'd19607, 16'd32427, 16'd4900, 16'd42074, 16'd29725, 16'd48511});
	test_expansion(128'h4b723738e5e7b3a7488ccb6ba6dce4ec, {16'd11672, 16'd26682, 16'd29982, 16'd36741, 16'd42118, 16'd7991, 16'd54462, 16'd31876, 16'd27328, 16'd51665, 16'd38032, 16'd58510, 16'd17278, 16'd19157, 16'd46438, 16'd52880, 16'd1774, 16'd48721, 16'd18632, 16'd48762, 16'd24089, 16'd27846, 16'd36680, 16'd20919, 16'd61933, 16'd49654});
	test_expansion(128'h9882d0328e6546b0054a490a75cb4b17, {16'd19068, 16'd10431, 16'd44212, 16'd3460, 16'd21201, 16'd36001, 16'd11036, 16'd34118, 16'd49319, 16'd9421, 16'd57871, 16'd53301, 16'd30113, 16'd25234, 16'd59294, 16'd45394, 16'd14151, 16'd60341, 16'd9216, 16'd15114, 16'd38242, 16'd31803, 16'd18092, 16'd27236, 16'd12897, 16'd13528});
	test_expansion(128'h7c4bb2bad0245a6fc25596961ab87aa0, {16'd25793, 16'd59416, 16'd21721, 16'd17161, 16'd42996, 16'd64509, 16'd63956, 16'd19343, 16'd16911, 16'd42364, 16'd37737, 16'd25092, 16'd38407, 16'd9604, 16'd10854, 16'd15936, 16'd15337, 16'd25730, 16'd57825, 16'd17794, 16'd5817, 16'd34340, 16'd11442, 16'd57001, 16'd17944, 16'd6201});
	test_expansion(128'h3dd9d38bcf3f289c84796c164c9b8629, {16'd46290, 16'd3028, 16'd38158, 16'd55594, 16'd13561, 16'd19507, 16'd62253, 16'd53333, 16'd54834, 16'd15662, 16'd11157, 16'd38748, 16'd62109, 16'd22534, 16'd28223, 16'd30755, 16'd23556, 16'd4545, 16'd58396, 16'd32264, 16'd47356, 16'd45833, 16'd23276, 16'd40880, 16'd53725, 16'd4839});
	test_expansion(128'h94489147e751c3c5a7dac7dbf91a696c, {16'd59550, 16'd2352, 16'd2798, 16'd10000, 16'd7843, 16'd37475, 16'd52521, 16'd19907, 16'd6215, 16'd5817, 16'd25404, 16'd52614, 16'd60393, 16'd222, 16'd55106, 16'd45741, 16'd25377, 16'd31557, 16'd15918, 16'd23752, 16'd57342, 16'd46199, 16'd11811, 16'd37828, 16'd29425, 16'd30925});
	test_expansion(128'ha2aa69e0f184f8980a20f92a9467fe94, {16'd31467, 16'd56475, 16'd33263, 16'd62824, 16'd60186, 16'd37053, 16'd64716, 16'd15982, 16'd6722, 16'd64115, 16'd26780, 16'd52377, 16'd2504, 16'd60262, 16'd338, 16'd27828, 16'd51550, 16'd20357, 16'd32555, 16'd26427, 16'd46968, 16'd7587, 16'd55736, 16'd28045, 16'd39088, 16'd54963});
	test_expansion(128'h6791b9f3f45bda572e345059c7f5fb23, {16'd62896, 16'd9009, 16'd61313, 16'd60143, 16'd37431, 16'd36652, 16'd7290, 16'd56665, 16'd40718, 16'd23923, 16'd39319, 16'd60985, 16'd30464, 16'd53375, 16'd51352, 16'd30213, 16'd28009, 16'd44284, 16'd42959, 16'd14727, 16'd24264, 16'd26402, 16'd52093, 16'd11244, 16'd62980, 16'd43674});
	test_expansion(128'hdd1d3ccba7b62634d6544194cbce79f6, {16'd34475, 16'd40330, 16'd31861, 16'd35836, 16'd35536, 16'd61526, 16'd24948, 16'd45785, 16'd45672, 16'd15914, 16'd46614, 16'd53254, 16'd8970, 16'd9635, 16'd2430, 16'd34639, 16'd51062, 16'd19806, 16'd51657, 16'd3577, 16'd51019, 16'd4550, 16'd29810, 16'd3682, 16'd35706, 16'd40929});
	test_expansion(128'hd1707c2844903d6d39d9acf3949a12e2, {16'd53682, 16'd65176, 16'd25001, 16'd11467, 16'd58148, 16'd9417, 16'd8888, 16'd40347, 16'd28554, 16'd4631, 16'd10287, 16'd61226, 16'd62454, 16'd18536, 16'd64318, 16'd16363, 16'd51788, 16'd50416, 16'd14006, 16'd58520, 16'd36809, 16'd15551, 16'd28388, 16'd20612, 16'd2791, 16'd58888});
	test_expansion(128'h0c752ae1fc68ffa264624cde7aa36115, {16'd25400, 16'd3011, 16'd50148, 16'd29293, 16'd47546, 16'd29881, 16'd40427, 16'd11816, 16'd23486, 16'd46829, 16'd64312, 16'd13802, 16'd63088, 16'd11343, 16'd4662, 16'd32887, 16'd15845, 16'd8184, 16'd62343, 16'd43925, 16'd25889, 16'd59421, 16'd8251, 16'd29350, 16'd54907, 16'd53424});
	test_expansion(128'hc044179e5192336c133d4a1fe9f1281f, {16'd525, 16'd58401, 16'd59710, 16'd47263, 16'd46353, 16'd46003, 16'd28374, 16'd192, 16'd3563, 16'd20618, 16'd21404, 16'd29232, 16'd1220, 16'd30054, 16'd41286, 16'd40858, 16'd19487, 16'd30499, 16'd52406, 16'd61073, 16'd30946, 16'd38905, 16'd53916, 16'd43842, 16'd7582, 16'd52976});
	test_expansion(128'h189afada225cd4ad559edf39b58649b8, {16'd28722, 16'd58564, 16'd45274, 16'd30927, 16'd47615, 16'd20084, 16'd29855, 16'd55813, 16'd11583, 16'd29329, 16'd8491, 16'd22423, 16'd63030, 16'd45552, 16'd7052, 16'd6112, 16'd19963, 16'd41264, 16'd22663, 16'd53830, 16'd29950, 16'd44799, 16'd18512, 16'd41679, 16'd33770, 16'd9006});
	test_expansion(128'he3c4134bd419d857ab926cd9f809254e, {16'd59559, 16'd7431, 16'd41974, 16'd59701, 16'd51108, 16'd59277, 16'd22162, 16'd40446, 16'd16020, 16'd50199, 16'd14324, 16'd14516, 16'd2373, 16'd63404, 16'd20540, 16'd6466, 16'd27318, 16'd47553, 16'd49012, 16'd48618, 16'd10012, 16'd30538, 16'd14151, 16'd12317, 16'd63484, 16'd50758});
	test_expansion(128'hf100de0e56b1a49ce6468d319799b27c, {16'd33160, 16'd7854, 16'd17780, 16'd8317, 16'd26383, 16'd27783, 16'd41779, 16'd15998, 16'd54929, 16'd62482, 16'd44868, 16'd61151, 16'd22928, 16'd50589, 16'd35841, 16'd65375, 16'd64152, 16'd63729, 16'd53211, 16'd41445, 16'd59368, 16'd2580, 16'd36490, 16'd13523, 16'd39199, 16'd9769});
	test_expansion(128'hc9102b6e34b04ec7280855291ea372e4, {16'd31226, 16'd39339, 16'd30867, 16'd22549, 16'd50997, 16'd53802, 16'd18054, 16'd38821, 16'd62728, 16'd24702, 16'd37589, 16'd8704, 16'd55645, 16'd34824, 16'd37331, 16'd42981, 16'd8289, 16'd49049, 16'd3646, 16'd35869, 16'd46952, 16'd40799, 16'd2826, 16'd27618, 16'd30417, 16'd21685});
	test_expansion(128'h7b2794a744da5eeb1b5d252b641b12d8, {16'd29465, 16'd59217, 16'd16774, 16'd23268, 16'd5481, 16'd13303, 16'd18033, 16'd9967, 16'd59423, 16'd64605, 16'd27816, 16'd32987, 16'd44898, 16'd31089, 16'd1189, 16'd28762, 16'd22135, 16'd22433, 16'd58759, 16'd925, 16'd64013, 16'd36746, 16'd16638, 16'd60592, 16'd19995, 16'd7375});
	test_expansion(128'h50886c3587d2d6ae76a274affbf6d31d, {16'd9143, 16'd31270, 16'd24537, 16'd9589, 16'd44771, 16'd48527, 16'd61547, 16'd50449, 16'd62692, 16'd53555, 16'd18375, 16'd35586, 16'd56891, 16'd43239, 16'd62306, 16'd12251, 16'd48837, 16'd24122, 16'd62160, 16'd37490, 16'd40105, 16'd44184, 16'd7276, 16'd16947, 16'd2151, 16'd59817});
	test_expansion(128'h2239da6664ff71f60289272334843fb8, {16'd31842, 16'd11154, 16'd36815, 16'd34412, 16'd25095, 16'd16708, 16'd23048, 16'd133, 16'd26027, 16'd4294, 16'd64999, 16'd62951, 16'd8014, 16'd8445, 16'd40324, 16'd14671, 16'd6161, 16'd47689, 16'd1184, 16'd60033, 16'd63061, 16'd14410, 16'd21921, 16'd54074, 16'd45486, 16'd4514});
	test_expansion(128'h185912e21d7f0690da1cd988c49fde94, {16'd8760, 16'd16990, 16'd5663, 16'd61337, 16'd16847, 16'd27685, 16'd7385, 16'd59965, 16'd47919, 16'd42840, 16'd40177, 16'd32410, 16'd29212, 16'd11717, 16'd45183, 16'd23731, 16'd2085, 16'd64883, 16'd1098, 16'd32457, 16'd47491, 16'd32840, 16'd57593, 16'd52963, 16'd62599, 16'd18069});
	test_expansion(128'h0333b1390c9ffa69a07a9afd5eb63ed3, {16'd49514, 16'd8918, 16'd6963, 16'd5230, 16'd43654, 16'd17707, 16'd16861, 16'd42770, 16'd28335, 16'd45840, 16'd62814, 16'd20137, 16'd52876, 16'd50722, 16'd31311, 16'd22423, 16'd28287, 16'd19460, 16'd35240, 16'd38713, 16'd35716, 16'd4199, 16'd22118, 16'd39291, 16'd5923, 16'd9602});
	test_expansion(128'h22c652b0e72be584f7bb521e1ea0fdca, {16'd52845, 16'd35722, 16'd63872, 16'd30408, 16'd58906, 16'd20343, 16'd20186, 16'd52745, 16'd34061, 16'd26540, 16'd8287, 16'd10442, 16'd56723, 16'd36230, 16'd33590, 16'd52074, 16'd33077, 16'd57290, 16'd64012, 16'd19841, 16'd43044, 16'd38745, 16'd27636, 16'd12199, 16'd2887, 16'd15824});
	test_expansion(128'h36b959a81ec1ca7368b4131cf2e3a214, {16'd20667, 16'd37483, 16'd43475, 16'd2777, 16'd61402, 16'd19911, 16'd50851, 16'd58662, 16'd34366, 16'd25738, 16'd57429, 16'd7381, 16'd46063, 16'd49841, 16'd42985, 16'd48916, 16'd6662, 16'd30073, 16'd16306, 16'd54615, 16'd4326, 16'd60107, 16'd26030, 16'd26973, 16'd43980, 16'd38803});
	test_expansion(128'h5fbf62f4c19a3d6097fe27e615d88791, {16'd48674, 16'd19060, 16'd42334, 16'd36892, 16'd52943, 16'd20915, 16'd21999, 16'd33640, 16'd12680, 16'd955, 16'd37584, 16'd25533, 16'd65028, 16'd42897, 16'd53037, 16'd3320, 16'd57955, 16'd33377, 16'd33714, 16'd49427, 16'd41181, 16'd7790, 16'd11735, 16'd51058, 16'd35618, 16'd8268});
	test_expansion(128'h9f3b7e02f028498bbdbdd34b121fa81c, {16'd30019, 16'd31913, 16'd60351, 16'd11200, 16'd24154, 16'd54561, 16'd7653, 16'd64038, 16'd44054, 16'd46810, 16'd1994, 16'd23892, 16'd57514, 16'd38214, 16'd48903, 16'd54364, 16'd31299, 16'd45482, 16'd15260, 16'd62255, 16'd4822, 16'd53461, 16'd3608, 16'd2959, 16'd20391, 16'd62863});
	test_expansion(128'hf7637147c926bb7653d0c6180cf49ff1, {16'd1544, 16'd10896, 16'd41124, 16'd60848, 16'd60123, 16'd488, 16'd8331, 16'd34144, 16'd27426, 16'd23645, 16'd41534, 16'd9462, 16'd63386, 16'd16242, 16'd55989, 16'd59051, 16'd14358, 16'd23871, 16'd20173, 16'd2896, 16'd60632, 16'd50801, 16'd60174, 16'd46919, 16'd18371, 16'd24990});
	test_expansion(128'h2296e1452fe9fa7674dc5449c95c2ddc, {16'd20097, 16'd13403, 16'd38002, 16'd23020, 16'd61149, 16'd26866, 16'd47686, 16'd53596, 16'd39696, 16'd60361, 16'd63400, 16'd23948, 16'd56188, 16'd30759, 16'd61569, 16'd38051, 16'd19270, 16'd7862, 16'd60293, 16'd58942, 16'd42590, 16'd29064, 16'd29624, 16'd49346, 16'd2146, 16'd51269});
	test_expansion(128'he67b672bc27dd470fd6e511f44f86d37, {16'd38947, 16'd2773, 16'd33570, 16'd49821, 16'd44591, 16'd37345, 16'd39598, 16'd30897, 16'd19547, 16'd26737, 16'd50578, 16'd32352, 16'd31207, 16'd4355, 16'd3363, 16'd29417, 16'd3244, 16'd29422, 16'd44859, 16'd39329, 16'd32593, 16'd61959, 16'd7101, 16'd22486, 16'd40257, 16'd9125});
	test_expansion(128'h1eff4e03d6ba00a9e05f775706ac8921, {16'd54797, 16'd55304, 16'd63275, 16'd57406, 16'd22004, 16'd14575, 16'd40043, 16'd42821, 16'd38277, 16'd61214, 16'd26886, 16'd29887, 16'd60522, 16'd55647, 16'd23473, 16'd18849, 16'd25825, 16'd7259, 16'd1197, 16'd11097, 16'd65135, 16'd60234, 16'd36624, 16'd46881, 16'd65147, 16'd28820});
	test_expansion(128'h46e295b96869f181c0e5aa76a839eb0c, {16'd25505, 16'd40959, 16'd50194, 16'd55103, 16'd37313, 16'd29943, 16'd41874, 16'd39722, 16'd7376, 16'd53169, 16'd23450, 16'd56774, 16'd56153, 16'd16041, 16'd50303, 16'd36708, 16'd22352, 16'd22247, 16'd38425, 16'd56066, 16'd5043, 16'd41745, 16'd53799, 16'd64301, 16'd45884, 16'd38787});
	test_expansion(128'h4ff7dee9a4bccf728f9afd8b1ad9ff6b, {16'd705, 16'd61674, 16'd20980, 16'd50220, 16'd30463, 16'd50590, 16'd57759, 16'd19161, 16'd29895, 16'd6994, 16'd25745, 16'd53553, 16'd55070, 16'd2521, 16'd50848, 16'd14945, 16'd52428, 16'd17092, 16'd52662, 16'd48437, 16'd19352, 16'd60431, 16'd17578, 16'd14767, 16'd43110, 16'd7612});
	test_expansion(128'he132acb5e6562d71aca44500f0e57924, {16'd19428, 16'd41254, 16'd32232, 16'd28208, 16'd2993, 16'd58583, 16'd63920, 16'd13170, 16'd50196, 16'd57485, 16'd61341, 16'd10952, 16'd30109, 16'd61998, 16'd58369, 16'd26015, 16'd23883, 16'd27503, 16'd63275, 16'd22494, 16'd57987, 16'd63893, 16'd28154, 16'd39295, 16'd9738, 16'd33223});
	test_expansion(128'h836ce6b78d3d17b729b0eab4271c3a35, {16'd23588, 16'd57343, 16'd25689, 16'd52930, 16'd20322, 16'd60726, 16'd25216, 16'd37306, 16'd56512, 16'd26910, 16'd17959, 16'd14115, 16'd39981, 16'd42883, 16'd32871, 16'd53521, 16'd60474, 16'd64598, 16'd27715, 16'd42340, 16'd8421, 16'd22515, 16'd15826, 16'd62533, 16'd47598, 16'd2589});
	test_expansion(128'ha915598fc6d12d7eaac03bce8084684c, {16'd541, 16'd17632, 16'd50918, 16'd17133, 16'd713, 16'd23125, 16'd48258, 16'd26645, 16'd49214, 16'd12850, 16'd59730, 16'd3081, 16'd49742, 16'd62149, 16'd15393, 16'd19784, 16'd58160, 16'd38260, 16'd44303, 16'd59378, 16'd2727, 16'd5446, 16'd52173, 16'd25055, 16'd13529, 16'd30095});
	test_expansion(128'h0ad49f5831c6adbaaf4db47ae8147deb, {16'd26961, 16'd40270, 16'd62640, 16'd19792, 16'd48556, 16'd5052, 16'd29745, 16'd61993, 16'd11701, 16'd39803, 16'd23064, 16'd55884, 16'd60297, 16'd65430, 16'd47599, 16'd30002, 16'd34910, 16'd25586, 16'd44470, 16'd28256, 16'd19345, 16'd548, 16'd44075, 16'd61323, 16'd65013, 16'd39795});
	test_expansion(128'h2f174d9ace5b3cff4b8a359658f86c25, {16'd24548, 16'd42352, 16'd21948, 16'd17408, 16'd2385, 16'd14574, 16'd37672, 16'd55816, 16'd17654, 16'd36413, 16'd7177, 16'd16345, 16'd57503, 16'd6250, 16'd57597, 16'd9109, 16'd45776, 16'd19907, 16'd36789, 16'd64586, 16'd64864, 16'd64111, 16'd10070, 16'd16425, 16'd41280, 16'd34880});
	test_expansion(128'h91328ca73f2cf6944bb081cb714460eb, {16'd5502, 16'd28229, 16'd7800, 16'd49823, 16'd25523, 16'd15621, 16'd30004, 16'd10506, 16'd5703, 16'd40532, 16'd43529, 16'd3345, 16'd22105, 16'd7676, 16'd54295, 16'd27238, 16'd13871, 16'd58651, 16'd6719, 16'd35365, 16'd13734, 16'd6211, 16'd41926, 16'd61676, 16'd48843, 16'd26195});
	test_expansion(128'hf79c48689bc9688b3fd8fdf3aa4e6aed, {16'd2028, 16'd32278, 16'd64434, 16'd44503, 16'd4758, 16'd19239, 16'd43883, 16'd3458, 16'd64023, 16'd65323, 16'd1495, 16'd52718, 16'd43162, 16'd40964, 16'd32856, 16'd61160, 16'd50683, 16'd33113, 16'd15924, 16'd47451, 16'd41085, 16'd60048, 16'd27784, 16'd18959, 16'd30119, 16'd13223});
	test_expansion(128'h08e7d4a69680a68e52b30d27ee5b2b37, {16'd4227, 16'd36146, 16'd18270, 16'd34565, 16'd31938, 16'd19025, 16'd60624, 16'd1967, 16'd32952, 16'd5333, 16'd62389, 16'd44947, 16'd37408, 16'd64326, 16'd8697, 16'd50517, 16'd36021, 16'd22087, 16'd55148, 16'd7064, 16'd13273, 16'd49273, 16'd35056, 16'd26232, 16'd24007, 16'd20464});
	test_expansion(128'h298cfcd2b508aac899bd2c50d74d56f7, {16'd38484, 16'd47651, 16'd18314, 16'd8303, 16'd3620, 16'd41935, 16'd11415, 16'd10822, 16'd54583, 16'd16267, 16'd10129, 16'd29663, 16'd57722, 16'd58594, 16'd24, 16'd23873, 16'd53975, 16'd35921, 16'd38874, 16'd32060, 16'd40485, 16'd46872, 16'd41105, 16'd35004, 16'd25636, 16'd45377});
	test_expansion(128'hda39371b226156a27ad9cb1c5618cc71, {16'd19329, 16'd48353, 16'd36778, 16'd18395, 16'd29163, 16'd13250, 16'd14836, 16'd39707, 16'd25802, 16'd41684, 16'd11870, 16'd31500, 16'd3088, 16'd2491, 16'd38723, 16'd19392, 16'd23717, 16'd12507, 16'd36150, 16'd25426, 16'd59356, 16'd51340, 16'd8951, 16'd48608, 16'd25148, 16'd62505});
	test_expansion(128'h543975810ead16c94475ae083861642f, {16'd52303, 16'd30080, 16'd32487, 16'd21118, 16'd46328, 16'd32867, 16'd11071, 16'd12430, 16'd28465, 16'd32702, 16'd36381, 16'd41801, 16'd44591, 16'd53333, 16'd30239, 16'd59765, 16'd43074, 16'd18623, 16'd17744, 16'd23826, 16'd46506, 16'd51859, 16'd54325, 16'd23021, 16'd25976, 16'd13130});
	test_expansion(128'hdeb661697014d1d8adb3b4e42fa4973f, {16'd28797, 16'd59712, 16'd11599, 16'd34504, 16'd19458, 16'd15184, 16'd61138, 16'd64909, 16'd62933, 16'd24810, 16'd55738, 16'd8391, 16'd49761, 16'd59271, 16'd43866, 16'd32547, 16'd28577, 16'd18828, 16'd38468, 16'd22778, 16'd58422, 16'd15953, 16'd33120, 16'd42376, 16'd5954, 16'd51277});
	test_expansion(128'h9d17c084c5ad7439be7818fb3d18bb46, {16'd12356, 16'd38633, 16'd41080, 16'd45156, 16'd33567, 16'd20586, 16'd1293, 16'd15865, 16'd19423, 16'd35453, 16'd33674, 16'd15476, 16'd58092, 16'd44834, 16'd49906, 16'd13578, 16'd26991, 16'd53659, 16'd60671, 16'd16580, 16'd41554, 16'd24428, 16'd43449, 16'd16604, 16'd62429, 16'd26930});
	test_expansion(128'h527c3b43e5b9ab07e4115634fe94dfea, {16'd38459, 16'd45547, 16'd35855, 16'd11512, 16'd22066, 16'd10942, 16'd34590, 16'd40914, 16'd63265, 16'd15044, 16'd50643, 16'd20686, 16'd25650, 16'd54336, 16'd46861, 16'd7243, 16'd51023, 16'd4070, 16'd53209, 16'd14935, 16'd46363, 16'd34461, 16'd49165, 16'd5524, 16'd63812, 16'd28280});
	test_expansion(128'h585c85ba579be0c7ec3b028dae2f2574, {16'd29992, 16'd55127, 16'd54807, 16'd28049, 16'd28397, 16'd39939, 16'd55964, 16'd53447, 16'd57098, 16'd36557, 16'd29613, 16'd32069, 16'd23409, 16'd10390, 16'd38986, 16'd31967, 16'd43105, 16'd38477, 16'd40685, 16'd37705, 16'd25618, 16'd22202, 16'd44019, 16'd41564, 16'd28358, 16'd41285});
	test_expansion(128'hd65a64e86ea5510bf35d82a08b8ddf1f, {16'd2353, 16'd40750, 16'd14965, 16'd61712, 16'd24697, 16'd32533, 16'd17981, 16'd32835, 16'd62964, 16'd39848, 16'd790, 16'd48061, 16'd3868, 16'd35030, 16'd22500, 16'd50481, 16'd26909, 16'd58977, 16'd51617, 16'd55641, 16'd10810, 16'd10048, 16'd24506, 16'd42174, 16'd40539, 16'd14513});
	test_expansion(128'haf91eec28e9a651f44cdd625904e1ca3, {16'd41639, 16'd54737, 16'd16912, 16'd26033, 16'd42220, 16'd29977, 16'd20207, 16'd11064, 16'd46129, 16'd28246, 16'd56781, 16'd2722, 16'd58650, 16'd57237, 16'd55022, 16'd21205, 16'd40522, 16'd44983, 16'd63339, 16'd793, 16'd43367, 16'd35157, 16'd55729, 16'd24782, 16'd24238, 16'd40700});
	test_expansion(128'h364801d574b2476bfafb2176e73e72a8, {16'd23934, 16'd24169, 16'd13035, 16'd4025, 16'd26418, 16'd56668, 16'd7385, 16'd11569, 16'd45089, 16'd15022, 16'd5386, 16'd4458, 16'd55723, 16'd7607, 16'd50718, 16'd2792, 16'd38436, 16'd51941, 16'd24995, 16'd60700, 16'd50820, 16'd51726, 16'd41721, 16'd36329, 16'd4932, 16'd62424});
	test_expansion(128'h578aa35773c4374f62c32b60c811cc76, {16'd30115, 16'd15443, 16'd39535, 16'd55134, 16'd35438, 16'd33643, 16'd13420, 16'd9417, 16'd46300, 16'd26477, 16'd42283, 16'd32712, 16'd63862, 16'd22688, 16'd56957, 16'd30273, 16'd36643, 16'd63576, 16'd10520, 16'd27907, 16'd64015, 16'd38975, 16'd53821, 16'd42208, 16'd43666, 16'd6919});
	test_expansion(128'h34bdf10fb743d044b0e0f7ba10961da7, {16'd28155, 16'd21179, 16'd17868, 16'd7652, 16'd37062, 16'd26862, 16'd13751, 16'd27940, 16'd20678, 16'd35964, 16'd5994, 16'd40361, 16'd44070, 16'd54101, 16'd59342, 16'd63213, 16'd13175, 16'd37843, 16'd50968, 16'd26694, 16'd47710, 16'd5241, 16'd38782, 16'd62799, 16'd17254, 16'd64056});
	test_expansion(128'h748c6bb08a44989220dc6770dbc43fd6, {16'd54395, 16'd10369, 16'd57152, 16'd63229, 16'd22444, 16'd34850, 16'd11451, 16'd34691, 16'd6101, 16'd22810, 16'd17462, 16'd10586, 16'd42780, 16'd7349, 16'd53196, 16'd30641, 16'd3557, 16'd30340, 16'd30776, 16'd4434, 16'd52727, 16'd5551, 16'd53069, 16'd36539, 16'd49226, 16'd24897});
	test_expansion(128'ha6e48bb5df6f73e79bc282b0e02c9623, {16'd15545, 16'd21101, 16'd40372, 16'd29759, 16'd41262, 16'd8609, 16'd28165, 16'd25746, 16'd62612, 16'd63981, 16'd1478, 16'd26420, 16'd55062, 16'd50753, 16'd9696, 16'd26423, 16'd31034, 16'd42357, 16'd3843, 16'd1075, 16'd63340, 16'd5848, 16'd45038, 16'd56870, 16'd42977, 16'd9597});
	test_expansion(128'h65574e40599df4f51f8217e1bd7bd3d1, {16'd44669, 16'd45943, 16'd30296, 16'd34036, 16'd29724, 16'd12963, 16'd5659, 16'd48638, 16'd43070, 16'd27790, 16'd44592, 16'd27937, 16'd63472, 16'd21986, 16'd16112, 16'd15476, 16'd1527, 16'd19975, 16'd34581, 16'd1414, 16'd10356, 16'd62687, 16'd21407, 16'd32701, 16'd7018, 16'd10643});
	test_expansion(128'hb31a69364a5bd16a0fa058bd0d93e496, {16'd17891, 16'd61626, 16'd18401, 16'd21951, 16'd49880, 16'd1528, 16'd45554, 16'd60360, 16'd8487, 16'd16677, 16'd28535, 16'd29094, 16'd1076, 16'd7344, 16'd15753, 16'd20183, 16'd17508, 16'd20006, 16'd50929, 16'd64154, 16'd13029, 16'd29040, 16'd59869, 16'd54370, 16'd44721, 16'd32788});
	test_expansion(128'hb2ae85164f2b8574fd7935bb34dc8c5b, {16'd923, 16'd4750, 16'd63551, 16'd25822, 16'd10990, 16'd60372, 16'd61106, 16'd37065, 16'd33561, 16'd57563, 16'd32286, 16'd422, 16'd6580, 16'd25765, 16'd58833, 16'd30213, 16'd52436, 16'd37853, 16'd26832, 16'd52914, 16'd27469, 16'd43318, 16'd53160, 16'd12745, 16'd28845, 16'd39895});
	test_expansion(128'hb6687d1034d05a0fe14c715738acd034, {16'd38063, 16'd53510, 16'd59876, 16'd59364, 16'd41761, 16'd59892, 16'd34346, 16'd43458, 16'd49669, 16'd40757, 16'd50067, 16'd40980, 16'd17181, 16'd25142, 16'd29214, 16'd32757, 16'd43280, 16'd28689, 16'd52716, 16'd40247, 16'd16900, 16'd33009, 16'd34606, 16'd816, 16'd62190, 16'd9367});
	test_expansion(128'h6c961b3b5816193a73f6094ef149f8d8, {16'd2994, 16'd60173, 16'd50225, 16'd55521, 16'd54583, 16'd21501, 16'd49329, 16'd7936, 16'd63455, 16'd46144, 16'd59957, 16'd55424, 16'd5762, 16'd35675, 16'd42899, 16'd33052, 16'd47342, 16'd20712, 16'd8035, 16'd26197, 16'd10841, 16'd36309, 16'd18407, 16'd49201, 16'd51793, 16'd18194});
	test_expansion(128'hed1534eea396d8e17a98bf551233b020, {16'd16167, 16'd62391, 16'd62747, 16'd34809, 16'd34837, 16'd31876, 16'd6657, 16'd60202, 16'd4389, 16'd42521, 16'd41960, 16'd44361, 16'd48692, 16'd32115, 16'd18174, 16'd24041, 16'd10047, 16'd19215, 16'd20872, 16'd31725, 16'd19831, 16'd19381, 16'd64239, 16'd52855, 16'd14387, 16'd20885});
	test_expansion(128'h363486d12e75fa114c97d4a0fdbb28bd, {16'd13891, 16'd23390, 16'd35219, 16'd2610, 16'd39313, 16'd26601, 16'd7297, 16'd54586, 16'd17337, 16'd33964, 16'd61772, 16'd9280, 16'd1780, 16'd46933, 16'd1346, 16'd17796, 16'd42617, 16'd7157, 16'd34626, 16'd13166, 16'd45244, 16'd43937, 16'd7666, 16'd57186, 16'd30961, 16'd45910});
	test_expansion(128'h51377ef7d2fa67e5261e2d4134aad1b7, {16'd26790, 16'd5601, 16'd44951, 16'd58915, 16'd58675, 16'd56285, 16'd56006, 16'd4940, 16'd7606, 16'd12203, 16'd25603, 16'd13773, 16'd19406, 16'd22380, 16'd52546, 16'd3201, 16'd14580, 16'd7120, 16'd18722, 16'd53502, 16'd51577, 16'd18033, 16'd6173, 16'd12129, 16'd16481, 16'd52911});
	test_expansion(128'h82b50fe6d9d1a70ef898c64076951f75, {16'd2648, 16'd19885, 16'd36676, 16'd60169, 16'd32230, 16'd29638, 16'd48527, 16'd57559, 16'd57622, 16'd30461, 16'd65185, 16'd63727, 16'd55637, 16'd54845, 16'd39747, 16'd51645, 16'd11951, 16'd59404, 16'd6839, 16'd54960, 16'd32269, 16'd36257, 16'd51680, 16'd53692, 16'd10581, 16'd15515});
	test_expansion(128'hc0d403e422c94851a46ba921a9bde06a, {16'd19928, 16'd6913, 16'd52816, 16'd26699, 16'd22891, 16'd3120, 16'd52652, 16'd23133, 16'd48193, 16'd29593, 16'd53753, 16'd53148, 16'd2110, 16'd46500, 16'd11120, 16'd35760, 16'd43939, 16'd62977, 16'd64786, 16'd39879, 16'd47071, 16'd33228, 16'd29552, 16'd39631, 16'd51294, 16'd32853});
	test_expansion(128'hec6b89e876446f51d11cc6dbfcd45a94, {16'd59944, 16'd22255, 16'd41802, 16'd23392, 16'd55694, 16'd30033, 16'd39363, 16'd13178, 16'd18490, 16'd26892, 16'd57036, 16'd40912, 16'd28247, 16'd50509, 16'd58798, 16'd53758, 16'd33863, 16'd21766, 16'd11475, 16'd37902, 16'd51158, 16'd47259, 16'd31857, 16'd21517, 16'd33720, 16'd31755});
	test_expansion(128'h985b9fd9043ada6524aff432e9a6f4bd, {16'd20810, 16'd18231, 16'd55489, 16'd43823, 16'd34128, 16'd10240, 16'd56174, 16'd58574, 16'd41401, 16'd22466, 16'd24610, 16'd37837, 16'd45293, 16'd27921, 16'd63827, 16'd18814, 16'd19981, 16'd8592, 16'd57374, 16'd4100, 16'd36949, 16'd41887, 16'd52738, 16'd8877, 16'd51217, 16'd34244});
	test_expansion(128'he5e11e0c6925671b3092f4e3e04d6f4c, {16'd6002, 16'd8811, 16'd54439, 16'd57343, 16'd14880, 16'd17802, 16'd62370, 16'd13437, 16'd37300, 16'd41180, 16'd5529, 16'd44372, 16'd49702, 16'd43353, 16'd50151, 16'd65397, 16'd14433, 16'd54053, 16'd37796, 16'd1171, 16'd63830, 16'd3904, 16'd31290, 16'd43397, 16'd35655, 16'd10410});
	test_expansion(128'h2d1158e390e09bea15f5152dbb4bf9fd, {16'd12853, 16'd49689, 16'd34994, 16'd56486, 16'd51986, 16'd4757, 16'd33033, 16'd6424, 16'd48917, 16'd61859, 16'd18254, 16'd53356, 16'd16550, 16'd5512, 16'd59096, 16'd61980, 16'd13560, 16'd24921, 16'd55041, 16'd64047, 16'd43946, 16'd54088, 16'd58585, 16'd59400, 16'd20894, 16'd54783});
	test_expansion(128'ha895953c13dddba40c27c0389583ead4, {16'd8893, 16'd63609, 16'd31119, 16'd64341, 16'd20701, 16'd17370, 16'd64061, 16'd35822, 16'd20633, 16'd8382, 16'd23386, 16'd25622, 16'd55826, 16'd23220, 16'd30630, 16'd21868, 16'd42833, 16'd34227, 16'd43240, 16'd36677, 16'd10849, 16'd26646, 16'd9013, 16'd63488, 16'd22613, 16'd41472});
	test_expansion(128'h9f18b84228ee13bf3c5075bf9be097bd, {16'd46036, 16'd58016, 16'd9310, 16'd52447, 16'd37316, 16'd16649, 16'd48128, 16'd57826, 16'd14337, 16'd23124, 16'd36238, 16'd28608, 16'd13733, 16'd64160, 16'd19029, 16'd63525, 16'd34418, 16'd37833, 16'd54879, 16'd22362, 16'd5242, 16'd47777, 16'd34051, 16'd24420, 16'd57021, 16'd15272});
	test_expansion(128'haf9a96bc355297d4540d600d3bb74d95, {16'd8462, 16'd31715, 16'd44930, 16'd25079, 16'd28852, 16'd8753, 16'd60594, 16'd1174, 16'd11783, 16'd28174, 16'd48352, 16'd30119, 16'd49486, 16'd33421, 16'd62511, 16'd12823, 16'd17009, 16'd21263, 16'd5579, 16'd32097, 16'd11073, 16'd50666, 16'd19170, 16'd28802, 16'd39275, 16'd4966});
	test_expansion(128'h16f926910fd9438925ed6534decdb2b3, {16'd53748, 16'd20248, 16'd24224, 16'd594, 16'd25719, 16'd27665, 16'd26857, 16'd51811, 16'd42166, 16'd23101, 16'd48298, 16'd8467, 16'd34083, 16'd62252, 16'd45553, 16'd9903, 16'd45101, 16'd26957, 16'd13696, 16'd21658, 16'd1372, 16'd22628, 16'd44992, 16'd28093, 16'd61845, 16'd34469});
	test_expansion(128'hfa2c6ccb4d7c718ab5e79a3627c2cee9, {16'd44530, 16'd28406, 16'd26452, 16'd17544, 16'd30516, 16'd2290, 16'd36891, 16'd58185, 16'd54742, 16'd37313, 16'd64532, 16'd63038, 16'd30218, 16'd38802, 16'd12748, 16'd8855, 16'd47877, 16'd19170, 16'd33004, 16'd19383, 16'd31402, 16'd13735, 16'd65315, 16'd4902, 16'd26928, 16'd59373});
	test_expansion(128'h12b54aa897c09d0f6b4814459b306bb4, {16'd36643, 16'd22115, 16'd46755, 16'd44758, 16'd63330, 16'd24645, 16'd57680, 16'd22182, 16'd9997, 16'd51816, 16'd17566, 16'd8099, 16'd25992, 16'd45625, 16'd25306, 16'd57436, 16'd17536, 16'd19135, 16'd33655, 16'd57920, 16'd6770, 16'd57679, 16'd59818, 16'd23796, 16'd55737, 16'd60206});
	test_expansion(128'ha46398a1a0255b8981de3215857ed600, {16'd12779, 16'd63380, 16'd5254, 16'd48278, 16'd29959, 16'd50389, 16'd64726, 16'd57723, 16'd20002, 16'd40082, 16'd32102, 16'd35348, 16'd8207, 16'd48986, 16'd43234, 16'd12900, 16'd11343, 16'd6325, 16'd34147, 16'd29029, 16'd28167, 16'd15024, 16'd43212, 16'd52292, 16'd29326, 16'd49922});
	test_expansion(128'h846746209d952b3d605faf97e1001495, {16'd50612, 16'd2179, 16'd26208, 16'd5330, 16'd598, 16'd60026, 16'd9502, 16'd65091, 16'd210, 16'd29554, 16'd28072, 16'd36199, 16'd14831, 16'd26160, 16'd33735, 16'd3082, 16'd1470, 16'd18484, 16'd48987, 16'd17126, 16'd57769, 16'd29731, 16'd22635, 16'd51459, 16'd48110, 16'd29516});
	test_expansion(128'h83805f4ebce2dbaa4e9cd56d317fc469, {16'd1642, 16'd13245, 16'd60480, 16'd35606, 16'd21484, 16'd62901, 16'd22619, 16'd55025, 16'd5208, 16'd1443, 16'd9668, 16'd33837, 16'd11396, 16'd61151, 16'd40020, 16'd19595, 16'd38702, 16'd10440, 16'd46861, 16'd36009, 16'd3230, 16'd51829, 16'd19294, 16'd58830, 16'd14885, 16'd20471});
	test_expansion(128'h8ea5d90a82f59e5ba3c50b608998d54a, {16'd62429, 16'd56086, 16'd11867, 16'd4047, 16'd15052, 16'd18609, 16'd56930, 16'd27851, 16'd11319, 16'd63183, 16'd38466, 16'd25999, 16'd17104, 16'd11343, 16'd20247, 16'd21260, 16'd15598, 16'd35217, 16'd53611, 16'd52934, 16'd2276, 16'd14177, 16'd4953, 16'd41311, 16'd16289, 16'd9391});
	test_expansion(128'h6a1d2226a767a7cbed143239b821c6be, {16'd9192, 16'd30339, 16'd35981, 16'd41224, 16'd13494, 16'd60570, 16'd61144, 16'd57356, 16'd14944, 16'd44991, 16'd43696, 16'd14443, 16'd18925, 16'd21956, 16'd23773, 16'd35974, 16'd53744, 16'd50244, 16'd6379, 16'd40465, 16'd12583, 16'd43741, 16'd14101, 16'd9391, 16'd63612, 16'd34313});
	test_expansion(128'ha7dfb01a5038736bfde76280f5c741ed, {16'd33271, 16'd55591, 16'd49514, 16'd17545, 16'd35851, 16'd16096, 16'd51071, 16'd21868, 16'd40397, 16'd18081, 16'd2644, 16'd7432, 16'd55949, 16'd26399, 16'd13574, 16'd20690, 16'd40184, 16'd23082, 16'd41172, 16'd23664, 16'd42685, 16'd24118, 16'd55909, 16'd26867, 16'd52864, 16'd22468});
	test_expansion(128'h076d66714dfbd24c850788dd883da50a, {16'd60889, 16'd3362, 16'd45865, 16'd37876, 16'd63978, 16'd11797, 16'd50554, 16'd60811, 16'd63417, 16'd20760, 16'd4165, 16'd35099, 16'd43956, 16'd33164, 16'd62952, 16'd4801, 16'd19576, 16'd47790, 16'd58165, 16'd24799, 16'd45806, 16'd37922, 16'd30903, 16'd41530, 16'd35314, 16'd52081});
	test_expansion(128'h4c9f74be290c0ca45142147594e53e88, {16'd12307, 16'd42015, 16'd59464, 16'd7521, 16'd44434, 16'd15008, 16'd52685, 16'd28432, 16'd32324, 16'd1664, 16'd7152, 16'd23987, 16'd58782, 16'd7417, 16'd30545, 16'd32820, 16'd44965, 16'd54184, 16'd55950, 16'd4953, 16'd55064, 16'd44996, 16'd60945, 16'd44349, 16'd43640, 16'd40630});
	test_expansion(128'h196e0d8b2c666601b7b3984c5eb6442f, {16'd1846, 16'd2749, 16'd33902, 16'd30225, 16'd25094, 16'd56144, 16'd29395, 16'd44253, 16'd7923, 16'd47056, 16'd57291, 16'd7070, 16'd29604, 16'd61033, 16'd25271, 16'd61725, 16'd4966, 16'd39200, 16'd6334, 16'd56202, 16'd18761, 16'd38112, 16'd21741, 16'd1985, 16'd8802, 16'd31403});
	test_expansion(128'h6c4073da8ef1c4bc65c705e1a301a3ea, {16'd33141, 16'd47364, 16'd57147, 16'd56844, 16'd5335, 16'd42088, 16'd34472, 16'd28414, 16'd62994, 16'd44809, 16'd49308, 16'd20714, 16'd52952, 16'd38394, 16'd43413, 16'd60494, 16'd48711, 16'd53706, 16'd25013, 16'd49586, 16'd49789, 16'd40735, 16'd49754, 16'd23066, 16'd42557, 16'd60476});
	test_expansion(128'heda675019ff82de8133630383dbe7d59, {16'd39624, 16'd38520, 16'd29349, 16'd8929, 16'd61638, 16'd55231, 16'd38174, 16'd7334, 16'd44117, 16'd1953, 16'd62865, 16'd42798, 16'd49209, 16'd6280, 16'd54040, 16'd15829, 16'd36087, 16'd63267, 16'd7959, 16'd47196, 16'd25943, 16'd22833, 16'd35478, 16'd36381, 16'd64009, 16'd27428});
	test_expansion(128'h35b6395eea5fded1526669cbb3a28058, {16'd33096, 16'd42235, 16'd1598, 16'd5981, 16'd54404, 16'd20338, 16'd17046, 16'd12962, 16'd55939, 16'd44398, 16'd27606, 16'd43649, 16'd46927, 16'd39183, 16'd42546, 16'd37031, 16'd22343, 16'd46549, 16'd40566, 16'd8550, 16'd1779, 16'd60163, 16'd53299, 16'd42180, 16'd59628, 16'd61389});
	test_expansion(128'h58560457f841c82130b837bcc01398dd, {16'd45304, 16'd11005, 16'd61872, 16'd34560, 16'd13304, 16'd37923, 16'd49984, 16'd25217, 16'd6210, 16'd37492, 16'd5198, 16'd40612, 16'd7814, 16'd19593, 16'd8558, 16'd61147, 16'd56171, 16'd31403, 16'd16364, 16'd33047, 16'd29756, 16'd10984, 16'd51643, 16'd23782, 16'd32725, 16'd63920});
	test_expansion(128'h6bbd73d33974c7274669dcaea302b278, {16'd48189, 16'd35323, 16'd52001, 16'd16354, 16'd7905, 16'd62857, 16'd60968, 16'd10196, 16'd39825, 16'd286, 16'd46576, 16'd29866, 16'd5813, 16'd32935, 16'd37584, 16'd44496, 16'd15289, 16'd50450, 16'd39682, 16'd32071, 16'd49503, 16'd51016, 16'd3613, 16'd49648, 16'd49486, 16'd22442});
	test_expansion(128'h5be543bfdc17917ce21bec8d0e4c9d12, {16'd19082, 16'd64346, 16'd30306, 16'd7122, 16'd36235, 16'd18551, 16'd29361, 16'd8245, 16'd54934, 16'd57056, 16'd53549, 16'd1186, 16'd12659, 16'd47753, 16'd1430, 16'd14304, 16'd68, 16'd26863, 16'd41628, 16'd41418, 16'd23801, 16'd20577, 16'd8269, 16'd52667, 16'd23840, 16'd49151});
	test_expansion(128'h59f8959a1e72467b3caf14e72135a20d, {16'd55968, 16'd34457, 16'd55856, 16'd17954, 16'd35097, 16'd6346, 16'd48299, 16'd38774, 16'd26352, 16'd4651, 16'd35501, 16'd52261, 16'd21317, 16'd25933, 16'd34061, 16'd15698, 16'd20821, 16'd48512, 16'd48960, 16'd51860, 16'd33766, 16'd64929, 16'd43115, 16'd20391, 16'd43682, 16'd40721});
	test_expansion(128'h6cc44cdd358a47cd0a8edbc0f974b74d, {16'd39955, 16'd5987, 16'd30948, 16'd33235, 16'd3750, 16'd32077, 16'd46166, 16'd63021, 16'd14018, 16'd63697, 16'd27731, 16'd59905, 16'd55783, 16'd40268, 16'd23958, 16'd11463, 16'd29811, 16'd12359, 16'd48830, 16'd54058, 16'd14148, 16'd29790, 16'd7804, 16'd47143, 16'd49358, 16'd59541});
	test_expansion(128'he9b4fc1caf15b4956df24542620e298f, {16'd63209, 16'd25098, 16'd49409, 16'd35640, 16'd49470, 16'd33185, 16'd14353, 16'd30150, 16'd6435, 16'd39965, 16'd27437, 16'd3604, 16'd9896, 16'd48893, 16'd37939, 16'd50188, 16'd15161, 16'd28235, 16'd63349, 16'd48130, 16'd49576, 16'd15760, 16'd57562, 16'd37485, 16'd60335, 16'd5619});
	test_expansion(128'hb29d77a46d95e0ad384b6fd10bd3b5ce, {16'd23522, 16'd15574, 16'd16832, 16'd24798, 16'd33961, 16'd33812, 16'd23286, 16'd63379, 16'd43802, 16'd20144, 16'd59447, 16'd17508, 16'd35746, 16'd61795, 16'd60787, 16'd4578, 16'd5568, 16'd10749, 16'd42179, 16'd42298, 16'd16970, 16'd56867, 16'd39754, 16'd27074, 16'd39973, 16'd61371});
	test_expansion(128'hb8bdd90affad31adf7d916fc58238da8, {16'd55174, 16'd952, 16'd13042, 16'd39002, 16'd62152, 16'd53343, 16'd24516, 16'd36499, 16'd35699, 16'd57821, 16'd25629, 16'd15485, 16'd31592, 16'd45531, 16'd13473, 16'd23961, 16'd45411, 16'd47839, 16'd29904, 16'd63706, 16'd3896, 16'd30539, 16'd48529, 16'd10010, 16'd48934, 16'd45776});
	test_expansion(128'h9025079abb7979d74432d18ca1374677, {16'd9100, 16'd18450, 16'd37987, 16'd3954, 16'd31365, 16'd38369, 16'd41817, 16'd4039, 16'd53319, 16'd27468, 16'd2041, 16'd49667, 16'd2680, 16'd36183, 16'd33149, 16'd17061, 16'd5190, 16'd40533, 16'd4553, 16'd46651, 16'd6007, 16'd21358, 16'd18827, 16'd31603, 16'd8354, 16'd15418});
	test_expansion(128'h2e24310e3078995a29672caa6250f5d6, {16'd2896, 16'd21111, 16'd46788, 16'd47667, 16'd24554, 16'd11846, 16'd26026, 16'd42648, 16'd65510, 16'd12253, 16'd54109, 16'd18633, 16'd49122, 16'd2362, 16'd21315, 16'd8594, 16'd30053, 16'd28706, 16'd59288, 16'd61936, 16'd64496, 16'd4027, 16'd31073, 16'd42876, 16'd27645, 16'd9924});
	test_expansion(128'h8bfb58a1de88228be72e826e5daffeb6, {16'd6128, 16'd33466, 16'd22923, 16'd6294, 16'd35395, 16'd15362, 16'd2870, 16'd34196, 16'd11093, 16'd28473, 16'd10606, 16'd711, 16'd25950, 16'd4375, 16'd32119, 16'd43011, 16'd29593, 16'd36612, 16'd10158, 16'd1540, 16'd54586, 16'd35997, 16'd45598, 16'd37679, 16'd20743, 16'd62922});
	test_expansion(128'hd114ffd6f66c7d82ab42d31a8bb9ab0e, {16'd2822, 16'd51002, 16'd32790, 16'd26759, 16'd2409, 16'd37227, 16'd51773, 16'd32371, 16'd57893, 16'd64860, 16'd2436, 16'd61574, 16'd391, 16'd46512, 16'd53112, 16'd65158, 16'd25249, 16'd7619, 16'd62190, 16'd57597, 16'd51022, 16'd45807, 16'd46310, 16'd39786, 16'd28236, 16'd19735});
	test_expansion(128'h74d8936f1025a58d4e1852a28ca5245d, {16'd37028, 16'd5649, 16'd46279, 16'd22438, 16'd23968, 16'd7026, 16'd54098, 16'd57127, 16'd5470, 16'd29922, 16'd60024, 16'd31269, 16'd54709, 16'd1066, 16'd55124, 16'd37662, 16'd9357, 16'd53849, 16'd34754, 16'd35749, 16'd34325, 16'd64580, 16'd44939, 16'd59548, 16'd58402, 16'd25317});
	test_expansion(128'hc7a6ba0176bcc3920409d10cfda540fa, {16'd52091, 16'd57454, 16'd23120, 16'd27619, 16'd16100, 16'd13928, 16'd54472, 16'd39374, 16'd7602, 16'd6411, 16'd17219, 16'd19759, 16'd19580, 16'd44734, 16'd43484, 16'd66, 16'd10900, 16'd59751, 16'd3811, 16'd17257, 16'd50785, 16'd38453, 16'd28457, 16'd41797, 16'd49130, 16'd46206});
	test_expansion(128'h4b79927a49cf932ba6800e1fdbdeeeb7, {16'd12289, 16'd16718, 16'd61119, 16'd44816, 16'd24969, 16'd2330, 16'd2685, 16'd7110, 16'd29936, 16'd35003, 16'd51741, 16'd22421, 16'd17225, 16'd57780, 16'd1048, 16'd15787, 16'd32470, 16'd1727, 16'd11623, 16'd22870, 16'd10813, 16'd60412, 16'd40754, 16'd35199, 16'd32436, 16'd2208});
	test_expansion(128'h868247dd78631eb18042d03b640674cf, {16'd10633, 16'd6694, 16'd34181, 16'd1872, 16'd25973, 16'd62033, 16'd44542, 16'd50257, 16'd36779, 16'd44057, 16'd39849, 16'd43350, 16'd65237, 16'd27955, 16'd24816, 16'd56465, 16'd64296, 16'd56096, 16'd49032, 16'd8352, 16'd22958, 16'd13268, 16'd22654, 16'd64390, 16'd5116, 16'd3725});
	test_expansion(128'h3cf7a144666c16b155ca98cee7e41288, {16'd55775, 16'd48786, 16'd64780, 16'd10999, 16'd17472, 16'd31538, 16'd761, 16'd9566, 16'd45260, 16'd46104, 16'd4972, 16'd49519, 16'd17809, 16'd5967, 16'd49153, 16'd12634, 16'd61813, 16'd17176, 16'd34986, 16'd3573, 16'd4354, 16'd44546, 16'd32796, 16'd56728, 16'd29978, 16'd29629});
	test_expansion(128'h3d6428bf254a2e2ded633c0dd75a4f6b, {16'd3131, 16'd3967, 16'd60004, 16'd4320, 16'd23896, 16'd60989, 16'd16532, 16'd34854, 16'd54216, 16'd49482, 16'd7513, 16'd9819, 16'd57538, 16'd23603, 16'd35896, 16'd30689, 16'd61083, 16'd13291, 16'd13067, 16'd29807, 16'd62190, 16'd59415, 16'd10976, 16'd17176, 16'd44479, 16'd65141});
	test_expansion(128'h0a4996c0bf476f7b83b466e2fd25a445, {16'd1780, 16'd14344, 16'd21911, 16'd27440, 16'd36124, 16'd26533, 16'd37280, 16'd35981, 16'd26054, 16'd4352, 16'd41468, 16'd32837, 16'd50386, 16'd59939, 16'd2444, 16'd46959, 16'd62561, 16'd11090, 16'd50632, 16'd30313, 16'd25361, 16'd52476, 16'd27690, 16'd36074, 16'd46817, 16'd25740});
	test_expansion(128'hec3544de8e87730bb852f97894a79b04, {16'd6357, 16'd24082, 16'd11555, 16'd12909, 16'd20938, 16'd37530, 16'd41008, 16'd7388, 16'd30107, 16'd34873, 16'd50903, 16'd7921, 16'd58299, 16'd18066, 16'd44273, 16'd1639, 16'd58698, 16'd17643, 16'd34747, 16'd8967, 16'd55625, 16'd39088, 16'd61059, 16'd24508, 16'd4922, 16'd62431});
	test_expansion(128'hed89a975ea2664ddcdeef34bdde2c1e2, {16'd4823, 16'd54471, 16'd62218, 16'd3903, 16'd25200, 16'd48130, 16'd63231, 16'd41627, 16'd41000, 16'd63202, 16'd63647, 16'd23616, 16'd53361, 16'd38648, 16'd20101, 16'd7731, 16'd36999, 16'd27, 16'd52588, 16'd55761, 16'd64587, 16'd9001, 16'd44878, 16'd16498, 16'd29939, 16'd248});
	test_expansion(128'h0b394858aaba209eb22aba5df0dc1da9, {16'd10066, 16'd23254, 16'd44561, 16'd11606, 16'd61080, 16'd30188, 16'd35730, 16'd40916, 16'd60119, 16'd3850, 16'd32850, 16'd30512, 16'd31712, 16'd14, 16'd50890, 16'd57738, 16'd22184, 16'd55693, 16'd45462, 16'd45445, 16'd42786, 16'd49654, 16'd61942, 16'd12932, 16'd11779, 16'd41327});
	test_expansion(128'h6931291bc2a0cd9258e5d6d6f466408e, {16'd116, 16'd37149, 16'd12879, 16'd49699, 16'd25566, 16'd30619, 16'd14872, 16'd6709, 16'd31031, 16'd34696, 16'd62361, 16'd24092, 16'd23469, 16'd63620, 16'd55331, 16'd5524, 16'd35575, 16'd49587, 16'd55879, 16'd34196, 16'd11781, 16'd4569, 16'd53586, 16'd54024, 16'd25569, 16'd3020});
	test_expansion(128'h6980534af6b9249af5009c833b27e457, {16'd7384, 16'd52587, 16'd53083, 16'd48136, 16'd5734, 16'd4614, 16'd32884, 16'd23778, 16'd51136, 16'd18669, 16'd8242, 16'd52565, 16'd53505, 16'd35257, 16'd61537, 16'd49680, 16'd46117, 16'd57849, 16'd10686, 16'd28621, 16'd46374, 16'd48950, 16'd39372, 16'd7149, 16'd54948, 16'd19380});
	test_expansion(128'h85f6a1b9979a8fe052f133a8b8c8113a, {16'd37132, 16'd32913, 16'd48238, 16'd58634, 16'd56696, 16'd30588, 16'd34146, 16'd48808, 16'd18001, 16'd5443, 16'd4577, 16'd5659, 16'd43641, 16'd21535, 16'd9117, 16'd61954, 16'd54933, 16'd5148, 16'd41280, 16'd59053, 16'd10561, 16'd60104, 16'd11434, 16'd24408, 16'd59355, 16'd15474});
	test_expansion(128'h3f393e9de5e74e0eccefb0ef549eedc3, {16'd13072, 16'd18160, 16'd61955, 16'd1513, 16'd18546, 16'd4843, 16'd56215, 16'd60044, 16'd53706, 16'd57255, 16'd8578, 16'd2511, 16'd15294, 16'd31953, 16'd41319, 16'd40153, 16'd49759, 16'd47746, 16'd1919, 16'd50746, 16'd16996, 16'd4904, 16'd53437, 16'd29973, 16'd37346, 16'd33113});
	test_expansion(128'h9c81dcff5b01b3fcc0a6949039c9cc62, {16'd57505, 16'd53020, 16'd31187, 16'd23523, 16'd37078, 16'd45035, 16'd62611, 16'd19334, 16'd46005, 16'd55903, 16'd6631, 16'd4730, 16'd62375, 16'd33701, 16'd22789, 16'd17043, 16'd61812, 16'd26757, 16'd13450, 16'd51306, 16'd15820, 16'd39401, 16'd23273, 16'd58071, 16'd63090, 16'd18779});
	test_expansion(128'h0b715de47e751e1a44b44fd10e9d4364, {16'd64057, 16'd63365, 16'd51990, 16'd38269, 16'd35408, 16'd33753, 16'd5278, 16'd22848, 16'd48908, 16'd55982, 16'd9423, 16'd53604, 16'd33070, 16'd56162, 16'd14871, 16'd301, 16'd439, 16'd35361, 16'd19987, 16'd62995, 16'd32704, 16'd248, 16'd40931, 16'd58538, 16'd32327, 16'd44878});
	test_expansion(128'h54288b80c5b846fb371373a0c429afe8, {16'd29247, 16'd62451, 16'd39823, 16'd33933, 16'd34744, 16'd25353, 16'd25998, 16'd12424, 16'd10353, 16'd48091, 16'd31114, 16'd36420, 16'd9640, 16'd8740, 16'd11710, 16'd21627, 16'd64478, 16'd7624, 16'd27569, 16'd64486, 16'd64859, 16'd16652, 16'd39008, 16'd33441, 16'd27585, 16'd2315});
	test_expansion(128'h03bd5f8c315a61018f29f99074f98332, {16'd17071, 16'd28550, 16'd36765, 16'd7590, 16'd21357, 16'd40190, 16'd46295, 16'd26716, 16'd36987, 16'd26436, 16'd2555, 16'd64490, 16'd47707, 16'd6898, 16'd6995, 16'd44954, 16'd44849, 16'd10380, 16'd59117, 16'd63108, 16'd26907, 16'd58160, 16'd29017, 16'd28967, 16'd10212, 16'd55544});
	test_expansion(128'h2dbaee5b9e4d5118c80ddefcf0fef35c, {16'd58660, 16'd7015, 16'd44042, 16'd34938, 16'd32455, 16'd32064, 16'd59817, 16'd50712, 16'd49727, 16'd25963, 16'd45274, 16'd30950, 16'd51087, 16'd63269, 16'd14824, 16'd1062, 16'd61854, 16'd21451, 16'd1092, 16'd36860, 16'd14301, 16'd16919, 16'd7886, 16'd53508, 16'd14156, 16'd64404});
	test_expansion(128'h6be2d42e4b7496e580369c94a2403871, {16'd26829, 16'd7229, 16'd2044, 16'd60512, 16'd29662, 16'd78, 16'd40659, 16'd64699, 16'd59428, 16'd49378, 16'd55192, 16'd40773, 16'd31897, 16'd23543, 16'd19575, 16'd63298, 16'd49265, 16'd16702, 16'd7767, 16'd42147, 16'd56739, 16'd43591, 16'd64824, 16'd20348, 16'd52748, 16'd59369});
	test_expansion(128'hcbfdaea4f7c5ae9f6dea266448ef6bba, {16'd32266, 16'd32729, 16'd56854, 16'd8088, 16'd55900, 16'd11542, 16'd48474, 16'd55937, 16'd22929, 16'd33831, 16'd63124, 16'd42744, 16'd17198, 16'd14234, 16'd17479, 16'd48344, 16'd45228, 16'd41950, 16'd17365, 16'd21671, 16'd15454, 16'd26713, 16'd39986, 16'd31893, 16'd57600, 16'd1609});
	test_expansion(128'h4edd4b6adcd8318fe1d53076ea21c251, {16'd16381, 16'd37705, 16'd33910, 16'd46379, 16'd59685, 16'd43025, 16'd57400, 16'd38157, 16'd9039, 16'd40113, 16'd44122, 16'd7106, 16'd25300, 16'd16556, 16'd25094, 16'd60843, 16'd25638, 16'd56433, 16'd59520, 16'd53083, 16'd14930, 16'd8696, 16'd45631, 16'd38034, 16'd38310, 16'd41296});
	test_expansion(128'h453cb767ebe1ea4879cd21708b09ac9e, {16'd35468, 16'd27896, 16'd14508, 16'd32640, 16'd52276, 16'd54283, 16'd17817, 16'd31988, 16'd55836, 16'd6994, 16'd18277, 16'd41182, 16'd63501, 16'd64254, 16'd10016, 16'd32773, 16'd6844, 16'd60044, 16'd28004, 16'd54525, 16'd19813, 16'd60408, 16'd9776, 16'd1410, 16'd56176, 16'd59123});
	test_expansion(128'h73befb551e61c2f449d958bd783f2528, {16'd21375, 16'd12976, 16'd21314, 16'd9393, 16'd14381, 16'd33446, 16'd22543, 16'd55760, 16'd39983, 16'd49770, 16'd62269, 16'd51821, 16'd21825, 16'd56523, 16'd36475, 16'd26337, 16'd52271, 16'd23758, 16'd39776, 16'd27699, 16'd1585, 16'd49906, 16'd54219, 16'd40233, 16'd54730, 16'd46468});
	test_expansion(128'hc612bf3e9ba99c5454ffcef85618d444, {16'd3078, 16'd56907, 16'd18151, 16'd61319, 16'd64531, 16'd11609, 16'd45416, 16'd30038, 16'd12979, 16'd34769, 16'd16862, 16'd6041, 16'd51473, 16'd19670, 16'd53611, 16'd41972, 16'd65501, 16'd13518, 16'd32445, 16'd15021, 16'd4062, 16'd63069, 16'd47065, 16'd43406, 16'd52855, 16'd32069});
	test_expansion(128'h1f10e1f502ade1c22fe1bf517304a060, {16'd59186, 16'd56909, 16'd48680, 16'd38019, 16'd45836, 16'd12359, 16'd44225, 16'd4881, 16'd42697, 16'd31233, 16'd6678, 16'd8036, 16'd28364, 16'd37000, 16'd21543, 16'd59205, 16'd42558, 16'd31339, 16'd47001, 16'd39727, 16'd7393, 16'd55435, 16'd60202, 16'd51117, 16'd63135, 16'd14368});
	test_expansion(128'hc82719cdfeea2b6aefb59bd0ef4579b6, {16'd51560, 16'd4006, 16'd16514, 16'd41754, 16'd29637, 16'd28890, 16'd12875, 16'd17677, 16'd29537, 16'd31374, 16'd36774, 16'd50611, 16'd49562, 16'd44200, 16'd33377, 16'd57231, 16'd11209, 16'd24785, 16'd63004, 16'd38951, 16'd42881, 16'd49711, 16'd39507, 16'd44571, 16'd62133, 16'd45808});
	test_expansion(128'ha8ece4261fd04c88a1029d3477319c5d, {16'd18027, 16'd47075, 16'd28590, 16'd25443, 16'd54660, 16'd34749, 16'd64917, 16'd30021, 16'd60299, 16'd29414, 16'd59136, 16'd31509, 16'd27378, 16'd5105, 16'd63825, 16'd63277, 16'd51072, 16'd37775, 16'd23567, 16'd50013, 16'd5937, 16'd15126, 16'd27963, 16'd45869, 16'd46402, 16'd41963});
	test_expansion(128'hcce1d031e6cd92b9a75e495bf27ac597, {16'd14250, 16'd53633, 16'd30729, 16'd17429, 16'd51337, 16'd10082, 16'd60745, 16'd2996, 16'd39971, 16'd7617, 16'd38466, 16'd7189, 16'd51552, 16'd1887, 16'd47393, 16'd20407, 16'd99, 16'd31888, 16'd16970, 16'd52798, 16'd7364, 16'd10061, 16'd52957, 16'd44200, 16'd6490, 16'd58495});
	test_expansion(128'h6c6397d7ab2981aba6fa487133bb7bce, {16'd33101, 16'd14782, 16'd18591, 16'd20350, 16'd38469, 16'd11549, 16'd10830, 16'd43199, 16'd30144, 16'd3969, 16'd48770, 16'd1993, 16'd42369, 16'd2007, 16'd6038, 16'd14880, 16'd50028, 16'd30311, 16'd4868, 16'd36369, 16'd3298, 16'd324, 16'd56833, 16'd31876, 16'd21958, 16'd4746});
	test_expansion(128'habaed8c29a2cd2ff1723d4f99c179766, {16'd22720, 16'd42427, 16'd36014, 16'd53740, 16'd38507, 16'd50054, 16'd61922, 16'd10527, 16'd31053, 16'd63773, 16'd47296, 16'd12803, 16'd53894, 16'd10558, 16'd53762, 16'd928, 16'd21943, 16'd51109, 16'd45210, 16'd31516, 16'd24727, 16'd56885, 16'd41622, 16'd35305, 16'd46612, 16'd7336});
	test_expansion(128'hca11e3ba9cf204cdd38543570752fc78, {16'd22850, 16'd34246, 16'd4939, 16'd31300, 16'd28371, 16'd36271, 16'd24827, 16'd324, 16'd15815, 16'd53489, 16'd7757, 16'd2000, 16'd54653, 16'd10920, 16'd2438, 16'd18333, 16'd37145, 16'd14192, 16'd51187, 16'd63927, 16'd11516, 16'd10345, 16'd12597, 16'd21332, 16'd36493, 16'd41604});
	test_expansion(128'h92f95a54b57f39784fa00cb5cd81c8c2, {16'd48909, 16'd35404, 16'd25785, 16'd36971, 16'd15678, 16'd23403, 16'd963, 16'd58551, 16'd42188, 16'd62917, 16'd23110, 16'd38780, 16'd61447, 16'd56236, 16'd24119, 16'd23537, 16'd40714, 16'd52161, 16'd61102, 16'd58653, 16'd1574, 16'd17822, 16'd46985, 16'd3203, 16'd57353, 16'd29582});
	test_expansion(128'hcdf17e1abd99886516bd116ae671b3f9, {16'd47109, 16'd21162, 16'd41595, 16'd34495, 16'd41635, 16'd1094, 16'd27953, 16'd2770, 16'd44571, 16'd9591, 16'd5809, 16'd4822, 16'd64147, 16'd21316, 16'd45225, 16'd20320, 16'd51430, 16'd53842, 16'd24753, 16'd35199, 16'd2548, 16'd18868, 16'd32980, 16'd27192, 16'd24887, 16'd60133});
	test_expansion(128'h6c149fea81078e668eea556f8dabcfa7, {16'd56677, 16'd57094, 16'd58315, 16'd38789, 16'd6007, 16'd5245, 16'd43102, 16'd12573, 16'd8003, 16'd40603, 16'd16746, 16'd38995, 16'd9317, 16'd49454, 16'd10078, 16'd22322, 16'd3954, 16'd52387, 16'd6580, 16'd21383, 16'd23266, 16'd33449, 16'd20301, 16'd22317, 16'd17069, 16'd54279});
	test_expansion(128'hef503784f13a110e56beb6ac41eac0b0, {16'd47147, 16'd16388, 16'd11439, 16'd17250, 16'd27136, 16'd48803, 16'd58296, 16'd16484, 16'd31010, 16'd46016, 16'd38314, 16'd55651, 16'd57504, 16'd3578, 16'd33643, 16'd10376, 16'd17893, 16'd47119, 16'd39423, 16'd63498, 16'd3817, 16'd30044, 16'd40736, 16'd11509, 16'd43574, 16'd2432});
	test_expansion(128'hc96403d4a4bfb420d911c24156b0c981, {16'd64480, 16'd15982, 16'd21971, 16'd51393, 16'd49657, 16'd40490, 16'd44115, 16'd18856, 16'd11398, 16'd18301, 16'd18348, 16'd62886, 16'd8077, 16'd28693, 16'd7231, 16'd45106, 16'd13038, 16'd62364, 16'd16143, 16'd35406, 16'd60279, 16'd27741, 16'd16065, 16'd29247, 16'd38205, 16'd41858});
	test_expansion(128'hdb70e84cf331ed4f1b184a1a9c05bb9b, {16'd5679, 16'd51808, 16'd51097, 16'd26721, 16'd62508, 16'd25996, 16'd35547, 16'd56106, 16'd30488, 16'd27167, 16'd63240, 16'd48967, 16'd65170, 16'd65462, 16'd41028, 16'd25618, 16'd28187, 16'd2685, 16'd30932, 16'd54354, 16'd30606, 16'd30589, 16'd18497, 16'd13392, 16'd36216, 16'd9790});
	test_expansion(128'h3194dee2391c60fa72929a2c5938b3e5, {16'd10358, 16'd27392, 16'd44310, 16'd62245, 16'd60598, 16'd33690, 16'd64728, 16'd28687, 16'd13775, 16'd29063, 16'd2715, 16'd45645, 16'd19246, 16'd23771, 16'd11354, 16'd38191, 16'd1482, 16'd29544, 16'd58546, 16'd21565, 16'd38099, 16'd20951, 16'd52564, 16'd40209, 16'd9627, 16'd34783});
	test_expansion(128'h348236a8cf1cfc125eb3259e82c81cb5, {16'd30759, 16'd39054, 16'd60604, 16'd22557, 16'd42106, 16'd57796, 16'd29818, 16'd55950, 16'd6460, 16'd16404, 16'd4901, 16'd20022, 16'd32222, 16'd34661, 16'd61009, 16'd26666, 16'd31990, 16'd43216, 16'd50658, 16'd22589, 16'd65461, 16'd27463, 16'd64793, 16'd59429, 16'd41306, 16'd46432});
	test_expansion(128'h53a744783d3ce97af9046c3ad52eaf3c, {16'd53008, 16'd4437, 16'd26920, 16'd28407, 16'd63030, 16'd14988, 16'd48786, 16'd19080, 16'd65004, 16'd52288, 16'd59589, 16'd25509, 16'd40668, 16'd6660, 16'd45896, 16'd60028, 16'd62159, 16'd63501, 16'd31167, 16'd62495, 16'd53304, 16'd16545, 16'd47439, 16'd3840, 16'd62867, 16'd8412});
	test_expansion(128'hddbcd51109542ba83776c59984a823a3, {16'd49285, 16'd61336, 16'd16387, 16'd62674, 16'd30734, 16'd61237, 16'd39944, 16'd19711, 16'd20141, 16'd26119, 16'd35279, 16'd58364, 16'd28029, 16'd10690, 16'd36494, 16'd15895, 16'd60522, 16'd16245, 16'd3149, 16'd37928, 16'd7119, 16'd29077, 16'd3111, 16'd54016, 16'd10866, 16'd65115});
	test_expansion(128'h13c5efc2f0e51d83e7de6e2d6faa6555, {16'd8079, 16'd25968, 16'd36093, 16'd11351, 16'd15303, 16'd40670, 16'd34888, 16'd47986, 16'd64505, 16'd62594, 16'd45876, 16'd8012, 16'd62112, 16'd16908, 16'd32319, 16'd32354, 16'd3091, 16'd44651, 16'd39085, 16'd62326, 16'd52850, 16'd43930, 16'd43663, 16'd999, 16'd34109, 16'd7070});
	test_expansion(128'h9d62e677f407825db1f742749282f6e7, {16'd49646, 16'd28072, 16'd11525, 16'd4914, 16'd54553, 16'd51156, 16'd21169, 16'd51135, 16'd15302, 16'd12658, 16'd44390, 16'd30366, 16'd34268, 16'd32466, 16'd26047, 16'd27716, 16'd16335, 16'd36141, 16'd20969, 16'd26067, 16'd63581, 16'd27326, 16'd21491, 16'd40856, 16'd57017, 16'd52199});
	test_expansion(128'h583bf418a45c5eedb35ba1f6e2d3f0d9, {16'd61025, 16'd26560, 16'd51275, 16'd10791, 16'd8382, 16'd47501, 16'd9501, 16'd40445, 16'd59556, 16'd57100, 16'd31597, 16'd59859, 16'd2030, 16'd59339, 16'd26626, 16'd20772, 16'd50797, 16'd46281, 16'd27001, 16'd24643, 16'd22233, 16'd49251, 16'd57942, 16'd33933, 16'd55697, 16'd47808});
	test_expansion(128'h0c1b0f4d8f6cff2ff9fd091970ab51d0, {16'd35538, 16'd47424, 16'd48344, 16'd21470, 16'd64983, 16'd53857, 16'd50446, 16'd11095, 16'd21060, 16'd24369, 16'd60100, 16'd52713, 16'd38016, 16'd6812, 16'd34025, 16'd7059, 16'd21595, 16'd26155, 16'd37384, 16'd4821, 16'd15124, 16'd17543, 16'd54661, 16'd24880, 16'd47015, 16'd43867});
	test_expansion(128'h18b085708cd84941ea139c1242e75605, {16'd41686, 16'd47462, 16'd17617, 16'd23708, 16'd39739, 16'd38532, 16'd24707, 16'd47853, 16'd23114, 16'd21097, 16'd42621, 16'd11548, 16'd43731, 16'd31993, 16'd17785, 16'd18734, 16'd28649, 16'd54800, 16'd32665, 16'd43593, 16'd17852, 16'd28240, 16'd5806, 16'd60911, 16'd26668, 16'd12691});
	test_expansion(128'hde6039cfb1d576dc7c15e3ef75351f43, {16'd26180, 16'd50629, 16'd41834, 16'd33351, 16'd63075, 16'd29074, 16'd3419, 16'd43703, 16'd1617, 16'd41416, 16'd13095, 16'd18901, 16'd20764, 16'd27156, 16'd34759, 16'd6901, 16'd57714, 16'd23334, 16'd50841, 16'd65366, 16'd17547, 16'd39270, 16'd38036, 16'd21756, 16'd16761, 16'd12587});
	test_expansion(128'he569a76337e3d803be337a14c239a935, {16'd25651, 16'd26083, 16'd29696, 16'd3140, 16'd37885, 16'd11161, 16'd1800, 16'd36954, 16'd25489, 16'd12331, 16'd55429, 16'd49431, 16'd14374, 16'd52772, 16'd33443, 16'd7067, 16'd5336, 16'd29840, 16'd27588, 16'd58607, 16'd17307, 16'd54810, 16'd44156, 16'd19169, 16'd54335, 16'd48682});
	test_expansion(128'hc9c90d6dfd67723288e5cc73e7dfa86f, {16'd27309, 16'd3792, 16'd49079, 16'd17724, 16'd17829, 16'd13016, 16'd11146, 16'd17790, 16'd47369, 16'd28751, 16'd57927, 16'd41715, 16'd44129, 16'd368, 16'd50506, 16'd24898, 16'd59446, 16'd40124, 16'd50528, 16'd61244, 16'd18255, 16'd4959, 16'd26977, 16'd10069, 16'd64309, 16'd51003});
	test_expansion(128'h987ae09089560c29e980000a8cd7e966, {16'd57643, 16'd12571, 16'd44737, 16'd5833, 16'd55099, 16'd16, 16'd58652, 16'd29972, 16'd60474, 16'd44672, 16'd22528, 16'd6741, 16'd58422, 16'd54271, 16'd34168, 16'd17500, 16'd60917, 16'd36665, 16'd51563, 16'd5951, 16'd7979, 16'd17180, 16'd50653, 16'd58289, 16'd27757, 16'd19351});
	test_expansion(128'hd84bfdf036f657a8e38f9f540471458d, {16'd61472, 16'd46341, 16'd49441, 16'd4468, 16'd22882, 16'd53821, 16'd370, 16'd37619, 16'd31038, 16'd30482, 16'd21362, 16'd28504, 16'd48210, 16'd40045, 16'd48273, 16'd50072, 16'd50587, 16'd13082, 16'd12248, 16'd35473, 16'd62961, 16'd26750, 16'd38878, 16'd34785, 16'd63750, 16'd52737});
	test_expansion(128'h3a5dddd7a3d8c691d4536c5f68ce3ad8, {16'd58366, 16'd51181, 16'd26669, 16'd47676, 16'd3439, 16'd11164, 16'd17197, 16'd22783, 16'd12793, 16'd41940, 16'd28118, 16'd12101, 16'd24131, 16'd29781, 16'd47080, 16'd37398, 16'd21578, 16'd2709, 16'd19850, 16'd39613, 16'd41406, 16'd56782, 16'd37419, 16'd7406, 16'd52363, 16'd53384});
	test_expansion(128'h88e008a0488ce9e66d70a2bdc9b238e6, {16'd176, 16'd2386, 16'd60529, 16'd38124, 16'd58360, 16'd26886, 16'd29197, 16'd41955, 16'd41429, 16'd1926, 16'd34071, 16'd13607, 16'd42698, 16'd7129, 16'd54711, 16'd45170, 16'd1081, 16'd43576, 16'd47781, 16'd6072, 16'd1601, 16'd8675, 16'd20473, 16'd13590, 16'd28098, 16'd3092});
	test_expansion(128'h2dec6d304419b9a860d45e8996d16397, {16'd12306, 16'd1444, 16'd3035, 16'd52568, 16'd9739, 16'd41626, 16'd23095, 16'd21533, 16'd7869, 16'd7305, 16'd52774, 16'd24978, 16'd8357, 16'd5617, 16'd49900, 16'd52251, 16'd29056, 16'd33993, 16'd42282, 16'd1332, 16'd63748, 16'd54116, 16'd32432, 16'd28700, 16'd65434, 16'd30209});
	test_expansion(128'h4b8f888b9e70a64db3441c6eace32fb1, {16'd51552, 16'd61949, 16'd60362, 16'd35042, 16'd12675, 16'd48498, 16'd65509, 16'd7145, 16'd19041, 16'd57252, 16'd51024, 16'd64270, 16'd60488, 16'd57235, 16'd27523, 16'd21047, 16'd26196, 16'd9289, 16'd15544, 16'd11757, 16'd56089, 16'd53779, 16'd15556, 16'd23832, 16'd4937, 16'd13240});
	test_expansion(128'h76a1e89cbe17b5879665f75074fc9807, {16'd27729, 16'd35726, 16'd17907, 16'd27228, 16'd43062, 16'd11281, 16'd54799, 16'd10102, 16'd42538, 16'd31917, 16'd37855, 16'd27481, 16'd40563, 16'd34879, 16'd14461, 16'd35132, 16'd7959, 16'd62941, 16'd55614, 16'd45277, 16'd41034, 16'd31687, 16'd19700, 16'd53505, 16'd2933, 16'd4372});
	test_expansion(128'h116806ff6c1de7065490cbe2e7091b49, {16'd2169, 16'd62962, 16'd1704, 16'd46034, 16'd62282, 16'd28048, 16'd20488, 16'd48028, 16'd6687, 16'd24651, 16'd35745, 16'd18567, 16'd62439, 16'd39649, 16'd56125, 16'd25600, 16'd25887, 16'd44474, 16'd13965, 16'd34627, 16'd31710, 16'd59442, 16'd63459, 16'd1894, 16'd39108, 16'd21946});
	test_expansion(128'h73921e3430dff7a1a889d3e24b7f8ba9, {16'd14050, 16'd24976, 16'd55049, 16'd7697, 16'd8654, 16'd41927, 16'd33688, 16'd61235, 16'd49799, 16'd4447, 16'd20392, 16'd33514, 16'd24477, 16'd26675, 16'd27457, 16'd45451, 16'd10413, 16'd20476, 16'd17910, 16'd44689, 16'd36893, 16'd20724, 16'd43788, 16'd30399, 16'd20478, 16'd65423});
	test_expansion(128'h8e49cd1bbf22844ee801758979c1a057, {16'd1040, 16'd25181, 16'd26571, 16'd46454, 16'd31476, 16'd61847, 16'd14962, 16'd16049, 16'd63543, 16'd27943, 16'd25206, 16'd54369, 16'd45211, 16'd4965, 16'd50202, 16'd36995, 16'd64702, 16'd7863, 16'd41785, 16'd32516, 16'd43413, 16'd53440, 16'd11293, 16'd13644, 16'd16899, 16'd31880});
	test_expansion(128'h6aa21548bc1b40275dbd0084e5ddab50, {16'd41637, 16'd32059, 16'd45873, 16'd6539, 16'd19473, 16'd34064, 16'd34564, 16'd13569, 16'd63346, 16'd29384, 16'd30346, 16'd17361, 16'd59935, 16'd39234, 16'd49313, 16'd63644, 16'd55523, 16'd7983, 16'd27579, 16'd39393, 16'd36440, 16'd5754, 16'd56608, 16'd50514, 16'd42297, 16'd8878});
	test_expansion(128'h4f873847b8dc50cb6ade1cf9f18ba813, {16'd25154, 16'd49054, 16'd21743, 16'd30081, 16'd2990, 16'd10624, 16'd59700, 16'd62480, 16'd40543, 16'd10544, 16'd55925, 16'd6588, 16'd16778, 16'd54281, 16'd122, 16'd41736, 16'd16884, 16'd34067, 16'd61318, 16'd20273, 16'd23981, 16'd18976, 16'd50122, 16'd51812, 16'd226, 16'd16224});
	test_expansion(128'h20b142d458f3ac930c40ee3658e89eef, {16'd42964, 16'd8948, 16'd22651, 16'd38406, 16'd8796, 16'd6126, 16'd21171, 16'd64804, 16'd6492, 16'd58016, 16'd43985, 16'd36127, 16'd44358, 16'd19924, 16'd17468, 16'd3179, 16'd38325, 16'd25251, 16'd2947, 16'd10363, 16'd17423, 16'd18641, 16'd46100, 16'd44942, 16'd7613, 16'd39881});
	test_expansion(128'h1901aef1908245588c103176df240c18, {16'd44504, 16'd59814, 16'd49810, 16'd48348, 16'd7466, 16'd30109, 16'd17890, 16'd2320, 16'd29331, 16'd29220, 16'd30976, 16'd62913, 16'd4257, 16'd50702, 16'd43633, 16'd24866, 16'd33293, 16'd5518, 16'd58687, 16'd54704, 16'd25732, 16'd3654, 16'd8498, 16'd44623, 16'd8783, 16'd34870});
	test_expansion(128'hfb31bdc9587185179ef30b629a238eeb, {16'd65077, 16'd3908, 16'd55965, 16'd12902, 16'd37373, 16'd57728, 16'd10198, 16'd45189, 16'd65466, 16'd9741, 16'd42364, 16'd47417, 16'd32722, 16'd484, 16'd26425, 16'd31983, 16'd22869, 16'd28038, 16'd28165, 16'd4354, 16'd64978, 16'd8441, 16'd20508, 16'd34583, 16'd51709, 16'd1858});
	test_expansion(128'h1c573f2f977bbd38af98d45e60af9cbd, {16'd37692, 16'd59900, 16'd35701, 16'd31291, 16'd62447, 16'd59800, 16'd2240, 16'd15799, 16'd22245, 16'd37572, 16'd40787, 16'd49493, 16'd31188, 16'd33333, 16'd28666, 16'd54398, 16'd4749, 16'd28714, 16'd4411, 16'd65403, 16'd7206, 16'd44275, 16'd41722, 16'd4668, 16'd62051, 16'd29826});
	test_expansion(128'hc2e7075af827fab13fc903895726f014, {16'd49668, 16'd15872, 16'd50447, 16'd33474, 16'd26189, 16'd30106, 16'd55838, 16'd19299, 16'd56649, 16'd10062, 16'd38455, 16'd40712, 16'd50176, 16'd58784, 16'd28800, 16'd53509, 16'd31163, 16'd8048, 16'd5365, 16'd26200, 16'd32895, 16'd255, 16'd39772, 16'd1509, 16'd46798, 16'd42079});
	test_expansion(128'hd4a8bba9efad443456f8475e010f2061, {16'd49461, 16'd28297, 16'd28518, 16'd3685, 16'd31924, 16'd6196, 16'd42485, 16'd7242, 16'd63649, 16'd9937, 16'd9459, 16'd18539, 16'd43220, 16'd13204, 16'd27282, 16'd59680, 16'd8244, 16'd59896, 16'd34964, 16'd45296, 16'd32243, 16'd13881, 16'd24310, 16'd33533, 16'd32318, 16'd6076});
	test_expansion(128'he81ced116ac113e1c9ac4698e8e222d7, {16'd63600, 16'd64086, 16'd20341, 16'd52433, 16'd61758, 16'd54101, 16'd63672, 16'd47159, 16'd38098, 16'd58500, 16'd494, 16'd49318, 16'd61549, 16'd59262, 16'd17142, 16'd15192, 16'd60025, 16'd53318, 16'd51509, 16'd45354, 16'd7482, 16'd64717, 16'd15148, 16'd11979, 16'd50542, 16'd7330});
	test_expansion(128'h9b2047cb1d6cf8f08a270e85ee6594b3, {16'd65161, 16'd48758, 16'd11801, 16'd20075, 16'd62317, 16'd47667, 16'd25825, 16'd47035, 16'd5945, 16'd16787, 16'd60343, 16'd15018, 16'd38179, 16'd34059, 16'd11377, 16'd13201, 16'd9664, 16'd5534, 16'd22883, 16'd47114, 16'd21996, 16'd24087, 16'd7615, 16'd10637, 16'd2712, 16'd58655});
	test_expansion(128'h4d41d370026b24cdc6c088701d6c2c88, {16'd28665, 16'd58300, 16'd37874, 16'd64099, 16'd14133, 16'd7129, 16'd30658, 16'd5133, 16'd14803, 16'd42037, 16'd46233, 16'd59984, 16'd17817, 16'd41502, 16'd49657, 16'd8907, 16'd37053, 16'd35599, 16'd63708, 16'd17104, 16'd48910, 16'd48121, 16'd54253, 16'd38642, 16'd47347, 16'd60122});
	test_expansion(128'hc2f6b5afd259f93e1afed58c8bc64d8b, {16'd18610, 16'd50805, 16'd35063, 16'd54705, 16'd23531, 16'd41085, 16'd12245, 16'd55950, 16'd33534, 16'd40510, 16'd22982, 16'd29251, 16'd35523, 16'd34523, 16'd39134, 16'd30021, 16'd5434, 16'd55864, 16'd44099, 16'd48279, 16'd64688, 16'd4982, 16'd61841, 16'd4844, 16'd33021, 16'd38843});
	test_expansion(128'hf3046a5ea6c58bcab1a60127b9aff8f7, {16'd11175, 16'd23366, 16'd6587, 16'd61031, 16'd57524, 16'd24893, 16'd39365, 16'd32141, 16'd21654, 16'd63771, 16'd54082, 16'd37780, 16'd37879, 16'd52373, 16'd41613, 16'd48643, 16'd64708, 16'd14296, 16'd47988, 16'd45901, 16'd48104, 16'd64365, 16'd7031, 16'd10865, 16'd31422, 16'd32543});
	test_expansion(128'h536a5a40af1429959c16bf60f24fb1db, {16'd44448, 16'd47897, 16'd555, 16'd43935, 16'd17231, 16'd9804, 16'd40581, 16'd30232, 16'd57069, 16'd16936, 16'd32155, 16'd39718, 16'd56302, 16'd58394, 16'd18643, 16'd58534, 16'd47141, 16'd49039, 16'd9290, 16'd51131, 16'd2470, 16'd8242, 16'd47002, 16'd8673, 16'd40695, 16'd3686});
	test_expansion(128'hdfa3ec568f5345444362a64d30c66712, {16'd9251, 16'd24887, 16'd17949, 16'd14151, 16'd47961, 16'd29492, 16'd25713, 16'd39134, 16'd57881, 16'd21336, 16'd11838, 16'd47578, 16'd21712, 16'd1154, 16'd6183, 16'd32587, 16'd52055, 16'd396, 16'd7651, 16'd31240, 16'd21501, 16'd47455, 16'd65213, 16'd58051, 16'd37004, 16'd53191});
	test_expansion(128'h77942154444cef929f20512f08ecc50c, {16'd47963, 16'd61555, 16'd30185, 16'd39364, 16'd45123, 16'd34019, 16'd23114, 16'd20781, 16'd57221, 16'd6110, 16'd59367, 16'd62129, 16'd26280, 16'd52540, 16'd24343, 16'd13863, 16'd59329, 16'd25230, 16'd64531, 16'd16772, 16'd44510, 16'd14669, 16'd55212, 16'd37467, 16'd22613, 16'd26262});
	test_expansion(128'h37da5034697a76c3f961b23772252156, {16'd37476, 16'd6407, 16'd33377, 16'd19070, 16'd60733, 16'd20703, 16'd58543, 16'd4775, 16'd49563, 16'd41029, 16'd37066, 16'd49531, 16'd53669, 16'd17024, 16'd34122, 16'd40582, 16'd15386, 16'd5378, 16'd2978, 16'd21044, 16'd53374, 16'd1551, 16'd14894, 16'd26891, 16'd45259, 16'd467});
	test_expansion(128'h0dee744e3cb30397b03eb9a9dcdf5fea, {16'd28767, 16'd1620, 16'd47415, 16'd65187, 16'd33682, 16'd38479, 16'd30282, 16'd29873, 16'd8457, 16'd8414, 16'd21875, 16'd479, 16'd14690, 16'd59857, 16'd63033, 16'd16183, 16'd9952, 16'd31257, 16'd30702, 16'd61010, 16'd43297, 16'd37371, 16'd37948, 16'd8028, 16'd39660, 16'd16427});
	test_expansion(128'h92f85819b86f1430b3776458a469065d, {16'd36526, 16'd57399, 16'd6668, 16'd60038, 16'd38021, 16'd56882, 16'd46690, 16'd64798, 16'd28004, 16'd14474, 16'd47307, 16'd43328, 16'd35803, 16'd38096, 16'd53112, 16'd59922, 16'd34383, 16'd39955, 16'd23166, 16'd57614, 16'd7062, 16'd8829, 16'd12622, 16'd48630, 16'd4393, 16'd4070});
	test_expansion(128'h9fb1ad08babf1af6bf9796cdac29031a, {16'd18588, 16'd4109, 16'd42685, 16'd51230, 16'd24139, 16'd29782, 16'd215, 16'd5621, 16'd17702, 16'd63551, 16'd39004, 16'd64026, 16'd37158, 16'd45803, 16'd60874, 16'd47196, 16'd28584, 16'd9567, 16'd11532, 16'd61146, 16'd16146, 16'd25633, 16'd48891, 16'd22849, 16'd48571, 16'd12693});
	test_expansion(128'h9fe400a7876b2e524c5f4610e99afce5, {16'd29514, 16'd63670, 16'd15663, 16'd23021, 16'd34661, 16'd18645, 16'd1848, 16'd7025, 16'd33497, 16'd36752, 16'd10540, 16'd37258, 16'd1722, 16'd13884, 16'd58765, 16'd17234, 16'd39441, 16'd9040, 16'd54369, 16'd17880, 16'd10007, 16'd12548, 16'd39828, 16'd37184, 16'd55833, 16'd53337});
	test_expansion(128'hce379f0caaa5807fcd5c5a819a8fd756, {16'd11356, 16'd17262, 16'd45701, 16'd24460, 16'd52096, 16'd59189, 16'd45732, 16'd4510, 16'd31504, 16'd4711, 16'd31878, 16'd49365, 16'd32149, 16'd57763, 16'd47512, 16'd531, 16'd29554, 16'd21618, 16'd20700, 16'd62066, 16'd13171, 16'd58778, 16'd12651, 16'd52161, 16'd61281, 16'd44106});
	test_expansion(128'h17199c49e37d1e38b888bc6129d2223a, {16'd36101, 16'd27590, 16'd48333, 16'd33861, 16'd42583, 16'd24676, 16'd24000, 16'd21920, 16'd15792, 16'd38034, 16'd52410, 16'd3794, 16'd53646, 16'd28273, 16'd2029, 16'd43314, 16'd46898, 16'd3853, 16'd34134, 16'd1972, 16'd28191, 16'd63266, 16'd688, 16'd49618, 16'd22182, 16'd33108});
	test_expansion(128'hc89eddd83e21754206eb3917e653e78c, {16'd57510, 16'd10009, 16'd52697, 16'd43203, 16'd1930, 16'd40504, 16'd61217, 16'd61889, 16'd58867, 16'd35687, 16'd35571, 16'd26928, 16'd2848, 16'd25867, 16'd28660, 16'd45987, 16'd36665, 16'd55033, 16'd30251, 16'd57012, 16'd27765, 16'd22301, 16'd10827, 16'd32379, 16'd2190, 16'd26408});
	test_expansion(128'h00e2e76a9e79daa7b45511a1e711c466, {16'd60936, 16'd44972, 16'd57116, 16'd26279, 16'd49074, 16'd39374, 16'd21933, 16'd21077, 16'd54198, 16'd14726, 16'd3538, 16'd24120, 16'd36632, 16'd13655, 16'd3494, 16'd50942, 16'd8958, 16'd20400, 16'd55781, 16'd43627, 16'd29232, 16'd62849, 16'd12706, 16'd2518, 16'd49959, 16'd25471});
	test_expansion(128'h98ef27435762f63cf887a15f68d1538d, {16'd18618, 16'd15547, 16'd10198, 16'd6651, 16'd53431, 16'd27771, 16'd59533, 16'd24469, 16'd46779, 16'd73, 16'd32949, 16'd13279, 16'd33073, 16'd63184, 16'd41306, 16'd6719, 16'd6515, 16'd35735, 16'd39693, 16'd16093, 16'd36028, 16'd42305, 16'd47734, 16'd27099, 16'd19688, 16'd54078});
	test_expansion(128'h8dcdf3ce0d7952332519aa9b3ed52513, {16'd15668, 16'd20881, 16'd7137, 16'd40421, 16'd62711, 16'd54205, 16'd41070, 16'd38842, 16'd20367, 16'd33788, 16'd39350, 16'd33263, 16'd23153, 16'd41620, 16'd31823, 16'd49992, 16'd38786, 16'd16772, 16'd59614, 16'd3720, 16'd15152, 16'd5556, 16'd55293, 16'd54323, 16'd58912, 16'd47851});
	test_expansion(128'h101af1b2c54179dcf46b1208db36463d, {16'd61261, 16'd31433, 16'd30292, 16'd52243, 16'd1547, 16'd57304, 16'd53338, 16'd31895, 16'd8567, 16'd49445, 16'd25602, 16'd57863, 16'd56490, 16'd31755, 16'd42805, 16'd38776, 16'd40799, 16'd39643, 16'd27929, 16'd17866, 16'd20305, 16'd63408, 16'd4469, 16'd22103, 16'd59129, 16'd17259});
	test_expansion(128'h1ed6d2cdedea2f9f037ee8c5a84061a8, {16'd21299, 16'd39762, 16'd59896, 16'd42820, 16'd38909, 16'd28556, 16'd18235, 16'd38408, 16'd4361, 16'd63494, 16'd26867, 16'd3050, 16'd11838, 16'd51262, 16'd25259, 16'd54242, 16'd19571, 16'd59635, 16'd26709, 16'd17103, 16'd23955, 16'd29999, 16'd1306, 16'd31219, 16'd40979, 16'd51206});
	test_expansion(128'h3bba88dd83d546073dfb2523bf875dcb, {16'd19807, 16'd41517, 16'd36143, 16'd32456, 16'd47225, 16'd25040, 16'd56273, 16'd16620, 16'd28784, 16'd61600, 16'd23233, 16'd44023, 16'd20323, 16'd9381, 16'd36007, 16'd10350, 16'd51348, 16'd45478, 16'd21451, 16'd11090, 16'd62745, 16'd59117, 16'd1914, 16'd33685, 16'd57294, 16'd39235});
	test_expansion(128'hc85d8d58b3c3875fbd51be28b51ed401, {16'd60860, 16'd13720, 16'd41656, 16'd26900, 16'd39329, 16'd56840, 16'd61136, 16'd8718, 16'd38170, 16'd37431, 16'd5989, 16'd63372, 16'd16866, 16'd50033, 16'd5245, 16'd34991, 16'd30485, 16'd20526, 16'd18501, 16'd14807, 16'd60842, 16'd45046, 16'd11607, 16'd23454, 16'd23701, 16'd45807});
	test_expansion(128'h99892c7c5868415e1bf73340dd50c7d7, {16'd58187, 16'd32080, 16'd20594, 16'd53593, 16'd8793, 16'd59900, 16'd29338, 16'd15188, 16'd4236, 16'd12078, 16'd46354, 16'd64854, 16'd52372, 16'd58265, 16'd12600, 16'd44193, 16'd65429, 16'd53550, 16'd35902, 16'd31472, 16'd65047, 16'd15491, 16'd9327, 16'd29407, 16'd52863, 16'd4310});
	test_expansion(128'h9623de7705aed5454bc89f5c784b27f1, {16'd22945, 16'd18124, 16'd42381, 16'd27660, 16'd1104, 16'd30798, 16'd845, 16'd42412, 16'd1956, 16'd63331, 16'd46723, 16'd60563, 16'd1226, 16'd56671, 16'd40474, 16'd46883, 16'd33699, 16'd37349, 16'd48323, 16'd39794, 16'd63401, 16'd210, 16'd3149, 16'd58132, 16'd46156, 16'd53015});
	test_expansion(128'h8195a4838543373a23e40ac207ea4445, {16'd25295, 16'd15053, 16'd8178, 16'd47326, 16'd37888, 16'd52414, 16'd26001, 16'd35960, 16'd36375, 16'd36485, 16'd37333, 16'd48369, 16'd31629, 16'd35973, 16'd27741, 16'd22941, 16'd42640, 16'd55144, 16'd32439, 16'd25468, 16'd23454, 16'd43590, 16'd26960, 16'd22202, 16'd33667, 16'd26056});
	test_expansion(128'hee269b2f10ebb275da2cf51fc82cfe52, {16'd63923, 16'd39155, 16'd12650, 16'd4994, 16'd64390, 16'd52690, 16'd8621, 16'd36155, 16'd6783, 16'd52335, 16'd64156, 16'd49226, 16'd60551, 16'd57554, 16'd49512, 16'd38383, 16'd19117, 16'd24499, 16'd45982, 16'd3035, 16'd36416, 16'd3700, 16'd26834, 16'd30739, 16'd52842, 16'd30214});
	test_expansion(128'h2250f77b84d5c51146471c394d3c28a5, {16'd38903, 16'd9927, 16'd32573, 16'd26360, 16'd59525, 16'd15179, 16'd32624, 16'd10560, 16'd37127, 16'd63079, 16'd40538, 16'd37592, 16'd25280, 16'd17253, 16'd34129, 16'd1605, 16'd40686, 16'd20884, 16'd61545, 16'd26674, 16'd23716, 16'd61910, 16'd42957, 16'd47219, 16'd49853, 16'd33346});
	test_expansion(128'h889570252654f1218aa392584779e5f6, {16'd12645, 16'd40963, 16'd15182, 16'd16687, 16'd63498, 16'd50149, 16'd28648, 16'd64840, 16'd15198, 16'd63851, 16'd18022, 16'd41797, 16'd35492, 16'd8520, 16'd41682, 16'd32791, 16'd15667, 16'd30650, 16'd761, 16'd5417, 16'd35034, 16'd53489, 16'd15950, 16'd10492, 16'd60529, 16'd53746});
	test_expansion(128'hefdd377096aef7ff3b87630212f6bf19, {16'd61657, 16'd50682, 16'd18109, 16'd62177, 16'd52066, 16'd60786, 16'd26639, 16'd14776, 16'd6991, 16'd33915, 16'd47005, 16'd27792, 16'd37410, 16'd38760, 16'd6846, 16'd9459, 16'd40616, 16'd13714, 16'd61565, 16'd55278, 16'd39346, 16'd53668, 16'd29284, 16'd35809, 16'd54569, 16'd1749});
	test_expansion(128'h14417fe8f70c9c4ba37b8844d9f20f53, {16'd20906, 16'd15729, 16'd5795, 16'd61146, 16'd22324, 16'd41344, 16'd63455, 16'd58629, 16'd7207, 16'd3915, 16'd41191, 16'd57331, 16'd3628, 16'd1755, 16'd5490, 16'd10512, 16'd64856, 16'd13734, 16'd58973, 16'd63277, 16'd26452, 16'd64200, 16'd21664, 16'd34506, 16'd36698, 16'd33823});
	test_expansion(128'h606478601ab641d704fd44c7874bbf30, {16'd48762, 16'd783, 16'd313, 16'd11176, 16'd40909, 16'd37715, 16'd30222, 16'd59252, 16'd61046, 16'd32483, 16'd16818, 16'd48549, 16'd27773, 16'd61587, 16'd31760, 16'd48279, 16'd36859, 16'd8723, 16'd62274, 16'd34670, 16'd61142, 16'd39633, 16'd34024, 16'd44771, 16'd21603, 16'd6159});
	test_expansion(128'h42694aaf8eb3e5f24d679842e65cba74, {16'd36583, 16'd27030, 16'd59799, 16'd34481, 16'd53835, 16'd24724, 16'd34971, 16'd50133, 16'd23546, 16'd30063, 16'd62358, 16'd18318, 16'd4825, 16'd42232, 16'd40861, 16'd7057, 16'd56718, 16'd14458, 16'd14368, 16'd39754, 16'd44654, 16'd20176, 16'd5266, 16'd32569, 16'd7233, 16'd16088});
	test_expansion(128'h078862a3956b90470e0c6bd9963677c2, {16'd16077, 16'd36913, 16'd54976, 16'd5146, 16'd53196, 16'd17652, 16'd10083, 16'd62285, 16'd33243, 16'd52741, 16'd41679, 16'd53438, 16'd56307, 16'd8517, 16'd50398, 16'd30165, 16'd6937, 16'd29473, 16'd34658, 16'd55018, 16'd35923, 16'd26378, 16'd1976, 16'd28416, 16'd41481, 16'd33260});
	test_expansion(128'he392b0440903b4ef2e46ac5524afaa9d, {16'd26352, 16'd19711, 16'd51731, 16'd48213, 16'd45312, 16'd15920, 16'd39838, 16'd40413, 16'd7463, 16'd50909, 16'd1892, 16'd8431, 16'd48424, 16'd59272, 16'd43495, 16'd10796, 16'd50184, 16'd5295, 16'd5943, 16'd26002, 16'd29638, 16'd15296, 16'd33705, 16'd11606, 16'd58970, 16'd19086});
	test_expansion(128'h54c764bd7c115d3317a92b3a4b4dceae, {16'd44869, 16'd47825, 16'd7550, 16'd36907, 16'd10632, 16'd5281, 16'd46594, 16'd23968, 16'd55159, 16'd35324, 16'd62109, 16'd11381, 16'd54105, 16'd38802, 16'd25678, 16'd1680, 16'd16564, 16'd11423, 16'd9770, 16'd40417, 16'd34433, 16'd63946, 16'd51811, 16'd35749, 16'd57114, 16'd59388});
	test_expansion(128'h312597be2a989db6cfc516149caf1c34, {16'd36199, 16'd40536, 16'd21453, 16'd14558, 16'd17991, 16'd43065, 16'd2442, 16'd20806, 16'd9706, 16'd9362, 16'd20274, 16'd57016, 16'd56028, 16'd58396, 16'd8712, 16'd8711, 16'd50314, 16'd49922, 16'd29175, 16'd18852, 16'd6991, 16'd39718, 16'd5063, 16'd10426, 16'd47983, 16'd46172});
	test_expansion(128'h40d125e46db1c62c7c91891aa97d2a9b, {16'd1842, 16'd41527, 16'd40519, 16'd19286, 16'd20122, 16'd53886, 16'd55135, 16'd44475, 16'd35645, 16'd18944, 16'd16681, 16'd62542, 16'd64297, 16'd55603, 16'd35728, 16'd64909, 16'd35280, 16'd20646, 16'd51815, 16'd29595, 16'd6386, 16'd17250, 16'd55058, 16'd15762, 16'd59368, 16'd28361});
	test_expansion(128'hddd1bfc03bf353731895ce15d7a2a7e6, {16'd15489, 16'd51480, 16'd31594, 16'd29324, 16'd62668, 16'd13934, 16'd58260, 16'd52007, 16'd63447, 16'd13463, 16'd52905, 16'd19692, 16'd24298, 16'd42259, 16'd50353, 16'd35951, 16'd2295, 16'd2461, 16'd11185, 16'd6210, 16'd45360, 16'd38052, 16'd58543, 16'd59441, 16'd50598, 16'd48706});
	test_expansion(128'h3dc3ed9be4956e26bb2c6a885b9527b9, {16'd50961, 16'd52622, 16'd31952, 16'd32259, 16'd4057, 16'd47677, 16'd55926, 16'd16069, 16'd23605, 16'd5137, 16'd30932, 16'd28274, 16'd64548, 16'd44770, 16'd6571, 16'd59466, 16'd64916, 16'd33958, 16'd58442, 16'd31325, 16'd49659, 16'd62153, 16'd16355, 16'd58761, 16'd1567, 16'd42854});
	test_expansion(128'h63dc9c25b21a1b921f393626b5f75abc, {16'd51198, 16'd4581, 16'd27955, 16'd55548, 16'd452, 16'd49764, 16'd15034, 16'd39822, 16'd18766, 16'd14896, 16'd7802, 16'd36659, 16'd31951, 16'd61058, 16'd47967, 16'd51072, 16'd31870, 16'd48907, 16'd50775, 16'd18454, 16'd61323, 16'd44528, 16'd31853, 16'd18184, 16'd19665, 16'd28815});
	test_expansion(128'h0041553315bb93105e8e615a2c0a4530, {16'd56492, 16'd45004, 16'd29904, 16'd5231, 16'd39753, 16'd7136, 16'd22295, 16'd63398, 16'd31816, 16'd5140, 16'd20781, 16'd43946, 16'd14865, 16'd18256, 16'd5831, 16'd43649, 16'd13318, 16'd37133, 16'd38980, 16'd39505, 16'd33100, 16'd51435, 16'd36018, 16'd6227, 16'd56249, 16'd22128});
	test_expansion(128'h69caaa0d3835d0168da0f4d5ffe01f61, {16'd32253, 16'd11152, 16'd55529, 16'd4594, 16'd8397, 16'd25695, 16'd11344, 16'd55041, 16'd43546, 16'd35882, 16'd54698, 16'd346, 16'd42427, 16'd3970, 16'd63263, 16'd49112, 16'd11593, 16'd25520, 16'd57306, 16'd22595, 16'd18411, 16'd43836, 16'd51014, 16'd21114, 16'd23037, 16'd45030});
	test_expansion(128'h99edbe20b8b78d10e682ad186d1935e6, {16'd55910, 16'd55374, 16'd45180, 16'd57501, 16'd29883, 16'd54211, 16'd6451, 16'd11920, 16'd32259, 16'd54586, 16'd52479, 16'd11833, 16'd10749, 16'd33893, 16'd32043, 16'd47319, 16'd35467, 16'd51177, 16'd23650, 16'd11525, 16'd60815, 16'd3366, 16'd47864, 16'd7861, 16'd63752, 16'd17768});
	test_expansion(128'h8adf79ec5f5e3e21467a6ab054b3f3f9, {16'd50823, 16'd43319, 16'd29115, 16'd18002, 16'd36580, 16'd26270, 16'd26940, 16'd20794, 16'd37218, 16'd54101, 16'd5065, 16'd47985, 16'd26629, 16'd17263, 16'd19042, 16'd11622, 16'd58899, 16'd29169, 16'd52773, 16'd50760, 16'd44982, 16'd23942, 16'd26052, 16'd37651, 16'd30862, 16'd20396});
	test_expansion(128'h87d0f82a972028e115c27094058a4e55, {16'd41893, 16'd49487, 16'd30568, 16'd29761, 16'd33502, 16'd25916, 16'd25618, 16'd64120, 16'd62731, 16'd15387, 16'd38028, 16'd47646, 16'd18470, 16'd30908, 16'd25094, 16'd46272, 16'd34342, 16'd42820, 16'd35623, 16'd5338, 16'd19185, 16'd62956, 16'd13188, 16'd36956, 16'd35914, 16'd61104});
	test_expansion(128'h32305aebc367a42cdb502fb68c11add6, {16'd33596, 16'd28569, 16'd30064, 16'd60627, 16'd9169, 16'd1755, 16'd10210, 16'd33518, 16'd57805, 16'd54010, 16'd43318, 16'd27209, 16'd48239, 16'd19567, 16'd58838, 16'd14392, 16'd4855, 16'd47600, 16'd15763, 16'd11521, 16'd18090, 16'd36106, 16'd48421, 16'd32551, 16'd608, 16'd48782});
	test_expansion(128'hedb73df40362de4d09220eb32b6a2c3d, {16'd62461, 16'd8277, 16'd31008, 16'd32021, 16'd63299, 16'd21019, 16'd52748, 16'd42792, 16'd30840, 16'd54215, 16'd33369, 16'd42742, 16'd60134, 16'd25537, 16'd6936, 16'd5711, 16'd2696, 16'd2548, 16'd55825, 16'd19547, 16'd9520, 16'd19595, 16'd8725, 16'd198, 16'd65475, 16'd22065});
	test_expansion(128'h400f18bc1e63e46c62b774c71753d018, {16'd13248, 16'd30702, 16'd27713, 16'd28979, 16'd61704, 16'd55939, 16'd19745, 16'd18541, 16'd43604, 16'd22242, 16'd43603, 16'd30561, 16'd12843, 16'd40246, 16'd65383, 16'd23760, 16'd39563, 16'd28840, 16'd48898, 16'd29823, 16'd23416, 16'd49664, 16'd61500, 16'd30878, 16'd20565, 16'd18755});
	test_expansion(128'h6f628a8ffc8872fbd4b9761edca9e9ce, {16'd38016, 16'd64186, 16'd59829, 16'd16215, 16'd39867, 16'd2916, 16'd20715, 16'd22103, 16'd48810, 16'd31425, 16'd31491, 16'd33712, 16'd21130, 16'd10565, 16'd46139, 16'd13879, 16'd59687, 16'd44108, 16'd30, 16'd18166, 16'd7698, 16'd5493, 16'd7734, 16'd41395, 16'd25644, 16'd49192});
	test_expansion(128'h2ae8e8028f9f1e3f1044062a24913b74, {16'd44694, 16'd18511, 16'd29995, 16'd5633, 16'd19209, 16'd39156, 16'd43183, 16'd31606, 16'd24939, 16'd49834, 16'd61212, 16'd50263, 16'd39604, 16'd12705, 16'd56646, 16'd57924, 16'd12544, 16'd65348, 16'd64952, 16'd44204, 16'd26881, 16'd21276, 16'd51213, 16'd3109, 16'd55267, 16'd27551});
	test_expansion(128'h9323414d5bc1c94e542d95104f2a809f, {16'd61061, 16'd45257, 16'd13116, 16'd63860, 16'd42211, 16'd8679, 16'd55550, 16'd13383, 16'd11088, 16'd58074, 16'd6891, 16'd42699, 16'd65067, 16'd54511, 16'd26716, 16'd58596, 16'd63225, 16'd23986, 16'd40041, 16'd27763, 16'd9208, 16'd6052, 16'd1882, 16'd48970, 16'd9167, 16'd33015});
	test_expansion(128'h312231d2416af6e12942536f2704a96b, {16'd10832, 16'd25488, 16'd33612, 16'd2337, 16'd53758, 16'd3557, 16'd16394, 16'd22464, 16'd9254, 16'd43224, 16'd40820, 16'd13688, 16'd20240, 16'd45584, 16'd50594, 16'd19040, 16'd58599, 16'd17109, 16'd31078, 16'd17766, 16'd61791, 16'd21856, 16'd42034, 16'd2257, 16'd7048, 16'd31074});
	test_expansion(128'h0f8b32cfffdcdaac69b42a7747f2ffc8, {16'd48995, 16'd20058, 16'd16475, 16'd45022, 16'd22884, 16'd36235, 16'd12462, 16'd15217, 16'd33452, 16'd53719, 16'd53296, 16'd43815, 16'd13185, 16'd33122, 16'd52045, 16'd62744, 16'd2420, 16'd34378, 16'd36896, 16'd52736, 16'd33071, 16'd46062, 16'd22914, 16'd26428, 16'd10010, 16'd2683});
	test_expansion(128'h33476136b80cb0f23ed163a01c86caae, {16'd17566, 16'd1394, 16'd45816, 16'd32933, 16'd47972, 16'd5173, 16'd65512, 16'd51223, 16'd45529, 16'd42050, 16'd56870, 16'd3305, 16'd36536, 16'd36978, 16'd6855, 16'd58351, 16'd6596, 16'd65208, 16'd52678, 16'd54307, 16'd64722, 16'd27806, 16'd5430, 16'd49788, 16'd30206, 16'd10836});
	test_expansion(128'h93ac04f2f31eef25933584ee01016eca, {16'd47382, 16'd20889, 16'd44420, 16'd13579, 16'd57347, 16'd20263, 16'd38616, 16'd42179, 16'd63784, 16'd1400, 16'd19316, 16'd27651, 16'd43324, 16'd7213, 16'd45324, 16'd52028, 16'd19378, 16'd18924, 16'd3941, 16'd62582, 16'd37906, 16'd56963, 16'd63890, 16'd101, 16'd59219, 16'd64231});
	test_expansion(128'ha4b092d3467712ce4387989a3595f330, {16'd7201, 16'd43065, 16'd65402, 16'd44598, 16'd16975, 16'd8315, 16'd28811, 16'd47602, 16'd63932, 16'd55623, 16'd35539, 16'd47846, 16'd61082, 16'd44911, 16'd25513, 16'd41254, 16'd61973, 16'd18778, 16'd44640, 16'd57210, 16'd10898, 16'd1732, 16'd60415, 16'd39071, 16'd58800, 16'd7784});
	test_expansion(128'h59e597210ab1ac70924ea7308976d6d0, {16'd55719, 16'd23866, 16'd65384, 16'd28162, 16'd63588, 16'd62697, 16'd20791, 16'd44746, 16'd48952, 16'd14782, 16'd16528, 16'd8538, 16'd54, 16'd98, 16'd52878, 16'd13936, 16'd31022, 16'd43079, 16'd28043, 16'd58781, 16'd16060, 16'd6579, 16'd32103, 16'd63381, 16'd16771, 16'd54515});
	test_expansion(128'h994922c5a16b3ca0bb950a71048849a4, {16'd44884, 16'd30224, 16'd48469, 16'd65088, 16'd20990, 16'd20702, 16'd14378, 16'd2758, 16'd45566, 16'd65106, 16'd59046, 16'd36289, 16'd3477, 16'd10825, 16'd44217, 16'd38263, 16'd50565, 16'd5524, 16'd51341, 16'd20440, 16'd35353, 16'd52075, 16'd17531, 16'd18671, 16'd46838, 16'd17455});
	test_expansion(128'h1311aff855ca12762c34e6895b8cfedc, {16'd23973, 16'd39580, 16'd61032, 16'd31377, 16'd52007, 16'd46992, 16'd46534, 16'd26911, 16'd24556, 16'd65068, 16'd56107, 16'd44255, 16'd59949, 16'd35075, 16'd49202, 16'd48432, 16'd10868, 16'd61221, 16'd7235, 16'd9901, 16'd10677, 16'd52365, 16'd31291, 16'd11887, 16'd21996, 16'd62778});
	test_expansion(128'hc32f1161944f986a7423c75c5e9afd97, {16'd39634, 16'd52075, 16'd31895, 16'd38398, 16'd7726, 16'd55056, 16'd21683, 16'd55123, 16'd57325, 16'd34254, 16'd61982, 16'd836, 16'd54097, 16'd31316, 16'd24772, 16'd29189, 16'd50787, 16'd9669, 16'd58650, 16'd1648, 16'd52875, 16'd26996, 16'd25985, 16'd43926, 16'd43662, 16'd65104});
	test_expansion(128'hd5879de63540b0b1a57ac11249385cf1, {16'd18420, 16'd17624, 16'd56141, 16'd24495, 16'd13370, 16'd29003, 16'd50284, 16'd8955, 16'd1520, 16'd10152, 16'd12387, 16'd11235, 16'd60548, 16'd47531, 16'd41789, 16'd25265, 16'd7569, 16'd6574, 16'd40620, 16'd57400, 16'd11430, 16'd21597, 16'd9594, 16'd38387, 16'd17568, 16'd12200});
	test_expansion(128'h7c128f3eef58480329c14c0a8ac15783, {16'd44215, 16'd14216, 16'd4556, 16'd36710, 16'd61533, 16'd38379, 16'd17997, 16'd11086, 16'd33847, 16'd5820, 16'd61383, 16'd44630, 16'd64417, 16'd62856, 16'd32100, 16'd45960, 16'd59634, 16'd17145, 16'd53842, 16'd16230, 16'd8983, 16'd8682, 16'd62605, 16'd11447, 16'd54051, 16'd13776});
	test_expansion(128'hf999f58c4bb17097cf139c7fe9f27711, {16'd48876, 16'd29294, 16'd46923, 16'd44429, 16'd53161, 16'd22820, 16'd35853, 16'd61595, 16'd25420, 16'd37259, 16'd17062, 16'd7162, 16'd49417, 16'd19166, 16'd40507, 16'd2261, 16'd44250, 16'd20558, 16'd59860, 16'd51921, 16'd27844, 16'd2431, 16'd21078, 16'd44629, 16'd58120, 16'd56713});
	test_expansion(128'hdf6e2c9689d83574374b78bf70657bef, {16'd38319, 16'd57033, 16'd60775, 16'd44952, 16'd36314, 16'd18621, 16'd57493, 16'd40527, 16'd45659, 16'd16749, 16'd27863, 16'd4278, 16'd38619, 16'd4040, 16'd19414, 16'd51488, 16'd15743, 16'd11763, 16'd64474, 16'd63639, 16'd21422, 16'd18987, 16'd47587, 16'd34927, 16'd52362, 16'd42766});
	test_expansion(128'h4b5895641467905c33fa655e833c88ad, {16'd56717, 16'd22928, 16'd27171, 16'd31798, 16'd1079, 16'd46972, 16'd48268, 16'd1867, 16'd14393, 16'd9331, 16'd25305, 16'd55297, 16'd45064, 16'd38428, 16'd49215, 16'd20866, 16'd33001, 16'd31948, 16'd54115, 16'd19314, 16'd33556, 16'd64356, 16'd38461, 16'd12304, 16'd23352, 16'd34525});
	test_expansion(128'h7d364b4ba52fce10340b0fd30f51785e, {16'd28529, 16'd3665, 16'd28514, 16'd38790, 16'd63928, 16'd11733, 16'd30436, 16'd15373, 16'd24365, 16'd26616, 16'd44831, 16'd46563, 16'd36832, 16'd12045, 16'd51666, 16'd57209, 16'd1131, 16'd27276, 16'd63329, 16'd37795, 16'd21540, 16'd13234, 16'd20314, 16'd49138, 16'd25177, 16'd13285});
	test_expansion(128'h9002473c081c0228b8fa60e09a132dc3, {16'd61887, 16'd49185, 16'd18585, 16'd7041, 16'd26230, 16'd46331, 16'd36280, 16'd4318, 16'd11703, 16'd13216, 16'd46515, 16'd34833, 16'd1425, 16'd8273, 16'd19565, 16'd33301, 16'd47641, 16'd46225, 16'd65502, 16'd17688, 16'd5717, 16'd62404, 16'd31495, 16'd29887, 16'd3590, 16'd9025});
	test_expansion(128'h3dd300c46d54ccd2ae57e22a21e1640c, {16'd55725, 16'd15422, 16'd11666, 16'd22956, 16'd22509, 16'd54666, 16'd45682, 16'd52191, 16'd61093, 16'd8733, 16'd30349, 16'd24496, 16'd30348, 16'd28510, 16'd40468, 16'd56714, 16'd24197, 16'd51118, 16'd55677, 16'd14591, 16'd44348, 16'd16309, 16'd899, 16'd26986, 16'd52735, 16'd4916});
	test_expansion(128'h73dd0f94ea323e8f8e64e06d1396fc02, {16'd4203, 16'd4627, 16'd37890, 16'd37302, 16'd65253, 16'd25184, 16'd28454, 16'd29858, 16'd57793, 16'd47902, 16'd46728, 16'd65347, 16'd48580, 16'd32995, 16'd12464, 16'd9919, 16'd22138, 16'd38037, 16'd1109, 16'd8154, 16'd25981, 16'd52764, 16'd31514, 16'd53595, 16'd48100, 16'd29105});
	test_expansion(128'h49e3a262f6541bfae9d918f1653126e0, {16'd22820, 16'd36071, 16'd49139, 16'd7701, 16'd39921, 16'd58573, 16'd27727, 16'd63435, 16'd8469, 16'd18884, 16'd10448, 16'd10477, 16'd20597, 16'd21135, 16'd45290, 16'd10980, 16'd50731, 16'd61158, 16'd22622, 16'd40010, 16'd5718, 16'd3148, 16'd35360, 16'd17108, 16'd64091, 16'd54405});
	test_expansion(128'h9901d2f7a27712bf3644a5dab6afb9d1, {16'd49343, 16'd47041, 16'd36209, 16'd55241, 16'd43062, 16'd4190, 16'd26635, 16'd36257, 16'd2900, 16'd31123, 16'd10173, 16'd12156, 16'd48188, 16'd6752, 16'd46772, 16'd28970, 16'd28571, 16'd41092, 16'd24571, 16'd19322, 16'd40804, 16'd54883, 16'd22975, 16'd1386, 16'd6155, 16'd1090});
	test_expansion(128'ha1a6ad490cb88f9bde5d2f056b99ff33, {16'd41455, 16'd20398, 16'd61473, 16'd61182, 16'd17536, 16'd6141, 16'd12654, 16'd3143, 16'd56468, 16'd26191, 16'd41554, 16'd27853, 16'd1182, 16'd29235, 16'd49893, 16'd18735, 16'd21250, 16'd10999, 16'd49925, 16'd62756, 16'd51584, 16'd64306, 16'd22870, 16'd37914, 16'd46312, 16'd8179});
	test_expansion(128'hd2eb1f95384150ddb1f206aa268253ca, {16'd18743, 16'd37741, 16'd14550, 16'd54031, 16'd34274, 16'd49503, 16'd61636, 16'd47601, 16'd16295, 16'd14709, 16'd20337, 16'd1732, 16'd22131, 16'd3502, 16'd22088, 16'd56964, 16'd39550, 16'd48846, 16'd65395, 16'd28903, 16'd59212, 16'd4503, 16'd13413, 16'd12709, 16'd36975, 16'd65443});
	test_expansion(128'hb01079e02e4de68de820c4e80559e17e, {16'd22573, 16'd61778, 16'd20271, 16'd7742, 16'd40671, 16'd25661, 16'd59365, 16'd52553, 16'd27428, 16'd22280, 16'd56067, 16'd7011, 16'd28121, 16'd12590, 16'd45529, 16'd50544, 16'd1286, 16'd26757, 16'd42193, 16'd49665, 16'd1829, 16'd37539, 16'd11727, 16'd52581, 16'd27682, 16'd25880});
	test_expansion(128'hc56d15268358ec5adfa4b61a9871a74c, {16'd20452, 16'd57148, 16'd52054, 16'd13532, 16'd12455, 16'd64178, 16'd6578, 16'd2811, 16'd62791, 16'd29542, 16'd45950, 16'd51203, 16'd44524, 16'd21085, 16'd35465, 16'd60313, 16'd29223, 16'd58075, 16'd38728, 16'd55678, 16'd27957, 16'd37263, 16'd35327, 16'd43761, 16'd17355, 16'd9357});
	test_expansion(128'h4c21a324bafef5140e7bb5ed0161fd0c, {16'd54161, 16'd51456, 16'd14687, 16'd9417, 16'd53691, 16'd43510, 16'd30121, 16'd1683, 16'd13311, 16'd42912, 16'd41079, 16'd24741, 16'd18825, 16'd2922, 16'd19592, 16'd44731, 16'd7827, 16'd50947, 16'd17197, 16'd25794, 16'd27061, 16'd56929, 16'd36980, 16'd21862, 16'd46378, 16'd25322});
	test_expansion(128'hf37aef451fb1ef90ce8a8f6e6e825b41, {16'd46229, 16'd8615, 16'd23577, 16'd5003, 16'd46257, 16'd8139, 16'd266, 16'd21370, 16'd4786, 16'd20893, 16'd34446, 16'd38047, 16'd35185, 16'd55501, 16'd19898, 16'd65398, 16'd43637, 16'd61504, 16'd61122, 16'd2331, 16'd35613, 16'd44827, 16'd11690, 16'd8957, 16'd18591, 16'd29963});
	test_expansion(128'h8f2e814f2a5b0347b2adc24295af1ae0, {16'd49368, 16'd54377, 16'd5448, 16'd11715, 16'd65044, 16'd46313, 16'd23636, 16'd2737, 16'd20107, 16'd57084, 16'd1500, 16'd10482, 16'd52108, 16'd42470, 16'd35716, 16'd58279, 16'd38381, 16'd18125, 16'd14192, 16'd41231, 16'd31829, 16'd47163, 16'd10450, 16'd34088, 16'd42259, 16'd34312});
	test_expansion(128'hea28409cd54709a39e63bc96db62d37d, {16'd5530, 16'd60819, 16'd30763, 16'd7768, 16'd48528, 16'd13180, 16'd36050, 16'd31625, 16'd11170, 16'd51403, 16'd31412, 16'd40090, 16'd6626, 16'd40570, 16'd30272, 16'd57198, 16'd19847, 16'd53704, 16'd58904, 16'd64785, 16'd45229, 16'd8559, 16'd17989, 16'd60217, 16'd27017, 16'd41716});
	test_expansion(128'hc4857964d7864bb23a0ab7546ce6208b, {16'd39994, 16'd33703, 16'd30252, 16'd6824, 16'd63134, 16'd49464, 16'd39534, 16'd64532, 16'd52075, 16'd34479, 16'd64580, 16'd22373, 16'd2932, 16'd856, 16'd6415, 16'd27552, 16'd12679, 16'd35963, 16'd35647, 16'd61895, 16'd6798, 16'd37390, 16'd31688, 16'd35233, 16'd13612, 16'd30600});
	test_expansion(128'h5fcec5e5af53620d80f691e5ad16208a, {16'd33498, 16'd34932, 16'd31453, 16'd2860, 16'd17251, 16'd10912, 16'd25583, 16'd23453, 16'd60617, 16'd57521, 16'd57313, 16'd60005, 16'd3754, 16'd32883, 16'd1421, 16'd32368, 16'd61064, 16'd17272, 16'd49088, 16'd1696, 16'd26549, 16'd1023, 16'd98, 16'd45563, 16'd56149, 16'd29661});
	test_expansion(128'h980e1bca0e79f3eff9a586272cdc14c6, {16'd53217, 16'd3291, 16'd40313, 16'd22086, 16'd41738, 16'd22385, 16'd31837, 16'd42448, 16'd60293, 16'd19854, 16'd6039, 16'd13936, 16'd532, 16'd52975, 16'd46643, 16'd35064, 16'd41565, 16'd5384, 16'd43913, 16'd21185, 16'd55167, 16'd9693, 16'd33165, 16'd32031, 16'd27293, 16'd7588});
	test_expansion(128'h9987d7cd10a7946e378461ab6c5c1bd0, {16'd24899, 16'd32481, 16'd8315, 16'd49558, 16'd23053, 16'd49954, 16'd17722, 16'd32342, 16'd61739, 16'd44232, 16'd12439, 16'd37902, 16'd51927, 16'd34701, 16'd4558, 16'd34643, 16'd31962, 16'd32226, 16'd51995, 16'd43912, 16'd25003, 16'd41867, 16'd28921, 16'd61306, 16'd3089, 16'd63764});
	test_expansion(128'hab18c5adf5d35a11a643dd86abca5c58, {16'd49612, 16'd47739, 16'd62662, 16'd17509, 16'd15387, 16'd35442, 16'd34505, 16'd33847, 16'd13258, 16'd35459, 16'd6819, 16'd7107, 16'd52868, 16'd45826, 16'd65394, 16'd46283, 16'd55497, 16'd16004, 16'd15246, 16'd6193, 16'd730, 16'd55342, 16'd57871, 16'd16806, 16'd2643, 16'd10837});
	test_expansion(128'h3d9788764bac8ce536956fe24df0f3aa, {16'd31054, 16'd17209, 16'd59631, 16'd25557, 16'd826, 16'd16988, 16'd57460, 16'd19591, 16'd5663, 16'd11498, 16'd47238, 16'd42057, 16'd7129, 16'd40475, 16'd45396, 16'd58546, 16'd30401, 16'd35519, 16'd62930, 16'd38690, 16'd17632, 16'd32275, 16'd62441, 16'd44173, 16'd10670, 16'd25445});
	test_expansion(128'h43c6f866b9831f8191be81a6899e0757, {16'd31715, 16'd15756, 16'd29694, 16'd65228, 16'd52122, 16'd16386, 16'd27774, 16'd61970, 16'd7489, 16'd13703, 16'd20960, 16'd29657, 16'd11986, 16'd58281, 16'd24026, 16'd26369, 16'd15064, 16'd17115, 16'd34527, 16'd30493, 16'd27538, 16'd42513, 16'd33197, 16'd32837, 16'd52421, 16'd10716});
	test_expansion(128'h4eb34d19f5a11067b0f378ec85c291d3, {16'd62943, 16'd55672, 16'd13458, 16'd36902, 16'd46082, 16'd54998, 16'd51563, 16'd33339, 16'd25054, 16'd26114, 16'd27007, 16'd16686, 16'd42625, 16'd30667, 16'd35914, 16'd35386, 16'd51298, 16'd52969, 16'd20034, 16'd51892, 16'd14531, 16'd56995, 16'd9680, 16'd48839, 16'd15050, 16'd37823});
	test_expansion(128'had1510f35d5c21741b3ba99ddeed09d5, {16'd58791, 16'd37391, 16'd1786, 16'd21922, 16'd8573, 16'd37060, 16'd11054, 16'd11281, 16'd4893, 16'd40802, 16'd30586, 16'd35445, 16'd44843, 16'd41531, 16'd731, 16'd19955, 16'd22843, 16'd58738, 16'd25861, 16'd17260, 16'd29829, 16'd50555, 16'd20330, 16'd9902, 16'd61060, 16'd49926});
	test_expansion(128'h326f3ff9ba6a1848014d32e967a240e1, {16'd12970, 16'd2945, 16'd15385, 16'd52665, 16'd64222, 16'd51385, 16'd35053, 16'd60034, 16'd6388, 16'd64958, 16'd50642, 16'd57429, 16'd26709, 16'd43372, 16'd12930, 16'd63196, 16'd14024, 16'd24533, 16'd6206, 16'd23946, 16'd55168, 16'd21156, 16'd65119, 16'd19765, 16'd60433, 16'd65044});
	test_expansion(128'h393da5663ce92c042b082abdd63efc46, {16'd47491, 16'd52616, 16'd22413, 16'd60106, 16'd26531, 16'd33427, 16'd37528, 16'd21198, 16'd8776, 16'd11681, 16'd48986, 16'd27616, 16'd60634, 16'd36953, 16'd49105, 16'd30779, 16'd22106, 16'd42424, 16'd21293, 16'd46226, 16'd33504, 16'd62434, 16'd17937, 16'd18262, 16'd27538, 16'd4486});
	test_expansion(128'h3d05b172c7dac48ac4be195b6276a52c, {16'd40031, 16'd10655, 16'd48684, 16'd9801, 16'd40829, 16'd17411, 16'd27286, 16'd2, 16'd64966, 16'd1754, 16'd2738, 16'd17402, 16'd22682, 16'd2808, 16'd254, 16'd28193, 16'd65209, 16'd28894, 16'd11245, 16'd43901, 16'd53701, 16'd12907, 16'd29200, 16'd8549, 16'd63048, 16'd10230});
	test_expansion(128'h15de97f16b5b2909841aca0cf37ab877, {16'd42964, 16'd11056, 16'd42620, 16'd47539, 16'd7445, 16'd64591, 16'd42661, 16'd36197, 16'd5924, 16'd34290, 16'd31327, 16'd40673, 16'd7640, 16'd52573, 16'd156, 16'd17044, 16'd3672, 16'd22033, 16'd23213, 16'd2098, 16'd51004, 16'd23519, 16'd64534, 16'd16756, 16'd55978, 16'd16583});
	test_expansion(128'h0cf8dbdd8fef2f59da1b0bbc9cd0881d, {16'd28257, 16'd4375, 16'd23324, 16'd38033, 16'd10583, 16'd39144, 16'd32908, 16'd38940, 16'd50911, 16'd46599, 16'd5966, 16'd14788, 16'd22426, 16'd47307, 16'd65217, 16'd12956, 16'd50122, 16'd45588, 16'd32345, 16'd50994, 16'd48294, 16'd56627, 16'd16647, 16'd4607, 16'd24853, 16'd11574});
	test_expansion(128'h5b8b629381412a426e0f083bb56031c5, {16'd28051, 16'd24658, 16'd23924, 16'd17468, 16'd59288, 16'd9018, 16'd27197, 16'd39638, 16'd56303, 16'd61577, 16'd21814, 16'd52768, 16'd60646, 16'd11395, 16'd33239, 16'd1999, 16'd31408, 16'd43045, 16'd8949, 16'd4295, 16'd1818, 16'd43312, 16'd30086, 16'd11625, 16'd61356, 16'd6462});
	test_expansion(128'h6fdc34462bad6af184d6d124e19f3730, {16'd62180, 16'd50339, 16'd34666, 16'd22081, 16'd14072, 16'd48115, 16'd57128, 16'd148, 16'd14378, 16'd6997, 16'd37485, 16'd62454, 16'd11327, 16'd41240, 16'd2918, 16'd36099, 16'd41306, 16'd2441, 16'd62925, 16'd14008, 16'd25506, 16'd30335, 16'd65022, 16'd51752, 16'd16793, 16'd18350});
	test_expansion(128'h4192bbf39e6576e270ea4ff9fc92c973, {16'd16100, 16'd17779, 16'd31046, 16'd57018, 16'd38832, 16'd60286, 16'd8055, 16'd13526, 16'd21171, 16'd19262, 16'd23584, 16'd48736, 16'd52343, 16'd35686, 16'd37363, 16'd47466, 16'd25631, 16'd46959, 16'd64013, 16'd18237, 16'd41613, 16'd56612, 16'd15948, 16'd216, 16'd45479, 16'd32470});
	test_expansion(128'h13df4995e565200250616ee3b645b2c4, {16'd60733, 16'd42698, 16'd35386, 16'd64342, 16'd11976, 16'd29442, 16'd6470, 16'd5085, 16'd38139, 16'd53079, 16'd62798, 16'd1760, 16'd191, 16'd33015, 16'd18825, 16'd62992, 16'd52062, 16'd41818, 16'd2059, 16'd8205, 16'd16972, 16'd16214, 16'd17034, 16'd64163, 16'd49201, 16'd18555});
	test_expansion(128'h600297514a75539e928f60f867ee9507, {16'd14068, 16'd32823, 16'd34085, 16'd1702, 16'd60274, 16'd6307, 16'd28622, 16'd40394, 16'd646, 16'd38540, 16'd7724, 16'd28336, 16'd54710, 16'd26195, 16'd61701, 16'd15834, 16'd28512, 16'd11514, 16'd192, 16'd57960, 16'd38683, 16'd52780, 16'd13986, 16'd40596, 16'd3272, 16'd10808});
	test_expansion(128'h07ed83d4fed83e638fa9d8e9dd38805b, {16'd20919, 16'd47068, 16'd16228, 16'd64088, 16'd57350, 16'd32735, 16'd5427, 16'd37921, 16'd31189, 16'd38838, 16'd37880, 16'd39737, 16'd46812, 16'd18301, 16'd60501, 16'd10391, 16'd45103, 16'd57333, 16'd23894, 16'd53336, 16'd6188, 16'd54239, 16'd43165, 16'd53872, 16'd57978, 16'd18959});
	test_expansion(128'h12e944328ef18fc56d2f69ccca32c54a, {16'd58397, 16'd26661, 16'd64909, 16'd62068, 16'd47718, 16'd64711, 16'd21690, 16'd37325, 16'd10607, 16'd35510, 16'd60624, 16'd2997, 16'd54075, 16'd17147, 16'd43803, 16'd15475, 16'd62235, 16'd27910, 16'd17133, 16'd32690, 16'd3501, 16'd55674, 16'd48221, 16'd42832, 16'd32838, 16'd50580});
	test_expansion(128'hfaea9899954f5da85e4f3436c03f6679, {16'd5142, 16'd11105, 16'd9639, 16'd3561, 16'd41482, 16'd21100, 16'd1595, 16'd1370, 16'd208, 16'd63827, 16'd45014, 16'd41905, 16'd53238, 16'd33258, 16'd57413, 16'd52200, 16'd50727, 16'd16641, 16'd3735, 16'd51075, 16'd10561, 16'd38443, 16'd62650, 16'd55940, 16'd15812, 16'd49123});
	test_expansion(128'hcc80582702314c91057acbab73ff370f, {16'd33081, 16'd34479, 16'd26084, 16'd12824, 16'd39975, 16'd22648, 16'd26256, 16'd5202, 16'd3011, 16'd45953, 16'd61900, 16'd64175, 16'd15609, 16'd39564, 16'd36469, 16'd13244, 16'd48085, 16'd16286, 16'd35713, 16'd29232, 16'd62561, 16'd15003, 16'd12691, 16'd49194, 16'd3710, 16'd45194});
	test_expansion(128'h99dc201cf7b4ca45ce72371e4a74833b, {16'd11134, 16'd3552, 16'd12315, 16'd33736, 16'd15203, 16'd27379, 16'd54606, 16'd59455, 16'd35849, 16'd12265, 16'd22300, 16'd16899, 16'd47908, 16'd47306, 16'd2421, 16'd55455, 16'd27858, 16'd59243, 16'd2932, 16'd20829, 16'd38201, 16'd4997, 16'd14651, 16'd33654, 16'd36694, 16'd51812});
	test_expansion(128'hfc4a8df6fa2cc27c7ddffa3dda720a11, {16'd36427, 16'd60140, 16'd1613, 16'd1315, 16'd14973, 16'd22019, 16'd20104, 16'd3472, 16'd44001, 16'd15221, 16'd31506, 16'd17880, 16'd14949, 16'd15277, 16'd49641, 16'd12989, 16'd53847, 16'd18519, 16'd55998, 16'd22027, 16'd39268, 16'd6526, 16'd56640, 16'd30381, 16'd18711, 16'd39654});
	test_expansion(128'h6da5df04ade77482a1e54d2171bd34b0, {16'd45148, 16'd50113, 16'd48948, 16'd46763, 16'd12953, 16'd1297, 16'd12651, 16'd20588, 16'd5374, 16'd40250, 16'd29145, 16'd16960, 16'd43805, 16'd12329, 16'd63839, 16'd43323, 16'd27327, 16'd15773, 16'd44356, 16'd53847, 16'd63753, 16'd9807, 16'd4175, 16'd18567, 16'd4684, 16'd27632});
	test_expansion(128'h150039156d56cbf735e8ae48e319c73b, {16'd38836, 16'd22591, 16'd11473, 16'd27462, 16'd36567, 16'd54399, 16'd9592, 16'd4472, 16'd13866, 16'd5452, 16'd20881, 16'd7499, 16'd56051, 16'd6341, 16'd31345, 16'd519, 16'd5083, 16'd3809, 16'd61541, 16'd6698, 16'd45450, 16'd41111, 16'd37479, 16'd11949, 16'd39407, 16'd17578});
	test_expansion(128'h41b02e749765ac961828201596515258, {16'd16352, 16'd39570, 16'd30377, 16'd13404, 16'd40522, 16'd9261, 16'd33270, 16'd15472, 16'd3712, 16'd14623, 16'd31536, 16'd61784, 16'd24201, 16'd18673, 16'd14094, 16'd20629, 16'd64641, 16'd61650, 16'd9607, 16'd7303, 16'd21910, 16'd65138, 16'd2189, 16'd1791, 16'd35450, 16'd58219});
	test_expansion(128'h1d3147e0fc77a3a9979455903e2d1e88, {16'd58831, 16'd22447, 16'd42021, 16'd30953, 16'd63436, 16'd914, 16'd48334, 16'd22040, 16'd22235, 16'd5697, 16'd30269, 16'd27107, 16'd46898, 16'd62577, 16'd22951, 16'd47046, 16'd35239, 16'd45957, 16'd51726, 16'd1613, 16'd51005, 16'd32395, 16'd27315, 16'd18331, 16'd49894, 16'd55865});
	test_expansion(128'hde5ac22d1288781382dc275f8681d4a9, {16'd26756, 16'd47368, 16'd39909, 16'd5005, 16'd5524, 16'd13237, 16'd13145, 16'd3445, 16'd57810, 16'd38829, 16'd7483, 16'd44391, 16'd13782, 16'd44630, 16'd33779, 16'd22831, 16'd17069, 16'd47728, 16'd21641, 16'd54554, 16'd35596, 16'd47915, 16'd46948, 16'd62468, 16'd47251, 16'd22584});
	test_expansion(128'h47d8e624d8d05d5c8ee877dee63ef32c, {16'd39125, 16'd44180, 16'd36930, 16'd55855, 16'd53676, 16'd54452, 16'd53835, 16'd36963, 16'd50578, 16'd21343, 16'd6848, 16'd2665, 16'd42227, 16'd29287, 16'd63271, 16'd65160, 16'd7651, 16'd39497, 16'd58907, 16'd60712, 16'd60047, 16'd2751, 16'd53705, 16'd47271, 16'd58641, 16'd36273});
	test_expansion(128'h158316cfdf28757b1cfe65726483383a, {16'd3827, 16'd32711, 16'd53634, 16'd46899, 16'd16780, 16'd56557, 16'd35264, 16'd18208, 16'd46240, 16'd6334, 16'd64659, 16'd54198, 16'd25013, 16'd57118, 16'd8688, 16'd20921, 16'd44582, 16'd55326, 16'd42693, 16'd13867, 16'd60393, 16'd59101, 16'd50558, 16'd39353, 16'd27438, 16'd50775});
	test_expansion(128'h2e032eb3daaf4af12fc928f4c48c94e3, {16'd16060, 16'd22054, 16'd23988, 16'd2617, 16'd43293, 16'd42884, 16'd8474, 16'd9795, 16'd40537, 16'd38102, 16'd44061, 16'd58657, 16'd11999, 16'd19137, 16'd3611, 16'd7613, 16'd60954, 16'd13607, 16'd13443, 16'd42981, 16'd64300, 16'd48700, 16'd47267, 16'd14227, 16'd53324, 16'd32939});
	test_expansion(128'hee8dbd9b4889cf416c4327fec8146320, {16'd43228, 16'd45197, 16'd36660, 16'd25002, 16'd32529, 16'd33659, 16'd9532, 16'd31266, 16'd17023, 16'd51825, 16'd53739, 16'd55793, 16'd47593, 16'd64848, 16'd42758, 16'd57043, 16'd8807, 16'd23879, 16'd26330, 16'd14247, 16'd864, 16'd64692, 16'd1366, 16'd44715, 16'd28839, 16'd42744});
	test_expansion(128'h8d0bd86b60e297b67ac6ffbe3c66bbc9, {16'd44558, 16'd17768, 16'd33744, 16'd59210, 16'd50704, 16'd60581, 16'd32986, 16'd13429, 16'd47030, 16'd63696, 16'd18489, 16'd28708, 16'd61284, 16'd52607, 16'd1300, 16'd53594, 16'd41416, 16'd9810, 16'd13553, 16'd4234, 16'd804, 16'd34180, 16'd37155, 16'd16416, 16'd21289, 16'd63966});
	test_expansion(128'hffa52a56a11178780c3da74379c7a584, {16'd60771, 16'd13173, 16'd1829, 16'd27921, 16'd49103, 16'd63631, 16'd48697, 16'd17410, 16'd24475, 16'd939, 16'd1201, 16'd40912, 16'd22877, 16'd48283, 16'd45171, 16'd51521, 16'd20512, 16'd43030, 16'd5905, 16'd21086, 16'd13914, 16'd32137, 16'd6766, 16'd35291, 16'd55005, 16'd55844});
	test_expansion(128'h3b714757eb89eb7eb7628e537130fc8a, {16'd51870, 16'd43956, 16'd44686, 16'd31533, 16'd27430, 16'd39582, 16'd16245, 16'd28608, 16'd60452, 16'd23458, 16'd33944, 16'd44822, 16'd27446, 16'd32222, 16'd53424, 16'd53601, 16'd40507, 16'd61007, 16'd14554, 16'd44554, 16'd37311, 16'd39354, 16'd23431, 16'd58787, 16'd26507, 16'd62408});
	test_expansion(128'h9f1cc233dab8b029a33a1a3bc6bc3094, {16'd65422, 16'd28138, 16'd3574, 16'd54624, 16'd5806, 16'd36897, 16'd33542, 16'd20339, 16'd55520, 16'd30385, 16'd52146, 16'd26651, 16'd19373, 16'd57908, 16'd38464, 16'd30970, 16'd27107, 16'd58923, 16'd62060, 16'd32486, 16'd46880, 16'd45892, 16'd29075, 16'd27411, 16'd17216, 16'd29135});
	test_expansion(128'h0fb8e60a37fb2a0de0aa42417749e751, {16'd53760, 16'd17808, 16'd50900, 16'd13979, 16'd30000, 16'd36898, 16'd51202, 16'd32522, 16'd1772, 16'd9428, 16'd26958, 16'd58030, 16'd26628, 16'd3589, 16'd62049, 16'd20711, 16'd26342, 16'd62785, 16'd20041, 16'd37546, 16'd29598, 16'd23969, 16'd24118, 16'd60715, 16'd35233, 16'd29763});
	test_expansion(128'ha3c2d74f46f105f1e8a1acddfa9dce72, {16'd38696, 16'd29470, 16'd15123, 16'd49161, 16'd57877, 16'd46202, 16'd50628, 16'd32175, 16'd30723, 16'd9273, 16'd41650, 16'd37863, 16'd45090, 16'd40201, 16'd61959, 16'd1657, 16'd24240, 16'd59822, 16'd5212, 16'd12993, 16'd28838, 16'd46447, 16'd9651, 16'd32152, 16'd17273, 16'd4208});
	test_expansion(128'h80ca159fe3367316a28971ac01597f60, {16'd55603, 16'd38728, 16'd12586, 16'd46829, 16'd29743, 16'd9638, 16'd25210, 16'd55442, 16'd38843, 16'd22979, 16'd38866, 16'd3543, 16'd61597, 16'd1069, 16'd25780, 16'd18889, 16'd45251, 16'd49189, 16'd58733, 16'd57462, 16'd36890, 16'd20467, 16'd51963, 16'd33906, 16'd50185, 16'd42625});
	test_expansion(128'h4dc8c8ddb7f51755fa9cbeddce533a2a, {16'd2757, 16'd15282, 16'd33063, 16'd46471, 16'd58862, 16'd2388, 16'd56027, 16'd26842, 16'd10584, 16'd34417, 16'd11573, 16'd20787, 16'd1496, 16'd21637, 16'd46291, 16'd50131, 16'd58202, 16'd43217, 16'd62814, 16'd30811, 16'd57642, 16'd43691, 16'd37398, 16'd14331, 16'd19008, 16'd44909});
	test_expansion(128'h245947f70573862a3c823d25025fb96b, {16'd15902, 16'd25926, 16'd19067, 16'd6401, 16'd41336, 16'd18514, 16'd43680, 16'd16615, 16'd58377, 16'd35349, 16'd23844, 16'd24288, 16'd31876, 16'd62950, 16'd57359, 16'd24615, 16'd37110, 16'd60482, 16'd28315, 16'd38024, 16'd55171, 16'd20539, 16'd1246, 16'd3272, 16'd19047, 16'd58968});
	test_expansion(128'h7f639897740ee2169486c2f9b09e8743, {16'd52354, 16'd59927, 16'd58186, 16'd61853, 16'd21414, 16'd25314, 16'd48562, 16'd26037, 16'd28953, 16'd47519, 16'd44145, 16'd21813, 16'd22251, 16'd61770, 16'd51992, 16'd57482, 16'd50922, 16'd50453, 16'd15359, 16'd46404, 16'd18493, 16'd61654, 16'd13535, 16'd44321, 16'd25746, 16'd30415});
	test_expansion(128'h3f9784cb249f30cdb7fb82564d7dc85b, {16'd920, 16'd6, 16'd23241, 16'd12824, 16'd2384, 16'd46075, 16'd18307, 16'd34171, 16'd14568, 16'd20247, 16'd48373, 16'd39725, 16'd29566, 16'd50124, 16'd20490, 16'd61446, 16'd3170, 16'd28728, 16'd45616, 16'd1118, 16'd45013, 16'd2254, 16'd21946, 16'd10538, 16'd7585, 16'd31063});
	test_expansion(128'h313215f5629681f47e664e94441c63e7, {16'd11586, 16'd22866, 16'd48936, 16'd7846, 16'd18478, 16'd49601, 16'd25493, 16'd25062, 16'd55181, 16'd33113, 16'd58009, 16'd30305, 16'd49411, 16'd12776, 16'd40101, 16'd49367, 16'd41504, 16'd9824, 16'd6952, 16'd4999, 16'd29085, 16'd28111, 16'd64386, 16'd61953, 16'd45033, 16'd11927});
	test_expansion(128'h6ca5a6a213fc50aff447df5b089966d1, {16'd30368, 16'd64963, 16'd54635, 16'd32777, 16'd15278, 16'd30781, 16'd61773, 16'd42413, 16'd32098, 16'd56558, 16'd17053, 16'd31700, 16'd41402, 16'd43064, 16'd37793, 16'd32975, 16'd65047, 16'd16426, 16'd49746, 16'd24417, 16'd24295, 16'd47113, 16'd14150, 16'd34701, 16'd27648, 16'd22320});
	test_expansion(128'hdc94d4cb5ce2c44d2e3446f91a92260d, {16'd53320, 16'd50458, 16'd43473, 16'd32641, 16'd61623, 16'd1628, 16'd56299, 16'd18395, 16'd30422, 16'd55359, 16'd50069, 16'd31330, 16'd1515, 16'd38933, 16'd13560, 16'd36204, 16'd64067, 16'd36147, 16'd60461, 16'd32363, 16'd24833, 16'd18908, 16'd65353, 16'd6916, 16'd49647, 16'd25495});
	test_expansion(128'h3b0d330a8000afd5af7fe9ed9f8c7901, {16'd41863, 16'd50987, 16'd55480, 16'd230, 16'd54447, 16'd36823, 16'd57370, 16'd10826, 16'd61099, 16'd55694, 16'd15517, 16'd49192, 16'd11495, 16'd33119, 16'd32326, 16'd4562, 16'd11663, 16'd18447, 16'd21328, 16'd8554, 16'd18423, 16'd26546, 16'd42401, 16'd62402, 16'd27915, 16'd42837});
	test_expansion(128'hb9021e52d858ef3d937d758c379fa115, {16'd24197, 16'd38868, 16'd12015, 16'd22110, 16'd23473, 16'd18455, 16'd37528, 16'd55222, 16'd56288, 16'd41319, 16'd1480, 16'd40484, 16'd12523, 16'd18245, 16'd4842, 16'd25186, 16'd2947, 16'd33641, 16'd2215, 16'd22314, 16'd39982, 16'd14134, 16'd53675, 16'd21594, 16'd44519, 16'd14152});
	test_expansion(128'hacdea55cf65d6a8f72cb839fd0b82332, {16'd50210, 16'd41793, 16'd23553, 16'd45545, 16'd43539, 16'd30787, 16'd35106, 16'd21268, 16'd21645, 16'd31936, 16'd7804, 16'd59187, 16'd10468, 16'd6608, 16'd9906, 16'd1744, 16'd21027, 16'd53331, 16'd102, 16'd16891, 16'd32279, 16'd64601, 16'd22403, 16'd62373, 16'd1218, 16'd27614});
	test_expansion(128'h84753926b089a43aa24f4a51d10322c5, {16'd2514, 16'd47678, 16'd39600, 16'd44941, 16'd16214, 16'd59043, 16'd39279, 16'd34689, 16'd45888, 16'd35081, 16'd15316, 16'd60333, 16'd884, 16'd19583, 16'd34269, 16'd42606, 16'd804, 16'd5616, 16'd31794, 16'd2161, 16'd52015, 16'd47817, 16'd64806, 16'd46375, 16'd15763, 16'd51495});
	test_expansion(128'h9de55e7c525715521416eaec1fae3829, {16'd3488, 16'd13422, 16'd16699, 16'd62366, 16'd54505, 16'd31376, 16'd11127, 16'd30089, 16'd61515, 16'd15951, 16'd24565, 16'd60330, 16'd35519, 16'd31452, 16'd2524, 16'd30537, 16'd50556, 16'd973, 16'd51930, 16'd54288, 16'd45496, 16'd9759, 16'd38828, 16'd36768, 16'd682, 16'd10772});
	test_expansion(128'hbc72a3e3354861d4fe43d80e1a4cf447, {16'd43505, 16'd1406, 16'd58200, 16'd39962, 16'd31819, 16'd54574, 16'd61890, 16'd10879, 16'd42791, 16'd54807, 16'd65422, 16'd43784, 16'd59579, 16'd47257, 16'd5949, 16'd62105, 16'd12603, 16'd31371, 16'd4611, 16'd37251, 16'd63619, 16'd6118, 16'd17853, 16'd41904, 16'd22127, 16'd18807});
	test_expansion(128'hbea65a3cb107c98509854818b7801545, {16'd492, 16'd28348, 16'd2740, 16'd45339, 16'd36272, 16'd7640, 16'd43232, 16'd50418, 16'd4622, 16'd50501, 16'd35346, 16'd57973, 16'd56779, 16'd29481, 16'd53130, 16'd354, 16'd46195, 16'd60196, 16'd60005, 16'd11140, 16'd21843, 16'd16883, 16'd62506, 16'd2011, 16'd53524, 16'd28942});
	test_expansion(128'h7cdc8545f68c14a770a19edf2caa50d1, {16'd50074, 16'd53095, 16'd13440, 16'd7241, 16'd52362, 16'd39514, 16'd90, 16'd24868, 16'd4507, 16'd46797, 16'd47184, 16'd1064, 16'd33204, 16'd8246, 16'd14515, 16'd55448, 16'd16511, 16'd41054, 16'd54311, 16'd61481, 16'd9032, 16'd32509, 16'd29732, 16'd40203, 16'd20704, 16'd10972});
	test_expansion(128'h3f731f056ea0a4c05d204d8742526849, {16'd19171, 16'd41992, 16'd33139, 16'd17483, 16'd21513, 16'd17621, 16'd54214, 16'd18120, 16'd21595, 16'd33268, 16'd35708, 16'd16299, 16'd12290, 16'd65304, 16'd58312, 16'd29275, 16'd37131, 16'd47992, 16'd22145, 16'd34866, 16'd57330, 16'd42687, 16'd40977, 16'd13370, 16'd61387, 16'd37288});
	test_expansion(128'h04891d74c88f2a5eb8fa2c5b9043567c, {16'd15209, 16'd41781, 16'd57452, 16'd3795, 16'd56307, 16'd35773, 16'd24862, 16'd6606, 16'd47288, 16'd27989, 16'd15596, 16'd44371, 16'd29319, 16'd12680, 16'd51293, 16'd651, 16'd20872, 16'd17460, 16'd6379, 16'd60203, 16'd22807, 16'd26620, 16'd47280, 16'd55255, 16'd7647, 16'd27764});
	test_expansion(128'h7a1393d5c9b2cdd637d7d6f93c96909b, {16'd59207, 16'd14828, 16'd48330, 16'd43520, 16'd37647, 16'd911, 16'd1381, 16'd11374, 16'd58420, 16'd50635, 16'd51992, 16'd24327, 16'd35765, 16'd34587, 16'd12355, 16'd51632, 16'd36503, 16'd47403, 16'd9627, 16'd31482, 16'd31197, 16'd18447, 16'd23484, 16'd35429, 16'd43036, 16'd51028});
	test_expansion(128'h822c4ba9ef0125797a23debde01864e3, {16'd54469, 16'd3046, 16'd3239, 16'd41086, 16'd32987, 16'd4694, 16'd18743, 16'd4870, 16'd59197, 16'd19945, 16'd29596, 16'd19907, 16'd26172, 16'd60408, 16'd12299, 16'd58677, 16'd56713, 16'd55214, 16'd9271, 16'd43432, 16'd24798, 16'd3666, 16'd12683, 16'd9896, 16'd45576, 16'd59826});
	test_expansion(128'haae39972a5e10a7291ea70804276196d, {16'd39990, 16'd51451, 16'd56455, 16'd24129, 16'd1807, 16'd13878, 16'd9655, 16'd361, 16'd54025, 16'd15715, 16'd55847, 16'd32180, 16'd60363, 16'd27966, 16'd21707, 16'd25921, 16'd50194, 16'd16251, 16'd39522, 16'd43998, 16'd5627, 16'd60685, 16'd50394, 16'd22915, 16'd43346, 16'd38669});
	test_expansion(128'h1d6e00da0792bc2a38bf3871eeb4f42a, {16'd28572, 16'd49873, 16'd63753, 16'd19807, 16'd32576, 16'd62922, 16'd43922, 16'd60616, 16'd17581, 16'd53306, 16'd13851, 16'd12159, 16'd37188, 16'd13708, 16'd50785, 16'd20348, 16'd13421, 16'd39621, 16'd29735, 16'd18448, 16'd10816, 16'd15026, 16'd62009, 16'd33616, 16'd8553, 16'd47524});
	test_expansion(128'hd25a7894b084d6ecf7af2808809a2326, {16'd41462, 16'd55390, 16'd8342, 16'd42255, 16'd33226, 16'd19694, 16'd27744, 16'd25265, 16'd10191, 16'd30175, 16'd57425, 16'd46629, 16'd32488, 16'd19642, 16'd55882, 16'd14945, 16'd23413, 16'd32573, 16'd29999, 16'd25037, 16'd57424, 16'd47210, 16'd43349, 16'd19121, 16'd10482, 16'd19313});
	test_expansion(128'hebec895dd64d2f40869a1f3c1d989fd9, {16'd47572, 16'd52939, 16'd12063, 16'd31159, 16'd34342, 16'd65533, 16'd798, 16'd39346, 16'd41298, 16'd21366, 16'd51424, 16'd4115, 16'd22646, 16'd62184, 16'd51763, 16'd2588, 16'd41851, 16'd40205, 16'd3518, 16'd42296, 16'd62412, 16'd30355, 16'd26238, 16'd32291, 16'd27965, 16'd14743});
	test_expansion(128'hcdb9ad80bb943d3e0aad7d2a9ae48fc2, {16'd62658, 16'd39914, 16'd59136, 16'd3670, 16'd59318, 16'd28544, 16'd29507, 16'd2785, 16'd61993, 16'd26, 16'd55521, 16'd53884, 16'd9996, 16'd16021, 16'd59116, 16'd14360, 16'd56, 16'd54440, 16'd23662, 16'd35888, 16'd10995, 16'd22815, 16'd54212, 16'd426, 16'd33133, 16'd41814});
	test_expansion(128'h7a8026c02a2f871ef370c4931d4cbfd9, {16'd21201, 16'd56591, 16'd28840, 16'd39339, 16'd63307, 16'd18109, 16'd12850, 16'd34252, 16'd51232, 16'd49089, 16'd43990, 16'd42638, 16'd29642, 16'd45216, 16'd24616, 16'd59242, 16'd8956, 16'd24810, 16'd37083, 16'd56974, 16'd1499, 16'd1193, 16'd1254, 16'd45199, 16'd10945, 16'd44240});
	test_expansion(128'h488804a6f1e4c3524f200ffb781470ad, {16'd19910, 16'd65060, 16'd11579, 16'd22412, 16'd62521, 16'd47952, 16'd36039, 16'd62613, 16'd17967, 16'd27284, 16'd42562, 16'd48209, 16'd4866, 16'd2788, 16'd23890, 16'd38496, 16'd49026, 16'd49897, 16'd36262, 16'd38743, 16'd60550, 16'd50900, 16'd8377, 16'd4552, 16'd43872, 16'd54620});
	test_expansion(128'hbd7ec1fb4628e9e93c3a832ecf010eb7, {16'd50267, 16'd3311, 16'd323, 16'd1040, 16'd63625, 16'd59799, 16'd34518, 16'd47497, 16'd33871, 16'd50466, 16'd27111, 16'd29602, 16'd28627, 16'd57967, 16'd61120, 16'd40324, 16'd29449, 16'd22278, 16'd16756, 16'd49624, 16'd58840, 16'd5460, 16'd33183, 16'd59462, 16'd48082, 16'd19381});
	test_expansion(128'he45a573a5c59508cb30667efe10f3034, {16'd40985, 16'd44337, 16'd29422, 16'd52849, 16'd41908, 16'd5349, 16'd65097, 16'd26410, 16'd36441, 16'd28227, 16'd10149, 16'd12170, 16'd19804, 16'd23232, 16'd63395, 16'd48210, 16'd44987, 16'd21121, 16'd35684, 16'd50046, 16'd43751, 16'd21603, 16'd57770, 16'd18253, 16'd40590, 16'd33114});
	test_expansion(128'h11f1cfff8ecee2dc747308eec388ef15, {16'd33443, 16'd14118, 16'd64389, 16'd63812, 16'd54640, 16'd8046, 16'd17413, 16'd50361, 16'd3674, 16'd62181, 16'd23948, 16'd26881, 16'd34687, 16'd53129, 16'd63417, 16'd23094, 16'd45839, 16'd56200, 16'd47833, 16'd12083, 16'd37751, 16'd38238, 16'd17885, 16'd36446, 16'd33152, 16'd51095});
	test_expansion(128'h3a53d3f5ca1e03b55d321bf1578debf4, {16'd61584, 16'd30061, 16'd47018, 16'd44445, 16'd44542, 16'd61278, 16'd52264, 16'd24589, 16'd39976, 16'd59838, 16'd47800, 16'd64930, 16'd16353, 16'd50978, 16'd34658, 16'd27444, 16'd27254, 16'd63261, 16'd51430, 16'd43780, 16'd48812, 16'd33883, 16'd59423, 16'd46845, 16'd30381, 16'd25596});
	test_expansion(128'hcd4036808a58f4352901dcd2b1e38af9, {16'd43650, 16'd40546, 16'd16562, 16'd36255, 16'd50637, 16'd18887, 16'd37169, 16'd22989, 16'd61965, 16'd27839, 16'd11478, 16'd24369, 16'd7569, 16'd23593, 16'd2983, 16'd63651, 16'd10195, 16'd37016, 16'd26569, 16'd8527, 16'd15300, 16'd11057, 16'd35019, 16'd52643, 16'd31701, 16'd47726});
	test_expansion(128'h6499adecedb181d31fc4fa35fdb289a8, {16'd39755, 16'd35512, 16'd56953, 16'd62009, 16'd55756, 16'd52587, 16'd60065, 16'd37169, 16'd48119, 16'd54917, 16'd29684, 16'd25354, 16'd46611, 16'd36128, 16'd26708, 16'd26534, 16'd8370, 16'd4813, 16'd19793, 16'd11223, 16'd48061, 16'd56778, 16'd40592, 16'd16692, 16'd21533, 16'd6971});
	test_expansion(128'h828623788de2743e8e7faae3392d90fe, {16'd21662, 16'd3785, 16'd50746, 16'd18919, 16'd23087, 16'd60011, 16'd18024, 16'd10568, 16'd52719, 16'd49925, 16'd11043, 16'd9585, 16'd17547, 16'd53385, 16'd3091, 16'd46283, 16'd3750, 16'd44658, 16'd44934, 16'd15599, 16'd7416, 16'd3695, 16'd5619, 16'd59527, 16'd12992, 16'd57169});
	test_expansion(128'hd134903b6188ad3a2dbfa049683e2e5a, {16'd27604, 16'd32337, 16'd44592, 16'd9962, 16'd52659, 16'd44662, 16'd8159, 16'd17285, 16'd40692, 16'd22700, 16'd21776, 16'd3495, 16'd63959, 16'd54178, 16'd34984, 16'd34469, 16'd36998, 16'd14223, 16'd47239, 16'd50582, 16'd42719, 16'd21903, 16'd1545, 16'd38455, 16'd50656, 16'd24252});
	test_expansion(128'h32597835784a041b539190777c67be62, {16'd32435, 16'd15657, 16'd58620, 16'd23065, 16'd44191, 16'd23157, 16'd35163, 16'd30539, 16'd19820, 16'd43347, 16'd24164, 16'd42924, 16'd40660, 16'd19687, 16'd47483, 16'd43257, 16'd17666, 16'd12591, 16'd32601, 16'd28212, 16'd4379, 16'd13646, 16'd7236, 16'd41388, 16'd19358, 16'd682});
	test_expansion(128'hf56934f9df02d73b349bf3bb3835c7d2, {16'd51520, 16'd57081, 16'd47954, 16'd48449, 16'd14135, 16'd12515, 16'd52722, 16'd17177, 16'd24448, 16'd11968, 16'd13627, 16'd44479, 16'd45222, 16'd27836, 16'd1835, 16'd64551, 16'd59521, 16'd17031, 16'd2133, 16'd13525, 16'd54987, 16'd15089, 16'd6777, 16'd17403, 16'd36086, 16'd13613});
	test_expansion(128'h7d71833ae88a87cbf53c43196f2f0411, {16'd13065, 16'd14494, 16'd50114, 16'd40232, 16'd40177, 16'd54437, 16'd164, 16'd63670, 16'd10541, 16'd50332, 16'd9148, 16'd49768, 16'd17354, 16'd54591, 16'd33223, 16'd22656, 16'd51467, 16'd3378, 16'd64889, 16'd45768, 16'd55674, 16'd34737, 16'd55297, 16'd49481, 16'd33375, 16'd49669});
	test_expansion(128'h82db413399a218d60e929defee7e1b03, {16'd62376, 16'd60901, 16'd10332, 16'd26247, 16'd28016, 16'd44254, 16'd2228, 16'd44932, 16'd61032, 16'd45745, 16'd6359, 16'd32616, 16'd14344, 16'd29956, 16'd32057, 16'd64603, 16'd36230, 16'd22169, 16'd26925, 16'd8989, 16'd12110, 16'd19542, 16'd38969, 16'd14875, 16'd31294, 16'd64209});
	test_expansion(128'h2fcbd0b8f4f2c95a12152abe6853546b, {16'd7254, 16'd3491, 16'd53127, 16'd16353, 16'd27223, 16'd27137, 16'd13195, 16'd9685, 16'd47737, 16'd14952, 16'd17465, 16'd61750, 16'd10740, 16'd40860, 16'd12473, 16'd7856, 16'd49366, 16'd7717, 16'd42220, 16'd32028, 16'd56388, 16'd24771, 16'd58046, 16'd20443, 16'd13751, 16'd28343});
	test_expansion(128'h165f9e42d945d253d0f47ce60ba93a44, {16'd8732, 16'd12032, 16'd40828, 16'd57282, 16'd16377, 16'd17446, 16'd1295, 16'd3650, 16'd7602, 16'd33374, 16'd21039, 16'd61980, 16'd33772, 16'd47964, 16'd41503, 16'd64545, 16'd24680, 16'd54673, 16'd44157, 16'd12835, 16'd41402, 16'd2723, 16'd17165, 16'd8257, 16'd34012, 16'd52179});
	test_expansion(128'h6be965880031fc744c08509db3f71f57, {16'd53386, 16'd56630, 16'd10086, 16'd12629, 16'd34406, 16'd35404, 16'd16569, 16'd35751, 16'd26127, 16'd54815, 16'd6942, 16'd59980, 16'd27492, 16'd5265, 16'd41449, 16'd11822, 16'd27686, 16'd55801, 16'd57769, 16'd64594, 16'd59242, 16'd48042, 16'd51470, 16'd29961, 16'd41598, 16'd59542});
	test_expansion(128'h994e0eb63163f7679b74a8547d875cd6, {16'd473, 16'd63472, 16'd65386, 16'd45495, 16'd17417, 16'd14052, 16'd55784, 16'd57309, 16'd62059, 16'd51060, 16'd4989, 16'd64810, 16'd64971, 16'd16453, 16'd42078, 16'd13938, 16'd33113, 16'd18634, 16'd9248, 16'd36913, 16'd6835, 16'd64612, 16'd30708, 16'd56429, 16'd61463, 16'd63296});
	test_expansion(128'hf4df1776ec00f2f2b02619bd9e1b3652, {16'd43683, 16'd8502, 16'd50749, 16'd46666, 16'd42458, 16'd30021, 16'd6652, 16'd63884, 16'd35863, 16'd63347, 16'd14730, 16'd28969, 16'd61598, 16'd25508, 16'd25157, 16'd45675, 16'd26356, 16'd54798, 16'd10676, 16'd2684, 16'd13680, 16'd36553, 16'd48249, 16'd22921, 16'd5742, 16'd46209});
	test_expansion(128'he919d8378a0e25d5cc95adfd40ae1eb5, {16'd24764, 16'd52386, 16'd23624, 16'd33718, 16'd20192, 16'd4651, 16'd49759, 16'd56117, 16'd43977, 16'd19054, 16'd59089, 16'd56034, 16'd4447, 16'd2078, 16'd14840, 16'd64054, 16'd18873, 16'd36734, 16'd12647, 16'd52935, 16'd264, 16'd12384, 16'd37348, 16'd27121, 16'd53686, 16'd21069});
	test_expansion(128'h6cf33c4d05c7cba4ab8b4b0c3293eb7f, {16'd19819, 16'd17852, 16'd29633, 16'd4536, 16'd27764, 16'd36903, 16'd14943, 16'd53526, 16'd29553, 16'd22824, 16'd45975, 16'd6011, 16'd46498, 16'd31679, 16'd47224, 16'd21142, 16'd47942, 16'd47359, 16'd13737, 16'd2375, 16'd55448, 16'd27714, 16'd34725, 16'd11726, 16'd28057, 16'd39381});
	test_expansion(128'hca95544c564d6b38ef1591696b70df90, {16'd45957, 16'd20338, 16'd65240, 16'd46742, 16'd22198, 16'd52902, 16'd17088, 16'd26452, 16'd678, 16'd51814, 16'd16383, 16'd857, 16'd28339, 16'd50683, 16'd24094, 16'd6852, 16'd60832, 16'd65074, 16'd12600, 16'd34501, 16'd43415, 16'd35767, 16'd30635, 16'd4533, 16'd34581, 16'd44423});
	test_expansion(128'h1a5df50ca442739ccad1de2060f1b97a, {16'd41552, 16'd9184, 16'd7946, 16'd14930, 16'd11741, 16'd13786, 16'd28130, 16'd19581, 16'd65496, 16'd18044, 16'd64011, 16'd51214, 16'd56132, 16'd4617, 16'd57318, 16'd64051, 16'd20008, 16'd55856, 16'd43279, 16'd44605, 16'd38759, 16'd31445, 16'd52532, 16'd51311, 16'd59362, 16'd34233});
	test_expansion(128'h2e44cdcbdc0c7995dc8bf2a8b4718476, {16'd45999, 16'd14833, 16'd14825, 16'd7183, 16'd8690, 16'd16820, 16'd44091, 16'd4567, 16'd32443, 16'd32226, 16'd51481, 16'd12101, 16'd39581, 16'd36255, 16'd56524, 16'd31730, 16'd46132, 16'd2057, 16'd52937, 16'd23832, 16'd15631, 16'd17630, 16'd50701, 16'd18543, 16'd35641, 16'd45966});
	test_expansion(128'heba20490568f852d71c1e1b1b5a91c34, {16'd23137, 16'd9852, 16'd48292, 16'd64428, 16'd61571, 16'd51107, 16'd35441, 16'd25678, 16'd64548, 16'd45188, 16'd35109, 16'd39595, 16'd3971, 16'd29132, 16'd49277, 16'd24328, 16'd29833, 16'd6043, 16'd56860, 16'd41725, 16'd4465, 16'd59398, 16'd52871, 16'd32930, 16'd55087, 16'd23404});
	test_expansion(128'h60b70926f52f92188808db4046e8a1de, {16'd31034, 16'd7438, 16'd38948, 16'd25533, 16'd64989, 16'd48171, 16'd57850, 16'd43575, 16'd13884, 16'd56732, 16'd38664, 16'd36916, 16'd42668, 16'd65481, 16'd51684, 16'd56722, 16'd42471, 16'd38659, 16'd16356, 16'd25636, 16'd32150, 16'd44135, 16'd14368, 16'd49281, 16'd65485, 16'd49245});
	test_expansion(128'hcddef13ebf70ce527643f6456e786a84, {16'd51361, 16'd26061, 16'd3003, 16'd308, 16'd10977, 16'd37717, 16'd24167, 16'd39111, 16'd9916, 16'd13063, 16'd10420, 16'd57140, 16'd13774, 16'd21543, 16'd1877, 16'd57237, 16'd29136, 16'd21500, 16'd39289, 16'd44345, 16'd62193, 16'd23028, 16'd23496, 16'd336, 16'd18690, 16'd16230});
	test_expansion(128'hdf7c87d1adcef14cedfb4d9aab8125eb, {16'd47707, 16'd58454, 16'd14499, 16'd16587, 16'd8900, 16'd60813, 16'd63881, 16'd23372, 16'd27779, 16'd53134, 16'd10740, 16'd22904, 16'd59614, 16'd8797, 16'd55926, 16'd3525, 16'd8049, 16'd5289, 16'd1577, 16'd13567, 16'd59021, 16'd23587, 16'd29032, 16'd64517, 16'd53204, 16'd10632});
	test_expansion(128'h504dbb2c43d4f081ab0ffb50fb3607dd, {16'd1156, 16'd21745, 16'd61430, 16'd28539, 16'd52168, 16'd44217, 16'd28432, 16'd60439, 16'd27154, 16'd57602, 16'd23956, 16'd23193, 16'd54276, 16'd5458, 16'd7265, 16'd63944, 16'd37268, 16'd18892, 16'd57245, 16'd62709, 16'd61762, 16'd3624, 16'd60204, 16'd25854, 16'd23237, 16'd40802});
	test_expansion(128'hb042b560d18170290969bd894154b0aa, {16'd60246, 16'd6239, 16'd1381, 16'd19478, 16'd6972, 16'd59906, 16'd53246, 16'd56872, 16'd54831, 16'd55967, 16'd24910, 16'd41246, 16'd34868, 16'd19567, 16'd22472, 16'd57905, 16'd33115, 16'd27063, 16'd52298, 16'd30414, 16'd60115, 16'd41004, 16'd52102, 16'd25817, 16'd32799, 16'd16953});
	test_expansion(128'h09ba48dd88a3904a18f52e8e0ed5e790, {16'd63055, 16'd10881, 16'd826, 16'd54270, 16'd50914, 16'd14060, 16'd7620, 16'd61092, 16'd23314, 16'd49219, 16'd42837, 16'd39967, 16'd21056, 16'd62605, 16'd45715, 16'd3381, 16'd2694, 16'd17865, 16'd21728, 16'd40052, 16'd2925, 16'd58126, 16'd23900, 16'd54735, 16'd34837, 16'd293});
	test_expansion(128'h9149ae3038ddcd0eda62dab4416398da, {16'd53055, 16'd27465, 16'd59858, 16'd2023, 16'd45481, 16'd64769, 16'd40913, 16'd11257, 16'd16711, 16'd24287, 16'd38562, 16'd23656, 16'd5693, 16'd46605, 16'd53280, 16'd49304, 16'd4859, 16'd45927, 16'd39393, 16'd11302, 16'd53433, 16'd26525, 16'd8638, 16'd23169, 16'd18974, 16'd14030});
	test_expansion(128'h1d8520fa7b26576b7b71b3d09450adff, {16'd48513, 16'd53642, 16'd59170, 16'd18644, 16'd18399, 16'd9880, 16'd58172, 16'd13956, 16'd47103, 16'd26174, 16'd3418, 16'd39359, 16'd63855, 16'd4905, 16'd18538, 16'd33006, 16'd63173, 16'd48024, 16'd13367, 16'd45509, 16'd53148, 16'd60185, 16'd21347, 16'd46050, 16'd20162, 16'd34355});
	test_expansion(128'h8a95aeb147b690eb79fd0996ce742225, {16'd47058, 16'd22482, 16'd55015, 16'd990, 16'd45512, 16'd54691, 16'd9360, 16'd59024, 16'd10374, 16'd1665, 16'd10980, 16'd34163, 16'd8044, 16'd18031, 16'd28492, 16'd63851, 16'd14434, 16'd61744, 16'd31829, 16'd17343, 16'd41407, 16'd46580, 16'd37638, 16'd15897, 16'd18047, 16'd61522});
	test_expansion(128'hfab9fd09960a25178cbcd2deb7b5315c, {16'd35404, 16'd29915, 16'd19630, 16'd36844, 16'd16783, 16'd38328, 16'd54715, 16'd64560, 16'd38051, 16'd23049, 16'd42563, 16'd57035, 16'd60655, 16'd48518, 16'd24586, 16'd2341, 16'd5976, 16'd13257, 16'd47601, 16'd16898, 16'd41025, 16'd61714, 16'd24823, 16'd30132, 16'd29587, 16'd64506});
	test_expansion(128'hc2c308422ce7e35111718a972eebeee2, {16'd65250, 16'd35016, 16'd17631, 16'd57499, 16'd41770, 16'd64251, 16'd57501, 16'd12772, 16'd23361, 16'd33161, 16'd64784, 16'd35199, 16'd43342, 16'd20418, 16'd57335, 16'd50121, 16'd17456, 16'd52916, 16'd52293, 16'd34789, 16'd60442, 16'd38105, 16'd33944, 16'd28287, 16'd37465, 16'd19397});
	test_expansion(128'hcb479850d3d9d49195d92a0b7c12872d, {16'd40447, 16'd22934, 16'd22933, 16'd38675, 16'd26185, 16'd51567, 16'd64975, 16'd7223, 16'd11104, 16'd61485, 16'd37835, 16'd44238, 16'd10367, 16'd20787, 16'd8481, 16'd8037, 16'd44120, 16'd61225, 16'd6877, 16'd29358, 16'd33164, 16'd50580, 16'd5684, 16'd18248, 16'd50091, 16'd35772});
	test_expansion(128'h7baf76a2de89f01f4584b529710157d2, {16'd4436, 16'd6515, 16'd15427, 16'd56253, 16'd30565, 16'd6555, 16'd559, 16'd51777, 16'd338, 16'd38117, 16'd28012, 16'd14337, 16'd22380, 16'd13966, 16'd57627, 16'd24738, 16'd31811, 16'd62978, 16'd6640, 16'd6815, 16'd21306, 16'd53781, 16'd60239, 16'd29566, 16'd36038, 16'd7197});
	test_expansion(128'hc26d608368bb440dcec420413cf3f5d3, {16'd18449, 16'd53810, 16'd28520, 16'd47116, 16'd58635, 16'd52214, 16'd13290, 16'd20236, 16'd48466, 16'd54737, 16'd5242, 16'd22498, 16'd37169, 16'd37565, 16'd59522, 16'd58248, 16'd53940, 16'd9185, 16'd45126, 16'd524, 16'd10275, 16'd2812, 16'd51303, 16'd12045, 16'd10825, 16'd44393});
	test_expansion(128'h858dc7d8dcf0bfdd7dab4b5d8749de62, {16'd62902, 16'd42501, 16'd28657, 16'd5728, 16'd20535, 16'd64079, 16'd61060, 16'd61460, 16'd20631, 16'd38048, 16'd43456, 16'd55199, 16'd17533, 16'd12538, 16'd32926, 16'd33733, 16'd21753, 16'd14302, 16'd45562, 16'd39437, 16'd64734, 16'd61438, 16'd28076, 16'd37868, 16'd59926, 16'd42753});
	test_expansion(128'hfae7478b7a6362c5c11ea7f32ef1c615, {16'd56759, 16'd41209, 16'd57184, 16'd49713, 16'd50083, 16'd48874, 16'd56945, 16'd10952, 16'd9559, 16'd19190, 16'd15237, 16'd63970, 16'd20152, 16'd7024, 16'd2745, 16'd64575, 16'd51864, 16'd58102, 16'd13642, 16'd20007, 16'd8711, 16'd10628, 16'd31103, 16'd55373, 16'd34777, 16'd56218});
	test_expansion(128'hffff638ed4601764df9d62354321e012, {16'd19681, 16'd29649, 16'd40286, 16'd59602, 16'd40939, 16'd53312, 16'd46361, 16'd46054, 16'd58597, 16'd7128, 16'd47918, 16'd61833, 16'd38004, 16'd53635, 16'd59714, 16'd44684, 16'd23729, 16'd45876, 16'd7127, 16'd64341, 16'd60243, 16'd2217, 16'd40630, 16'd55088, 16'd30014, 16'd18265});
	test_expansion(128'h4aff745f1c546c3a22baf1444c89265d, {16'd19359, 16'd47441, 16'd63850, 16'd15881, 16'd34104, 16'd53125, 16'd234, 16'd55497, 16'd13457, 16'd51362, 16'd40658, 16'd3892, 16'd64469, 16'd14255, 16'd8845, 16'd41974, 16'd38366, 16'd58849, 16'd18671, 16'd15975, 16'd30819, 16'd40474, 16'd54849, 16'd30256, 16'd27072, 16'd40658});
	test_expansion(128'h3d10536bcfe113a65468d9bae1232e41, {16'd63751, 16'd5610, 16'd58996, 16'd27991, 16'd33173, 16'd16035, 16'd48669, 16'd20204, 16'd24615, 16'd11286, 16'd19200, 16'd28813, 16'd10196, 16'd36361, 16'd31173, 16'd47856, 16'd9165, 16'd61156, 16'd21627, 16'd25238, 16'd8137, 16'd39731, 16'd27171, 16'd61374, 16'd22828, 16'd10428});
	test_expansion(128'ha4b9202ca25b3c97456ae0857ff2b476, {16'd54559, 16'd32290, 16'd51443, 16'd11614, 16'd36569, 16'd61221, 16'd3134, 16'd54291, 16'd56134, 16'd7386, 16'd15874, 16'd53501, 16'd25765, 16'd57531, 16'd31493, 16'd11040, 16'd31740, 16'd52273, 16'd62590, 16'd2133, 16'd56137, 16'd54356, 16'd23213, 16'd54346, 16'd29024, 16'd13839});
	test_expansion(128'h837d65c9869a5ac0d84eef9af70770b6, {16'd865, 16'd26200, 16'd15172, 16'd21083, 16'd15143, 16'd18603, 16'd46330, 16'd14584, 16'd57163, 16'd54712, 16'd49265, 16'd37404, 16'd32882, 16'd53585, 16'd27352, 16'd5468, 16'd22069, 16'd37732, 16'd32755, 16'd58368, 16'd49881, 16'd16829, 16'd1229, 16'd37697, 16'd13713, 16'd50819});
	test_expansion(128'hae4b98df083e8a5d40d15a6b36f991e8, {16'd43144, 16'd15503, 16'd1277, 16'd30718, 16'd51092, 16'd44021, 16'd60214, 16'd52637, 16'd6023, 16'd10306, 16'd38686, 16'd22667, 16'd23719, 16'd46004, 16'd26024, 16'd34218, 16'd59293, 16'd34867, 16'd42867, 16'd42495, 16'd54908, 16'd26690, 16'd46101, 16'd20716, 16'd36038, 16'd51634});
	test_expansion(128'h798cfcb7f6f439f4e62ec996f47ab79e, {16'd58272, 16'd7613, 16'd53947, 16'd50391, 16'd56687, 16'd39237, 16'd25013, 16'd29516, 16'd58217, 16'd61791, 16'd34397, 16'd11338, 16'd25578, 16'd10718, 16'd20546, 16'd52001, 16'd48612, 16'd17523, 16'd17838, 16'd63402, 16'd46169, 16'd13604, 16'd3083, 16'd2835, 16'd35857, 16'd23480});
	test_expansion(128'h9a20ef024416f537ec13c19bc97449fd, {16'd48517, 16'd49643, 16'd2268, 16'd65413, 16'd8589, 16'd58997, 16'd17018, 16'd9068, 16'd31700, 16'd35694, 16'd33894, 16'd28194, 16'd41545, 16'd25237, 16'd64817, 16'd58633, 16'd13668, 16'd17862, 16'd56339, 16'd25676, 16'd23889, 16'd54489, 16'd30876, 16'd57714, 16'd262, 16'd30121});
	test_expansion(128'h2565aadaa863115b1ab7b6bec4d026ef, {16'd2578, 16'd44467, 16'd42779, 16'd55225, 16'd44219, 16'd52172, 16'd23865, 16'd37484, 16'd8118, 16'd41971, 16'd11586, 16'd3289, 16'd37560, 16'd2377, 16'd27953, 16'd58566, 16'd57755, 16'd9389, 16'd28620, 16'd28556, 16'd32910, 16'd33038, 16'd21988, 16'd51791, 16'd4609, 16'd41904});
	test_expansion(128'h0844502c15f368a6c019959831f03e3b, {16'd8681, 16'd25410, 16'd45177, 16'd59189, 16'd10329, 16'd23834, 16'd30950, 16'd58416, 16'd48154, 16'd36567, 16'd40060, 16'd31677, 16'd8513, 16'd35025, 16'd6290, 16'd50060, 16'd16339, 16'd13469, 16'd46248, 16'd61630, 16'd51919, 16'd34469, 16'd39738, 16'd17409, 16'd39875, 16'd58554});
	test_expansion(128'h6648eaa11a383896c71a09454f8c6999, {16'd39471, 16'd10205, 16'd5448, 16'd17818, 16'd50495, 16'd16280, 16'd2380, 16'd64180, 16'd44822, 16'd29848, 16'd23178, 16'd30911, 16'd48938, 16'd50227, 16'd40375, 16'd32526, 16'd53546, 16'd58318, 16'd48038, 16'd1163, 16'd8158, 16'd62815, 16'd2811, 16'd27368, 16'd52727, 16'd58303});
	test_expansion(128'ha0663b3c6c1d2440e3554d2705b5f7c7, {16'd52800, 16'd2252, 16'd18036, 16'd53789, 16'd58272, 16'd45287, 16'd13191, 16'd48791, 16'd10529, 16'd30823, 16'd50840, 16'd26532, 16'd1900, 16'd933, 16'd32788, 16'd50383, 16'd40420, 16'd24543, 16'd38047, 16'd60788, 16'd22148, 16'd21995, 16'd34397, 16'd6910, 16'd29164, 16'd5733});
	test_expansion(128'h7d0750163decb5b72e544ba9b48fa333, {16'd47425, 16'd2470, 16'd39087, 16'd27920, 16'd7413, 16'd17581, 16'd53341, 16'd41878, 16'd6202, 16'd13023, 16'd6760, 16'd45487, 16'd63639, 16'd7128, 16'd60031, 16'd39699, 16'd2899, 16'd56029, 16'd44697, 16'd54771, 16'd12320, 16'd17337, 16'd30551, 16'd5534, 16'd47665, 16'd31322});
	test_expansion(128'hcc76787b07b25271b402220f3893a21f, {16'd34565, 16'd5882, 16'd5949, 16'd28514, 16'd47610, 16'd4815, 16'd33292, 16'd14067, 16'd32499, 16'd56124, 16'd10637, 16'd30582, 16'd61599, 16'd40261, 16'd42609, 16'd61207, 16'd54939, 16'd44587, 16'd22401, 16'd34773, 16'd31445, 16'd48409, 16'd35909, 16'd4793, 16'd58081, 16'd32680});
	test_expansion(128'h0794adda90d2bc238df26fc869eed635, {16'd9181, 16'd21913, 16'd59955, 16'd62964, 16'd37316, 16'd33257, 16'd43793, 16'd19796, 16'd5249, 16'd38697, 16'd4035, 16'd53058, 16'd26538, 16'd45679, 16'd10740, 16'd52541, 16'd17622, 16'd8541, 16'd51106, 16'd32071, 16'd499, 16'd58233, 16'd37709, 16'd10779, 16'd19662, 16'd53768});
	test_expansion(128'ha4d2e3caac4dce102e6d9d6c7f826140, {16'd59503, 16'd15856, 16'd22750, 16'd63435, 16'd20120, 16'd49185, 16'd16380, 16'd31311, 16'd18472, 16'd61761, 16'd33248, 16'd26563, 16'd64898, 16'd63948, 16'd12753, 16'd59969, 16'd27925, 16'd36926, 16'd55521, 16'd59363, 16'd51175, 16'd36182, 16'd13413, 16'd17140, 16'd2774, 16'd1852});
	test_expansion(128'ha20977f6077fb37a00226bd8b0acebdd, {16'd29478, 16'd23237, 16'd7100, 16'd2694, 16'd34262, 16'd55925, 16'd32106, 16'd41030, 16'd9624, 16'd62882, 16'd53472, 16'd5802, 16'd50815, 16'd36779, 16'd57199, 16'd8455, 16'd36406, 16'd9126, 16'd32028, 16'd22863, 16'd15099, 16'd45397, 16'd10650, 16'd30584, 16'd27132, 16'd26054});
	test_expansion(128'hafc1d18e4f8cddff4c6d49e464710262, {16'd48535, 16'd6898, 16'd58068, 16'd11001, 16'd35125, 16'd27290, 16'd36934, 16'd31721, 16'd17188, 16'd58421, 16'd32752, 16'd22792, 16'd61230, 16'd27426, 16'd50716, 16'd14718, 16'd49017, 16'd40542, 16'd38071, 16'd3648, 16'd2401, 16'd22332, 16'd59298, 16'd44088, 16'd44004, 16'd1630});
	test_expansion(128'h654a148d8cfb17aba82e11602c2576a2, {16'd60230, 16'd10957, 16'd45466, 16'd21492, 16'd43337, 16'd14456, 16'd55998, 16'd56276, 16'd23356, 16'd44745, 16'd8035, 16'd34242, 16'd41085, 16'd18691, 16'd55974, 16'd36256, 16'd64135, 16'd54243, 16'd49221, 16'd27669, 16'd13387, 16'd14658, 16'd28303, 16'd52474, 16'd8726, 16'd28960});
	test_expansion(128'h3aaa58fe55114eec3910449146d454c1, {16'd44659, 16'd40424, 16'd23550, 16'd41581, 16'd62471, 16'd63849, 16'd30371, 16'd9213, 16'd8066, 16'd19384, 16'd23504, 16'd42610, 16'd19799, 16'd39331, 16'd3666, 16'd17189, 16'd19325, 16'd12396, 16'd49486, 16'd32948, 16'd40146, 16'd28802, 16'd40547, 16'd2786, 16'd40474, 16'd44903});
	test_expansion(128'h081317a5ce6175d51a52f799e4e8d9ff, {16'd2116, 16'd52855, 16'd10610, 16'd12704, 16'd5977, 16'd12813, 16'd34583, 16'd48408, 16'd2647, 16'd23950, 16'd6223, 16'd56877, 16'd16541, 16'd55200, 16'd7910, 16'd5494, 16'd50632, 16'd8090, 16'd53892, 16'd32176, 16'd3954, 16'd39895, 16'd32527, 16'd62205, 16'd10944, 16'd55300});
	test_expansion(128'h741dd125467a839d1302248a6cc07728, {16'd8607, 16'd55028, 16'd32803, 16'd55226, 16'd16293, 16'd62950, 16'd24767, 16'd64837, 16'd32115, 16'd12651, 16'd55905, 16'd62702, 16'd15779, 16'd18191, 16'd872, 16'd24885, 16'd13565, 16'd27398, 16'd17279, 16'd32838, 16'd50408, 16'd49557, 16'd63525, 16'd57051, 16'd30266, 16'd23868});
	test_expansion(128'ha3b96209978a7cf5ebf8ed0f6915212e, {16'd64936, 16'd11537, 16'd8568, 16'd11523, 16'd62928, 16'd23608, 16'd59106, 16'd22854, 16'd17125, 16'd9873, 16'd3322, 16'd12742, 16'd3098, 16'd12564, 16'd63263, 16'd40292, 16'd17792, 16'd52618, 16'd56071, 16'd48781, 16'd22302, 16'd23238, 16'd29337, 16'd55469, 16'd56339, 16'd17599});
	test_expansion(128'hf1444788ab0b4adb06ae2b1d3f1bd68d, {16'd44245, 16'd60611, 16'd44181, 16'd58542, 16'd61262, 16'd60340, 16'd47072, 16'd1894, 16'd16146, 16'd60298, 16'd23537, 16'd7734, 16'd58398, 16'd37467, 16'd55679, 16'd44720, 16'd27501, 16'd21333, 16'd60547, 16'd24747, 16'd31312, 16'd37984, 16'd64101, 16'd26659, 16'd59234, 16'd14235});
	test_expansion(128'h2e784e716348c18cc3acc97c04ae1557, {16'd17331, 16'd31841, 16'd8850, 16'd47299, 16'd21230, 16'd53810, 16'd20095, 16'd50662, 16'd13823, 16'd51371, 16'd52684, 16'd25755, 16'd9184, 16'd19656, 16'd20758, 16'd49434, 16'd41973, 16'd13457, 16'd434, 16'd48014, 16'd61712, 16'd1893, 16'd7586, 16'd20760, 16'd55193, 16'd39169});
	test_expansion(128'h9a52d15c3ffba95f50334df9246589cc, {16'd52492, 16'd62837, 16'd65250, 16'd37504, 16'd52271, 16'd8892, 16'd25834, 16'd38037, 16'd37227, 16'd62218, 16'd6967, 16'd21117, 16'd18204, 16'd43210, 16'd44219, 16'd33782, 16'd34911, 16'd9359, 16'd10997, 16'd21208, 16'd357, 16'd44520, 16'd62345, 16'd50373, 16'd50909, 16'd26199});
	test_expansion(128'h7b8674dae7bba524620d5013de3953ae, {16'd6288, 16'd48983, 16'd40369, 16'd31999, 16'd35475, 16'd45015, 16'd8731, 16'd55381, 16'd27899, 16'd15511, 16'd59865, 16'd32227, 16'd11217, 16'd26612, 16'd37021, 16'd17958, 16'd34283, 16'd65191, 16'd29406, 16'd17, 16'd23323, 16'd62671, 16'd47816, 16'd28963, 16'd8099, 16'd52790});
	test_expansion(128'h2b5cc21bdd997c1ec81e8cb08fe22ce5, {16'd20385, 16'd64458, 16'd53862, 16'd30498, 16'd24328, 16'd13416, 16'd21236, 16'd56525, 16'd52148, 16'd29770, 16'd20050, 16'd37993, 16'd22668, 16'd52670, 16'd28449, 16'd24102, 16'd52262, 16'd39289, 16'd27612, 16'd29709, 16'd10291, 16'd40623, 16'd41186, 16'd14752, 16'd29408, 16'd36589});
	test_expansion(128'h523b7c3e3e7823a8b5482a2146ef5234, {16'd24456, 16'd45630, 16'd1209, 16'd62480, 16'd8897, 16'd49843, 16'd62494, 16'd42645, 16'd12038, 16'd14807, 16'd20492, 16'd30517, 16'd58189, 16'd27994, 16'd27386, 16'd34356, 16'd5693, 16'd4367, 16'd49822, 16'd28602, 16'd48609, 16'd14174, 16'd11858, 16'd63778, 16'd41519, 16'd54439});
	test_expansion(128'hdcceadfb4d49353a9c0cd74ef80b19f5, {16'd42050, 16'd10765, 16'd39064, 16'd17830, 16'd11214, 16'd18985, 16'd35070, 16'd7843, 16'd39011, 16'd1076, 16'd25086, 16'd55000, 16'd28305, 16'd56096, 16'd33082, 16'd37876, 16'd37372, 16'd16827, 16'd57294, 16'd52419, 16'd29533, 16'd41114, 16'd42137, 16'd33006, 16'd51180, 16'd20002});
	test_expansion(128'h108f0bb90ff3d8764e3af1673725ac41, {16'd22302, 16'd50101, 16'd29884, 16'd62021, 16'd43768, 16'd3007, 16'd19603, 16'd36139, 16'd12189, 16'd62246, 16'd1840, 16'd27627, 16'd4012, 16'd27328, 16'd33419, 16'd35333, 16'd36889, 16'd17358, 16'd15925, 16'd57984, 16'd26770, 16'd43357, 16'd17653, 16'd56306, 16'd11750, 16'd52177});
	test_expansion(128'hcfa45deaa2642d2cf1b61226022c57e1, {16'd38343, 16'd57848, 16'd39185, 16'd9601, 16'd24050, 16'd59372, 16'd49935, 16'd10275, 16'd20664, 16'd30496, 16'd6290, 16'd35565, 16'd8909, 16'd57560, 16'd37511, 16'd11608, 16'd39437, 16'd2658, 16'd16584, 16'd26408, 16'd11403, 16'd53459, 16'd55800, 16'd43753, 16'd47043, 16'd8867});
	test_expansion(128'h80ed430492910248cee4bdc444580ce3, {16'd47976, 16'd41123, 16'd36522, 16'd63593, 16'd29092, 16'd15991, 16'd17864, 16'd42524, 16'd6830, 16'd50939, 16'd45788, 16'd37030, 16'd53592, 16'd57936, 16'd57760, 16'd6521, 16'd27573, 16'd22502, 16'd11382, 16'd50494, 16'd63455, 16'd44560, 16'd27414, 16'd22053, 16'd4042, 16'd21965});
	test_expansion(128'h4e66d6a4542f4a951a9872561dbf5e8d, {16'd166, 16'd2082, 16'd30250, 16'd4015, 16'd38142, 16'd15284, 16'd64789, 16'd58384, 16'd30801, 16'd23613, 16'd22841, 16'd25688, 16'd27099, 16'd48695, 16'd38987, 16'd22608, 16'd48272, 16'd55311, 16'd11887, 16'd61066, 16'd36560, 16'd5660, 16'd16927, 16'd15653, 16'd48228, 16'd55284});
	test_expansion(128'h76e9ce847a85ce0cb7fc3295d7f01b2f, {16'd53987, 16'd59688, 16'd9140, 16'd29632, 16'd6474, 16'd29623, 16'd60503, 16'd53018, 16'd24107, 16'd42127, 16'd36327, 16'd10695, 16'd40129, 16'd24302, 16'd13369, 16'd16747, 16'd49181, 16'd5253, 16'd10989, 16'd2192, 16'd24803, 16'd31036, 16'd16861, 16'd563, 16'd10276, 16'd39364});
	test_expansion(128'he1480c42d6c56f1292fc0c8a559fd2ee, {16'd36797, 16'd54070, 16'd50066, 16'd47082, 16'd9747, 16'd32065, 16'd32588, 16'd57100, 16'd18005, 16'd41382, 16'd6739, 16'd54494, 16'd12944, 16'd13519, 16'd38435, 16'd3626, 16'd2763, 16'd25871, 16'd26744, 16'd57333, 16'd21243, 16'd17454, 16'd47806, 16'd8874, 16'd15587, 16'd24628});
	test_expansion(128'h1c6b455c39b80345195519fd76d34ec7, {16'd38556, 16'd56671, 16'd65496, 16'd30613, 16'd777, 16'd24374, 16'd64555, 16'd13545, 16'd38600, 16'd64122, 16'd25646, 16'd12992, 16'd6907, 16'd50575, 16'd5461, 16'd60549, 16'd45190, 16'd45574, 16'd14504, 16'd64926, 16'd8719, 16'd19377, 16'd37925, 16'd18665, 16'd55736, 16'd20074});
	test_expansion(128'hefe8233cdb58dcc7c104aefa4c8e6329, {16'd739, 16'd10359, 16'd40101, 16'd34035, 16'd52109, 16'd9425, 16'd32916, 16'd60928, 16'd8013, 16'd56767, 16'd51306, 16'd36992, 16'd38039, 16'd61438, 16'd61957, 16'd24555, 16'd37594, 16'd52892, 16'd13886, 16'd20992, 16'd28589, 16'd1046, 16'd58774, 16'd28339, 16'd39705, 16'd175});
	test_expansion(128'hecf423482523f32d332b5c1e32a84ecf, {16'd43281, 16'd7461, 16'd45999, 16'd2584, 16'd60262, 16'd63063, 16'd9560, 16'd753, 16'd48038, 16'd48586, 16'd7465, 16'd55536, 16'd54698, 16'd3331, 16'd2717, 16'd43830, 16'd21306, 16'd58835, 16'd4071, 16'd20666, 16'd46461, 16'd36087, 16'd26629, 16'd44531, 16'd17890, 16'd64767});
	test_expansion(128'h01be69a94c9486c661df4d4dcc7605ec, {16'd15223, 16'd57040, 16'd22744, 16'd19187, 16'd37708, 16'd39055, 16'd35612, 16'd35049, 16'd26686, 16'd10654, 16'd15307, 16'd14763, 16'd1225, 16'd39418, 16'd18726, 16'd21875, 16'd28337, 16'd34396, 16'd32273, 16'd50278, 16'd4020, 16'd31521, 16'd59262, 16'd30261, 16'd43787, 16'd43957});
	test_expansion(128'haa6c2d0bc4926cc0f81714234b728e7b, {16'd33360, 16'd57485, 16'd59328, 16'd31458, 16'd46727, 16'd50928, 16'd48960, 16'd37525, 16'd4054, 16'd50188, 16'd17265, 16'd23663, 16'd18349, 16'd13436, 16'd61896, 16'd2832, 16'd63191, 16'd36632, 16'd37986, 16'd8077, 16'd23553, 16'd1490, 16'd48503, 16'd30715, 16'd16725, 16'd54153});
	test_expansion(128'hc94899713184d7dc0868ac79fe0010ef, {16'd26736, 16'd31919, 16'd26476, 16'd36722, 16'd32189, 16'd17028, 16'd46404, 16'd37993, 16'd13694, 16'd8624, 16'd61266, 16'd43586, 16'd59252, 16'd30485, 16'd40984, 16'd5012, 16'd60589, 16'd50255, 16'd43515, 16'd7888, 16'd33663, 16'd52171, 16'd48459, 16'd12407, 16'd47978, 16'd60847});
	test_expansion(128'h85c0e766cbc72e8d1ed0c4dceeafc6a9, {16'd36492, 16'd61823, 16'd32125, 16'd37400, 16'd64034, 16'd54516, 16'd41132, 16'd51570, 16'd19284, 16'd44574, 16'd47221, 16'd59606, 16'd25029, 16'd61586, 16'd13766, 16'd15908, 16'd49377, 16'd47813, 16'd4110, 16'd28180, 16'd32387, 16'd45501, 16'd1067, 16'd12135, 16'd7191, 16'd50359});
	test_expansion(128'hb18cb933e9819a704376e440ba3bfb14, {16'd44522, 16'd2586, 16'd49675, 16'd57597, 16'd38492, 16'd56893, 16'd4059, 16'd43384, 16'd2635, 16'd57984, 16'd12454, 16'd61454, 16'd26572, 16'd7950, 16'd62304, 16'd47418, 16'd734, 16'd51034, 16'd22902, 16'd59927, 16'd17980, 16'd29174, 16'd33415, 16'd39549, 16'd50373, 16'd45152});
	test_expansion(128'h240238098653ebbc5ac4c779026de70d, {16'd59595, 16'd32368, 16'd33471, 16'd42200, 16'd56093, 16'd47318, 16'd6206, 16'd30847, 16'd55899, 16'd64437, 16'd47560, 16'd52748, 16'd14298, 16'd32874, 16'd40084, 16'd7340, 16'd42282, 16'd8482, 16'd485, 16'd54477, 16'd41178, 16'd44394, 16'd44313, 16'd9138, 16'd44158, 16'd759});
	test_expansion(128'hc179f5cd459b0a52e6375374280d79cf, {16'd56601, 16'd12170, 16'd6801, 16'd31916, 16'd19603, 16'd50624, 16'd3504, 16'd28271, 16'd25084, 16'd7115, 16'd29184, 16'd21087, 16'd23374, 16'd61173, 16'd58872, 16'd264, 16'd62753, 16'd14154, 16'd8215, 16'd51175, 16'd29592, 16'd60458, 16'd7900, 16'd48518, 16'd46495, 16'd39084});
	test_expansion(128'hc65d9a5e40130ca73b4aa4452e73fe20, {16'd45607, 16'd56789, 16'd54448, 16'd23411, 16'd43210, 16'd11971, 16'd51750, 16'd47566, 16'd52761, 16'd36991, 16'd32090, 16'd49472, 16'd39162, 16'd44304, 16'd17430, 16'd1692, 16'd3832, 16'd746, 16'd43539, 16'd3272, 16'd26497, 16'd2865, 16'd3160, 16'd32704, 16'd3974, 16'd15673});
	test_expansion(128'hdd1021a32f0bd304f265bedfc318eb98, {16'd59499, 16'd56142, 16'd37735, 16'd15273, 16'd27, 16'd58554, 16'd57226, 16'd6623, 16'd41081, 16'd41177, 16'd14703, 16'd28247, 16'd52749, 16'd4847, 16'd7366, 16'd22994, 16'd48235, 16'd16613, 16'd40629, 16'd42499, 16'd61838, 16'd64579, 16'd55890, 16'd58569, 16'd41731, 16'd4263});
	test_expansion(128'h464e2da7b995fefcb0d3088e461f559d, {16'd22706, 16'd60401, 16'd46010, 16'd10360, 16'd48047, 16'd34780, 16'd28790, 16'd8711, 16'd26003, 16'd12561, 16'd35685, 16'd46775, 16'd40918, 16'd62566, 16'd13545, 16'd41279, 16'd7732, 16'd23825, 16'd51569, 16'd61801, 16'd20269, 16'd60743, 16'd7112, 16'd46449, 16'd58719, 16'd57309});
	test_expansion(128'hbf1b33b9d7627a5fabb1ed5e00216903, {16'd16671, 16'd59703, 16'd20351, 16'd19800, 16'd60551, 16'd4825, 16'd11886, 16'd47277, 16'd21678, 16'd40559, 16'd64794, 16'd17742, 16'd22608, 16'd37971, 16'd47885, 16'd30415, 16'd25200, 16'd64004, 16'd48928, 16'd38951, 16'd10090, 16'd30056, 16'd37136, 16'd23298, 16'd7805, 16'd12167});
	test_expansion(128'h5fdff825d9b7d139e62537ca3663faf0, {16'd9762, 16'd50828, 16'd23068, 16'd41045, 16'd30711, 16'd13025, 16'd15333, 16'd30628, 16'd17307, 16'd42182, 16'd40098, 16'd62540, 16'd2881, 16'd46664, 16'd8173, 16'd49041, 16'd900, 16'd56952, 16'd26666, 16'd6596, 16'd52350, 16'd41849, 16'd36036, 16'd51808, 16'd52726, 16'd57527});
	test_expansion(128'h229538bf8ebce3fce322997bc26e0cda, {16'd3465, 16'd10417, 16'd45690, 16'd2949, 16'd59570, 16'd281, 16'd46131, 16'd59538, 16'd11959, 16'd28045, 16'd17211, 16'd27933, 16'd7838, 16'd25757, 16'd49272, 16'd52302, 16'd49691, 16'd35583, 16'd6614, 16'd30513, 16'd23064, 16'd63866, 16'd29429, 16'd30753, 16'd8361, 16'd25640});
	test_expansion(128'h076d1aedaac7ed210852b2a210202ea6, {16'd44594, 16'd19423, 16'd58448, 16'd8177, 16'd59108, 16'd28932, 16'd47035, 16'd19257, 16'd25290, 16'd60241, 16'd33714, 16'd4143, 16'd8235, 16'd50510, 16'd2845, 16'd59221, 16'd21029, 16'd9989, 16'd55194, 16'd44237, 16'd12263, 16'd61304, 16'd17216, 16'd38299, 16'd14707, 16'd40473});
	test_expansion(128'he8cb41f05dd860482e5772c3f25594f2, {16'd15152, 16'd44358, 16'd16174, 16'd23079, 16'd26451, 16'd42873, 16'd60385, 16'd11621, 16'd61413, 16'd62300, 16'd52718, 16'd26467, 16'd16652, 16'd28835, 16'd4786, 16'd10162, 16'd14188, 16'd6738, 16'd41135, 16'd40229, 16'd8130, 16'd26997, 16'd57744, 16'd19167, 16'd51172, 16'd38139});
	test_expansion(128'h198bcaae7cdba5740935f3dde0699c6c, {16'd19777, 16'd48092, 16'd24557, 16'd20483, 16'd35636, 16'd47606, 16'd4146, 16'd1261, 16'd20071, 16'd17168, 16'd7100, 16'd44770, 16'd50179, 16'd37702, 16'd46973, 16'd33231, 16'd35676, 16'd4232, 16'd3762, 16'd44280, 16'd30524, 16'd36529, 16'd17801, 16'd32293, 16'd1936, 16'd45000});
	test_expansion(128'h4247d01f861debf3c92c47cd402c0c68, {16'd58210, 16'd60553, 16'd34245, 16'd11452, 16'd31651, 16'd46917, 16'd34847, 16'd47652, 16'd38615, 16'd35541, 16'd2951, 16'd1007, 16'd13999, 16'd38964, 16'd8210, 16'd45977, 16'd26498, 16'd46644, 16'd23592, 16'd17930, 16'd31938, 16'd62131, 16'd8140, 16'd31219, 16'd212, 16'd52898});
	test_expansion(128'h822acd1bac50c7f931b02d9f1ebeafee, {16'd39049, 16'd62458, 16'd45916, 16'd33651, 16'd50094, 16'd13334, 16'd37969, 16'd54923, 16'd43485, 16'd35973, 16'd52416, 16'd52045, 16'd15046, 16'd12110, 16'd16643, 16'd5029, 16'd9301, 16'd58363, 16'd56743, 16'd50591, 16'd28469, 16'd62724, 16'd12109, 16'd47518, 16'd62753, 16'd49303});
	test_expansion(128'h174a985fc313ff3ed283e0b6fb3b839a, {16'd27930, 16'd27753, 16'd11994, 16'd7215, 16'd9929, 16'd54106, 16'd54528, 16'd6589, 16'd4800, 16'd58814, 16'd43187, 16'd42218, 16'd61931, 16'd19805, 16'd34171, 16'd2086, 16'd14595, 16'd3745, 16'd35191, 16'd6303, 16'd61162, 16'd65273, 16'd31872, 16'd63173, 16'd27072, 16'd55617});
	test_expansion(128'h3ed04805a94ac5f5c41ac650d5a37dee, {16'd17600, 16'd55969, 16'd11914, 16'd8393, 16'd34140, 16'd64690, 16'd29640, 16'd56164, 16'd33149, 16'd15287, 16'd46742, 16'd32391, 16'd40867, 16'd12705, 16'd9003, 16'd6857, 16'd52149, 16'd23924, 16'd11142, 16'd57958, 16'd59139, 16'd63474, 16'd21139, 16'd37344, 16'd36396, 16'd12189});
	test_expansion(128'hef2aa4182a2c648d0e09dc8d24678740, {16'd24793, 16'd14942, 16'd53165, 16'd47882, 16'd19643, 16'd62224, 16'd55336, 16'd46343, 16'd42003, 16'd28291, 16'd41104, 16'd31077, 16'd52142, 16'd22013, 16'd58429, 16'd27754, 16'd61722, 16'd25906, 16'd22804, 16'd47232, 16'd26078, 16'd48332, 16'd62452, 16'd59537, 16'd43383, 16'd54587});
	test_expansion(128'h987d383c59316c5a441eacb68f2783f1, {16'd43225, 16'd10762, 16'd42436, 16'd25728, 16'd37272, 16'd32689, 16'd59053, 16'd3159, 16'd43625, 16'd17188, 16'd27093, 16'd5999, 16'd63583, 16'd65024, 16'd36727, 16'd9852, 16'd48389, 16'd14558, 16'd39619, 16'd38769, 16'd20255, 16'd33284, 16'd54440, 16'd8264, 16'd44035, 16'd19058});
	test_expansion(128'hac5a3fb76727b796b4a419df43168241, {16'd15359, 16'd46411, 16'd20572, 16'd35705, 16'd60838, 16'd299, 16'd29941, 16'd37289, 16'd12567, 16'd49322, 16'd6004, 16'd6941, 16'd25457, 16'd36353, 16'd57473, 16'd29809, 16'd8473, 16'd53346, 16'd47232, 16'd64614, 16'd17318, 16'd24458, 16'd45574, 16'd36800, 16'd27426, 16'd2597});
	test_expansion(128'hd8a4bf283abbd917cb5e7edc539a3e24, {16'd54007, 16'd52405, 16'd3180, 16'd52794, 16'd24757, 16'd8134, 16'd9136, 16'd46052, 16'd40890, 16'd15153, 16'd30174, 16'd59570, 16'd24351, 16'd27291, 16'd34776, 16'd4196, 16'd42684, 16'd562, 16'd7966, 16'd29866, 16'd45559, 16'd39959, 16'd16024, 16'd24942, 16'd51908, 16'd52054});
	test_expansion(128'h8a1b8647cd58db001190774aa7641f62, {16'd41763, 16'd60192, 16'd20919, 16'd4555, 16'd45493, 16'd52817, 16'd42176, 16'd44860, 16'd45265, 16'd57667, 16'd15164, 16'd27213, 16'd43549, 16'd13333, 16'd38169, 16'd49234, 16'd28149, 16'd51817, 16'd45866, 16'd3233, 16'd57834, 16'd33347, 16'd48387, 16'd25059, 16'd6328, 16'd7468});
	test_expansion(128'hf19afa7d722f8fc7d2264e4be5c79583, {16'd14679, 16'd12917, 16'd7531, 16'd34961, 16'd38961, 16'd51817, 16'd41698, 16'd58083, 16'd14817, 16'd40569, 16'd42528, 16'd63938, 16'd19188, 16'd26245, 16'd58576, 16'd20594, 16'd23563, 16'd13682, 16'd37902, 16'd46047, 16'd41807, 16'd40733, 16'd21933, 16'd60345, 16'd11250, 16'd20277});
	test_expansion(128'h8ce99df457583332b8437936e8d56958, {16'd48088, 16'd14549, 16'd51426, 16'd58267, 16'd56061, 16'd47226, 16'd58437, 16'd40340, 16'd62880, 16'd21291, 16'd46578, 16'd48219, 16'd35061, 16'd57423, 16'd39620, 16'd58380, 16'd31392, 16'd12671, 16'd36091, 16'd22361, 16'd25097, 16'd54890, 16'd19626, 16'd12936, 16'd50471, 16'd50165});
	test_expansion(128'h6b2a28815b3563569a0cd23aad0e36ee, {16'd13699, 16'd16437, 16'd40893, 16'd39154, 16'd20328, 16'd21346, 16'd22711, 16'd52656, 16'd7979, 16'd14592, 16'd31950, 16'd12901, 16'd50453, 16'd55412, 16'd6606, 16'd43414, 16'd35149, 16'd62383, 16'd43862, 16'd39400, 16'd35754, 16'd20269, 16'd40050, 16'd13587, 16'd21173, 16'd15937});
	test_expansion(128'h8e79fd09b88ee3157760d827e91bbf39, {16'd42592, 16'd32159, 16'd36764, 16'd22378, 16'd53563, 16'd64243, 16'd29489, 16'd12799, 16'd49243, 16'd21124, 16'd42272, 16'd46316, 16'd43054, 16'd7274, 16'd10104, 16'd18928, 16'd15821, 16'd12784, 16'd43927, 16'd33227, 16'd32092, 16'd46200, 16'd53143, 16'd27759, 16'd65130, 16'd40384});
	test_expansion(128'hc3acfe5d19784b095c4de5cb4442dd5a, {16'd36596, 16'd8729, 16'd9138, 16'd22800, 16'd42548, 16'd53597, 16'd58655, 16'd27512, 16'd61985, 16'd54129, 16'd58074, 16'd26006, 16'd10871, 16'd32509, 16'd57242, 16'd46007, 16'd22553, 16'd3907, 16'd51659, 16'd20726, 16'd34669, 16'd9563, 16'd18505, 16'd417, 16'd59566, 16'd60600});
	test_expansion(128'h4fa10c5d352b7aa8576c93597cb6ced8, {16'd9928, 16'd26509, 16'd59729, 16'd31664, 16'd20202, 16'd43263, 16'd6642, 16'd1946, 16'd16918, 16'd64002, 16'd30774, 16'd451, 16'd6979, 16'd47563, 16'd9721, 16'd27075, 16'd855, 16'd20968, 16'd60842, 16'd55807, 16'd46344, 16'd54549, 16'd20670, 16'd23843, 16'd63320, 16'd27250});
	test_expansion(128'he09f047288b293ef53697699fd4bcba3, {16'd54143, 16'd55205, 16'd26587, 16'd27384, 16'd48351, 16'd25415, 16'd4197, 16'd40488, 16'd2966, 16'd2352, 16'd35410, 16'd43132, 16'd42809, 16'd3272, 16'd20556, 16'd60704, 16'd843, 16'd21960, 16'd13158, 16'd47232, 16'd7893, 16'd2930, 16'd15442, 16'd33007, 16'd3966, 16'd59269});
	test_expansion(128'h7abf37ddd3072a90da38dc8921a410e6, {16'd56459, 16'd58538, 16'd14302, 16'd10806, 16'd56619, 16'd24158, 16'd51081, 16'd4833, 16'd10639, 16'd54259, 16'd59388, 16'd51876, 16'd35077, 16'd57855, 16'd62537, 16'd32746, 16'd28012, 16'd49278, 16'd23560, 16'd38231, 16'd20417, 16'd56121, 16'd9700, 16'd16303, 16'd61851, 16'd25967});
	test_expansion(128'he2dc0f943b064eeba4e751f1cd0aa077, {16'd59368, 16'd25646, 16'd16063, 16'd51581, 16'd2810, 16'd55420, 16'd27432, 16'd30871, 16'd23492, 16'd20435, 16'd52283, 16'd22509, 16'd53852, 16'd41020, 16'd9914, 16'd18272, 16'd47797, 16'd60164, 16'd40236, 16'd8875, 16'd55047, 16'd27101, 16'd63714, 16'd40531, 16'd44124, 16'd11215});
	test_expansion(128'hcd12003b218fde9674525b4b482e2305, {16'd17499, 16'd41848, 16'd25315, 16'd50482, 16'd28447, 16'd16639, 16'd14196, 16'd412, 16'd12098, 16'd55172, 16'd44897, 16'd47068, 16'd14990, 16'd13945, 16'd64720, 16'd33104, 16'd47584, 16'd54527, 16'd61189, 16'd23251, 16'd57984, 16'd41132, 16'd45045, 16'd20100, 16'd55102, 16'd10271});
	test_expansion(128'h968629594c9645f54595fd1e076a7d63, {16'd11525, 16'd44001, 16'd32666, 16'd25578, 16'd8990, 16'd11212, 16'd42024, 16'd8888, 16'd29109, 16'd33634, 16'd60888, 16'd28598, 16'd61036, 16'd37939, 16'd38007, 16'd39819, 16'd33194, 16'd27489, 16'd27423, 16'd27182, 16'd53065, 16'd63492, 16'd34069, 16'd8036, 16'd48303, 16'd56128});
	test_expansion(128'h41d453d4759d1380145ecc7ca210e156, {16'd378, 16'd37488, 16'd30858, 16'd29934, 16'd28080, 16'd37887, 16'd40422, 16'd11039, 16'd50946, 16'd35834, 16'd8902, 16'd6184, 16'd54064, 16'd22930, 16'd9563, 16'd42167, 16'd49639, 16'd19139, 16'd47960, 16'd12410, 16'd44863, 16'd14394, 16'd35641, 16'd3933, 16'd44570, 16'd20846});
	test_expansion(128'h163f4f9c13624e5b420692f27166c263, {16'd38894, 16'd40923, 16'd61505, 16'd13519, 16'd34001, 16'd414, 16'd25207, 16'd6179, 16'd62562, 16'd1434, 16'd11012, 16'd60510, 16'd13119, 16'd186, 16'd49760, 16'd34406, 16'd39536, 16'd16256, 16'd32256, 16'd25286, 16'd48300, 16'd49945, 16'd53043, 16'd5939, 16'd39293, 16'd40417});
	test_expansion(128'h94fac1f51eb6acf10f2965e11f03c299, {16'd49511, 16'd28135, 16'd1489, 16'd51950, 16'd63196, 16'd64450, 16'd60938, 16'd36940, 16'd64901, 16'd22223, 16'd11080, 16'd49438, 16'd16175, 16'd38646, 16'd51713, 16'd40960, 16'd22081, 16'd8004, 16'd3743, 16'd43497, 16'd4731, 16'd30599, 16'd27572, 16'd21482, 16'd15483, 16'd8277});
	test_expansion(128'h22d03dce3c89fff09d04615b514490d2, {16'd45142, 16'd26281, 16'd13818, 16'd11214, 16'd36758, 16'd65497, 16'd2821, 16'd32170, 16'd58603, 16'd58701, 16'd58622, 16'd54050, 16'd17173, 16'd22860, 16'd51182, 16'd15163, 16'd59606, 16'd46364, 16'd45966, 16'd33132, 16'd41282, 16'd4405, 16'd34186, 16'd49380, 16'd31859, 16'd62460});
	test_expansion(128'h0ca88d6ceaadd18f1830d070197b1837, {16'd62166, 16'd54894, 16'd20448, 16'd54740, 16'd38584, 16'd8015, 16'd54531, 16'd55174, 16'd53716, 16'd13716, 16'd34762, 16'd64402, 16'd20231, 16'd5394, 16'd31091, 16'd61462, 16'd10129, 16'd22651, 16'd35053, 16'd40484, 16'd50054, 16'd20771, 16'd33355, 16'd30659, 16'd30450, 16'd29677});
	test_expansion(128'hf0ddcc27ac23f8cc5aeb4ea6f7a241c1, {16'd50245, 16'd18292, 16'd56443, 16'd36256, 16'd21695, 16'd14907, 16'd39141, 16'd9941, 16'd35200, 16'd11273, 16'd42825, 16'd22781, 16'd50626, 16'd27762, 16'd59156, 16'd54703, 16'd51107, 16'd843, 16'd34244, 16'd58878, 16'd34030, 16'd21436, 16'd49329, 16'd54983, 16'd47430, 16'd46570});
	test_expansion(128'hdf8b70fcdfe20d686d07385e32ac53f6, {16'd18727, 16'd16922, 16'd23115, 16'd35121, 16'd32028, 16'd37307, 16'd50912, 16'd13378, 16'd7693, 16'd62874, 16'd5706, 16'd6349, 16'd305, 16'd28573, 16'd9620, 16'd11071, 16'd17326, 16'd5690, 16'd52129, 16'd45245, 16'd32929, 16'd19362, 16'd42661, 16'd56784, 16'd36149, 16'd14287});
	test_expansion(128'h6e0e614be3bb5212e6e1998f09374fc3, {16'd27761, 16'd26478, 16'd63037, 16'd11193, 16'd7680, 16'd1090, 16'd13702, 16'd6390, 16'd7688, 16'd6297, 16'd3990, 16'd45658, 16'd39824, 16'd32038, 16'd32678, 16'd15199, 16'd25186, 16'd26716, 16'd32670, 16'd59291, 16'd3691, 16'd30928, 16'd64212, 16'd2833, 16'd36256, 16'd10348});
	test_expansion(128'h436a417fca863bb6d4f6192cb98fac87, {16'd36276, 16'd29104, 16'd24319, 16'd14561, 16'd1610, 16'd50570, 16'd681, 16'd44086, 16'd64228, 16'd42671, 16'd65145, 16'd17746, 16'd60346, 16'd46414, 16'd55577, 16'd27304, 16'd26442, 16'd3996, 16'd47725, 16'd5589, 16'd15820, 16'd55531, 16'd39850, 16'd2457, 16'd2562, 16'd10849});
	test_expansion(128'hfe1ab1f8b07669dc987ae91bdfb68910, {16'd24721, 16'd38174, 16'd17799, 16'd2774, 16'd33219, 16'd60305, 16'd27347, 16'd56882, 16'd50131, 16'd43194, 16'd45111, 16'd15761, 16'd15645, 16'd42628, 16'd47375, 16'd20166, 16'd7620, 16'd62348, 16'd18557, 16'd38386, 16'd58503, 16'd58659, 16'd14332, 16'd17318, 16'd33649, 16'd38888});
	test_expansion(128'hab6de2707b64c2178c264f7ac44285b2, {16'd27199, 16'd40518, 16'd39408, 16'd10955, 16'd31397, 16'd37912, 16'd26850, 16'd11268, 16'd65269, 16'd17932, 16'd9426, 16'd52223, 16'd56955, 16'd63218, 16'd19893, 16'd60092, 16'd33411, 16'd16808, 16'd49149, 16'd40536, 16'd23033, 16'd64580, 16'd22299, 16'd12153, 16'd51029, 16'd15236});
	test_expansion(128'h0e02e0786098ae58af25aac23fec999e, {16'd48909, 16'd25122, 16'd41179, 16'd62308, 16'd22634, 16'd26226, 16'd38163, 16'd36574, 16'd56901, 16'd17227, 16'd7565, 16'd36655, 16'd16035, 16'd12149, 16'd49795, 16'd36250, 16'd38137, 16'd20708, 16'd8524, 16'd41063, 16'd58218, 16'd11213, 16'd60201, 16'd7229, 16'd61051, 16'd30469});
	test_expansion(128'h595d74df45c0d8bdf0f0b08fa8502168, {16'd32515, 16'd11808, 16'd48679, 16'd29052, 16'd42188, 16'd51242, 16'd11924, 16'd32235, 16'd45551, 16'd21997, 16'd11671, 16'd6056, 16'd34913, 16'd20867, 16'd25306, 16'd36463, 16'd61651, 16'd11243, 16'd61580, 16'd18236, 16'd4831, 16'd45135, 16'd16076, 16'd37664, 16'd19231, 16'd49082});
	test_expansion(128'hb54a5103a12b968db2194645f5c291ad, {16'd50595, 16'd1594, 16'd52057, 16'd20097, 16'd42573, 16'd5955, 16'd43830, 16'd10988, 16'd54132, 16'd10524, 16'd4239, 16'd46981, 16'd22950, 16'd8413, 16'd43433, 16'd15693, 16'd25813, 16'd29884, 16'd62619, 16'd49968, 16'd14025, 16'd20695, 16'd45104, 16'd18468, 16'd57386, 16'd2399});
	test_expansion(128'hbae4ee2168c1c4ad33c6f828626329d8, {16'd17526, 16'd16950, 16'd600, 16'd20632, 16'd2631, 16'd58350, 16'd18154, 16'd11185, 16'd1176, 16'd4058, 16'd62398, 16'd8790, 16'd17152, 16'd38106, 16'd31017, 16'd26390, 16'd54529, 16'd4180, 16'd59424, 16'd23283, 16'd26873, 16'd37439, 16'd2692, 16'd23516, 16'd31211, 16'd20802});
	test_expansion(128'h059788ffaf05ae356bb3cd293c35658e, {16'd20545, 16'd63688, 16'd63465, 16'd10634, 16'd19742, 16'd65054, 16'd64841, 16'd5187, 16'd56505, 16'd15030, 16'd7649, 16'd10821, 16'd27723, 16'd9967, 16'd36686, 16'd47076, 16'd30236, 16'd33906, 16'd20547, 16'd56536, 16'd6680, 16'd57115, 16'd1819, 16'd16869, 16'd3640, 16'd49581});
	test_expansion(128'hfcde3112554cb294d55f465539ffa2c4, {16'd53610, 16'd22524, 16'd39856, 16'd8462, 16'd23714, 16'd16027, 16'd50694, 16'd27302, 16'd25947, 16'd28994, 16'd29807, 16'd43257, 16'd63709, 16'd58899, 16'd40718, 16'd64038, 16'd17989, 16'd38397, 16'd34265, 16'd26609, 16'd63284, 16'd60180, 16'd3968, 16'd46111, 16'd16163, 16'd20026});
	test_expansion(128'h1afcad078aaa658c32719ec4eff81ade, {16'd62210, 16'd32847, 16'd7784, 16'd42448, 16'd23273, 16'd33108, 16'd12593, 16'd47698, 16'd18013, 16'd27263, 16'd12098, 16'd60186, 16'd7385, 16'd48809, 16'd12570, 16'd17257, 16'd11129, 16'd28075, 16'd3924, 16'd15799, 16'd6884, 16'd57490, 16'd21427, 16'd20002, 16'd14903, 16'd63366});
	test_expansion(128'hc48d3111121dac1d94af19a849b30dda, {16'd55480, 16'd60585, 16'd34362, 16'd57197, 16'd55515, 16'd22538, 16'd36887, 16'd30534, 16'd32529, 16'd47009, 16'd17956, 16'd56685, 16'd1648, 16'd62920, 16'd63965, 16'd12354, 16'd60478, 16'd52277, 16'd43779, 16'd42801, 16'd12652, 16'd51674, 16'd47115, 16'd17743, 16'd20360, 16'd8477});
	test_expansion(128'h8aac7ff9e2a63ef2a3652ed63748395b, {16'd41193, 16'd33728, 16'd11171, 16'd33672, 16'd27553, 16'd53009, 16'd32456, 16'd42428, 16'd32777, 16'd61898, 16'd43047, 16'd24870, 16'd44764, 16'd45891, 16'd4152, 16'd41651, 16'd1392, 16'd30096, 16'd33480, 16'd53181, 16'd40337, 16'd65357, 16'd59161, 16'd54750, 16'd17411, 16'd10573});
	test_expansion(128'he8a55f899161fa51629e71b01dea953f, {16'd60572, 16'd14451, 16'd42741, 16'd42102, 16'd49012, 16'd65534, 16'd30695, 16'd11179, 16'd7520, 16'd212, 16'd33209, 16'd42533, 16'd28539, 16'd6681, 16'd23921, 16'd8098, 16'd38283, 16'd9413, 16'd52714, 16'd39797, 16'd63334, 16'd7515, 16'd45549, 16'd61301, 16'd10830, 16'd63263});
	test_expansion(128'hfb0cda3e6a34b196bbea9818892617d4, {16'd46754, 16'd44201, 16'd3269, 16'd2863, 16'd9456, 16'd62993, 16'd6654, 16'd14740, 16'd64738, 16'd60515, 16'd30916, 16'd50472, 16'd24538, 16'd2646, 16'd50288, 16'd10431, 16'd39397, 16'd39631, 16'd63731, 16'd6742, 16'd16709, 16'd31171, 16'd60019, 16'd7482, 16'd50718, 16'd34847});
	test_expansion(128'h2026f59e126b3ab84b00e715674cdf3b, {16'd14341, 16'd5607, 16'd5354, 16'd48746, 16'd53363, 16'd49919, 16'd57021, 16'd31484, 16'd7661, 16'd37031, 16'd16088, 16'd12285, 16'd2419, 16'd36145, 16'd48433, 16'd47152, 16'd51963, 16'd25775, 16'd242, 16'd20604, 16'd55139, 16'd48111, 16'd24543, 16'd11964, 16'd13790, 16'd39174});
	test_expansion(128'hbc496c9683b29599cb9b777602fc96b3, {16'd45539, 16'd31829, 16'd37872, 16'd41615, 16'd14074, 16'd42140, 16'd64763, 16'd48834, 16'd38440, 16'd9039, 16'd33320, 16'd31450, 16'd57751, 16'd64990, 16'd59281, 16'd12887, 16'd55526, 16'd9617, 16'd3665, 16'd15984, 16'd19267, 16'd8665, 16'd55492, 16'd45678, 16'd60177, 16'd15289});
	test_expansion(128'h46b83a0562abdd53a100e2cce5ce50af, {16'd10580, 16'd60653, 16'd49439, 16'd27481, 16'd4379, 16'd51750, 16'd12381, 16'd56763, 16'd38798, 16'd608, 16'd20532, 16'd54495, 16'd12066, 16'd184, 16'd62976, 16'd55013, 16'd36000, 16'd6250, 16'd2538, 16'd38899, 16'd64289, 16'd35274, 16'd2977, 16'd31210, 16'd42662, 16'd55389});
	test_expansion(128'h2e9cd960a9c2860611a087693d67bf6a, {16'd65077, 16'd24609, 16'd12960, 16'd10602, 16'd49164, 16'd8962, 16'd58546, 16'd8486, 16'd19796, 16'd14697, 16'd39860, 16'd26262, 16'd12249, 16'd10202, 16'd41774, 16'd49772, 16'd18506, 16'd1288, 16'd58473, 16'd12343, 16'd58604, 16'd31771, 16'd56353, 16'd40312, 16'd63436, 16'd48598});
	test_expansion(128'h07f8b1fe3a6dda74009ca632d9626961, {16'd26642, 16'd55595, 16'd38636, 16'd8925, 16'd51880, 16'd50382, 16'd51965, 16'd55676, 16'd14458, 16'd37793, 16'd51482, 16'd30678, 16'd18390, 16'd56728, 16'd11779, 16'd36303, 16'd35387, 16'd53761, 16'd9743, 16'd29290, 16'd37639, 16'd48578, 16'd38800, 16'd3920, 16'd9428, 16'd1088});
	test_expansion(128'h7e6a770ca43af47ed53774284320a55c, {16'd46917, 16'd61926, 16'd20976, 16'd49088, 16'd11405, 16'd57764, 16'd8067, 16'd11242, 16'd9996, 16'd58158, 16'd10310, 16'd63904, 16'd55352, 16'd24768, 16'd27472, 16'd32645, 16'd55239, 16'd27742, 16'd50243, 16'd1309, 16'd12885, 16'd1733, 16'd7730, 16'd8357, 16'd47538, 16'd15107});
	test_expansion(128'h0029f9b74b39ea96008ce5c430c0f609, {16'd52504, 16'd30758, 16'd19792, 16'd12863, 16'd56909, 16'd44101, 16'd58441, 16'd518, 16'd61808, 16'd59928, 16'd58001, 16'd3436, 16'd19366, 16'd30628, 16'd27363, 16'd2432, 16'd57400, 16'd55938, 16'd64659, 16'd31202, 16'd13639, 16'd39971, 16'd45998, 16'd55287, 16'd52686, 16'd8846});
	test_expansion(128'hfd7ec537e2ef343c09f81dd4467f56a9, {16'd28392, 16'd44101, 16'd60909, 16'd32826, 16'd37592, 16'd64393, 16'd30712, 16'd6445, 16'd39116, 16'd50532, 16'd37076, 16'd26200, 16'd47888, 16'd50702, 16'd22539, 16'd29541, 16'd37615, 16'd47385, 16'd24234, 16'd54111, 16'd10602, 16'd41761, 16'd28749, 16'd23693, 16'd27460, 16'd45599});
	test_expansion(128'hac5c4c911a182cf5f0403192d0bd4287, {16'd56010, 16'd1906, 16'd48524, 16'd21626, 16'd15055, 16'd6386, 16'd12825, 16'd17239, 16'd41362, 16'd25571, 16'd3653, 16'd41938, 16'd52848, 16'd44827, 16'd57553, 16'd50453, 16'd65269, 16'd2524, 16'd54768, 16'd39241, 16'd8861, 16'd21828, 16'd59398, 16'd59403, 16'd8337, 16'd61790});
	test_expansion(128'h81453a30bdb12510bdbb7cff114de271, {16'd49329, 16'd47833, 16'd10887, 16'd60404, 16'd8062, 16'd15113, 16'd34739, 16'd65457, 16'd1381, 16'd47587, 16'd42159, 16'd8743, 16'd47777, 16'd17454, 16'd43566, 16'd20269, 16'd62850, 16'd7993, 16'd47454, 16'd12142, 16'd35919, 16'd51157, 16'd10, 16'd27246, 16'd61344, 16'd60027});
	test_expansion(128'h1c0b94b367b5ba7e0161e6076447c586, {16'd55034, 16'd9953, 16'd58828, 16'd55198, 16'd20077, 16'd19031, 16'd17917, 16'd50922, 16'd26120, 16'd16062, 16'd58907, 16'd35035, 16'd40481, 16'd25657, 16'd58573, 16'd3160, 16'd22349, 16'd44828, 16'd16887, 16'd54339, 16'd51692, 16'd19890, 16'd52, 16'd31488, 16'd20060, 16'd32331});
	test_expansion(128'h001deb89d288b75473573a1d5cda09bf, {16'd9982, 16'd15709, 16'd61221, 16'd9222, 16'd25400, 16'd15274, 16'd36723, 16'd65345, 16'd27120, 16'd9190, 16'd48361, 16'd56862, 16'd13506, 16'd94, 16'd56619, 16'd31130, 16'd50415, 16'd25720, 16'd7049, 16'd18955, 16'd16360, 16'd42297, 16'd6842, 16'd61051, 16'd53850, 16'd15419});
	test_expansion(128'h1d915ef4d7ae156a6fefc0ca4e4c5f8d, {16'd56954, 16'd12427, 16'd11324, 16'd4944, 16'd27118, 16'd37895, 16'd19607, 16'd57849, 16'd17063, 16'd34821, 16'd6523, 16'd27882, 16'd64134, 16'd51717, 16'd12115, 16'd16735, 16'd55209, 16'd27072, 16'd26712, 16'd28936, 16'd42886, 16'd1564, 16'd25562, 16'd47581, 16'd23727, 16'd34134});
	test_expansion(128'h0614573770088471f64bacb1209babe3, {16'd3859, 16'd33360, 16'd28293, 16'd30179, 16'd16063, 16'd26032, 16'd65403, 16'd15119, 16'd37602, 16'd14453, 16'd51007, 16'd51553, 16'd30614, 16'd23085, 16'd10943, 16'd37143, 16'd39695, 16'd60154, 16'd53701, 16'd35239, 16'd49302, 16'd18701, 16'd2963, 16'd5435, 16'd59506, 16'd8875});
	test_expansion(128'h428394f6e0c08ee34e2fec914e6d59db, {16'd12313, 16'd49381, 16'd37335, 16'd45891, 16'd41746, 16'd19845, 16'd5522, 16'd41297, 16'd16700, 16'd56908, 16'd3787, 16'd33610, 16'd61783, 16'd38519, 16'd42604, 16'd59661, 16'd16585, 16'd63849, 16'd14788, 16'd51253, 16'd63300, 16'd52906, 16'd34300, 16'd18532, 16'd54380, 16'd65353});
	test_expansion(128'h12fbed524b7328d11a1ee0db99ca467d, {16'd44769, 16'd26453, 16'd1922, 16'd35063, 16'd121, 16'd38583, 16'd36894, 16'd18336, 16'd9828, 16'd15805, 16'd35294, 16'd29936, 16'd15532, 16'd49, 16'd15778, 16'd28486, 16'd6020, 16'd51233, 16'd62893, 16'd39016, 16'd13664, 16'd55955, 16'd60957, 16'd40192, 16'd35197, 16'd22783});
	test_expansion(128'h63a247e1553bba91b02b5c0f024e34b6, {16'd61991, 16'd63334, 16'd62426, 16'd62264, 16'd53612, 16'd23453, 16'd33117, 16'd60908, 16'd21607, 16'd9913, 16'd61473, 16'd25492, 16'd7315, 16'd15569, 16'd49826, 16'd214, 16'd61603, 16'd57981, 16'd11497, 16'd22682, 16'd18042, 16'd44010, 16'd8592, 16'd54515, 16'd7471, 16'd38394});
	test_expansion(128'h400a541e018c6095719defac395bee2a, {16'd36088, 16'd5504, 16'd26667, 16'd62455, 16'd1109, 16'd35702, 16'd17276, 16'd45573, 16'd50199, 16'd50903, 16'd47196, 16'd65139, 16'd13290, 16'd21598, 16'd2653, 16'd25892, 16'd27688, 16'd28984, 16'd26742, 16'd50223, 16'd26931, 16'd33111, 16'd27036, 16'd5922, 16'd21193, 16'd4427});
	test_expansion(128'hd54afeebeab15865f6ad5feabf91930d, {16'd77, 16'd27659, 16'd12976, 16'd8723, 16'd2207, 16'd23841, 16'd46387, 16'd7656, 16'd61430, 16'd37893, 16'd45117, 16'd58640, 16'd31462, 16'd9602, 16'd3213, 16'd51902, 16'd36280, 16'd56390, 16'd8479, 16'd61740, 16'd4420, 16'd21934, 16'd16599, 16'd17989, 16'd13650, 16'd51103});
	test_expansion(128'hcddd9e125ce29d74aaf2fd031cf9e10f, {16'd64703, 16'd65479, 16'd5245, 16'd49821, 16'd33696, 16'd11076, 16'd22325, 16'd45258, 16'd25286, 16'd47270, 16'd63238, 16'd58046, 16'd2472, 16'd38840, 16'd39299, 16'd61718, 16'd17468, 16'd1592, 16'd27719, 16'd49314, 16'd48157, 16'd53492, 16'd64451, 16'd13057, 16'd20570, 16'd25969});
	test_expansion(128'h29bb5067e708a0e189d61cc47a55f8f7, {16'd57618, 16'd40567, 16'd32794, 16'd6856, 16'd8536, 16'd43681, 16'd19993, 16'd28136, 16'd10527, 16'd48965, 16'd4688, 16'd47528, 16'd46315, 16'd14367, 16'd43247, 16'd34853, 16'd59168, 16'd65187, 16'd28737, 16'd12446, 16'd50630, 16'd21173, 16'd31593, 16'd6566, 16'd28224, 16'd8613});
	test_expansion(128'h68348ddac1a758f477d4e1778b699c60, {16'd33043, 16'd18547, 16'd24806, 16'd46282, 16'd52676, 16'd7645, 16'd62433, 16'd57575, 16'd48428, 16'd16453, 16'd1018, 16'd3482, 16'd12454, 16'd17554, 16'd45, 16'd42468, 16'd41097, 16'd16091, 16'd44780, 16'd4827, 16'd28899, 16'd23882, 16'd49339, 16'd11833, 16'd53889, 16'd24326});
	test_expansion(128'h857964fb6d05e739554a0201980a5a25, {16'd12698, 16'd57721, 16'd38587, 16'd33655, 16'd31183, 16'd24920, 16'd49627, 16'd15279, 16'd9772, 16'd2085, 16'd3577, 16'd11928, 16'd42650, 16'd13406, 16'd8987, 16'd63691, 16'd28070, 16'd46333, 16'd61868, 16'd55657, 16'd8507, 16'd49043, 16'd18342, 16'd41572, 16'd65294, 16'd64798});
	test_expansion(128'h97f72a81a246a7e83f61f8af431045e9, {16'd55661, 16'd16225, 16'd41191, 16'd40493, 16'd8061, 16'd19429, 16'd32893, 16'd28634, 16'd31507, 16'd54077, 16'd40467, 16'd12341, 16'd44989, 16'd50734, 16'd21705, 16'd4076, 16'd26604, 16'd26304, 16'd2319, 16'd20391, 16'd5776, 16'd23889, 16'd33350, 16'd47229, 16'd61855, 16'd8671});
	test_expansion(128'h84023fda44a7298ae61306407cffbe18, {16'd40835, 16'd37778, 16'd25749, 16'd21972, 16'd25943, 16'd54058, 16'd33385, 16'd24266, 16'd12989, 16'd26658, 16'd6716, 16'd35989, 16'd29326, 16'd54575, 16'd56624, 16'd3922, 16'd53205, 16'd28161, 16'd4713, 16'd56070, 16'd15515, 16'd46452, 16'd44433, 16'd1432, 16'd39335, 16'd22940});
	test_expansion(128'hb253fc4f13baecf006600e794f813cdd, {16'd22414, 16'd39892, 16'd32574, 16'd31284, 16'd30984, 16'd21556, 16'd11043, 16'd30109, 16'd16369, 16'd52253, 16'd21818, 16'd25275, 16'd49008, 16'd46335, 16'd6070, 16'd20518, 16'd31867, 16'd14254, 16'd49826, 16'd56501, 16'd4943, 16'd62769, 16'd62859, 16'd42574, 16'd33457, 16'd23001});
	test_expansion(128'h1c4e8eb5b472de7a35901c5c49dcd383, {16'd22493, 16'd47537, 16'd4884, 16'd62182, 16'd49367, 16'd14817, 16'd42147, 16'd11572, 16'd2474, 16'd61236, 16'd32320, 16'd63040, 16'd13838, 16'd56322, 16'd35404, 16'd54209, 16'd40657, 16'd13389, 16'd37839, 16'd27611, 16'd40733, 16'd39006, 16'd41788, 16'd20169, 16'd43432, 16'd60388});
	test_expansion(128'h4114ee588ef3c5ec4680a432a0274ac1, {16'd54831, 16'd42615, 16'd36603, 16'd32109, 16'd45734, 16'd26981, 16'd60277, 16'd16655, 16'd9098, 16'd10163, 16'd28043, 16'd8241, 16'd63285, 16'd24051, 16'd49329, 16'd21892, 16'd8925, 16'd28764, 16'd9226, 16'd39105, 16'd29014, 16'd56161, 16'd17780, 16'd63817, 16'd8522, 16'd26352});
	test_expansion(128'h966a2365cd1d683a444f437af00813fd, {16'd59647, 16'd41600, 16'd37948, 16'd62503, 16'd53299, 16'd18315, 16'd23911, 16'd5494, 16'd42347, 16'd34561, 16'd10332, 16'd55974, 16'd31880, 16'd19901, 16'd9689, 16'd38111, 16'd15597, 16'd33541, 16'd17286, 16'd34543, 16'd43543, 16'd23653, 16'd1219, 16'd49160, 16'd64024, 16'd43028});
	test_expansion(128'hb7d4cf67c9f430ed654d513ffd29f7d5, {16'd27036, 16'd51184, 16'd32, 16'd53050, 16'd17162, 16'd23517, 16'd2078, 16'd61929, 16'd39578, 16'd12495, 16'd32806, 16'd53092, 16'd44131, 16'd7931, 16'd62483, 16'd52463, 16'd43321, 16'd10012, 16'd56140, 16'd1609, 16'd29448, 16'd9175, 16'd64790, 16'd13304, 16'd38742, 16'd62763});
	test_expansion(128'h1bcea1484d065234b4614a31515d381b, {16'd54959, 16'd41883, 16'd34043, 16'd35032, 16'd23014, 16'd9636, 16'd6887, 16'd5576, 16'd13657, 16'd35307, 16'd22875, 16'd29043, 16'd32698, 16'd15428, 16'd64661, 16'd41713, 16'd56002, 16'd17862, 16'd43960, 16'd32480, 16'd35619, 16'd36190, 16'd50669, 16'd62076, 16'd34421, 16'd34591});
	test_expansion(128'hc01f52598f5a1d3ba92ae6c837c19aa2, {16'd3956, 16'd32634, 16'd31102, 16'd46610, 16'd7929, 16'd1504, 16'd35219, 16'd43634, 16'd49118, 16'd30107, 16'd22720, 16'd25433, 16'd20434, 16'd4282, 16'd57626, 16'd34240, 16'd44295, 16'd44771, 16'd13132, 16'd22128, 16'd45880, 16'd13940, 16'd24934, 16'd22869, 16'd24926, 16'd41626});
	test_expansion(128'h71e923d7c2d1cb6f5bcff093a12e9a81, {16'd16322, 16'd51950, 16'd37850, 16'd6220, 16'd2499, 16'd31491, 16'd5980, 16'd18, 16'd47732, 16'd18027, 16'd57918, 16'd4537, 16'd56725, 16'd12795, 16'd61926, 16'd34824, 16'd15701, 16'd37644, 16'd47299, 16'd52179, 16'd1627, 16'd34865, 16'd28424, 16'd29738, 16'd24374, 16'd1723});
	test_expansion(128'h11b213d937cafa2cc3542328cf3345ff, {16'd54614, 16'd24795, 16'd40171, 16'd28873, 16'd54140, 16'd58403, 16'd25326, 16'd23358, 16'd54632, 16'd4035, 16'd2429, 16'd10089, 16'd18167, 16'd23811, 16'd56918, 16'd16454, 16'd6195, 16'd42652, 16'd21389, 16'd61868, 16'd62344, 16'd44903, 16'd7323, 16'd4616, 16'd56565, 16'd13035});
	test_expansion(128'ha071e30bdeb04525e9c73f2bba88c4d1, {16'd15899, 16'd38892, 16'd41582, 16'd14921, 16'd57600, 16'd18888, 16'd30166, 16'd58537, 16'd2302, 16'd58664, 16'd63846, 16'd30641, 16'd54647, 16'd13204, 16'd11760, 16'd35499, 16'd37105, 16'd24288, 16'd39100, 16'd64311, 16'd51730, 16'd26958, 16'd30664, 16'd45109, 16'd37625, 16'd64010});
	test_expansion(128'hb09578008a2227f93b74a99188b899b2, {16'd40473, 16'd14318, 16'd58018, 16'd59589, 16'd15359, 16'd59621, 16'd51658, 16'd2878, 16'd16199, 16'd8153, 16'd55396, 16'd16928, 16'd20559, 16'd9376, 16'd24292, 16'd18954, 16'd46256, 16'd11068, 16'd53422, 16'd43128, 16'd737, 16'd63239, 16'd46266, 16'd16639, 16'd53795, 16'd25000});
	test_expansion(128'h47f029e3ede35bf8f4b282ef131e8321, {16'd20392, 16'd19836, 16'd46454, 16'd34660, 16'd41710, 16'd32794, 16'd19839, 16'd18726, 16'd49157, 16'd57950, 16'd28539, 16'd38550, 16'd48646, 16'd27654, 16'd30931, 16'd47679, 16'd24896, 16'd58039, 16'd28525, 16'd34657, 16'd30988, 16'd35368, 16'd17703, 16'd515, 16'd53260, 16'd3872});
	test_expansion(128'h392fadaaafac1484909a702ac6c26e38, {16'd16611, 16'd38282, 16'd40316, 16'd39334, 16'd29094, 16'd7169, 16'd23398, 16'd25414, 16'd16848, 16'd48440, 16'd25761, 16'd60424, 16'd28852, 16'd39143, 16'd25932, 16'd60909, 16'd3658, 16'd13039, 16'd63051, 16'd42388, 16'd36257, 16'd46366, 16'd24593, 16'd33764, 16'd7234, 16'd33940});
	test_expansion(128'h9544d919e44148d2d55e0f115e7772ad, {16'd41230, 16'd5866, 16'd33366, 16'd30, 16'd39846, 16'd54894, 16'd63046, 16'd11865, 16'd6227, 16'd38684, 16'd3705, 16'd23901, 16'd32063, 16'd52702, 16'd53440, 16'd61247, 16'd40573, 16'd54940, 16'd1211, 16'd21031, 16'd6439, 16'd59442, 16'd10960, 16'd41066, 16'd16987, 16'd19015});
	test_expansion(128'h20128bed17e7a89e7f248870f80106c3, {16'd17023, 16'd27925, 16'd16092, 16'd63245, 16'd48377, 16'd43965, 16'd54256, 16'd65006, 16'd37599, 16'd39911, 16'd29911, 16'd44278, 16'd56155, 16'd19454, 16'd62220, 16'd58558, 16'd59671, 16'd22508, 16'd5747, 16'd56974, 16'd4163, 16'd51341, 16'd28102, 16'd6784, 16'd61111, 16'd59419});
	test_expansion(128'hdb2c7ff342d6ee13948860fc8248492b, {16'd58738, 16'd27731, 16'd43296, 16'd34244, 16'd41873, 16'd56425, 16'd8119, 16'd12416, 16'd48239, 16'd44655, 16'd38979, 16'd24090, 16'd43138, 16'd49938, 16'd35071, 16'd1001, 16'd45106, 16'd2170, 16'd55197, 16'd10708, 16'd9303, 16'd29813, 16'd18026, 16'd53290, 16'd7645, 16'd26168});
	test_expansion(128'h3c5c39f30643f68cd9de61ebd058acc3, {16'd60538, 16'd54780, 16'd17458, 16'd55307, 16'd54971, 16'd4333, 16'd5848, 16'd35696, 16'd27648, 16'd40133, 16'd22837, 16'd29656, 16'd46823, 16'd26280, 16'd40889, 16'd58876, 16'd45991, 16'd4678, 16'd41730, 16'd25072, 16'd79, 16'd4743, 16'd14825, 16'd56015, 16'd50118, 16'd38780});
	test_expansion(128'haf6c4d38a12f43f5435939b0a52774a5, {16'd10323, 16'd52399, 16'd7848, 16'd44866, 16'd32231, 16'd36664, 16'd12700, 16'd11974, 16'd2231, 16'd1780, 16'd15052, 16'd58153, 16'd7889, 16'd46857, 16'd8896, 16'd497, 16'd23131, 16'd54931, 16'd46949, 16'd12777, 16'd9832, 16'd32394, 16'd57518, 16'd16338, 16'd1548, 16'd26420});
	test_expansion(128'h2003e8436aeb6d9bee6febb38b45f14d, {16'd48100, 16'd50690, 16'd37183, 16'd64976, 16'd38034, 16'd27717, 16'd10410, 16'd26037, 16'd56571, 16'd65161, 16'd50360, 16'd31767, 16'd21041, 16'd1843, 16'd17189, 16'd39993, 16'd60634, 16'd50551, 16'd26508, 16'd33776, 16'd33103, 16'd32392, 16'd24631, 16'd54050, 16'd876, 16'd42329});
	test_expansion(128'h960213323ee1f17253b7574ab7f27e3d, {16'd31630, 16'd30702, 16'd13359, 16'd3360, 16'd14111, 16'd49478, 16'd3476, 16'd62484, 16'd59159, 16'd29692, 16'd4799, 16'd48718, 16'd17657, 16'd43649, 16'd43062, 16'd62512, 16'd22919, 16'd29030, 16'd46843, 16'd54582, 16'd43781, 16'd23103, 16'd50568, 16'd36464, 16'd62032, 16'd55876});
	test_expansion(128'h353826f92aae7d10466c5c022c0bd6a1, {16'd5959, 16'd4915, 16'd46213, 16'd3240, 16'd43363, 16'd20811, 16'd6508, 16'd45339, 16'd62552, 16'd39117, 16'd37751, 16'd4127, 16'd63618, 16'd53320, 16'd25691, 16'd42382, 16'd37619, 16'd48313, 16'd30892, 16'd26397, 16'd60118, 16'd6308, 16'd24849, 16'd59571, 16'd12326, 16'd55828});
	test_expansion(128'hb7949b285dc51b3a64be336c1fc1703c, {16'd49373, 16'd16214, 16'd19713, 16'd44210, 16'd38207, 16'd12052, 16'd39682, 16'd59153, 16'd56573, 16'd48360, 16'd3828, 16'd30353, 16'd11601, 16'd20177, 16'd34870, 16'd55874, 16'd64727, 16'd1136, 16'd16760, 16'd6830, 16'd42242, 16'd50064, 16'd42643, 16'd33362, 16'd1239, 16'd3255});
	test_expansion(128'h1186f559f2ac138353de5585f7512a84, {16'd23646, 16'd53120, 16'd41530, 16'd60930, 16'd55733, 16'd20456, 16'd40059, 16'd59080, 16'd56502, 16'd3593, 16'd53320, 16'd18380, 16'd49263, 16'd42897, 16'd33525, 16'd43464, 16'd38989, 16'd34985, 16'd48062, 16'd54172, 16'd28493, 16'd13394, 16'd42908, 16'd25916, 16'd2149, 16'd61450});
	test_expansion(128'hae78c47f0fa6e3fae6ba1e6b7fd88a20, {16'd7748, 16'd36267, 16'd52960, 16'd56854, 16'd24820, 16'd22122, 16'd14194, 16'd10327, 16'd64642, 16'd59950, 16'd33561, 16'd20208, 16'd29395, 16'd18386, 16'd25694, 16'd33830, 16'd11885, 16'd41276, 16'd19850, 16'd21174, 16'd61978, 16'd43041, 16'd55146, 16'd37574, 16'd53150, 16'd10052});
	test_expansion(128'ha36632dd84aa05a46c20334b7f09d76e, {16'd51988, 16'd52683, 16'd31857, 16'd55535, 16'd675, 16'd45780, 16'd50392, 16'd18136, 16'd32560, 16'd50648, 16'd60682, 16'd47040, 16'd45033, 16'd34076, 16'd24824, 16'd23987, 16'd22576, 16'd22853, 16'd35178, 16'd19596, 16'd5467, 16'd11432, 16'd34977, 16'd6998, 16'd1349, 16'd28614});
	test_expansion(128'h1b2eb4c98bb7f6117f590aa62209d6ce, {16'd59370, 16'd31828, 16'd8683, 16'd44880, 16'd53222, 16'd24838, 16'd22341, 16'd58372, 16'd31806, 16'd16071, 16'd1776, 16'd52568, 16'd5134, 16'd63375, 16'd35974, 16'd28494, 16'd11533, 16'd38242, 16'd36974, 16'd38953, 16'd37699, 16'd43110, 16'd35917, 16'd46233, 16'd64543, 16'd60918});
	test_expansion(128'h80cd562c48aa2c1c0fb30510c5d94e9b, {16'd56795, 16'd41607, 16'd26992, 16'd47300, 16'd64964, 16'd24208, 16'd16896, 16'd39523, 16'd22199, 16'd28020, 16'd53093, 16'd16322, 16'd18604, 16'd51851, 16'd25351, 16'd3309, 16'd44258, 16'd10413, 16'd26539, 16'd25999, 16'd43500, 16'd21102, 16'd26713, 16'd1790, 16'd58493, 16'd59758});
	test_expansion(128'h12d550b60ec921fcda0f1a01c349793c, {16'd63828, 16'd20790, 16'd45362, 16'd40684, 16'd53355, 16'd32319, 16'd18801, 16'd57761, 16'd31531, 16'd8990, 16'd34626, 16'd45266, 16'd50149, 16'd26349, 16'd33186, 16'd47887, 16'd47796, 16'd17718, 16'd57742, 16'd9903, 16'd63240, 16'd41792, 16'd7932, 16'd18264, 16'd51208, 16'd4297});
	test_expansion(128'hdef0d2a4770b469b015c05db0e8987b6, {16'd8482, 16'd10322, 16'd35432, 16'd8369, 16'd4536, 16'd42546, 16'd33076, 16'd63545, 16'd14020, 16'd20103, 16'd45846, 16'd43621, 16'd56883, 16'd45558, 16'd1622, 16'd2826, 16'd55898, 16'd63852, 16'd23801, 16'd62733, 16'd6649, 16'd43113, 16'd64459, 16'd11833, 16'd15974, 16'd31769});
	test_expansion(128'h7a905c0285bfbb91884ae9145d9fd8a8, {16'd47809, 16'd48739, 16'd49848, 16'd24088, 16'd54657, 16'd59872, 16'd43048, 16'd7454, 16'd51267, 16'd49208, 16'd58573, 16'd58312, 16'd10462, 16'd1475, 16'd3920, 16'd53876, 16'd60343, 16'd63829, 16'd12459, 16'd48092, 16'd51504, 16'd51849, 16'd64016, 16'd22620, 16'd63011, 16'd56099});
	test_expansion(128'h64dc885130778fb80064bdae17201d86, {16'd24173, 16'd23627, 16'd43009, 16'd24860, 16'd40423, 16'd48123, 16'd7034, 16'd55182, 16'd60793, 16'd2855, 16'd27557, 16'd10894, 16'd29267, 16'd24769, 16'd50354, 16'd38116, 16'd5267, 16'd48340, 16'd50658, 16'd10727, 16'd43709, 16'd30162, 16'd54534, 16'd44652, 16'd6083, 16'd30264});
	test_expansion(128'hbaca77fa297b341c66e48a0f98367bea, {16'd21407, 16'd18116, 16'd36790, 16'd63363, 16'd28504, 16'd44136, 16'd18069, 16'd36131, 16'd59646, 16'd63491, 16'd25706, 16'd61823, 16'd49634, 16'd44868, 16'd13846, 16'd52509, 16'd40773, 16'd24452, 16'd51234, 16'd54544, 16'd57318, 16'd26107, 16'd45775, 16'd7887, 16'd57905, 16'd10701});
	test_expansion(128'h5c20c9e18532ef322c7aaeb77d003b92, {16'd59736, 16'd48937, 16'd36820, 16'd14805, 16'd16226, 16'd3816, 16'd37506, 16'd8869, 16'd28514, 16'd9044, 16'd40780, 16'd22267, 16'd64810, 16'd42525, 16'd34931, 16'd50385, 16'd59712, 16'd11363, 16'd8923, 16'd43275, 16'd37154, 16'd11474, 16'd26628, 16'd62463, 16'd62609, 16'd26734});
	test_expansion(128'hd892589a81bc2ae84971a125168ee9bf, {16'd39757, 16'd38509, 16'd64791, 16'd41209, 16'd48330, 16'd843, 16'd7062, 16'd59654, 16'd60626, 16'd4343, 16'd36602, 16'd27112, 16'd61880, 16'd60884, 16'd334, 16'd3972, 16'd51209, 16'd11400, 16'd59756, 16'd50735, 16'd19707, 16'd23088, 16'd57062, 16'd4132, 16'd50687, 16'd59339});
	test_expansion(128'ha1629979394fd7f9db9042078e91e747, {16'd63173, 16'd50116, 16'd27296, 16'd600, 16'd59956, 16'd56429, 16'd46217, 16'd14563, 16'd43108, 16'd63622, 16'd63290, 16'd26762, 16'd29495, 16'd53076, 16'd24965, 16'd18871, 16'd57187, 16'd45704, 16'd26805, 16'd32571, 16'd16938, 16'd1873, 16'd57790, 16'd9057, 16'd11917, 16'd3280});
	test_expansion(128'h877edd29e28b22aca6a7bf22523b5ab2, {16'd49618, 16'd20447, 16'd9776, 16'd8935, 16'd10464, 16'd51294, 16'd60764, 16'd56914, 16'd1993, 16'd59043, 16'd61988, 16'd13565, 16'd64690, 16'd36615, 16'd45644, 16'd7623, 16'd48597, 16'd12112, 16'd58712, 16'd6621, 16'd49412, 16'd7395, 16'd12150, 16'd4189, 16'd24145, 16'd13303});
	test_expansion(128'hd72295b392c1c897400f4beccd4ac2b6, {16'd45429, 16'd46890, 16'd12276, 16'd11499, 16'd46222, 16'd53654, 16'd49517, 16'd5050, 16'd31263, 16'd20078, 16'd18507, 16'd20245, 16'd25718, 16'd37086, 16'd34309, 16'd4987, 16'd44196, 16'd8286, 16'd61527, 16'd57607, 16'd54658, 16'd17834, 16'd48156, 16'd41166, 16'd35699, 16'd1357});
	test_expansion(128'hea50f547f0a15d0e02f0e76188e13eeb, {16'd50399, 16'd9966, 16'd28036, 16'd32348, 16'd24504, 16'd45505, 16'd33756, 16'd31962, 16'd20694, 16'd15637, 16'd28388, 16'd64899, 16'd259, 16'd23332, 16'd29176, 16'd41230, 16'd39807, 16'd28502, 16'd44043, 16'd42920, 16'd13972, 16'd9671, 16'd43440, 16'd51164, 16'd670, 16'd33669});
	test_expansion(128'h55d6b74b1b5cc3b1eaf6195d97dd5b3e, {16'd38610, 16'd45166, 16'd10652, 16'd4395, 16'd2738, 16'd62047, 16'd44857, 16'd43723, 16'd25424, 16'd35404, 16'd15240, 16'd29856, 16'd47080, 16'd6048, 16'd17111, 16'd25059, 16'd44388, 16'd34430, 16'd35027, 16'd18864, 16'd7202, 16'd10476, 16'd12693, 16'd63818, 16'd11730, 16'd22606});
	test_expansion(128'hce7ff8a4bd72b22db1d3efc9cd103bcd, {16'd46073, 16'd49096, 16'd7001, 16'd41845, 16'd58592, 16'd52534, 16'd3815, 16'd4504, 16'd13976, 16'd53563, 16'd3594, 16'd6200, 16'd10645, 16'd43873, 16'd34647, 16'd49179, 16'd26566, 16'd33049, 16'd47171, 16'd17044, 16'd50778, 16'd17500, 16'd55801, 16'd47479, 16'd25067, 16'd16148});
	test_expansion(128'h886661f0e3ebed1510dd355df79b02a8, {16'd6829, 16'd54026, 16'd50005, 16'd7011, 16'd16361, 16'd24935, 16'd25188, 16'd16674, 16'd26103, 16'd24066, 16'd19436, 16'd65290, 16'd53684, 16'd10238, 16'd62191, 16'd27857, 16'd54643, 16'd40134, 16'd32199, 16'd27078, 16'd38028, 16'd39616, 16'd25942, 16'd14779, 16'd25627, 16'd28081});
	test_expansion(128'he7a0b2e276f68fd5d2180f3ded5ee766, {16'd29294, 16'd56655, 16'd35327, 16'd57160, 16'd39212, 16'd3729, 16'd51593, 16'd5567, 16'd21390, 16'd58502, 16'd6351, 16'd64564, 16'd7073, 16'd45391, 16'd22707, 16'd26182, 16'd61778, 16'd34812, 16'd56198, 16'd32796, 16'd39313, 16'd52606, 16'd58157, 16'd34840, 16'd19503, 16'd50918});
	test_expansion(128'h1b64bac343e4873ceb2b8be0024154bb, {16'd25480, 16'd46019, 16'd41380, 16'd26573, 16'd31737, 16'd10386, 16'd23920, 16'd33410, 16'd20320, 16'd24448, 16'd52880, 16'd27578, 16'd16317, 16'd29771, 16'd40611, 16'd53320, 16'd58397, 16'd34633, 16'd61182, 16'd34360, 16'd5964, 16'd48864, 16'd19287, 16'd49091, 16'd12200, 16'd38989});
	test_expansion(128'h86acd352b32fe0d7d173081877944e0d, {16'd49112, 16'd5170, 16'd36001, 16'd1842, 16'd61944, 16'd65288, 16'd61517, 16'd27161, 16'd1904, 16'd12240, 16'd5242, 16'd27022, 16'd64581, 16'd36999, 16'd10715, 16'd31796, 16'd27271, 16'd35281, 16'd47682, 16'd43295, 16'd44720, 16'd56156, 16'd62257, 16'd63298, 16'd59728, 16'd27315});
	test_expansion(128'h35eb6d2d331c8638609d271c919eea20, {16'd873, 16'd29571, 16'd19461, 16'd7910, 16'd47042, 16'd7980, 16'd56850, 16'd54561, 16'd15400, 16'd31277, 16'd27258, 16'd14810, 16'd5614, 16'd41759, 16'd35711, 16'd50013, 16'd63922, 16'd11505, 16'd60742, 16'd33016, 16'd7708, 16'd56088, 16'd21851, 16'd9605, 16'd63429, 16'd60559});
	test_expansion(128'ha57b9e9d32337d7348b864269879c85d, {16'd30149, 16'd2692, 16'd9271, 16'd41039, 16'd30720, 16'd974, 16'd14332, 16'd52395, 16'd45267, 16'd58582, 16'd61928, 16'd5313, 16'd18991, 16'd41592, 16'd44560, 16'd1417, 16'd33981, 16'd63862, 16'd36318, 16'd63503, 16'd43436, 16'd20052, 16'd22370, 16'd57216, 16'd54134, 16'd59193});
	test_expansion(128'hd53c5fe15c8038569ac3b672529e5d9f, {16'd3167, 16'd45622, 16'd60185, 16'd43546, 16'd6418, 16'd28912, 16'd59347, 16'd45494, 16'd2763, 16'd29995, 16'd13957, 16'd12294, 16'd27929, 16'd40044, 16'd6857, 16'd36783, 16'd55690, 16'd25388, 16'd64162, 16'd26309, 16'd18462, 16'd16343, 16'd45126, 16'd38514, 16'd30633, 16'd19299});
	test_expansion(128'h0110180b4e43926ee005e30ae323b0d1, {16'd45584, 16'd241, 16'd8060, 16'd20713, 16'd21486, 16'd8017, 16'd57034, 16'd2932, 16'd33988, 16'd23965, 16'd30093, 16'd46750, 16'd1891, 16'd23568, 16'd48840, 16'd756, 16'd17835, 16'd37777, 16'd36410, 16'd28957, 16'd2881, 16'd25620, 16'd47388, 16'd49641, 16'd42702, 16'd34186});
	test_expansion(128'h58715f5a148ba6a12e206442d8b5b165, {16'd4839, 16'd54009, 16'd56569, 16'd50535, 16'd63538, 16'd2790, 16'd38872, 16'd17364, 16'd33075, 16'd31400, 16'd40327, 16'd3626, 16'd16523, 16'd46765, 16'd24094, 16'd56580, 16'd53846, 16'd34216, 16'd7809, 16'd57667, 16'd60553, 16'd23434, 16'd8876, 16'd8966, 16'd14952, 16'd39525});
	test_expansion(128'h8f6a1c02056b6b269eb0c88cd0d77d58, {16'd23878, 16'd47338, 16'd46448, 16'd36488, 16'd59467, 16'd45449, 16'd33380, 16'd30374, 16'd13177, 16'd54384, 16'd58649, 16'd27956, 16'd43157, 16'd1903, 16'd5123, 16'd59007, 16'd50960, 16'd24014, 16'd40297, 16'd36254, 16'd17212, 16'd19136, 16'd1712, 16'd59445, 16'd5589, 16'd45867});
	test_expansion(128'ha9a35a72cbf9cc62ebada13b049dccc9, {16'd62902, 16'd52957, 16'd5206, 16'd59133, 16'd65168, 16'd5931, 16'd42589, 16'd46144, 16'd20667, 16'd11628, 16'd13148, 16'd4633, 16'd24782, 16'd48992, 16'd15930, 16'd2868, 16'd28975, 16'd24492, 16'd9331, 16'd53400, 16'd6231, 16'd10297, 16'd30913, 16'd37432, 16'd7632, 16'd15687});
	test_expansion(128'h0892cbf58011d6e486c73f913daad49e, {16'd22300, 16'd23516, 16'd39348, 16'd22845, 16'd30471, 16'd52820, 16'd26226, 16'd3568, 16'd43060, 16'd53830, 16'd32566, 16'd53163, 16'd23234, 16'd2433, 16'd22786, 16'd52235, 16'd6105, 16'd4457, 16'd7664, 16'd50498, 16'd63489, 16'd9830, 16'd12566, 16'd21526, 16'd3380, 16'd50023});
	test_expansion(128'he40ad3d5df7dfa7804b3adfafa79711c, {16'd41889, 16'd41725, 16'd32624, 16'd46054, 16'd63816, 16'd1821, 16'd47755, 16'd42616, 16'd18413, 16'd43439, 16'd37103, 16'd41553, 16'd20933, 16'd18279, 16'd53259, 16'd59752, 16'd9590, 16'd63930, 16'd58093, 16'd42799, 16'd36377, 16'd49149, 16'd48128, 16'd47186, 16'd10022, 16'd43230});
	test_expansion(128'h670ccbb49ee460a8f7d3b40b8adfde4d, {16'd11270, 16'd1499, 16'd2316, 16'd24948, 16'd28887, 16'd25850, 16'd7461, 16'd51216, 16'd17111, 16'd62761, 16'd1750, 16'd8514, 16'd40475, 16'd58611, 16'd26250, 16'd62295, 16'd46506, 16'd54397, 16'd7859, 16'd45713, 16'd39960, 16'd12590, 16'd57890, 16'd48670, 16'd51575, 16'd43225});
	test_expansion(128'he7107f7838e2ae5f37cf0efe92b50a1c, {16'd20463, 16'd48516, 16'd56346, 16'd56463, 16'd34092, 16'd43116, 16'd41142, 16'd19409, 16'd52738, 16'd54526, 16'd17177, 16'd46261, 16'd10733, 16'd767, 16'd43543, 16'd53905, 16'd59495, 16'd51191, 16'd19473, 16'd26467, 16'd2266, 16'd10298, 16'd4282, 16'd16867, 16'd36555, 16'd4899});
	test_expansion(128'hc373caf8eebfbaa8cfbba55324984c55, {16'd57287, 16'd14949, 16'd61140, 16'd58470, 16'd33694, 16'd38054, 16'd4247, 16'd63808, 16'd61556, 16'd47768, 16'd57654, 16'd8233, 16'd25742, 16'd21553, 16'd62954, 16'd49743, 16'd30508, 16'd49338, 16'd23213, 16'd4890, 16'd26786, 16'd59684, 16'd7537, 16'd34463, 16'd45309, 16'd20588});
	test_expansion(128'he7d1590b1380a839ba001fe2cf156769, {16'd62596, 16'd56127, 16'd41599, 16'd17445, 16'd958, 16'd4055, 16'd43004, 16'd37318, 16'd41837, 16'd63324, 16'd26856, 16'd47521, 16'd1438, 16'd49636, 16'd62982, 16'd65453, 16'd11596, 16'd28119, 16'd20646, 16'd58295, 16'd10653, 16'd25502, 16'd29064, 16'd15745, 16'd33470, 16'd37406});
	test_expansion(128'h14a4c5bb31a3a7b64c1dddcd7f353f6d, {16'd34343, 16'd31774, 16'd30149, 16'd58540, 16'd54791, 16'd488, 16'd11220, 16'd41997, 16'd24803, 16'd40555, 16'd55468, 16'd35982, 16'd38300, 16'd63010, 16'd45833, 16'd51823, 16'd51419, 16'd13152, 16'd31075, 16'd4950, 16'd34751, 16'd51916, 16'd50239, 16'd8106, 16'd22521, 16'd8967});
	test_expansion(128'hef38522ae036e42a8c7edb36fe8492b0, {16'd46310, 16'd12007, 16'd28926, 16'd58628, 16'd56442, 16'd1716, 16'd62742, 16'd33678, 16'd25905, 16'd15430, 16'd63018, 16'd3565, 16'd34884, 16'd61428, 16'd28287, 16'd24631, 16'd62753, 16'd8472, 16'd31937, 16'd14758, 16'd16936, 16'd65514, 16'd48613, 16'd32294, 16'd61056, 16'd16170});
	test_expansion(128'h066bbe98f00677e093286e9e0af0f786, {16'd43204, 16'd34842, 16'd27828, 16'd28697, 16'd65372, 16'd58755, 16'd9601, 16'd7849, 16'd8543, 16'd20416, 16'd26662, 16'd28176, 16'd14525, 16'd25346, 16'd56262, 16'd20302, 16'd61664, 16'd53955, 16'd11022, 16'd41289, 16'd3659, 16'd25804, 16'd45477, 16'd52652, 16'd47902, 16'd42742});
	test_expansion(128'h9bf04353be07bae314edabf443b32b5b, {16'd43876, 16'd12959, 16'd36027, 16'd26036, 16'd47721, 16'd12976, 16'd49568, 16'd13166, 16'd41710, 16'd35906, 16'd32968, 16'd38650, 16'd58433, 16'd61846, 16'd52797, 16'd59261, 16'd37035, 16'd15831, 16'd19151, 16'd26433, 16'd4482, 16'd50978, 16'd28054, 16'd6297, 16'd41164, 16'd57349});
	test_expansion(128'h3fb73f4d6f3dcf0a564c6fbed69fea48, {16'd40547, 16'd48440, 16'd42381, 16'd45411, 16'd32678, 16'd34506, 16'd47589, 16'd48236, 16'd21500, 16'd38870, 16'd15059, 16'd40942, 16'd970, 16'd15218, 16'd38432, 16'd40632, 16'd49288, 16'd61667, 16'd62855, 16'd4536, 16'd23189, 16'd41284, 16'd52585, 16'd22602, 16'd3466, 16'd22614});
	test_expansion(128'h68aeefbe3098214bf55ef7a98ccc8cea, {16'd32793, 16'd15734, 16'd12789, 16'd20122, 16'd60504, 16'd21664, 16'd5498, 16'd63243, 16'd19323, 16'd48148, 16'd49461, 16'd37710, 16'd19840, 16'd53617, 16'd12228, 16'd34459, 16'd53471, 16'd33930, 16'd4660, 16'd13118, 16'd46969, 16'd60833, 16'd11051, 16'd32360, 16'd24370, 16'd29832});
	test_expansion(128'heaeebea3736257ae22b6c086144589e2, {16'd23285, 16'd57750, 16'd61876, 16'd56344, 16'd43236, 16'd7764, 16'd18816, 16'd9134, 16'd50985, 16'd63919, 16'd2584, 16'd21120, 16'd51039, 16'd32215, 16'd30172, 16'd12430, 16'd33063, 16'd43724, 16'd9193, 16'd7621, 16'd40611, 16'd5183, 16'd43669, 16'd18233, 16'd10360, 16'd32545});
	test_expansion(128'hb19f1a4ae562dfe6d0a0383ba5835ebc, {16'd24815, 16'd2336, 16'd35833, 16'd35098, 16'd47806, 16'd57361, 16'd8547, 16'd40078, 16'd18540, 16'd53797, 16'd23564, 16'd50497, 16'd4675, 16'd64014, 16'd28099, 16'd1472, 16'd3185, 16'd9678, 16'd29782, 16'd2769, 16'd53510, 16'd47093, 16'd55445, 16'd61120, 16'd26954, 16'd47425});
	test_expansion(128'h3e5f68ed9c3852a2fdafbd34533bdda9, {16'd22076, 16'd40275, 16'd12843, 16'd25175, 16'd56228, 16'd18258, 16'd39998, 16'd25098, 16'd43179, 16'd2557, 16'd15630, 16'd10256, 16'd61759, 16'd51844, 16'd37252, 16'd25975, 16'd6582, 16'd31474, 16'd26508, 16'd49932, 16'd20365, 16'd25996, 16'd35197, 16'd50763, 16'd38358, 16'd15070});
	test_expansion(128'ha05568622ff84d15e54f8b9952d23eab, {16'd25352, 16'd10115, 16'd56716, 16'd17807, 16'd31257, 16'd59736, 16'd27593, 16'd50964, 16'd55888, 16'd54760, 16'd15928, 16'd3642, 16'd32449, 16'd49567, 16'd28163, 16'd7784, 16'd45652, 16'd36028, 16'd35532, 16'd54667, 16'd38539, 16'd25676, 16'd27771, 16'd23470, 16'd30743, 16'd3541});
	test_expansion(128'h9b5bf785a6cd917a180ef5db644f68bc, {16'd32584, 16'd14539, 16'd52104, 16'd12803, 16'd64495, 16'd53490, 16'd35098, 16'd42514, 16'd38395, 16'd39487, 16'd15608, 16'd12947, 16'd14331, 16'd2018, 16'd33335, 16'd28887, 16'd27240, 16'd14896, 16'd47305, 16'd55011, 16'd44219, 16'd42623, 16'd49323, 16'd41899, 16'd57228, 16'd3315});
	test_expansion(128'hfdd2cb75129445d6963758fd1f59cf6f, {16'd39977, 16'd61652, 16'd5301, 16'd58297, 16'd11555, 16'd50867, 16'd13399, 16'd183, 16'd32897, 16'd64678, 16'd45053, 16'd26279, 16'd3142, 16'd54840, 16'd25583, 16'd47850, 16'd38165, 16'd61546, 16'd6557, 16'd10822, 16'd38705, 16'd1311, 16'd54969, 16'd39087, 16'd11756, 16'd41461});
	test_expansion(128'hd908f495ecef9488079f1794ad61108d, {16'd19837, 16'd9859, 16'd26993, 16'd53478, 16'd26880, 16'd9227, 16'd62498, 16'd56661, 16'd55635, 16'd17625, 16'd51986, 16'd41190, 16'd39606, 16'd24093, 16'd53632, 16'd4191, 16'd38430, 16'd340, 16'd15864, 16'd2022, 16'd1767, 16'd46988, 16'd47652, 16'd27088, 16'd25705, 16'd55275});
	test_expansion(128'h12dab6b4bd1d5e44b39c129ac7bb8ac1, {16'd59990, 16'd5044, 16'd57097, 16'd34349, 16'd2265, 16'd10436, 16'd24150, 16'd6024, 16'd61889, 16'd8454, 16'd20604, 16'd32983, 16'd90, 16'd9473, 16'd14103, 16'd15799, 16'd56033, 16'd46248, 16'd55292, 16'd42780, 16'd18874, 16'd45388, 16'd10261, 16'd32967, 16'd21880, 16'd17595});
	test_expansion(128'hdec397b7dc1054d2e4afce7717cd126f, {16'd64805, 16'd22002, 16'd62072, 16'd14435, 16'd55721, 16'd1725, 16'd54078, 16'd34213, 16'd62560, 16'd30318, 16'd25493, 16'd52069, 16'd3860, 16'd18849, 16'd47827, 16'd6286, 16'd10359, 16'd61329, 16'd65534, 16'd58399, 16'd37449, 16'd63672, 16'd14964, 16'd46690, 16'd32938, 16'd44490});
	test_expansion(128'hb672875e539882733c9d983b22cdad35, {16'd44906, 16'd1415, 16'd51171, 16'd64561, 16'd6427, 16'd31111, 16'd23209, 16'd32693, 16'd38154, 16'd41843, 16'd64341, 16'd42635, 16'd17391, 16'd58932, 16'd47600, 16'd64478, 16'd62466, 16'd18399, 16'd53585, 16'd54425, 16'd53511, 16'd62325, 16'd8813, 16'd57366, 16'd9706, 16'd30336});
	test_expansion(128'h52019ae06b51382a70a5518e4db8d8d2, {16'd7874, 16'd38930, 16'd59409, 16'd1415, 16'd15486, 16'd3684, 16'd40837, 16'd15488, 16'd50529, 16'd41416, 16'd8338, 16'd22555, 16'd60677, 16'd7984, 16'd17568, 16'd33620, 16'd13286, 16'd5802, 16'd57614, 16'd5498, 16'd45502, 16'd5540, 16'd4407, 16'd53043, 16'd64785, 16'd48912});
	test_expansion(128'hc6f022fa5d6e3fb69be10bf027c54219, {16'd26433, 16'd45902, 16'd14036, 16'd39820, 16'd60623, 16'd25245, 16'd57882, 16'd40615, 16'd29855, 16'd58068, 16'd61988, 16'd46706, 16'd61018, 16'd5087, 16'd24516, 16'd34830, 16'd14841, 16'd24264, 16'd49238, 16'd43272, 16'd10601, 16'd53923, 16'd3246, 16'd48456, 16'd32960, 16'd27985});
	test_expansion(128'h2bd64ffcf42935ceae9259196c9dcf71, {16'd10390, 16'd49706, 16'd38804, 16'd55382, 16'd16280, 16'd23855, 16'd35048, 16'd10640, 16'd63368, 16'd56130, 16'd57290, 16'd42336, 16'd58647, 16'd44167, 16'd25852, 16'd29571, 16'd62854, 16'd20585, 16'd29536, 16'd50229, 16'd27351, 16'd48578, 16'd1882, 16'd20411, 16'd31664, 16'd19640});
	test_expansion(128'h91b24b75dc06cd4a2c56470828ada7e5, {16'd13001, 16'd31565, 16'd12472, 16'd36154, 16'd63245, 16'd14198, 16'd6696, 16'd7299, 16'd44900, 16'd34686, 16'd51768, 16'd60206, 16'd36718, 16'd43419, 16'd37402, 16'd41799, 16'd8460, 16'd9097, 16'd41796, 16'd32228, 16'd19338, 16'd58465, 16'd1114, 16'd40651, 16'd40181, 16'd33542});
	test_expansion(128'h82af4451f0befe5b5878f09fc2abe732, {16'd57416, 16'd46842, 16'd18591, 16'd49477, 16'd31445, 16'd42337, 16'd35714, 16'd32454, 16'd53924, 16'd24370, 16'd36738, 16'd15582, 16'd16206, 16'd26406, 16'd14338, 16'd50266, 16'd45118, 16'd36680, 16'd62997, 16'd10346, 16'd26636, 16'd60969, 16'd50091, 16'd15404, 16'd26825, 16'd37020});
	test_expansion(128'h6c4d2f294a7f503dc0bbf20d3f047c7b, {16'd22666, 16'd11640, 16'd60527, 16'd51668, 16'd35714, 16'd23452, 16'd38716, 16'd2266, 16'd10514, 16'd63844, 16'd41946, 16'd48389, 16'd21309, 16'd42423, 16'd49290, 16'd58442, 16'd2818, 16'd7968, 16'd39401, 16'd13666, 16'd39562, 16'd57220, 16'd20509, 16'd51495, 16'd15479, 16'd52837});
	test_expansion(128'ha2030de5e6a4e9fc4409499c862c43d9, {16'd11455, 16'd62143, 16'd43894, 16'd3105, 16'd35719, 16'd27165, 16'd30374, 16'd57277, 16'd11310, 16'd18190, 16'd13734, 16'd14020, 16'd24888, 16'd43706, 16'd32481, 16'd16858, 16'd36838, 16'd22268, 16'd35627, 16'd60801, 16'd15549, 16'd14023, 16'd38962, 16'd36506, 16'd11790, 16'd46203});
	test_expansion(128'ha5dbae6704814cf30a9988556bd3ed7b, {16'd25632, 16'd47612, 16'd18224, 16'd5822, 16'd16092, 16'd23268, 16'd10851, 16'd49299, 16'd9720, 16'd38255, 16'd40336, 16'd14589, 16'd17309, 16'd39846, 16'd60268, 16'd51580, 16'd45268, 16'd57773, 16'd25836, 16'd60535, 16'd34757, 16'd2173, 16'd19163, 16'd53358, 16'd29753, 16'd29654});
	test_expansion(128'h393593dd3c505327f9dab2b2e6943d7b, {16'd12557, 16'd31119, 16'd59176, 16'd27292, 16'd50179, 16'd62049, 16'd55460, 16'd63432, 16'd39853, 16'd27086, 16'd34310, 16'd44680, 16'd65326, 16'd21745, 16'd11956, 16'd62476, 16'd36047, 16'd35861, 16'd35260, 16'd2514, 16'd63909, 16'd39577, 16'd1569, 16'd41777, 16'd15427, 16'd56641});
	test_expansion(128'h1959e7caca3cf94a788aa0668c38466a, {16'd3395, 16'd49103, 16'd24653, 16'd53232, 16'd30843, 16'd20625, 16'd8990, 16'd27312, 16'd65090, 16'd43737, 16'd1505, 16'd40773, 16'd15009, 16'd13430, 16'd2755, 16'd9797, 16'd62045, 16'd24004, 16'd37985, 16'd49936, 16'd59054, 16'd5699, 16'd32487, 16'd36789, 16'd60546, 16'd4403});
	test_expansion(128'h76b54fa1ac8e39aa584393ca06b8c0e0, {16'd49211, 16'd51685, 16'd55496, 16'd63838, 16'd8047, 16'd50672, 16'd8814, 16'd13945, 16'd33407, 16'd59273, 16'd4264, 16'd46084, 16'd31785, 16'd14663, 16'd20186, 16'd7843, 16'd29171, 16'd14336, 16'd56707, 16'd54245, 16'd52801, 16'd32877, 16'd64738, 16'd5530, 16'd65048, 16'd59222});
	test_expansion(128'he508304e9004a84c7e103a91cd69383b, {16'd31637, 16'd43993, 16'd34779, 16'd64910, 16'd24155, 16'd17887, 16'd50563, 16'd11884, 16'd13935, 16'd25649, 16'd38704, 16'd9166, 16'd29636, 16'd5977, 16'd29102, 16'd5096, 16'd11798, 16'd26646, 16'd58220, 16'd54140, 16'd1222, 16'd36726, 16'd30001, 16'd50419, 16'd11847, 16'd39657});
	test_expansion(128'h3e9fa32c4a5d6778c30713ee6ba51f99, {16'd54507, 16'd12001, 16'd1538, 16'd38388, 16'd9332, 16'd60884, 16'd8340, 16'd61114, 16'd25597, 16'd37049, 16'd52736, 16'd62564, 16'd26575, 16'd13095, 16'd19754, 16'd31805, 16'd41792, 16'd49870, 16'd28979, 16'd8399, 16'd44074, 16'd25533, 16'd43542, 16'd23406, 16'd41230, 16'd55126});
	test_expansion(128'h34827ca32da7102d9569627158db2cbd, {16'd37680, 16'd13119, 16'd58556, 16'd55119, 16'd26189, 16'd54966, 16'd10662, 16'd18578, 16'd57807, 16'd9214, 16'd46315, 16'd54167, 16'd27727, 16'd4541, 16'd63384, 16'd44805, 16'd13474, 16'd52615, 16'd54464, 16'd31006, 16'd57118, 16'd6888, 16'd51792, 16'd58300, 16'd26057, 16'd62332});
	test_expansion(128'h127d519a8b7cf07c702ecaa63cbdcfc8, {16'd7477, 16'd1570, 16'd20220, 16'd19206, 16'd38780, 16'd7219, 16'd21185, 16'd64485, 16'd1762, 16'd3106, 16'd13559, 16'd39994, 16'd42861, 16'd43315, 16'd41249, 16'd1679, 16'd19384, 16'd235, 16'd18966, 16'd4818, 16'd23357, 16'd45953, 16'd38490, 16'd22465, 16'd51446, 16'd5117});
	test_expansion(128'h99df517baf3502ecdde1553b37fbb276, {16'd57290, 16'd36807, 16'd43807, 16'd37553, 16'd37170, 16'd10788, 16'd4025, 16'd46932, 16'd39528, 16'd23546, 16'd50711, 16'd56218, 16'd257, 16'd11539, 16'd8508, 16'd52403, 16'd46292, 16'd40427, 16'd27359, 16'd27576, 16'd51111, 16'd44295, 16'd45657, 16'd63012, 16'd21334, 16'd26519});
	test_expansion(128'h0fcd9c4fdf9a8d57bb36af17e9e0ce58, {16'd57581, 16'd28233, 16'd55157, 16'd2113, 16'd52494, 16'd35011, 16'd46141, 16'd28817, 16'd43819, 16'd12743, 16'd7484, 16'd43904, 16'd51799, 16'd37900, 16'd39003, 16'd25608, 16'd27538, 16'd54519, 16'd21781, 16'd17588, 16'd19932, 16'd39794, 16'd5416, 16'd31069, 16'd47879, 16'd27106});
	test_expansion(128'hc65fdd8ef2825cad09a8440666cbbb60, {16'd38934, 16'd65086, 16'd5918, 16'd27161, 16'd19970, 16'd60236, 16'd16525, 16'd34477, 16'd40386, 16'd63916, 16'd10394, 16'd971, 16'd57995, 16'd22914, 16'd44069, 16'd12382, 16'd47748, 16'd49795, 16'd52580, 16'd19658, 16'd14959, 16'd33690, 16'd60704, 16'd643, 16'd8364, 16'd64443});
	test_expansion(128'h347704a46b6be3e77e5e6fe772bb02f8, {16'd34853, 16'd16617, 16'd6609, 16'd2079, 16'd36909, 16'd58546, 16'd15755, 16'd48926, 16'd3620, 16'd31508, 16'd1403, 16'd31986, 16'd47842, 16'd10105, 16'd59725, 16'd35022, 16'd24684, 16'd32902, 16'd42416, 16'd31782, 16'd27742, 16'd57643, 16'd41055, 16'd45999, 16'd23432, 16'd9149});
	test_expansion(128'h948f61da14649da92abb65996086d1b6, {16'd11379, 16'd35323, 16'd38664, 16'd33828, 16'd33933, 16'd5204, 16'd28267, 16'd46716, 16'd46412, 16'd35594, 16'd37783, 16'd12804, 16'd15064, 16'd36273, 16'd16776, 16'd14821, 16'd19763, 16'd20838, 16'd39327, 16'd17320, 16'd60936, 16'd32425, 16'd64485, 16'd6881, 16'd56106, 16'd48973});
	test_expansion(128'h3211923967a3710017fc299b58a2127b, {16'd52406, 16'd38709, 16'd42673, 16'd535, 16'd9846, 16'd49285, 16'd53277, 16'd13103, 16'd32240, 16'd23428, 16'd53194, 16'd19819, 16'd7767, 16'd34365, 16'd37600, 16'd49424, 16'd3545, 16'd5753, 16'd32744, 16'd25113, 16'd6837, 16'd33637, 16'd23509, 16'd27165, 16'd34375, 16'd24251});
	test_expansion(128'h921d2936a48ad11fe5d273129798346e, {16'd42539, 16'd61284, 16'd34039, 16'd17818, 16'd14419, 16'd18435, 16'd34330, 16'd48142, 16'd4140, 16'd36056, 16'd8628, 16'd55024, 16'd27838, 16'd41723, 16'd37779, 16'd30673, 16'd30603, 16'd3943, 16'd16717, 16'd43076, 16'd15795, 16'd43908, 16'd44679, 16'd25860, 16'd5629, 16'd63951});
	test_expansion(128'hb8e8056953c50fa9115c9db67cbd742f, {16'd55594, 16'd57729, 16'd38264, 16'd22466, 16'd15637, 16'd32731, 16'd54658, 16'd61301, 16'd55918, 16'd18057, 16'd43783, 16'd28363, 16'd17463, 16'd54637, 16'd27431, 16'd23162, 16'd53622, 16'd23876, 16'd49384, 16'd10899, 16'd24210, 16'd13744, 16'd54, 16'd44689, 16'd43739, 16'd50990});
	test_expansion(128'h3bebad16fceeb31056b713801182c2ce, {16'd1882, 16'd60215, 16'd52188, 16'd48047, 16'd33080, 16'd22062, 16'd6745, 16'd44648, 16'd27050, 16'd12821, 16'd2331, 16'd47475, 16'd45313, 16'd52082, 16'd10623, 16'd19225, 16'd49726, 16'd31298, 16'd50567, 16'd13433, 16'd31432, 16'd63270, 16'd20943, 16'd16420, 16'd42796, 16'd4154});
	test_expansion(128'h7efa6512c91745cf714ba9feee33f3ab, {16'd51030, 16'd23222, 16'd30395, 16'd36982, 16'd56543, 16'd39642, 16'd25663, 16'd63070, 16'd8475, 16'd21493, 16'd53085, 16'd8889, 16'd14542, 16'd25314, 16'd14434, 16'd2936, 16'd65000, 16'd42720, 16'd35329, 16'd48061, 16'd61373, 16'd39819, 16'd8785, 16'd21100, 16'd55425, 16'd50574});
	test_expansion(128'hfd0e58d0ff8af8f4582dfee240f8bd31, {16'd34624, 16'd61779, 16'd33339, 16'd10102, 16'd27339, 16'd57500, 16'd60670, 16'd37553, 16'd65100, 16'd37060, 16'd5956, 16'd42991, 16'd1073, 16'd10919, 16'd51594, 16'd39176, 16'd48346, 16'd8733, 16'd55632, 16'd58941, 16'd52002, 16'd27826, 16'd53323, 16'd53283, 16'd33657, 16'd26288});
	test_expansion(128'hd559e80ebd8071d6bacceee065369757, {16'd51367, 16'd43620, 16'd24384, 16'd36973, 16'd51054, 16'd31427, 16'd28162, 16'd38682, 16'd9829, 16'd57752, 16'd51615, 16'd61850, 16'd11730, 16'd48683, 16'd64824, 16'd7002, 16'd42519, 16'd40521, 16'd19369, 16'd60064, 16'd10615, 16'd30713, 16'd20555, 16'd58492, 16'd48564, 16'd24081});
	test_expansion(128'hdbef741ddff94819777467a29084676a, {16'd20270, 16'd7111, 16'd19345, 16'd65506, 16'd23804, 16'd55767, 16'd22189, 16'd57638, 16'd38741, 16'd43588, 16'd9441, 16'd39142, 16'd31172, 16'd46166, 16'd10159, 16'd52139, 16'd18109, 16'd47470, 16'd26646, 16'd44361, 16'd8633, 16'd14003, 16'd51137, 16'd16004, 16'd35926, 16'd18706});
	test_expansion(128'h26fdb6913db27634d6ea3bbd95759c23, {16'd27590, 16'd23254, 16'd19960, 16'd9005, 16'd30161, 16'd59594, 16'd22824, 16'd276, 16'd20999, 16'd11760, 16'd5569, 16'd13456, 16'd38600, 16'd43516, 16'd37252, 16'd57426, 16'd25311, 16'd34966, 16'd20408, 16'd17992, 16'd7884, 16'd2403, 16'd46177, 16'd35352, 16'd850, 16'd54928});
	test_expansion(128'h6b1636bfc68777d80b2576b7ec8747bd, {16'd47469, 16'd40983, 16'd3902, 16'd4946, 16'd33920, 16'd56931, 16'd53196, 16'd22355, 16'd36152, 16'd45587, 16'd57020, 16'd45608, 16'd25723, 16'd22106, 16'd60105, 16'd9376, 16'd63729, 16'd15153, 16'd24752, 16'd43948, 16'd29874, 16'd34778, 16'd18968, 16'd31749, 16'd26208, 16'd10736});
	test_expansion(128'h98a9566d48e68c9dbacdbf832546e2c2, {16'd47072, 16'd60205, 16'd49604, 16'd60122, 16'd5747, 16'd29286, 16'd51413, 16'd23861, 16'd64580, 16'd4487, 16'd25104, 16'd47057, 16'd25462, 16'd16311, 16'd39349, 16'd2706, 16'd41677, 16'd33560, 16'd55829, 16'd25024, 16'd1606, 16'd19588, 16'd64500, 16'd42487, 16'd31830, 16'd42576});
	test_expansion(128'had3696ca48d1ca0c7225fb04bf8ff62e, {16'd39220, 16'd23755, 16'd39788, 16'd15960, 16'd27732, 16'd17736, 16'd31363, 16'd47997, 16'd18656, 16'd2534, 16'd5341, 16'd60395, 16'd54048, 16'd43611, 16'd58934, 16'd37568, 16'd22930, 16'd21951, 16'd21399, 16'd45959, 16'd27041, 16'd62028, 16'd45323, 16'd64712, 16'd51646, 16'd41026});
	test_expansion(128'ha6ddb545f74d3c2a26f3e8c372d241b1, {16'd65435, 16'd41402, 16'd61805, 16'd50431, 16'd48573, 16'd61271, 16'd13264, 16'd25848, 16'd50134, 16'd35290, 16'd38103, 16'd43015, 16'd51359, 16'd44917, 16'd16361, 16'd28431, 16'd30809, 16'd16315, 16'd22637, 16'd59920, 16'd60614, 16'd58587, 16'd61875, 16'd7827, 16'd56117, 16'd19269});
	test_expansion(128'h4545567392b1955c6333d7c550d7cd63, {16'd9644, 16'd2596, 16'd42881, 16'd49074, 16'd35578, 16'd43743, 16'd50463, 16'd52375, 16'd58972, 16'd59652, 16'd16139, 16'd43287, 16'd12470, 16'd8757, 16'd32833, 16'd50597, 16'd21824, 16'd54459, 16'd10055, 16'd39888, 16'd1610, 16'd16355, 16'd63924, 16'd47390, 16'd62683, 16'd13789});
	test_expansion(128'h8559f2ed5e94967dce2164cf9d1e9cfe, {16'd15897, 16'd25751, 16'd50642, 16'd12099, 16'd13720, 16'd34983, 16'd867, 16'd22026, 16'd26186, 16'd45923, 16'd37306, 16'd36715, 16'd21907, 16'd63382, 16'd37770, 16'd52390, 16'd36439, 16'd61414, 16'd61209, 16'd2733, 16'd61756, 16'd30987, 16'd42049, 16'd47678, 16'd18963, 16'd14926});
	test_expansion(128'hccda4b97d8a5194cc5db08a792db24c8, {16'd17729, 16'd2805, 16'd37524, 16'd9647, 16'd36575, 16'd56861, 16'd14624, 16'd60892, 16'd33032, 16'd53724, 16'd39247, 16'd36244, 16'd11901, 16'd50628, 16'd11290, 16'd24705, 16'd46515, 16'd45253, 16'd24983, 16'd36855, 16'd2326, 16'd38716, 16'd38443, 16'd19274, 16'd34952, 16'd25393});
	test_expansion(128'h1e09bf6bbe55fce2953ba832abce0912, {16'd1658, 16'd44532, 16'd31890, 16'd16698, 16'd26412, 16'd20447, 16'd58650, 16'd42721, 16'd49737, 16'd65070, 16'd39640, 16'd34278, 16'd47097, 16'd24258, 16'd38494, 16'd51656, 16'd31845, 16'd21471, 16'd35114, 16'd16613, 16'd5428, 16'd18215, 16'd59095, 16'd9487, 16'd52947, 16'd60931});
	test_expansion(128'h5593dca0173f48860cae8bf8e407e4f4, {16'd19513, 16'd59291, 16'd13986, 16'd50019, 16'd35608, 16'd21203, 16'd7754, 16'd1477, 16'd19027, 16'd54972, 16'd18336, 16'd27092, 16'd11374, 16'd34576, 16'd63256, 16'd5979, 16'd23294, 16'd62, 16'd49230, 16'd62822, 16'd24125, 16'd37812, 16'd33820, 16'd35214, 16'd29839, 16'd24973});
	test_expansion(128'h0b58a276e2866f344ee526ad4126f831, {16'd9050, 16'd60957, 16'd48789, 16'd59520, 16'd58087, 16'd27690, 16'd38813, 16'd55006, 16'd38279, 16'd15443, 16'd51332, 16'd3921, 16'd37887, 16'd36198, 16'd51496, 16'd62870, 16'd32228, 16'd24727, 16'd59885, 16'd62900, 16'd17172, 16'd20680, 16'd39365, 16'd53103, 16'd43843, 16'd40639});
	test_expansion(128'h7f8f97f18bb8b2d4ea665dfc252047bd, {16'd55016, 16'd35136, 16'd61638, 16'd43951, 16'd55102, 16'd45613, 16'd44787, 16'd25625, 16'd21876, 16'd30358, 16'd17359, 16'd53755, 16'd51516, 16'd1168, 16'd65108, 16'd61659, 16'd23899, 16'd53541, 16'd39784, 16'd42523, 16'd62273, 16'd18613, 16'd46629, 16'd22450, 16'd34554, 16'd3461});
	test_expansion(128'h2fcfe538860afa5682e305cdded05967, {16'd32906, 16'd36467, 16'd6416, 16'd58506, 16'd44504, 16'd27291, 16'd55897, 16'd41862, 16'd28615, 16'd8706, 16'd39182, 16'd30351, 16'd15440, 16'd17011, 16'd50165, 16'd14650, 16'd64931, 16'd14897, 16'd49325, 16'd43816, 16'd39883, 16'd48004, 16'd410, 16'd9310, 16'd47240, 16'd58406});
	test_expansion(128'he55ac664d8af3474a39d90c72ebbefc5, {16'd38245, 16'd26721, 16'd6806, 16'd35898, 16'd57197, 16'd22387, 16'd64626, 16'd29935, 16'd47819, 16'd48927, 16'd32689, 16'd7958, 16'd13783, 16'd55190, 16'd61494, 16'd62201, 16'd35387, 16'd15076, 16'd64705, 16'd28929, 16'd39259, 16'd63752, 16'd17443, 16'd47693, 16'd58314, 16'd15404});
	test_expansion(128'h86ace388a3a63feb3e747c958fdfd135, {16'd30306, 16'd18781, 16'd7044, 16'd44248, 16'd49946, 16'd59166, 16'd11487, 16'd23708, 16'd25821, 16'd19234, 16'd7103, 16'd33703, 16'd65278, 16'd37446, 16'd23660, 16'd11742, 16'd60174, 16'd59593, 16'd55968, 16'd43218, 16'd35326, 16'd34611, 16'd46307, 16'd44658, 16'd29100, 16'd58767});
	test_expansion(128'hf346dcd17880b77b67575c25699882f8, {16'd20947, 16'd9671, 16'd20457, 16'd41287, 16'd63105, 16'd61903, 16'd33745, 16'd55486, 16'd56483, 16'd58977, 16'd28157, 16'd16765, 16'd36597, 16'd56530, 16'd32290, 16'd5759, 16'd26570, 16'd43198, 16'd46834, 16'd45387, 16'd39618, 16'd30298, 16'd55978, 16'd50773, 16'd27447, 16'd9453});
	test_expansion(128'h14944514de4879d9b7619057c9fbfbb6, {16'd43491, 16'd54430, 16'd54813, 16'd30969, 16'd16748, 16'd3566, 16'd45249, 16'd12383, 16'd21402, 16'd42617, 16'd59416, 16'd5871, 16'd8430, 16'd55051, 16'd63674, 16'd14083, 16'd30231, 16'd52305, 16'd52268, 16'd61047, 16'd10403, 16'd35202, 16'd27065, 16'd8775, 16'd10308, 16'd57826});
	test_expansion(128'hd783691978357d172039253a7130b1ed, {16'd11226, 16'd22248, 16'd58004, 16'd13483, 16'd37040, 16'd57348, 16'd7532, 16'd47624, 16'd30633, 16'd2003, 16'd4527, 16'd33848, 16'd39937, 16'd10182, 16'd31103, 16'd34386, 16'd22320, 16'd18020, 16'd43318, 16'd36524, 16'd28604, 16'd40546, 16'd18606, 16'd9659, 16'd55212, 16'd53646});
	test_expansion(128'h1f2c18e365850d5350431d219b10a270, {16'd19497, 16'd29253, 16'd36518, 16'd56834, 16'd50947, 16'd47225, 16'd39101, 16'd44552, 16'd60352, 16'd35550, 16'd107, 16'd35518, 16'd12283, 16'd23, 16'd40203, 16'd49092, 16'd1623, 16'd36295, 16'd23558, 16'd3516, 16'd64976, 16'd32492, 16'd7446, 16'd16747, 16'd62679, 16'd12});
	test_expansion(128'h73ee0e087374068c2567190522256eb0, {16'd9827, 16'd1781, 16'd34867, 16'd837, 16'd5469, 16'd44389, 16'd54840, 16'd41390, 16'd42689, 16'd44282, 16'd2685, 16'd18882, 16'd58572, 16'd65310, 16'd17853, 16'd23651, 16'd43340, 16'd49760, 16'd17080, 16'd61110, 16'd24821, 16'd15999, 16'd31267, 16'd19013, 16'd56692, 16'd16918});
	test_expansion(128'h15f0770d51c865e008eddcb23fa59203, {16'd41811, 16'd50071, 16'd37770, 16'd61784, 16'd60682, 16'd33808, 16'd6406, 16'd209, 16'd11772, 16'd50013, 16'd32501, 16'd8579, 16'd23008, 16'd768, 16'd31003, 16'd64401, 16'd8157, 16'd20558, 16'd57472, 16'd43286, 16'd26797, 16'd26610, 16'd65001, 16'd56748, 16'd1498, 16'd31485});
	test_expansion(128'hc85d27d4e17ea54a3f404e252701a522, {16'd18848, 16'd26249, 16'd52624, 16'd37271, 16'd16883, 16'd31727, 16'd11336, 16'd52581, 16'd53153, 16'd8134, 16'd56608, 16'd37410, 16'd61056, 16'd19868, 16'd42214, 16'd35258, 16'd41758, 16'd20146, 16'd38116, 16'd28330, 16'd52577, 16'd36558, 16'd45163, 16'd47208, 16'd2359, 16'd13219});
	test_expansion(128'hdea751ffeb549771dc00af67f468c1bf, {16'd27922, 16'd30089, 16'd14200, 16'd17636, 16'd38234, 16'd4314, 16'd61324, 16'd17319, 16'd39205, 16'd48922, 16'd39461, 16'd55440, 16'd3767, 16'd62941, 16'd32049, 16'd14082, 16'd59794, 16'd6584, 16'd38064, 16'd2336, 16'd22333, 16'd26470, 16'd21034, 16'd41829, 16'd8454, 16'd28022});
	test_expansion(128'h17f25ef10a2c5307c923d26777d84d5b, {16'd64674, 16'd3110, 16'd37836, 16'd38204, 16'd63555, 16'd26568, 16'd18999, 16'd34711, 16'd43617, 16'd22701, 16'd62483, 16'd9088, 16'd48716, 16'd57963, 16'd64590, 16'd57961, 16'd54678, 16'd26172, 16'd44668, 16'd18034, 16'd15596, 16'd32697, 16'd62203, 16'd29857, 16'd2264, 16'd39904});
	test_expansion(128'h750f277545f8973f717491fe16e62f9e, {16'd3308, 16'd25810, 16'd10516, 16'd50423, 16'd2394, 16'd59613, 16'd39898, 16'd63638, 16'd38810, 16'd55833, 16'd24480, 16'd4615, 16'd55913, 16'd17304, 16'd45036, 16'd41800, 16'd58698, 16'd18265, 16'd31652, 16'd63750, 16'd4241, 16'd52321, 16'd26942, 16'd50063, 16'd16758, 16'd55923});
	test_expansion(128'hf225f5d883ffc903d52d3a6b89ce275f, {16'd2743, 16'd40324, 16'd26177, 16'd15723, 16'd44208, 16'd30766, 16'd44303, 16'd64977, 16'd35279, 16'd26246, 16'd33570, 16'd39174, 16'd56688, 16'd51424, 16'd62610, 16'd61937, 16'd5338, 16'd14585, 16'd24602, 16'd6999, 16'd31260, 16'd62766, 16'd34669, 16'd8773, 16'd20631, 16'd9693});
	test_expansion(128'hb07e36c36fadff8a4890bac6770136e6, {16'd12071, 16'd42808, 16'd45863, 16'd51835, 16'd28372, 16'd58502, 16'd36090, 16'd3602, 16'd26608, 16'd9331, 16'd39726, 16'd14209, 16'd9814, 16'd32061, 16'd5888, 16'd21918, 16'd39726, 16'd24050, 16'd59012, 16'd39071, 16'd5674, 16'd30979, 16'd62386, 16'd19243, 16'd14820, 16'd2923});
	test_expansion(128'he025b812d76bb6e9350f53c6c589b97c, {16'd8881, 16'd52440, 16'd29066, 16'd62496, 16'd64781, 16'd61464, 16'd45216, 16'd2369, 16'd51743, 16'd3477, 16'd17425, 16'd34921, 16'd63645, 16'd30198, 16'd11176, 16'd8594, 16'd25464, 16'd12966, 16'd23145, 16'd24268, 16'd52306, 16'd47254, 16'd9500, 16'd9733, 16'd60690, 16'd29252});
	test_expansion(128'hc83b44a3c532c1aaa512666575e7ae9c, {16'd61761, 16'd3143, 16'd27212, 16'd10584, 16'd52202, 16'd4125, 16'd26906, 16'd2482, 16'd43553, 16'd22048, 16'd9609, 16'd23318, 16'd16085, 16'd39580, 16'd15905, 16'd26356, 16'd64311, 16'd60407, 16'd50240, 16'd40676, 16'd15360, 16'd1802, 16'd54045, 16'd58302, 16'd13744, 16'd20781});
	test_expansion(128'h92bdc76b830a96097528bce012f1e0df, {16'd11864, 16'd11673, 16'd3285, 16'd64277, 16'd14212, 16'd19108, 16'd50125, 16'd60140, 16'd18673, 16'd21920, 16'd65450, 16'd9828, 16'd28107, 16'd23076, 16'd50700, 16'd59394, 16'd29856, 16'd47929, 16'd61394, 16'd9568, 16'd17004, 16'd11385, 16'd7311, 16'd57455, 16'd63428, 16'd50821});
	test_expansion(128'h241948a4a023e3a873e2695c4eeb175d, {16'd60034, 16'd34534, 16'd54116, 16'd8998, 16'd56613, 16'd30697, 16'd61050, 16'd52619, 16'd18018, 16'd34890, 16'd33646, 16'd10895, 16'd54701, 16'd50920, 16'd13138, 16'd53545, 16'd23385, 16'd64341, 16'd58322, 16'd14993, 16'd5941, 16'd1882, 16'd48863, 16'd31144, 16'd38877, 16'd42962});
	test_expansion(128'he707fef90cc71aee28471ba3c725aef4, {16'd27738, 16'd24595, 16'd36319, 16'd6084, 16'd42159, 16'd48778, 16'd14386, 16'd7184, 16'd15683, 16'd21278, 16'd10369, 16'd32217, 16'd36470, 16'd32796, 16'd64144, 16'd51348, 16'd42373, 16'd28076, 16'd775, 16'd13552, 16'd31065, 16'd22125, 16'd46059, 16'd36892, 16'd27369, 16'd8936});
	test_expansion(128'h8c7ac50c10789831df734976ff0d7dfc, {16'd14345, 16'd7581, 16'd4147, 16'd9062, 16'd43587, 16'd43895, 16'd52855, 16'd64932, 16'd9403, 16'd35212, 16'd18684, 16'd65024, 16'd64223, 16'd45890, 16'd23457, 16'd16820, 16'd63254, 16'd24768, 16'd25503, 16'd2410, 16'd10562, 16'd32788, 16'd29228, 16'd4406, 16'd23538, 16'd56231});
	test_expansion(128'hfa2cd213d941c572b5c5c11182a14b8c, {16'd54768, 16'd32724, 16'd62790, 16'd62349, 16'd36955, 16'd31572, 16'd13690, 16'd1486, 16'd5578, 16'd35306, 16'd19749, 16'd24952, 16'd16124, 16'd10648, 16'd32102, 16'd20249, 16'd55369, 16'd45007, 16'd29120, 16'd57879, 16'd15863, 16'd63657, 16'd61831, 16'd26812, 16'd49315, 16'd64407});
	test_expansion(128'hb52c245103aaf8f41098791ba5422f37, {16'd35599, 16'd54617, 16'd3064, 16'd50386, 16'd32271, 16'd57281, 16'd50546, 16'd885, 16'd58406, 16'd33741, 16'd52617, 16'd51667, 16'd21338, 16'd9041, 16'd5925, 16'd36423, 16'd14941, 16'd40684, 16'd38064, 16'd35336, 16'd34128, 16'd44789, 16'd11219, 16'd41326, 16'd46623, 16'd5455});
	test_expansion(128'h2b683f6ebf2d1003e2ee3080152c39fa, {16'd64537, 16'd28628, 16'd55111, 16'd33730, 16'd28059, 16'd29401, 16'd11446, 16'd48658, 16'd58643, 16'd25263, 16'd17250, 16'd52415, 16'd43184, 16'd7003, 16'd11517, 16'd21984, 16'd49461, 16'd28525, 16'd43236, 16'd61074, 16'd23522, 16'd12307, 16'd44670, 16'd37847, 16'd18466, 16'd9137});
	test_expansion(128'h8cdfb17d42bbaf75483eb7f39495a0d7, {16'd12412, 16'd24589, 16'd34427, 16'd32786, 16'd22452, 16'd54951, 16'd50259, 16'd16219, 16'd3309, 16'd62615, 16'd20679, 16'd19389, 16'd16232, 16'd39275, 16'd52603, 16'd16361, 16'd55859, 16'd11157, 16'd30174, 16'd25790, 16'd28100, 16'd60288, 16'd30278, 16'd11865, 16'd61976, 16'd39591});
	test_expansion(128'h4c659d3ab77a82246a3a08ed7fefa976, {16'd15510, 16'd33640, 16'd45746, 16'd13417, 16'd37549, 16'd24456, 16'd30666, 16'd22359, 16'd645, 16'd61986, 16'd17198, 16'd13315, 16'd20547, 16'd57269, 16'd30866, 16'd7618, 16'd42768, 16'd41285, 16'd20209, 16'd40378, 16'd54433, 16'd54357, 16'd1219, 16'd27729, 16'd50902, 16'd38617});
	test_expansion(128'hdaf85b3fc0de77bc208438b01c01eb7a, {16'd11516, 16'd51421, 16'd44449, 16'd38585, 16'd33565, 16'd8584, 16'd55024, 16'd31703, 16'd5893, 16'd40592, 16'd62631, 16'd40708, 16'd46036, 16'd59573, 16'd29892, 16'd2518, 16'd54044, 16'd32929, 16'd55040, 16'd38593, 16'd63820, 16'd41025, 16'd55251, 16'd61591, 16'd12564, 16'd18919});
	test_expansion(128'h671a57fc391cefcb17cb733b8524c786, {16'd57773, 16'd30194, 16'd2995, 16'd60881, 16'd46820, 16'd56482, 16'd33596, 16'd42252, 16'd14491, 16'd52781, 16'd57270, 16'd25939, 16'd28359, 16'd12914, 16'd18487, 16'd56388, 16'd14832, 16'd12179, 16'd15057, 16'd17835, 16'd15297, 16'd23263, 16'd24733, 16'd34836, 16'd888, 16'd36100});
	test_expansion(128'h94a92c16f6dbacb8553d39bc34b38831, {16'd41847, 16'd61529, 16'd50776, 16'd14757, 16'd5442, 16'd46136, 16'd17042, 16'd27518, 16'd27585, 16'd14775, 16'd22705, 16'd14661, 16'd45830, 16'd1853, 16'd30035, 16'd47964, 16'd41977, 16'd62615, 16'd26555, 16'd64509, 16'd13538, 16'd34769, 16'd58307, 16'd48641, 16'd16057, 16'd35500});
	test_expansion(128'h56a0486547924a0d057b5af3dede246c, {16'd47664, 16'd4162, 16'd27480, 16'd47940, 16'd47153, 16'd51817, 16'd23470, 16'd62884, 16'd18164, 16'd46982, 16'd23855, 16'd23495, 16'd60381, 16'd49688, 16'd65108, 16'd34492, 16'd35209, 16'd323, 16'd23496, 16'd46688, 16'd57311, 16'd25549, 16'd61539, 16'd12768, 16'd22935, 16'd39932});
	test_expansion(128'h9537940182e60d575cd9eb1371dc3bce, {16'd40388, 16'd53459, 16'd17137, 16'd8001, 16'd45389, 16'd21189, 16'd59295, 16'd22999, 16'd36621, 16'd17409, 16'd43261, 16'd46387, 16'd23653, 16'd5732, 16'd54304, 16'd2431, 16'd53303, 16'd15231, 16'd38649, 16'd15365, 16'd25723, 16'd60883, 16'd44801, 16'd51705, 16'd26347, 16'd19085});
	test_expansion(128'h3e5a4c32389f7a0556e97ff03cd33d93, {16'd63734, 16'd51800, 16'd54572, 16'd51469, 16'd19810, 16'd13828, 16'd48889, 16'd29823, 16'd47178, 16'd59843, 16'd2189, 16'd51304, 16'd51414, 16'd50112, 16'd38814, 16'd25144, 16'd18190, 16'd44011, 16'd25176, 16'd12692, 16'd20923, 16'd18144, 16'd61552, 16'd43330, 16'd36488, 16'd2595});
	test_expansion(128'h6c1b41458f0e8fd536eea56661ea82fb, {16'd14911, 16'd7598, 16'd12, 16'd10599, 16'd55568, 16'd902, 16'd15766, 16'd13505, 16'd19258, 16'd35093, 16'd32031, 16'd17502, 16'd19067, 16'd16157, 16'd33488, 16'd9042, 16'd16034, 16'd41874, 16'd47613, 16'd55227, 16'd7215, 16'd32493, 16'd7325, 16'd64165, 16'd31215, 16'd34828});
	test_expansion(128'ha7634d49c62f14c1d2d059272ec04de1, {16'd59288, 16'd45541, 16'd16745, 16'd15375, 16'd7090, 16'd13124, 16'd49104, 16'd63197, 16'd20193, 16'd60543, 16'd38304, 16'd18270, 16'd12979, 16'd44473, 16'd26290, 16'd40441, 16'd14306, 16'd38516, 16'd10502, 16'd44799, 16'd24833, 16'd1674, 16'd30135, 16'd61467, 16'd13820, 16'd63544});
	test_expansion(128'h3b21dd5404c853033876a98ca6a2a964, {16'd56251, 16'd56894, 16'd35521, 16'd26728, 16'd16688, 16'd26931, 16'd6338, 16'd39903, 16'd38150, 16'd37622, 16'd37330, 16'd23844, 16'd36707, 16'd52465, 16'd29101, 16'd3841, 16'd41057, 16'd41884, 16'd61076, 16'd48823, 16'd49652, 16'd35459, 16'd31014, 16'd41734, 16'd2691, 16'd7762});
	test_expansion(128'ha63cca5ac9ab1dfc3bf458034ac3c685, {16'd29315, 16'd60225, 16'd9218, 16'd21931, 16'd11793, 16'd62592, 16'd6412, 16'd1635, 16'd15232, 16'd5237, 16'd44883, 16'd38157, 16'd16150, 16'd7936, 16'd58218, 16'd36363, 16'd39653, 16'd41508, 16'd9465, 16'd41424, 16'd41061, 16'd36472, 16'd57138, 16'd42621, 16'd63209, 16'd33462});
	test_expansion(128'hed55475eea665b9d55dc6cace9030e8f, {16'd16437, 16'd29628, 16'd33582, 16'd26536, 16'd23471, 16'd31198, 16'd32432, 16'd44933, 16'd56249, 16'd27800, 16'd53688, 16'd33676, 16'd50314, 16'd34563, 16'd16719, 16'd36523, 16'd42080, 16'd25475, 16'd53432, 16'd37726, 16'd18131, 16'd24118, 16'd3107, 16'd1700, 16'd55367, 16'd32427});
	test_expansion(128'hf0dd389fc924e0ced4343376f5b6ac1d, {16'd57374, 16'd38346, 16'd58373, 16'd20056, 16'd57356, 16'd33142, 16'd64735, 16'd22311, 16'd16239, 16'd18903, 16'd34346, 16'd27401, 16'd5772, 16'd36937, 16'd34320, 16'd23795, 16'd26334, 16'd16294, 16'd58109, 16'd7911, 16'd1230, 16'd60403, 16'd31120, 16'd27605, 16'd497, 16'd1019});
	test_expansion(128'h0f257b529dcf9afb44a9541dec255b35, {16'd47490, 16'd13143, 16'd37548, 16'd8835, 16'd62213, 16'd40648, 16'd30114, 16'd12827, 16'd4055, 16'd55033, 16'd55622, 16'd49104, 16'd12576, 16'd848, 16'd9022, 16'd1547, 16'd12257, 16'd52066, 16'd21332, 16'd57263, 16'd22365, 16'd36335, 16'd52103, 16'd150, 16'd24116, 16'd10144});
	test_expansion(128'hc8229505aa9c373c23a5231f9afddc72, {16'd51597, 16'd39608, 16'd28420, 16'd33698, 16'd8294, 16'd12988, 16'd7832, 16'd64627, 16'd64906, 16'd61072, 16'd31053, 16'd22890, 16'd35528, 16'd8109, 16'd60381, 16'd47294, 16'd488, 16'd20926, 16'd22599, 16'd38996, 16'd50305, 16'd53001, 16'd21789, 16'd17605, 16'd42691, 16'd49968});
	test_expansion(128'hb542ff33b8a6a4352821de1e0db23029, {16'd32205, 16'd21636, 16'd32032, 16'd31740, 16'd11140, 16'd47762, 16'd16118, 16'd39837, 16'd64071, 16'd24382, 16'd1821, 16'd335, 16'd3535, 16'd20009, 16'd36605, 16'd49427, 16'd1770, 16'd14552, 16'd50896, 16'd50260, 16'd43963, 16'd33254, 16'd18529, 16'd3627, 16'd8109, 16'd28620});
	test_expansion(128'h9e7ef9d2a5457a6c141671f40da62154, {16'd52049, 16'd4626, 16'd53598, 16'd6942, 16'd10690, 16'd2132, 16'd11742, 16'd50640, 16'd32855, 16'd29553, 16'd11405, 16'd47417, 16'd56575, 16'd20043, 16'd53452, 16'd45998, 16'd41314, 16'd6081, 16'd54872, 16'd48923, 16'd22866, 16'd13688, 16'd52805, 16'd8471, 16'd59405, 16'd18307});
	test_expansion(128'h079013c66b5aa99138f5d09930aaf276, {16'd50336, 16'd25850, 16'd10745, 16'd27076, 16'd13118, 16'd3026, 16'd24986, 16'd63475, 16'd37082, 16'd28422, 16'd57362, 16'd3478, 16'd20845, 16'd19111, 16'd43771, 16'd39320, 16'd41916, 16'd18768, 16'd12396, 16'd10684, 16'd65489, 16'd58940, 16'd18112, 16'd21, 16'd46326, 16'd37727});
	test_expansion(128'hac58e6e092fa81ded7ef24ad70d56f06, {16'd10316, 16'd50843, 16'd48034, 16'd28480, 16'd5196, 16'd50407, 16'd61618, 16'd30315, 16'd3001, 16'd34114, 16'd36602, 16'd52008, 16'd11988, 16'd15996, 16'd13962, 16'd34283, 16'd18873, 16'd50253, 16'd57364, 16'd63524, 16'd59826, 16'd20912, 16'd60183, 16'd23278, 16'd21103, 16'd25957});
	test_expansion(128'h3c158850a83a574500f3148a9f86a1a6, {16'd52802, 16'd45246, 16'd63147, 16'd46671, 16'd61283, 16'd65212, 16'd47386, 16'd31429, 16'd53937, 16'd57664, 16'd45267, 16'd50034, 16'd10176, 16'd29855, 16'd44476, 16'd22652, 16'd22219, 16'd28176, 16'd17601, 16'd14015, 16'd39430, 16'd26435, 16'd41338, 16'd31745, 16'd36464, 16'd44242});
	test_expansion(128'he58519a98f67dc42fc9085814f759659, {16'd52178, 16'd384, 16'd43863, 16'd37943, 16'd9124, 16'd60035, 16'd59190, 16'd41842, 16'd36228, 16'd16901, 16'd4180, 16'd6920, 16'd59106, 16'd5324, 16'd29459, 16'd56487, 16'd39583, 16'd50657, 16'd16568, 16'd23608, 16'd14064, 16'd61006, 16'd96, 16'd6379, 16'd57265, 16'd34308});
	test_expansion(128'hafb82d6b9a3f577a3eea1e08e0a32ab6, {16'd55109, 16'd31234, 16'd25092, 16'd62902, 16'd11607, 16'd43288, 16'd35247, 16'd29314, 16'd15659, 16'd13854, 16'd55644, 16'd58132, 16'd38652, 16'd54390, 16'd35473, 16'd10693, 16'd65273, 16'd15412, 16'd60980, 16'd13816, 16'd44743, 16'd911, 16'd29033, 16'd34284, 16'd41251, 16'd58558});
	test_expansion(128'h679447bd9e4bec03e9d80906468a5286, {16'd24131, 16'd28973, 16'd34726, 16'd29888, 16'd59622, 16'd15239, 16'd40133, 16'd31568, 16'd19683, 16'd54872, 16'd32564, 16'd49483, 16'd30393, 16'd42575, 16'd58116, 16'd33183, 16'd28289, 16'd64431, 16'd4828, 16'd33864, 16'd63445, 16'd7183, 16'd713, 16'd17604, 16'd39190, 16'd4655});
	test_expansion(128'hf92ced5799d8f7ec9c5b33ffc779c768, {16'd16491, 16'd13402, 16'd38353, 16'd254, 16'd10078, 16'd56220, 16'd511, 16'd42676, 16'd35449, 16'd52448, 16'd50573, 16'd6286, 16'd37699, 16'd50643, 16'd13792, 16'd55473, 16'd16316, 16'd3105, 16'd5007, 16'd47120, 16'd36129, 16'd18361, 16'd981, 16'd18374, 16'd46037, 16'd52275});
	test_expansion(128'h8fa2e9a40af50e5ce19f29345381ff78, {16'd45164, 16'd27943, 16'd40238, 16'd1147, 16'd46864, 16'd39606, 16'd33258, 16'd15004, 16'd38901, 16'd24051, 16'd50977, 16'd28137, 16'd41089, 16'd48355, 16'd57176, 16'd19920, 16'd63169, 16'd37293, 16'd52205, 16'd21736, 16'd41287, 16'd20587, 16'd6808, 16'd507, 16'd2405, 16'd45823});
	test_expansion(128'h52d70cf1b67eecf000f6a3bda65851e8, {16'd4883, 16'd16187, 16'd36014, 16'd16979, 16'd15230, 16'd18926, 16'd7970, 16'd17284, 16'd38261, 16'd22493, 16'd29166, 16'd248, 16'd59916, 16'd24166, 16'd39105, 16'd33272, 16'd11282, 16'd9764, 16'd37295, 16'd59692, 16'd59047, 16'd49163, 16'd40610, 16'd33182, 16'd16893, 16'd45435});
	test_expansion(128'h3c2f5455a1723b60b8e56d3f0748a5a0, {16'd15620, 16'd23322, 16'd40291, 16'd14380, 16'd34233, 16'd62076, 16'd30510, 16'd55195, 16'd17741, 16'd48454, 16'd35602, 16'd38758, 16'd19905, 16'd20596, 16'd27541, 16'd59214, 16'd12062, 16'd48205, 16'd62693, 16'd9829, 16'd11799, 16'd56248, 16'd51570, 16'd31725, 16'd9132, 16'd46713});
	test_expansion(128'h8205f0c1b572f312c7d7690f7c4095fc, {16'd6374, 16'd11787, 16'd39394, 16'd51358, 16'd44703, 16'd26722, 16'd37308, 16'd60262, 16'd48938, 16'd36875, 16'd874, 16'd57738, 16'd13773, 16'd27173, 16'd27969, 16'd62287, 16'd54283, 16'd8784, 16'd54644, 16'd23196, 16'd34771, 16'd8493, 16'd34496, 16'd56498, 16'd30103, 16'd19940});
	test_expansion(128'h747580ec2b7bc76d59338bd709ff2e77, {16'd58379, 16'd34802, 16'd52043, 16'd58025, 16'd53451, 16'd4735, 16'd11689, 16'd48481, 16'd5932, 16'd12762, 16'd18161, 16'd12277, 16'd30699, 16'd52002, 16'd3761, 16'd52330, 16'd46689, 16'd50906, 16'd47489, 16'd50106, 16'd63669, 16'd46207, 16'd5139, 16'd52773, 16'd38082, 16'd46811});
	test_expansion(128'hf9f80606c9b5c7ba2d5d19de8ad878e4, {16'd2325, 16'd1550, 16'd64387, 16'd40419, 16'd2394, 16'd29302, 16'd20691, 16'd21505, 16'd11110, 16'd2248, 16'd48318, 16'd519, 16'd21168, 16'd45588, 16'd27937, 16'd53432, 16'd41610, 16'd59175, 16'd57163, 16'd17693, 16'd39624, 16'd14136, 16'd31205, 16'd50810, 16'd57964, 16'd33535});
	test_expansion(128'h7767855cf2e763bea054e2ea9021b8af, {16'd30103, 16'd47929, 16'd61813, 16'd20649, 16'd18703, 16'd55448, 16'd51194, 16'd32704, 16'd21418, 16'd12272, 16'd46004, 16'd33355, 16'd50018, 16'd7924, 16'd56563, 16'd31816, 16'd45876, 16'd33593, 16'd51338, 16'd24309, 16'd32472, 16'd25594, 16'd50773, 16'd49636, 16'd8063, 16'd54110});
	test_expansion(128'hd05f39132fa3cc8e1e576e46f97e5cd3, {16'd56165, 16'd32045, 16'd48670, 16'd3925, 16'd28723, 16'd46267, 16'd1553, 16'd2795, 16'd41827, 16'd56767, 16'd35574, 16'd54263, 16'd4624, 16'd61018, 16'd49360, 16'd26602, 16'd29023, 16'd22940, 16'd30523, 16'd63797, 16'd61492, 16'd34004, 16'd9519, 16'd5429, 16'd62158, 16'd52758});
	test_expansion(128'h4c454d05af06119f22d5925826976818, {16'd22697, 16'd28949, 16'd557, 16'd32234, 16'd59090, 16'd44323, 16'd39583, 16'd36598, 16'd48433, 16'd11378, 16'd51566, 16'd33942, 16'd24186, 16'd23251, 16'd940, 16'd22797, 16'd64500, 16'd55648, 16'd1321, 16'd17236, 16'd51511, 16'd54376, 16'd49268, 16'd41268, 16'd7185, 16'd62985});
	test_expansion(128'h848553873816648457e1d0919f0dfc96, {16'd20731, 16'd34435, 16'd62482, 16'd46068, 16'd16836, 16'd60914, 16'd5417, 16'd29588, 16'd30234, 16'd28673, 16'd1977, 16'd9524, 16'd48503, 16'd2162, 16'd11758, 16'd53151, 16'd12228, 16'd17432, 16'd47943, 16'd61276, 16'd41368, 16'd27651, 16'd8640, 16'd28048, 16'd13173, 16'd31835});
	test_expansion(128'h85ee411c191b8e82df3ababafc675b58, {16'd16105, 16'd40924, 16'd56946, 16'd16375, 16'd59767, 16'd18833, 16'd31010, 16'd3782, 16'd12826, 16'd20700, 16'd46809, 16'd17416, 16'd15436, 16'd26272, 16'd52573, 16'd16530, 16'd23554, 16'd1962, 16'd51087, 16'd345, 16'd62471, 16'd34350, 16'd21492, 16'd15822, 16'd42679, 16'd54927});
	test_expansion(128'he5e2d31a85a656a26ec3272f875d634b, {16'd14386, 16'd34827, 16'd897, 16'd32014, 16'd14052, 16'd27720, 16'd31378, 16'd15144, 16'd59387, 16'd6821, 16'd13143, 16'd39015, 16'd42755, 16'd52466, 16'd44975, 16'd51542, 16'd52908, 16'd64222, 16'd47700, 16'd37922, 16'd56222, 16'd53611, 16'd56065, 16'd38910, 16'd5250, 16'd42871});
	test_expansion(128'h87d08ca052e0486d36d56be7819e82f8, {16'd10425, 16'd40984, 16'd40699, 16'd7931, 16'd51537, 16'd33961, 16'd41915, 16'd13297, 16'd26496, 16'd10200, 16'd20105, 16'd53459, 16'd11361, 16'd4593, 16'd9410, 16'd45466, 16'd39837, 16'd23167, 16'd12818, 16'd39344, 16'd61898, 16'd45957, 16'd4947, 16'd17801, 16'd33202, 16'd27301});
	test_expansion(128'h022d05774dc5e3f465c5049e73969d61, {16'd1223, 16'd8309, 16'd52714, 16'd38769, 16'd41799, 16'd1509, 16'd61967, 16'd57095, 16'd14302, 16'd17135, 16'd33537, 16'd2566, 16'd33590, 16'd27932, 16'd42460, 16'd16078, 16'd27246, 16'd56842, 16'd8051, 16'd15376, 16'd52790, 16'd29480, 16'd45747, 16'd49217, 16'd17124, 16'd53508});
	test_expansion(128'h73792d51a9e10174fe3633382649e194, {16'd21430, 16'd26253, 16'd17479, 16'd57160, 16'd28512, 16'd58332, 16'd509, 16'd28075, 16'd7448, 16'd28592, 16'd49605, 16'd43488, 16'd63525, 16'd23202, 16'd63412, 16'd289, 16'd22715, 16'd53033, 16'd23285, 16'd32984, 16'd44958, 16'd7742, 16'd2286, 16'd11212, 16'd36225, 16'd37172});
	test_expansion(128'hb63e593e53ad848c326901565f769bc8, {16'd26907, 16'd61590, 16'd20510, 16'd60697, 16'd45038, 16'd50052, 16'd337, 16'd3513, 16'd19353, 16'd39355, 16'd12925, 16'd7924, 16'd29316, 16'd21920, 16'd28283, 16'd37727, 16'd57525, 16'd39631, 16'd16466, 16'd23684, 16'd13246, 16'd56209, 16'd21060, 16'd2236, 16'd35317, 16'd15811});
	test_expansion(128'haf39f345d40749f1b864bffc8b68bb18, {16'd43032, 16'd23021, 16'd38889, 16'd59979, 16'd31965, 16'd48853, 16'd33075, 16'd32506, 16'd38672, 16'd61007, 16'd54964, 16'd39517, 16'd33481, 16'd23369, 16'd39221, 16'd9326, 16'd11814, 16'd14047, 16'd22369, 16'd18032, 16'd35153, 16'd5309, 16'd32152, 16'd62528, 16'd64925, 16'd48257});
	test_expansion(128'h6c2cd0df1f2ea97978ba17c476ffae6f, {16'd63287, 16'd30722, 16'd10613, 16'd27600, 16'd9439, 16'd18096, 16'd14797, 16'd50662, 16'd8955, 16'd25185, 16'd14133, 16'd48398, 16'd11485, 16'd10350, 16'd43027, 16'd17624, 16'd7142, 16'd8340, 16'd15403, 16'd38831, 16'd34564, 16'd50283, 16'd4920, 16'd6154, 16'd3220, 16'd65235});
	test_expansion(128'hfc25d5816f707175745c0e43826afd69, {16'd50273, 16'd64068, 16'd11102, 16'd49279, 16'd20266, 16'd38254, 16'd1382, 16'd27750, 16'd11948, 16'd22568, 16'd10420, 16'd49663, 16'd63699, 16'd17349, 16'd18272, 16'd47888, 16'd16342, 16'd10622, 16'd36263, 16'd34186, 16'd16268, 16'd23971, 16'd14575, 16'd56914, 16'd22488, 16'd16594});
	test_expansion(128'h693e1bf34b8f74fcb81622c369fa3ef6, {16'd59716, 16'd15032, 16'd16701, 16'd1849, 16'd53017, 16'd17414, 16'd9938, 16'd6862, 16'd13383, 16'd47926, 16'd16348, 16'd43980, 16'd27583, 16'd38802, 16'd47228, 16'd30156, 16'd33973, 16'd16570, 16'd10443, 16'd53757, 16'd26356, 16'd10125, 16'd27344, 16'd20742, 16'd63922, 16'd23529});
	test_expansion(128'hc357db9aebb1d1e12f5fad3666376d6b, {16'd146, 16'd18118, 16'd37147, 16'd64459, 16'd11869, 16'd752, 16'd3179, 16'd24978, 16'd39926, 16'd42762, 16'd8136, 16'd14644, 16'd52934, 16'd18773, 16'd30408, 16'd63929, 16'd61266, 16'd15389, 16'd16587, 16'd39761, 16'd28276, 16'd57328, 16'd45695, 16'd43023, 16'd43495, 16'd50423});
	test_expansion(128'h9dff5eb532fcd5de6da296296ae3fcbb, {16'd37557, 16'd65387, 16'd28033, 16'd61104, 16'd2031, 16'd5837, 16'd52417, 16'd14290, 16'd51600, 16'd24399, 16'd56386, 16'd15241, 16'd41767, 16'd25286, 16'd15784, 16'd48207, 16'd13434, 16'd37726, 16'd30750, 16'd48488, 16'd36842, 16'd29809, 16'd41460, 16'd46250, 16'd12116, 16'd14563});
	test_expansion(128'ha1097d88a183072aae6077c67a6f9dd2, {16'd7174, 16'd9374, 16'd7432, 16'd43483, 16'd65356, 16'd39883, 16'd30775, 16'd45148, 16'd61484, 16'd35968, 16'd9578, 16'd36938, 16'd17329, 16'd16656, 16'd11157, 16'd15634, 16'd31027, 16'd5090, 16'd56319, 16'd15352, 16'd64687, 16'd13552, 16'd60656, 16'd56334, 16'd56463, 16'd50589});
	test_expansion(128'h0656cb31c11ab5a13577aa0adc199469, {16'd1624, 16'd2217, 16'd57235, 16'd38514, 16'd14079, 16'd46662, 16'd28495, 16'd24184, 16'd52211, 16'd24376, 16'd41568, 16'd46392, 16'd702, 16'd13919, 16'd44676, 16'd41049, 16'd10153, 16'd11742, 16'd28481, 16'd5728, 16'd4186, 16'd50942, 16'd27533, 16'd3634, 16'd40610, 16'd56514});
	test_expansion(128'hadc3a780a28eb44a8d61525ead538663, {16'd5578, 16'd49904, 16'd61213, 16'd50069, 16'd32073, 16'd18455, 16'd21030, 16'd4816, 16'd47472, 16'd33845, 16'd27097, 16'd41414, 16'd28761, 16'd12519, 16'd48750, 16'd7558, 16'd28436, 16'd61949, 16'd5955, 16'd32202, 16'd9289, 16'd21920, 16'd64304, 16'd43133, 16'd65372, 16'd61492});
	test_expansion(128'hdab5f6d8c244d789a36023a72aa817ae, {16'd54196, 16'd58566, 16'd38516, 16'd5196, 16'd42148, 16'd15319, 16'd63031, 16'd36264, 16'd25183, 16'd31105, 16'd8562, 16'd39536, 16'd6157, 16'd14673, 16'd2687, 16'd12286, 16'd15735, 16'd56370, 16'd56726, 16'd29691, 16'd33774, 16'd15587, 16'd18524, 16'd33054, 16'd64837, 16'd36881});
	test_expansion(128'h6042502208b52176028656051591eeb2, {16'd51258, 16'd49828, 16'd11789, 16'd62621, 16'd29817, 16'd64789, 16'd13906, 16'd13838, 16'd31156, 16'd2703, 16'd8657, 16'd59097, 16'd7526, 16'd50736, 16'd35962, 16'd4570, 16'd59173, 16'd18923, 16'd47507, 16'd41671, 16'd8757, 16'd34475, 16'd147, 16'd32835, 16'd31432, 16'd63306});
	test_expansion(128'h347c50c4c5a846ff449da251248ac92c, {16'd13309, 16'd18659, 16'd19843, 16'd56694, 16'd56435, 16'd52454, 16'd58205, 16'd32587, 16'd55388, 16'd6536, 16'd61608, 16'd17314, 16'd61834, 16'd45949, 16'd19914, 16'd27945, 16'd59567, 16'd3721, 16'd51717, 16'd23415, 16'd2643, 16'd47742, 16'd40899, 16'd15183, 16'd55803, 16'd65341});
	test_expansion(128'h09d4fc5d8179a74ae30cdc36f40758e9, {16'd60749, 16'd3322, 16'd3556, 16'd52444, 16'd14586, 16'd37169, 16'd60559, 16'd34701, 16'd36753, 16'd51216, 16'd36383, 16'd46335, 16'd34975, 16'd15002, 16'd61979, 16'd12781, 16'd53805, 16'd43277, 16'd18810, 16'd31314, 16'd37126, 16'd63700, 16'd61443, 16'd8937, 16'd24864, 16'd6987});
	test_expansion(128'h04e3d0923c0bd8a780d8c9c678f47227, {16'd58959, 16'd22819, 16'd58799, 16'd38122, 16'd26352, 16'd19115, 16'd12520, 16'd3523, 16'd12333, 16'd6497, 16'd14025, 16'd37701, 16'd18853, 16'd2474, 16'd7107, 16'd8013, 16'd32825, 16'd33995, 16'd50900, 16'd36305, 16'd21105, 16'd38915, 16'd62114, 16'd33323, 16'd7981, 16'd25641});
	test_expansion(128'h678181608df7a8384f6d148587c0a3d1, {16'd1791, 16'd43371, 16'd1391, 16'd45920, 16'd30731, 16'd49205, 16'd35884, 16'd26274, 16'd20754, 16'd43796, 16'd54253, 16'd53998, 16'd15394, 16'd10995, 16'd38549, 16'd1222, 16'd15902, 16'd1882, 16'd30226, 16'd63778, 16'd51380, 16'd20416, 16'd13828, 16'd31054, 16'd19327, 16'd52599});
	test_expansion(128'h58832186b13f65e7e26916798db55e9e, {16'd20710, 16'd18761, 16'd44485, 16'd18379, 16'd12112, 16'd25908, 16'd2338, 16'd34179, 16'd34465, 16'd15134, 16'd47255, 16'd37537, 16'd39603, 16'd16012, 16'd6090, 16'd19031, 16'd39157, 16'd48601, 16'd38265, 16'd61405, 16'd55692, 16'd35011, 16'd54739, 16'd6373, 16'd20647, 16'd12203});
	test_expansion(128'h19a8ebd646e658cddee7f6c73a90831d, {16'd38599, 16'd41775, 16'd17607, 16'd18451, 16'd28867, 16'd29887, 16'd41010, 16'd2281, 16'd13506, 16'd27447, 16'd50713, 16'd30217, 16'd32548, 16'd52701, 16'd17796, 16'd43598, 16'd53638, 16'd59973, 16'd8944, 16'd6345, 16'd45260, 16'd20202, 16'd65201, 16'd47271, 16'd28855, 16'd36003});
	test_expansion(128'h732078d614c01f8d6ae4325e7e5d78de, {16'd54256, 16'd14695, 16'd8035, 16'd404, 16'd60978, 16'd31942, 16'd25897, 16'd50340, 16'd49374, 16'd7625, 16'd4198, 16'd42949, 16'd20925, 16'd26834, 16'd16641, 16'd59415, 16'd40528, 16'd49585, 16'd36538, 16'd62559, 16'd64970, 16'd24128, 16'd7474, 16'd54863, 16'd14882, 16'd49664});
	test_expansion(128'hc616b0788520e260d066a1475aa8bc3c, {16'd13787, 16'd51224, 16'd39624, 16'd48778, 16'd3227, 16'd27111, 16'd46141, 16'd19859, 16'd21160, 16'd33143, 16'd9461, 16'd45295, 16'd23265, 16'd2415, 16'd42333, 16'd43119, 16'd50712, 16'd39783, 16'd54650, 16'd32187, 16'd63151, 16'd46039, 16'd40442, 16'd35457, 16'd40650, 16'd2072});
	test_expansion(128'h7cbed21bf85294d256ece86e405a1ce5, {16'd62644, 16'd9675, 16'd41393, 16'd39904, 16'd19643, 16'd35531, 16'd24591, 16'd646, 16'd24747, 16'd17556, 16'd39675, 16'd54217, 16'd30043, 16'd33406, 16'd48340, 16'd59650, 16'd35905, 16'd6593, 16'd60101, 16'd6757, 16'd15530, 16'd41951, 16'd8413, 16'd30257, 16'd21017, 16'd40267});
	test_expansion(128'h5d594a4e9bdae94dc63c9d5f42b1becd, {16'd13293, 16'd5536, 16'd57921, 16'd54910, 16'd23118, 16'd63681, 16'd8388, 16'd6959, 16'd34302, 16'd43700, 16'd26045, 16'd8750, 16'd42282, 16'd58320, 16'd34885, 16'd38696, 16'd29593, 16'd43188, 16'd35690, 16'd6953, 16'd47204, 16'd13923, 16'd32252, 16'd37226, 16'd21364, 16'd64846});
	test_expansion(128'h301edc8fe58a38c1f8c86ba64ca45128, {16'd36656, 16'd27810, 16'd14955, 16'd34541, 16'd53662, 16'd6850, 16'd46584, 16'd15699, 16'd5720, 16'd49812, 16'd36870, 16'd12448, 16'd17472, 16'd64629, 16'd6297, 16'd16286, 16'd58540, 16'd57116, 16'd64808, 16'd35379, 16'd30866, 16'd61023, 16'd40808, 16'd4164, 16'd1273, 16'd23573});
	test_expansion(128'h5231af11090532018bf8785505112f55, {16'd32673, 16'd2741, 16'd64539, 16'd49430, 16'd22791, 16'd60531, 16'd40649, 16'd27396, 16'd19505, 16'd13401, 16'd26328, 16'd38303, 16'd11216, 16'd44456, 16'd26839, 16'd9075, 16'd13916, 16'd33244, 16'd6189, 16'd63631, 16'd51521, 16'd19625, 16'd8659, 16'd952, 16'd60758, 16'd58381});
	test_expansion(128'h25692198fa25e7c2f58e1d859c6fddee, {16'd3558, 16'd11024, 16'd59089, 16'd57923, 16'd42549, 16'd41228, 16'd39004, 16'd26672, 16'd48119, 16'd37867, 16'd18720, 16'd24564, 16'd48483, 16'd34003, 16'd28383, 16'd36167, 16'd46195, 16'd16668, 16'd60723, 16'd56050, 16'd58039, 16'd24144, 16'd41297, 16'd13440, 16'd47894, 16'd48221});
	test_expansion(128'h33a730050ff69f67d42ea9606e403ceb, {16'd24793, 16'd11448, 16'd37647, 16'd30385, 16'd62862, 16'd33553, 16'd62526, 16'd58839, 16'd65412, 16'd4491, 16'd44493, 16'd57850, 16'd6792, 16'd2204, 16'd10782, 16'd4946, 16'd38200, 16'd55557, 16'd2310, 16'd48831, 16'd19838, 16'd41921, 16'd64955, 16'd62877, 16'd37130, 16'd52222});
	test_expansion(128'hd86356be2d603343ce07449d6b80eacb, {16'd29569, 16'd29920, 16'd45307, 16'd27839, 16'd32933, 16'd18361, 16'd62865, 16'd23161, 16'd9610, 16'd57760, 16'd27548, 16'd55521, 16'd14417, 16'd31068, 16'd39115, 16'd57339, 16'd36291, 16'd50921, 16'd57584, 16'd64691, 16'd30532, 16'd21985, 16'd43284, 16'd25906, 16'd11621, 16'd34964});
	test_expansion(128'h9547c9edf4655afced1c58f0e83ea880, {16'd5816, 16'd47069, 16'd30768, 16'd44860, 16'd27829, 16'd54739, 16'd35050, 16'd25604, 16'd9487, 16'd2580, 16'd43329, 16'd47006, 16'd14388, 16'd12973, 16'd63084, 16'd54931, 16'd45607, 16'd21977, 16'd65362, 16'd42104, 16'd28171, 16'd52038, 16'd10910, 16'd12102, 16'd39938, 16'd14706});
	test_expansion(128'hf86d1c11b267136ebe85b95f24b473e3, {16'd63752, 16'd19852, 16'd46967, 16'd5051, 16'd9427, 16'd2116, 16'd41136, 16'd31290, 16'd14371, 16'd18889, 16'd28712, 16'd18103, 16'd12908, 16'd39155, 16'd16659, 16'd21484, 16'd30758, 16'd1941, 16'd12898, 16'd15254, 16'd5145, 16'd30740, 16'd859, 16'd57194, 16'd32328, 16'd46001});
	test_expansion(128'h30b2f26699dc48fc009d5a15267dbd3e, {16'd34708, 16'd51673, 16'd15794, 16'd48350, 16'd40326, 16'd21349, 16'd7540, 16'd62117, 16'd51709, 16'd38887, 16'd9516, 16'd83, 16'd30545, 16'd43062, 16'd25621, 16'd12084, 16'd43360, 16'd54681, 16'd27925, 16'd40392, 16'd51018, 16'd8489, 16'd4470, 16'd59230, 16'd1212, 16'd45303});
	test_expansion(128'hcb5cdb0ab2644cbb475d52bb15d65a55, {16'd33482, 16'd16148, 16'd16088, 16'd57768, 16'd20633, 16'd6317, 16'd15883, 16'd53618, 16'd57413, 16'd63642, 16'd8575, 16'd38659, 16'd12390, 16'd13957, 16'd24973, 16'd42836, 16'd15851, 16'd10551, 16'd26393, 16'd20282, 16'd8378, 16'd63429, 16'd62154, 16'd64147, 16'd45134, 16'd21507});
	test_expansion(128'h919bb7ca34f8cfcdd127e10db1da491c, {16'd1476, 16'd20775, 16'd22907, 16'd33446, 16'd14082, 16'd54052, 16'd55775, 16'd36726, 16'd13905, 16'd60716, 16'd6859, 16'd15663, 16'd49060, 16'd16436, 16'd9760, 16'd24281, 16'd18752, 16'd39446, 16'd25736, 16'd16542, 16'd41205, 16'd58222, 16'd38777, 16'd6652, 16'd24931, 16'd60195});
	test_expansion(128'hc0124ada8bdb4b1f1cc624bf118165ea, {16'd26025, 16'd58313, 16'd53134, 16'd33621, 16'd45634, 16'd8017, 16'd23848, 16'd20774, 16'd40303, 16'd12872, 16'd2881, 16'd19230, 16'd25596, 16'd15857, 16'd31914, 16'd59104, 16'd37845, 16'd663, 16'd39617, 16'd60108, 16'd48567, 16'd58557, 16'd31636, 16'd63560, 16'd19244, 16'd58983});
	test_expansion(128'h4a52b632bbe7fa03f24db5fd0fb458e1, {16'd10587, 16'd57188, 16'd24269, 16'd53502, 16'd14268, 16'd17886, 16'd41603, 16'd8603, 16'd13132, 16'd48613, 16'd33623, 16'd25156, 16'd50839, 16'd27421, 16'd7099, 16'd39104, 16'd9790, 16'd43502, 16'd2172, 16'd58024, 16'd64309, 16'd22179, 16'd34049, 16'd37798, 16'd20124, 16'd12564});
	test_expansion(128'ha6d28fa63c4257d73c79b2d8c468d7f1, {16'd58622, 16'd20553, 16'd52451, 16'd50799, 16'd22223, 16'd2474, 16'd13215, 16'd2010, 16'd5544, 16'd9252, 16'd34621, 16'd23059, 16'd48516, 16'd32842, 16'd379, 16'd3880, 16'd59606, 16'd56709, 16'd60990, 16'd24378, 16'd47616, 16'd33926, 16'd8103, 16'd402, 16'd40031, 16'd33691});
	test_expansion(128'h13186ebe7002b6853fa4752be6c2de40, {16'd28844, 16'd10975, 16'd59810, 16'd8510, 16'd6702, 16'd18878, 16'd22249, 16'd56210, 16'd461, 16'd52956, 16'd40721, 16'd41043, 16'd16094, 16'd7650, 16'd56541, 16'd5138, 16'd7835, 16'd59963, 16'd40806, 16'd50918, 16'd64337, 16'd11258, 16'd9436, 16'd59830, 16'd64157, 16'd36304});
	test_expansion(128'h732e133866ccce25bf9d89cb085d1b36, {16'd42296, 16'd19808, 16'd55396, 16'd65273, 16'd44858, 16'd13185, 16'd55645, 16'd3209, 16'd9909, 16'd29714, 16'd34990, 16'd49212, 16'd19999, 16'd37074, 16'd7691, 16'd13382, 16'd40716, 16'd56325, 16'd53661, 16'd43331, 16'd24992, 16'd28752, 16'd61330, 16'd36616, 16'd15114, 16'd29554});
	test_expansion(128'h1ea6910a1878644f85b91d26a97bf246, {16'd14200, 16'd29797, 16'd43853, 16'd23100, 16'd58738, 16'd59715, 16'd11541, 16'd18655, 16'd15590, 16'd64132, 16'd62975, 16'd23694, 16'd64476, 16'd16673, 16'd3866, 16'd12037, 16'd3861, 16'd42748, 16'd32950, 16'd22966, 16'd51457, 16'd32469, 16'd31237, 16'd8782, 16'd27753, 16'd29285});
	test_expansion(128'h8f0635bba97a1be0384d509d8cae1f34, {16'd53405, 16'd62949, 16'd41637, 16'd12248, 16'd10846, 16'd6278, 16'd34849, 16'd32386, 16'd42332, 16'd49303, 16'd22704, 16'd30860, 16'd56153, 16'd11832, 16'd39215, 16'd5247, 16'd23083, 16'd60630, 16'd25433, 16'd48927, 16'd14830, 16'd10056, 16'd12184, 16'd32319, 16'd37613, 16'd37082});
	test_expansion(128'h2409db46f9c5c18513a23d6783b01f6b, {16'd52982, 16'd22804, 16'd23753, 16'd63388, 16'd28255, 16'd52010, 16'd45058, 16'd15956, 16'd36915, 16'd46054, 16'd10081, 16'd25095, 16'd35616, 16'd4079, 16'd22508, 16'd16450, 16'd22422, 16'd39073, 16'd26737, 16'd59722, 16'd9899, 16'd60624, 16'd58386, 16'd44685, 16'd34531, 16'd31358});
	test_expansion(128'hb428b10dfaa9864a808b844534b84805, {16'd10012, 16'd56666, 16'd26867, 16'd35352, 16'd26687, 16'd61157, 16'd31604, 16'd10022, 16'd35054, 16'd2824, 16'd33376, 16'd18297, 16'd25811, 16'd38161, 16'd41241, 16'd11358, 16'd28574, 16'd31484, 16'd61385, 16'd27831, 16'd44882, 16'd48983, 16'd31429, 16'd41644, 16'd2479, 16'd21719});
	test_expansion(128'h7bfc5b44280e918ec09c8daa4dbeab17, {16'd33584, 16'd58371, 16'd51626, 16'd5148, 16'd43469, 16'd48623, 16'd15830, 16'd22858, 16'd32241, 16'd44753, 16'd61544, 16'd61972, 16'd63139, 16'd64231, 16'd45244, 16'd15013, 16'd17357, 16'd56442, 16'd65287, 16'd10987, 16'd62639, 16'd41871, 16'd52279, 16'd30485, 16'd51147, 16'd11510});
	test_expansion(128'h7cd7e4a3a6175e54a32ee3c766208ce7, {16'd47656, 16'd15281, 16'd31340, 16'd34822, 16'd41015, 16'd49120, 16'd61380, 16'd52352, 16'd36651, 16'd61676, 16'd62336, 16'd33393, 16'd16970, 16'd4603, 16'd21422, 16'd19249, 16'd33286, 16'd11541, 16'd31539, 16'd64330, 16'd57778, 16'd58803, 16'd13768, 16'd45210, 16'd31509, 16'd25140});
	test_expansion(128'hf5701af2a9585fb524f60ef1bb959434, {16'd2760, 16'd43784, 16'd14073, 16'd12792, 16'd63628, 16'd63140, 16'd53860, 16'd63229, 16'd4202, 16'd31278, 16'd19594, 16'd32398, 16'd51621, 16'd39684, 16'd61259, 16'd41006, 16'd15307, 16'd47486, 16'd48243, 16'd43091, 16'd62177, 16'd31746, 16'd31051, 16'd22434, 16'd55126, 16'd45644});
	test_expansion(128'h7255a7e0b73f85e271b1dd0e4eed3b21, {16'd15569, 16'd6976, 16'd16155, 16'd61628, 16'd64322, 16'd30200, 16'd37575, 16'd51972, 16'd39608, 16'd32580, 16'd35829, 16'd37430, 16'd55697, 16'd32423, 16'd11695, 16'd53346, 16'd13985, 16'd10825, 16'd63913, 16'd55461, 16'd22576, 16'd54733, 16'd9916, 16'd43203, 16'd48363, 16'd7640});
	test_expansion(128'h1818415d11acdfe40e6f5ed09f5b9bfc, {16'd65089, 16'd3470, 16'd60819, 16'd9609, 16'd53123, 16'd59272, 16'd23058, 16'd54896, 16'd24235, 16'd16986, 16'd36031, 16'd20700, 16'd3656, 16'd28471, 16'd59468, 16'd23672, 16'd13653, 16'd38968, 16'd12594, 16'd31505, 16'd51806, 16'd65428, 16'd62694, 16'd60218, 16'd34107, 16'd269});
	test_expansion(128'h8fde45e46328d8572b41071528dcf158, {16'd19449, 16'd51054, 16'd6119, 16'd21621, 16'd1737, 16'd9293, 16'd22242, 16'd11163, 16'd52670, 16'd22046, 16'd41060, 16'd38309, 16'd42405, 16'd32595, 16'd40230, 16'd25248, 16'd3188, 16'd20971, 16'd62940, 16'd9663, 16'd22256, 16'd19207, 16'd51773, 16'd6129, 16'd62194, 16'd8630});
	test_expansion(128'h51f5cf976ba271dddd1597d68707d50a, {16'd44245, 16'd16730, 16'd60939, 16'd48463, 16'd46705, 16'd29142, 16'd25151, 16'd30551, 16'd61382, 16'd58942, 16'd37388, 16'd51936, 16'd18737, 16'd50846, 16'd13925, 16'd15652, 16'd28241, 16'd48484, 16'd12665, 16'd18013, 16'd7622, 16'd49624, 16'd6274, 16'd54563, 16'd25447, 16'd47382});
	test_expansion(128'h130668aa0a4296fd03bd11c23724f6e9, {16'd61418, 16'd30313, 16'd20296, 16'd60997, 16'd16536, 16'd37444, 16'd12018, 16'd41749, 16'd13028, 16'd34920, 16'd29757, 16'd23881, 16'd45768, 16'd29487, 16'd33741, 16'd48396, 16'd61064, 16'd11350, 16'd58859, 16'd61610, 16'd48622, 16'd3557, 16'd13298, 16'd63125, 16'd5951, 16'd59788});
	test_expansion(128'h97dbc51ef36dcc0ea9e148029c917afd, {16'd43242, 16'd26130, 16'd54741, 16'd59338, 16'd58457, 16'd60850, 16'd36708, 16'd242, 16'd57165, 16'd12647, 16'd39530, 16'd2510, 16'd38027, 16'd54272, 16'd38505, 16'd22204, 16'd27487, 16'd44787, 16'd59989, 16'd19708, 16'd37333, 16'd39044, 16'd45498, 16'd29669, 16'd31397, 16'd33854});
	test_expansion(128'h42fd2b61cc9e1ed32ebd00fec94e2b1f, {16'd44153, 16'd52407, 16'd48164, 16'd7912, 16'd22807, 16'd46084, 16'd43797, 16'd18956, 16'd22708, 16'd32543, 16'd51827, 16'd61745, 16'd30461, 16'd59295, 16'd15183, 16'd65153, 16'd32980, 16'd4547, 16'd944, 16'd45551, 16'd19740, 16'd42991, 16'd1697, 16'd8735, 16'd58512, 16'd37752});
	test_expansion(128'h86d85ff40f9713f238bb5e931a8e8a54, {16'd62642, 16'd53958, 16'd59561, 16'd44662, 16'd19797, 16'd18779, 16'd60228, 16'd59802, 16'd40502, 16'd36118, 16'd6714, 16'd34750, 16'd61880, 16'd42120, 16'd46467, 16'd17977, 16'd25548, 16'd2563, 16'd11652, 16'd28975, 16'd28859, 16'd3013, 16'd47026, 16'd5167, 16'd1395, 16'd8923});
	test_expansion(128'h4526c07343896b7ef0af3f5ab453e2cf, {16'd33865, 16'd48263, 16'd19668, 16'd33873, 16'd57489, 16'd63709, 16'd6194, 16'd30029, 16'd12437, 16'd6570, 16'd46540, 16'd35827, 16'd58399, 16'd13025, 16'd17628, 16'd51184, 16'd60635, 16'd29446, 16'd2089, 16'd23515, 16'd45076, 16'd14113, 16'd32909, 16'd14653, 16'd20223, 16'd58952});
	test_expansion(128'hc20170709427eb74578a9d844fa26b87, {16'd51168, 16'd47796, 16'd51918, 16'd3732, 16'd6879, 16'd51606, 16'd20097, 16'd42142, 16'd32401, 16'd64881, 16'd1806, 16'd17875, 16'd59909, 16'd24669, 16'd23572, 16'd52220, 16'd20646, 16'd5812, 16'd38498, 16'd31789, 16'd26653, 16'd27090, 16'd20584, 16'd22198, 16'd10280, 16'd13416});
	test_expansion(128'h1abef658fb234faddc5bb162771cdfcf, {16'd29866, 16'd61154, 16'd11483, 16'd36147, 16'd51913, 16'd5087, 16'd34368, 16'd58084, 16'd63222, 16'd45511, 16'd12922, 16'd10021, 16'd12019, 16'd6387, 16'd34538, 16'd6383, 16'd60725, 16'd13572, 16'd46418, 16'd51895, 16'd27390, 16'd50462, 16'd52126, 16'd59125, 16'd6397, 16'd20746});
	test_expansion(128'h8edce513dac243032802960ea8d18735, {16'd62864, 16'd9446, 16'd34046, 16'd43798, 16'd4116, 16'd24808, 16'd32125, 16'd40790, 16'd13971, 16'd17659, 16'd58268, 16'd32451, 16'd51556, 16'd15680, 16'd60411, 16'd3226, 16'd601, 16'd29143, 16'd7461, 16'd27127, 16'd14156, 16'd62487, 16'd15546, 16'd37132, 16'd51506, 16'd56894});
	test_expansion(128'hf6e9dba3a5aa4445fa4fcb061d686ea2, {16'd23332, 16'd17603, 16'd51746, 16'd64533, 16'd43451, 16'd25758, 16'd35694, 16'd7960, 16'd35174, 16'd41205, 16'd20616, 16'd34216, 16'd17915, 16'd33976, 16'd37800, 16'd14382, 16'd50726, 16'd64624, 16'd34314, 16'd45042, 16'd46270, 16'd24212, 16'd31826, 16'd58625, 16'd27916, 16'd63112});
	test_expansion(128'h7d18317b91fb348c8b2fcc1fb3e00dd5, {16'd5953, 16'd47450, 16'd60378, 16'd63672, 16'd20281, 16'd22639, 16'd62675, 16'd42488, 16'd37281, 16'd29899, 16'd61319, 16'd54104, 16'd21004, 16'd37025, 16'd27410, 16'd7351, 16'd64174, 16'd46852, 16'd17772, 16'd54877, 16'd30179, 16'd51607, 16'd2970, 16'd10731, 16'd29973, 16'd18051});
	test_expansion(128'h6fc8451eb0c27229a395f7f549b7556b, {16'd28735, 16'd63038, 16'd51160, 16'd26821, 16'd25241, 16'd17565, 16'd45451, 16'd24436, 16'd59819, 16'd54431, 16'd61870, 16'd39411, 16'd37693, 16'd6216, 16'd1592, 16'd9114, 16'd44914, 16'd23253, 16'd46946, 16'd6648, 16'd35309, 16'd3178, 16'd30379, 16'd61413, 16'd14603, 16'd7574});
	test_expansion(128'h1b85235b0284e9de47016b9ebbfc8046, {16'd14399, 16'd5057, 16'd37403, 16'd1947, 16'd54483, 16'd17238, 16'd29017, 16'd59545, 16'd41982, 16'd41550, 16'd12139, 16'd52770, 16'd20150, 16'd43384, 16'd52090, 16'd3328, 16'd38737, 16'd64932, 16'd12726, 16'd52725, 16'd16635, 16'd14908, 16'd4923, 16'd20893, 16'd31441, 16'd25396});
	test_expansion(128'h35b8a11a2b399eae8596fbb2807d5e93, {16'd31871, 16'd32604, 16'd15004, 16'd34102, 16'd65181, 16'd32740, 16'd51077, 16'd45731, 16'd22681, 16'd3381, 16'd12184, 16'd13904, 16'd58733, 16'd17594, 16'd42359, 16'd65527, 16'd37950, 16'd39929, 16'd24969, 16'd45901, 16'd19434, 16'd44426, 16'd52319, 16'd48323, 16'd62834, 16'd35096});
	test_expansion(128'h0f592e0a025c1569371adfa7a055d099, {16'd1095, 16'd30523, 16'd39013, 16'd50058, 16'd21948, 16'd45070, 16'd34617, 16'd2145, 16'd51805, 16'd60727, 16'd10825, 16'd31902, 16'd37825, 16'd28527, 16'd8359, 16'd11473, 16'd1693, 16'd58293, 16'd4684, 16'd59033, 16'd59834, 16'd24705, 16'd9462, 16'd39131, 16'd54728, 16'd47894});
	test_expansion(128'h01e7e40975e23a221ddad1089e09300d, {16'd63652, 16'd34124, 16'd13532, 16'd27499, 16'd46411, 16'd2309, 16'd24496, 16'd59955, 16'd17270, 16'd27482, 16'd32706, 16'd50595, 16'd25526, 16'd6208, 16'd30702, 16'd33564, 16'd13277, 16'd29501, 16'd38389, 16'd43396, 16'd49727, 16'd62380, 16'd4698, 16'd14431, 16'd48653, 16'd43075});
	test_expansion(128'hf6708f3a9bd6b782447decd29491b755, {16'd8868, 16'd24218, 16'd3974, 16'd53297, 16'd42697, 16'd41013, 16'd58766, 16'd58918, 16'd3511, 16'd49161, 16'd5298, 16'd54048, 16'd41527, 16'd1332, 16'd63303, 16'd50670, 16'd20818, 16'd56156, 16'd54332, 16'd6318, 16'd18715, 16'd44931, 16'd31253, 16'd44996, 16'd33240, 16'd63984});
	test_expansion(128'h042cc13118c9be90b0c8e041f756c806, {16'd8921, 16'd42590, 16'd34714, 16'd47265, 16'd61230, 16'd53631, 16'd27258, 16'd16884, 16'd35930, 16'd12053, 16'd36359, 16'd39202, 16'd12559, 16'd18935, 16'd7524, 16'd54632, 16'd27131, 16'd18760, 16'd45894, 16'd24690, 16'd53989, 16'd36439, 16'd22950, 16'd19699, 16'd6053, 16'd35970});
	test_expansion(128'h7b4d803d60c95abb7dc61e33f3dcf8b6, {16'd13191, 16'd27186, 16'd36154, 16'd57701, 16'd52436, 16'd27599, 16'd56137, 16'd22885, 16'd55759, 16'd31641, 16'd31892, 16'd21084, 16'd37770, 16'd58248, 16'd59313, 16'd62060, 16'd1685, 16'd14831, 16'd10465, 16'd29733, 16'd20205, 16'd59059, 16'd9043, 16'd19946, 16'd36341, 16'd47672});
	test_expansion(128'hd5f0eb14bff3c9d39d64e20d5cafebed, {16'd63538, 16'd13777, 16'd54252, 16'd8324, 16'd8781, 16'd16760, 16'd5212, 16'd35367, 16'd52263, 16'd29500, 16'd62448, 16'd45246, 16'd37009, 16'd43795, 16'd5858, 16'd32079, 16'd25819, 16'd40630, 16'd22004, 16'd32977, 16'd41129, 16'd5632, 16'd45904, 16'd23848, 16'd21738, 16'd3931});
	test_expansion(128'h11dbc59c955c9af9c6e282ff3fc33d30, {16'd56133, 16'd62473, 16'd52232, 16'd63029, 16'd3878, 16'd64179, 16'd47956, 16'd58382, 16'd17407, 16'd38734, 16'd23776, 16'd52627, 16'd25159, 16'd18226, 16'd20083, 16'd17218, 16'd9611, 16'd1812, 16'd63836, 16'd57712, 16'd15894, 16'd5345, 16'd39542, 16'd46250, 16'd2185, 16'd25201});
	test_expansion(128'h56957e13c3804caf6814d2d909212ea3, {16'd2193, 16'd628, 16'd62183, 16'd50587, 16'd9835, 16'd22370, 16'd18178, 16'd31709, 16'd42170, 16'd49430, 16'd5417, 16'd41438, 16'd48647, 16'd19925, 16'd40370, 16'd43178, 16'd42032, 16'd54873, 16'd46196, 16'd14493, 16'd54474, 16'd25931, 16'd19759, 16'd25374, 16'd4084, 16'd36194});
	test_expansion(128'h69c36c631de6b663ba05a3770210e086, {16'd52396, 16'd42829, 16'd13692, 16'd42672, 16'd43904, 16'd26773, 16'd6299, 16'd14819, 16'd3868, 16'd8155, 16'd4272, 16'd11604, 16'd3885, 16'd61534, 16'd49707, 16'd42292, 16'd20406, 16'd49516, 16'd22863, 16'd50862, 16'd22516, 16'd54877, 16'd22261, 16'd25390, 16'd50620, 16'd60973});
	test_expansion(128'hb14c5f0bcf229297662e89a8496b8a65, {16'd33416, 16'd38671, 16'd51717, 16'd48814, 16'd6107, 16'd34577, 16'd29974, 16'd48927, 16'd38947, 16'd60245, 16'd41386, 16'd59288, 16'd61455, 16'd6275, 16'd22134, 16'd30608, 16'd7328, 16'd20185, 16'd8609, 16'd18586, 16'd27401, 16'd15959, 16'd19517, 16'd23801, 16'd17544, 16'd37614});
	test_expansion(128'h304199ae4218438ff10a6d0af89fdd3a, {16'd53289, 16'd27169, 16'd29040, 16'd14678, 16'd6992, 16'd62843, 16'd33733, 16'd39599, 16'd38171, 16'd28040, 16'd45140, 16'd28180, 16'd7866, 16'd2433, 16'd2112, 16'd31769, 16'd4985, 16'd37808, 16'd58689, 16'd51995, 16'd6113, 16'd49296, 16'd8648, 16'd13093, 16'd64664, 16'd48485});
	test_expansion(128'ha1dd2f42499670495a9ae96adcc2c654, {16'd61885, 16'd62587, 16'd10088, 16'd7148, 16'd38434, 16'd55514, 16'd12455, 16'd17689, 16'd63841, 16'd41587, 16'd43347, 16'd61998, 16'd12675, 16'd7346, 16'd29423, 16'd9600, 16'd35434, 16'd29363, 16'd54595, 16'd33273, 16'd1549, 16'd3936, 16'd19363, 16'd13003, 16'd35802, 16'd35739});
	test_expansion(128'ha673e1404abc2a990de57428976f5bdb, {16'd62143, 16'd28974, 16'd51176, 16'd1182, 16'd23132, 16'd57898, 16'd47615, 16'd35904, 16'd6809, 16'd31357, 16'd309, 16'd607, 16'd45907, 16'd23886, 16'd35079, 16'd20905, 16'd64838, 16'd9462, 16'd9314, 16'd1806, 16'd40964, 16'd12248, 16'd64899, 16'd13018, 16'd5252, 16'd18066});
	test_expansion(128'h8a60c07b8644b85d5c61297b5f6b3553, {16'd48597, 16'd53971, 16'd52758, 16'd62370, 16'd37270, 16'd58592, 16'd20732, 16'd26935, 16'd26186, 16'd42832, 16'd14138, 16'd3516, 16'd52366, 16'd30088, 16'd25312, 16'd45484, 16'd33692, 16'd59162, 16'd22161, 16'd61494, 16'd10371, 16'd27570, 16'd61753, 16'd15877, 16'd57310, 16'd34501});
	test_expansion(128'h000d4b7d1b6c299bd188cf06f3501f7d, {16'd22757, 16'd60014, 16'd16946, 16'd47173, 16'd28382, 16'd43193, 16'd34391, 16'd15705, 16'd937, 16'd56366, 16'd54512, 16'd26120, 16'd34843, 16'd48167, 16'd62891, 16'd46830, 16'd17729, 16'd1419, 16'd3704, 16'd31088, 16'd33956, 16'd38118, 16'd5082, 16'd23893, 16'd55875, 16'd27214});
	test_expansion(128'h758da4148cfd334990a0df117105bb9d, {16'd6540, 16'd16050, 16'd36699, 16'd17091, 16'd39027, 16'd59246, 16'd1571, 16'd52554, 16'd60169, 16'd63438, 16'd24324, 16'd13720, 16'd60480, 16'd27529, 16'd31909, 16'd43024, 16'd8929, 16'd22582, 16'd32994, 16'd29053, 16'd35359, 16'd3541, 16'd46904, 16'd48561, 16'd24907, 16'd10809});
	test_expansion(128'h22a10607a69391158a15882cf1976c4a, {16'd36548, 16'd48094, 16'd2352, 16'd39634, 16'd22425, 16'd12868, 16'd18397, 16'd25376, 16'd42690, 16'd35197, 16'd48080, 16'd35615, 16'd6154, 16'd54933, 16'd57566, 16'd28106, 16'd8833, 16'd48875, 16'd32210, 16'd64619, 16'd21165, 16'd9398, 16'd18047, 16'd44208, 16'd47020, 16'd42828});
	test_expansion(128'h21d47a00d30479f4019fd73ad578da2e, {16'd16488, 16'd46967, 16'd48304, 16'd57619, 16'd18377, 16'd59699, 16'd27797, 16'd31308, 16'd812, 16'd41133, 16'd39045, 16'd16360, 16'd40301, 16'd26598, 16'd38671, 16'd56439, 16'd7111, 16'd18571, 16'd7283, 16'd18252, 16'd29941, 16'd59912, 16'd62624, 16'd57987, 16'd1379, 16'd60967});
	test_expansion(128'h309f4ab192774807f3f98d010bdad29e, {16'd912, 16'd1940, 16'd55469, 16'd21814, 16'd58932, 16'd42775, 16'd38976, 16'd29602, 16'd60122, 16'd54327, 16'd25126, 16'd30461, 16'd38812, 16'd32390, 16'd31337, 16'd12292, 16'd6418, 16'd26612, 16'd38740, 16'd36276, 16'd1665, 16'd55617, 16'd55929, 16'd51347, 16'd24442, 16'd35954});
	test_expansion(128'hebb989082bdc76f84513f68d81e3bc92, {16'd64641, 16'd38644, 16'd6073, 16'd53584, 16'd46071, 16'd31896, 16'd27022, 16'd39530, 16'd23583, 16'd19924, 16'd38288, 16'd40689, 16'd40743, 16'd39232, 16'd38026, 16'd5752, 16'd1372, 16'd4675, 16'd62038, 16'd14022, 16'd60917, 16'd41914, 16'd16768, 16'd15053, 16'd59792, 16'd33803});
	test_expansion(128'h192198b3e5715d5ae0e8a6ab23ae26e7, {16'd39292, 16'd22960, 16'd63819, 16'd31678, 16'd10801, 16'd25434, 16'd27888, 16'd37549, 16'd37738, 16'd33788, 16'd896, 16'd881, 16'd7648, 16'd12549, 16'd2501, 16'd59080, 16'd46827, 16'd49276, 16'd22951, 16'd15652, 16'd52879, 16'd61301, 16'd61811, 16'd2403, 16'd39537, 16'd49445});
	test_expansion(128'haf4c29fe2e102cfad20cc65855a493c5, {16'd63913, 16'd38948, 16'd38364, 16'd30459, 16'd61702, 16'd28241, 16'd41422, 16'd25736, 16'd24548, 16'd45892, 16'd48308, 16'd2277, 16'd47390, 16'd29113, 16'd21454, 16'd28491, 16'd9536, 16'd12122, 16'd30659, 16'd61211, 16'd31994, 16'd4179, 16'd54979, 16'd38604, 16'd47793, 16'd62764});
	test_expansion(128'hc6256ebdb6290aca9dee3381a76c2903, {16'd7398, 16'd54707, 16'd7459, 16'd45763, 16'd12334, 16'd6070, 16'd26063, 16'd34016, 16'd22972, 16'd38692, 16'd29602, 16'd2235, 16'd54890, 16'd61452, 16'd32113, 16'd7294, 16'd47459, 16'd6468, 16'd1553, 16'd1058, 16'd5986, 16'd6877, 16'd31904, 16'd63565, 16'd65055, 16'd14182});
	test_expansion(128'h53dc971535aaf0961b7da66d831ef064, {16'd33792, 16'd31966, 16'd41118, 16'd10394, 16'd61746, 16'd10696, 16'd38651, 16'd31189, 16'd63986, 16'd45904, 16'd18468, 16'd576, 16'd54347, 16'd34085, 16'd34125, 16'd10592, 16'd55442, 16'd37015, 16'd22283, 16'd28323, 16'd4787, 16'd17492, 16'd34533, 16'd37587, 16'd46949, 16'd16654});
	test_expansion(128'hf199dba67b9f90521fe792ebd17e93e0, {16'd36082, 16'd16282, 16'd65178, 16'd16251, 16'd19608, 16'd3329, 16'd30649, 16'd58498, 16'd61991, 16'd61461, 16'd18254, 16'd63452, 16'd62170, 16'd14130, 16'd32146, 16'd18009, 16'd34778, 16'd1914, 16'd24328, 16'd63211, 16'd47401, 16'd6051, 16'd38582, 16'd45238, 16'd52358, 16'd40299});
	test_expansion(128'h6f9260eb90c103bdc249c0e368de884b, {16'd58966, 16'd23911, 16'd50913, 16'd45066, 16'd14085, 16'd42575, 16'd50976, 16'd19028, 16'd30709, 16'd49261, 16'd11874, 16'd37564, 16'd27743, 16'd12539, 16'd39431, 16'd8673, 16'd65356, 16'd35442, 16'd8830, 16'd37835, 16'd47870, 16'd34746, 16'd62085, 16'd56432, 16'd37553, 16'd37303});
	test_expansion(128'h5419d3c382a4fc534be10d7842e5a5a1, {16'd47840, 16'd16848, 16'd40513, 16'd40841, 16'd5899, 16'd41381, 16'd38988, 16'd44751, 16'd46395, 16'd61493, 16'd7221, 16'd21363, 16'd50406, 16'd36391, 16'd27016, 16'd48164, 16'd63833, 16'd56820, 16'd18491, 16'd62584, 16'd33092, 16'd21428, 16'd31792, 16'd26342, 16'd45619, 16'd8413});
	test_expansion(128'he000e42ab28f15fe17abcfdcda74982e, {16'd6080, 16'd31622, 16'd5520, 16'd49809, 16'd47454, 16'd58670, 16'd5693, 16'd61274, 16'd37409, 16'd18310, 16'd2067, 16'd35262, 16'd51881, 16'd59794, 16'd60306, 16'd50345, 16'd44380, 16'd19762, 16'd26332, 16'd65108, 16'd1802, 16'd29000, 16'd55248, 16'd50307, 16'd2385, 16'd20176});
	test_expansion(128'h5cb43bf9d9cffedd63296217f11d697e, {16'd3525, 16'd12015, 16'd65067, 16'd38310, 16'd57070, 16'd8631, 16'd3852, 16'd21883, 16'd10997, 16'd31137, 16'd15288, 16'd22850, 16'd56874, 16'd21114, 16'd50518, 16'd24940, 16'd38609, 16'd24100, 16'd6777, 16'd17904, 16'd9020, 16'd6093, 16'd10181, 16'd47524, 16'd45178, 16'd43029});
	test_expansion(128'h6fa5654e5d32a618d46ecbacf2493c67, {16'd1017, 16'd41525, 16'd36533, 16'd36231, 16'd36344, 16'd20294, 16'd7278, 16'd60632, 16'd56583, 16'd36247, 16'd50412, 16'd36816, 16'd20542, 16'd27719, 16'd56931, 16'd5385, 16'd24904, 16'd9885, 16'd32699, 16'd57419, 16'd8047, 16'd4828, 16'd4056, 16'd8515, 16'd31345, 16'd51700});
	test_expansion(128'h6f4f9a54e1a64ff09f3c36af737b8ec8, {16'd57919, 16'd26805, 16'd26894, 16'd46469, 16'd11223, 16'd39034, 16'd22358, 16'd25431, 16'd47182, 16'd15080, 16'd44822, 16'd39552, 16'd58872, 16'd33621, 16'd23917, 16'd30270, 16'd61287, 16'd50188, 16'd54419, 16'd44863, 16'd63059, 16'd50307, 16'd27052, 16'd53078, 16'd36136, 16'd50080});
	test_expansion(128'hf4cfd33b30c12b5dcea8befacf9c0e31, {16'd20896, 16'd59991, 16'd13289, 16'd55164, 16'd61127, 16'd49193, 16'd9574, 16'd50852, 16'd45199, 16'd9892, 16'd54074, 16'd6228, 16'd55564, 16'd31835, 16'd12261, 16'd20887, 16'd54812, 16'd31691, 16'd17648, 16'd33221, 16'd45218, 16'd21090, 16'd19115, 16'd44724, 16'd17772, 16'd3851});
	test_expansion(128'h835fc7c3c35782172678f4cdc1bcfb08, {16'd38633, 16'd60956, 16'd26332, 16'd50182, 16'd29312, 16'd9750, 16'd1844, 16'd35065, 16'd27661, 16'd62721, 16'd35515, 16'd50997, 16'd58569, 16'd41697, 16'd62226, 16'd61716, 16'd20832, 16'd60238, 16'd33425, 16'd13056, 16'd18921, 16'd41551, 16'd2747, 16'd37246, 16'd40124, 16'd47288});
	test_expansion(128'ha1b9829604e98394d5c361e1fadbe25c, {16'd64562, 16'd59606, 16'd16381, 16'd55360, 16'd49687, 16'd3397, 16'd12598, 16'd48714, 16'd33375, 16'd57899, 16'd29552, 16'd16748, 16'd55638, 16'd1596, 16'd42718, 16'd5915, 16'd48790, 16'd8225, 16'd22110, 16'd36703, 16'd51721, 16'd15652, 16'd57270, 16'd22300, 16'd52233, 16'd23270});
	test_expansion(128'hc9b067a0b8033b788ceab96369ee9cfe, {16'd11459, 16'd25626, 16'd51923, 16'd39958, 16'd43298, 16'd39207, 16'd49939, 16'd4220, 16'd53588, 16'd63317, 16'd54566, 16'd43769, 16'd15716, 16'd40302, 16'd19617, 16'd47799, 16'd39190, 16'd44813, 16'd40774, 16'd10648, 16'd18396, 16'd54246, 16'd65404, 16'd10978, 16'd47986, 16'd59560});
	test_expansion(128'h084c1c901f0231ba9435e83223163b11, {16'd38991, 16'd19140, 16'd20470, 16'd41120, 16'd52689, 16'd36385, 16'd34697, 16'd46914, 16'd9242, 16'd832, 16'd28189, 16'd33710, 16'd44498, 16'd42165, 16'd56957, 16'd47208, 16'd31705, 16'd2802, 16'd19449, 16'd55915, 16'd55202, 16'd26115, 16'd20816, 16'd62581, 16'd28137, 16'd19621});
	test_expansion(128'h36e198ed72bca8b0e1584b4b76d193fe, {16'd33732, 16'd47440, 16'd15322, 16'd28217, 16'd9399, 16'd48813, 16'd47225, 16'd51084, 16'd52205, 16'd36513, 16'd33137, 16'd58769, 16'd42552, 16'd22927, 16'd46279, 16'd28901, 16'd46470, 16'd3896, 16'd39076, 16'd10659, 16'd22479, 16'd61047, 16'd61451, 16'd45207, 16'd59492, 16'd11808});
	test_expansion(128'h6f4650edab276a061512c6efafafc95a, {16'd53378, 16'd51087, 16'd21920, 16'd32724, 16'd5844, 16'd42522, 16'd20722, 16'd52984, 16'd44004, 16'd10981, 16'd37407, 16'd60676, 16'd29593, 16'd42272, 16'd3676, 16'd35587, 16'd64648, 16'd54221, 16'd5070, 16'd54469, 16'd53461, 16'd47689, 16'd6305, 16'd38132, 16'd34467, 16'd44825});
	test_expansion(128'hcd5c81c59910054823dfe4c05a9c1c66, {16'd18516, 16'd48287, 16'd54328, 16'd30954, 16'd45355, 16'd50947, 16'd28128, 16'd12123, 16'd2566, 16'd17052, 16'd54745, 16'd7988, 16'd40006, 16'd6680, 16'd31188, 16'd4602, 16'd49171, 16'd8581, 16'd14697, 16'd15974, 16'd43813, 16'd11982, 16'd2064, 16'd31027, 16'd33751, 16'd30142});
	test_expansion(128'h4056f66ceaecb1abad5d67794314915c, {16'd38243, 16'd29713, 16'd6537, 16'd55799, 16'd54562, 16'd7196, 16'd17905, 16'd52320, 16'd58313, 16'd26267, 16'd739, 16'd4385, 16'd1560, 16'd63641, 16'd64919, 16'd47091, 16'd59865, 16'd19162, 16'd2857, 16'd2868, 16'd37299, 16'd33610, 16'd20806, 16'd6197, 16'd46706, 16'd51541});
	test_expansion(128'h05cb493e06130127e45c9db458de19ea, {16'd17094, 16'd41474, 16'd53169, 16'd37587, 16'd59133, 16'd40135, 16'd49911, 16'd27043, 16'd29536, 16'd40936, 16'd57541, 16'd41750, 16'd30264, 16'd29162, 16'd7855, 16'd33817, 16'd24966, 16'd58283, 16'd39938, 16'd31722, 16'd1841, 16'd36391, 16'd63232, 16'd33654, 16'd15398, 16'd57741});
	test_expansion(128'ha6ccabd0688ccf05b833e8e829445f6c, {16'd27925, 16'd60209, 16'd27629, 16'd13177, 16'd8229, 16'd45287, 16'd64920, 16'd64797, 16'd1067, 16'd30746, 16'd64501, 16'd55209, 16'd65528, 16'd54708, 16'd27562, 16'd40917, 16'd42806, 16'd51623, 16'd62552, 16'd27028, 16'd60903, 16'd28687, 16'd39583, 16'd5303, 16'd11810, 16'd6749});
	test_expansion(128'h8a5c84f27ab9a5245ae22ffdb6a74bca, {16'd62934, 16'd6453, 16'd20740, 16'd48651, 16'd64046, 16'd6412, 16'd4228, 16'd27734, 16'd13668, 16'd40691, 16'd34555, 16'd56279, 16'd46397, 16'd58387, 16'd5395, 16'd19923, 16'd34950, 16'd3304, 16'd6755, 16'd8031, 16'd36051, 16'd34522, 16'd25285, 16'd27341, 16'd9330, 16'd1153});
	test_expansion(128'h3b5ad9424efe1289ebd19d5b7eac6215, {16'd9538, 16'd37085, 16'd60763, 16'd39571, 16'd57402, 16'd43887, 16'd52376, 16'd51551, 16'd28500, 16'd57253, 16'd19869, 16'd40293, 16'd6898, 16'd51316, 16'd35388, 16'd6237, 16'd5112, 16'd10946, 16'd2813, 16'd43971, 16'd48831, 16'd46543, 16'd50438, 16'd26634, 16'd15576, 16'd20007});
	test_expansion(128'hf2d0b541fc896a5c1f467098dc37cc61, {16'd48077, 16'd61822, 16'd20980, 16'd36315, 16'd48702, 16'd60323, 16'd55704, 16'd33956, 16'd65515, 16'd53923, 16'd61550, 16'd15512, 16'd2821, 16'd4625, 16'd20301, 16'd8678, 16'd62106, 16'd56564, 16'd13368, 16'd5328, 16'd51803, 16'd27934, 16'd37137, 16'd8054, 16'd56572, 16'd47814});
	test_expansion(128'hbaacc9583ea7092123b9dd02df2ba040, {16'd40645, 16'd64884, 16'd5510, 16'd45957, 16'd2328, 16'd24571, 16'd28951, 16'd6349, 16'd37575, 16'd35050, 16'd41161, 16'd62401, 16'd1533, 16'd44695, 16'd24097, 16'd38522, 16'd51510, 16'd47983, 16'd1685, 16'd4691, 16'd64764, 16'd59310, 16'd3725, 16'd40142, 16'd23599, 16'd58614});
	test_expansion(128'h92befc42fc2bca000694cfbd815cde04, {16'd50852, 16'd59587, 16'd41179, 16'd32245, 16'd15980, 16'd42253, 16'd12289, 16'd39505, 16'd22802, 16'd49868, 16'd57122, 16'd61262, 16'd63746, 16'd34761, 16'd30581, 16'd12458, 16'd56866, 16'd64787, 16'd12997, 16'd62456, 16'd20692, 16'd60915, 16'd52479, 16'd32825, 16'd63293, 16'd33317});
	test_expansion(128'h24e39f884e13e36dc9f04ceabcce775e, {16'd3813, 16'd15735, 16'd28199, 16'd39980, 16'd8747, 16'd24346, 16'd5583, 16'd27867, 16'd16060, 16'd25445, 16'd16066, 16'd17650, 16'd3744, 16'd100, 16'd65245, 16'd8591, 16'd21388, 16'd25526, 16'd64249, 16'd16213, 16'd17806, 16'd24737, 16'd46878, 16'd21832, 16'd9670, 16'd3709});
	test_expansion(128'h67ba0b1ed66f8227fb241aea1946b745, {16'd58683, 16'd5801, 16'd52445, 16'd16255, 16'd5202, 16'd61326, 16'd52503, 16'd61886, 16'd40911, 16'd38117, 16'd31447, 16'd57239, 16'd29339, 16'd31760, 16'd31056, 16'd55387, 16'd30637, 16'd53391, 16'd13537, 16'd7136, 16'd55093, 16'd8394, 16'd7246, 16'd27852, 16'd23316, 16'd54285});
	test_expansion(128'h867096f7a4dcf82f47865ae01475e968, {16'd56769, 16'd60751, 16'd1632, 16'd25157, 16'd20851, 16'd37938, 16'd56211, 16'd13162, 16'd25356, 16'd1609, 16'd34725, 16'd37350, 16'd48520, 16'd7455, 16'd55815, 16'd11296, 16'd29248, 16'd55800, 16'd24451, 16'd31209, 16'd34230, 16'd63637, 16'd59568, 16'd31310, 16'd53509, 16'd11034});
	test_expansion(128'h88dc6658e3f7eece60429902bb1cbb23, {16'd57929, 16'd28789, 16'd2897, 16'd25555, 16'd25673, 16'd9728, 16'd5020, 16'd59777, 16'd54642, 16'd19043, 16'd43818, 16'd42626, 16'd41349, 16'd10314, 16'd1992, 16'd52233, 16'd61876, 16'd61589, 16'd6382, 16'd28670, 16'd39456, 16'd28875, 16'd58331, 16'd5957, 16'd27524, 16'd64860});
	test_expansion(128'h17062dbfd148fc3a838302beeeb4278c, {16'd228, 16'd4213, 16'd20927, 16'd41810, 16'd44388, 16'd25106, 16'd25764, 16'd45233, 16'd11757, 16'd22091, 16'd19684, 16'd36805, 16'd11416, 16'd56676, 16'd25243, 16'd52663, 16'd56091, 16'd37587, 16'd9467, 16'd53045, 16'd47202, 16'd35877, 16'd18885, 16'd34555, 16'd589, 16'd22012});
	test_expansion(128'h9150aadaed7948896772d6cbfc430c04, {16'd36103, 16'd17319, 16'd35598, 16'd31447, 16'd18048, 16'd3677, 16'd21292, 16'd40421, 16'd61059, 16'd7846, 16'd53193, 16'd7705, 16'd18741, 16'd53938, 16'd29109, 16'd5601, 16'd20250, 16'd6351, 16'd34602, 16'd27550, 16'd3383, 16'd39847, 16'd52453, 16'd49309, 16'd63338, 16'd45775});
	test_expansion(128'h710041ce13efcd4264d3c25a02981bd6, {16'd45044, 16'd54427, 16'd18659, 16'd6476, 16'd17059, 16'd15969, 16'd31624, 16'd22045, 16'd43907, 16'd28014, 16'd59719, 16'd7948, 16'd30742, 16'd44103, 16'd55928, 16'd26403, 16'd59171, 16'd52453, 16'd55627, 16'd60784, 16'd32100, 16'd12518, 16'd63320, 16'd21201, 16'd26624, 16'd18606});
	test_expansion(128'hbc98f3ed89845c7959e5bfe484d55344, {16'd56108, 16'd7514, 16'd644, 16'd45320, 16'd955, 16'd42853, 16'd47126, 16'd14358, 16'd51166, 16'd17193, 16'd25335, 16'd64000, 16'd22632, 16'd29419, 16'd39537, 16'd19658, 16'd50620, 16'd11484, 16'd51799, 16'd31442, 16'd13999, 16'd39858, 16'd11856, 16'd35367, 16'd62786, 16'd33979});
	test_expansion(128'h6c2d88a80e501032b31ac8cdaa94d33c, {16'd18747, 16'd57970, 16'd1004, 16'd63126, 16'd62843, 16'd65154, 16'd54336, 16'd360, 16'd37092, 16'd30828, 16'd26445, 16'd31184, 16'd38404, 16'd5887, 16'd4062, 16'd5592, 16'd18324, 16'd6848, 16'd35903, 16'd35405, 16'd40645, 16'd41463, 16'd63594, 16'd29152, 16'd16440, 16'd26553});
	test_expansion(128'h47481d70884bd6cd3622cfd9ccbbfd29, {16'd60276, 16'd47706, 16'd4752, 16'd3282, 16'd59042, 16'd50615, 16'd24159, 16'd59421, 16'd8271, 16'd26631, 16'd37118, 16'd19131, 16'd59158, 16'd51644, 16'd64366, 16'd44776, 16'd26084, 16'd41217, 16'd39570, 16'd45725, 16'd34773, 16'd10842, 16'd42243, 16'd47570, 16'd25757, 16'd27792});
	test_expansion(128'ha35f8aa971cbf27fcaa7e53fd1c08711, {16'd60212, 16'd30308, 16'd58047, 16'd60176, 16'd4030, 16'd47874, 16'd44043, 16'd11810, 16'd34714, 16'd41360, 16'd62936, 16'd3092, 16'd4999, 16'd48420, 16'd5952, 16'd53702, 16'd61173, 16'd2506, 16'd16485, 16'd50776, 16'd34783, 16'd6207, 16'd30535, 16'd33245, 16'd54305, 16'd16395});
	test_expansion(128'h66eca84001382f822cef4187669336e5, {16'd23598, 16'd782, 16'd58009, 16'd46230, 16'd6455, 16'd42241, 16'd45011, 16'd4508, 16'd44671, 16'd46964, 16'd16697, 16'd727, 16'd65211, 16'd57635, 16'd10791, 16'd26804, 16'd45796, 16'd58841, 16'd16222, 16'd26389, 16'd49529, 16'd29422, 16'd14787, 16'd5495, 16'd14156, 16'd2230});
	test_expansion(128'h0d316e8480e659054256037ccd1bab38, {16'd33527, 16'd21756, 16'd23909, 16'd54073, 16'd27092, 16'd11107, 16'd53341, 16'd7194, 16'd43690, 16'd5093, 16'd61919, 16'd26723, 16'd52291, 16'd57191, 16'd46102, 16'd43359, 16'd3595, 16'd18858, 16'd58020, 16'd45341, 16'd47287, 16'd34709, 16'd31779, 16'd15577, 16'd56853, 16'd15017});
	test_expansion(128'ha089f497fd3c6fc69902efaf9f91380c, {16'd209, 16'd30632, 16'd36318, 16'd59592, 16'd90, 16'd34432, 16'd55359, 16'd28719, 16'd42261, 16'd35436, 16'd50548, 16'd32187, 16'd51783, 16'd22313, 16'd60465, 16'd14811, 16'd53524, 16'd31206, 16'd32332, 16'd18878, 16'd12955, 16'd60954, 16'd21904, 16'd4498, 16'd55958, 16'd35895});
	test_expansion(128'hffa27d5df63a896562914e2b1a6a7a81, {16'd42621, 16'd50869, 16'd6987, 16'd43375, 16'd43919, 16'd22020, 16'd19691, 16'd15742, 16'd32253, 16'd16512, 16'd22977, 16'd38019, 16'd37839, 16'd58264, 16'd42504, 16'd18715, 16'd49219, 16'd58027, 16'd60538, 16'd45074, 16'd57186, 16'd49203, 16'd52019, 16'd17207, 16'd54126, 16'd16990});
	test_expansion(128'h2d2a4bd6625dd64d322d036207494298, {16'd4038, 16'd22261, 16'd47802, 16'd49026, 16'd64852, 16'd60350, 16'd51728, 16'd39277, 16'd30974, 16'd58910, 16'd53443, 16'd19260, 16'd35667, 16'd27697, 16'd36045, 16'd21305, 16'd25697, 16'd46750, 16'd14825, 16'd50546, 16'd16717, 16'd44234, 16'd57953, 16'd8137, 16'd60246, 16'd41380});
	test_expansion(128'hc011508e8065fd3a8aa097cf31e03cea, {16'd5877, 16'd30899, 16'd46295, 16'd63670, 16'd10965, 16'd3564, 16'd32469, 16'd45357, 16'd46827, 16'd35716, 16'd6087, 16'd16460, 16'd32654, 16'd55334, 16'd8875, 16'd21010, 16'd57433, 16'd18002, 16'd29088, 16'd53753, 16'd3876, 16'd24045, 16'd32695, 16'd53978, 16'd60114, 16'd63654});
	test_expansion(128'hb169619845cc1fd3f7699d0533a20f03, {16'd4339, 16'd6902, 16'd34008, 16'd54230, 16'd14490, 16'd38569, 16'd12860, 16'd64791, 16'd10675, 16'd33546, 16'd28434, 16'd54567, 16'd60094, 16'd31084, 16'd20410, 16'd31688, 16'd7738, 16'd1049, 16'd16562, 16'd46750, 16'd46690, 16'd6703, 16'd33410, 16'd55133, 16'd20420, 16'd21001});
	test_expansion(128'h1ff480beb245bf37e4257693d5794d06, {16'd18792, 16'd58189, 16'd15925, 16'd37605, 16'd62409, 16'd2255, 16'd25705, 16'd38921, 16'd31932, 16'd57403, 16'd4404, 16'd53065, 16'd60192, 16'd15250, 16'd11209, 16'd51989, 16'd6113, 16'd31758, 16'd34265, 16'd14537, 16'd5508, 16'd1816, 16'd21327, 16'd7390, 16'd27146, 16'd53614});
	test_expansion(128'ha9087050a698d779ca22ece6a3cf60c6, {16'd47642, 16'd16305, 16'd15988, 16'd4902, 16'd42920, 16'd28800, 16'd62931, 16'd20454, 16'd15678, 16'd10720, 16'd43269, 16'd63349, 16'd12098, 16'd11081, 16'd23790, 16'd47739, 16'd622, 16'd20957, 16'd26245, 16'd49637, 16'd4621, 16'd34584, 16'd55750, 16'd56955, 16'd3793, 16'd60954});
	test_expansion(128'h90b751f0d012aeb61afc8e1e753c6767, {16'd45418, 16'd26245, 16'd41783, 16'd29126, 16'd4842, 16'd50148, 16'd63239, 16'd43262, 16'd28032, 16'd30639, 16'd13459, 16'd53365, 16'd47505, 16'd50197, 16'd9749, 16'd132, 16'd36704, 16'd48636, 16'd57204, 16'd20515, 16'd33071, 16'd58543, 16'd20462, 16'd64787, 16'd14521, 16'd3637});
	test_expansion(128'h52b2f962432c0d98d22bc77c105527a1, {16'd27323, 16'd31523, 16'd59459, 16'd40794, 16'd39876, 16'd41424, 16'd10893, 16'd16395, 16'd22819, 16'd58390, 16'd53773, 16'd63541, 16'd45854, 16'd18778, 16'd21425, 16'd14753, 16'd58957, 16'd53279, 16'd33848, 16'd17981, 16'd25815, 16'd53272, 16'd40036, 16'd40429, 16'd10067, 16'd24299});
	test_expansion(128'h37a170d1f64e0b0996213750456c9413, {16'd4639, 16'd29663, 16'd18668, 16'd59519, 16'd53054, 16'd57164, 16'd41330, 16'd59100, 16'd12997, 16'd22534, 16'd33619, 16'd51421, 16'd30446, 16'd54370, 16'd43859, 16'd56179, 16'd8862, 16'd20277, 16'd64934, 16'd49778, 16'd36009, 16'd58800, 16'd18890, 16'd28483, 16'd27511, 16'd2213});
	test_expansion(128'ha445448bc00894489b00b15caf48a2ec, {16'd45365, 16'd29746, 16'd52486, 16'd65269, 16'd18833, 16'd242, 16'd5397, 16'd49263, 16'd19043, 16'd48217, 16'd55416, 16'd64458, 16'd38940, 16'd52461, 16'd10782, 16'd29528, 16'd1215, 16'd40485, 16'd35638, 16'd51449, 16'd63092, 16'd45907, 16'd61281, 16'd47395, 16'd24994, 16'd20776});
	test_expansion(128'hc62251b3fda79ba39d956fb1e894b2a4, {16'd96, 16'd42659, 16'd678, 16'd28100, 16'd25093, 16'd20835, 16'd53576, 16'd46314, 16'd64828, 16'd33734, 16'd17275, 16'd35532, 16'd64645, 16'd5906, 16'd49442, 16'd26157, 16'd42372, 16'd65305, 16'd28028, 16'd60861, 16'd53377, 16'd36728, 16'd8022, 16'd54708, 16'd3699, 16'd42481});
	test_expansion(128'h9dfd4f3668fcc35d82380a86bb6ac427, {16'd48046, 16'd41409, 16'd62071, 16'd33223, 16'd16254, 16'd41670, 16'd16374, 16'd53808, 16'd51844, 16'd15569, 16'd19473, 16'd11558, 16'd21046, 16'd47620, 16'd55753, 16'd41316, 16'd5998, 16'd42357, 16'd57117, 16'd9795, 16'd49121, 16'd19941, 16'd8999, 16'd6216, 16'd21883, 16'd51336});
	test_expansion(128'h77e5da42c785128d3f81e9783af4ce46, {16'd8166, 16'd31623, 16'd9631, 16'd58634, 16'd640, 16'd42474, 16'd19497, 16'd41093, 16'd50177, 16'd5217, 16'd49351, 16'd57044, 16'd44547, 16'd2159, 16'd55770, 16'd8251, 16'd28293, 16'd30602, 16'd18411, 16'd64634, 16'd38729, 16'd38666, 16'd20535, 16'd18393, 16'd10253, 16'd7708});
	test_expansion(128'h5ee87c52724654b67d4e86f1b65153aa, {16'd6575, 16'd11705, 16'd14903, 16'd9619, 16'd34493, 16'd32490, 16'd29710, 16'd38819, 16'd50341, 16'd26682, 16'd61894, 16'd40417, 16'd26840, 16'd51275, 16'd49395, 16'd59131, 16'd36582, 16'd45128, 16'd37882, 16'd38109, 16'd58897, 16'd31511, 16'd51003, 16'd12510, 16'd54585, 16'd30929});
	test_expansion(128'hfae60d01f480e88e5d57f326e6081791, {16'd64846, 16'd31766, 16'd3942, 16'd21487, 16'd46753, 16'd61287, 16'd359, 16'd4477, 16'd21358, 16'd8317, 16'd65006, 16'd28104, 16'd58503, 16'd7727, 16'd41354, 16'd49781, 16'd31807, 16'd11608, 16'd28856, 16'd17932, 16'd46395, 16'd31435, 16'd34629, 16'd36818, 16'd11326, 16'd15565});
	test_expansion(128'h91b798dfaaf805c88eadd3ba604f6e00, {16'd38254, 16'd18858, 16'd21261, 16'd9065, 16'd48248, 16'd28009, 16'd29854, 16'd35745, 16'd1188, 16'd64177, 16'd8494, 16'd13383, 16'd46232, 16'd39845, 16'd52888, 16'd16589, 16'd23404, 16'd40838, 16'd18084, 16'd21904, 16'd38741, 16'd17156, 16'd59920, 16'd21907, 16'd14743, 16'd27713});
	test_expansion(128'h99936b9742ea4c72ae144cdc9dd2bbeb, {16'd32742, 16'd31531, 16'd516, 16'd23749, 16'd50060, 16'd16326, 16'd18531, 16'd13008, 16'd54051, 16'd5305, 16'd50366, 16'd22435, 16'd42081, 16'd29705, 16'd3500, 16'd16382, 16'd12314, 16'd42851, 16'd48839, 16'd45250, 16'd44369, 16'd60057, 16'd3433, 16'd7019, 16'd40112, 16'd18006});
	test_expansion(128'haf12560e803c49ac6077b5907942d3f9, {16'd39994, 16'd27455, 16'd11523, 16'd2278, 16'd1581, 16'd27174, 16'd25060, 16'd34094, 16'd58487, 16'd37482, 16'd29960, 16'd9294, 16'd44609, 16'd12166, 16'd55800, 16'd15392, 16'd34351, 16'd54004, 16'd46273, 16'd52976, 16'd23778, 16'd13612, 16'd3938, 16'd24974, 16'd27734, 16'd41550});
	test_expansion(128'he01eef63d0bb1c368398c1abc14d00aa, {16'd64134, 16'd56921, 16'd40039, 16'd6522, 16'd9351, 16'd31669, 16'd63250, 16'd15296, 16'd56601, 16'd51839, 16'd37307, 16'd54257, 16'd3663, 16'd58463, 16'd63911, 16'd53815, 16'd43756, 16'd52107, 16'd21952, 16'd14338, 16'd54575, 16'd49868, 16'd63897, 16'd36593, 16'd49552, 16'd33036});
	test_expansion(128'h422cc6774d3470799e917da2c8b9a649, {16'd43962, 16'd607, 16'd9061, 16'd12812, 16'd42223, 16'd19632, 16'd44506, 16'd24393, 16'd41425, 16'd52618, 16'd61158, 16'd10292, 16'd62640, 16'd17793, 16'd48264, 16'd31207, 16'd21457, 16'd5250, 16'd29956, 16'd13419, 16'd54714, 16'd277, 16'd5188, 16'd42990, 16'd62189, 16'd36783});
	test_expansion(128'h025354ef2c4906387eb171ecfa81d9e7, {16'd27118, 16'd8112, 16'd62108, 16'd10135, 16'd26808, 16'd36245, 16'd46375, 16'd59017, 16'd14259, 16'd35561, 16'd5906, 16'd12746, 16'd52496, 16'd8095, 16'd28046, 16'd30844, 16'd3240, 16'd13435, 16'd30020, 16'd40948, 16'd58023, 16'd41241, 16'd50164, 16'd4890, 16'd31129, 16'd59627});
	test_expansion(128'h66d6dfdf01e4110f3924f4139e5d4e0a, {16'd47557, 16'd40313, 16'd34008, 16'd977, 16'd16587, 16'd30467, 16'd43303, 16'd44004, 16'd19431, 16'd59376, 16'd38201, 16'd3964, 16'd7888, 16'd19635, 16'd41264, 16'd24223, 16'd64711, 16'd22455, 16'd1049, 16'd13938, 16'd1602, 16'd52804, 16'd24534, 16'd1827, 16'd2200, 16'd56289});
	test_expansion(128'h0e0ed05fbe9596cb8d65ed46470f21f8, {16'd44405, 16'd65514, 16'd35656, 16'd46469, 16'd875, 16'd23175, 16'd17791, 16'd43209, 16'd27965, 16'd10252, 16'd58340, 16'd57338, 16'd20658, 16'd7744, 16'd14323, 16'd51634, 16'd38642, 16'd35514, 16'd19787, 16'd31295, 16'd30848, 16'd46013, 16'd54401, 16'd58969, 16'd52455, 16'd29039});
	test_expansion(128'h202d1918561cacfa6a43c00cd987d375, {16'd64021, 16'd34727, 16'd47195, 16'd9496, 16'd6065, 16'd9339, 16'd29674, 16'd32890, 16'd2930, 16'd45479, 16'd23525, 16'd27085, 16'd36575, 16'd48040, 16'd34275, 16'd44640, 16'd61392, 16'd8261, 16'd11019, 16'd58390, 16'd29014, 16'd38384, 16'd26619, 16'd62421, 16'd46811, 16'd41894});
	test_expansion(128'h74129d832036fd4929436d569f42c92f, {16'd36475, 16'd49232, 16'd1860, 16'd39628, 16'd7849, 16'd45511, 16'd56153, 16'd36201, 16'd15664, 16'd34415, 16'd35923, 16'd55448, 16'd42870, 16'd48708, 16'd4184, 16'd56101, 16'd60497, 16'd35095, 16'd25786, 16'd11672, 16'd17866, 16'd63797, 16'd63304, 16'd48273, 16'd26727, 16'd39342});
	test_expansion(128'h7a6b9a8cae32706ae013c8541fd6645f, {16'd54959, 16'd28099, 16'd30448, 16'd60667, 16'd55947, 16'd20758, 16'd25144, 16'd56342, 16'd59101, 16'd27954, 16'd28244, 16'd36907, 16'd48791, 16'd18369, 16'd44008, 16'd58644, 16'd45324, 16'd36972, 16'd33267, 16'd50421, 16'd33498, 16'd7678, 16'd57830, 16'd10311, 16'd15595, 16'd60034});
	test_expansion(128'h6fa4b23c01fda6f105ae701dc11e3b15, {16'd17963, 16'd31028, 16'd29792, 16'd55685, 16'd38864, 16'd29593, 16'd20762, 16'd16232, 16'd56012, 16'd5485, 16'd51926, 16'd11304, 16'd49161, 16'd50515, 16'd15129, 16'd62552, 16'd24041, 16'd54966, 16'd5050, 16'd57624, 16'd65274, 16'd25772, 16'd43532, 16'd59644, 16'd54413, 16'd50897});
	test_expansion(128'h08389b043e5a7c6771780e15548cad1e, {16'd49751, 16'd28494, 16'd59218, 16'd20130, 16'd45238, 16'd53102, 16'd45259, 16'd30830, 16'd56372, 16'd47144, 16'd49734, 16'd41317, 16'd46972, 16'd45668, 16'd62347, 16'd47935, 16'd43729, 16'd55089, 16'd47819, 16'd52248, 16'd29690, 16'd60093, 16'd31294, 16'd29963, 16'd15956, 16'd37132});
	test_expansion(128'h0b3ceb34415a40f674788066a328c709, {16'd3923, 16'd54948, 16'd11211, 16'd19169, 16'd14537, 16'd60736, 16'd64046, 16'd3895, 16'd11818, 16'd64638, 16'd36022, 16'd39084, 16'd27743, 16'd5858, 16'd46294, 16'd23718, 16'd2419, 16'd34401, 16'd54747, 16'd33050, 16'd30527, 16'd30866, 16'd47693, 16'd20587, 16'd58634, 16'd23476});
	test_expansion(128'h412133ec1d5551e34ea316a5bc0db112, {16'd38436, 16'd20304, 16'd18984, 16'd44332, 16'd44201, 16'd14383, 16'd52291, 16'd49093, 16'd16275, 16'd13773, 16'd1034, 16'd58029, 16'd36961, 16'd3927, 16'd48398, 16'd61062, 16'd51243, 16'd48487, 16'd11591, 16'd29474, 16'd50654, 16'd10400, 16'd7861, 16'd8741, 16'd62854, 16'd48894});
	test_expansion(128'h76f3b6a7576b4103f1afbcd99138ddb9, {16'd24547, 16'd51524, 16'd25748, 16'd50634, 16'd51488, 16'd4178, 16'd62831, 16'd31588, 16'd10256, 16'd33028, 16'd15079, 16'd26795, 16'd38443, 16'd14403, 16'd15782, 16'd57260, 16'd37748, 16'd3692, 16'd25040, 16'd21171, 16'd43735, 16'd26638, 16'd9477, 16'd34475, 16'd5834, 16'd24223});
	test_expansion(128'h9a1e102655295c93cce7e41adddc7b0d, {16'd25794, 16'd5915, 16'd35, 16'd32611, 16'd63418, 16'd51542, 16'd26604, 16'd44317, 16'd20932, 16'd42116, 16'd39548, 16'd12683, 16'd34614, 16'd26104, 16'd47509, 16'd13804, 16'd48152, 16'd14746, 16'd30653, 16'd24831, 16'd5786, 16'd55614, 16'd34169, 16'd63548, 16'd30002, 16'd336});
	test_expansion(128'h81b4fbf6a0179ef5e48b3185e8d078b9, {16'd45835, 16'd41923, 16'd9541, 16'd56400, 16'd6318, 16'd54537, 16'd33986, 16'd7153, 16'd62028, 16'd57893, 16'd25239, 16'd27482, 16'd52284, 16'd19768, 16'd57297, 16'd2574, 16'd47725, 16'd18640, 16'd41563, 16'd57751, 16'd47656, 16'd571, 16'd45814, 16'd7239, 16'd34929, 16'd36412});
	test_expansion(128'h0ecf69a46a20d9a371fd9cf8ca208cd1, {16'd22711, 16'd60173, 16'd14302, 16'd24888, 16'd11790, 16'd42547, 16'd34416, 16'd11221, 16'd63317, 16'd4334, 16'd41252, 16'd4426, 16'd12029, 16'd13948, 16'd16354, 16'd18856, 16'd11571, 16'd25340, 16'd63192, 16'd19012, 16'd61115, 16'd39707, 16'd14739, 16'd52452, 16'd30794, 16'd40064});
	test_expansion(128'h0526ea2c4cada66b111590ad870aa46f, {16'd55127, 16'd58935, 16'd53016, 16'd55040, 16'd30370, 16'd57761, 16'd60149, 16'd945, 16'd28867, 16'd20223, 16'd42821, 16'd14993, 16'd43957, 16'd58695, 16'd53292, 16'd59786, 16'd43803, 16'd34307, 16'd48416, 16'd31066, 16'd39528, 16'd22316, 16'd18339, 16'd5580, 16'd63178, 16'd7229});
	test_expansion(128'h7cf3ec87122d78573824911ea1cb5ae5, {16'd8253, 16'd9651, 16'd12657, 16'd28151, 16'd30370, 16'd35656, 16'd22456, 16'd22286, 16'd37314, 16'd381, 16'd38728, 16'd51099, 16'd63599, 16'd29468, 16'd27792, 16'd44723, 16'd54240, 16'd27463, 16'd57547, 16'd27125, 16'd13478, 16'd7170, 16'd53242, 16'd36903, 16'd8550, 16'd11809});
	test_expansion(128'hc233c35c27f63ab4d7a73bbdeb38728e, {16'd38439, 16'd26104, 16'd57891, 16'd59082, 16'd25005, 16'd29438, 16'd65060, 16'd8695, 16'd39344, 16'd60541, 16'd8172, 16'd42586, 16'd44123, 16'd15884, 16'd29617, 16'd38689, 16'd60726, 16'd58936, 16'd34519, 16'd42760, 16'd22485, 16'd47565, 16'd43785, 16'd15161, 16'd56196, 16'd58495});
	test_expansion(128'hb838ec4b1baa1786190e0524cfcef53d, {16'd35372, 16'd58474, 16'd36209, 16'd37796, 16'd16093, 16'd65082, 16'd14573, 16'd32484, 16'd18029, 16'd1477, 16'd8749, 16'd42562, 16'd25862, 16'd65214, 16'd19935, 16'd30808, 16'd33587, 16'd27529, 16'd47319, 16'd54618, 16'd42613, 16'd14740, 16'd30291, 16'd32595, 16'd45978, 16'd11695});
	test_expansion(128'h97dc3275966526243d4a85c8dd4b3673, {16'd30094, 16'd58237, 16'd40566, 16'd55064, 16'd19743, 16'd25825, 16'd14501, 16'd23514, 16'd24137, 16'd45378, 16'd39868, 16'd23546, 16'd14458, 16'd9834, 16'd14362, 16'd64210, 16'd16185, 16'd44948, 16'd57794, 16'd46365, 16'd61460, 16'd4448, 16'd12498, 16'd249, 16'd53249, 16'd13753});
	test_expansion(128'h25c7f83ab80e7554486c134a0f6db684, {16'd10949, 16'd34522, 16'd35172, 16'd62270, 16'd45079, 16'd57096, 16'd31976, 16'd63588, 16'd17594, 16'd13903, 16'd52778, 16'd57732, 16'd63024, 16'd53854, 16'd52436, 16'd9851, 16'd52559, 16'd1761, 16'd9642, 16'd9383, 16'd24901, 16'd65298, 16'd2164, 16'd26833, 16'd32765, 16'd47443});
	test_expansion(128'h5fecdc35abb9139df583c298b1149191, {16'd41739, 16'd45860, 16'd25737, 16'd55559, 16'd32379, 16'd18049, 16'd30701, 16'd42372, 16'd18743, 16'd31711, 16'd54199, 16'd48589, 16'd62283, 16'd9135, 16'd6642, 16'd15156, 16'd37589, 16'd58589, 16'd60458, 16'd45778, 16'd37323, 16'd55913, 16'd34428, 16'd14412, 16'd64669, 16'd25425});
	test_expansion(128'hb0abd09283104e5e7dace1e08eadc6e8, {16'd51336, 16'd30462, 16'd31491, 16'd55578, 16'd50742, 16'd56919, 16'd40088, 16'd61863, 16'd30064, 16'd37306, 16'd7365, 16'd37476, 16'd54694, 16'd36510, 16'd30808, 16'd39326, 16'd5995, 16'd29595, 16'd60671, 16'd616, 16'd47779, 16'd61451, 16'd22905, 16'd41063, 16'd53654, 16'd194});
	test_expansion(128'h2a794a687f1eb137611f41edb74afdfb, {16'd11231, 16'd4274, 16'd22893, 16'd16478, 16'd6303, 16'd50419, 16'd26185, 16'd52817, 16'd31004, 16'd15960, 16'd34139, 16'd58883, 16'd1297, 16'd23307, 16'd9951, 16'd33587, 16'd36711, 16'd26874, 16'd4273, 16'd34981, 16'd7281, 16'd52588, 16'd21479, 16'd42783, 16'd8080, 16'd52550});
	test_expansion(128'hb99279b1aa5641b7ea0bec98be79832f, {16'd26208, 16'd44904, 16'd60603, 16'd7115, 16'd64417, 16'd48936, 16'd19009, 16'd36478, 16'd60712, 16'd17732, 16'd30800, 16'd32374, 16'd8128, 16'd12952, 16'd40073, 16'd48083, 16'd7974, 16'd44298, 16'd50521, 16'd59631, 16'd17647, 16'd3623, 16'd15752, 16'd18813, 16'd16667, 16'd26967});
	test_expansion(128'h67d782c56bfb6805050c6e916f42440a, {16'd24566, 16'd55762, 16'd28640, 16'd52643, 16'd1117, 16'd34931, 16'd39108, 16'd8875, 16'd21390, 16'd51797, 16'd32947, 16'd58330, 16'd18074, 16'd4990, 16'd22851, 16'd17527, 16'd5774, 16'd38019, 16'd7467, 16'd50639, 16'd50954, 16'd46605, 16'd54542, 16'd53580, 16'd40839, 16'd25882});
	test_expansion(128'he74dc6252623e3a5e686286076e5c325, {16'd20739, 16'd20197, 16'd2836, 16'd22764, 16'd51978, 16'd2860, 16'd54044, 16'd63573, 16'd3764, 16'd62147, 16'd40282, 16'd29616, 16'd28691, 16'd37625, 16'd29599, 16'd63992, 16'd45488, 16'd56250, 16'd60829, 16'd1215, 16'd62391, 16'd22453, 16'd5817, 16'd56799, 16'd58059, 16'd38926});
	test_expansion(128'h44eae28b1401cb2539545dd73526876f, {16'd44372, 16'd59879, 16'd14719, 16'd17724, 16'd37326, 16'd20522, 16'd56443, 16'd34595, 16'd2489, 16'd16306, 16'd51669, 16'd8814, 16'd25974, 16'd21863, 16'd3240, 16'd47283, 16'd3537, 16'd45692, 16'd32882, 16'd4329, 16'd34407, 16'd8729, 16'd2659, 16'd64717, 16'd49082, 16'd50694});
	test_expansion(128'h35cccdd82697fc3d1e2b1f35c5a176de, {16'd19186, 16'd57647, 16'd39833, 16'd13279, 16'd41230, 16'd43244, 16'd3229, 16'd58073, 16'd9084, 16'd41355, 16'd48427, 16'd47363, 16'd64830, 16'd56117, 16'd43347, 16'd23153, 16'd25153, 16'd60059, 16'd23834, 16'd57958, 16'd37917, 16'd64443, 16'd25901, 16'd1860, 16'd7707, 16'd8571});
	test_expansion(128'hb94b7b1b3d558580f76566d7880c2fd4, {16'd24814, 16'd43050, 16'd10959, 16'd6648, 16'd11014, 16'd57847, 16'd43207, 16'd57018, 16'd28254, 16'd53203, 16'd45665, 16'd26152, 16'd42135, 16'd54436, 16'd62133, 16'd8134, 16'd27845, 16'd58133, 16'd20004, 16'd8363, 16'd56208, 16'd8090, 16'd51816, 16'd40791, 16'd4739, 16'd12106});
	test_expansion(128'h32abf1e1bda393afc934fa2dd5ea6d3c, {16'd58382, 16'd13622, 16'd16887, 16'd58589, 16'd13080, 16'd22478, 16'd45360, 16'd27695, 16'd40373, 16'd54488, 16'd21188, 16'd43254, 16'd4567, 16'd18153, 16'd32453, 16'd7418, 16'd33702, 16'd8363, 16'd58893, 16'd64975, 16'd35273, 16'd37798, 16'd29960, 16'd28777, 16'd23054, 16'd7343});
	test_expansion(128'h34214af9b1ec716f4d9944e30b6f6935, {16'd50036, 16'd25560, 16'd62662, 16'd2897, 16'd3022, 16'd58040, 16'd21316, 16'd21067, 16'd28555, 16'd38610, 16'd17113, 16'd62931, 16'd8529, 16'd52343, 16'd62131, 16'd31017, 16'd29744, 16'd15042, 16'd7959, 16'd8673, 16'd37713, 16'd43742, 16'd16807, 16'd432, 16'd7466, 16'd47643});
	test_expansion(128'h610f83434738f67745a4f9760e611dc6, {16'd4685, 16'd23602, 16'd40048, 16'd33780, 16'd14641, 16'd26988, 16'd16098, 16'd31832, 16'd51824, 16'd29529, 16'd44731, 16'd55199, 16'd9369, 16'd37971, 16'd57585, 16'd44045, 16'd1815, 16'd4189, 16'd19199, 16'd21482, 16'd36483, 16'd19353, 16'd10974, 16'd737, 16'd52421, 16'd41853});
	test_expansion(128'h8e7e4c86c2fd6ef38f5f3d8c1e1a6770, {16'd14329, 16'd40547, 16'd7262, 16'd2170, 16'd14839, 16'd49189, 16'd23047, 16'd38481, 16'd12585, 16'd56595, 16'd42470, 16'd22628, 16'd52542, 16'd15610, 16'd30201, 16'd1257, 16'd29919, 16'd7136, 16'd45985, 16'd52707, 16'd26501, 16'd45453, 16'd54287, 16'd42793, 16'd2015, 16'd31470});
	test_expansion(128'he630e60ec79a24c19d2e5edf3c60de67, {16'd8465, 16'd32093, 16'd49663, 16'd20573, 16'd36928, 16'd62149, 16'd53747, 16'd63006, 16'd49855, 16'd17805, 16'd10741, 16'd26146, 16'd57782, 16'd45193, 16'd57474, 16'd29331, 16'd13835, 16'd26123, 16'd27696, 16'd54388, 16'd57936, 16'd62897, 16'd22752, 16'd55484, 16'd54253, 16'd57329});
	test_expansion(128'h6297434e84c3ff5de323488276fdd6f8, {16'd15848, 16'd10024, 16'd39275, 16'd37856, 16'd18414, 16'd10136, 16'd59404, 16'd9505, 16'd36057, 16'd62944, 16'd24784, 16'd51993, 16'd43416, 16'd16327, 16'd37866, 16'd38160, 16'd89, 16'd4858, 16'd64924, 16'd40980, 16'd5570, 16'd12967, 16'd28058, 16'd32781, 16'd26598, 16'd14582});
	test_expansion(128'h15fec5f53923269598c50e1f0cdc51d6, {16'd14039, 16'd14899, 16'd384, 16'd23459, 16'd27992, 16'd61234, 16'd43106, 16'd31541, 16'd15383, 16'd40452, 16'd49320, 16'd19304, 16'd51340, 16'd55744, 16'd33439, 16'd22869, 16'd65233, 16'd64624, 16'd9191, 16'd11880, 16'd12680, 16'd14547, 16'd58636, 16'd12164, 16'd138, 16'd63256});
	test_expansion(128'he1f7009a520c20309be70d77f13c228c, {16'd37325, 16'd52713, 16'd21598, 16'd5115, 16'd15175, 16'd51673, 16'd43606, 16'd16450, 16'd61136, 16'd31876, 16'd57378, 16'd7917, 16'd59964, 16'd39231, 16'd26630, 16'd41547, 16'd31940, 16'd151, 16'd20521, 16'd24623, 16'd21722, 16'd14105, 16'd50935, 16'd48088, 16'd3121, 16'd42116});
	test_expansion(128'h0a8cb86017f6f795c875cf52ec912de4, {16'd37295, 16'd29961, 16'd872, 16'd44722, 16'd36488, 16'd31811, 16'd55856, 16'd52062, 16'd12476, 16'd34599, 16'd23183, 16'd14540, 16'd30050, 16'd45873, 16'd11268, 16'd13596, 16'd26767, 16'd37828, 16'd12196, 16'd6233, 16'd15971, 16'd64207, 16'd59167, 16'd13384, 16'd29203, 16'd38690});
	test_expansion(128'h4cb25b77e19d04142483cb517f68e2f5, {16'd46644, 16'd14193, 16'd58953, 16'd5395, 16'd20900, 16'd42936, 16'd12295, 16'd57039, 16'd53293, 16'd33101, 16'd6863, 16'd2285, 16'd50307, 16'd11662, 16'd39828, 16'd25585, 16'd23006, 16'd35471, 16'd230, 16'd19071, 16'd23697, 16'd14656, 16'd9582, 16'd24721, 16'd30686, 16'd39258});
	test_expansion(128'h74f69d819e2b82ff0a2fd75d9ad1774b, {16'd36321, 16'd27186, 16'd10429, 16'd58915, 16'd57229, 16'd29995, 16'd26589, 16'd56975, 16'd38587, 16'd17411, 16'd53749, 16'd62930, 16'd27290, 16'd28159, 16'd47617, 16'd9497, 16'd14261, 16'd35598, 16'd56501, 16'd5942, 16'd30538, 16'd32377, 16'd26180, 16'd29023, 16'd63648, 16'd25969});
	test_expansion(128'h0bb67ffb0dccc29713873d1a83716340, {16'd42461, 16'd36721, 16'd7918, 16'd10664, 16'd53783, 16'd5268, 16'd62259, 16'd6966, 16'd57081, 16'd9773, 16'd52152, 16'd59224, 16'd40496, 16'd1159, 16'd33611, 16'd16629, 16'd59359, 16'd33308, 16'd55986, 16'd23033, 16'd5916, 16'd63427, 16'd35187, 16'd50366, 16'd44468, 16'd62621});
	test_expansion(128'heeab47328fc2671c25a20186bf99f236, {16'd61497, 16'd23149, 16'd60538, 16'd17169, 16'd1452, 16'd14199, 16'd57102, 16'd32475, 16'd55208, 16'd31292, 16'd9869, 16'd48941, 16'd42951, 16'd63544, 16'd24545, 16'd48733, 16'd24569, 16'd33536, 16'd47587, 16'd47726, 16'd56630, 16'd51014, 16'd50506, 16'd54582, 16'd56985, 16'd34064});
	test_expansion(128'h53072cbd1349d2cf5e3392b472ef9d8c, {16'd13275, 16'd40360, 16'd51154, 16'd44303, 16'd60392, 16'd30297, 16'd64975, 16'd32404, 16'd16711, 16'd41069, 16'd35438, 16'd26452, 16'd17369, 16'd37793, 16'd53789, 16'd17699, 16'd50315, 16'd33436, 16'd17831, 16'd20209, 16'd8196, 16'd22350, 16'd51325, 16'd28890, 16'd38331, 16'd37583});
	test_expansion(128'hc164c44bb51ad56c28b4b9074eff8c3e, {16'd14625, 16'd10977, 16'd12830, 16'd31350, 16'd25953, 16'd18041, 16'd24187, 16'd14, 16'd32446, 16'd14269, 16'd61968, 16'd22317, 16'd32224, 16'd20428, 16'd42781, 16'd32450, 16'd48447, 16'd32722, 16'd35904, 16'd29979, 16'd51480, 16'd63053, 16'd50731, 16'd59529, 16'd7976, 16'd12569});
	test_expansion(128'h8a1692e1d895bb3c1b0dfe14438fad2f, {16'd26071, 16'd27744, 16'd60345, 16'd28761, 16'd28116, 16'd39350, 16'd26511, 16'd36366, 16'd8515, 16'd35245, 16'd32643, 16'd62536, 16'd30103, 16'd52641, 16'd1038, 16'd21707, 16'd25464, 16'd61217, 16'd20831, 16'd5012, 16'd44293, 16'd56776, 16'd48861, 16'd52885, 16'd48830, 16'd54994});
	test_expansion(128'h76719f85862de267ac4e27dce09c8df5, {16'd11789, 16'd52637, 16'd32491, 16'd38885, 16'd41076, 16'd60738, 16'd35184, 16'd56083, 16'd45776, 16'd1660, 16'd14908, 16'd18623, 16'd31301, 16'd22616, 16'd32234, 16'd3027, 16'd11381, 16'd59562, 16'd50646, 16'd50605, 16'd11981, 16'd3927, 16'd49220, 16'd44891, 16'd5509, 16'd46507});
	test_expansion(128'h3d5ff25ff2896a47a4097b8ccca4d60b, {16'd30576, 16'd26434, 16'd643, 16'd35106, 16'd15542, 16'd18244, 16'd45665, 16'd43853, 16'd50135, 16'd13316, 16'd64963, 16'd3641, 16'd47815, 16'd62459, 16'd45058, 16'd34170, 16'd1974, 16'd23535, 16'd16261, 16'd2417, 16'd4128, 16'd17786, 16'd3072, 16'd7399, 16'd21878, 16'd39127});
	test_expansion(128'hb3d0eeb5aa069c166d0d1b14adb692fa, {16'd42914, 16'd41769, 16'd56339, 16'd52698, 16'd9908, 16'd11282, 16'd2925, 16'd50057, 16'd58492, 16'd58655, 16'd49079, 16'd35475, 16'd16624, 16'd45695, 16'd49646, 16'd62274, 16'd4731, 16'd8781, 16'd50636, 16'd8263, 16'd60061, 16'd31834, 16'd51359, 16'd52944, 16'd28539, 16'd53950});
	test_expansion(128'h0bd90cadf486ac2616733b0f3985b220, {16'd16261, 16'd27273, 16'd50854, 16'd16066, 16'd64196, 16'd17984, 16'd3775, 16'd19602, 16'd43206, 16'd4516, 16'd28256, 16'd54756, 16'd59878, 16'd49787, 16'd25389, 16'd45491, 16'd57241, 16'd46542, 16'd17227, 16'd55926, 16'd63984, 16'd15616, 16'd45311, 16'd35085, 16'd58932, 16'd31902});
	test_expansion(128'h63c60b33d66a125981727fa03f6b4a01, {16'd31890, 16'd8560, 16'd31300, 16'd21179, 16'd55220, 16'd22601, 16'd16241, 16'd42107, 16'd32841, 16'd7504, 16'd39940, 16'd52666, 16'd25914, 16'd52653, 16'd12489, 16'd5144, 16'd46982, 16'd4215, 16'd53928, 16'd60158, 16'd23894, 16'd61153, 16'd43821, 16'd521, 16'd65303, 16'd17869});
	test_expansion(128'h958820bf4ed434e9a1531392dcab9c14, {16'd32633, 16'd35315, 16'd741, 16'd24168, 16'd62774, 16'd30622, 16'd25735, 16'd65230, 16'd33788, 16'd2301, 16'd19204, 16'd14176, 16'd47228, 16'd65528, 16'd9588, 16'd60663, 16'd4152, 16'd21328, 16'd12611, 16'd50181, 16'd61504, 16'd11244, 16'd5753, 16'd59147, 16'd53441, 16'd43946});
	test_expansion(128'h7e0bb6659e5426dafcbc76b49fd98689, {16'd57963, 16'd58290, 16'd40905, 16'd10633, 16'd61153, 16'd15364, 16'd7684, 16'd41702, 16'd53959, 16'd2021, 16'd52816, 16'd62838, 16'd56135, 16'd20958, 16'd55141, 16'd48206, 16'd50563, 16'd64253, 16'd65208, 16'd5611, 16'd39645, 16'd26700, 16'd1459, 16'd41470, 16'd25468, 16'd563});
	test_expansion(128'hf4bf6d42fc968dceeb8269081ffd4e22, {16'd16013, 16'd56242, 16'd7184, 16'd1927, 16'd18397, 16'd29720, 16'd26680, 16'd13541, 16'd59630, 16'd10068, 16'd13337, 16'd37623, 16'd26421, 16'd22105, 16'd24614, 16'd56690, 16'd15030, 16'd31986, 16'd14002, 16'd46474, 16'd20025, 16'd28586, 16'd53179, 16'd21777, 16'd32369, 16'd31922});
	test_expansion(128'ha77e76a6f7c62e9bad4187a5ebe4f784, {16'd14042, 16'd13681, 16'd51323, 16'd51046, 16'd11279, 16'd16109, 16'd54250, 16'd25072, 16'd24973, 16'd7139, 16'd22764, 16'd32337, 16'd44490, 16'd2839, 16'd50647, 16'd59823, 16'd34429, 16'd26868, 16'd59208, 16'd54709, 16'd17198, 16'd58898, 16'd26009, 16'd44622, 16'd39145, 16'd49439});
	test_expansion(128'h395a670fe7e0faf68487c9e1f0bd0979, {16'd61777, 16'd3658, 16'd47423, 16'd61935, 16'd420, 16'd3920, 16'd63688, 16'd12508, 16'd36646, 16'd26073, 16'd27238, 16'd36684, 16'd64527, 16'd52694, 16'd9511, 16'd55753, 16'd13373, 16'd39160, 16'd57354, 16'd22067, 16'd6475, 16'd49718, 16'd50004, 16'd57238, 16'd48118, 16'd10311});
	test_expansion(128'h9618a0348f59d648c384726a3a5929f2, {16'd24444, 16'd42235, 16'd40307, 16'd7015, 16'd9218, 16'd65354, 16'd44826, 16'd4205, 16'd2933, 16'd31498, 16'd11269, 16'd2611, 16'd39084, 16'd21264, 16'd21145, 16'd43954, 16'd44717, 16'd28025, 16'd35465, 16'd39295, 16'd33206, 16'd63508, 16'd16689, 16'd62885, 16'd39329, 16'd22149});
	test_expansion(128'ha94cd7e99a78d3396880cde8913e627a, {16'd23551, 16'd11638, 16'd10395, 16'd20003, 16'd26027, 16'd41566, 16'd64240, 16'd50950, 16'd5444, 16'd58419, 16'd9611, 16'd19357, 16'd2070, 16'd38843, 16'd13720, 16'd21208, 16'd12085, 16'd64045, 16'd48123, 16'd49135, 16'd9325, 16'd19264, 16'd47760, 16'd44838, 16'd64972, 16'd39939});
	test_expansion(128'h48bcf3d89b4d439197512e8ce36767bb, {16'd43346, 16'd64409, 16'd18504, 16'd16192, 16'd25345, 16'd28292, 16'd39183, 16'd9494, 16'd42509, 16'd62304, 16'd41933, 16'd16137, 16'd38054, 16'd59719, 16'd26345, 16'd2730, 16'd25942, 16'd65031, 16'd39171, 16'd19565, 16'd26075, 16'd22378, 16'd57970, 16'd22636, 16'd46416, 16'd9646});
	test_expansion(128'h0683ebba65ad687dbdd7b12af1c834d5, {16'd24271, 16'd28629, 16'd26209, 16'd53218, 16'd65087, 16'd32463, 16'd65206, 16'd8596, 16'd22046, 16'd4644, 16'd64810, 16'd36073, 16'd53901, 16'd22670, 16'd4776, 16'd26792, 16'd12263, 16'd45160, 16'd23240, 16'd21778, 16'd56995, 16'd42757, 16'd40940, 16'd65140, 16'd16640, 16'd32348});
	test_expansion(128'hd6dedab9772909fc89264628dfcbf1f2, {16'd52323, 16'd11691, 16'd12082, 16'd15460, 16'd40959, 16'd30605, 16'd45236, 16'd26284, 16'd60139, 16'd35491, 16'd53997, 16'd28561, 16'd50151, 16'd29823, 16'd4922, 16'd50428, 16'd32825, 16'd64549, 16'd44613, 16'd40833, 16'd41585, 16'd29015, 16'd15544, 16'd49757, 16'd19920, 16'd31782});
	test_expansion(128'he8286aa14f00b9237f7e9089473537ef, {16'd123, 16'd7465, 16'd64497, 16'd60650, 16'd8453, 16'd51094, 16'd26221, 16'd18463, 16'd55273, 16'd3634, 16'd8347, 16'd12685, 16'd32364, 16'd7883, 16'd50893, 16'd59941, 16'd56413, 16'd53613, 16'd31159, 16'd19165, 16'd10991, 16'd53716, 16'd35940, 16'd16439, 16'd26747, 16'd8443});
	test_expansion(128'h896e0168b93792e51080824690b1df42, {16'd3048, 16'd39161, 16'd41513, 16'd6022, 16'd61218, 16'd7253, 16'd33487, 16'd2100, 16'd22979, 16'd24811, 16'd50485, 16'd45802, 16'd59875, 16'd23572, 16'd29370, 16'd45397, 16'd63964, 16'd55773, 16'd29495, 16'd57661, 16'd12087, 16'd58421, 16'd62679, 16'd63031, 16'd50142, 16'd25971});
	test_expansion(128'ha1775024b495a02ca2f21a5afa65fc46, {16'd37086, 16'd47713, 16'd24711, 16'd8243, 16'd30819, 16'd25732, 16'd19410, 16'd9172, 16'd41659, 16'd46099, 16'd10835, 16'd53815, 16'd26678, 16'd1667, 16'd22576, 16'd54880, 16'd7885, 16'd28815, 16'd42113, 16'd44916, 16'd7167, 16'd50420, 16'd19029, 16'd34080, 16'd25445, 16'd10416});
	test_expansion(128'h873329ba99d84ffd22a215a8727a8633, {16'd11024, 16'd51680, 16'd25836, 16'd56694, 16'd40471, 16'd35656, 16'd35147, 16'd2591, 16'd10338, 16'd59791, 16'd47075, 16'd24621, 16'd32955, 16'd34707, 16'd53886, 16'd25832, 16'd18975, 16'd983, 16'd9237, 16'd45140, 16'd52608, 16'd27302, 16'd58633, 16'd41415, 16'd1469, 16'd7373});
	test_expansion(128'h4b694656c0e9c7478ae5dd28e5b19c25, {16'd23606, 16'd17232, 16'd8108, 16'd3071, 16'd23668, 16'd7338, 16'd18060, 16'd16107, 16'd14227, 16'd46432, 16'd12240, 16'd6086, 16'd33385, 16'd25335, 16'd62422, 16'd52016, 16'd32588, 16'd22567, 16'd32257, 16'd44474, 16'd42532, 16'd65426, 16'd64915, 16'd34985, 16'd44306, 16'd8662});
	test_expansion(128'hdbd6de2ac04d2c8748a317ba20140d0a, {16'd43509, 16'd65026, 16'd54203, 16'd15267, 16'd26625, 16'd31976, 16'd27975, 16'd26625, 16'd1308, 16'd58250, 16'd60464, 16'd882, 16'd36911, 16'd53605, 16'd63675, 16'd52093, 16'd23348, 16'd36867, 16'd24844, 16'd7459, 16'd6946, 16'd53839, 16'd38780, 16'd65292, 16'd29979, 16'd58988});
	test_expansion(128'h3cc0ff4af2ca33826c218646332f4786, {16'd41567, 16'd59671, 16'd1372, 16'd62308, 16'd7561, 16'd60932, 16'd30078, 16'd27258, 16'd37313, 16'd3376, 16'd50457, 16'd58143, 16'd34453, 16'd9906, 16'd43975, 16'd64730, 16'd36100, 16'd42628, 16'd50207, 16'd10771, 16'd29850, 16'd64058, 16'd2277, 16'd1393, 16'd53935, 16'd58900});
	test_expansion(128'ha5f765e464370b5d638848cb0d865834, {16'd40951, 16'd58064, 16'd52139, 16'd19273, 16'd44757, 16'd58111, 16'd11641, 16'd51081, 16'd39563, 16'd13788, 16'd27176, 16'd8880, 16'd1094, 16'd30009, 16'd43444, 16'd20663, 16'd10816, 16'd35940, 16'd9212, 16'd9231, 16'd8130, 16'd9551, 16'd31893, 16'd28026, 16'd58207, 16'd36651});
	test_expansion(128'hf9ce7aadd6b532229b8913e5a87c407d, {16'd14348, 16'd45522, 16'd19175, 16'd30818, 16'd45064, 16'd10094, 16'd46107, 16'd39048, 16'd517, 16'd25927, 16'd13336, 16'd8125, 16'd20947, 16'd43815, 16'd8004, 16'd48163, 16'd21651, 16'd2883, 16'd1661, 16'd32317, 16'd19381, 16'd61511, 16'd914, 16'd38963, 16'd35146, 16'd23062});
	test_expansion(128'h44450f9365a4ce5c44c6ed634942fe4f, {16'd51387, 16'd61142, 16'd32933, 16'd38304, 16'd33807, 16'd34759, 16'd29034, 16'd15033, 16'd56629, 16'd33510, 16'd13857, 16'd50066, 16'd43797, 16'd46635, 16'd52292, 16'd22285, 16'd46440, 16'd29665, 16'd11534, 16'd39111, 16'd39068, 16'd58154, 16'd64860, 16'd64648, 16'd52403, 16'd24514});
	test_expansion(128'h5603ffd06358628ae2097dc86a5752be, {16'd56063, 16'd59864, 16'd57863, 16'd17260, 16'd31347, 16'd27626, 16'd39161, 16'd39880, 16'd5327, 16'd37459, 16'd42529, 16'd56196, 16'd355, 16'd33777, 16'd36394, 16'd25180, 16'd25816, 16'd33010, 16'd28115, 16'd20732, 16'd42000, 16'd16788, 16'd18985, 16'd28862, 16'd56252, 16'd49123});
	test_expansion(128'h455cd2100b720e9094c1149249ce92ee, {16'd45577, 16'd59796, 16'd13497, 16'd29064, 16'd4624, 16'd33648, 16'd12625, 16'd37404, 16'd10598, 16'd57264, 16'd45726, 16'd51511, 16'd65026, 16'd35131, 16'd35302, 16'd37474, 16'd30955, 16'd60477, 16'd11584, 16'd47895, 16'd19052, 16'd36442, 16'd6948, 16'd6289, 16'd22501, 16'd58200});
	test_expansion(128'h00fbcc7cdecf21274ddb5e3b92a03ff1, {16'd64032, 16'd28050, 16'd50141, 16'd17616, 16'd37543, 16'd44225, 16'd6870, 16'd47393, 16'd55178, 16'd27012, 16'd40820, 16'd42303, 16'd35446, 16'd61973, 16'd17486, 16'd52271, 16'd37037, 16'd56740, 16'd1045, 16'd49757, 16'd57052, 16'd40577, 16'd60848, 16'd6612, 16'd62348, 16'd44004});
	test_expansion(128'hd6088584fc72c2155f7dfa7fa6e5c9af, {16'd34871, 16'd26614, 16'd9920, 16'd409, 16'd47592, 16'd11040, 16'd23085, 16'd56095, 16'd64387, 16'd16147, 16'd33033, 16'd11376, 16'd14818, 16'd22905, 16'd34743, 16'd13936, 16'd12447, 16'd18000, 16'd53598, 16'd47608, 16'd6945, 16'd57344, 16'd59898, 16'd37082, 16'd20720, 16'd61143});
	test_expansion(128'hf49763a20e31a4b9e8c4548154ff59f1, {16'd25458, 16'd16514, 16'd53588, 16'd14620, 16'd25976, 16'd19033, 16'd38100, 16'd8456, 16'd39939, 16'd57186, 16'd57006, 16'd50889, 16'd23815, 16'd36712, 16'd28113, 16'd3527, 16'd37298, 16'd40241, 16'd59520, 16'd36317, 16'd29482, 16'd62262, 16'd56279, 16'd45102, 16'd17759, 16'd25629});
	test_expansion(128'h1176c416811fc023ef345e6cf69e6803, {16'd16845, 16'd46406, 16'd6060, 16'd60199, 16'd48921, 16'd34672, 16'd47114, 16'd560, 16'd57234, 16'd59750, 16'd19914, 16'd6956, 16'd14580, 16'd11148, 16'd36705, 16'd3117, 16'd10599, 16'd39847, 16'd27352, 16'd6499, 16'd2923, 16'd20784, 16'd44878, 16'd44619, 16'd23247, 16'd41915});
	test_expansion(128'hd5c2c658d7770d681d15a499cbab36d0, {16'd49247, 16'd14402, 16'd31075, 16'd55073, 16'd54908, 16'd5261, 16'd54526, 16'd62466, 16'd27813, 16'd40196, 16'd53142, 16'd10190, 16'd56891, 16'd43723, 16'd41051, 16'd40001, 16'd2266, 16'd24322, 16'd3803, 16'd491, 16'd48974, 16'd47819, 16'd51991, 16'd38294, 16'd45462, 16'd31919});
	test_expansion(128'hd5139a946af2fd1ba8bf0cca10831f6b, {16'd19672, 16'd18627, 16'd57181, 16'd20283, 16'd1138, 16'd12614, 16'd17483, 16'd8238, 16'd1415, 16'd21469, 16'd24250, 16'd35420, 16'd18566, 16'd23273, 16'd17845, 16'd16721, 16'd29126, 16'd33047, 16'd23924, 16'd1803, 16'd65251, 16'd52307, 16'd18086, 16'd24421, 16'd19881, 16'd5941});
	test_expansion(128'h101aa8265fe072a42bd9ff45c1d20d55, {16'd1007, 16'd55448, 16'd47850, 16'd15794, 16'd46474, 16'd30271, 16'd61683, 16'd4248, 16'd21542, 16'd24951, 16'd57201, 16'd9450, 16'd29187, 16'd39083, 16'd30741, 16'd34300, 16'd56624, 16'd4423, 16'd48115, 16'd53284, 16'd43880, 16'd63796, 16'd61225, 16'd42133, 16'd33990, 16'd16962});
	test_expansion(128'hef348cc0f3551393c2c4878b38439fc8, {16'd10521, 16'd7550, 16'd8953, 16'd11475, 16'd8323, 16'd64044, 16'd48883, 16'd11613, 16'd53566, 16'd14004, 16'd61669, 16'd56483, 16'd32208, 16'd65150, 16'd17487, 16'd51779, 16'd59293, 16'd58109, 16'd10706, 16'd50082, 16'd16634, 16'd30756, 16'd10767, 16'd12589, 16'd2442, 16'd52858});
	test_expansion(128'h40f84bc4a99835d1285eea686ac3c104, {16'd10993, 16'd40353, 16'd27687, 16'd22549, 16'd61631, 16'd60482, 16'd21438, 16'd17662, 16'd21259, 16'd10264, 16'd57877, 16'd26215, 16'd58200, 16'd13033, 16'd1908, 16'd1949, 16'd4036, 16'd57829, 16'd49738, 16'd36578, 16'd42847, 16'd47520, 16'd52579, 16'd1577, 16'd53030, 16'd61641});
	test_expansion(128'hf3dc499c606ee530897099e4b733a15e, {16'd58032, 16'd19226, 16'd19593, 16'd62072, 16'd24693, 16'd18296, 16'd54603, 16'd11446, 16'd37590, 16'd46935, 16'd14666, 16'd3485, 16'd474, 16'd59828, 16'd62751, 16'd63729, 16'd41776, 16'd62029, 16'd40395, 16'd8024, 16'd52032, 16'd15273, 16'd46746, 16'd48212, 16'd31908, 16'd51046});
	test_expansion(128'hf959a6f9412cc683580154cfe114262a, {16'd61234, 16'd1072, 16'd65502, 16'd18255, 16'd41195, 16'd950, 16'd15774, 16'd37635, 16'd24340, 16'd59033, 16'd1435, 16'd23420, 16'd16087, 16'd40586, 16'd46213, 16'd57314, 16'd48285, 16'd18198, 16'd32239, 16'd41172, 16'd15374, 16'd40950, 16'd58103, 16'd17231, 16'd16449, 16'd54929});
	test_expansion(128'hb3989c91f52e828874d28ea2272ac23b, {16'd32347, 16'd2674, 16'd33273, 16'd57140, 16'd19338, 16'd64186, 16'd64663, 16'd59080, 16'd45899, 16'd47900, 16'd46965, 16'd63260, 16'd8717, 16'd64790, 16'd25384, 16'd31889, 16'd56281, 16'd10237, 16'd24714, 16'd36912, 16'd62550, 16'd13333, 16'd2264, 16'd36021, 16'd12958, 16'd35875});
	test_expansion(128'h046108a7d139606f9d84cbd563a7df9d, {16'd61044, 16'd54697, 16'd42089, 16'd31607, 16'd14711, 16'd56250, 16'd30246, 16'd40907, 16'd34231, 16'd20386, 16'd29850, 16'd33661, 16'd52121, 16'd65174, 16'd28211, 16'd27538, 16'd45869, 16'd45479, 16'd48238, 16'd59250, 16'd53204, 16'd21360, 16'd57297, 16'd65237, 16'd297, 16'd61828});
	test_expansion(128'h5a965596b70b8d5f5724cc737111801a, {16'd7134, 16'd50865, 16'd16595, 16'd6065, 16'd45504, 16'd49522, 16'd29335, 16'd45298, 16'd55035, 16'd17705, 16'd42193, 16'd1769, 16'd39004, 16'd10781, 16'd59067, 16'd33215, 16'd8320, 16'd22158, 16'd43289, 16'd65263, 16'd30781, 16'd53324, 16'd24005, 16'd235, 16'd40579, 16'd42438});
	test_expansion(128'hbdba9e2b4200f0be2b5eeed42130e7ac, {16'd2524, 16'd53842, 16'd24267, 16'd58086, 16'd58504, 16'd34802, 16'd54740, 16'd46411, 16'd24643, 16'd57984, 16'd31579, 16'd22882, 16'd52901, 16'd10128, 16'd47008, 16'd5011, 16'd37283, 16'd35557, 16'd10085, 16'd48016, 16'd39959, 16'd27968, 16'd27944, 16'd32262, 16'd51176, 16'd14076});
	test_expansion(128'h499cc5c79f30c7ce2a5b9b89510a845a, {16'd6523, 16'd16509, 16'd52837, 16'd44275, 16'd27760, 16'd44286, 16'd3126, 16'd47735, 16'd8386, 16'd45846, 16'd56130, 16'd21503, 16'd45740, 16'd46702, 16'd46940, 16'd61857, 16'd32375, 16'd43071, 16'd35306, 16'd12822, 16'd23498, 16'd47735, 16'd63402, 16'd1835, 16'd28848, 16'd16079});
	test_expansion(128'h1a9dee823a2e58113c15c741f3f4e530, {16'd23349, 16'd286, 16'd50247, 16'd40467, 16'd60438, 16'd903, 16'd53650, 16'd57386, 16'd12916, 16'd43586, 16'd45258, 16'd31383, 16'd43763, 16'd60203, 16'd38856, 16'd52713, 16'd44981, 16'd33122, 16'd40242, 16'd30663, 16'd31525, 16'd9730, 16'd61376, 16'd25928, 16'd4644, 16'd14695});
	test_expansion(128'hf4321464a72ac6af9cf69a090409c824, {16'd45610, 16'd23348, 16'd37532, 16'd9015, 16'd51318, 16'd22332, 16'd31133, 16'd44383, 16'd40501, 16'd1547, 16'd57321, 16'd20775, 16'd43728, 16'd11935, 16'd53996, 16'd55277, 16'd34272, 16'd61774, 16'd50441, 16'd52839, 16'd21103, 16'd54161, 16'd34155, 16'd10010, 16'd13684, 16'd54873});
	test_expansion(128'h5558571283ee19d2ef65846a0bd4a127, {16'd51813, 16'd33786, 16'd23643, 16'd17113, 16'd28704, 16'd45103, 16'd59582, 16'd39425, 16'd51209, 16'd25613, 16'd19974, 16'd33471, 16'd45654, 16'd51754, 16'd50174, 16'd7883, 16'd52567, 16'd34906, 16'd7512, 16'd2230, 16'd59267, 16'd8258, 16'd46111, 16'd18735, 16'd29158, 16'd51701});
	test_expansion(128'hbfd9a56b424e6a2f3574fb36d89ba3a3, {16'd41328, 16'd12200, 16'd15835, 16'd992, 16'd45218, 16'd4856, 16'd16386, 16'd49263, 16'd35565, 16'd7031, 16'd48029, 16'd50468, 16'd12036, 16'd29118, 16'd33631, 16'd38455, 16'd39325, 16'd38231, 16'd12489, 16'd46413, 16'd20371, 16'd5091, 16'd52029, 16'd17989, 16'd61260, 16'd8861});
	test_expansion(128'h9d84790e0f52087080a2336c356769f7, {16'd57475, 16'd21624, 16'd41251, 16'd24516, 16'd23318, 16'd44903, 16'd45922, 16'd43976, 16'd22376, 16'd29678, 16'd21976, 16'd57913, 16'd7035, 16'd62288, 16'd7160, 16'd3905, 16'd6343, 16'd38323, 16'd27085, 16'd40246, 16'd59296, 16'd55273, 16'd51138, 16'd44074, 16'd37828, 16'd41953});
	test_expansion(128'h2825033e7bda607783fd22bc50a5e81c, {16'd35955, 16'd10420, 16'd56677, 16'd52653, 16'd42948, 16'd5171, 16'd27861, 16'd44157, 16'd25835, 16'd260, 16'd22730, 16'd28830, 16'd34302, 16'd17854, 16'd46257, 16'd30005, 16'd15551, 16'd23641, 16'd5902, 16'd5320, 16'd36910, 16'd11885, 16'd38949, 16'd27287, 16'd64572, 16'd53139});
	test_expansion(128'ha342ed67b3ab829c3ee7b98df4be0b77, {16'd26567, 16'd42875, 16'd39153, 16'd12354, 16'd34114, 16'd48809, 16'd9480, 16'd19117, 16'd44046, 16'd40029, 16'd18272, 16'd19460, 16'd27100, 16'd32517, 16'd1656, 16'd2084, 16'd1532, 16'd43252, 16'd25077, 16'd26060, 16'd49095, 16'd40105, 16'd14150, 16'd13528, 16'd52806, 16'd9511});
	test_expansion(128'h45dfc949c9c1327afc720540ef410906, {16'd49339, 16'd20218, 16'd55768, 16'd43007, 16'd40189, 16'd31858, 16'd53035, 16'd26494, 16'd61625, 16'd5448, 16'd20822, 16'd9118, 16'd3826, 16'd10084, 16'd49778, 16'd24509, 16'd54849, 16'd61546, 16'd46445, 16'd1884, 16'd33261, 16'd27154, 16'd33186, 16'd60090, 16'd18968, 16'd56914});
	test_expansion(128'h369658582ffd0b3a3f100b34e3a9818e, {16'd50695, 16'd25055, 16'd57364, 16'd19086, 16'd58625, 16'd9865, 16'd34039, 16'd30162, 16'd61152, 16'd64582, 16'd60464, 16'd41946, 16'd36461, 16'd34926, 16'd28626, 16'd48376, 16'd10857, 16'd63454, 16'd37608, 16'd7444, 16'd59632, 16'd60856, 16'd62868, 16'd18215, 16'd46566, 16'd36911});
	test_expansion(128'h1490e203eea4f27f2c76e359c11ff3f9, {16'd58482, 16'd51587, 16'd30315, 16'd44454, 16'd32377, 16'd8470, 16'd9629, 16'd14122, 16'd11748, 16'd62070, 16'd12324, 16'd60598, 16'd11531, 16'd9233, 16'd2176, 16'd8551, 16'd7876, 16'd44552, 16'd29859, 16'd29269, 16'd61048, 16'd15805, 16'd3338, 16'd53632, 16'd5168, 16'd33422});
	test_expansion(128'h71c8b6d8441c1958ef73d86e9ec44f5b, {16'd57341, 16'd63496, 16'd47754, 16'd8617, 16'd45245, 16'd56591, 16'd35939, 16'd35829, 16'd46266, 16'd60808, 16'd45648, 16'd15515, 16'd55212, 16'd60559, 16'd13161, 16'd8765, 16'd45350, 16'd22456, 16'd7118, 16'd665, 16'd4292, 16'd15197, 16'd36093, 16'd58730, 16'd58772, 16'd6606});
	test_expansion(128'h8657805969ff62922cca59aa95e05e95, {16'd36445, 16'd1231, 16'd48563, 16'd54497, 16'd7384, 16'd35022, 16'd57995, 16'd12552, 16'd49207, 16'd5136, 16'd46546, 16'd31070, 16'd59295, 16'd59251, 16'd59326, 16'd34767, 16'd19384, 16'd47284, 16'd62169, 16'd46203, 16'd35308, 16'd1500, 16'd56331, 16'd32664, 16'd42816, 16'd15744});
	test_expansion(128'h7e14de409e80db168f01dbfc608968f8, {16'd26022, 16'd44536, 16'd39709, 16'd23752, 16'd5096, 16'd12257, 16'd61844, 16'd20491, 16'd37654, 16'd58469, 16'd59585, 16'd18884, 16'd25544, 16'd23922, 16'd52287, 16'd62483, 16'd451, 16'd5692, 16'd36572, 16'd2496, 16'd5300, 16'd29351, 16'd35521, 16'd50914, 16'd33160, 16'd723});
	test_expansion(128'ha7486b0eda385da701f4bcb41a618be3, {16'd16163, 16'd4153, 16'd35850, 16'd22006, 16'd34105, 16'd20281, 16'd3375, 16'd31717, 16'd33768, 16'd28628, 16'd63606, 16'd27325, 16'd6085, 16'd5326, 16'd23066, 16'd34794, 16'd3685, 16'd41681, 16'd36806, 16'd18850, 16'd3449, 16'd52830, 16'd57675, 16'd35484, 16'd19574, 16'd14134});
	test_expansion(128'hed09608e7c8093dd9ee91fd474fc770f, {16'd61951, 16'd27840, 16'd56354, 16'd35573, 16'd57197, 16'd13166, 16'd48458, 16'd58188, 16'd58024, 16'd53331, 16'd55725, 16'd21077, 16'd3765, 16'd10085, 16'd30921, 16'd22993, 16'd29613, 16'd21671, 16'd40542, 16'd19333, 16'd41360, 16'd65041, 16'd32031, 16'd21759, 16'd29822, 16'd31455});
	test_expansion(128'hc2a51990d507bb98752788f8e01c9454, {16'd9982, 16'd56740, 16'd60142, 16'd47176, 16'd9300, 16'd55850, 16'd6116, 16'd52102, 16'd56864, 16'd26859, 16'd5692, 16'd35376, 16'd18618, 16'd40440, 16'd52415, 16'd7334, 16'd18261, 16'd57683, 16'd50535, 16'd46993, 16'd50753, 16'd39320, 16'd38909, 16'd52670, 16'd47732, 16'd48020});
	test_expansion(128'hee2412550f65fcb7b5f76cc48d5fbcba, {16'd46007, 16'd51904, 16'd34371, 16'd13885, 16'd4109, 16'd56331, 16'd42183, 16'd26339, 16'd19890, 16'd19907, 16'd17266, 16'd14114, 16'd51293, 16'd21776, 16'd41017, 16'd62440, 16'd52882, 16'd24691, 16'd20890, 16'd30770, 16'd62239, 16'd31557, 16'd10584, 16'd51265, 16'd17006, 16'd24358});
	test_expansion(128'h8ae7e47e051c275b3a2e35dc5def0ad9, {16'd2578, 16'd1699, 16'd31025, 16'd14332, 16'd42001, 16'd6544, 16'd10127, 16'd58407, 16'd39512, 16'd20128, 16'd18117, 16'd36712, 16'd26834, 16'd26902, 16'd11845, 16'd41390, 16'd36647, 16'd56885, 16'd29859, 16'd34984, 16'd9747, 16'd21896, 16'd49698, 16'd40694, 16'd28156, 16'd16524});
	test_expansion(128'h9313417a157863ca23d576355a7c316b, {16'd59754, 16'd37613, 16'd9234, 16'd28791, 16'd14149, 16'd39423, 16'd31140, 16'd28708, 16'd29857, 16'd53453, 16'd54239, 16'd14553, 16'd16600, 16'd11069, 16'd11435, 16'd13190, 16'd13481, 16'd34689, 16'd22659, 16'd39659, 16'd50230, 16'd27734, 16'd32861, 16'd38801, 16'd39297, 16'd4101});
	test_expansion(128'h6ffc17a6ab345b8648c458d28cd9cf2f, {16'd26796, 16'd4414, 16'd28292, 16'd11996, 16'd8751, 16'd43257, 16'd31748, 16'd13500, 16'd26894, 16'd35274, 16'd13354, 16'd47741, 16'd35849, 16'd42383, 16'd29317, 16'd36539, 16'd39870, 16'd44028, 16'd60703, 16'd27795, 16'd62364, 16'd60941, 16'd21604, 16'd62454, 16'd53709, 16'd223});
	test_expansion(128'hfc00c2ebb8686a7f11f7e5a9fa19fa88, {16'd30873, 16'd50579, 16'd9471, 16'd2024, 16'd55914, 16'd64976, 16'd62630, 16'd33495, 16'd6100, 16'd48978, 16'd9943, 16'd7241, 16'd3496, 16'd44499, 16'd39477, 16'd35726, 16'd49732, 16'd61334, 16'd35188, 16'd1411, 16'd63434, 16'd5101, 16'd1615, 16'd16769, 16'd31822, 16'd41514});
	test_expansion(128'hb990b8b3bdcade869386c45ef9693beb, {16'd26313, 16'd22309, 16'd16675, 16'd56748, 16'd47673, 16'd540, 16'd35397, 16'd30740, 16'd19064, 16'd23081, 16'd12461, 16'd30210, 16'd33046, 16'd51684, 16'd45771, 16'd23619, 16'd38709, 16'd63722, 16'd855, 16'd28419, 16'd7869, 16'd55462, 16'd64961, 16'd22381, 16'd17025, 16'd52891});
	test_expansion(128'hc48757e9a7ef0af5353757c071bfc06a, {16'd13426, 16'd57736, 16'd2461, 16'd60336, 16'd38975, 16'd41276, 16'd29792, 16'd8320, 16'd7266, 16'd41744, 16'd41675, 16'd43887, 16'd3618, 16'd63541, 16'd47600, 16'd12712, 16'd1707, 16'd46067, 16'd64395, 16'd57197, 16'd62558, 16'd64576, 16'd38135, 16'd37200, 16'd40136, 16'd54128});
	test_expansion(128'h72a659cce23b8c905bdfbb8b66d5255d, {16'd9041, 16'd29837, 16'd51965, 16'd57827, 16'd15685, 16'd61716, 16'd41835, 16'd26750, 16'd53063, 16'd18399, 16'd3043, 16'd45260, 16'd12518, 16'd35781, 16'd41925, 16'd47895, 16'd45309, 16'd20462, 16'd60970, 16'd21042, 16'd42051, 16'd33242, 16'd21996, 16'd11576, 16'd8893, 16'd6735});
	test_expansion(128'h58eba18b23768e55b8f32fc327260c29, {16'd8703, 16'd53124, 16'd51256, 16'd4707, 16'd42717, 16'd61788, 16'd34485, 16'd56879, 16'd1748, 16'd21799, 16'd36380, 16'd58810, 16'd52122, 16'd52072, 16'd59518, 16'd61634, 16'd45572, 16'd62339, 16'd33319, 16'd61779, 16'd65164, 16'd2372, 16'd47339, 16'd4802, 16'd8602, 16'd35752});
	test_expansion(128'h2a636da4005de456820fb0e4e704297a, {16'd26426, 16'd4479, 16'd55909, 16'd24350, 16'd987, 16'd50163, 16'd33874, 16'd49563, 16'd61100, 16'd60412, 16'd34012, 16'd32302, 16'd113, 16'd31630, 16'd30245, 16'd62470, 16'd9501, 16'd48135, 16'd2079, 16'd19752, 16'd36730, 16'd63606, 16'd15017, 16'd43213, 16'd5246, 16'd57510});
	test_expansion(128'hd0e13d3fdb4a8de429a612633608766c, {16'd5420, 16'd7302, 16'd56711, 16'd60850, 16'd47596, 16'd13671, 16'd23444, 16'd64502, 16'd4725, 16'd27910, 16'd61395, 16'd17661, 16'd40846, 16'd12013, 16'd45717, 16'd7547, 16'd7101, 16'd64591, 16'd27896, 16'd3437, 16'd46877, 16'd36443, 16'd22345, 16'd60563, 16'd52051, 16'd48750});
	test_expansion(128'hd332b686cc20130aadb2b7a57f318bb1, {16'd24977, 16'd7099, 16'd61475, 16'd30999, 16'd57347, 16'd24928, 16'd10567, 16'd60602, 16'd7697, 16'd8140, 16'd1262, 16'd14097, 16'd605, 16'd64686, 16'd58910, 16'd56728, 16'd40384, 16'd24805, 16'd38765, 16'd43723, 16'd19793, 16'd10134, 16'd10610, 16'd23706, 16'd28453, 16'd19157});
	test_expansion(128'hf4b5a73a56a22772a1b8115372f13c8f, {16'd62551, 16'd31691, 16'd6836, 16'd10100, 16'd63682, 16'd5862, 16'd40462, 16'd62544, 16'd39571, 16'd48150, 16'd50159, 16'd11937, 16'd10044, 16'd56806, 16'd58761, 16'd44260, 16'd34267, 16'd20927, 16'd29381, 16'd53784, 16'd12832, 16'd33074, 16'd19283, 16'd35698, 16'd42643, 16'd32893});
	test_expansion(128'h9cc89e3b5be8413cb0b514d1062186c7, {16'd19569, 16'd64227, 16'd24114, 16'd12156, 16'd54743, 16'd24660, 16'd22560, 16'd63852, 16'd14294, 16'd52090, 16'd38214, 16'd30777, 16'd10135, 16'd30009, 16'd53367, 16'd41463, 16'd37400, 16'd48520, 16'd40171, 16'd58917, 16'd51489, 16'd27245, 16'd14754, 16'd62376, 16'd57485, 16'd9806});
	test_expansion(128'h2191b91b881f53e54ef7a172af287552, {16'd6070, 16'd42737, 16'd29202, 16'd49494, 16'd667, 16'd47550, 16'd42263, 16'd54271, 16'd10965, 16'd28073, 16'd14807, 16'd42176, 16'd10819, 16'd6165, 16'd12808, 16'd56506, 16'd35834, 16'd47092, 16'd59800, 16'd49428, 16'd43684, 16'd19551, 16'd2604, 16'd21316, 16'd7919, 16'd9852});
	test_expansion(128'h9ec345b67dcf87814cb5f53023f0cfaf, {16'd28262, 16'd39815, 16'd11588, 16'd33391, 16'd49534, 16'd63124, 16'd34191, 16'd54185, 16'd42475, 16'd46877, 16'd9316, 16'd3958, 16'd1761, 16'd31547, 16'd20853, 16'd7891, 16'd39281, 16'd25262, 16'd33638, 16'd1619, 16'd25327, 16'd30557, 16'd34979, 16'd16325, 16'd32748, 16'd18943});
	test_expansion(128'hb188b898a52cddfd31c2ec79757b02fc, {16'd47862, 16'd59943, 16'd55029, 16'd5967, 16'd46019, 16'd59739, 16'd40726, 16'd4472, 16'd7627, 16'd47720, 16'd60324, 16'd4935, 16'd52025, 16'd46519, 16'd34266, 16'd55062, 16'd48021, 16'd12438, 16'd50251, 16'd23195, 16'd3549, 16'd11656, 16'd13679, 16'd51721, 16'd45119, 16'd40045});
	test_expansion(128'h96713e7dfb48a68505555d17555b58af, {16'd40202, 16'd37782, 16'd51122, 16'd62157, 16'd42338, 16'd4598, 16'd59666, 16'd14590, 16'd376, 16'd341, 16'd54346, 16'd25282, 16'd42949, 16'd46585, 16'd2357, 16'd24874, 16'd30550, 16'd65255, 16'd26476, 16'd38942, 16'd50202, 16'd60516, 16'd20209, 16'd54771, 16'd40621, 16'd23380});
	test_expansion(128'h5395d0110e616e71a74912fbef834fd4, {16'd6851, 16'd32683, 16'd38683, 16'd16736, 16'd49099, 16'd44271, 16'd6556, 16'd361, 16'd53075, 16'd55193, 16'd16984, 16'd25829, 16'd49878, 16'd7420, 16'd47103, 16'd2614, 16'd61632, 16'd58491, 16'd23878, 16'd42509, 16'd60600, 16'd2690, 16'd49195, 16'd25738, 16'd45218, 16'd17891});
	test_expansion(128'h5c19b3da7d133af6a1b21e4e17b051a9, {16'd27928, 16'd31449, 16'd293, 16'd46032, 16'd820, 16'd53967, 16'd34116, 16'd29070, 16'd4626, 16'd21185, 16'd15386, 16'd1233, 16'd15340, 16'd21824, 16'd28217, 16'd24031, 16'd54917, 16'd22266, 16'd9279, 16'd61571, 16'd21688, 16'd17941, 16'd12019, 16'd34317, 16'd21084, 16'd56045});
	test_expansion(128'h7ee4fd1a5eb928881984b05f9ceed33b, {16'd14651, 16'd1364, 16'd3544, 16'd19042, 16'd11877, 16'd1194, 16'd49283, 16'd12691, 16'd18159, 16'd10303, 16'd11219, 16'd26977, 16'd19363, 16'd35600, 16'd60307, 16'd26694, 16'd24569, 16'd11705, 16'd35593, 16'd38112, 16'd2088, 16'd6216, 16'd31324, 16'd18141, 16'd45700, 16'd42038});
	test_expansion(128'hfbe615fe58f5c1a1865fddd3eb779ac4, {16'd25502, 16'd42309, 16'd63519, 16'd63682, 16'd29431, 16'd9938, 16'd40672, 16'd36966, 16'd27054, 16'd60671, 16'd18139, 16'd49418, 16'd17, 16'd63783, 16'd63085, 16'd9286, 16'd5039, 16'd10824, 16'd58660, 16'd19917, 16'd41512, 16'd38646, 16'd14604, 16'd42580, 16'd60708, 16'd45749});
	test_expansion(128'h81e17ed56e3a14c126ba11c52110aa96, {16'd50540, 16'd49648, 16'd60348, 16'd10020, 16'd35395, 16'd20927, 16'd38217, 16'd53741, 16'd14129, 16'd29259, 16'd872, 16'd52239, 16'd29199, 16'd41069, 16'd50323, 16'd29750, 16'd29104, 16'd27890, 16'd38653, 16'd5928, 16'd13887, 16'd62538, 16'd17817, 16'd15327, 16'd9403, 16'd39076});
	test_expansion(128'he0a313a631c730596e2ab7e150700b29, {16'd31166, 16'd62466, 16'd42808, 16'd31369, 16'd30142, 16'd65244, 16'd11252, 16'd39536, 16'd50823, 16'd11906, 16'd46734, 16'd3831, 16'd33771, 16'd40314, 16'd57012, 16'd61259, 16'd41428, 16'd23056, 16'd30102, 16'd41753, 16'd56824, 16'd38512, 16'd7713, 16'd43353, 16'd1345, 16'd21363});
	test_expansion(128'h9101c38d408b4827e4fad94fc86d1e65, {16'd26034, 16'd11109, 16'd58320, 16'd10589, 16'd6121, 16'd19066, 16'd10759, 16'd26859, 16'd11907, 16'd13889, 16'd59381, 16'd52195, 16'd2381, 16'd63866, 16'd61745, 16'd37701, 16'd43691, 16'd33076, 16'd6996, 16'd7310, 16'd45185, 16'd26360, 16'd14101, 16'd40379, 16'd63704, 16'd39461});
	test_expansion(128'h6f141343df0e50cbc928f02f8054cbbc, {16'd61257, 16'd58416, 16'd65255, 16'd31388, 16'd19936, 16'd9365, 16'd36340, 16'd46950, 16'd14566, 16'd25724, 16'd33528, 16'd46531, 16'd49727, 16'd41683, 16'd14491, 16'd11972, 16'd7343, 16'd20483, 16'd32221, 16'd21765, 16'd25953, 16'd60026, 16'd60431, 16'd57328, 16'd61477, 16'd63208});
	test_expansion(128'h861202ca414cf62f0d1f2752345fe6ff, {16'd61790, 16'd13214, 16'd63061, 16'd32318, 16'd36426, 16'd46593, 16'd44285, 16'd61229, 16'd28361, 16'd51320, 16'd53019, 16'd5007, 16'd44948, 16'd31363, 16'd40767, 16'd56036, 16'd54278, 16'd22372, 16'd27992, 16'd40604, 16'd13463, 16'd46042, 16'd8347, 16'd29573, 16'd978, 16'd44876});
	test_expansion(128'h5ee9799ac55273eac0b71afa57d59d19, {16'd15296, 16'd55181, 16'd43610, 16'd20872, 16'd22355, 16'd20183, 16'd25388, 16'd8192, 16'd27022, 16'd42839, 16'd18915, 16'd59343, 16'd30736, 16'd49372, 16'd27716, 16'd53595, 16'd16394, 16'd13630, 16'd35688, 16'd28127, 16'd56618, 16'd59473, 16'd23326, 16'd39903, 16'd52222, 16'd50686});
	test_expansion(128'h185ab12fe9c7833d2b1e2cf2c6a26273, {16'd39823, 16'd1830, 16'd23989, 16'd48099, 16'd1442, 16'd3277, 16'd44114, 16'd18752, 16'd41929, 16'd52891, 16'd32244, 16'd41513, 16'd52703, 16'd13189, 16'd22947, 16'd23460, 16'd11810, 16'd46530, 16'd30162, 16'd58704, 16'd56266, 16'd30343, 16'd19502, 16'd51238, 16'd22185, 16'd55336});
	test_expansion(128'h8b8848ef885da57e3ee42f186367283a, {16'd24736, 16'd17532, 16'd55249, 16'd55448, 16'd43390, 16'd23910, 16'd44842, 16'd61283, 16'd30462, 16'd41220, 16'd20145, 16'd17369, 16'd54809, 16'd7783, 16'd35837, 16'd32315, 16'd29802, 16'd6765, 16'd24577, 16'd6831, 16'd7121, 16'd34332, 16'd45353, 16'd62087, 16'd10223, 16'd22004});
	test_expansion(128'h7c8b5fe4e79f7693ddf5d16bc2a4213f, {16'd4802, 16'd2518, 16'd65145, 16'd54264, 16'd11393, 16'd65415, 16'd38347, 16'd34441, 16'd5829, 16'd38726, 16'd52354, 16'd13405, 16'd51399, 16'd26490, 16'd34153, 16'd4666, 16'd55245, 16'd23299, 16'd54107, 16'd16873, 16'd19040, 16'd52760, 16'd47856, 16'd13888, 16'd25297, 16'd49698});
	test_expansion(128'hba2d80959f703032954c269eb7db3017, {16'd24318, 16'd34248, 16'd12281, 16'd15035, 16'd29965, 16'd27948, 16'd23257, 16'd22660, 16'd56070, 16'd22331, 16'd53022, 16'd6916, 16'd27036, 16'd16993, 16'd56466, 16'd35755, 16'd56447, 16'd52278, 16'd24111, 16'd12181, 16'd49026, 16'd51258, 16'd3876, 16'd17298, 16'd42184, 16'd47020});
	test_expansion(128'hb224926d25bd49178f15a58a495e524a, {16'd731, 16'd51364, 16'd51397, 16'd53048, 16'd41810, 16'd54802, 16'd11981, 16'd3936, 16'd7770, 16'd14459, 16'd18412, 16'd22234, 16'd24681, 16'd48612, 16'd26208, 16'd57112, 16'd18845, 16'd51192, 16'd52208, 16'd7461, 16'd32946, 16'd51222, 16'd7144, 16'd36939, 16'd59709, 16'd9032});
	test_expansion(128'hc14c26ee55776aa82a479ade2453f4d0, {16'd23529, 16'd22522, 16'd40625, 16'd52059, 16'd60763, 16'd30905, 16'd49647, 16'd56092, 16'd29671, 16'd54606, 16'd15513, 16'd33650, 16'd44775, 16'd50733, 16'd46736, 16'd20913, 16'd11143, 16'd39292, 16'd59311, 16'd4935, 16'd28432, 16'd28754, 16'd64352, 16'd19577, 16'd25736, 16'd58461});
	test_expansion(128'hc2cd483a2d6c1a9c40c069e7a7f79e19, {16'd27424, 16'd14554, 16'd23507, 16'd27111, 16'd43207, 16'd49235, 16'd26733, 16'd54967, 16'd9050, 16'd11414, 16'd11058, 16'd64484, 16'd608, 16'd64422, 16'd64232, 16'd9791, 16'd60534, 16'd265, 16'd56628, 16'd49011, 16'd28921, 16'd34039, 16'd46716, 16'd1207, 16'd37186, 16'd45949});
	test_expansion(128'haff823bf442123e310de9409504578d5, {16'd62663, 16'd9919, 16'd25965, 16'd26803, 16'd48083, 16'd1764, 16'd17101, 16'd25111, 16'd7638, 16'd19203, 16'd18128, 16'd52193, 16'd36636, 16'd40906, 16'd11141, 16'd36382, 16'd40788, 16'd14622, 16'd38288, 16'd35462, 16'd935, 16'd63560, 16'd18995, 16'd28689, 16'd62166, 16'd14328});
	test_expansion(128'hfd487bbed727782cfaef455aaa33745b, {16'd22650, 16'd4409, 16'd14358, 16'd54190, 16'd45768, 16'd43180, 16'd30006, 16'd21213, 16'd64528, 16'd16870, 16'd46549, 16'd2417, 16'd19736, 16'd39340, 16'd23588, 16'd48131, 16'd24223, 16'd44910, 16'd8373, 16'd31135, 16'd44710, 16'd43361, 16'd34437, 16'd54089, 16'd22864, 16'd64967});
	test_expansion(128'he2c9fd06eca1e0f02e0e7e2e59e5fbbf, {16'd14597, 16'd61662, 16'd32961, 16'd60097, 16'd31186, 16'd9392, 16'd53027, 16'd24983, 16'd44345, 16'd10503, 16'd46780, 16'd54095, 16'd50723, 16'd15417, 16'd3012, 16'd31215, 16'd18552, 16'd36737, 16'd30293, 16'd7920, 16'd7853, 16'd44455, 16'd40104, 16'd40903, 16'd13028, 16'd59872});
	test_expansion(128'hdbefccd351c2304463da6dadf26b2395, {16'd62577, 16'd47858, 16'd61023, 16'd49692, 16'd18532, 16'd15951, 16'd49237, 16'd63574, 16'd57951, 16'd16610, 16'd54821, 16'd12280, 16'd24269, 16'd55486, 16'd37418, 16'd6079, 16'd37401, 16'd58061, 16'd16394, 16'd36180, 16'd45639, 16'd9451, 16'd57973, 16'd60198, 16'd1031, 16'd37989});
	test_expansion(128'he9959a4762fe0dbaa16f2e57ff9c5bfc, {16'd56859, 16'd41751, 16'd14521, 16'd30642, 16'd941, 16'd15847, 16'd52577, 16'd58210, 16'd44787, 16'd15832, 16'd44615, 16'd53867, 16'd44853, 16'd55609, 16'd64998, 16'd56383, 16'd42473, 16'd8570, 16'd20554, 16'd38497, 16'd36835, 16'd61472, 16'd42806, 16'd751, 16'd43761, 16'd41804});
	test_expansion(128'hc8c47db19840c0422a813f51351f7b30, {16'd34537, 16'd41915, 16'd62711, 16'd32422, 16'd21368, 16'd25732, 16'd15832, 16'd12581, 16'd34698, 16'd18861, 16'd53210, 16'd11300, 16'd37041, 16'd25251, 16'd24905, 16'd33157, 16'd9554, 16'd32442, 16'd63020, 16'd65074, 16'd22630, 16'd12954, 16'd63200, 16'd6790, 16'd3424, 16'd4262});
	test_expansion(128'h370d92baca923e0584e93cd7dab582e9, {16'd10895, 16'd7041, 16'd31961, 16'd48543, 16'd64412, 16'd34181, 16'd4224, 16'd26780, 16'd62922, 16'd36875, 16'd21404, 16'd52496, 16'd12431, 16'd3119, 16'd4374, 16'd17866, 16'd59768, 16'd1207, 16'd32580, 16'd44566, 16'd14919, 16'd64177, 16'd24762, 16'd22503, 16'd57824, 16'd23949});
	test_expansion(128'h046042a0997ed0b61bfbe587df2d10ad, {16'd61425, 16'd2225, 16'd2837, 16'd44434, 16'd56046, 16'd60128, 16'd54124, 16'd51428, 16'd16741, 16'd19773, 16'd49702, 16'd5934, 16'd58239, 16'd58817, 16'd10693, 16'd24170, 16'd4820, 16'd15092, 16'd26778, 16'd26203, 16'd31418, 16'd15987, 16'd31554, 16'd12843, 16'd42984, 16'd23246});
	test_expansion(128'he14614f1657ae48955ea9dd7a2f11e58, {16'd49277, 16'd50706, 16'd53847, 16'd34770, 16'd15068, 16'd48638, 16'd46773, 16'd25592, 16'd14156, 16'd4724, 16'd7778, 16'd57156, 16'd3131, 16'd2706, 16'd19893, 16'd19822, 16'd33768, 16'd31620, 16'd26930, 16'd12348, 16'd22559, 16'd38190, 16'd37757, 16'd14252, 16'd12393, 16'd44324});
	test_expansion(128'h7939c5a9cbb8b9866b3eb62d5b18a55d, {16'd28655, 16'd14790, 16'd35308, 16'd38005, 16'd31772, 16'd11452, 16'd6401, 16'd16769, 16'd34282, 16'd9119, 16'd18542, 16'd21689, 16'd31714, 16'd13854, 16'd40396, 16'd45010, 16'd29857, 16'd27775, 16'd17790, 16'd29327, 16'd17021, 16'd41618, 16'd29351, 16'd21908, 16'd57524, 16'd24743});
	test_expansion(128'h65c07bb874a5ef833d0ee56b452db1f8, {16'd18436, 16'd62709, 16'd29291, 16'd33058, 16'd7869, 16'd49409, 16'd9284, 16'd6906, 16'd54987, 16'd46922, 16'd64646, 16'd47518, 16'd12832, 16'd27033, 16'd52204, 16'd39656, 16'd4309, 16'd58849, 16'd33031, 16'd30296, 16'd1364, 16'd53185, 16'd5476, 16'd26507, 16'd17704, 16'd42597});
	test_expansion(128'h996b643a90b73c352e42607145facfb2, {16'd32269, 16'd65012, 16'd23695, 16'd11250, 16'd34345, 16'd60921, 16'd53921, 16'd51009, 16'd57030, 16'd57054, 16'd30137, 16'd59026, 16'd36013, 16'd31866, 16'd47119, 16'd24535, 16'd45414, 16'd51320, 16'd23104, 16'd14595, 16'd15921, 16'd11236, 16'd27617, 16'd23721, 16'd26159, 16'd62843});
	test_expansion(128'h2dfe9ce5a9457c9d793845f693ab8085, {16'd30205, 16'd16892, 16'd11543, 16'd18182, 16'd38660, 16'd24991, 16'd16838, 16'd1232, 16'd43285, 16'd11134, 16'd5332, 16'd6441, 16'd24662, 16'd16753, 16'd55012, 16'd62475, 16'd34567, 16'd35539, 16'd65209, 16'd47122, 16'd33387, 16'd61116, 16'd15648, 16'd63430, 16'd4687, 16'd39102});
	test_expansion(128'h54a93bf18cac23435ed5d7e99b2c175b, {16'd1225, 16'd41049, 16'd43404, 16'd64729, 16'd57569, 16'd39511, 16'd39511, 16'd1515, 16'd6038, 16'd26402, 16'd747, 16'd11884, 16'd50272, 16'd59389, 16'd1352, 16'd35778, 16'd24590, 16'd40884, 16'd39662, 16'd58959, 16'd36420, 16'd13912, 16'd10632, 16'd44494, 16'd6282, 16'd19688});
	test_expansion(128'h2eda7e46c80cfe6a0dcca70f29716477, {16'd7110, 16'd34598, 16'd10403, 16'd42008, 16'd46252, 16'd13565, 16'd61916, 16'd19120, 16'd10776, 16'd23859, 16'd43759, 16'd39136, 16'd21955, 16'd8349, 16'd2968, 16'd26603, 16'd51430, 16'd26945, 16'd26042, 16'd62795, 16'd65382, 16'd20976, 16'd18295, 16'd3600, 16'd46183, 16'd11291});
	test_expansion(128'h310787cf8502a2c790ea8ab688580e9d, {16'd42996, 16'd15910, 16'd41977, 16'd16400, 16'd6472, 16'd45303, 16'd17953, 16'd2277, 16'd47843, 16'd64255, 16'd21076, 16'd33081, 16'd30266, 16'd37377, 16'd42250, 16'd30760, 16'd14353, 16'd484, 16'd32227, 16'd51174, 16'd6701, 16'd18521, 16'd53906, 16'd9379, 16'd11141, 16'd44921});
	test_expansion(128'h6c48dc84144e9410d09b65b8ab547459, {16'd27210, 16'd62820, 16'd52570, 16'd37296, 16'd64004, 16'd45934, 16'd40607, 16'd7893, 16'd54114, 16'd47176, 16'd21697, 16'd26397, 16'd62163, 16'd41176, 16'd43255, 16'd57719, 16'd49362, 16'd7340, 16'd59484, 16'd14648, 16'd5662, 16'd14289, 16'd47063, 16'd18182, 16'd1532, 16'd53096});
	test_expansion(128'hf379bb34fb6604972ed52a41a32e1541, {16'd48479, 16'd53833, 16'd1597, 16'd51474, 16'd4853, 16'd58793, 16'd29847, 16'd13615, 16'd14146, 16'd48136, 16'd51783, 16'd29489, 16'd57577, 16'd40606, 16'd43655, 16'd10579, 16'd16386, 16'd19532, 16'd57583, 16'd2056, 16'd16236, 16'd6199, 16'd22721, 16'd64998, 16'd64783, 16'd42276});
	test_expansion(128'h788d50818b60811badc474bab0deb64e, {16'd28151, 16'd2307, 16'd17516, 16'd56979, 16'd5319, 16'd38508, 16'd30290, 16'd24559, 16'd38231, 16'd46297, 16'd2216, 16'd64581, 16'd5630, 16'd1716, 16'd48894, 16'd11786, 16'd6327, 16'd7813, 16'd42729, 16'd63499, 16'd42833, 16'd45022, 16'd783, 16'd24401, 16'd42401, 16'd15329});
	test_expansion(128'h4010c31722130c84545340773facefa1, {16'd8201, 16'd26454, 16'd44734, 16'd1638, 16'd524, 16'd19386, 16'd45921, 16'd21182, 16'd35828, 16'd51050, 16'd28546, 16'd18455, 16'd35297, 16'd12888, 16'd29467, 16'd51297, 16'd14654, 16'd29892, 16'd59261, 16'd52599, 16'd55971, 16'd28329, 16'd43776, 16'd35062, 16'd30801, 16'd40778});
	test_expansion(128'hee6692c8dd044bb7336a80365d72a753, {16'd16483, 16'd50148, 16'd5647, 16'd45573, 16'd62340, 16'd22857, 16'd46814, 16'd42444, 16'd65032, 16'd25488, 16'd33957, 16'd46503, 16'd21593, 16'd7130, 16'd17992, 16'd47416, 16'd52042, 16'd11899, 16'd56821, 16'd49247, 16'd17481, 16'd43579, 16'd32763, 16'd58511, 16'd19592, 16'd39517});
	test_expansion(128'ha81f0a8b2fa82e5245979fff206a1fda, {16'd59096, 16'd3712, 16'd52566, 16'd1615, 16'd5816, 16'd25782, 16'd9486, 16'd12732, 16'd25120, 16'd44758, 16'd65107, 16'd28304, 16'd58970, 16'd55637, 16'd11341, 16'd37570, 16'd20133, 16'd31004, 16'd5517, 16'd14666, 16'd6284, 16'd52109, 16'd56337, 16'd39154, 16'd33234, 16'd58686});
	test_expansion(128'h7ed43df70e0a06a40f5dc28c453a06c4, {16'd36091, 16'd47281, 16'd783, 16'd37300, 16'd29059, 16'd6571, 16'd39178, 16'd62463, 16'd58098, 16'd42243, 16'd9872, 16'd26301, 16'd31411, 16'd12016, 16'd32517, 16'd29824, 16'd9314, 16'd58766, 16'd30607, 16'd47902, 16'd30891, 16'd30960, 16'd18216, 16'd43837, 16'd54240, 16'd21565});
	test_expansion(128'hafd0ab5be4a9f5112ed2581a7627a3bd, {16'd6105, 16'd54607, 16'd1457, 16'd62899, 16'd60020, 16'd19032, 16'd58777, 16'd5041, 16'd56696, 16'd45466, 16'd50079, 16'd59311, 16'd33856, 16'd41230, 16'd20974, 16'd55568, 16'd2443, 16'd21332, 16'd25608, 16'd12257, 16'd348, 16'd13189, 16'd51329, 16'd12746, 16'd26401, 16'd54083});
	test_expansion(128'h67603fa9c42ef5d525687f26e28be07d, {16'd50489, 16'd56823, 16'd31394, 16'd53955, 16'd37567, 16'd60899, 16'd11521, 16'd49211, 16'd35506, 16'd61359, 16'd16904, 16'd47009, 16'd8522, 16'd20804, 16'd65473, 16'd11609, 16'd16660, 16'd52312, 16'd28522, 16'd44528, 16'd3154, 16'd49446, 16'd46658, 16'd35039, 16'd8957, 16'd39512});
	test_expansion(128'hcc2726d5542dc798e6e8a25f696d2ce5, {16'd55005, 16'd20971, 16'd19479, 16'd24077, 16'd42686, 16'd12636, 16'd20679, 16'd49411, 16'd55183, 16'd29531, 16'd28474, 16'd31843, 16'd6879, 16'd50338, 16'd20645, 16'd53212, 16'd52880, 16'd48725, 16'd59158, 16'd11464, 16'd11230, 16'd15060, 16'd15856, 16'd26427, 16'd63373, 16'd58800});
	test_expansion(128'h9fd2953894b39e20dff652bb3bac1d53, {16'd34244, 16'd29474, 16'd12523, 16'd23763, 16'd65257, 16'd33890, 16'd16639, 16'd30340, 16'd5518, 16'd16364, 16'd40052, 16'd28532, 16'd56719, 16'd31329, 16'd18733, 16'd22401, 16'd16285, 16'd15691, 16'd58217, 16'd41443, 16'd7137, 16'd64581, 16'd44286, 16'd58145, 16'd5574, 16'd8939});
	test_expansion(128'h81ff6e12d634d6f93b1e44fb1e396d83, {16'd52687, 16'd23524, 16'd12259, 16'd18183, 16'd49763, 16'd50672, 16'd37595, 16'd58312, 16'd4724, 16'd4379, 16'd27964, 16'd52410, 16'd49998, 16'd41934, 16'd7989, 16'd7274, 16'd1126, 16'd61458, 16'd27002, 16'd31192, 16'd59864, 16'd3895, 16'd11444, 16'd35084, 16'd33919, 16'd6097});
	test_expansion(128'h65dd1be4cd08313afe4cdadb36058f15, {16'd60027, 16'd59895, 16'd17654, 16'd21610, 16'd40220, 16'd52363, 16'd44301, 16'd7947, 16'd13774, 16'd6662, 16'd25411, 16'd21941, 16'd59065, 16'd38291, 16'd60614, 16'd52703, 16'd50181, 16'd21183, 16'd29610, 16'd1508, 16'd50481, 16'd3992, 16'd34689, 16'd979, 16'd60570, 16'd15215});
	test_expansion(128'h6e3b77fe221a1cbe2fd3aba78d13f00e, {16'd64070, 16'd27383, 16'd31683, 16'd59377, 16'd24413, 16'd33987, 16'd23251, 16'd16288, 16'd58472, 16'd7698, 16'd26322, 16'd26540, 16'd44793, 16'd37614, 16'd28086, 16'd32595, 16'd15293, 16'd29741, 16'd28860, 16'd27365, 16'd34188, 16'd5721, 16'd18841, 16'd62291, 16'd32738, 16'd48797});
	test_expansion(128'h6b2a7ac31798e0bbcd8cef702a948e4f, {16'd25978, 16'd41658, 16'd62806, 16'd59944, 16'd12379, 16'd50305, 16'd13138, 16'd25610, 16'd49998, 16'd44179, 16'd23279, 16'd64256, 16'd56828, 16'd49345, 16'd33142, 16'd55926, 16'd22255, 16'd60896, 16'd24698, 16'd34889, 16'd54300, 16'd63846, 16'd32850, 16'd54368, 16'd64335, 16'd19286});
	test_expansion(128'h491e672fe048872eff782ce77070c94a, {16'd33333, 16'd46602, 16'd59450, 16'd47707, 16'd43057, 16'd29562, 16'd564, 16'd52701, 16'd14559, 16'd24633, 16'd30975, 16'd62081, 16'd15071, 16'd65472, 16'd64438, 16'd882, 16'd37911, 16'd50020, 16'd33860, 16'd27452, 16'd45907, 16'd54205, 16'd9867, 16'd26794, 16'd30460, 16'd33792});
	test_expansion(128'h164af319b3d366066157e0fe1d8d8d42, {16'd47070, 16'd45169, 16'd25687, 16'd4685, 16'd1048, 16'd23594, 16'd8352, 16'd61458, 16'd46141, 16'd11289, 16'd61305, 16'd52223, 16'd15311, 16'd53232, 16'd34720, 16'd13240, 16'd59362, 16'd7788, 16'd38619, 16'd18135, 16'd13241, 16'd34115, 16'd13638, 16'd6188, 16'd15725, 16'd15967});
	test_expansion(128'h7a9702e9e04e2c95f8e53c0c2d37a49e, {16'd13684, 16'd37833, 16'd32734, 16'd27440, 16'd49353, 16'd64528, 16'd37411, 16'd29788, 16'd11507, 16'd29022, 16'd23621, 16'd9999, 16'd60139, 16'd2361, 16'd57851, 16'd43707, 16'd32997, 16'd8958, 16'd44338, 16'd41480, 16'd30424, 16'd26828, 16'd49485, 16'd23308, 16'd24469, 16'd6214});
	test_expansion(128'h6f3410801a0d53cdfe3b18f9b1f75336, {16'd49430, 16'd4545, 16'd36348, 16'd9375, 16'd25307, 16'd27791, 16'd55118, 16'd42008, 16'd34874, 16'd38321, 16'd49230, 16'd32406, 16'd29920, 16'd27846, 16'd33726, 16'd37073, 16'd6968, 16'd31315, 16'd63796, 16'd11415, 16'd46528, 16'd17687, 16'd54863, 16'd46408, 16'd3627, 16'd43748});
	test_expansion(128'h024ba0a2b9a5df1034ac78f90bcd0f99, {16'd20524, 16'd63048, 16'd8487, 16'd34561, 16'd33923, 16'd34921, 16'd55815, 16'd12739, 16'd50446, 16'd18249, 16'd47582, 16'd28486, 16'd37243, 16'd7258, 16'd31760, 16'd26472, 16'd30858, 16'd34277, 16'd60802, 16'd5068, 16'd9862, 16'd11072, 16'd58044, 16'd35397, 16'd21528, 16'd30389});
	test_expansion(128'h9baaac0f67e376657ad0226dd62b7321, {16'd63199, 16'd61908, 16'd35280, 16'd52375, 16'd45011, 16'd22956, 16'd6767, 16'd32026, 16'd62683, 16'd27520, 16'd40382, 16'd19119, 16'd37295, 16'd45897, 16'd48982, 16'd807, 16'd65082, 16'd12369, 16'd46975, 16'd17223, 16'd21309, 16'd2469, 16'd21940, 16'd55147, 16'd35896, 16'd46292});
	test_expansion(128'h1e35935ed5622013ced5b414c0ae7658, {16'd49177, 16'd49313, 16'd58021, 16'd4731, 16'd62066, 16'd28984, 16'd6367, 16'd64432, 16'd11676, 16'd38204, 16'd58250, 16'd1030, 16'd49350, 16'd54206, 16'd39575, 16'd60471, 16'd52531, 16'd20244, 16'd53691, 16'd14494, 16'd54891, 16'd57301, 16'd2818, 16'd45986, 16'd31304, 16'd14913});
	test_expansion(128'ha9e18dd957d090dd1978fd4a4c0c11cd, {16'd43685, 16'd65282, 16'd61194, 16'd63158, 16'd59862, 16'd63937, 16'd50008, 16'd55197, 16'd41331, 16'd34998, 16'd39757, 16'd9556, 16'd27860, 16'd13425, 16'd51921, 16'd7079, 16'd50452, 16'd27073, 16'd40845, 16'd39072, 16'd24630, 16'd21416, 16'd6744, 16'd5707, 16'd28049, 16'd9720});
	test_expansion(128'h418684591f6164a1efacc52402c6fcbc, {16'd10918, 16'd1500, 16'd47227, 16'd40663, 16'd18474, 16'd24264, 16'd34805, 16'd56943, 16'd39916, 16'd8944, 16'd31578, 16'd1733, 16'd52021, 16'd46740, 16'd31710, 16'd51371, 16'd34701, 16'd55208, 16'd39734, 16'd32967, 16'd56471, 16'd23140, 16'd13238, 16'd36365, 16'd300, 16'd4892});
	test_expansion(128'h59085b7cb5978b2a100135bb48a80dfe, {16'd4417, 16'd56805, 16'd45155, 16'd16022, 16'd28094, 16'd39407, 16'd46755, 16'd15828, 16'd41257, 16'd20135, 16'd23663, 16'd39929, 16'd1026, 16'd65226, 16'd5394, 16'd54959, 16'd64910, 16'd34872, 16'd33886, 16'd17535, 16'd11075, 16'd32588, 16'd22587, 16'd48453, 16'd64192, 16'd52421});
	test_expansion(128'h5f607d0b2ed4f2c440b1bb51e60df77f, {16'd7993, 16'd41350, 16'd4946, 16'd23711, 16'd22710, 16'd31088, 16'd42151, 16'd60772, 16'd3460, 16'd44234, 16'd38830, 16'd24451, 16'd46461, 16'd60052, 16'd65022, 16'd55481, 16'd11754, 16'd21240, 16'd20136, 16'd55362, 16'd27754, 16'd24334, 16'd39932, 16'd10118, 16'd28937, 16'd23172});
	test_expansion(128'h8d0373e1fac735d2c672e0d037fafa18, {16'd38528, 16'd1772, 16'd58054, 16'd6238, 16'd53565, 16'd11933, 16'd21873, 16'd64618, 16'd40152, 16'd54019, 16'd23674, 16'd12941, 16'd508, 16'd10934, 16'd18348, 16'd54724, 16'd12956, 16'd58138, 16'd6043, 16'd29241, 16'd15304, 16'd64043, 16'd52557, 16'd57229, 16'd39710, 16'd33431});
	test_expansion(128'hc95e76efdb936f42ff7b618b719d7c6a, {16'd21837, 16'd28800, 16'd38746, 16'd91, 16'd12454, 16'd61367, 16'd29605, 16'd34890, 16'd15338, 16'd9504, 16'd39105, 16'd37090, 16'd32530, 16'd62352, 16'd49201, 16'd35706, 16'd21052, 16'd59764, 16'd1523, 16'd37327, 16'd57128, 16'd10185, 16'd57954, 16'd10888, 16'd43717, 16'd36217});
	test_expansion(128'h433529dc28a90dbc02400fe14b913251, {16'd23455, 16'd6852, 16'd42636, 16'd43584, 16'd6158, 16'd4502, 16'd37382, 16'd32854, 16'd30486, 16'd25137, 16'd4759, 16'd15831, 16'd29770, 16'd12657, 16'd224, 16'd56689, 16'd35419, 16'd27239, 16'd9772, 16'd52400, 16'd16128, 16'd48500, 16'd43980, 16'd5986, 16'd60702, 16'd55558});
	test_expansion(128'he583749d165f0e69bbbbaa12f4a10cb9, {16'd56078, 16'd64126, 16'd58054, 16'd32587, 16'd1439, 16'd37017, 16'd35394, 16'd45603, 16'd39195, 16'd9371, 16'd6180, 16'd20086, 16'd6613, 16'd24425, 16'd2767, 16'd29014, 16'd33243, 16'd64074, 16'd63162, 16'd18957, 16'd39175, 16'd42300, 16'd20557, 16'd1052, 16'd64885, 16'd36990});
	test_expansion(128'h08bfd908567089b49ce7c5da5a4e2673, {16'd63966, 16'd50967, 16'd32624, 16'd38782, 16'd28640, 16'd6599, 16'd29287, 16'd16078, 16'd49663, 16'd4219, 16'd3105, 16'd55348, 16'd39090, 16'd10384, 16'd7570, 16'd13413, 16'd9795, 16'd34080, 16'd51167, 16'd44559, 16'd42343, 16'd53502, 16'd13154, 16'd5693, 16'd39343, 16'd15867});
	test_expansion(128'hc5ea8810da589b98fa1b39a2cdfa282a, {16'd57430, 16'd16041, 16'd31811, 16'd12276, 16'd617, 16'd5047, 16'd46526, 16'd50599, 16'd2526, 16'd23558, 16'd8344, 16'd18283, 16'd29176, 16'd34853, 16'd64788, 16'd34979, 16'd34722, 16'd60677, 16'd3186, 16'd10305, 16'd25025, 16'd41613, 16'd63874, 16'd42132, 16'd57397, 16'd63080});
	test_expansion(128'hdec4fcbda0074ef67ecee993f6920cec, {16'd42175, 16'd43834, 16'd59887, 16'd4184, 16'd10476, 16'd16384, 16'd2151, 16'd29687, 16'd33964, 16'd16152, 16'd51888, 16'd12985, 16'd10532, 16'd5495, 16'd51385, 16'd63457, 16'd25711, 16'd23204, 16'd35699, 16'd20762, 16'd54232, 16'd4680, 16'd22919, 16'd15277, 16'd1251, 16'd56854});
	test_expansion(128'h0eab762713b5c9dcb11728251cbd18c9, {16'd2116, 16'd31083, 16'd54, 16'd64567, 16'd27457, 16'd56238, 16'd31455, 16'd63463, 16'd7343, 16'd21619, 16'd5052, 16'd28171, 16'd16207, 16'd39073, 16'd37236, 16'd27754, 16'd26653, 16'd57606, 16'd50753, 16'd1449, 16'd10934, 16'd18777, 16'd9020, 16'd61743, 16'd52551, 16'd61095});
	test_expansion(128'h041e72b0817f52ea40453167d05357ea, {16'd48942, 16'd23274, 16'd12317, 16'd59295, 16'd16904, 16'd1320, 16'd55006, 16'd15411, 16'd58441, 16'd8702, 16'd64905, 16'd56581, 16'd50641, 16'd24869, 16'd53575, 16'd19618, 16'd60418, 16'd2813, 16'd63335, 16'd8532, 16'd35533, 16'd18946, 16'd56597, 16'd19297, 16'd37242, 16'd48824});
	test_expansion(128'h3098c307a81ab623eef19993c98c6753, {16'd50469, 16'd58186, 16'd34116, 16'd49314, 16'd21845, 16'd49622, 16'd34836, 16'd33080, 16'd24067, 16'd41974, 16'd44183, 16'd53549, 16'd3337, 16'd11563, 16'd30233, 16'd12145, 16'd56588, 16'd37975, 16'd17364, 16'd30795, 16'd18423, 16'd1435, 16'd869, 16'd23801, 16'd44055, 16'd43740});
	test_expansion(128'h7d386fcfb90234e9f59c664c2894d00f, {16'd29501, 16'd51563, 16'd11443, 16'd60510, 16'd56917, 16'd54959, 16'd10171, 16'd52923, 16'd16341, 16'd26149, 16'd10502, 16'd28531, 16'd57968, 16'd49482, 16'd15373, 16'd31562, 16'd61490, 16'd8369, 16'd5151, 16'd20721, 16'd38779, 16'd46704, 16'd57477, 16'd11962, 16'd12958, 16'd985});
	test_expansion(128'heb95357396fbbfe378fb0ba5f4e4f5d0, {16'd24422, 16'd47188, 16'd61896, 16'd50068, 16'd21668, 16'd45182, 16'd51418, 16'd43592, 16'd55727, 16'd26794, 16'd33896, 16'd51836, 16'd27989, 16'd62073, 16'd43552, 16'd51337, 16'd63011, 16'd43041, 16'd60342, 16'd42849, 16'd27391, 16'd6865, 16'd56354, 16'd30124, 16'd22999, 16'd28125});
	test_expansion(128'h8a66430a5c57c289761ff3e932b4ecf8, {16'd53189, 16'd9433, 16'd44414, 16'd10133, 16'd41966, 16'd10412, 16'd45378, 16'd29457, 16'd48561, 16'd50392, 16'd36685, 16'd55463, 16'd57302, 16'd25684, 16'd23194, 16'd20438, 16'd35268, 16'd13340, 16'd23905, 16'd62688, 16'd40739, 16'd47919, 16'd40812, 16'd36495, 16'd13586, 16'd39816});
	test_expansion(128'h3d0c621d1f0ad2d39d19b0f7291f3827, {16'd49591, 16'd58268, 16'd62399, 16'd22629, 16'd19632, 16'd44852, 16'd28509, 16'd11502, 16'd20328, 16'd53116, 16'd48239, 16'd21618, 16'd30898, 16'd51558, 16'd53768, 16'd28923, 16'd54729, 16'd11316, 16'd36878, 16'd21687, 16'd48506, 16'd39311, 16'd36588, 16'd41828, 16'd26557, 16'd63740});
	test_expansion(128'h496315214eac9044955eac7122023aaa, {16'd19498, 16'd58754, 16'd16974, 16'd23057, 16'd64532, 16'd29946, 16'd529, 16'd5692, 16'd39826, 16'd10439, 16'd832, 16'd38209, 16'd50552, 16'd15868, 16'd41395, 16'd42821, 16'd63918, 16'd63561, 16'd61266, 16'd33155, 16'd21405, 16'd45286, 16'd39971, 16'd58480, 16'd22414, 16'd18776});
	test_expansion(128'hac1e8b0a9d7ef5e4045058edd46f230c, {16'd34148, 16'd63127, 16'd41796, 16'd56132, 16'd41914, 16'd9016, 16'd33072, 16'd42026, 16'd57224, 16'd60475, 16'd1133, 16'd23218, 16'd53828, 16'd44170, 16'd37098, 16'd30878, 16'd16486, 16'd6010, 16'd28706, 16'd4339, 16'd46969, 16'd3513, 16'd9564, 16'd53544, 16'd62004, 16'd15332});
	test_expansion(128'h3a7997ab2ca6c2902c225fa1177f6b46, {16'd44280, 16'd52459, 16'd53691, 16'd61749, 16'd56142, 16'd5997, 16'd26130, 16'd60305, 16'd16648, 16'd65509, 16'd19125, 16'd34103, 16'd50299, 16'd24734, 16'd51058, 16'd9021, 16'd17706, 16'd40919, 16'd37793, 16'd21058, 16'd18932, 16'd46596, 16'd37392, 16'd48087, 16'd55448, 16'd23080});
	test_expansion(128'hf5d870a77c26f4ec128c342d4abd3fbb, {16'd64009, 16'd53140, 16'd32776, 16'd61683, 16'd53138, 16'd37483, 16'd28822, 16'd45393, 16'd13450, 16'd60935, 16'd24160, 16'd19003, 16'd15074, 16'd64213, 16'd45594, 16'd6526, 16'd54590, 16'd39366, 16'd40687, 16'd43443, 16'd29581, 16'd11657, 16'd7787, 16'd13033, 16'd30234, 16'd14916});
	test_expansion(128'hb225574a59a588b5f497aa5a241c98f5, {16'd50797, 16'd57223, 16'd9444, 16'd12039, 16'd55740, 16'd4400, 16'd15043, 16'd43431, 16'd34293, 16'd41185, 16'd16715, 16'd48903, 16'd61825, 16'd59727, 16'd45148, 16'd45577, 16'd42521, 16'd63548, 16'd7767, 16'd52321, 16'd3636, 16'd16059, 16'd28597, 16'd52443, 16'd22314, 16'd23810});
	test_expansion(128'heb8c4a4a1d4f1d0f25cb4e420a41e700, {16'd23899, 16'd36907, 16'd14409, 16'd6788, 16'd64087, 16'd5731, 16'd11077, 16'd5358, 16'd17089, 16'd17254, 16'd63694, 16'd48964, 16'd47029, 16'd26811, 16'd43653, 16'd60943, 16'd12630, 16'd52844, 16'd29954, 16'd29791, 16'd54615, 16'd24099, 16'd23748, 16'd13462, 16'd51114, 16'd19793});
	test_expansion(128'h386620706586faf600134d9c0c299f48, {16'd51496, 16'd43325, 16'd15742, 16'd7664, 16'd10056, 16'd9973, 16'd52949, 16'd7829, 16'd33424, 16'd7743, 16'd26177, 16'd7358, 16'd37125, 16'd53847, 16'd55760, 16'd18567, 16'd20125, 16'd31564, 16'd59601, 16'd54511, 16'd52518, 16'd32291, 16'd13490, 16'd11036, 16'd54201, 16'd32681});
	test_expansion(128'h8736564cf732a39a25968e40fec21e44, {16'd38889, 16'd38443, 16'd61916, 16'd64113, 16'd31517, 16'd18892, 16'd33646, 16'd27633, 16'd37952, 16'd41914, 16'd2344, 16'd39809, 16'd39108, 16'd33704, 16'd51245, 16'd4729, 16'd33626, 16'd61306, 16'd23946, 16'd25792, 16'd28713, 16'd18876, 16'd48465, 16'd57303, 16'd12877, 16'd34773});
	test_expansion(128'hb98c7bc6f5ae6223e3a958e8aef284ff, {16'd18500, 16'd33057, 16'd19372, 16'd29192, 16'd60900, 16'd41137, 16'd22999, 16'd40669, 16'd38532, 16'd17779, 16'd44097, 16'd32422, 16'd54319, 16'd38912, 16'd50075, 16'd38402, 16'd17923, 16'd62238, 16'd55851, 16'd62571, 16'd41081, 16'd2579, 16'd8497, 16'd17337, 16'd35568, 16'd65457});
	test_expansion(128'h97fa194a67563d1fabf5bf9de57a5e73, {16'd42947, 16'd63656, 16'd13128, 16'd38554, 16'd45332, 16'd27909, 16'd53658, 16'd56098, 16'd47439, 16'd36975, 16'd15497, 16'd6950, 16'd37954, 16'd14904, 16'd55128, 16'd32630, 16'd35374, 16'd35315, 16'd6374, 16'd17052, 16'd32982, 16'd27267, 16'd2867, 16'd22598, 16'd10838, 16'd10970});
	test_expansion(128'h22638c7411814b86c80bb8e240d799de, {16'd26252, 16'd56482, 16'd33458, 16'd54271, 16'd40791, 16'd36705, 16'd64087, 16'd16430, 16'd42135, 16'd42738, 16'd57064, 16'd60813, 16'd47327, 16'd39779, 16'd10599, 16'd20711, 16'd15071, 16'd100, 16'd25014, 16'd46885, 16'd20981, 16'd19048, 16'd56482, 16'd33173, 16'd34927, 16'd41702});
	test_expansion(128'he8e98c3485e87d3d18dcf61c65489685, {16'd31537, 16'd36329, 16'd12760, 16'd8737, 16'd19889, 16'd56370, 16'd45277, 16'd57995, 16'd40604, 16'd51811, 16'd22510, 16'd26579, 16'd56398, 16'd18913, 16'd43643, 16'd18420, 16'd26802, 16'd7809, 16'd55892, 16'd48418, 16'd39512, 16'd10131, 16'd35717, 16'd50582, 16'd52802, 16'd56107});
	test_expansion(128'h5b5c9c20346c8db958223bd9422868ba, {16'd35512, 16'd60907, 16'd27713, 16'd22447, 16'd1168, 16'd55139, 16'd65202, 16'd57567, 16'd21485, 16'd47684, 16'd35933, 16'd36760, 16'd41158, 16'd3903, 16'd54512, 16'd7809, 16'd12587, 16'd8488, 16'd21066, 16'd39906, 16'd53767, 16'd18020, 16'd22440, 16'd3349, 16'd37770, 16'd58262});
	test_expansion(128'hafa20212ceb9180931d290194145728d, {16'd23465, 16'd2531, 16'd44132, 16'd26487, 16'd13122, 16'd31498, 16'd323, 16'd57542, 16'd17043, 16'd4286, 16'd22491, 16'd17887, 16'd59870, 16'd35942, 16'd1878, 16'd10229, 16'd54510, 16'd9354, 16'd22440, 16'd15324, 16'd8063, 16'd34040, 16'd20477, 16'd34847, 16'd9710, 16'd43997});
	test_expansion(128'h14cf0f42748071f4f6efe919857aac89, {16'd4417, 16'd10439, 16'd49963, 16'd24199, 16'd58386, 16'd64397, 16'd41263, 16'd58485, 16'd7656, 16'd32154, 16'd207, 16'd6985, 16'd2697, 16'd45480, 16'd26426, 16'd16467, 16'd33947, 16'd38956, 16'd4020, 16'd59793, 16'd60235, 16'd59290, 16'd24862, 16'd47902, 16'd44795, 16'd38827});
	test_expansion(128'h629f4866169140f43c0894f0da2e6907, {16'd44619, 16'd2370, 16'd46615, 16'd32517, 16'd6339, 16'd11337, 16'd39481, 16'd5457, 16'd46262, 16'd62898, 16'd49059, 16'd30755, 16'd62931, 16'd44167, 16'd41854, 16'd1254, 16'd15798, 16'd10779, 16'd37723, 16'd61178, 16'd8968, 16'd33916, 16'd40451, 16'd18542, 16'd54268, 16'd7686});
	test_expansion(128'hb3899c6045c2885fefef530ea7b740ba, {16'd3116, 16'd52054, 16'd6793, 16'd27828, 16'd29089, 16'd30957, 16'd59420, 16'd129, 16'd23326, 16'd44968, 16'd43027, 16'd35772, 16'd41399, 16'd44061, 16'd65071, 16'd8793, 16'd24600, 16'd38810, 16'd22775, 16'd35106, 16'd24413, 16'd27096, 16'd48842, 16'd51224, 16'd64948, 16'd60785});
	test_expansion(128'h168fe37c0da1c2e632579b188ffd7932, {16'd61619, 16'd26358, 16'd33766, 16'd20923, 16'd56640, 16'd21476, 16'd35828, 16'd58636, 16'd6419, 16'd39334, 16'd49627, 16'd17838, 16'd36560, 16'd15945, 16'd37400, 16'd39132, 16'd28617, 16'd22527, 16'd20765, 16'd51887, 16'd21212, 16'd21567, 16'd29393, 16'd20237, 16'd13619, 16'd62601});
	test_expansion(128'hff5a5d2fdf5173819ca2eb5631f2e282, {16'd54045, 16'd10133, 16'd58552, 16'd43863, 16'd17230, 16'd1787, 16'd4526, 16'd35049, 16'd20988, 16'd57225, 16'd30410, 16'd2143, 16'd5159, 16'd9320, 16'd22048, 16'd31407, 16'd58100, 16'd32580, 16'd19723, 16'd28249, 16'd8588, 16'd33762, 16'd62347, 16'd25415, 16'd13081, 16'd19798});
	test_expansion(128'hec225f9fdff60ce7b5be623292167878, {16'd65093, 16'd10172, 16'd44153, 16'd23771, 16'd18925, 16'd55446, 16'd27303, 16'd16945, 16'd37027, 16'd63360, 16'd42130, 16'd11153, 16'd41900, 16'd20128, 16'd17663, 16'd19086, 16'd47723, 16'd11734, 16'd3721, 16'd25916, 16'd24973, 16'd52987, 16'd42223, 16'd48775, 16'd41509, 16'd22570});
	test_expansion(128'h7c64f96264a9162b0a7a104bddd1f22e, {16'd61265, 16'd59392, 16'd53077, 16'd10920, 16'd48237, 16'd28503, 16'd65264, 16'd49782, 16'd43278, 16'd51924, 16'd41552, 16'd46549, 16'd37938, 16'd4896, 16'd58500, 16'd24379, 16'd42155, 16'd7158, 16'd39676, 16'd9760, 16'd61022, 16'd29488, 16'd18046, 16'd39573, 16'd55594, 16'd17116});
	test_expansion(128'h62c521e3ee22e227d97504f97f14cbbc, {16'd51458, 16'd63394, 16'd53266, 16'd15561, 16'd4482, 16'd27497, 16'd15941, 16'd59074, 16'd49972, 16'd50319, 16'd59601, 16'd7942, 16'd22778, 16'd33578, 16'd30684, 16'd56661, 16'd58653, 16'd5246, 16'd12057, 16'd50853, 16'd64010, 16'd56327, 16'd62111, 16'd54728, 16'd49222, 16'd37647});
	test_expansion(128'h9d7ee4befd51714fcd6599908cfa3e5f, {16'd40342, 16'd4091, 16'd44262, 16'd49550, 16'd25446, 16'd62043, 16'd8485, 16'd63475, 16'd11326, 16'd22696, 16'd51720, 16'd36678, 16'd57575, 16'd125, 16'd61098, 16'd2147, 16'd16785, 16'd48713, 16'd56647, 16'd49866, 16'd19101, 16'd55593, 16'd39421, 16'd53519, 16'd27279, 16'd49530});
	test_expansion(128'hec9d71660c7c9b4363a99850b8fd4f76, {16'd38033, 16'd31817, 16'd2054, 16'd30111, 16'd39416, 16'd7116, 16'd45033, 16'd26755, 16'd13644, 16'd60142, 16'd45154, 16'd17090, 16'd24461, 16'd8342, 16'd23462, 16'd19092, 16'd31175, 16'd8993, 16'd10936, 16'd12321, 16'd54455, 16'd16067, 16'd56528, 16'd17422, 16'd3104, 16'd23756});
	test_expansion(128'h9bf239e101c8f34dcb6609d7a422edc6, {16'd43448, 16'd63198, 16'd21447, 16'd59203, 16'd18001, 16'd10804, 16'd1157, 16'd61519, 16'd18917, 16'd30356, 16'd54906, 16'd62378, 16'd53270, 16'd29585, 16'd5698, 16'd20646, 16'd27339, 16'd52810, 16'd52929, 16'd49567, 16'd38353, 16'd39730, 16'd27420, 16'd3623, 16'd36176, 16'd14590});
	test_expansion(128'h030a0e5f5c349e9902a2ea8f0bc99f95, {16'd2145, 16'd44893, 16'd41304, 16'd48601, 16'd18683, 16'd27412, 16'd20414, 16'd44547, 16'd12408, 16'd36576, 16'd7103, 16'd19347, 16'd31538, 16'd23487, 16'd26557, 16'd38119, 16'd38603, 16'd36926, 16'd36396, 16'd44740, 16'd20087, 16'd33146, 16'd2112, 16'd62162, 16'd44465, 16'd14095});
	test_expansion(128'h68b4d53783a74daf877d2a5798e72ae3, {16'd4268, 16'd40853, 16'd19460, 16'd20538, 16'd17760, 16'd14626, 16'd7541, 16'd44879, 16'd24150, 16'd61507, 16'd38904, 16'd15396, 16'd5012, 16'd27376, 16'd1070, 16'd41923, 16'd7689, 16'd14120, 16'd17384, 16'd11371, 16'd63430, 16'd43880, 16'd22230, 16'd54186, 16'd46086, 16'd42135});
	test_expansion(128'h93d072fbfc36c5432fc75a05f006ee0b, {16'd43447, 16'd56736, 16'd7647, 16'd16923, 16'd41010, 16'd48415, 16'd13504, 16'd28125, 16'd6612, 16'd55446, 16'd52205, 16'd43970, 16'd6711, 16'd21466, 16'd40604, 16'd25108, 16'd41248, 16'd60228, 16'd4024, 16'd304, 16'd43623, 16'd23722, 16'd39752, 16'd64379, 16'd3711, 16'd35894});
	test_expansion(128'haf4e6f97cba474161d2d6ab340685ea0, {16'd19930, 16'd9698, 16'd23964, 16'd1412, 16'd4381, 16'd45475, 16'd55727, 16'd59163, 16'd13768, 16'd28006, 16'd29779, 16'd38975, 16'd14966, 16'd36983, 16'd27865, 16'd38219, 16'd15747, 16'd14007, 16'd31613, 16'd3064, 16'd57925, 16'd63040, 16'd36396, 16'd55942, 16'd1926, 16'd34258});
	test_expansion(128'h57f6983b9288f1f5fca288265b39b627, {16'd22445, 16'd19587, 16'd42099, 16'd17048, 16'd22375, 16'd44723, 16'd60856, 16'd33686, 16'd27321, 16'd40659, 16'd51689, 16'd42013, 16'd7239, 16'd61626, 16'd3279, 16'd38624, 16'd3781, 16'd31340, 16'd23470, 16'd19555, 16'd62149, 16'd506, 16'd13795, 16'd40991, 16'd6093, 16'd26861});
	test_expansion(128'h505cf6232c49a871d1449a18d780470e, {16'd28925, 16'd31971, 16'd48086, 16'd17871, 16'd30601, 16'd41654, 16'd39301, 16'd49582, 16'd39099, 16'd28949, 16'd33470, 16'd63084, 16'd51907, 16'd45198, 16'd17122, 16'd14937, 16'd15196, 16'd56028, 16'd30984, 16'd5496, 16'd51137, 16'd4328, 16'd59169, 16'd26956, 16'd16338, 16'd49069});
	test_expansion(128'hbf7fdd3275ac79805080836c633fa8b7, {16'd20079, 16'd21602, 16'd43052, 16'd61910, 16'd39324, 16'd8877, 16'd16055, 16'd30341, 16'd59451, 16'd36180, 16'd36513, 16'd58898, 16'd64703, 16'd28372, 16'd18990, 16'd18512, 16'd28547, 16'd46374, 16'd11030, 16'd45952, 16'd8950, 16'd37114, 16'd44378, 16'd8286, 16'd9019, 16'd16837});
	test_expansion(128'h8f04698260788483babc4736dbd1c4b9, {16'd9546, 16'd51867, 16'd22562, 16'd16357, 16'd25171, 16'd22229, 16'd36867, 16'd50150, 16'd57729, 16'd58095, 16'd42741, 16'd63507, 16'd50344, 16'd56796, 16'd6626, 16'd62701, 16'd21674, 16'd45787, 16'd52584, 16'd34844, 16'd6101, 16'd14395, 16'd43092, 16'd33622, 16'd36846, 16'd60850});
	test_expansion(128'h2af9df1865e75e6f3d7b7e0dd40847e2, {16'd34120, 16'd58406, 16'd19677, 16'd38866, 16'd62096, 16'd47523, 16'd28572, 16'd13333, 16'd50112, 16'd58547, 16'd39502, 16'd19428, 16'd6281, 16'd24040, 16'd61781, 16'd41721, 16'd48775, 16'd41436, 16'd36068, 16'd25254, 16'd59181, 16'd33393, 16'd30821, 16'd38781, 16'd19805, 16'd58383});
	test_expansion(128'hb726059faca58b6e51b055b128cee921, {16'd28895, 16'd16098, 16'd4179, 16'd28933, 16'd5945, 16'd30687, 16'd39516, 16'd53209, 16'd34156, 16'd57406, 16'd62727, 16'd35918, 16'd35065, 16'd14231, 16'd14752, 16'd41888, 16'd51565, 16'd33090, 16'd4195, 16'd29751, 16'd62150, 16'd39718, 16'd33396, 16'd33038, 16'd48413, 16'd14250});
	test_expansion(128'h83049bef11600f3d4e344239cd92361e, {16'd19611, 16'd34525, 16'd59596, 16'd27230, 16'd7719, 16'd47367, 16'd14154, 16'd12259, 16'd22557, 16'd16425, 16'd11051, 16'd62475, 16'd29596, 16'd40151, 16'd37674, 16'd39203, 16'd47245, 16'd59413, 16'd13259, 16'd56771, 16'd38236, 16'd34861, 16'd53266, 16'd17754, 16'd40620, 16'd35118});
	test_expansion(128'hed5a99cc8fa186afe2fdaebab01e828a, {16'd55272, 16'd31571, 16'd65339, 16'd46625, 16'd29246, 16'd43693, 16'd8535, 16'd64106, 16'd42561, 16'd35820, 16'd58457, 16'd43217, 16'd5635, 16'd50372, 16'd10854, 16'd2767, 16'd49054, 16'd57397, 16'd56011, 16'd47722, 16'd22723, 16'd35557, 16'd47582, 16'd1876, 16'd4706, 16'd28622});
	test_expansion(128'h6111da4cc2801d1d6b6b20e73a00debe, {16'd65362, 16'd35366, 16'd37493, 16'd27755, 16'd46874, 16'd44664, 16'd9778, 16'd41715, 16'd15516, 16'd14595, 16'd22874, 16'd63162, 16'd63795, 16'd51158, 16'd58203, 16'd39840, 16'd32682, 16'd39543, 16'd64102, 16'd60198, 16'd11653, 16'd7450, 16'd3636, 16'd3214, 16'd5123, 16'd20623});
	test_expansion(128'hdbc1fcdab851aa7717fd6a8758e70b62, {16'd11475, 16'd51594, 16'd622, 16'd15426, 16'd6244, 16'd47440, 16'd36550, 16'd33675, 16'd65038, 16'd50711, 16'd35582, 16'd41883, 16'd3445, 16'd39936, 16'd31601, 16'd59021, 16'd551, 16'd9196, 16'd22153, 16'd57149, 16'd41344, 16'd34093, 16'd24033, 16'd30236, 16'd49457, 16'd61764});
	test_expansion(128'hc040b58c9cc84462c4153a74d3ec96ea, {16'd22367, 16'd60441, 16'd61522, 16'd31225, 16'd38345, 16'd36404, 16'd64590, 16'd4922, 16'd55036, 16'd23555, 16'd58283, 16'd36134, 16'd10658, 16'd20641, 16'd63860, 16'd54417, 16'd18032, 16'd36002, 16'd41983, 16'd58176, 16'd5037, 16'd45540, 16'd35606, 16'd65007, 16'd6170, 16'd31185});
	test_expansion(128'h7b90c952ab85d9fc3198f1819318f04f, {16'd4561, 16'd3862, 16'd43565, 16'd9690, 16'd593, 16'd49622, 16'd44260, 16'd9445, 16'd44675, 16'd42859, 16'd41005, 16'd39298, 16'd29684, 16'd57908, 16'd38550, 16'd47912, 16'd13012, 16'd2934, 16'd36212, 16'd40510, 16'd54696, 16'd13710, 16'd4413, 16'd31555, 16'd18681, 16'd41263});
	test_expansion(128'h7d91e098c993a9ac6fc7603400663e44, {16'd11780, 16'd18079, 16'd31778, 16'd47204, 16'd24022, 16'd7685, 16'd60553, 16'd46829, 16'd40476, 16'd8541, 16'd28271, 16'd9207, 16'd49568, 16'd29236, 16'd57929, 16'd32565, 16'd40691, 16'd51771, 16'd51615, 16'd50243, 16'd1642, 16'd48805, 16'd49040, 16'd11599, 16'd8279, 16'd22621});
	test_expansion(128'hfb52db8aafb8ad224218af42d52f9ac1, {16'd35820, 16'd29974, 16'd63541, 16'd9760, 16'd17606, 16'd33136, 16'd7060, 16'd2196, 16'd55623, 16'd28379, 16'd17529, 16'd8988, 16'd34358, 16'd65348, 16'd6689, 16'd56684, 16'd40398, 16'd30527, 16'd16938, 16'd44601, 16'd8568, 16'd460, 16'd59365, 16'd21924, 16'd30053, 16'd52070});
	test_expansion(128'h6cde1f6f1224bd66c768226bdfaccc55, {16'd42116, 16'd1262, 16'd29918, 16'd47180, 16'd57382, 16'd18637, 16'd710, 16'd29542, 16'd10939, 16'd28704, 16'd53664, 16'd7619, 16'd51495, 16'd33793, 16'd1752, 16'd20889, 16'd5329, 16'd11239, 16'd46895, 16'd55786, 16'd50607, 16'd41949, 16'd40547, 16'd29561, 16'd56251, 16'd21705});
	test_expansion(128'h20c907ebadc0ff9db2fc02a0119a9f6b, {16'd23282, 16'd24102, 16'd24478, 16'd43999, 16'd54107, 16'd2552, 16'd39329, 16'd26398, 16'd44532, 16'd29263, 16'd13238, 16'd19473, 16'd25920, 16'd49282, 16'd32238, 16'd51273, 16'd60780, 16'd52423, 16'd14287, 16'd40598, 16'd5393, 16'd5895, 16'd32402, 16'd42250, 16'd28278, 16'd4112});
	test_expansion(128'h82604f42be92975c76e2b6b6b0d7bd8d, {16'd24845, 16'd55394, 16'd46328, 16'd38222, 16'd13039, 16'd46071, 16'd42105, 16'd44014, 16'd35562, 16'd56078, 16'd64270, 16'd30228, 16'd11893, 16'd32913, 16'd50365, 16'd53462, 16'd30637, 16'd15358, 16'd6152, 16'd29740, 16'd57987, 16'd54818, 16'd62622, 16'd50370, 16'd12412, 16'd9052});
	test_expansion(128'h6be08aeb467262f4a292b114089ef2c1, {16'd44148, 16'd53768, 16'd19969, 16'd3078, 16'd30094, 16'd7598, 16'd50160, 16'd39101, 16'd48115, 16'd24845, 16'd45777, 16'd45575, 16'd27277, 16'd49685, 16'd20402, 16'd45453, 16'd47878, 16'd42919, 16'd17327, 16'd40031, 16'd64026, 16'd29284, 16'd34204, 16'd47343, 16'd31026, 16'd29727});
	test_expansion(128'h073380e6cd7ccbfc634901629e2247e3, {16'd51382, 16'd47090, 16'd44607, 16'd2097, 16'd16457, 16'd52326, 16'd9592, 16'd40744, 16'd45289, 16'd45470, 16'd12023, 16'd28168, 16'd54250, 16'd60084, 16'd15937, 16'd2915, 16'd18643, 16'd5107, 16'd34001, 16'd29403, 16'd25870, 16'd38314, 16'd35753, 16'd20922, 16'd26740, 16'd46901});
	test_expansion(128'h5fff34e35b1a7121e7ea9b01bc01da6b, {16'd21957, 16'd17223, 16'd31455, 16'd22357, 16'd23318, 16'd21859, 16'd7046, 16'd62400, 16'd62194, 16'd8140, 16'd41332, 16'd12136, 16'd10801, 16'd46866, 16'd12813, 16'd52748, 16'd23108, 16'd21338, 16'd32511, 16'd59169, 16'd52275, 16'd16506, 16'd2423, 16'd28421, 16'd34022, 16'd40662});
	test_expansion(128'h14eed167d2a10dc234b51db6f323299e, {16'd18800, 16'd46816, 16'd23367, 16'd33063, 16'd61949, 16'd37300, 16'd57151, 16'd25106, 16'd33317, 16'd11532, 16'd36179, 16'd38583, 16'd34394, 16'd3774, 16'd13868, 16'd14825, 16'd48267, 16'd53997, 16'd12846, 16'd33614, 16'd4104, 16'd36722, 16'd46876, 16'd55296, 16'd21002, 16'd33039});
	test_expansion(128'hb4b87bc14c43a98db96a469b0ca86509, {16'd62417, 16'd22569, 16'd35005, 16'd14171, 16'd25243, 16'd31619, 16'd60746, 16'd38747, 16'd16508, 16'd30278, 16'd62561, 16'd49448, 16'd57696, 16'd42375, 16'd3464, 16'd23895, 16'd50620, 16'd41923, 16'd14726, 16'd5283, 16'd9417, 16'd33735, 16'd3364, 16'd46762, 16'd60302, 16'd11289});
	test_expansion(128'hc39bcdcc5dc81d703e15f9e53aa84bdf, {16'd4219, 16'd61955, 16'd3902, 16'd5509, 16'd44841, 16'd29799, 16'd5613, 16'd10430, 16'd3480, 16'd6647, 16'd2037, 16'd6829, 16'd2266, 16'd42371, 16'd45239, 16'd14480, 16'd1891, 16'd17793, 16'd42508, 16'd559, 16'd42592, 16'd23078, 16'd44458, 16'd21903, 16'd35241, 16'd39209});
	test_expansion(128'h12c1f387fb21a6f0de46236e48743fc2, {16'd38772, 16'd27615, 16'd27666, 16'd25389, 16'd10662, 16'd31814, 16'd6895, 16'd4234, 16'd2127, 16'd43013, 16'd55360, 16'd65210, 16'd58940, 16'd21825, 16'd44760, 16'd61323, 16'd12559, 16'd44637, 16'd19347, 16'd46669, 16'd7654, 16'd31795, 16'd6052, 16'd36273, 16'd38352, 16'd53738});
	test_expansion(128'h95511186e44a79cf41b96f34a9342d94, {16'd9904, 16'd22663, 16'd14228, 16'd64333, 16'd7134, 16'd23688, 16'd5370, 16'd48179, 16'd32841, 16'd24382, 16'd38835, 16'd21918, 16'd11746, 16'd55102, 16'd40520, 16'd17171, 16'd65138, 16'd38868, 16'd31597, 16'd53669, 16'd18518, 16'd63185, 16'd63720, 16'd30393, 16'd44793, 16'd54412});
	test_expansion(128'h3c115110e1558b828756d967fae0e6c9, {16'd37413, 16'd46065, 16'd55738, 16'd51388, 16'd29982, 16'd45240, 16'd57779, 16'd65142, 16'd37804, 16'd30725, 16'd63047, 16'd35044, 16'd59278, 16'd60996, 16'd48503, 16'd7794, 16'd39510, 16'd25774, 16'd52351, 16'd51105, 16'd29050, 16'd63362, 16'd25888, 16'd1365, 16'd36765, 16'd6549});
	test_expansion(128'h3f651f3179a3489011f3fd1d734adf4e, {16'd30339, 16'd24988, 16'd34213, 16'd38815, 16'd50793, 16'd42527, 16'd65225, 16'd32065, 16'd11872, 16'd64134, 16'd55335, 16'd39683, 16'd28529, 16'd11759, 16'd60049, 16'd45046, 16'd24100, 16'd1335, 16'd59730, 16'd62818, 16'd30854, 16'd30976, 16'd8718, 16'd48767, 16'd41051, 16'd43184});
	test_expansion(128'he00c058abd1e011dabb516aeeb9a74d2, {16'd55130, 16'd25667, 16'd16901, 16'd15324, 16'd33298, 16'd34048, 16'd31007, 16'd2190, 16'd53066, 16'd64186, 16'd38019, 16'd2226, 16'd2543, 16'd26965, 16'd48510, 16'd45177, 16'd38568, 16'd28014, 16'd31053, 16'd42723, 16'd19394, 16'd63259, 16'd49660, 16'd19413, 16'd32528, 16'd38712});
	test_expansion(128'h5198c32143e4eac80f5b65a8167e926c, {16'd31897, 16'd17179, 16'd3337, 16'd41991, 16'd28895, 16'd12313, 16'd47703, 16'd25104, 16'd36394, 16'd25708, 16'd22926, 16'd12064, 16'd38454, 16'd39208, 16'd34881, 16'd59116, 16'd64362, 16'd446, 16'd4919, 16'd47178, 16'd18644, 16'd23093, 16'd38948, 16'd8763, 16'd21831, 16'd2545});
	test_expansion(128'h1e6f5b5005d044ab568568dd32640141, {16'd11945, 16'd4558, 16'd14833, 16'd17078, 16'd45784, 16'd36777, 16'd358, 16'd53239, 16'd63519, 16'd61273, 16'd24621, 16'd52263, 16'd17807, 16'd48906, 16'd21983, 16'd38204, 16'd17916, 16'd54055, 16'd39890, 16'd18275, 16'd17021, 16'd11430, 16'd28399, 16'd17700, 16'd14757, 16'd56624});
	test_expansion(128'h13b03b894e9f599a14e3fde36b323ff5, {16'd51018, 16'd17197, 16'd37900, 16'd26084, 16'd58128, 16'd35292, 16'd11677, 16'd20625, 16'd1398, 16'd36508, 16'd43246, 16'd8816, 16'd9362, 16'd16483, 16'd12868, 16'd19037, 16'd56796, 16'd789, 16'd33262, 16'd49396, 16'd24147, 16'd22628, 16'd31099, 16'd20836, 16'd64991, 16'd20100});
	test_expansion(128'h8e7ab181de2f2c653170051aeac35189, {16'd34855, 16'd31870, 16'd44939, 16'd26664, 16'd40931, 16'd34263, 16'd47363, 16'd42078, 16'd12080, 16'd13017, 16'd28256, 16'd36983, 16'd23907, 16'd43994, 16'd49694, 16'd29051, 16'd1348, 16'd43965, 16'd53117, 16'd33577, 16'd37417, 16'd34283, 16'd17191, 16'd48018, 16'd8720, 16'd41458});
	test_expansion(128'hcab456693f8eec075d5984423776a104, {16'd8723, 16'd13468, 16'd22728, 16'd13076, 16'd12676, 16'd36548, 16'd11546, 16'd47352, 16'd26103, 16'd19069, 16'd3521, 16'd26468, 16'd22255, 16'd17397, 16'd6293, 16'd55108, 16'd24704, 16'd41605, 16'd39618, 16'd2787, 16'd35219, 16'd3862, 16'd51722, 16'd26767, 16'd11757, 16'd4683});
	test_expansion(128'hba15651a98c712871a21c421a66a5360, {16'd34856, 16'd19384, 16'd16712, 16'd9922, 16'd2147, 16'd49889, 16'd50465, 16'd21439, 16'd55258, 16'd8547, 16'd43321, 16'd4146, 16'd15646, 16'd27756, 16'd20642, 16'd46221, 16'd15367, 16'd57436, 16'd14158, 16'd7231, 16'd20262, 16'd35394, 16'd34047, 16'd56088, 16'd50577, 16'd22807});
	test_expansion(128'h312c297626237355528782694fc6d3ac, {16'd22860, 16'd51120, 16'd12663, 16'd21642, 16'd20028, 16'd63260, 16'd53196, 16'd51027, 16'd5641, 16'd40872, 16'd53229, 16'd53461, 16'd58746, 16'd6941, 16'd61460, 16'd51262, 16'd37583, 16'd24224, 16'd36968, 16'd37493, 16'd39473, 16'd3989, 16'd56583, 16'd22888, 16'd24362, 16'd40730});
	test_expansion(128'h80c32052fe5b7eefe774e5afadc80381, {16'd54054, 16'd3871, 16'd25571, 16'd4913, 16'd57031, 16'd17864, 16'd64858, 16'd54574, 16'd23617, 16'd18936, 16'd53969, 16'd60463, 16'd6865, 16'd26318, 16'd2944, 16'd60452, 16'd16713, 16'd53258, 16'd1927, 16'd28987, 16'd21592, 16'd18396, 16'd44883, 16'd25047, 16'd24959, 16'd48326});
	test_expansion(128'he7546ed4c1a329805aa01969283641cf, {16'd25247, 16'd45930, 16'd29959, 16'd28016, 16'd15947, 16'd21190, 16'd6418, 16'd43804, 16'd61273, 16'd65290, 16'd18974, 16'd7878, 16'd26848, 16'd28849, 16'd30101, 16'd13170, 16'd51033, 16'd12519, 16'd39324, 16'd47399, 16'd27382, 16'd18405, 16'd44097, 16'd44230, 16'd27207, 16'd24899});
	test_expansion(128'h091b549122d4c808cd6714d06c9afe68, {16'd29457, 16'd2587, 16'd59407, 16'd19204, 16'd48468, 16'd3265, 16'd3673, 16'd60625, 16'd14193, 16'd60489, 16'd23567, 16'd573, 16'd47831, 16'd12604, 16'd195, 16'd15048, 16'd48300, 16'd58966, 16'd18697, 16'd7023, 16'd27955, 16'd59973, 16'd27328, 16'd51248, 16'd754, 16'd6770});
	test_expansion(128'h3cbc95a68f48a0f7ac3f709201d898b8, {16'd55912, 16'd50802, 16'd39804, 16'd57459, 16'd31920, 16'd7485, 16'd37874, 16'd3395, 16'd35878, 16'd14846, 16'd23707, 16'd58478, 16'd53518, 16'd47481, 16'd49830, 16'd5382, 16'd61322, 16'd12498, 16'd9389, 16'd1038, 16'd29839, 16'd27844, 16'd42488, 16'd9057, 16'd2940, 16'd399});
	test_expansion(128'haaa3d70a977ab5762ce19b8a4bb890a6, {16'd50066, 16'd44961, 16'd38941, 16'd15450, 16'd14478, 16'd14444, 16'd13173, 16'd50607, 16'd25290, 16'd49553, 16'd18901, 16'd385, 16'd7497, 16'd45069, 16'd51990, 16'd5695, 16'd33978, 16'd13402, 16'd56368, 16'd39771, 16'd15871, 16'd51258, 16'd16503, 16'd36285, 16'd51918, 16'd40993});
	test_expansion(128'hcb07d666a63dc373c29cf8ce0a3f3617, {16'd30564, 16'd8812, 16'd3988, 16'd32678, 16'd43693, 16'd24420, 16'd29884, 16'd9230, 16'd22299, 16'd30284, 16'd54542, 16'd36330, 16'd28246, 16'd26930, 16'd62704, 16'd4387, 16'd4323, 16'd63278, 16'd22390, 16'd60612, 16'd14964, 16'd62186, 16'd51556, 16'd33900, 16'd19052, 16'd22024});
	test_expansion(128'hec827b09c80d021374d45ff000684287, {16'd37785, 16'd15281, 16'd45380, 16'd7659, 16'd3782, 16'd6715, 16'd49752, 16'd3009, 16'd47906, 16'd40041, 16'd4271, 16'd16604, 16'd28186, 16'd45151, 16'd53030, 16'd41875, 16'd39256, 16'd31154, 16'd64868, 16'd9189, 16'd12289, 16'd54688, 16'd8006, 16'd11377, 16'd59949, 16'd17894});
	test_expansion(128'h114c5148aada900e52882655a2211de2, {16'd3635, 16'd3163, 16'd10531, 16'd25605, 16'd57837, 16'd17612, 16'd14820, 16'd1583, 16'd8063, 16'd2614, 16'd59092, 16'd16237, 16'd17976, 16'd18186, 16'd28668, 16'd8335, 16'd64206, 16'd64459, 16'd174, 16'd32565, 16'd28643, 16'd8585, 16'd5525, 16'd26979, 16'd62889, 16'd14609});
	test_expansion(128'h1fe534575d360799a661d124392e2f8e, {16'd21933, 16'd54382, 16'd39634, 16'd65201, 16'd6436, 16'd13902, 16'd8037, 16'd24612, 16'd52384, 16'd30903, 16'd2778, 16'd42055, 16'd48818, 16'd17419, 16'd61853, 16'd15705, 16'd59553, 16'd49425, 16'd63056, 16'd58519, 16'd63435, 16'd61857, 16'd40921, 16'd19824, 16'd60398, 16'd33474});
	test_expansion(128'h4eefac193b1a250125196f9dd63b2e8c, {16'd59182, 16'd46401, 16'd6863, 16'd19008, 16'd53874, 16'd23129, 16'd53200, 16'd25098, 16'd60495, 16'd31397, 16'd34841, 16'd56378, 16'd14400, 16'd43422, 16'd12127, 16'd62210, 16'd53176, 16'd7354, 16'd46708, 16'd36966, 16'd7418, 16'd24984, 16'd37885, 16'd37083, 16'd52589, 16'd58015});
	test_expansion(128'h5a9346c14771834c166eff8df33efecc, {16'd57423, 16'd20063, 16'd45313, 16'd25070, 16'd62792, 16'd57426, 16'd61415, 16'd34231, 16'd24747, 16'd17038, 16'd11985, 16'd7237, 16'd41343, 16'd7757, 16'd59129, 16'd56076, 16'd46834, 16'd49981, 16'd21878, 16'd22949, 16'd5489, 16'd22545, 16'd5257, 16'd19018, 16'd51377, 16'd16552});
	test_expansion(128'h8074365ef6b976e17e2400b58d593df5, {16'd64970, 16'd62116, 16'd52021, 16'd9269, 16'd49562, 16'd59368, 16'd62797, 16'd5539, 16'd63511, 16'd22020, 16'd14915, 16'd60709, 16'd10240, 16'd20927, 16'd49681, 16'd25366, 16'd21440, 16'd48461, 16'd38856, 16'd5697, 16'd64452, 16'd13479, 16'd39197, 16'd25613, 16'd15208, 16'd38170});
	test_expansion(128'h311d6b398a211d773834022bde91e6ee, {16'd20555, 16'd30635, 16'd64819, 16'd35339, 16'd25729, 16'd17480, 16'd30848, 16'd38427, 16'd19017, 16'd16817, 16'd24439, 16'd5552, 16'd44505, 16'd43726, 16'd18330, 16'd37654, 16'd44145, 16'd60881, 16'd21513, 16'd17596, 16'd40621, 16'd38232, 16'd58677, 16'd49298, 16'd20637, 16'd55098});
	test_expansion(128'ha01bd22ff2aa733f06f1ae6993c2bf04, {16'd59244, 16'd54775, 16'd57271, 16'd40665, 16'd45284, 16'd28100, 16'd20019, 16'd28931, 16'd4845, 16'd42860, 16'd60893, 16'd22326, 16'd52334, 16'd61173, 16'd40972, 16'd61627, 16'd51570, 16'd51752, 16'd47537, 16'd23531, 16'd52514, 16'd15724, 16'd11661, 16'd18795, 16'd20322, 16'd41732});
	test_expansion(128'h1b0225d080342460d10055db6b86785f, {16'd14642, 16'd6106, 16'd63831, 16'd39988, 16'd24987, 16'd49223, 16'd42653, 16'd55400, 16'd44669, 16'd53133, 16'd54651, 16'd40791, 16'd19767, 16'd9918, 16'd58971, 16'd48035, 16'd34227, 16'd51485, 16'd65185, 16'd58236, 16'd13152, 16'd33311, 16'd33699, 16'd57929, 16'd345, 16'd7663});
	test_expansion(128'hddcc29e0d9a2f0a65866abbeee81af42, {16'd6517, 16'd64873, 16'd38030, 16'd11560, 16'd53907, 16'd54682, 16'd16500, 16'd55007, 16'd21601, 16'd24552, 16'd61938, 16'd10951, 16'd9508, 16'd6429, 16'd33548, 16'd1402, 16'd27543, 16'd15777, 16'd60722, 16'd34258, 16'd2555, 16'd43230, 16'd22621, 16'd51273, 16'd44993, 16'd5342});
	test_expansion(128'h74002d55597cb904c347c2d7d0e2a965, {16'd64504, 16'd55148, 16'd59343, 16'd23499, 16'd46720, 16'd16756, 16'd29261, 16'd16114, 16'd9549, 16'd8886, 16'd27319, 16'd5742, 16'd40078, 16'd49102, 16'd1639, 16'd45205, 16'd23065, 16'd47872, 16'd3054, 16'd35537, 16'd14735, 16'd8746, 16'd10902, 16'd21264, 16'd14352, 16'd63427});
	test_expansion(128'h3031e3b7b1d17bfd0c998ff693b9f167, {16'd16786, 16'd25321, 16'd29964, 16'd16063, 16'd14156, 16'd28642, 16'd28538, 16'd49821, 16'd54105, 16'd31806, 16'd25861, 16'd50638, 16'd9966, 16'd57603, 16'd3290, 16'd44140, 16'd60451, 16'd23016, 16'd41791, 16'd46735, 16'd49082, 16'd23309, 16'd57512, 16'd45592, 16'd30338, 16'd50909});
	test_expansion(128'ha6d1a13832bb706b832563703e0cd8c4, {16'd26960, 16'd7922, 16'd31186, 16'd34721, 16'd4887, 16'd38724, 16'd41957, 16'd48273, 16'd31730, 16'd37234, 16'd28151, 16'd15162, 16'd42909, 16'd58541, 16'd9312, 16'd7021, 16'd6439, 16'd34404, 16'd2670, 16'd43331, 16'd44314, 16'd56966, 16'd3982, 16'd956, 16'd37219, 16'd53776});
	test_expansion(128'hce6f1ba932deab74786daabf9a45b636, {16'd6375, 16'd62499, 16'd39745, 16'd16617, 16'd49626, 16'd63718, 16'd53731, 16'd37113, 16'd46014, 16'd7182, 16'd8243, 16'd57603, 16'd23964, 16'd34863, 16'd4597, 16'd37453, 16'd12674, 16'd26811, 16'd9272, 16'd16945, 16'd27272, 16'd37913, 16'd27287, 16'd33388, 16'd23152, 16'd47711});
	test_expansion(128'ha7e0368fec774a8279587e0799b975a4, {16'd56496, 16'd43479, 16'd21015, 16'd64080, 16'd6220, 16'd65020, 16'd62407, 16'd64570, 16'd61126, 16'd15066, 16'd32367, 16'd60002, 16'd60992, 16'd4208, 16'd7763, 16'd13332, 16'd16779, 16'd33866, 16'd42369, 16'd60835, 16'd19729, 16'd41587, 16'd13209, 16'd57470, 16'd7848, 16'd60265});
	test_expansion(128'hb705f8518c2c4a720053302ef45375a0, {16'd17148, 16'd21560, 16'd23727, 16'd14021, 16'd16131, 16'd29209, 16'd3968, 16'd30532, 16'd11353, 16'd42446, 16'd24571, 16'd27633, 16'd25148, 16'd36918, 16'd22800, 16'd19576, 16'd48802, 16'd60193, 16'd31608, 16'd29717, 16'd61923, 16'd62576, 16'd5366, 16'd22493, 16'd25852, 16'd63759});
	test_expansion(128'h9bb29998784f40f9513ff74035b88245, {16'd60325, 16'd58702, 16'd3655, 16'd10465, 16'd12179, 16'd44426, 16'd24487, 16'd64170, 16'd40891, 16'd15542, 16'd49691, 16'd53474, 16'd51459, 16'd15609, 16'd56375, 16'd8748, 16'd22832, 16'd17753, 16'd37972, 16'd43163, 16'd58876, 16'd22144, 16'd13956, 16'd17561, 16'd22612, 16'd47082});
	test_expansion(128'h6522c44db083475396a8f88e6e7921f1, {16'd9163, 16'd61905, 16'd58949, 16'd39105, 16'd57126, 16'd65241, 16'd20785, 16'd44170, 16'd39148, 16'd1549, 16'd28994, 16'd62435, 16'd17273, 16'd13237, 16'd54114, 16'd59387, 16'd54895, 16'd12671, 16'd58879, 16'd15239, 16'd4211, 16'd13173, 16'd56499, 16'd34858, 16'd6419, 16'd64634});
	test_expansion(128'h5a2695ab9c2d30a09efdba71d7bc7704, {16'd27190, 16'd33310, 16'd25405, 16'd55633, 16'd62188, 16'd38495, 16'd46944, 16'd27817, 16'd3873, 16'd5494, 16'd28041, 16'd37652, 16'd44148, 16'd28117, 16'd37631, 16'd11288, 16'd13098, 16'd34401, 16'd36044, 16'd50338, 16'd63192, 16'd55174, 16'd12525, 16'd14699, 16'd12131, 16'd49160});
	test_expansion(128'h69cfc1cc4fb1d186025813853d8a1eb5, {16'd32642, 16'd605, 16'd5439, 16'd16171, 16'd63981, 16'd16859, 16'd42816, 16'd39349, 16'd2062, 16'd18949, 16'd34760, 16'd63840, 16'd45418, 16'd58043, 16'd2628, 16'd16040, 16'd37921, 16'd43783, 16'd54594, 16'd8722, 16'd26178, 16'd59942, 16'd54478, 16'd20801, 16'd34702, 16'd19158});
	test_expansion(128'hfe0e3e7eff047cdc40ff61ff2b7e8909, {16'd27980, 16'd45065, 16'd41694, 16'd32872, 16'd44400, 16'd39139, 16'd50408, 16'd29348, 16'd60965, 16'd63461, 16'd22293, 16'd28405, 16'd61836, 16'd36664, 16'd10159, 16'd53746, 16'd15356, 16'd42508, 16'd5540, 16'd9485, 16'd30898, 16'd34582, 16'd56679, 16'd23352, 16'd11122, 16'd39472});
	test_expansion(128'h3ae4b52defc18384799e1e54d2a45c3a, {16'd60004, 16'd63078, 16'd54694, 16'd5430, 16'd23793, 16'd55032, 16'd5194, 16'd13175, 16'd33226, 16'd39029, 16'd56992, 16'd5099, 16'd46604, 16'd8125, 16'd63530, 16'd20464, 16'd39100, 16'd26498, 16'd38677, 16'd60670, 16'd37155, 16'd49631, 16'd37690, 16'd40948, 16'd20069, 16'd50916});
	test_expansion(128'ha56c876ccf2d5c13ecd7dccaaebaf460, {16'd1511, 16'd34087, 16'd16884, 16'd41507, 16'd2884, 16'd37434, 16'd45470, 16'd34728, 16'd50935, 16'd59067, 16'd34908, 16'd27317, 16'd42169, 16'd62381, 16'd33892, 16'd55939, 16'd31309, 16'd41950, 16'd10651, 16'd57424, 16'd42427, 16'd27014, 16'd22165, 16'd11000, 16'd15990, 16'd24516});
	test_expansion(128'h1b559bf131566b250643fb77620c92fc, {16'd52775, 16'd42875, 16'd44775, 16'd31221, 16'd36121, 16'd21395, 16'd45323, 16'd15007, 16'd6971, 16'd61237, 16'd50147, 16'd25461, 16'd57866, 16'd5245, 16'd33299, 16'd19431, 16'd30690, 16'd61238, 16'd59002, 16'd38065, 16'd41584, 16'd38137, 16'd28718, 16'd32347, 16'd28211, 16'd8903});
	test_expansion(128'hc35bf657d5b1a829b223e7ba2ef77b66, {16'd2853, 16'd50306, 16'd38820, 16'd13298, 16'd35326, 16'd2760, 16'd15762, 16'd33316, 16'd26963, 16'd7827, 16'd33636, 16'd56968, 16'd31194, 16'd5549, 16'd11959, 16'd5623, 16'd47954, 16'd51379, 16'd56301, 16'd16294, 16'd55529, 16'd11457, 16'd22908, 16'd23707, 16'd31462, 16'd22122});
	test_expansion(128'h5812ceb326b4ab6a7f6b6711b48ca123, {16'd13546, 16'd63579, 16'd54813, 16'd49432, 16'd22969, 16'd22742, 16'd53690, 16'd34435, 16'd29108, 16'd27230, 16'd9070, 16'd31002, 16'd4583, 16'd3383, 16'd26645, 16'd7270, 16'd62230, 16'd19218, 16'd10648, 16'd28987, 16'd47320, 16'd46114, 16'd41589, 16'd11386, 16'd2975, 16'd13257});
	test_expansion(128'hbe50fcadb32606fa5b8099820f28c894, {16'd37428, 16'd30433, 16'd42279, 16'd40692, 16'd32895, 16'd7994, 16'd56017, 16'd44886, 16'd56366, 16'd16600, 16'd40795, 16'd44087, 16'd60773, 16'd42368, 16'd24424, 16'd32679, 16'd43042, 16'd2180, 16'd646, 16'd30486, 16'd3716, 16'd44558, 16'd38655, 16'd62586, 16'd23393, 16'd31532});
	test_expansion(128'hd95c2bd78c0014e65fd1b2bee7766f42, {16'd58934, 16'd5483, 16'd4109, 16'd63608, 16'd28340, 16'd18745, 16'd21326, 16'd28619, 16'd10625, 16'd23003, 16'd60164, 16'd15895, 16'd60508, 16'd5089, 16'd48138, 16'd38468, 16'd11050, 16'd46424, 16'd228, 16'd42466, 16'd44797, 16'd1452, 16'd13612, 16'd38019, 16'd33208, 16'd52528});
	test_expansion(128'hf0028630995979c7832200bd9711098d, {16'd14445, 16'd42865, 16'd14469, 16'd60320, 16'd57905, 16'd42788, 16'd38637, 16'd61289, 16'd18793, 16'd62529, 16'd22055, 16'd60542, 16'd11498, 16'd33168, 16'd13544, 16'd29248, 16'd39149, 16'd3697, 16'd46039, 16'd22878, 16'd9291, 16'd20186, 16'd37093, 16'd7170, 16'd64254, 16'd50887});
	test_expansion(128'h63c636f717729f67e8bf1105e878f5bd, {16'd11236, 16'd30793, 16'd2164, 16'd65317, 16'd6472, 16'd45526, 16'd12155, 16'd46755, 16'd44068, 16'd39753, 16'd41335, 16'd23553, 16'd2015, 16'd40614, 16'd19440, 16'd53878, 16'd12651, 16'd38878, 16'd55244, 16'd60778, 16'd12077, 16'd1883, 16'd22805, 16'd20700, 16'd46333, 16'd3633});
	test_expansion(128'he48acb3d63b214358c469b3abaca6c46, {16'd23777, 16'd18289, 16'd3705, 16'd38605, 16'd51768, 16'd64247, 16'd1748, 16'd40444, 16'd52324, 16'd22126, 16'd34572, 16'd43219, 16'd60289, 16'd24391, 16'd40697, 16'd31681, 16'd32341, 16'd20267, 16'd57536, 16'd29787, 16'd34882, 16'd44364, 16'd9669, 16'd27716, 16'd52401, 16'd64763});
	test_expansion(128'h993e026c745cd685de1644b71738e4d6, {16'd24426, 16'd65411, 16'd25474, 16'd6012, 16'd29739, 16'd2189, 16'd57225, 16'd63348, 16'd48091, 16'd2996, 16'd16808, 16'd10340, 16'd60017, 16'd5621, 16'd54285, 16'd2434, 16'd32315, 16'd48127, 16'd4502, 16'd14470, 16'd38646, 16'd30210, 16'd11929, 16'd59863, 16'd3392, 16'd4974});
	test_expansion(128'h8ba65f490d063a8ae0fc2a68fc481bc8, {16'd31423, 16'd34223, 16'd10229, 16'd33655, 16'd22889, 16'd48482, 16'd44717, 16'd62369, 16'd14501, 16'd28920, 16'd62973, 16'd51206, 16'd14246, 16'd65308, 16'd41185, 16'd11962, 16'd3313, 16'd12852, 16'd63160, 16'd11323, 16'd61598, 16'd12061, 16'd41131, 16'd9803, 16'd22422, 16'd63876});
	test_expansion(128'h5a6e20ee1ef5aac8e641cf1a90887822, {16'd49212, 16'd16704, 16'd21713, 16'd21955, 16'd36272, 16'd39108, 16'd2525, 16'd34154, 16'd45559, 16'd52252, 16'd32803, 16'd38095, 16'd18525, 16'd6185, 16'd18785, 16'd25475, 16'd23973, 16'd51188, 16'd42406, 16'd2919, 16'd8081, 16'd18525, 16'd59983, 16'd59894, 16'd17999, 16'd21584});
	test_expansion(128'h6236544ebd7874b77cbcd55150320ca1, {16'd6192, 16'd1812, 16'd16901, 16'd36299, 16'd3541, 16'd20046, 16'd34509, 16'd59714, 16'd50049, 16'd29567, 16'd36656, 16'd39981, 16'd51128, 16'd44249, 16'd50447, 16'd45282, 16'd22207, 16'd64189, 16'd820, 16'd15844, 16'd59755, 16'd7238, 16'd55361, 16'd55757, 16'd63227, 16'd28908});
	test_expansion(128'he921b2c4c80d948520a63684b30a8498, {16'd56013, 16'd56182, 16'd58789, 16'd13671, 16'd9390, 16'd5117, 16'd52789, 16'd1901, 16'd42227, 16'd41000, 16'd4902, 16'd16159, 16'd21316, 16'd48962, 16'd9838, 16'd36489, 16'd22111, 16'd35546, 16'd50056, 16'd4058, 16'd17772, 16'd64013, 16'd432, 16'd23446, 16'd13533, 16'd3437});
	test_expansion(128'hd2559dd8281bd4496b14af6319f19446, {16'd57430, 16'd1561, 16'd19938, 16'd21857, 16'd19930, 16'd63011, 16'd46087, 16'd30526, 16'd44638, 16'd35525, 16'd64243, 16'd37430, 16'd58994, 16'd24380, 16'd8218, 16'd19152, 16'd29949, 16'd60208, 16'd59448, 16'd22440, 16'd24596, 16'd54504, 16'd59528, 16'd37205, 16'd35715, 16'd21670});
	test_expansion(128'h33f284c64a781c33495900f3a659b83f, {16'd45906, 16'd54378, 16'd33751, 16'd39936, 16'd49663, 16'd27801, 16'd13044, 16'd24663, 16'd40443, 16'd19420, 16'd45697, 16'd22958, 16'd60038, 16'd54077, 16'd8, 16'd9202, 16'd35596, 16'd28241, 16'd58023, 16'd20170, 16'd48185, 16'd4829, 16'd12628, 16'd23888, 16'd45565, 16'd5352});
	test_expansion(128'h73082f5e696d92593b6361eea2cb650e, {16'd30976, 16'd22952, 16'd40748, 16'd23093, 16'd60630, 16'd59551, 16'd1662, 16'd2561, 16'd5421, 16'd35323, 16'd64105, 16'd15190, 16'd27866, 16'd52372, 16'd56934, 16'd35728, 16'd39249, 16'd974, 16'd26473, 16'd20504, 16'd7942, 16'd21778, 16'd59935, 16'd61126, 16'd51870, 16'd19579});
	test_expansion(128'hf002fb01ccf8b97d724898d706c3857e, {16'd17906, 16'd48891, 16'd55661, 16'd58464, 16'd53752, 16'd4381, 16'd57795, 16'd7056, 16'd61635, 16'd47555, 16'd20640, 16'd34378, 16'd40564, 16'd42676, 16'd18184, 16'd38103, 16'd14035, 16'd28980, 16'd25291, 16'd17169, 16'd17119, 16'd39101, 16'd13421, 16'd5116, 16'd13528, 16'd6898});
	test_expansion(128'h419a6adaf0c42725908f45e6f7aa9378, {16'd23615, 16'd40865, 16'd35326, 16'd17890, 16'd64812, 16'd6490, 16'd59131, 16'd5715, 16'd39468, 16'd28758, 16'd59602, 16'd38958, 16'd64447, 16'd59168, 16'd29458, 16'd16865, 16'd19998, 16'd59821, 16'd21366, 16'd47271, 16'd53906, 16'd46220, 16'd47850, 16'd48138, 16'd32755, 16'd45287});
	test_expansion(128'h186e253276500f06c042befa0c54417a, {16'd32710, 16'd38320, 16'd14242, 16'd36726, 16'd14310, 16'd65191, 16'd8950, 16'd47651, 16'd13762, 16'd11697, 16'd39529, 16'd52306, 16'd63012, 16'd43351, 16'd62586, 16'd18974, 16'd63596, 16'd24654, 16'd2059, 16'd9314, 16'd10506, 16'd13695, 16'd51722, 16'd64358, 16'd50152, 16'd17688});
	test_expansion(128'h1bc0d1111943544e9b16c232e93169b9, {16'd58418, 16'd8751, 16'd61517, 16'd61172, 16'd48995, 16'd18715, 16'd14329, 16'd27283, 16'd50116, 16'd11262, 16'd26409, 16'd44052, 16'd55618, 16'd18063, 16'd6603, 16'd4510, 16'd35367, 16'd24850, 16'd38209, 16'd57957, 16'd4531, 16'd7378, 16'd31339, 16'd49410, 16'd8338, 16'd47182});
	test_expansion(128'h2120fd6f57eb9d70f8fc6836b4f128d3, {16'd36338, 16'd2735, 16'd3451, 16'd45766, 16'd16762, 16'd19438, 16'd11248, 16'd7390, 16'd25136, 16'd3416, 16'd5058, 16'd36884, 16'd37051, 16'd38390, 16'd51435, 16'd64849, 16'd51680, 16'd6269, 16'd50772, 16'd53891, 16'd9619, 16'd14177, 16'd57005, 16'd36489, 16'd14494, 16'd18776});
	test_expansion(128'hea6f1d1a52319ef5976b136bcb8e134b, {16'd17754, 16'd37490, 16'd41745, 16'd34962, 16'd8866, 16'd65103, 16'd43984, 16'd54470, 16'd24853, 16'd11463, 16'd21907, 16'd18926, 16'd11194, 16'd60572, 16'd43418, 16'd1154, 16'd9949, 16'd54268, 16'd52428, 16'd30124, 16'd43170, 16'd57360, 16'd32010, 16'd31360, 16'd26674, 16'd35573});
	test_expansion(128'h9f065ee34240df318d13538356165168, {16'd31193, 16'd56974, 16'd47326, 16'd927, 16'd34987, 16'd16261, 16'd35181, 16'd38718, 16'd50772, 16'd63212, 16'd61075, 16'd38525, 16'd34372, 16'd26136, 16'd53978, 16'd37277, 16'd13780, 16'd4779, 16'd42111, 16'd52646, 16'd63252, 16'd11842, 16'd47707, 16'd17505, 16'd62114, 16'd59114});
	test_expansion(128'hd63ef3a3e99058849ff184a81edb8180, {16'd27113, 16'd40696, 16'd32897, 16'd59617, 16'd17536, 16'd62130, 16'd12387, 16'd1491, 16'd14290, 16'd8689, 16'd32376, 16'd55850, 16'd44050, 16'd38465, 16'd40175, 16'd57968, 16'd11359, 16'd4907, 16'd51396, 16'd11824, 16'd14737, 16'd22366, 16'd50845, 16'd42726, 16'd48236, 16'd6180});
	test_expansion(128'h35fca98ded6e7180d785a0fb147df9c8, {16'd5617, 16'd53827, 16'd50320, 16'd16416, 16'd29889, 16'd42855, 16'd60981, 16'd44877, 16'd1544, 16'd36692, 16'd40192, 16'd1650, 16'd59945, 16'd5515, 16'd48243, 16'd55854, 16'd54883, 16'd18525, 16'd585, 16'd54238, 16'd29478, 16'd44663, 16'd37338, 16'd9021, 16'd13621, 16'd42548});
	test_expansion(128'hf8fab049560d54d3ccd20461375267f2, {16'd62106, 16'd46472, 16'd54336, 16'd54333, 16'd40896, 16'd22120, 16'd62553, 16'd41484, 16'd16085, 16'd43199, 16'd35138, 16'd13796, 16'd20130, 16'd3102, 16'd59958, 16'd20080, 16'd10086, 16'd19070, 16'd10670, 16'd24546, 16'd63254, 16'd61808, 16'd30875, 16'd19143, 16'd58753, 16'd24810});
	test_expansion(128'hc064d84f520c85b30b6458d0ba55a839, {16'd63837, 16'd9996, 16'd12355, 16'd49859, 16'd46913, 16'd7721, 16'd32442, 16'd8506, 16'd18792, 16'd35229, 16'd24075, 16'd62174, 16'd3109, 16'd41812, 16'd56052, 16'd4274, 16'd41733, 16'd4637, 16'd7919, 16'd32677, 16'd61922, 16'd48150, 16'd1024, 16'd29614, 16'd42348, 16'd60665});
	test_expansion(128'hf1117248457659d749ce186b6d4f75f7, {16'd1632, 16'd53934, 16'd38270, 16'd27726, 16'd50374, 16'd11297, 16'd40757, 16'd62606, 16'd20116, 16'd53543, 16'd64785, 16'd50874, 16'd633, 16'd8172, 16'd41705, 16'd43192, 16'd3098, 16'd52239, 16'd6343, 16'd7606, 16'd58072, 16'd13045, 16'd58006, 16'd30861, 16'd11436, 16'd39879});
	test_expansion(128'hbf3d6fb2e8c9fbd9b8bd3c8b6cd1c947, {16'd50157, 16'd55877, 16'd50964, 16'd54061, 16'd46257, 16'd1961, 16'd42984, 16'd5421, 16'd29429, 16'd60045, 16'd3898, 16'd17834, 16'd1196, 16'd57281, 16'd56576, 16'd37386, 16'd40587, 16'd28914, 16'd59228, 16'd61768, 16'd45768, 16'd17113, 16'd10166, 16'd52690, 16'd32796, 16'd51783});
	test_expansion(128'h2f04024d32bcbf1b81ecc014f1d4216f, {16'd20328, 16'd6411, 16'd61709, 16'd28310, 16'd11998, 16'd52665, 16'd9100, 16'd55048, 16'd40423, 16'd25621, 16'd51817, 16'd62127, 16'd43982, 16'd22072, 16'd2897, 16'd20746, 16'd61983, 16'd36690, 16'd23878, 16'd54619, 16'd27771, 16'd9069, 16'd54225, 16'd45011, 16'd57639, 16'd44456});
	test_expansion(128'h91ec696905007c843a31235805b2b5b5, {16'd47000, 16'd31178, 16'd24158, 16'd62716, 16'd49565, 16'd62567, 16'd62621, 16'd23615, 16'd35345, 16'd54060, 16'd19669, 16'd7163, 16'd13712, 16'd37669, 16'd9378, 16'd12418, 16'd2734, 16'd41524, 16'd56922, 16'd906, 16'd55918, 16'd21159, 16'd9777, 16'd24420, 16'd38478, 16'd3170});
	test_expansion(128'h88061459743a67301bb2401f5d6246d1, {16'd60450, 16'd46722, 16'd33258, 16'd303, 16'd4132, 16'd8726, 16'd9225, 16'd338, 16'd43110, 16'd44952, 16'd59310, 16'd50811, 16'd40568, 16'd33246, 16'd24922, 16'd26600, 16'd45439, 16'd42570, 16'd38872, 16'd39169, 16'd6166, 16'd60006, 16'd15441, 16'd26637, 16'd3100, 16'd9405});
	test_expansion(128'h48de015bc9ce6ab2a1b8ae296c93e8fd, {16'd29560, 16'd23130, 16'd2509, 16'd51764, 16'd57359, 16'd51560, 16'd19368, 16'd43215, 16'd4472, 16'd38246, 16'd59769, 16'd38903, 16'd54067, 16'd49591, 16'd13148, 16'd46672, 16'd47999, 16'd36291, 16'd27958, 16'd19769, 16'd12909, 16'd14356, 16'd41580, 16'd44094, 16'd9919, 16'd23358});
	test_expansion(128'h8d7f7a80f9662379455526104b933703, {16'd28838, 16'd36943, 16'd20541, 16'd3557, 16'd39750, 16'd42923, 16'd21385, 16'd23648, 16'd46282, 16'd34512, 16'd6951, 16'd256, 16'd59091, 16'd53453, 16'd11843, 16'd27250, 16'd60181, 16'd8577, 16'd12848, 16'd30846, 16'd12357, 16'd21627, 16'd7457, 16'd48774, 16'd46910, 16'd15359});
	test_expansion(128'h730dfa1935628e189ab2f52035e50d5e, {16'd49205, 16'd43970, 16'd61153, 16'd17626, 16'd60969, 16'd41813, 16'd39852, 16'd9846, 16'd33312, 16'd60472, 16'd721, 16'd35285, 16'd23576, 16'd32970, 16'd34016, 16'd10126, 16'd34602, 16'd39904, 16'd10031, 16'd42894, 16'd63303, 16'd64520, 16'd47231, 16'd50485, 16'd39658, 16'd16991});
	test_expansion(128'h19b98ddcf49073cf5945dfa0582f7488, {16'd60377, 16'd59229, 16'd12821, 16'd50309, 16'd22019, 16'd3324, 16'd56464, 16'd44704, 16'd64904, 16'd64161, 16'd15387, 16'd18567, 16'd56253, 16'd39938, 16'd15477, 16'd60348, 16'd59377, 16'd21306, 16'd25281, 16'd12072, 16'd56652, 16'd45701, 16'd22811, 16'd30974, 16'd40881, 16'd44876});
	test_expansion(128'h71fbfef54b850e6085107755d2228311, {16'd51842, 16'd60459, 16'd7022, 16'd53611, 16'd26768, 16'd26512, 16'd64287, 16'd40040, 16'd46229, 16'd38514, 16'd22644, 16'd43063, 16'd9245, 16'd52225, 16'd20291, 16'd34915, 16'd51263, 16'd41319, 16'd50029, 16'd46771, 16'd29470, 16'd3743, 16'd6928, 16'd41899, 16'd47572, 16'd9042});
	test_expansion(128'hb3025406727f2fa8614999f1f9579683, {16'd60438, 16'd42175, 16'd34505, 16'd26685, 16'd27032, 16'd31912, 16'd12945, 16'd63456, 16'd38728, 16'd47361, 16'd53609, 16'd50936, 16'd35366, 16'd1436, 16'd41599, 16'd21533, 16'd23366, 16'd46821, 16'd9743, 16'd10686, 16'd39662, 16'd38418, 16'd23433, 16'd29208, 16'd14647, 16'd501});
	test_expansion(128'heca0cd2120d03612298c0f161dce658b, {16'd52110, 16'd40827, 16'd28911, 16'd59815, 16'd16578, 16'd5368, 16'd60649, 16'd36170, 16'd48519, 16'd49402, 16'd17211, 16'd16706, 16'd62645, 16'd34309, 16'd20220, 16'd47025, 16'd51746, 16'd30011, 16'd29948, 16'd61730, 16'd18273, 16'd2519, 16'd56063, 16'd12029, 16'd46106, 16'd49779});
	test_expansion(128'hd5ce58a9070b8e155c9bf1669485ebf5, {16'd56454, 16'd6530, 16'd34658, 16'd5855, 16'd46129, 16'd53995, 16'd49630, 16'd19574, 16'd39853, 16'd62934, 16'd31778, 16'd39885, 16'd10757, 16'd37565, 16'd4126, 16'd6754, 16'd64903, 16'd16340, 16'd36057, 16'd23629, 16'd44928, 16'd26009, 16'd41930, 16'd55269, 16'd57504, 16'd9908});
	test_expansion(128'h7cc2d65049f6430434cc66357932ddc9, {16'd35857, 16'd63128, 16'd12890, 16'd64205, 16'd29647, 16'd55445, 16'd32011, 16'd35122, 16'd33007, 16'd27023, 16'd20663, 16'd64863, 16'd46225, 16'd27173, 16'd39694, 16'd51794, 16'd28055, 16'd40160, 16'd31998, 16'd37896, 16'd29508, 16'd46191, 16'd30644, 16'd19782, 16'd45027, 16'd54966});
	test_expansion(128'h1716b433d7d7b774489455477714a738, {16'd3306, 16'd34400, 16'd41656, 16'd59486, 16'd56922, 16'd48252, 16'd12382, 16'd38910, 16'd53629, 16'd18739, 16'd19631, 16'd32534, 16'd23904, 16'd28290, 16'd55258, 16'd43623, 16'd9067, 16'd56543, 16'd11711, 16'd29858, 16'd44563, 16'd27932, 16'd23912, 16'd37658, 16'd63867, 16'd31171});
	test_expansion(128'h9d1e5d33eb7d6d45fd6415ae9e803686, {16'd9, 16'd16523, 16'd45679, 16'd28433, 16'd63461, 16'd22920, 16'd18304, 16'd34534, 16'd45629, 16'd64338, 16'd32667, 16'd62285, 16'd30246, 16'd26506, 16'd7298, 16'd37572, 16'd10622, 16'd39162, 16'd63992, 16'd3754, 16'd38563, 16'd56844, 16'd39602, 16'd28740, 16'd21978, 16'd56694});
	test_expansion(128'hdd1360bb58eb7f9b9d15c41b66eb43b4, {16'd35019, 16'd5277, 16'd45734, 16'd63446, 16'd56147, 16'd6508, 16'd57123, 16'd54627, 16'd24693, 16'd64929, 16'd40901, 16'd49754, 16'd15540, 16'd30861, 16'd18519, 16'd47303, 16'd17472, 16'd12393, 16'd24240, 16'd13818, 16'd24530, 16'd25955, 16'd50100, 16'd44218, 16'd2085, 16'd1022});
	test_expansion(128'haf41102f95ab5a84f0ed476931efdc8c, {16'd32026, 16'd35639, 16'd30592, 16'd63020, 16'd7641, 16'd65391, 16'd23332, 16'd58988, 16'd22965, 16'd13177, 16'd16295, 16'd10434, 16'd62950, 16'd43705, 16'd16445, 16'd24274, 16'd17879, 16'd59593, 16'd18650, 16'd12038, 16'd40495, 16'd30430, 16'd24137, 16'd64848, 16'd60772, 16'd13204});
	test_expansion(128'h0e423f649d7b3a5b15a9678b987d0520, {16'd53775, 16'd30487, 16'd48032, 16'd41548, 16'd11547, 16'd31009, 16'd37960, 16'd40134, 16'd7571, 16'd3583, 16'd43728, 16'd3129, 16'd17172, 16'd42201, 16'd18103, 16'd32126, 16'd24190, 16'd18826, 16'd8314, 16'd54423, 16'd47327, 16'd45183, 16'd10815, 16'd42345, 16'd53606, 16'd16309});
	test_expansion(128'h2a8ceb80b9e3690b638fd2e97d0ee798, {16'd23323, 16'd51964, 16'd54704, 16'd42373, 16'd8632, 16'd56817, 16'd31088, 16'd2158, 16'd56908, 16'd32141, 16'd24064, 16'd41552, 16'd3388, 16'd37588, 16'd10034, 16'd12841, 16'd52057, 16'd38729, 16'd23599, 16'd37698, 16'd7083, 16'd5391, 16'd36352, 16'd64975, 16'd18876, 16'd37414});
	test_expansion(128'h1ba77dfc0481b9ab7925f33c33a207c3, {16'd11810, 16'd7254, 16'd22782, 16'd45521, 16'd54799, 16'd30632, 16'd60467, 16'd52374, 16'd35593, 16'd64056, 16'd6818, 16'd24930, 16'd60889, 16'd41900, 16'd35555, 16'd19743, 16'd34152, 16'd5789, 16'd65258, 16'd31935, 16'd18765, 16'd60842, 16'd56390, 16'd32201, 16'd56619, 16'd54764});
	test_expansion(128'h047a5db0a4b26a3712e643cd6dce0f18, {16'd23547, 16'd32049, 16'd3976, 16'd57203, 16'd1484, 16'd40085, 16'd56684, 16'd9569, 16'd8875, 16'd37441, 16'd22677, 16'd60802, 16'd27317, 16'd20526, 16'd61642, 16'd59597, 16'd42531, 16'd50540, 16'd64097, 16'd16485, 16'd18109, 16'd43502, 16'd5938, 16'd32723, 16'd33916, 16'd43291});
	test_expansion(128'hde3e986b1ee5d8600031e8d9a55474ed, {16'd20153, 16'd62142, 16'd41115, 16'd32827, 16'd49247, 16'd64758, 16'd3992, 16'd60746, 16'd33107, 16'd51756, 16'd21316, 16'd19373, 16'd54115, 16'd17057, 16'd1707, 16'd51035, 16'd1265, 16'd7803, 16'd24231, 16'd15753, 16'd2219, 16'd39748, 16'd31438, 16'd41955, 16'd18117, 16'd13766});
	test_expansion(128'h7b1818323ceb6ec5e1a2c6893c59e31c, {16'd37592, 16'd45117, 16'd19590, 16'd22518, 16'd32306, 16'd17305, 16'd3812, 16'd19005, 16'd34320, 16'd22084, 16'd21504, 16'd22010, 16'd10829, 16'd9164, 16'd28374, 16'd4088, 16'd14917, 16'd31245, 16'd47478, 16'd37806, 16'd50735, 16'd28643, 16'd18183, 16'd46215, 16'd62327, 16'd35753});
	test_expansion(128'h839bd6cdb722f599c73e1a31918f81c6, {16'd33829, 16'd32552, 16'd57514, 16'd17268, 16'd53220, 16'd18691, 16'd36778, 16'd57458, 16'd40570, 16'd44062, 16'd16819, 16'd45482, 16'd62356, 16'd24517, 16'd45301, 16'd44336, 16'd13053, 16'd42996, 16'd57430, 16'd21943, 16'd53794, 16'd28479, 16'd45838, 16'd64251, 16'd54703, 16'd6878});
	test_expansion(128'h829c38d511f48e7b9c4323d9c79895cc, {16'd48283, 16'd15876, 16'd4212, 16'd12932, 16'd65493, 16'd22865, 16'd12502, 16'd49653, 16'd53779, 16'd6638, 16'd26450, 16'd51782, 16'd32092, 16'd15305, 16'd55973, 16'd56577, 16'd27858, 16'd42428, 16'd64960, 16'd42397, 16'd17391, 16'd52505, 16'd41880, 16'd17805, 16'd22810, 16'd54125});
	test_expansion(128'ha26ba101b10f192c9288579ae029b207, {16'd26863, 16'd23333, 16'd26425, 16'd1107, 16'd46769, 16'd44398, 16'd3966, 16'd64525, 16'd23781, 16'd29086, 16'd62698, 16'd35537, 16'd34217, 16'd45028, 16'd58357, 16'd29635, 16'd2958, 16'd5062, 16'd63843, 16'd16971, 16'd26055, 16'd4344, 16'd42053, 16'd39767, 16'd45, 16'd60371});
	test_expansion(128'h1c2a895c86322502d4b582b148b19757, {16'd55351, 16'd10924, 16'd11575, 16'd24401, 16'd40731, 16'd42595, 16'd20685, 16'd35647, 16'd58652, 16'd39687, 16'd8607, 16'd43995, 16'd41173, 16'd41381, 16'd4649, 16'd23364, 16'd36195, 16'd29508, 16'd11117, 16'd34462, 16'd10563, 16'd35194, 16'd63555, 16'd6256, 16'd19038, 16'd55454});
	test_expansion(128'hf747bedfa21bddb326e45609e21631c5, {16'd41192, 16'd23223, 16'd26985, 16'd41703, 16'd11988, 16'd13288, 16'd15076, 16'd26895, 16'd37579, 16'd42020, 16'd8978, 16'd51104, 16'd58653, 16'd12793, 16'd56558, 16'd658, 16'd23301, 16'd30509, 16'd58402, 16'd29275, 16'd27389, 16'd26328, 16'd1003, 16'd24774, 16'd48668, 16'd17594});
	test_expansion(128'hb01c2ca257ec0241b2a7641e7419be56, {16'd58695, 16'd16985, 16'd44320, 16'd43608, 16'd51368, 16'd56301, 16'd33336, 16'd3339, 16'd65390, 16'd21707, 16'd8880, 16'd31187, 16'd28110, 16'd6479, 16'd10885, 16'd49534, 16'd22690, 16'd57574, 16'd41777, 16'd48672, 16'd13420, 16'd64309, 16'd8121, 16'd64729, 16'd1785, 16'd38485});
	test_expansion(128'hb280fe88249919a694bf979f0636fd08, {16'd64247, 16'd30425, 16'd20249, 16'd20787, 16'd13978, 16'd31644, 16'd44027, 16'd40020, 16'd42217, 16'd34065, 16'd43073, 16'd60424, 16'd29526, 16'd27585, 16'd7741, 16'd3995, 16'd29886, 16'd36964, 16'd54300, 16'd60774, 16'd36840, 16'd38666, 16'd9344, 16'd32044, 16'd47939, 16'd4371});
	test_expansion(128'h5866361118e76bacc6c1b61d00aaeb0b, {16'd64179, 16'd49769, 16'd31947, 16'd34752, 16'd52029, 16'd19084, 16'd11593, 16'd535, 16'd42664, 16'd35470, 16'd64571, 16'd63992, 16'd64784, 16'd30128, 16'd23274, 16'd50071, 16'd18544, 16'd28771, 16'd53197, 16'd5711, 16'd56536, 16'd27336, 16'd530, 16'd63652, 16'd46142, 16'd50973});
	test_expansion(128'h7c0c4473e8f9cccabf3ad0ef7ba9207d, {16'd62995, 16'd61097, 16'd40328, 16'd46803, 16'd20706, 16'd7209, 16'd9321, 16'd52446, 16'd46598, 16'd41474, 16'd47665, 16'd61097, 16'd63654, 16'd55877, 16'd54904, 16'd12083, 16'd35707, 16'd16061, 16'd20600, 16'd39061, 16'd3459, 16'd36308, 16'd25989, 16'd7447, 16'd42671, 16'd8757});
	test_expansion(128'h0d2b12436755e246cefee1ab27f665da, {16'd4464, 16'd35091, 16'd56453, 16'd17735, 16'd46762, 16'd25158, 16'd54237, 16'd53113, 16'd30911, 16'd30382, 16'd41513, 16'd46354, 16'd56978, 16'd64220, 16'd28658, 16'd39505, 16'd2651, 16'd33120, 16'd44891, 16'd19632, 16'd60203, 16'd62526, 16'd52223, 16'd953, 16'd15635, 16'd49764});
	test_expansion(128'he7c70a81cb2a83b49e154d646e32d22c, {16'd35515, 16'd34339, 16'd48662, 16'd38939, 16'd19316, 16'd53292, 16'd45236, 16'd53654, 16'd62199, 16'd50159, 16'd23901, 16'd1936, 16'd35176, 16'd43601, 16'd60199, 16'd31968, 16'd10888, 16'd9071, 16'd28473, 16'd37140, 16'd41579, 16'd39704, 16'd2282, 16'd7406, 16'd28662, 16'd14342});
	test_expansion(128'hb635543caf331e36a66d8d7c8fac22b0, {16'd37716, 16'd46708, 16'd49402, 16'd60678, 16'd43322, 16'd10704, 16'd36876, 16'd40380, 16'd44711, 16'd46512, 16'd59585, 16'd48425, 16'd63133, 16'd51524, 16'd17701, 16'd33697, 16'd42706, 16'd13474, 16'd30575, 16'd59164, 16'd51720, 16'd1559, 16'd14045, 16'd31286, 16'd41588, 16'd32735});
	test_expansion(128'h34ea3ccd7c12cd905fee2a9fe4354e63, {16'd33197, 16'd34454, 16'd53410, 16'd57707, 16'd32690, 16'd64454, 16'd9184, 16'd26251, 16'd10358, 16'd36831, 16'd16654, 16'd5485, 16'd4391, 16'd47927, 16'd48772, 16'd50982, 16'd23561, 16'd20201, 16'd25704, 16'd13499, 16'd39419, 16'd30776, 16'd64428, 16'd21211, 16'd63902, 16'd6546});
	test_expansion(128'hfc5591ea1cff7c30cfbd429269816a83, {16'd27334, 16'd49314, 16'd17648, 16'd3151, 16'd56720, 16'd7292, 16'd5054, 16'd11326, 16'd30771, 16'd51147, 16'd35670, 16'd37, 16'd15587, 16'd5654, 16'd28774, 16'd21832, 16'd61508, 16'd11311, 16'd15820, 16'd64392, 16'd5051, 16'd6729, 16'd40855, 16'd61376, 16'd15292, 16'd54202});
	test_expansion(128'hb1c88d41120ef8a2438c91fa51c27516, {16'd48665, 16'd6605, 16'd52415, 16'd52780, 16'd33702, 16'd24697, 16'd63998, 16'd50535, 16'd23517, 16'd22270, 16'd22758, 16'd56039, 16'd52749, 16'd22340, 16'd12420, 16'd24705, 16'd5092, 16'd7786, 16'd5286, 16'd58389, 16'd25165, 16'd35750, 16'd18097, 16'd62119, 16'd46387, 16'd55885});
	test_expansion(128'h45c9ca97d635e4abbf75d0f2e470ba6c, {16'd18039, 16'd31411, 16'd48859, 16'd23569, 16'd55811, 16'd9568, 16'd52101, 16'd9125, 16'd23005, 16'd6690, 16'd3883, 16'd40853, 16'd61566, 16'd27045, 16'd52703, 16'd38220, 16'd24126, 16'd12089, 16'd29161, 16'd55222, 16'd27619, 16'd30039, 16'd199, 16'd19687, 16'd2853, 16'd57374});
	test_expansion(128'h9d3d6064d4db16b685a550b2bcf02b96, {16'd24558, 16'd24722, 16'd1522, 16'd61342, 16'd14222, 16'd49185, 16'd5639, 16'd5560, 16'd14022, 16'd12848, 16'd21777, 16'd18029, 16'd44422, 16'd51195, 16'd57625, 16'd60820, 16'd41336, 16'd60360, 16'd26157, 16'd62319, 16'd23267, 16'd42208, 16'd57821, 16'd15095, 16'd47519, 16'd2472});
	test_expansion(128'h47a92389d43aba2b87147306a44a1cf9, {16'd37664, 16'd24729, 16'd9796, 16'd5727, 16'd22583, 16'd48967, 16'd25696, 16'd7289, 16'd13210, 16'd24673, 16'd6872, 16'd44304, 16'd44048, 16'd21732, 16'd61062, 16'd16236, 16'd60546, 16'd49, 16'd51668, 16'd1174, 16'd3253, 16'd27321, 16'd12779, 16'd64246, 16'd35477, 16'd22187});
	test_expansion(128'hea09da035096dfbcd158f8536567041a, {16'd44974, 16'd26547, 16'd61197, 16'd47855, 16'd12254, 16'd39258, 16'd54931, 16'd58428, 16'd50615, 16'd20997, 16'd14597, 16'd43607, 16'd38455, 16'd26761, 16'd1042, 16'd46752, 16'd9587, 16'd31638, 16'd55379, 16'd46405, 16'd4005, 16'd30740, 16'd55603, 16'd64693, 16'd50541, 16'd7424});
	test_expansion(128'h20f469cbe916a3d97d74e6c02d5b60b4, {16'd11827, 16'd15413, 16'd24223, 16'd14404, 16'd26688, 16'd45441, 16'd46592, 16'd53073, 16'd41972, 16'd47625, 16'd50791, 16'd7717, 16'd9173, 16'd26645, 16'd64204, 16'd43096, 16'd21423, 16'd24015, 16'd1938, 16'd12667, 16'd3865, 16'd39349, 16'd18634, 16'd48616, 16'd16045, 16'd2703});
	test_expansion(128'h0e0f440aa4915925ddbf885a58c71c33, {16'd28276, 16'd50464, 16'd61179, 16'd4650, 16'd51213, 16'd9414, 16'd45263, 16'd7655, 16'd1323, 16'd35969, 16'd130, 16'd65213, 16'd37972, 16'd47953, 16'd12685, 16'd11149, 16'd41727, 16'd11805, 16'd35970, 16'd3460, 16'd10906, 16'd22150, 16'd8147, 16'd54722, 16'd56210, 16'd33798});
	test_expansion(128'he20bb0167e2ba14fa68587bbd7ca0bab, {16'd61100, 16'd39507, 16'd63229, 16'd5212, 16'd10306, 16'd40660, 16'd14948, 16'd15080, 16'd64111, 16'd34096, 16'd15401, 16'd46555, 16'd57086, 16'd26974, 16'd2111, 16'd34796, 16'd58828, 16'd62314, 16'd55571, 16'd65149, 16'd13865, 16'd4587, 16'd7535, 16'd34870, 16'd10831, 16'd37817});
	test_expansion(128'hfa287fac0e64cc86650f6219fdcf2a6e, {16'd48284, 16'd63969, 16'd33265, 16'd59509, 16'd29244, 16'd5708, 16'd51595, 16'd1400, 16'd30139, 16'd5031, 16'd61619, 16'd49190, 16'd19154, 16'd45862, 16'd20623, 16'd24353, 16'd45448, 16'd56631, 16'd34120, 16'd63612, 16'd65084, 16'd19422, 16'd6716, 16'd51026, 16'd52591, 16'd46244});
	test_expansion(128'hf9b57551fdb8a9bb62df7cae98fe7887, {16'd13678, 16'd19777, 16'd38264, 16'd6512, 16'd54374, 16'd39812, 16'd39006, 16'd11181, 16'd8037, 16'd11369, 16'd55823, 16'd33158, 16'd8589, 16'd3958, 16'd49275, 16'd47112, 16'd16187, 16'd23214, 16'd54050, 16'd50261, 16'd6649, 16'd53566, 16'd21389, 16'd28446, 16'd35160, 16'd45046});
	test_expansion(128'hd3cd39431f780c093cccf5ee0d1d60a7, {16'd19058, 16'd41456, 16'd40461, 16'd15678, 16'd31381, 16'd6924, 16'd31722, 16'd16706, 16'd43801, 16'd27201, 16'd20889, 16'd34671, 16'd53674, 16'd29322, 16'd9392, 16'd37951, 16'd44683, 16'd54556, 16'd55684, 16'd21488, 16'd53786, 16'd11962, 16'd23115, 16'd44925, 16'd17562, 16'd47092});
	test_expansion(128'hf36044f384975ffc9cb6051a2a9bb3cc, {16'd2308, 16'd22992, 16'd53973, 16'd44719, 16'd1054, 16'd27545, 16'd33371, 16'd31969, 16'd23125, 16'd52836, 16'd39844, 16'd8624, 16'd42330, 16'd738, 16'd45663, 16'd35086, 16'd1558, 16'd56136, 16'd31675, 16'd34294, 16'd27155, 16'd22439, 16'd18361, 16'd44244, 16'd63884, 16'd23755});
	test_expansion(128'h842313516da2f1217494e3898b0e5082, {16'd56658, 16'd47586, 16'd21841, 16'd17956, 16'd58387, 16'd39835, 16'd2308, 16'd58056, 16'd40240, 16'd50760, 16'd61373, 16'd51992, 16'd9121, 16'd3933, 16'd47025, 16'd15035, 16'd15272, 16'd21048, 16'd46499, 16'd14044, 16'd15021, 16'd7544, 16'd45339, 16'd32491, 16'd14744, 16'd13057});
	test_expansion(128'hd79e85ebfddaeb1e319b38c064f4ee72, {16'd45914, 16'd48970, 16'd27146, 16'd13674, 16'd5661, 16'd46333, 16'd1817, 16'd14462, 16'd1422, 16'd22740, 16'd28244, 16'd63483, 16'd26007, 16'd28582, 16'd39164, 16'd17975, 16'd11994, 16'd46029, 16'd34535, 16'd15185, 16'd57143, 16'd7474, 16'd23817, 16'd41801, 16'd52842, 16'd26064});
	test_expansion(128'h64a11b957e7a595731942bb670807d64, {16'd60175, 16'd30409, 16'd63496, 16'd56388, 16'd48979, 16'd47203, 16'd9792, 16'd13889, 16'd55634, 16'd31770, 16'd53636, 16'd9902, 16'd24106, 16'd20799, 16'd35115, 16'd48499, 16'd61911, 16'd63749, 16'd37423, 16'd19861, 16'd50414, 16'd7381, 16'd30981, 16'd45503, 16'd6006, 16'd36261});
	test_expansion(128'hd01c7b08def4d0cfafe78c9781903a34, {16'd8171, 16'd9711, 16'd24475, 16'd30340, 16'd32222, 16'd55185, 16'd35975, 16'd18358, 16'd3522, 16'd3025, 16'd55188, 16'd34092, 16'd30756, 16'd15231, 16'd14893, 16'd10514, 16'd32179, 16'd40844, 16'd19035, 16'd57488, 16'd54954, 16'd4466, 16'd28296, 16'd64786, 16'd17609, 16'd55395});
	test_expansion(128'hce25671b4e9fb4c218efd4df747d53f0, {16'd19405, 16'd27549, 16'd28069, 16'd42099, 16'd44435, 16'd32681, 16'd59578, 16'd38795, 16'd19099, 16'd848, 16'd47076, 16'd29766, 16'd38922, 16'd9419, 16'd19185, 16'd41739, 16'd63424, 16'd49046, 16'd36114, 16'd49462, 16'd25883, 16'd9714, 16'd1831, 16'd7292, 16'd35367, 16'd40657});
	test_expansion(128'h1724ff9215e77f253910222fee0c0886, {16'd27821, 16'd38947, 16'd57818, 16'd3176, 16'd23517, 16'd38914, 16'd11395, 16'd39364, 16'd34259, 16'd4562, 16'd60995, 16'd44567, 16'd63998, 16'd57201, 16'd35716, 16'd61105, 16'd59773, 16'd52749, 16'd3997, 16'd39841, 16'd41755, 16'd40911, 16'd57045, 16'd14154, 16'd14025, 16'd18672});
	test_expansion(128'hc5513a4ce4fd7e29d47d02f0b1b05c2d, {16'd9414, 16'd46590, 16'd62336, 16'd6561, 16'd45301, 16'd25235, 16'd13249, 16'd987, 16'd27831, 16'd39912, 16'd44418, 16'd62960, 16'd8953, 16'd40236, 16'd31796, 16'd44607, 16'd13111, 16'd10256, 16'd13358, 16'd16625, 16'd28989, 16'd56108, 16'd55234, 16'd57904, 16'd44738, 16'd24600});
	test_expansion(128'hd10244070588668c9f2852e300402c7a, {16'd63555, 16'd54020, 16'd38608, 16'd33054, 16'd22153, 16'd41810, 16'd64865, 16'd18316, 16'd34544, 16'd38308, 16'd4649, 16'd12725, 16'd33935, 16'd28613, 16'd27833, 16'd48757, 16'd21400, 16'd13993, 16'd22579, 16'd20502, 16'd15810, 16'd30367, 16'd7853, 16'd2904, 16'd64270, 16'd764});
	test_expansion(128'hd4447c08975e6adda0908b6b2674e485, {16'd52696, 16'd51183, 16'd16656, 16'd61525, 16'd5638, 16'd28846, 16'd41961, 16'd44920, 16'd11924, 16'd2242, 16'd56671, 16'd48053, 16'd11180, 16'd25390, 16'd22789, 16'd14428, 16'd38715, 16'd46028, 16'd1553, 16'd62242, 16'd44082, 16'd63629, 16'd59074, 16'd35459, 16'd42851, 16'd24890});
	test_expansion(128'hff4655f092f2574c644ceb85569c35bd, {16'd31186, 16'd55918, 16'd3488, 16'd48295, 16'd47863, 16'd49624, 16'd17216, 16'd40358, 16'd28896, 16'd32896, 16'd1199, 16'd45423, 16'd8066, 16'd42361, 16'd52444, 16'd46167, 16'd31295, 16'd56801, 16'd33203, 16'd6438, 16'd40584, 16'd54306, 16'd13607, 16'd2320, 16'd23699, 16'd41449});
	test_expansion(128'h0b19d78d991f4cf994ec68dc1289f819, {16'd3073, 16'd59041, 16'd16129, 16'd21468, 16'd12865, 16'd57122, 16'd35074, 16'd1097, 16'd51545, 16'd1541, 16'd183, 16'd21126, 16'd16760, 16'd34214, 16'd50054, 16'd15556, 16'd6426, 16'd60811, 16'd43502, 16'd62429, 16'd27667, 16'd44249, 16'd38158, 16'd24473, 16'd40570, 16'd33687});
	test_expansion(128'h4b6b6d214c46e7683825304074f57ffe, {16'd44991, 16'd52565, 16'd9992, 16'd49862, 16'd57305, 16'd364, 16'd42206, 16'd26990, 16'd36053, 16'd1129, 16'd36662, 16'd51161, 16'd35561, 16'd46338, 16'd31394, 16'd56056, 16'd12907, 16'd52869, 16'd14669, 16'd37200, 16'd65336, 16'd13774, 16'd45082, 16'd2927, 16'd24594, 16'd47230});
	test_expansion(128'h573e88b1b7f6bff0df5b5200794aa28e, {16'd39191, 16'd36053, 16'd63446, 16'd18885, 16'd6166, 16'd23613, 16'd3046, 16'd1261, 16'd45430, 16'd33067, 16'd28281, 16'd18894, 16'd3032, 16'd53888, 16'd61085, 16'd14263, 16'd1561, 16'd60896, 16'd55253, 16'd29832, 16'd27170, 16'd28180, 16'd9815, 16'd35065, 16'd27822, 16'd44339});
	test_expansion(128'h41197a3b67cee1befcfbf617942a4984, {16'd34084, 16'd18451, 16'd64846, 16'd60117, 16'd49269, 16'd49942, 16'd37785, 16'd44899, 16'd7585, 16'd11056, 16'd42504, 16'd58479, 16'd4440, 16'd38243, 16'd4329, 16'd13462, 16'd49894, 16'd54966, 16'd58930, 16'd15334, 16'd45567, 16'd10660, 16'd6316, 16'd32488, 16'd34843, 16'd37117});
	test_expansion(128'ha51619615a39eef202fb3aeb124406aa, {16'd30371, 16'd2407, 16'd13738, 16'd16814, 16'd11269, 16'd62770, 16'd36810, 16'd2479, 16'd53832, 16'd59293, 16'd19006, 16'd50565, 16'd22090, 16'd61031, 16'd62679, 16'd65410, 16'd15997, 16'd17520, 16'd1396, 16'd18667, 16'd49839, 16'd35877, 16'd12681, 16'd62370, 16'd40949, 16'd23178});
	test_expansion(128'h0806e59fa2efcc95cbe5ec25b52908a4, {16'd27161, 16'd59272, 16'd54868, 16'd9164, 16'd38296, 16'd54160, 16'd2702, 16'd62172, 16'd12112, 16'd21949, 16'd8078, 16'd13293, 16'd51304, 16'd17950, 16'd5922, 16'd20261, 16'd52574, 16'd6339, 16'd57603, 16'd6026, 16'd17176, 16'd39138, 16'd11739, 16'd54678, 16'd18977, 16'd62829});
	test_expansion(128'h445bf08ab7b5feb16ebc996ed3d9a633, {16'd60532, 16'd36331, 16'd56764, 16'd25947, 16'd1492, 16'd52958, 16'd21682, 16'd33615, 16'd59748, 16'd50606, 16'd14157, 16'd10211, 16'd20093, 16'd2756, 16'd24064, 16'd39595, 16'd303, 16'd16772, 16'd58385, 16'd41318, 16'd47393, 16'd51389, 16'd46065, 16'd63296, 16'd15314, 16'd42203});
	test_expansion(128'h59beb2b8b114b7a16f1ab8fa336d46a9, {16'd28963, 16'd1782, 16'd21135, 16'd16933, 16'd39110, 16'd9798, 16'd2462, 16'd42435, 16'd33639, 16'd55302, 16'd56620, 16'd11689, 16'd37456, 16'd20453, 16'd39636, 16'd63136, 16'd35886, 16'd38956, 16'd38547, 16'd54087, 16'd56275, 16'd60378, 16'd34200, 16'd12408, 16'd58091, 16'd26883});
	test_expansion(128'hf8f944bbc168a6a444a8e76e44c72712, {16'd22941, 16'd39772, 16'd6318, 16'd434, 16'd48649, 16'd17143, 16'd27564, 16'd57967, 16'd14116, 16'd12888, 16'd14947, 16'd48877, 16'd55704, 16'd58587, 16'd64349, 16'd8415, 16'd33267, 16'd62137, 16'd36871, 16'd24090, 16'd7828, 16'd55110, 16'd39725, 16'd55844, 16'd63182, 16'd61051});
	test_expansion(128'h1dc57fd61b1c0f52c14c58808bcfd8fc, {16'd47676, 16'd9169, 16'd33080, 16'd16674, 16'd39716, 16'd56685, 16'd24220, 16'd31253, 16'd10530, 16'd28592, 16'd21681, 16'd6824, 16'd11776, 16'd2039, 16'd34179, 16'd23610, 16'd24282, 16'd4932, 16'd30780, 16'd22874, 16'd33892, 16'd16564, 16'd279, 16'd19781, 16'd18646, 16'd28905});
	test_expansion(128'hd73609febd5f3ab10cf6b1332f97b6b3, {16'd61118, 16'd10952, 16'd219, 16'd28362, 16'd64413, 16'd21837, 16'd22189, 16'd12566, 16'd15982, 16'd45061, 16'd6459, 16'd45431, 16'd26046, 16'd31731, 16'd8207, 16'd13174, 16'd42477, 16'd36720, 16'd8144, 16'd33055, 16'd34176, 16'd47895, 16'd55514, 16'd33271, 16'd48280, 16'd30372});
	test_expansion(128'hc38bd1be8676bb78fa859ecd99a952b5, {16'd34344, 16'd40670, 16'd33643, 16'd22295, 16'd7104, 16'd18908, 16'd9810, 16'd11867, 16'd50949, 16'd19516, 16'd16812, 16'd34438, 16'd27117, 16'd56086, 16'd37655, 16'd44415, 16'd3105, 16'd3851, 16'd62523, 16'd44581, 16'd52142, 16'd56144, 16'd28404, 16'd64635, 16'd14786, 16'd38928});
	test_expansion(128'hcf24e81953eff1a36168ddcaa3d6ef91, {16'd34548, 16'd14964, 16'd54626, 16'd42494, 16'd54998, 16'd18826, 16'd65089, 16'd11573, 16'd49410, 16'd41259, 16'd30468, 16'd6423, 16'd58517, 16'd53294, 16'd34479, 16'd6979, 16'd62398, 16'd52295, 16'd8958, 16'd61228, 16'd27717, 16'd63022, 16'd2285, 16'd22972, 16'd52853, 16'd17804});
	test_expansion(128'h4d34a44e430af3d561c2ec1f88e38d00, {16'd54649, 16'd27005, 16'd46242, 16'd32472, 16'd26724, 16'd8203, 16'd41948, 16'd29861, 16'd6541, 16'd46716, 16'd63887, 16'd16189, 16'd32427, 16'd29812, 16'd36109, 16'd37425, 16'd63649, 16'd51819, 16'd35381, 16'd52582, 16'd59730, 16'd3985, 16'd13154, 16'd46875, 16'd15074, 16'd64558});
	test_expansion(128'h9d001201ff3cd9680b4527cdd5a80a89, {16'd58154, 16'd44728, 16'd6150, 16'd17615, 16'd57237, 16'd31425, 16'd58191, 16'd44009, 16'd52112, 16'd4254, 16'd34517, 16'd51639, 16'd34182, 16'd63906, 16'd51926, 16'd23894, 16'd9523, 16'd16179, 16'd42587, 16'd21232, 16'd45596, 16'd4562, 16'd8091, 16'd1654, 16'd58092, 16'd64782});
	test_expansion(128'h14bc2118217951eb7883a9869267036d, {16'd52581, 16'd39519, 16'd25812, 16'd18618, 16'd54472, 16'd46601, 16'd8978, 16'd9556, 16'd29404, 16'd43885, 16'd40146, 16'd35283, 16'd26101, 16'd58758, 16'd63820, 16'd12804, 16'd22194, 16'd37675, 16'd49630, 16'd45220, 16'd58595, 16'd2267, 16'd48992, 16'd29038, 16'd35852, 16'd40110});
	test_expansion(128'h84f7ee86b51ea081d3c196cabc7f3190, {16'd51020, 16'd17959, 16'd42960, 16'd2998, 16'd32098, 16'd9287, 16'd44905, 16'd26099, 16'd54406, 16'd44261, 16'd17710, 16'd1398, 16'd42265, 16'd25545, 16'd51952, 16'd20347, 16'd58600, 16'd2310, 16'd60949, 16'd7704, 16'd5970, 16'd59095, 16'd26768, 16'd45307, 16'd12514, 16'd63169});
	test_expansion(128'h8880d663d4d6c9721cb5eaaf30abd89d, {16'd30079, 16'd22137, 16'd41627, 16'd16175, 16'd13745, 16'd40264, 16'd16452, 16'd22826, 16'd47876, 16'd8600, 16'd5726, 16'd20014, 16'd4596, 16'd56582, 16'd11485, 16'd40117, 16'd43918, 16'd24684, 16'd33255, 16'd19783, 16'd34513, 16'd48630, 16'd27409, 16'd63566, 16'd17618, 16'd6046});
	test_expansion(128'ha5dd8520a4e4889441b4031440da0049, {16'd36603, 16'd4618, 16'd62784, 16'd52084, 16'd2100, 16'd51641, 16'd65092, 16'd13053, 16'd46183, 16'd42699, 16'd34460, 16'd12887, 16'd16241, 16'd9214, 16'd20297, 16'd27114, 16'd1455, 16'd47945, 16'd32873, 16'd20297, 16'd31858, 16'd3979, 16'd49616, 16'd16749, 16'd60417, 16'd32230});
	test_expansion(128'h0d30b20bee870120e789dec9cd9bbf38, {16'd34714, 16'd58075, 16'd62079, 16'd8630, 16'd13009, 16'd34930, 16'd49967, 16'd12108, 16'd47639, 16'd5815, 16'd43572, 16'd4419, 16'd19727, 16'd39020, 16'd55779, 16'd65317, 16'd22799, 16'd29380, 16'd28803, 16'd3220, 16'd37084, 16'd1176, 16'd29452, 16'd44725, 16'd43174, 16'd47542});
	test_expansion(128'h6d0f94bfd6c8d8f7a60b8df33bdd005b, {16'd64399, 16'd36371, 16'd6733, 16'd53465, 16'd46734, 16'd7535, 16'd11055, 16'd41357, 16'd57114, 16'd58793, 16'd16865, 16'd53208, 16'd44699, 16'd9543, 16'd22505, 16'd51942, 16'd47330, 16'd49755, 16'd59513, 16'd29353, 16'd17300, 16'd43039, 16'd59143, 16'd26278, 16'd21612, 16'd43004});
	test_expansion(128'h93ceb9bb23c0579c603cd1ef3948bcc6, {16'd6829, 16'd18935, 16'd24650, 16'd44362, 16'd6816, 16'd60776, 16'd23929, 16'd17532, 16'd25104, 16'd40895, 16'd36809, 16'd5300, 16'd43180, 16'd38672, 16'd550, 16'd34673, 16'd51297, 16'd57759, 16'd62488, 16'd61795, 16'd37198, 16'd49682, 16'd6622, 16'd62430, 16'd6087, 16'd35654});
	test_expansion(128'hb3ca716e92e3d653631ecfc994a9567c, {16'd23446, 16'd34277, 16'd6022, 16'd46603, 16'd51393, 16'd63081, 16'd27653, 16'd11018, 16'd26711, 16'd47396, 16'd31436, 16'd28470, 16'd6535, 16'd34769, 16'd65388, 16'd37739, 16'd28026, 16'd40248, 16'd63655, 16'd13191, 16'd57631, 16'd35021, 16'd22184, 16'd7543, 16'd10167, 16'd42038});
	test_expansion(128'h38dc3c98fbbcbc574db1719752ae327c, {16'd21148, 16'd26155, 16'd51169, 16'd55274, 16'd47876, 16'd11722, 16'd56766, 16'd27223, 16'd64656, 16'd27575, 16'd9693, 16'd14085, 16'd40256, 16'd53381, 16'd54989, 16'd52365, 16'd48194, 16'd312, 16'd38229, 16'd6671, 16'd62025, 16'd30324, 16'd55369, 16'd59828, 16'd41882, 16'd30033});
	test_expansion(128'h6a6fcd17c3cdc74b2956ad9d6ca5b72f, {16'd11906, 16'd29412, 16'd32217, 16'd45401, 16'd4108, 16'd55762, 16'd44455, 16'd8967, 16'd48064, 16'd44767, 16'd38909, 16'd46865, 16'd5535, 16'd16168, 16'd18871, 16'd62275, 16'd27512, 16'd59970, 16'd44671, 16'd57687, 16'd61445, 16'd34672, 16'd4656, 16'd50850, 16'd33807, 16'd1726});
	test_expansion(128'hffac413368725fd025188024301cad6b, {16'd13300, 16'd36156, 16'd26391, 16'd48118, 16'd31203, 16'd2491, 16'd16609, 16'd58435, 16'd26079, 16'd43438, 16'd7572, 16'd56305, 16'd48802, 16'd46581, 16'd25394, 16'd24602, 16'd14350, 16'd10882, 16'd35653, 16'd49015, 16'd35680, 16'd29525, 16'd40550, 16'd42116, 16'd5205, 16'd11926});
	test_expansion(128'h1d7cb8cbd47cc5a0d1377578242a9203, {16'd1158, 16'd46540, 16'd20926, 16'd42466, 16'd44319, 16'd37164, 16'd51509, 16'd17573, 16'd55220, 16'd22449, 16'd9043, 16'd158, 16'd37011, 16'd45943, 16'd25181, 16'd4150, 16'd6227, 16'd16326, 16'd51192, 16'd52767, 16'd23782, 16'd23699, 16'd12357, 16'd1027, 16'd34196, 16'd19760});
	test_expansion(128'h1bfd3c927d518ac22512b673e1101604, {16'd25017, 16'd15680, 16'd46041, 16'd45295, 16'd16673, 16'd57860, 16'd14269, 16'd48247, 16'd35749, 16'd7297, 16'd14238, 16'd46329, 16'd35686, 16'd43917, 16'd54704, 16'd55486, 16'd19920, 16'd43082, 16'd62942, 16'd22111, 16'd2052, 16'd54201, 16'd32545, 16'd7891, 16'd95, 16'd47174});
	test_expansion(128'hff9570ff4abed88805182bb998cc289c, {16'd14248, 16'd56697, 16'd12080, 16'd15273, 16'd1335, 16'd12706, 16'd53381, 16'd4758, 16'd20076, 16'd16529, 16'd21441, 16'd34099, 16'd5508, 16'd23200, 16'd28703, 16'd18582, 16'd33732, 16'd4170, 16'd63610, 16'd4082, 16'd54790, 16'd44393, 16'd39892, 16'd16610, 16'd38066, 16'd20009});
	test_expansion(128'h8af6bb943dbd28f6fec66989f7fbc8fa, {16'd8843, 16'd7128, 16'd25649, 16'd59147, 16'd3299, 16'd14526, 16'd17742, 16'd2301, 16'd19637, 16'd24780, 16'd45203, 16'd30852, 16'd25480, 16'd45848, 16'd63977, 16'd34533, 16'd559, 16'd33741, 16'd49351, 16'd41918, 16'd56760, 16'd24283, 16'd5189, 16'd24555, 16'd9849, 16'd7149});
	test_expansion(128'h81e87eccc9b9ef154e10d6b213280fab, {16'd43407, 16'd23752, 16'd58900, 16'd4939, 16'd44086, 16'd25027, 16'd44588, 16'd15475, 16'd20510, 16'd29972, 16'd48096, 16'd54561, 16'd22058, 16'd3895, 16'd17709, 16'd51455, 16'd6645, 16'd45860, 16'd50731, 16'd50303, 16'd54098, 16'd23168, 16'd828, 16'd14930, 16'd12537, 16'd6404});
	test_expansion(128'h7ec4147554d4c89e5ddd58afdf495ac2, {16'd36563, 16'd13676, 16'd7992, 16'd35308, 16'd8563, 16'd19492, 16'd12265, 16'd25995, 16'd2702, 16'd31461, 16'd3819, 16'd49101, 16'd63589, 16'd43001, 16'd11668, 16'd24906, 16'd13398, 16'd4841, 16'd52602, 16'd64729, 16'd43341, 16'd10475, 16'd63568, 16'd20263, 16'd4739, 16'd40915});
	test_expansion(128'h2409656ccbc41cc5df130992800c387e, {16'd61779, 16'd22145, 16'd61783, 16'd53504, 16'd41837, 16'd36871, 16'd39872, 16'd2558, 16'd13447, 16'd41278, 16'd59163, 16'd17698, 16'd2435, 16'd63773, 16'd14974, 16'd63566, 16'd55536, 16'd40612, 16'd61543, 16'd6372, 16'd28241, 16'd52474, 16'd22877, 16'd10843, 16'd33954, 16'd52975});
	test_expansion(128'h6337d405abe925cb18e8e7ac918efb2b, {16'd49680, 16'd18884, 16'd11115, 16'd36639, 16'd31487, 16'd40628, 16'd27951, 16'd48163, 16'd54221, 16'd4806, 16'd26251, 16'd2519, 16'd50603, 16'd25089, 16'd13683, 16'd61236, 16'd37468, 16'd44902, 16'd30360, 16'd30112, 16'd33115, 16'd15684, 16'd41862, 16'd10528, 16'd37549, 16'd19014});
	test_expansion(128'hc68e648064d13bf9f67433ec85ff8c77, {16'd64974, 16'd44984, 16'd52628, 16'd54487, 16'd19463, 16'd28741, 16'd33667, 16'd13910, 16'd21258, 16'd12344, 16'd20618, 16'd62154, 16'd3134, 16'd10399, 16'd427, 16'd34652, 16'd47948, 16'd49019, 16'd15406, 16'd723, 16'd21136, 16'd31541, 16'd44706, 16'd33093, 16'd58593, 16'd28610});
	test_expansion(128'h76f76c4d6600fbc019aeea3d94b96860, {16'd12804, 16'd33765, 16'd47182, 16'd27416, 16'd38525, 16'd5996, 16'd45585, 16'd61479, 16'd50645, 16'd27356, 16'd59382, 16'd5999, 16'd54671, 16'd63285, 16'd59673, 16'd44840, 16'd23142, 16'd14116, 16'd29923, 16'd53747, 16'd30637, 16'd31027, 16'd39737, 16'd51560, 16'd63680, 16'd15813});
	test_expansion(128'hbf8471f513132ef77078eb411f01b8b7, {16'd9706, 16'd21182, 16'd50198, 16'd15028, 16'd17409, 16'd55717, 16'd41580, 16'd49587, 16'd24423, 16'd14465, 16'd52034, 16'd53292, 16'd57398, 16'd43390, 16'd64738, 16'd54362, 16'd20445, 16'd44526, 16'd21728, 16'd18956, 16'd19435, 16'd60549, 16'd6592, 16'd26821, 16'd2708, 16'd39480});
	test_expansion(128'hf16866c4ba3ee1acc40f53f43a042400, {16'd28520, 16'd5564, 16'd16159, 16'd37986, 16'd11959, 16'd5252, 16'd28334, 16'd9666, 16'd32749, 16'd46439, 16'd46607, 16'd36139, 16'd59722, 16'd1792, 16'd45165, 16'd40753, 16'd32196, 16'd23906, 16'd46840, 16'd22013, 16'd22783, 16'd5248, 16'd16080, 16'd44885, 16'd51745, 16'd34572});
	test_expansion(128'h7cc7b73a351ac73d6b573ea5fa1c1bd2, {16'd37671, 16'd11688, 16'd16924, 16'd52207, 16'd11192, 16'd55788, 16'd34274, 16'd57394, 16'd22663, 16'd46309, 16'd29176, 16'd26786, 16'd23429, 16'd21931, 16'd47700, 16'd41624, 16'd1199, 16'd55194, 16'd27912, 16'd12982, 16'd52762, 16'd3829, 16'd46649, 16'd24831, 16'd62220, 16'd60038});
	test_expansion(128'h16ca7a9889c4d9ce03b95094fa2631bc, {16'd60380, 16'd48177, 16'd32440, 16'd43796, 16'd52174, 16'd10864, 16'd47844, 16'd20316, 16'd3188, 16'd53483, 16'd23483, 16'd3770, 16'd53676, 16'd2962, 16'd29404, 16'd62678, 16'd1868, 16'd50953, 16'd57758, 16'd49107, 16'd57456, 16'd24175, 16'd4244, 16'd54025, 16'd2925, 16'd32624});
	test_expansion(128'hf145ff45631d688f62578cd7dffde1e6, {16'd57080, 16'd10802, 16'd54553, 16'd19116, 16'd24171, 16'd22836, 16'd24019, 16'd26734, 16'd40400, 16'd27043, 16'd38003, 16'd21109, 16'd47840, 16'd16927, 16'd2136, 16'd52552, 16'd54837, 16'd45470, 16'd58973, 16'd34407, 16'd9289, 16'd40619, 16'd41426, 16'd63593, 16'd9984, 16'd14367});
	test_expansion(128'h4076a57b1b3e312de854655d9b132ce6, {16'd17482, 16'd54407, 16'd22074, 16'd60702, 16'd914, 16'd14651, 16'd64835, 16'd61537, 16'd38410, 16'd8232, 16'd27212, 16'd18035, 16'd57486, 16'd7185, 16'd12094, 16'd21397, 16'd16569, 16'd34155, 16'd52644, 16'd18521, 16'd45572, 16'd9756, 16'd38372, 16'd38620, 16'd42726, 16'd12522});
	test_expansion(128'h40fd2400fbb5433ea1c4484e93106517, {16'd62477, 16'd48816, 16'd49247, 16'd35643, 16'd27062, 16'd53088, 16'd20749, 16'd51501, 16'd11139, 16'd20607, 16'd49206, 16'd13342, 16'd13412, 16'd46597, 16'd18597, 16'd11742, 16'd12853, 16'd5784, 16'd4465, 16'd45204, 16'd55500, 16'd35395, 16'd32052, 16'd4458, 16'd2078, 16'd36042});
	test_expansion(128'h10c61593f68927b30c2676979cd98561, {16'd13339, 16'd1326, 16'd20068, 16'd64349, 16'd62058, 16'd17701, 16'd23604, 16'd27814, 16'd9202, 16'd19126, 16'd61173, 16'd64095, 16'd29348, 16'd40016, 16'd45629, 16'd27601, 16'd38312, 16'd12726, 16'd11407, 16'd54346, 16'd60945, 16'd34200, 16'd46559, 16'd50910, 16'd23601, 16'd32743});
	test_expansion(128'hc500a6a2876cfb2b134a2d5c27094905, {16'd13742, 16'd2231, 16'd30110, 16'd23871, 16'd42841, 16'd15731, 16'd29620, 16'd623, 16'd7123, 16'd45590, 16'd6432, 16'd14377, 16'd25903, 16'd17327, 16'd44769, 16'd52049, 16'd29367, 16'd60834, 16'd36824, 16'd63441, 16'd19091, 16'd22364, 16'd42248, 16'd65300, 16'd26387, 16'd29078});
	test_expansion(128'h70a99150139475aab7854205047074e8, {16'd39198, 16'd43968, 16'd46826, 16'd18714, 16'd27349, 16'd14962, 16'd7770, 16'd13216, 16'd18986, 16'd9566, 16'd35270, 16'd40736, 16'd35232, 16'd21561, 16'd24981, 16'd53768, 16'd46547, 16'd8144, 16'd33934, 16'd2280, 16'd51061, 16'd1965, 16'd14090, 16'd9228, 16'd38221, 16'd63532});
	test_expansion(128'hba951db52919f1f7bef709f5726b2c23, {16'd3953, 16'd34974, 16'd35218, 16'd23177, 16'd15014, 16'd46980, 16'd19677, 16'd15019, 16'd50552, 16'd49827, 16'd9893, 16'd19647, 16'd35733, 16'd6317, 16'd39480, 16'd59071, 16'd43168, 16'd54881, 16'd39491, 16'd61056, 16'd64305, 16'd16741, 16'd23602, 16'd34872, 16'd49603, 16'd13310});
	test_expansion(128'h7102b0c0ffd8ef87a0409da8bb719880, {16'd45415, 16'd53042, 16'd51353, 16'd12015, 16'd28173, 16'd62785, 16'd57736, 16'd36978, 16'd41311, 16'd19119, 16'd30750, 16'd7552, 16'd473, 16'd15084, 16'd644, 16'd12376, 16'd4920, 16'd61953, 16'd53114, 16'd18738, 16'd39215, 16'd10543, 16'd5585, 16'd48952, 16'd12716, 16'd17396});
	test_expansion(128'h70f9ca5a60768987058d959ff83d1e2f, {16'd33724, 16'd45071, 16'd42643, 16'd28526, 16'd5406, 16'd27708, 16'd49286, 16'd18835, 16'd13556, 16'd42904, 16'd22181, 16'd64283, 16'd55071, 16'd27462, 16'd33796, 16'd43601, 16'd8163, 16'd29784, 16'd41598, 16'd30755, 16'd3525, 16'd3842, 16'd7027, 16'd62152, 16'd41767, 16'd62803});
	test_expansion(128'hf4e1056e823a816e177ae1eb40137c7a, {16'd27863, 16'd24141, 16'd9218, 16'd16404, 16'd11228, 16'd61737, 16'd10177, 16'd10618, 16'd52524, 16'd46009, 16'd27322, 16'd17066, 16'd55590, 16'd30360, 16'd23672, 16'd18085, 16'd51895, 16'd49463, 16'd1910, 16'd34352, 16'd13141, 16'd55339, 16'd10341, 16'd4636, 16'd51702, 16'd28137});
	test_expansion(128'h6f43aacacfa417f78dc7ffbfe811f331, {16'd46854, 16'd16515, 16'd7932, 16'd10774, 16'd29654, 16'd63628, 16'd7148, 16'd63577, 16'd15202, 16'd9673, 16'd39459, 16'd11982, 16'd43120, 16'd58002, 16'd57847, 16'd13581, 16'd58844, 16'd23511, 16'd40891, 16'd6260, 16'd5038, 16'd6990, 16'd50912, 16'd10618, 16'd62716, 16'd64010});
	test_expansion(128'h23e6f38df60339dd13065c6118af5447, {16'd26805, 16'd53942, 16'd53691, 16'd4987, 16'd21793, 16'd51976, 16'd27692, 16'd60656, 16'd63020, 16'd55186, 16'd39385, 16'd37019, 16'd48779, 16'd14930, 16'd38961, 16'd32735, 16'd43443, 16'd41899, 16'd19293, 16'd39145, 16'd875, 16'd50031, 16'd34684, 16'd38215, 16'd39921, 16'd2540});
	test_expansion(128'he42bfc78392af06ab62f220a3c9e5f3d, {16'd28530, 16'd49501, 16'd42873, 16'd24959, 16'd63826, 16'd63259, 16'd51613, 16'd52499, 16'd31083, 16'd31472, 16'd8709, 16'd63086, 16'd29959, 16'd2978, 16'd5641, 16'd12846, 16'd15553, 16'd64080, 16'd24492, 16'd537, 16'd63808, 16'd64255, 16'd43046, 16'd49259, 16'd56424, 16'd3052});
	test_expansion(128'hfbc88ec904fc5dae2987334df0268abe, {16'd34964, 16'd9250, 16'd48088, 16'd23471, 16'd4802, 16'd11025, 16'd56612, 16'd42488, 16'd36322, 16'd33343, 16'd60918, 16'd45028, 16'd59156, 16'd28296, 16'd46095, 16'd11443, 16'd45353, 16'd3276, 16'd43561, 16'd40090, 16'd46253, 16'd9650, 16'd4696, 16'd10673, 16'd30359, 16'd26550});
	test_expansion(128'h47a6717d82a4fe36c02d42384a283cd9, {16'd879, 16'd25121, 16'd45558, 16'd59963, 16'd9522, 16'd34054, 16'd42060, 16'd3922, 16'd40987, 16'd26433, 16'd45225, 16'd6676, 16'd40380, 16'd14770, 16'd46637, 16'd26671, 16'd17710, 16'd49310, 16'd31385, 16'd49844, 16'd46188, 16'd3594, 16'd63562, 16'd15806, 16'd10558, 16'd22673});
	test_expansion(128'h552a14825bf05efee04214ee7dade40b, {16'd34887, 16'd48619, 16'd21431, 16'd26796, 16'd6625, 16'd20497, 16'd22010, 16'd62641, 16'd17795, 16'd51331, 16'd8994, 16'd30613, 16'd47663, 16'd16298, 16'd43132, 16'd26252, 16'd10303, 16'd19951, 16'd9988, 16'd23978, 16'd26108, 16'd31733, 16'd19350, 16'd20919, 16'd58484, 16'd39567});
	test_expansion(128'hc115d85a4ea55066c48947bde1e6a752, {16'd41423, 16'd19564, 16'd30972, 16'd53914, 16'd21875, 16'd61869, 16'd26978, 16'd57728, 16'd37764, 16'd6156, 16'd36252, 16'd24238, 16'd16569, 16'd14729, 16'd51584, 16'd58877, 16'd11300, 16'd46251, 16'd22862, 16'd3189, 16'd52519, 16'd31833, 16'd30617, 16'd29329, 16'd56191, 16'd25833});
	test_expansion(128'h404be6f4ef52ff13b4307624449b9586, {16'd56821, 16'd61228, 16'd10704, 16'd40877, 16'd41092, 16'd17801, 16'd9950, 16'd34787, 16'd54988, 16'd23223, 16'd57383, 16'd45033, 16'd40950, 16'd2685, 16'd58686, 16'd22900, 16'd11003, 16'd7161, 16'd2103, 16'd49233, 16'd1428, 16'd10316, 16'd5663, 16'd4732, 16'd61747, 16'd54490});
	test_expansion(128'h3f875a82a05100fe88fd793612e3be77, {16'd56714, 16'd26657, 16'd61355, 16'd2480, 16'd34554, 16'd62807, 16'd52749, 16'd5875, 16'd56044, 16'd14884, 16'd7038, 16'd50213, 16'd53251, 16'd51449, 16'd60755, 16'd58812, 16'd24157, 16'd48838, 16'd14823, 16'd45371, 16'd59181, 16'd64374, 16'd46245, 16'd47597, 16'd12700, 16'd25957});
	test_expansion(128'he7c9a06e05b45d349e8511eb5584d118, {16'd24009, 16'd9192, 16'd4504, 16'd64094, 16'd65149, 16'd53565, 16'd19859, 16'd44007, 16'd47300, 16'd1590, 16'd30656, 16'd31378, 16'd46085, 16'd64555, 16'd34338, 16'd13330, 16'd38742, 16'd37847, 16'd63725, 16'd24988, 16'd43627, 16'd36488, 16'd17285, 16'd42734, 16'd32331, 16'd64808});
	test_expansion(128'h64cc6089b7e6bd8894ad4f66b9468598, {16'd49847, 16'd8822, 16'd19618, 16'd13444, 16'd30834, 16'd40504, 16'd36365, 16'd21904, 16'd26359, 16'd11636, 16'd47552, 16'd509, 16'd16803, 16'd21526, 16'd61880, 16'd33337, 16'd27726, 16'd52716, 16'd24114, 16'd15878, 16'd10844, 16'd33205, 16'd12674, 16'd3778, 16'd62545, 16'd47166});
	test_expansion(128'h53b77774dd152fdbe2ecd3e4606ff10a, {16'd50497, 16'd22500, 16'd4308, 16'd58760, 16'd44063, 16'd9583, 16'd43973, 16'd28478, 16'd17628, 16'd58149, 16'd33383, 16'd51075, 16'd45581, 16'd57052, 16'd7046, 16'd19342, 16'd14170, 16'd28393, 16'd22796, 16'd22324, 16'd21161, 16'd9061, 16'd63766, 16'd26992, 16'd24529, 16'd37629});
	test_expansion(128'hd45b7a6e3f287caaf97afcb08c3f5991, {16'd12311, 16'd20243, 16'd60064, 16'd41414, 16'd15787, 16'd18217, 16'd25924, 16'd24332, 16'd7754, 16'd4195, 16'd61178, 16'd12022, 16'd12860, 16'd50814, 16'd64953, 16'd47558, 16'd8307, 16'd1352, 16'd8749, 16'd43929, 16'd52073, 16'd8841, 16'd11247, 16'd44236, 16'd3179, 16'd63528});
	test_expansion(128'hbf7e880cee0f5dce1f77716b481d76df, {16'd4222, 16'd26704, 16'd48009, 16'd32426, 16'd18460, 16'd25, 16'd47047, 16'd53950, 16'd15183, 16'd29855, 16'd47770, 16'd6020, 16'd54977, 16'd32208, 16'd28275, 16'd37022, 16'd61568, 16'd43931, 16'd64147, 16'd49300, 16'd35743, 16'd910, 16'd63896, 16'd25243, 16'd39970, 16'd63742});
	test_expansion(128'hc39024c71725a0766b406c1849266973, {16'd45317, 16'd35305, 16'd44303, 16'd22746, 16'd56754, 16'd51980, 16'd30522, 16'd5983, 16'd5163, 16'd21262, 16'd22916, 16'd6582, 16'd48562, 16'd33334, 16'd45797, 16'd30652, 16'd60639, 16'd41140, 16'd47971, 16'd39917, 16'd1707, 16'd11844, 16'd39967, 16'd1079, 16'd26474, 16'd8188});
	test_expansion(128'h6a9f62fbac9c949524f00ce444a73534, {16'd52499, 16'd6150, 16'd47384, 16'd53034, 16'd64692, 16'd51359, 16'd39622, 16'd17985, 16'd64617, 16'd42234, 16'd12789, 16'd8781, 16'd55898, 16'd21649, 16'd34927, 16'd15665, 16'd28543, 16'd53418, 16'd12493, 16'd50302, 16'd28455, 16'd31755, 16'd64876, 16'd55567, 16'd65176, 16'd21970});
	test_expansion(128'h77217e2ae445d6772720de945d3f5c8b, {16'd1165, 16'd10292, 16'd25322, 16'd58494, 16'd41183, 16'd63579, 16'd51338, 16'd60627, 16'd50345, 16'd49799, 16'd12107, 16'd30906, 16'd3929, 16'd53862, 16'd65438, 16'd25198, 16'd23414, 16'd19121, 16'd24682, 16'd40042, 16'd40128, 16'd52683, 16'd17649, 16'd40726, 16'd29958, 16'd10648});
	test_expansion(128'h622b2b7f19d0af3f481b6804ddbebe91, {16'd15829, 16'd51053, 16'd40840, 16'd18185, 16'd53164, 16'd40925, 16'd25919, 16'd5499, 16'd13276, 16'd20826, 16'd42026, 16'd17017, 16'd20339, 16'd37778, 16'd34667, 16'd30748, 16'd60362, 16'd35469, 16'd39740, 16'd53991, 16'd15675, 16'd62495, 16'd18441, 16'd21861, 16'd45468, 16'd26746});
	test_expansion(128'hfaa0e9f7434bf27c33c0e8aa395f3505, {16'd63857, 16'd51807, 16'd14648, 16'd21368, 16'd46189, 16'd27434, 16'd55712, 16'd37904, 16'd16572, 16'd54682, 16'd38192, 16'd13384, 16'd10669, 16'd5252, 16'd45983, 16'd11284, 16'd56951, 16'd49505, 16'd52096, 16'd1198, 16'd5225, 16'd30141, 16'd23191, 16'd12296, 16'd58022, 16'd60316});
	test_expansion(128'h0a498b339d761056d6d83ea98b6c9fba, {16'd65374, 16'd4454, 16'd39682, 16'd29498, 16'd42809, 16'd42019, 16'd11488, 16'd19639, 16'd5647, 16'd252, 16'd40673, 16'd23431, 16'd42390, 16'd23411, 16'd3721, 16'd26796, 16'd22679, 16'd53416, 16'd43547, 16'd17787, 16'd35524, 16'd25770, 16'd58079, 16'd28634, 16'd52912, 16'd63104});
	test_expansion(128'h40b0a4cdf68ec11546977daee17733f7, {16'd45566, 16'd40654, 16'd43265, 16'd43619, 16'd37376, 16'd17253, 16'd63399, 16'd25974, 16'd18743, 16'd26549, 16'd59066, 16'd17198, 16'd1323, 16'd19845, 16'd40767, 16'd63418, 16'd31232, 16'd16945, 16'd44651, 16'd626, 16'd24963, 16'd4761, 16'd62049, 16'd3053, 16'd14517, 16'd58476});
	test_expansion(128'h0ff85b68e87eba6a105ac28dcc0a3ff9, {16'd7571, 16'd3534, 16'd50085, 16'd45907, 16'd46701, 16'd65024, 16'd22230, 16'd21723, 16'd613, 16'd44078, 16'd9060, 16'd26973, 16'd14156, 16'd28241, 16'd24761, 16'd45253, 16'd57371, 16'd43873, 16'd30136, 16'd23370, 16'd51224, 16'd41011, 16'd46629, 16'd62397, 16'd8987, 16'd14878});
	test_expansion(128'h49860de8bfd868f8219ada953215f19e, {16'd51849, 16'd36675, 16'd19910, 16'd62303, 16'd42422, 16'd50484, 16'd16424, 16'd38966, 16'd36752, 16'd48226, 16'd50552, 16'd2867, 16'd43222, 16'd32053, 16'd30482, 16'd55017, 16'd22811, 16'd22138, 16'd15932, 16'd8218, 16'd20287, 16'd63975, 16'd24417, 16'd48078, 16'd33548, 16'd53104});
	test_expansion(128'hb02509346d1193ee16d71cb6baecb039, {16'd41240, 16'd55806, 16'd59720, 16'd25936, 16'd57257, 16'd12901, 16'd52066, 16'd50132, 16'd16575, 16'd802, 16'd41894, 16'd20637, 16'd6536, 16'd62146, 16'd45912, 16'd27831, 16'd51535, 16'd43806, 16'd64785, 16'd16418, 16'd1768, 16'd57444, 16'd32896, 16'd51381, 16'd47721, 16'd46818});
	test_expansion(128'hcc04d3d25962742cd763596481fe480e, {16'd11801, 16'd2627, 16'd55015, 16'd55047, 16'd25503, 16'd14991, 16'd36409, 16'd52318, 16'd14469, 16'd57850, 16'd25768, 16'd48434, 16'd61229, 16'd13661, 16'd31754, 16'd49101, 16'd30854, 16'd54336, 16'd29346, 16'd56879, 16'd7879, 16'd48423, 16'd12823, 16'd29880, 16'd28734, 16'd22065});
	test_expansion(128'h3eb54ebb90da8d8a151c59803d0b8042, {16'd33010, 16'd26454, 16'd49518, 16'd40832, 16'd52405, 16'd64602, 16'd61724, 16'd56061, 16'd56659, 16'd47383, 16'd16161, 16'd16921, 16'd11327, 16'd13464, 16'd42363, 16'd55424, 16'd14671, 16'd47433, 16'd31922, 16'd35325, 16'd55920, 16'd9171, 16'd16107, 16'd37163, 16'd19682, 16'd4658});
	test_expansion(128'h9b0a0d99b9348a0d24a68fb77d31b9b8, {16'd120, 16'd2295, 16'd58567, 16'd41668, 16'd58075, 16'd50159, 16'd53594, 16'd4770, 16'd27394, 16'd12531, 16'd31170, 16'd23684, 16'd44816, 16'd35933, 16'd16406, 16'd11617, 16'd17931, 16'd56972, 16'd53670, 16'd30691, 16'd17583, 16'd23724, 16'd3938, 16'd6906, 16'd11459, 16'd30170});
	test_expansion(128'hca7556840dd5e0df3e9cd87eaa972959, {16'd61612, 16'd22414, 16'd23626, 16'd19139, 16'd32683, 16'd30641, 16'd22070, 16'd32761, 16'd27535, 16'd30560, 16'd31050, 16'd10701, 16'd12335, 16'd57949, 16'd38302, 16'd42254, 16'd38990, 16'd21200, 16'd42265, 16'd61697, 16'd1429, 16'd61437, 16'd42230, 16'd30393, 16'd29468, 16'd7060});
	test_expansion(128'hf0c1dc4d6ff1f72fd0906db0fe454bb5, {16'd58847, 16'd33225, 16'd31927, 16'd6269, 16'd55385, 16'd6326, 16'd61269, 16'd23440, 16'd14023, 16'd51791, 16'd41567, 16'd46159, 16'd20368, 16'd31108, 16'd17602, 16'd49715, 16'd2088, 16'd11629, 16'd15836, 16'd50939, 16'd22630, 16'd51982, 16'd36167, 16'd28590, 16'd55555, 16'd16687});
	test_expansion(128'h02318783380b7b2391636923d2cf6595, {16'd30793, 16'd61323, 16'd59612, 16'd29774, 16'd37915, 16'd8139, 16'd55388, 16'd1928, 16'd41308, 16'd23911, 16'd51384, 16'd11748, 16'd41048, 16'd56936, 16'd53324, 16'd48368, 16'd37338, 16'd41403, 16'd63032, 16'd15881, 16'd792, 16'd22097, 16'd60422, 16'd50641, 16'd27272, 16'd1834});
	test_expansion(128'hb900c9e6078cea3db7c1d37d0678c257, {16'd63257, 16'd62799, 16'd17749, 16'd19354, 16'd24298, 16'd12412, 16'd25958, 16'd58372, 16'd64704, 16'd42806, 16'd36632, 16'd17165, 16'd6563, 16'd48128, 16'd17265, 16'd16590, 16'd24045, 16'd3994, 16'd39630, 16'd55176, 16'd33021, 16'd37662, 16'd34726, 16'd22331, 16'd33750, 16'd52471});
	test_expansion(128'hc3942c6b670bcc2bff0a047a365dd490, {16'd4467, 16'd47489, 16'd49360, 16'd2544, 16'd63624, 16'd24465, 16'd58911, 16'd32383, 16'd47242, 16'd16265, 16'd41150, 16'd35678, 16'd48407, 16'd26522, 16'd261, 16'd29420, 16'd33839, 16'd22744, 16'd22153, 16'd12831, 16'd33380, 16'd40199, 16'd32015, 16'd11856, 16'd1738, 16'd2077});
	test_expansion(128'hf61d53e6ccf9d7d9811ab3034fe343e7, {16'd16376, 16'd21113, 16'd6498, 16'd6950, 16'd12174, 16'd55815, 16'd15669, 16'd53252, 16'd36394, 16'd52454, 16'd46508, 16'd13388, 16'd49911, 16'd20364, 16'd19782, 16'd64735, 16'd12273, 16'd36970, 16'd59760, 16'd10385, 16'd8671, 16'd9873, 16'd53847, 16'd11361, 16'd10276, 16'd6575});
	test_expansion(128'h32b3c2231d5b999071cfa44eee5e7d1e, {16'd59186, 16'd21409, 16'd63862, 16'd14255, 16'd19356, 16'd6294, 16'd25953, 16'd11939, 16'd49096, 16'd32986, 16'd7098, 16'd17416, 16'd54372, 16'd42597, 16'd1306, 16'd62028, 16'd36788, 16'd14152, 16'd46252, 16'd23236, 16'd177, 16'd43743, 16'd43480, 16'd21733, 16'd3028, 16'd2098});
	test_expansion(128'h042fad58c1c1e725252548c696709ae5, {16'd30224, 16'd4549, 16'd34133, 16'd45452, 16'd11251, 16'd54556, 16'd16999, 16'd50135, 16'd51399, 16'd2263, 16'd16019, 16'd56911, 16'd19248, 16'd4101, 16'd60485, 16'd83, 16'd64124, 16'd56100, 16'd22679, 16'd3269, 16'd59970, 16'd27948, 16'd65190, 16'd36660, 16'd12305, 16'd38826});
	test_expansion(128'hc51c300d2549a3b9854df633b8a6bbf1, {16'd39060, 16'd58291, 16'd26806, 16'd46777, 16'd2894, 16'd52533, 16'd24455, 16'd21158, 16'd55061, 16'd22171, 16'd47998, 16'd62912, 16'd729, 16'd36089, 16'd23020, 16'd9240, 16'd49944, 16'd59331, 16'd48395, 16'd63317, 16'd54788, 16'd12295, 16'd43856, 16'd40810, 16'd29387, 16'd40738});
	test_expansion(128'hb493d504d630d68f6e13837f718462e0, {16'd1069, 16'd6598, 16'd3631, 16'd60085, 16'd17137, 16'd64738, 16'd3520, 16'd60855, 16'd50626, 16'd35348, 16'd23466, 16'd23178, 16'd43214, 16'd11305, 16'd47513, 16'd5712, 16'd9946, 16'd9459, 16'd23450, 16'd59266, 16'd20182, 16'd55599, 16'd54633, 16'd17084, 16'd19307, 16'd43433});
	test_expansion(128'hce7a0d429b598f875546def6314185c2, {16'd42470, 16'd60175, 16'd9218, 16'd46450, 16'd47236, 16'd60432, 16'd42425, 16'd54600, 16'd12113, 16'd12747, 16'd55145, 16'd52696, 16'd3028, 16'd5495, 16'd24534, 16'd61480, 16'd3138, 16'd43936, 16'd56048, 16'd40588, 16'd48332, 16'd56613, 16'd36736, 16'd28619, 16'd31897, 16'd29504});
	test_expansion(128'h5d0f6d6a05e2a53d7e2484f990402668, {16'd6906, 16'd20419, 16'd28452, 16'd38032, 16'd21102, 16'd61173, 16'd41944, 16'd4549, 16'd1248, 16'd43668, 16'd51715, 16'd35624, 16'd18146, 16'd23336, 16'd35154, 16'd36831, 16'd15382, 16'd28793, 16'd45151, 16'd30913, 16'd3084, 16'd26590, 16'd52703, 16'd46214, 16'd44707, 16'd16408});
	test_expansion(128'h9414bbd93af0dec342e1b076d4e4d516, {16'd32804, 16'd27783, 16'd39072, 16'd7990, 16'd30702, 16'd43186, 16'd31334, 16'd65128, 16'd32582, 16'd22009, 16'd43845, 16'd22209, 16'd33245, 16'd11692, 16'd8851, 16'd47705, 16'd57564, 16'd6457, 16'd61744, 16'd65369, 16'd26790, 16'd51171, 16'd58977, 16'd26866, 16'd42447, 16'd35694});
	test_expansion(128'h6fc4d883f19519112576f5467f6e29f7, {16'd32629, 16'd48690, 16'd49745, 16'd52428, 16'd23805, 16'd22112, 16'd39018, 16'd36991, 16'd33318, 16'd62124, 16'd48408, 16'd59278, 16'd37925, 16'd9751, 16'd20547, 16'd5055, 16'd20198, 16'd7671, 16'd2328, 16'd18351, 16'd48969, 16'd29838, 16'd55631, 16'd3633, 16'd16951, 16'd23263});
	test_expansion(128'h490969a43775a61078311cb2d0b20d3c, {16'd51060, 16'd52086, 16'd14610, 16'd2466, 16'd25503, 16'd31529, 16'd24885, 16'd10017, 16'd17195, 16'd50050, 16'd9368, 16'd41596, 16'd15962, 16'd4489, 16'd20026, 16'd56738, 16'd21160, 16'd4997, 16'd9624, 16'd15297, 16'd64342, 16'd19214, 16'd3359, 16'd38358, 16'd26630, 16'd65018});
	test_expansion(128'h55cfc5bf1be8621d9b15436da74203d1, {16'd55240, 16'd27720, 16'd58662, 16'd24152, 16'd63556, 16'd37234, 16'd26113, 16'd34761, 16'd35605, 16'd31030, 16'd64597, 16'd28170, 16'd61668, 16'd26049, 16'd5665, 16'd41719, 16'd24266, 16'd58656, 16'd32, 16'd65066, 16'd58341, 16'd51748, 16'd9011, 16'd9137, 16'd31716, 16'd4528});
	test_expansion(128'hbb11be9dd882c0800fe079db92631f4e, {16'd47474, 16'd2900, 16'd47221, 16'd25900, 16'd9504, 16'd6402, 16'd1930, 16'd37509, 16'd9389, 16'd61076, 16'd33870, 16'd33441, 16'd1440, 16'd19215, 16'd34717, 16'd2584, 16'd34472, 16'd2692, 16'd26685, 16'd35583, 16'd9068, 16'd57611, 16'd48924, 16'd14969, 16'd61077, 16'd29954});
	test_expansion(128'hc63710d955a323f9c252317911404807, {16'd2924, 16'd43955, 16'd15928, 16'd3201, 16'd38557, 16'd39291, 16'd21508, 16'd5510, 16'd62773, 16'd14865, 16'd29727, 16'd9868, 16'd3700, 16'd38659, 16'd12204, 16'd32149, 16'd19505, 16'd52694, 16'd1238, 16'd34574, 16'd49456, 16'd2814, 16'd23965, 16'd17277, 16'd26241, 16'd17426});
	test_expansion(128'h2c489579c6a2278b1d3ddcefa570686c, {16'd6727, 16'd6238, 16'd22175, 16'd57717, 16'd15292, 16'd24552, 16'd61450, 16'd59598, 16'd16077, 16'd18139, 16'd47127, 16'd31832, 16'd55768, 16'd22238, 16'd35369, 16'd33543, 16'd39046, 16'd60665, 16'd20822, 16'd43409, 16'd55343, 16'd21565, 16'd45282, 16'd13459, 16'd63398, 16'd19517});
	test_expansion(128'ha57add9c933a71a6fc6b5e2039f4065d, {16'd62948, 16'd39922, 16'd1008, 16'd38010, 16'd12647, 16'd8228, 16'd40364, 16'd39859, 16'd52430, 16'd45587, 16'd13914, 16'd14232, 16'd12129, 16'd51595, 16'd43963, 16'd62683, 16'd47776, 16'd4853, 16'd4655, 16'd2848, 16'd58410, 16'd40589, 16'd28163, 16'd55043, 16'd25544, 16'd65452});
	test_expansion(128'h1b18fdf8b26cda896f625a45be4a9ad5, {16'd34096, 16'd50539, 16'd58019, 16'd36395, 16'd2857, 16'd10739, 16'd64178, 16'd26729, 16'd37449, 16'd7402, 16'd18621, 16'd24626, 16'd31025, 16'd8989, 16'd19645, 16'd10174, 16'd51984, 16'd51399, 16'd11410, 16'd29237, 16'd8151, 16'd16492, 16'd6487, 16'd10344, 16'd41580, 16'd29784});
	test_expansion(128'hdb30f50029b7608e0586c6984c2d6906, {16'd37292, 16'd56684, 16'd7936, 16'd47417, 16'd41458, 16'd51002, 16'd33790, 16'd27653, 16'd41192, 16'd39702, 16'd6212, 16'd24441, 16'd54515, 16'd39298, 16'd19006, 16'd24926, 16'd16851, 16'd59457, 16'd51722, 16'd65483, 16'd62354, 16'd19248, 16'd55092, 16'd34530, 16'd65418, 16'd25733});
	test_expansion(128'hd61bf20382737b784b85c746c11421b6, {16'd10576, 16'd37336, 16'd64687, 16'd1572, 16'd46048, 16'd38441, 16'd13664, 16'd32966, 16'd18839, 16'd24623, 16'd60672, 16'd35664, 16'd47972, 16'd26231, 16'd51681, 16'd6792, 16'd50485, 16'd17548, 16'd8306, 16'd64744, 16'd28510, 16'd28425, 16'd40291, 16'd14364, 16'd31758, 16'd10571});
	test_expansion(128'hce1f18d699a8cd6d26d60ff484d80bcf, {16'd42737, 16'd34879, 16'd50666, 16'd27119, 16'd56478, 16'd62868, 16'd48140, 16'd9545, 16'd31890, 16'd17710, 16'd31587, 16'd49576, 16'd6710, 16'd28510, 16'd12611, 16'd62193, 16'd19444, 16'd9676, 16'd52369, 16'd34512, 16'd3082, 16'd24136, 16'd717, 16'd21976, 16'd2525, 16'd27508});
	test_expansion(128'h0ebd559a6860d9ccbb4104565f8ba62b, {16'd59728, 16'd54142, 16'd55224, 16'd22386, 16'd6533, 16'd5399, 16'd42491, 16'd19494, 16'd59115, 16'd15012, 16'd50799, 16'd37934, 16'd16559, 16'd21334, 16'd57932, 16'd17723, 16'd19042, 16'd62242, 16'd21709, 16'd21026, 16'd58565, 16'd50038, 16'd10936, 16'd10241, 16'd42269, 16'd30797});
	test_expansion(128'h879b046a0ef1ddba29b3f742e1ea8c6f, {16'd35865, 16'd16185, 16'd54710, 16'd38400, 16'd19375, 16'd30809, 16'd36387, 16'd50218, 16'd47231, 16'd1324, 16'd24147, 16'd39534, 16'd61445, 16'd63463, 16'd46952, 16'd60718, 16'd33432, 16'd61627, 16'd53352, 16'd56804, 16'd60914, 16'd32464, 16'd32697, 16'd57248, 16'd29851, 16'd55154});
	test_expansion(128'hb304dfb1c59d33d8020095b06aeb1790, {16'd59973, 16'd12648, 16'd38125, 16'd19865, 16'd60390, 16'd10060, 16'd42171, 16'd58273, 16'd46043, 16'd28701, 16'd22798, 16'd8484, 16'd36856, 16'd1862, 16'd30255, 16'd42740, 16'd1536, 16'd9233, 16'd17316, 16'd41457, 16'd49239, 16'd13195, 16'd10503, 16'd32923, 16'd41475, 16'd12468});
	test_expansion(128'h9fb783b5f42d19575ec95296e599eb8e, {16'd59177, 16'd456, 16'd34532, 16'd44947, 16'd28498, 16'd20222, 16'd12645, 16'd16444, 16'd6259, 16'd32073, 16'd54798, 16'd20290, 16'd17503, 16'd52648, 16'd32377, 16'd37744, 16'd32099, 16'd34497, 16'd1235, 16'd62127, 16'd64007, 16'd30310, 16'd29447, 16'd61605, 16'd31609, 16'd37143});
	test_expansion(128'h2644d31358cf6bd791dcc376d5e76850, {16'd12716, 16'd40390, 16'd7726, 16'd62980, 16'd8034, 16'd30554, 16'd6199, 16'd20012, 16'd7619, 16'd59533, 16'd22082, 16'd27656, 16'd25037, 16'd18583, 16'd2692, 16'd27458, 16'd24176, 16'd39571, 16'd52455, 16'd33159, 16'd37877, 16'd50468, 16'd6656, 16'd12148, 16'd44171, 16'd7035});
	test_expansion(128'hdde7859e623a35571ea5060469eac205, {16'd2324, 16'd4744, 16'd23435, 16'd27127, 16'd47610, 16'd17075, 16'd33590, 16'd25887, 16'd65408, 16'd27464, 16'd53389, 16'd30505, 16'd15013, 16'd55766, 16'd12806, 16'd47289, 16'd35808, 16'd6265, 16'd34438, 16'd38977, 16'd12741, 16'd62381, 16'd25071, 16'd16775, 16'd9434, 16'd24633});
	test_expansion(128'h0326f5269214db45304c1ba8a1b1e1cb, {16'd29874, 16'd18436, 16'd26746, 16'd23610, 16'd27102, 16'd55119, 16'd3617, 16'd44618, 16'd13112, 16'd2563, 16'd5871, 16'd44910, 16'd38276, 16'd7738, 16'd7379, 16'd60233, 16'd17527, 16'd62063, 16'd58865, 16'd38933, 16'd15016, 16'd41182, 16'd55617, 16'd56753, 16'd51875, 16'd35991});
	test_expansion(128'ha8bfa7b51ca046302bb8c285a7f3eb81, {16'd52663, 16'd43217, 16'd54859, 16'd11128, 16'd39498, 16'd57418, 16'd8229, 16'd45950, 16'd7783, 16'd36440, 16'd7092, 16'd53430, 16'd227, 16'd12278, 16'd55904, 16'd34166, 16'd58329, 16'd52992, 16'd56312, 16'd7604, 16'd3501, 16'd10218, 16'd43122, 16'd11723, 16'd15402, 16'd28914});
	test_expansion(128'h8a02d096afa1b50c5926febcabad5809, {16'd60313, 16'd64476, 16'd3111, 16'd48065, 16'd55435, 16'd56290, 16'd916, 16'd23848, 16'd33518, 16'd52563, 16'd32084, 16'd12832, 16'd24952, 16'd20565, 16'd60708, 16'd26498, 16'd4583, 16'd23522, 16'd62570, 16'd28090, 16'd46498, 16'd4752, 16'd54426, 16'd61959, 16'd32137, 16'd62538});
	test_expansion(128'h61bcddae3235aa90e0d556b4231c55a5, {16'd54626, 16'd634, 16'd708, 16'd28788, 16'd18822, 16'd58574, 16'd64546, 16'd48966, 16'd6131, 16'd63577, 16'd25333, 16'd45313, 16'd12372, 16'd57178, 16'd52243, 16'd65026, 16'd57669, 16'd8111, 16'd62103, 16'd44423, 16'd35550, 16'd9062, 16'd50672, 16'd32321, 16'd5032, 16'd34470});
	test_expansion(128'h5ca4621ebb363ceebf0569e8d73c54bf, {16'd25098, 16'd59923, 16'd40246, 16'd26176, 16'd16231, 16'd53914, 16'd64157, 16'd14171, 16'd10953, 16'd28738, 16'd19647, 16'd15618, 16'd34110, 16'd12321, 16'd20403, 16'd32123, 16'd32239, 16'd33534, 16'd29224, 16'd32527, 16'd23641, 16'd44291, 16'd60774, 16'd14920, 16'd52702, 16'd35031});
	test_expansion(128'h78bc0a22f6c8313db5092835f43b7a12, {16'd50111, 16'd26612, 16'd53431, 16'd12594, 16'd53746, 16'd43307, 16'd32105, 16'd17324, 16'd3238, 16'd14135, 16'd39673, 16'd51887, 16'd16401, 16'd17075, 16'd57282, 16'd30974, 16'd47928, 16'd41207, 16'd14582, 16'd49355, 16'd27027, 16'd19739, 16'd4227, 16'd22673, 16'd26395, 16'd3644});
	test_expansion(128'h351edf28bd1f17cb13cd5f26c5130944, {16'd21986, 16'd22580, 16'd51735, 16'd22400, 16'd48392, 16'd31518, 16'd64650, 16'd12380, 16'd42358, 16'd62048, 16'd63700, 16'd30092, 16'd48138, 16'd6318, 16'd64006, 16'd39063, 16'd2548, 16'd42161, 16'd63364, 16'd40601, 16'd2258, 16'd40885, 16'd40100, 16'd52392, 16'd4111, 16'd9245});
	test_expansion(128'h1a5af0aa99e3c791c469635880ac33e0, {16'd25513, 16'd24906, 16'd25101, 16'd35443, 16'd52118, 16'd34651, 16'd1478, 16'd64209, 16'd10558, 16'd65468, 16'd25727, 16'd37809, 16'd21635, 16'd27686, 16'd31812, 16'd54432, 16'd54225, 16'd26240, 16'd21139, 16'd887, 16'd21493, 16'd33256, 16'd7375, 16'd12986, 16'd515, 16'd1327});
	test_expansion(128'h62737898566981f2a36c75e6a21c502a, {16'd8219, 16'd47790, 16'd52407, 16'd19883, 16'd31099, 16'd33258, 16'd35434, 16'd43551, 16'd6882, 16'd21071, 16'd50620, 16'd63083, 16'd7541, 16'd23542, 16'd19306, 16'd54155, 16'd33858, 16'd4719, 16'd8518, 16'd14539, 16'd9532, 16'd48641, 16'd31289, 16'd53456, 16'd42306, 16'd29578});
	test_expansion(128'h0045ff043698263d15bd0849bd239c9e, {16'd36527, 16'd15607, 16'd42570, 16'd9317, 16'd61185, 16'd61246, 16'd57804, 16'd42168, 16'd4927, 16'd42829, 16'd17678, 16'd16995, 16'd58295, 16'd45450, 16'd55024, 16'd23999, 16'd35486, 16'd28691, 16'd58130, 16'd23456, 16'd11953, 16'd7438, 16'd37462, 16'd3954, 16'd29780, 16'd54666});
	test_expansion(128'hb50c7c1f1f941b0b787c49123a2b7cc8, {16'd5151, 16'd26861, 16'd41367, 16'd33612, 16'd21979, 16'd29459, 16'd16366, 16'd19900, 16'd4301, 16'd53563, 16'd52791, 16'd38927, 16'd7103, 16'd42249, 16'd2411, 16'd14938, 16'd19379, 16'd19408, 16'd7603, 16'd23756, 16'd42772, 16'd33253, 16'd28515, 16'd9700, 16'd33150, 16'd48032});
	test_expansion(128'he274cc7a9bf5c1d7d5caa8028f86ab42, {16'd62306, 16'd29512, 16'd25630, 16'd9779, 16'd28431, 16'd53713, 16'd4727, 16'd61221, 16'd46415, 16'd20146, 16'd51468, 16'd48835, 16'd14894, 16'd18552, 16'd48088, 16'd53198, 16'd33707, 16'd30349, 16'd9100, 16'd22147, 16'd53003, 16'd2595, 16'd19201, 16'd34246, 16'd45460, 16'd54412});
	test_expansion(128'h0ff3349c701559d6f7690886068a690b, {16'd27555, 16'd22366, 16'd2026, 16'd20105, 16'd12683, 16'd6825, 16'd39040, 16'd43149, 16'd32380, 16'd16074, 16'd37307, 16'd51272, 16'd41278, 16'd4008, 16'd36267, 16'd52924, 16'd20099, 16'd25249, 16'd51289, 16'd65523, 16'd60282, 16'd53482, 16'd51327, 16'd26859, 16'd48748, 16'd6987});
	test_expansion(128'he128daea475b2571510043f4f9c2f235, {16'd4688, 16'd28844, 16'd16514, 16'd6665, 16'd11662, 16'd20122, 16'd3978, 16'd39231, 16'd17425, 16'd6446, 16'd3278, 16'd16407, 16'd21099, 16'd45288, 16'd28102, 16'd33980, 16'd63388, 16'd57248, 16'd22082, 16'd40604, 16'd11267, 16'd42586, 16'd48919, 16'd60747, 16'd15173, 16'd10518});
	test_expansion(128'ha6f09f2e83f0ed30f8f93b1fec50ef1b, {16'd55532, 16'd28781, 16'd64652, 16'd44466, 16'd21398, 16'd64004, 16'd54619, 16'd17797, 16'd29751, 16'd43748, 16'd34179, 16'd36786, 16'd42682, 16'd31063, 16'd14061, 16'd25183, 16'd31248, 16'd62951, 16'd15520, 16'd48763, 16'd13990, 16'd36916, 16'd40857, 16'd51001, 16'd28828, 16'd65429});
	test_expansion(128'h63ff4f56eae158036a42f347c87f00e2, {16'd37062, 16'd22478, 16'd31895, 16'd64330, 16'd5202, 16'd47580, 16'd25556, 16'd53773, 16'd8806, 16'd5720, 16'd52644, 16'd15108, 16'd55295, 16'd23382, 16'd37231, 16'd52850, 16'd21870, 16'd18720, 16'd8115, 16'd50525, 16'd57763, 16'd7867, 16'd52898, 16'd41053, 16'd22145, 16'd37378});
	test_expansion(128'h5df0231283d3dd7440c795262d39b426, {16'd36172, 16'd37172, 16'd53077, 16'd30293, 16'd52357, 16'd36404, 16'd25072, 16'd55895, 16'd13999, 16'd58546, 16'd9201, 16'd40872, 16'd47998, 16'd16122, 16'd473, 16'd3760, 16'd2682, 16'd52637, 16'd38063, 16'd30589, 16'd33611, 16'd49951, 16'd33659, 16'd43111, 16'd22290, 16'd57404});
	test_expansion(128'h90316d0d41e19c636a63eb4555cd65a4, {16'd277, 16'd33788, 16'd36415, 16'd36512, 16'd33943, 16'd60173, 16'd831, 16'd25975, 16'd59873, 16'd50860, 16'd37184, 16'd7846, 16'd52014, 16'd41327, 16'd34953, 16'd28097, 16'd58524, 16'd46577, 16'd43984, 16'd31191, 16'd6032, 16'd4188, 16'd63920, 16'd49169, 16'd55928, 16'd1024});
	test_expansion(128'h787f56722725b9b3380e83b0add30925, {16'd18184, 16'd16571, 16'd48437, 16'd19236, 16'd5304, 16'd62269, 16'd4371, 16'd1234, 16'd57499, 16'd62478, 16'd7260, 16'd39437, 16'd5050, 16'd40495, 16'd20123, 16'd19957, 16'd56111, 16'd28223, 16'd15310, 16'd3170, 16'd22274, 16'd8971, 16'd23072, 16'd35087, 16'd17460, 16'd29332});
	test_expansion(128'h2752c4bae26e8f4bbcd5817eccbdbd0a, {16'd12225, 16'd57593, 16'd49360, 16'd2570, 16'd2013, 16'd42432, 16'd9414, 16'd49603, 16'd41792, 16'd54735, 16'd57820, 16'd12786, 16'd47161, 16'd15669, 16'd52761, 16'd38356, 16'd44377, 16'd2666, 16'd18314, 16'd21985, 16'd8082, 16'd32929, 16'd37353, 16'd60186, 16'd39443, 16'd61650});
	test_expansion(128'he100f893c52dcccc682c48f12bc6d01f, {16'd25800, 16'd28980, 16'd11967, 16'd1202, 16'd7941, 16'd63205, 16'd40520, 16'd27246, 16'd39275, 16'd57083, 16'd13420, 16'd37377, 16'd61511, 16'd32159, 16'd60003, 16'd12388, 16'd17486, 16'd31137, 16'd12557, 16'd63972, 16'd57624, 16'd22690, 16'd63757, 16'd34541, 16'd46618, 16'd40818});
	test_expansion(128'h2e3d31d229ee9c698476651d44cf683d, {16'd1698, 16'd58545, 16'd3385, 16'd42390, 16'd52293, 16'd17234, 16'd4233, 16'd58047, 16'd1935, 16'd42851, 16'd61077, 16'd816, 16'd35675, 16'd38138, 16'd40921, 16'd1156, 16'd17322, 16'd59657, 16'd58650, 16'd16498, 16'd24429, 16'd35880, 16'd14509, 16'd421, 16'd887, 16'd43039});
	test_expansion(128'hc9fa86802db7713e0d924ce64e231dbd, {16'd18388, 16'd58820, 16'd1473, 16'd95, 16'd39519, 16'd62987, 16'd40823, 16'd20005, 16'd42922, 16'd42669, 16'd42239, 16'd46680, 16'd29391, 16'd17691, 16'd63173, 16'd36058, 16'd38637, 16'd32979, 16'd15849, 16'd33930, 16'd43838, 16'd31569, 16'd1398, 16'd37043, 16'd2515, 16'd29788});
	test_expansion(128'he85bce3af0212bb409febeaf84910ec5, {16'd9216, 16'd53739, 16'd11215, 16'd1625, 16'd46485, 16'd19447, 16'd5536, 16'd11234, 16'd39413, 16'd42900, 16'd9631, 16'd1948, 16'd28370, 16'd1811, 16'd63487, 16'd28134, 16'd36352, 16'd21611, 16'd54726, 16'd45461, 16'd57224, 16'd8483, 16'd1169, 16'd44507, 16'd623, 16'd55700});
	test_expansion(128'h0ab7b12b908d750058dc764434a72050, {16'd38850, 16'd43086, 16'd6996, 16'd37828, 16'd32073, 16'd6894, 16'd26359, 16'd31798, 16'd61824, 16'd53767, 16'd26897, 16'd56998, 16'd41291, 16'd15199, 16'd38069, 16'd48287, 16'd57844, 16'd20151, 16'd21223, 16'd22280, 16'd30202, 16'd24108, 16'd34590, 16'd12932, 16'd42328, 16'd41899});
	test_expansion(128'h0e33dc71b5ca493eab4801b708d4b5b8, {16'd22093, 16'd43985, 16'd47777, 16'd12958, 16'd46726, 16'd56850, 16'd3059, 16'd22492, 16'd8976, 16'd38241, 16'd148, 16'd14696, 16'd36606, 16'd40049, 16'd35396, 16'd38105, 16'd45693, 16'd62560, 16'd15342, 16'd53894, 16'd11644, 16'd7945, 16'd19495, 16'd8426, 16'd29546, 16'd32164});
	test_expansion(128'h2353736e3ee126acc2c84a514c216977, {16'd7394, 16'd1828, 16'd61332, 16'd43945, 16'd8075, 16'd60601, 16'd7296, 16'd10066, 16'd248, 16'd29565, 16'd25114, 16'd21679, 16'd55841, 16'd21332, 16'd56799, 16'd14574, 16'd29503, 16'd21441, 16'd14743, 16'd18906, 16'd12451, 16'd2422, 16'd46032, 16'd30668, 16'd8600, 16'd36570});
	test_expansion(128'h4b3df853d299cabf2ef21c2bfeb00bbf, {16'd1033, 16'd44361, 16'd46076, 16'd34136, 16'd43775, 16'd28997, 16'd27112, 16'd6118, 16'd62755, 16'd38261, 16'd47631, 16'd6812, 16'd41058, 16'd7922, 16'd11703, 16'd28216, 16'd28665, 16'd61501, 16'd14828, 16'd62313, 16'd64524, 16'd15041, 16'd29808, 16'd16359, 16'd11192, 16'd39661});
	test_expansion(128'h81f53cce8b1e6d661513ef69d50f0acd, {16'd17707, 16'd2015, 16'd42521, 16'd33413, 16'd56157, 16'd59098, 16'd1540, 16'd36753, 16'd63606, 16'd56280, 16'd50457, 16'd11571, 16'd51981, 16'd43880, 16'd17175, 16'd15467, 16'd2223, 16'd17658, 16'd42078, 16'd38734, 16'd2401, 16'd61805, 16'd9330, 16'd35480, 16'd28681, 16'd31532});
	test_expansion(128'h3fa7f7e76c97cce1ece474865973852b, {16'd33725, 16'd38745, 16'd23612, 16'd2263, 16'd23338, 16'd60662, 16'd52109, 16'd34464, 16'd57914, 16'd51741, 16'd19130, 16'd50335, 16'd5604, 16'd50683, 16'd64726, 16'd64186, 16'd54629, 16'd29332, 16'd5544, 16'd26094, 16'd8852, 16'd55808, 16'd12289, 16'd46889, 16'd2650, 16'd40019});
	test_expansion(128'h72e8afa6ee562554e672d6949fa1a21f, {16'd18089, 16'd25326, 16'd41680, 16'd15334, 16'd7158, 16'd51791, 16'd19136, 16'd26979, 16'd39991, 16'd1534, 16'd62279, 16'd30864, 16'd62107, 16'd26828, 16'd16583, 16'd47574, 16'd21661, 16'd17479, 16'd12099, 16'd5592, 16'd20903, 16'd16385, 16'd2989, 16'd44404, 16'd11339, 16'd15803});
	test_expansion(128'h9305ce84dbc29eb4b555a8bbd8e16838, {16'd12111, 16'd37428, 16'd46550, 16'd39988, 16'd34995, 16'd59080, 16'd45904, 16'd63214, 16'd18123, 16'd6258, 16'd35047, 16'd15394, 16'd18771, 16'd33273, 16'd49942, 16'd26605, 16'd56723, 16'd43147, 16'd57242, 16'd5240, 16'd4132, 16'd33789, 16'd61507, 16'd50949, 16'd25517, 16'd38681});
	test_expansion(128'hd7045f7d103bd174718922c1d60f9f89, {16'd49972, 16'd16946, 16'd30647, 16'd63129, 16'd32291, 16'd39102, 16'd30287, 16'd6099, 16'd31428, 16'd35061, 16'd33449, 16'd24958, 16'd19828, 16'd2990, 16'd16020, 16'd60330, 16'd64238, 16'd13735, 16'd12993, 16'd31280, 16'd5999, 16'd24091, 16'd18592, 16'd4415, 16'd62909, 16'd38342});
	test_expansion(128'h60a561d93d00b044cfb8ad26b9d12f64, {16'd36247, 16'd47485, 16'd18175, 16'd55413, 16'd59645, 16'd42365, 16'd23513, 16'd62988, 16'd20776, 16'd56704, 16'd47167, 16'd47426, 16'd2486, 16'd19359, 16'd15350, 16'd15866, 16'd29721, 16'd36125, 16'd49639, 16'd24438, 16'd13559, 16'd54979, 16'd62729, 16'd53623, 16'd63426, 16'd511});
	test_expansion(128'h6c012c071ab468c3038ef3593430f4cc, {16'd18568, 16'd53879, 16'd48700, 16'd60403, 16'd58678, 16'd28394, 16'd43904, 16'd62844, 16'd62464, 16'd11758, 16'd110, 16'd176, 16'd19430, 16'd6219, 16'd34920, 16'd52467, 16'd21537, 16'd42079, 16'd35864, 16'd9545, 16'd41668, 16'd16029, 16'd53221, 16'd12654, 16'd49706, 16'd18619});
	test_expansion(128'h7c6a323cfde25157fa2fc0f95f78c04b, {16'd47314, 16'd14110, 16'd59493, 16'd45645, 16'd28836, 16'd3709, 16'd37106, 16'd5035, 16'd60267, 16'd19012, 16'd33885, 16'd3053, 16'd5922, 16'd38888, 16'd60102, 16'd12969, 16'd31185, 16'd13465, 16'd11268, 16'd7641, 16'd706, 16'd13590, 16'd16451, 16'd41409, 16'd14153, 16'd36677});
	test_expansion(128'h0d6dbc21bdd90d73c5a823f2f36b266e, {16'd37753, 16'd34113, 16'd18905, 16'd50599, 16'd15318, 16'd20746, 16'd40163, 16'd62049, 16'd22302, 16'd47382, 16'd37950, 16'd44793, 16'd6058, 16'd36296, 16'd53279, 16'd65283, 16'd40285, 16'd41511, 16'd38266, 16'd27657, 16'd49127, 16'd23243, 16'd24765, 16'd48239, 16'd52761, 16'd52598});
	test_expansion(128'h9c6aaa9d8060512cb770e1106e16174b, {16'd36385, 16'd27425, 16'd29019, 16'd45627, 16'd36084, 16'd33029, 16'd56324, 16'd24594, 16'd48838, 16'd33962, 16'd28136, 16'd59143, 16'd43686, 16'd6729, 16'd60385, 16'd17628, 16'd57298, 16'd5094, 16'd16948, 16'd45517, 16'd14145, 16'd39330, 16'd60128, 16'd3827, 16'd35888, 16'd38799});
	test_expansion(128'hd6a501f2988c418cf8e0699f54e2cf3c, {16'd5028, 16'd20169, 16'd17737, 16'd25460, 16'd2065, 16'd26575, 16'd34037, 16'd51857, 16'd12186, 16'd24727, 16'd61386, 16'd29646, 16'd5736, 16'd50873, 16'd17870, 16'd57145, 16'd45500, 16'd52499, 16'd41242, 16'd39178, 16'd22731, 16'd2881, 16'd29512, 16'd55138, 16'd55573, 16'd45998});
	test_expansion(128'hd027d6bf7705c4c8c18bf916b7ae56a1, {16'd40752, 16'd48639, 16'd12377, 16'd181, 16'd44677, 16'd14136, 16'd33031, 16'd27623, 16'd35621, 16'd63255, 16'd42738, 16'd65211, 16'd55317, 16'd11147, 16'd42888, 16'd32935, 16'd14380, 16'd36091, 16'd22636, 16'd53936, 16'd43850, 16'd54092, 16'd60556, 16'd10787, 16'd40310, 16'd65418});
	test_expansion(128'h80f1a9fbe32981246041f952ff55cefa, {16'd24390, 16'd33270, 16'd55275, 16'd48520, 16'd16280, 16'd35165, 16'd15424, 16'd32812, 16'd51329, 16'd15156, 16'd56088, 16'd105, 16'd33397, 16'd60674, 16'd46665, 16'd50905, 16'd55023, 16'd31357, 16'd50348, 16'd63592, 16'd59224, 16'd33536, 16'd64361, 16'd35731, 16'd65223, 16'd59771});
	test_expansion(128'h57b44614abb1280c8270ba22280b014f, {16'd35100, 16'd29208, 16'd54252, 16'd17648, 16'd27877, 16'd40707, 16'd41404, 16'd22735, 16'd59690, 16'd55501, 16'd18527, 16'd36481, 16'd19256, 16'd3661, 16'd29181, 16'd3243, 16'd36893, 16'd25144, 16'd50478, 16'd42008, 16'd28146, 16'd47785, 16'd51060, 16'd5052, 16'd948, 16'd5525});
	test_expansion(128'he31b55b327c54ab940d69c03d1d708ca, {16'd46678, 16'd63067, 16'd46395, 16'd9927, 16'd49356, 16'd48597, 16'd64226, 16'd22002, 16'd61625, 16'd14298, 16'd46969, 16'd57020, 16'd23585, 16'd41853, 16'd21172, 16'd26858, 16'd24782, 16'd41251, 16'd28375, 16'd13798, 16'd50286, 16'd6853, 16'd5235, 16'd60271, 16'd20310, 16'd30462});
	test_expansion(128'h820afd587ca69bfc2eb670f289ce0b59, {16'd38767, 16'd27382, 16'd63720, 16'd24206, 16'd50017, 16'd2213, 16'd4591, 16'd17053, 16'd20574, 16'd5571, 16'd4208, 16'd15334, 16'd51165, 16'd32107, 16'd36110, 16'd29308, 16'd59349, 16'd16123, 16'd62978, 16'd13798, 16'd22599, 16'd63640, 16'd14642, 16'd23317, 16'd2642, 16'd12601});
	test_expansion(128'h45f3966edaad92ee37dcb6bb057ce308, {16'd41519, 16'd21973, 16'd36716, 16'd39910, 16'd1783, 16'd58756, 16'd56658, 16'd13063, 16'd48169, 16'd64476, 16'd31392, 16'd24674, 16'd42677, 16'd39495, 16'd48584, 16'd53681, 16'd35249, 16'd9667, 16'd61338, 16'd16837, 16'd50998, 16'd37070, 16'd21113, 16'd16345, 16'd14597, 16'd53510});
	test_expansion(128'h1da919dc7e9f0813e8b17e583a32d5c0, {16'd47678, 16'd16957, 16'd62962, 16'd53793, 16'd63875, 16'd28494, 16'd26836, 16'd46564, 16'd50128, 16'd11767, 16'd65202, 16'd6616, 16'd59640, 16'd48144, 16'd30862, 16'd4908, 16'd60513, 16'd31710, 16'd13656, 16'd39247, 16'd23789, 16'd40810, 16'd27615, 16'd18255, 16'd9659, 16'd53830});
	test_expansion(128'h0b23337841997b38505571f2416fc6af, {16'd63796, 16'd51652, 16'd64464, 16'd38353, 16'd33629, 16'd7457, 16'd51089, 16'd18899, 16'd61321, 16'd24095, 16'd44156, 16'd50680, 16'd44570, 16'd41535, 16'd40210, 16'd6492, 16'd59176, 16'd32904, 16'd23579, 16'd28238, 16'd1343, 16'd8347, 16'd48914, 16'd55470, 16'd9380, 16'd49708});
	test_expansion(128'h16a6c609d970fba4f1440a8bb49d2536, {16'd59396, 16'd12058, 16'd41967, 16'd21111, 16'd763, 16'd13807, 16'd41147, 16'd16288, 16'd13935, 16'd1599, 16'd45205, 16'd20113, 16'd18668, 16'd36082, 16'd49345, 16'd62799, 16'd36905, 16'd32445, 16'd1495, 16'd59738, 16'd10551, 16'd5451, 16'd1870, 16'd59653, 16'd26078, 16'd17298});
	test_expansion(128'h371d1d95551a855956edfaf921faa95b, {16'd55848, 16'd16420, 16'd40319, 16'd42189, 16'd502, 16'd34083, 16'd56978, 16'd11255, 16'd12832, 16'd7122, 16'd42156, 16'd64668, 16'd58989, 16'd28390, 16'd16814, 16'd25263, 16'd44582, 16'd19871, 16'd51142, 16'd27848, 16'd17257, 16'd47468, 16'd32039, 16'd548, 16'd18830, 16'd29741});
	test_expansion(128'he5f896f5c884c6182cfe712887544c45, {16'd33029, 16'd49920, 16'd167, 16'd28506, 16'd26647, 16'd43121, 16'd63902, 16'd49118, 16'd6286, 16'd11807, 16'd20557, 16'd63925, 16'd28748, 16'd40822, 16'd13644, 16'd50876, 16'd22791, 16'd34670, 16'd10262, 16'd64383, 16'd21537, 16'd34734, 16'd57077, 16'd46574, 16'd6747, 16'd11782});
	test_expansion(128'h23ad5f14d49adc43b13d87d21a516bd2, {16'd19570, 16'd62101, 16'd51736, 16'd7217, 16'd22153, 16'd50494, 16'd27256, 16'd19218, 16'd41203, 16'd12631, 16'd4672, 16'd29378, 16'd30030, 16'd7195, 16'd56068, 16'd46218, 16'd36491, 16'd55282, 16'd28494, 16'd47320, 16'd56135, 16'd59905, 16'd48957, 16'd5127, 16'd23451, 16'd57835});
	test_expansion(128'h8f5692bfc3f301d25b01a6fb260290ff, {16'd57905, 16'd51011, 16'd8319, 16'd5677, 16'd19559, 16'd39507, 16'd60677, 16'd47102, 16'd11667, 16'd2058, 16'd42057, 16'd44557, 16'd29813, 16'd28846, 16'd21433, 16'd28617, 16'd45619, 16'd60112, 16'd42633, 16'd23696, 16'd38196, 16'd38785, 16'd57602, 16'd40501, 16'd17617, 16'd50985});
	test_expansion(128'h24d331061e1f03fe7fbb6d583a6cbe04, {16'd61320, 16'd60941, 16'd9264, 16'd57775, 16'd46179, 16'd41846, 16'd8057, 16'd2346, 16'd18319, 16'd30130, 16'd32851, 16'd31778, 16'd39244, 16'd3347, 16'd2183, 16'd10411, 16'd32963, 16'd10206, 16'd25157, 16'd41821, 16'd26257, 16'd18980, 16'd43324, 16'd30978, 16'd7747, 16'd8378});
	test_expansion(128'h9c0338c9c134624ded1898fb1ee9df0c, {16'd1579, 16'd43162, 16'd20978, 16'd13887, 16'd19444, 16'd28267, 16'd31284, 16'd23192, 16'd29145, 16'd18673, 16'd28102, 16'd34747, 16'd8715, 16'd64206, 16'd50590, 16'd15074, 16'd37319, 16'd28911, 16'd42733, 16'd22296, 16'd5218, 16'd41119, 16'd17879, 16'd52396, 16'd10028, 16'd51810});
	test_expansion(128'hd3db9517bc0b53eb9a1aa4bed1b233d4, {16'd36314, 16'd988, 16'd49286, 16'd43535, 16'd4255, 16'd11422, 16'd48250, 16'd48689, 16'd24235, 16'd21044, 16'd57692, 16'd14308, 16'd50454, 16'd35354, 16'd10074, 16'd20521, 16'd2640, 16'd2348, 16'd1037, 16'd49071, 16'd27244, 16'd48210, 16'd22913, 16'd38050, 16'd46234, 16'd61961});
	test_expansion(128'hb5aed7b6e73f069c13838ef26fdb2614, {16'd5946, 16'd56077, 16'd20624, 16'd29887, 16'd31212, 16'd25642, 16'd33594, 16'd5832, 16'd2892, 16'd48359, 16'd57530, 16'd5208, 16'd30281, 16'd64829, 16'd9366, 16'd47419, 16'd43771, 16'd48343, 16'd36630, 16'd29455, 16'd8149, 16'd24122, 16'd59495, 16'd56355, 16'd30066, 16'd45359});
	test_expansion(128'h83b2a55129bcbe5a4bde8ed7847f10e4, {16'd19695, 16'd45138, 16'd37680, 16'd3165, 16'd50571, 16'd32096, 16'd22737, 16'd35335, 16'd6981, 16'd942, 16'd28073, 16'd40188, 16'd43012, 16'd58503, 16'd47724, 16'd1033, 16'd52509, 16'd14685, 16'd10363, 16'd61483, 16'd55958, 16'd13282, 16'd13250, 16'd18107, 16'd20276, 16'd31289});
	test_expansion(128'hbb9eec35876010ea1c29225d99e632a4, {16'd32682, 16'd57481, 16'd51641, 16'd41646, 16'd51327, 16'd16192, 16'd5998, 16'd46670, 16'd54637, 16'd589, 16'd3893, 16'd34699, 16'd27064, 16'd58405, 16'd50693, 16'd34564, 16'd34338, 16'd20161, 16'd10529, 16'd25503, 16'd64419, 16'd43022, 16'd60116, 16'd28593, 16'd23290, 16'd43166});
	test_expansion(128'h2bdfea259458185ab555ff68992eb68a, {16'd38709, 16'd65529, 16'd674, 16'd12022, 16'd62231, 16'd13242, 16'd56895, 16'd14839, 16'd5087, 16'd4434, 16'd58702, 16'd1410, 16'd41594, 16'd35142, 16'd32217, 16'd18073, 16'd13758, 16'd29715, 16'd26502, 16'd30760, 16'd50819, 16'd54538, 16'd1660, 16'd55631, 16'd47535, 16'd5147});
	test_expansion(128'h3c39597269fde0cc1ec5fe5f9b3928e2, {16'd53371, 16'd47484, 16'd13096, 16'd47538, 16'd39597, 16'd2021, 16'd24165, 16'd31089, 16'd27453, 16'd33449, 16'd45162, 16'd35288, 16'd37845, 16'd61738, 16'd40396, 16'd10525, 16'd13018, 16'd21568, 16'd5636, 16'd18911, 16'd12359, 16'd50569, 16'd45142, 16'd38329, 16'd59183, 16'd31941});
	test_expansion(128'h291cf0ebb7d8625698b12ea2cc95fbc7, {16'd24540, 16'd514, 16'd41994, 16'd41221, 16'd47664, 16'd33739, 16'd51965, 16'd27439, 16'd35818, 16'd40123, 16'd5227, 16'd60216, 16'd19637, 16'd30702, 16'd151, 16'd51186, 16'd43636, 16'd26570, 16'd23601, 16'd2777, 16'd3043, 16'd51572, 16'd52764, 16'd27582, 16'd4676, 16'd50857});
	test_expansion(128'h7b673bebfea82ae1212ba791c553af45, {16'd22366, 16'd15945, 16'd15264, 16'd32140, 16'd57230, 16'd9476, 16'd6775, 16'd9178, 16'd62309, 16'd7026, 16'd63083, 16'd19033, 16'd8414, 16'd40790, 16'd56664, 16'd42186, 16'd51162, 16'd57977, 16'd28, 16'd42912, 16'd43748, 16'd59406, 16'd26406, 16'd15636, 16'd58782, 16'd9361});
	test_expansion(128'h8b00385ea90407f5ed23a42cf3ec7d88, {16'd48218, 16'd40170, 16'd48888, 16'd50889, 16'd18114, 16'd3972, 16'd65119, 16'd54499, 16'd42210, 16'd59335, 16'd15555, 16'd15644, 16'd1581, 16'd12972, 16'd61418, 16'd14543, 16'd39794, 16'd52013, 16'd43697, 16'd23348, 16'd5190, 16'd41094, 16'd22398, 16'd14459, 16'd40740, 16'd17660});
	test_expansion(128'heba4377ac10dba0e4cdf08e74800b87d, {16'd36367, 16'd61139, 16'd9856, 16'd41412, 16'd64717, 16'd21383, 16'd28673, 16'd3289, 16'd25772, 16'd6748, 16'd63560, 16'd8274, 16'd46179, 16'd33584, 16'd26889, 16'd44560, 16'd25059, 16'd64355, 16'd40122, 16'd62383, 16'd3766, 16'd43234, 16'd9646, 16'd44824, 16'd27064, 16'd678});
	test_expansion(128'hc98ec5d9145d1ce32a383285a451bf08, {16'd4185, 16'd28585, 16'd20459, 16'd18850, 16'd18671, 16'd12413, 16'd54945, 16'd12498, 16'd25660, 16'd33383, 16'd3422, 16'd43367, 16'd4539, 16'd11670, 16'd45460, 16'd9245, 16'd51941, 16'd39463, 16'd54354, 16'd4740, 16'd686, 16'd50412, 16'd64174, 16'd8012, 16'd45435, 16'd32951});
	test_expansion(128'h88859a87d88e4b1e03d139c385eac261, {16'd12634, 16'd57004, 16'd51883, 16'd9619, 16'd28692, 16'd33811, 16'd38191, 16'd2322, 16'd15284, 16'd44937, 16'd59018, 16'd55544, 16'd53694, 16'd44112, 16'd9749, 16'd32248, 16'd59682, 16'd37302, 16'd21888, 16'd31609, 16'd16464, 16'd18043, 16'd56669, 16'd5808, 16'd53793, 16'd15920});
	test_expansion(128'h9ff1b54c93358571f5cd5697830dd2a9, {16'd56745, 16'd19219, 16'd10065, 16'd24755, 16'd39681, 16'd47830, 16'd33645, 16'd25016, 16'd57406, 16'd64582, 16'd40475, 16'd1604, 16'd24244, 16'd50912, 16'd29031, 16'd37483, 16'd34426, 16'd28401, 16'd35819, 16'd46544, 16'd11175, 16'd53257, 16'd27357, 16'd42298, 16'd59656, 16'd17151});
	test_expansion(128'h49f2851e871866d99d773a408f7122cd, {16'd20900, 16'd52251, 16'd37095, 16'd45266, 16'd56541, 16'd58176, 16'd58206, 16'd27009, 16'd11645, 16'd19422, 16'd24768, 16'd61752, 16'd1040, 16'd47927, 16'd1249, 16'd62537, 16'd35645, 16'd22308, 16'd30743, 16'd65533, 16'd36165, 16'd33621, 16'd32229, 16'd1711, 16'd46159, 16'd28259});
	test_expansion(128'hd2c7d9af1040af02ee7bb81eeed61a80, {16'd13484, 16'd7826, 16'd31150, 16'd16182, 16'd17192, 16'd42448, 16'd46850, 16'd62299, 16'd42989, 16'd11732, 16'd17349, 16'd31685, 16'd11114, 16'd60500, 16'd52482, 16'd37482, 16'd48070, 16'd22414, 16'd58306, 16'd51877, 16'd2148, 16'd45504, 16'd58821, 16'd10112, 16'd48724, 16'd49765});
	test_expansion(128'hef0f95a9ae8d2a50174c47d23cfc38f9, {16'd7582, 16'd41096, 16'd317, 16'd39931, 16'd38813, 16'd63774, 16'd51659, 16'd65347, 16'd13994, 16'd58998, 16'd2027, 16'd45227, 16'd30190, 16'd64294, 16'd60227, 16'd44223, 16'd60927, 16'd4309, 16'd1872, 16'd52800, 16'd7229, 16'd37562, 16'd59963, 16'd11168, 16'd27196, 16'd7673});
	test_expansion(128'h7fd6072c04574306453ddcdcbcd651cb, {16'd55351, 16'd56736, 16'd24533, 16'd32763, 16'd9475, 16'd62019, 16'd62933, 16'd4303, 16'd24650, 16'd52073, 16'd50307, 16'd11051, 16'd43249, 16'd62884, 16'd39188, 16'd15767, 16'd53949, 16'd50432, 16'd32226, 16'd42665, 16'd20906, 16'd12812, 16'd39847, 16'd35822, 16'd18309, 16'd50966});
	test_expansion(128'h0108cccda755ff4d608b28a2822038dd, {16'd56099, 16'd45176, 16'd44520, 16'd19284, 16'd43419, 16'd52302, 16'd65100, 16'd12852, 16'd3262, 16'd46653, 16'd60653, 16'd31441, 16'd56123, 16'd42023, 16'd39067, 16'd21012, 16'd57076, 16'd19325, 16'd3389, 16'd20715, 16'd63819, 16'd413, 16'd35358, 16'd59202, 16'd30360, 16'd20010});
	test_expansion(128'h195bdf12ef95f21b480e1d88eb719159, {16'd24497, 16'd30536, 16'd64315, 16'd39859, 16'd51812, 16'd50451, 16'd22057, 16'd29697, 16'd23671, 16'd41090, 16'd22067, 16'd45950, 16'd44191, 16'd53852, 16'd45053, 16'd14749, 16'd45125, 16'd56250, 16'd699, 16'd3550, 16'd63936, 16'd33539, 16'd13921, 16'd17354, 16'd15028, 16'd50174});
	test_expansion(128'ha6b70606337a843305a3a50a27dc58ab, {16'd40444, 16'd43606, 16'd44086, 16'd33868, 16'd64130, 16'd58400, 16'd22174, 16'd4189, 16'd31609, 16'd60488, 16'd14978, 16'd2930, 16'd2542, 16'd18982, 16'd28520, 16'd57485, 16'd35577, 16'd10678, 16'd13589, 16'd54886, 16'd2640, 16'd17828, 16'd1850, 16'd28735, 16'd240, 16'd59820});
	test_expansion(128'h77ce1201d1ce8f3e92f624279ea676dc, {16'd49029, 16'd37683, 16'd45515, 16'd43224, 16'd56598, 16'd51790, 16'd62317, 16'd1697, 16'd29527, 16'd34678, 16'd48958, 16'd18459, 16'd62897, 16'd64889, 16'd17450, 16'd2122, 16'd11596, 16'd25162, 16'd52153, 16'd31795, 16'd35275, 16'd742, 16'd59222, 16'd15872, 16'd7670, 16'd28957});
	test_expansion(128'hd77e2f40e0c725b3e27e107a0223cd89, {16'd63335, 16'd19882, 16'd33276, 16'd35140, 16'd41022, 16'd23637, 16'd57317, 16'd64537, 16'd41783, 16'd44222, 16'd62158, 16'd25052, 16'd48918, 16'd17160, 16'd43950, 16'd29603, 16'd42030, 16'd59986, 16'd13637, 16'd49707, 16'd9585, 16'd19698, 16'd9674, 16'd60793, 16'd10396, 16'd54766});
	test_expansion(128'h6a70d3d7e1030d7a17976514a1f3de83, {16'd43831, 16'd40869, 16'd63035, 16'd2374, 16'd12071, 16'd32202, 16'd25856, 16'd52074, 16'd11490, 16'd29708, 16'd32528, 16'd12424, 16'd1129, 16'd64350, 16'd16627, 16'd11654, 16'd12186, 16'd11232, 16'd44186, 16'd5225, 16'd46101, 16'd55984, 16'd2238, 16'd49046, 16'd7574, 16'd11219});
	test_expansion(128'h13949b399fdb8cd57d5c2679bb2a73f3, {16'd36438, 16'd4605, 16'd42042, 16'd56138, 16'd49954, 16'd36383, 16'd25670, 16'd33165, 16'd55956, 16'd16469, 16'd35732, 16'd19562, 16'd39225, 16'd16100, 16'd12582, 16'd34839, 16'd43228, 16'd1067, 16'd19389, 16'd54636, 16'd33214, 16'd4078, 16'd36077, 16'd20846, 16'd65213, 16'd28987});
	test_expansion(128'h171c3cfda6772bac7e68652f77a3b5ab, {16'd51679, 16'd37419, 16'd59622, 16'd27887, 16'd32185, 16'd39285, 16'd5744, 16'd6164, 16'd60508, 16'd57159, 16'd50903, 16'd35345, 16'd32242, 16'd31785, 16'd11330, 16'd13879, 16'd48637, 16'd23938, 16'd20372, 16'd45027, 16'd57502, 16'd21264, 16'd1784, 16'd28949, 16'd27125, 16'd12306});
	test_expansion(128'h2cca2805232d3d1e63a1d8f2e6c14e1f, {16'd17188, 16'd47467, 16'd53384, 16'd55755, 16'd47707, 16'd60006, 16'd13562, 16'd18657, 16'd63816, 16'd64306, 16'd32582, 16'd55164, 16'd52276, 16'd6968, 16'd4455, 16'd31345, 16'd61656, 16'd51009, 16'd8072, 16'd7851, 16'd16214, 16'd9445, 16'd10305, 16'd29128, 16'd17552, 16'd63522});
	test_expansion(128'h4b50d01e2038645e39bd2b3804613a81, {16'd56092, 16'd27531, 16'd65488, 16'd5451, 16'd43149, 16'd58799, 16'd50097, 16'd5517, 16'd8363, 16'd13227, 16'd64931, 16'd53945, 16'd3010, 16'd21158, 16'd25344, 16'd57456, 16'd10971, 16'd22687, 16'd54680, 16'd20764, 16'd62484, 16'd49164, 16'd2771, 16'd35564, 16'd19048, 16'd28701});
	test_expansion(128'he2e2d2d1450d67f027ba1db52962cede, {16'd1864, 16'd12433, 16'd4912, 16'd9337, 16'd27234, 16'd30824, 16'd34025, 16'd1201, 16'd27788, 16'd56055, 16'd39512, 16'd38248, 16'd224, 16'd1915, 16'd55954, 16'd45631, 16'd12886, 16'd11232, 16'd51367, 16'd834, 16'd51849, 16'd60594, 16'd60500, 16'd34419, 16'd23449, 16'd46822});
	test_expansion(128'h97a2556e3ccd11b36891fe60fb9b9ec7, {16'd40282, 16'd16988, 16'd59727, 16'd54435, 16'd31017, 16'd13734, 16'd63859, 16'd14290, 16'd20667, 16'd18223, 16'd27790, 16'd22700, 16'd14189, 16'd46126, 16'd12232, 16'd59728, 16'd53309, 16'd23790, 16'd10438, 16'd55518, 16'd61481, 16'd60364, 16'd59424, 16'd7896, 16'd42338, 16'd53393});
	test_expansion(128'h8a47a356e33ddeddf89b44eeabd5ca37, {16'd14869, 16'd15080, 16'd55010, 16'd20068, 16'd33336, 16'd60577, 16'd13010, 16'd42082, 16'd9660, 16'd63131, 16'd18498, 16'd58713, 16'd31130, 16'd7335, 16'd2315, 16'd33538, 16'd19907, 16'd57095, 16'd17992, 16'd40301, 16'd23536, 16'd63965, 16'd24002, 16'd47937, 16'd52064, 16'd26250});
	test_expansion(128'h7b23ed576a36a82e06091e40e568ba28, {16'd16143, 16'd16735, 16'd54681, 16'd58180, 16'd62194, 16'd21051, 16'd47917, 16'd3084, 16'd8523, 16'd49451, 16'd17998, 16'd9069, 16'd939, 16'd54824, 16'd49309, 16'd58041, 16'd57676, 16'd65363, 16'd3737, 16'd31714, 16'd5512, 16'd24405, 16'd12551, 16'd34677, 16'd57544, 16'd38240});
	test_expansion(128'hcda8afa63f92f1f7ad79449c98b2a1f9, {16'd36518, 16'd15259, 16'd61951, 16'd2249, 16'd30849, 16'd9383, 16'd53207, 16'd37369, 16'd53999, 16'd42026, 16'd7677, 16'd47053, 16'd24141, 16'd37232, 16'd24565, 16'd38392, 16'd50018, 16'd22735, 16'd33690, 16'd15449, 16'd38069, 16'd63919, 16'd3164, 16'd40641, 16'd52456, 16'd59491});
	test_expansion(128'he0d42521ebf0922ede0eba30c380d563, {16'd59398, 16'd1797, 16'd37684, 16'd41242, 16'd43512, 16'd35037, 16'd46083, 16'd24573, 16'd29352, 16'd62697, 16'd3254, 16'd27614, 16'd49362, 16'd38223, 16'd54931, 16'd18606, 16'd6504, 16'd53159, 16'd44965, 16'd7182, 16'd54213, 16'd19655, 16'd46321, 16'd41958, 16'd777, 16'd65053});
	test_expansion(128'h473726f2a2404745a45a510552db0fc8, {16'd55593, 16'd14378, 16'd14899, 16'd2835, 16'd45834, 16'd53599, 16'd28936, 16'd11269, 16'd50575, 16'd29995, 16'd90, 16'd64834, 16'd4536, 16'd34472, 16'd10644, 16'd7886, 16'd37964, 16'd57164, 16'd39072, 16'd21957, 16'd25246, 16'd47004, 16'd11113, 16'd33042, 16'd42571, 16'd63593});
	test_expansion(128'h00bbb8b7ac0a06d20ff608e8e0dfef25, {16'd25400, 16'd50300, 16'd26237, 16'd13440, 16'd40180, 16'd23568, 16'd3823, 16'd31519, 16'd23358, 16'd28991, 16'd50724, 16'd6855, 16'd34810, 16'd22968, 16'd3477, 16'd55097, 16'd49932, 16'd36540, 16'd31843, 16'd34237, 16'd45660, 16'd23536, 16'd44590, 16'd7989, 16'd38126, 16'd54950});
	test_expansion(128'hc03778036e510e3ab02056ded33f15fd, {16'd10254, 16'd53824, 16'd28712, 16'd21045, 16'd11129, 16'd36433, 16'd21432, 16'd17212, 16'd9592, 16'd49310, 16'd18859, 16'd62762, 16'd56528, 16'd34931, 16'd44855, 16'd25650, 16'd303, 16'd36243, 16'd42144, 16'd46471, 16'd43477, 16'd63840, 16'd40109, 16'd51882, 16'd37957, 16'd15206});
	test_expansion(128'hd7ee94faad6891c7491cc1c93f93fa55, {16'd13482, 16'd30591, 16'd45819, 16'd31456, 16'd671, 16'd21602, 16'd42354, 16'd26639, 16'd35004, 16'd60368, 16'd55235, 16'd48930, 16'd48356, 16'd32655, 16'd14587, 16'd16181, 16'd53918, 16'd19595, 16'd61639, 16'd38916, 16'd51043, 16'd62592, 16'd15164, 16'd55859, 16'd1569, 16'd10671});
	test_expansion(128'h1854b283b57990fb551ad6129225a753, {16'd9291, 16'd34025, 16'd15258, 16'd16320, 16'd44634, 16'd25700, 16'd19887, 16'd24810, 16'd8675, 16'd46946, 16'd63935, 16'd42085, 16'd59871, 16'd60194, 16'd47972, 16'd21263, 16'd8630, 16'd48766, 16'd3083, 16'd58692, 16'd8192, 16'd23930, 16'd45343, 16'd59050, 16'd47472, 16'd7641});
	test_expansion(128'hfeeb7f7701e1324b93c1632ce8d5d82d, {16'd28659, 16'd31028, 16'd619, 16'd17975, 16'd10944, 16'd50531, 16'd7754, 16'd35128, 16'd62025, 16'd21785, 16'd25338, 16'd11694, 16'd29454, 16'd5286, 16'd26781, 16'd23779, 16'd15955, 16'd56812, 16'd14120, 16'd48034, 16'd44945, 16'd54037, 16'd7793, 16'd33673, 16'd6724, 16'd52125});
	test_expansion(128'hdf90343cf96a6eeb3beeb18d3c0a560f, {16'd49841, 16'd22570, 16'd1758, 16'd11316, 16'd2798, 16'd24967, 16'd12144, 16'd56962, 16'd13058, 16'd29533, 16'd8906, 16'd57958, 16'd5626, 16'd9995, 16'd28337, 16'd41883, 16'd13565, 16'd37184, 16'd23202, 16'd28747, 16'd32680, 16'd45217, 16'd17949, 16'd1353, 16'd44576, 16'd40171});
	test_expansion(128'h6c313efb88e64e882dd157188f162adc, {16'd51689, 16'd27777, 16'd55729, 16'd1689, 16'd11348, 16'd64759, 16'd18800, 16'd43175, 16'd42738, 16'd28417, 16'd62935, 16'd42408, 16'd27178, 16'd41612, 16'd45954, 16'd21828, 16'd33567, 16'd4695, 16'd59224, 16'd31919, 16'd42904, 16'd38066, 16'd23981, 16'd7484, 16'd27205, 16'd17052});
	test_expansion(128'h712b2a4392ab3f3d2a180a5c799e11aa, {16'd62632, 16'd45229, 16'd38081, 16'd28668, 16'd52819, 16'd46, 16'd23873, 16'd19745, 16'd60482, 16'd46379, 16'd46230, 16'd27549, 16'd23069, 16'd13001, 16'd63415, 16'd24605, 16'd25462, 16'd60534, 16'd10388, 16'd46997, 16'd34077, 16'd41467, 16'd8992, 16'd11183, 16'd54806, 16'd30482});
	test_expansion(128'h7ce3404c85cd1391744883bcf143250d, {16'd799, 16'd58635, 16'd40228, 16'd45166, 16'd1425, 16'd41190, 16'd63574, 16'd62253, 16'd31439, 16'd49152, 16'd11106, 16'd3253, 16'd7065, 16'd58196, 16'd48232, 16'd45942, 16'd36178, 16'd50075, 16'd9329, 16'd7066, 16'd26162, 16'd29943, 16'd42510, 16'd16497, 16'd10720, 16'd39332});
	test_expansion(128'hc76e782d5a03c1879becbcbf9651de2c, {16'd30231, 16'd53652, 16'd45966, 16'd43219, 16'd60849, 16'd64774, 16'd34184, 16'd64469, 16'd50438, 16'd56890, 16'd43883, 16'd55869, 16'd17367, 16'd26405, 16'd12886, 16'd33758, 16'd25452, 16'd12124, 16'd64092, 16'd34168, 16'd50253, 16'd56878, 16'd6907, 16'd50189, 16'd32785, 16'd38429});
	test_expansion(128'h3b873f0f84f1135369adcb2ddabc76d4, {16'd9475, 16'd28506, 16'd29264, 16'd10083, 16'd60647, 16'd4102, 16'd47587, 16'd21446, 16'd55401, 16'd30724, 16'd6863, 16'd12656, 16'd44311, 16'd57399, 16'd59905, 16'd50721, 16'd2402, 16'd44826, 16'd58714, 16'd521, 16'd7840, 16'd9263, 16'd7063, 16'd64050, 16'd46820, 16'd36840});
	test_expansion(128'h2ee63ef6bec1ea9f0f80ac6a6e90e00b, {16'd57531, 16'd9004, 16'd58204, 16'd1679, 16'd64720, 16'd43860, 16'd20429, 16'd14455, 16'd43928, 16'd62173, 16'd48609, 16'd5497, 16'd22974, 16'd51567, 16'd15764, 16'd10409, 16'd47232, 16'd37987, 16'd55514, 16'd25881, 16'd38490, 16'd21390, 16'd12272, 16'd36873, 16'd1368, 16'd33970});
	test_expansion(128'h4fcbd43841f7ebb8c1e8b60f6e30558b, {16'd12348, 16'd873, 16'd24109, 16'd61932, 16'd42480, 16'd42247, 16'd13123, 16'd38989, 16'd46097, 16'd5284, 16'd26173, 16'd18061, 16'd22329, 16'd36012, 16'd26954, 16'd28673, 16'd48502, 16'd41462, 16'd37276, 16'd45936, 16'd22971, 16'd942, 16'd48077, 16'd62676, 16'd19901, 16'd62831});
	test_expansion(128'h9171f1b9c52063abecc09433d7f399e9, {16'd23904, 16'd37316, 16'd25498, 16'd27851, 16'd61909, 16'd23049, 16'd3014, 16'd52650, 16'd29947, 16'd45433, 16'd9003, 16'd4591, 16'd48723, 16'd1797, 16'd16315, 16'd42285, 16'd65529, 16'd53011, 16'd19294, 16'd58994, 16'd31878, 16'd62201, 16'd56362, 16'd25952, 16'd55311, 16'd1563});
	test_expansion(128'hd467bde4b411cd14f3b40f48ac907683, {16'd3109, 16'd29892, 16'd51582, 16'd59774, 16'd45397, 16'd35773, 16'd26062, 16'd25557, 16'd841, 16'd12334, 16'd54677, 16'd28947, 16'd38781, 16'd28995, 16'd16758, 16'd50720, 16'd54353, 16'd38806, 16'd26375, 16'd32528, 16'd31830, 16'd23919, 16'd42708, 16'd56969, 16'd45446, 16'd46700});
	test_expansion(128'h8d5e0c65feb14d2d3df92448d3fa671c, {16'd58224, 16'd59333, 16'd12395, 16'd19157, 16'd54775, 16'd6405, 16'd11549, 16'd52349, 16'd23304, 16'd50067, 16'd32885, 16'd26781, 16'd55381, 16'd858, 16'd4339, 16'd55612, 16'd53594, 16'd43628, 16'd22291, 16'd49654, 16'd30618, 16'd22746, 16'd9750, 16'd59593, 16'd32702, 16'd58622});
	test_expansion(128'h479ab12f1350c7e308fe927de1e58d0f, {16'd61254, 16'd44697, 16'd13637, 16'd61761, 16'd14800, 16'd11216, 16'd49333, 16'd40269, 16'd30625, 16'd42910, 16'd23018, 16'd7128, 16'd40850, 16'd44866, 16'd5009, 16'd45370, 16'd4715, 16'd46965, 16'd56360, 16'd44665, 16'd24029, 16'd49206, 16'd39298, 16'd40438, 16'd21276, 16'd46253});
	test_expansion(128'h8959e933951d684483d90bee9269f3ee, {16'd29095, 16'd39681, 16'd47226, 16'd10280, 16'd53092, 16'd11407, 16'd21483, 16'd31064, 16'd4334, 16'd29439, 16'd17318, 16'd26080, 16'd26125, 16'd26011, 16'd51381, 16'd56517, 16'd39882, 16'd47741, 16'd54017, 16'd59502, 16'd10954, 16'd5175, 16'd45266, 16'd7802, 16'd20066, 16'd8632});
	test_expansion(128'haf71f160de4fffba996c2366be5e1892, {16'd58787, 16'd41984, 16'd53756, 16'd29033, 16'd39447, 16'd40309, 16'd4687, 16'd61241, 16'd40628, 16'd33163, 16'd8026, 16'd7532, 16'd41074, 16'd14077, 16'd39861, 16'd42852, 16'd60364, 16'd36373, 16'd18765, 16'd42799, 16'd13308, 16'd45201, 16'd5714, 16'd57673, 16'd50009, 16'd17596});
	test_expansion(128'h9aad41146e0fecbc8452b13fa8d18f27, {16'd941, 16'd28363, 16'd16129, 16'd47231, 16'd22537, 16'd13919, 16'd59227, 16'd56679, 16'd61016, 16'd42846, 16'd44367, 16'd49655, 16'd56964, 16'd5253, 16'd33865, 16'd26081, 16'd26536, 16'd48133, 16'd31624, 16'd57859, 16'd4142, 16'd17083, 16'd18615, 16'd61334, 16'd52378, 16'd9085});
	test_expansion(128'h9d87b0da29f9e978e30fcedff10fde23, {16'd60817, 16'd27509, 16'd28219, 16'd38635, 16'd36751, 16'd49616, 16'd22777, 16'd15101, 16'd43852, 16'd30860, 16'd46798, 16'd42886, 16'd61208, 16'd27251, 16'd8476, 16'd1232, 16'd29594, 16'd2810, 16'd11852, 16'd49906, 16'd10932, 16'd34134, 16'd60633, 16'd47686, 16'd55894, 16'd12513});
	test_expansion(128'h1ae2242d19cf5ee90e16762ca49d36e0, {16'd50369, 16'd63698, 16'd19077, 16'd6604, 16'd57013, 16'd19903, 16'd56417, 16'd54829, 16'd40811, 16'd43057, 16'd10315, 16'd64621, 16'd60721, 16'd20304, 16'd40517, 16'd2208, 16'd42729, 16'd41856, 16'd22239, 16'd20681, 16'd52862, 16'd41119, 16'd55582, 16'd55986, 16'd47963, 16'd63229});
	test_expansion(128'hbbde69a14cff3479e0006a13c2889a79, {16'd11090, 16'd57803, 16'd50718, 16'd26181, 16'd35391, 16'd65317, 16'd12979, 16'd58734, 16'd10043, 16'd36944, 16'd65440, 16'd8092, 16'd25997, 16'd55260, 16'd27158, 16'd56147, 16'd18178, 16'd60138, 16'd8404, 16'd16197, 16'd43774, 16'd55715, 16'd2736, 16'd44187, 16'd55206, 16'd25731});
	test_expansion(128'h61fd53747b8a072d7cf1cfaacc2c4c86, {16'd20281, 16'd21732, 16'd26695, 16'd2357, 16'd50546, 16'd48246, 16'd5277, 16'd29760, 16'd41926, 16'd2110, 16'd56280, 16'd5167, 16'd61151, 16'd16975, 16'd57828, 16'd60551, 16'd40370, 16'd32087, 16'd54412, 16'd32767, 16'd20079, 16'd6572, 16'd6898, 16'd7104, 16'd13053, 16'd2186});
	test_expansion(128'h2f5209a62fa753e5e87c222b8c6eea18, {16'd46727, 16'd27401, 16'd27232, 16'd59219, 16'd20916, 16'd35269, 16'd6447, 16'd43791, 16'd51014, 16'd55323, 16'd4200, 16'd3684, 16'd64457, 16'd22389, 16'd5809, 16'd43937, 16'd38757, 16'd30296, 16'd26357, 16'd47413, 16'd16006, 16'd58996, 16'd437, 16'd47988, 16'd22742, 16'd39929});
	test_expansion(128'h8071432b878cb35f7aabe13bfdada61d, {16'd4790, 16'd38151, 16'd55164, 16'd62866, 16'd10006, 16'd30699, 16'd37298, 16'd28800, 16'd44840, 16'd16763, 16'd64422, 16'd32203, 16'd14334, 16'd14205, 16'd5765, 16'd50549, 16'd19750, 16'd20161, 16'd17473, 16'd29434, 16'd10019, 16'd5658, 16'd19303, 16'd15834, 16'd8801, 16'd45133});
	test_expansion(128'hf57317f47c26366b2c79715c5893a3b7, {16'd42356, 16'd22065, 16'd45497, 16'd2043, 16'd47050, 16'd31217, 16'd43339, 16'd8203, 16'd31683, 16'd57731, 16'd26305, 16'd31092, 16'd3993, 16'd30498, 16'd5573, 16'd3582, 16'd19582, 16'd59518, 16'd41444, 16'd891, 16'd14235, 16'd55347, 16'd26835, 16'd13854, 16'd7103, 16'd22653});
	test_expansion(128'h97553ea5a9cf5f9204532449f4bbf8b8, {16'd41211, 16'd20607, 16'd46116, 16'd32296, 16'd37264, 16'd60381, 16'd57621, 16'd49701, 16'd2161, 16'd46483, 16'd34480, 16'd5502, 16'd37375, 16'd4990, 16'd44443, 16'd41598, 16'd9984, 16'd63818, 16'd41990, 16'd8751, 16'd1030, 16'd860, 16'd40628, 16'd55716, 16'd48177, 16'd41522});
	test_expansion(128'h2ddd66c52a87fc813d90bbc3ad3c0443, {16'd15372, 16'd51592, 16'd17985, 16'd37853, 16'd31223, 16'd1198, 16'd25947, 16'd26818, 16'd55283, 16'd18909, 16'd63885, 16'd17155, 16'd47314, 16'd14276, 16'd9494, 16'd7213, 16'd49789, 16'd43867, 16'd5066, 16'd37302, 16'd21158, 16'd2461, 16'd25076, 16'd2635, 16'd3371, 16'd5692});
	test_expansion(128'hdc82267f71064181a313dfa090fa69b8, {16'd7734, 16'd6403, 16'd22941, 16'd53637, 16'd63813, 16'd32468, 16'd5689, 16'd63605, 16'd16828, 16'd35631, 16'd35695, 16'd27547, 16'd55529, 16'd42523, 16'd46280, 16'd3931, 16'd4765, 16'd16750, 16'd34960, 16'd9390, 16'd48513, 16'd40617, 16'd33076, 16'd567, 16'd56855, 16'd51936});
	test_expansion(128'h38aacb31774586fefce6992fdb8447e4, {16'd3626, 16'd10091, 16'd65142, 16'd23726, 16'd15804, 16'd15659, 16'd19141, 16'd38596, 16'd48098, 16'd14197, 16'd56056, 16'd45768, 16'd63398, 16'd9436, 16'd10150, 16'd998, 16'd5049, 16'd56977, 16'd7335, 16'd59183, 16'd40102, 16'd54323, 16'd23586, 16'd53107, 16'd32860, 16'd4312});
	test_expansion(128'h3ae9ec6be72d944d0652f600b7ae68c7, {16'd22787, 16'd45072, 16'd14686, 16'd58418, 16'd12578, 16'd46143, 16'd18330, 16'd7536, 16'd27904, 16'd14983, 16'd51594, 16'd62330, 16'd14678, 16'd55562, 16'd59346, 16'd19133, 16'd17804, 16'd3290, 16'd64818, 16'd9685, 16'd41922, 16'd15462, 16'd62162, 16'd50497, 16'd55552, 16'd1065});
	test_expansion(128'hd1b79935624eb24d6423e19f9165f3fe, {16'd45814, 16'd33925, 16'd17513, 16'd34358, 16'd43601, 16'd9655, 16'd0, 16'd6698, 16'd36801, 16'd65527, 16'd1483, 16'd31411, 16'd35368, 16'd52128, 16'd35964, 16'd52462, 16'd39491, 16'd25901, 16'd51177, 16'd3293, 16'd24411, 16'd59577, 16'd32376, 16'd6243, 16'd35553, 16'd37368});
	test_expansion(128'h2c5bf12ce62a26539466855964dc0b7d, {16'd38555, 16'd21999, 16'd20294, 16'd10113, 16'd65389, 16'd40785, 16'd20916, 16'd19720, 16'd14933, 16'd49701, 16'd44443, 16'd20097, 16'd60807, 16'd36357, 16'd44648, 16'd42192, 16'd8633, 16'd14021, 16'd32533, 16'd16530, 16'd17595, 16'd153, 16'd1700, 16'd20669, 16'd11056, 16'd20072});
	test_expansion(128'h66c29c50537047a05480fd0b137f654f, {16'd2023, 16'd23878, 16'd47518, 16'd26913, 16'd21399, 16'd31893, 16'd44070, 16'd2355, 16'd42919, 16'd39884, 16'd45036, 16'd23708, 16'd47241, 16'd62152, 16'd60903, 16'd42769, 16'd29060, 16'd44029, 16'd26277, 16'd26012, 16'd36649, 16'd5747, 16'd55503, 16'd2255, 16'd2462, 16'd20770});
	test_expansion(128'h6eaf9969a981a75583a091206659a993, {16'd50259, 16'd17705, 16'd26890, 16'd2586, 16'd7901, 16'd15365, 16'd53412, 16'd34007, 16'd14233, 16'd11199, 16'd53241, 16'd9938, 16'd56621, 16'd49494, 16'd54190, 16'd5570, 16'd51348, 16'd38346, 16'd3945, 16'd28058, 16'd2602, 16'd10091, 16'd49537, 16'd51645, 16'd15162, 16'd49537});
	test_expansion(128'hb78b1e94c53eca0172af4bec64bf9a71, {16'd37342, 16'd3367, 16'd47363, 16'd24593, 16'd41826, 16'd45660, 16'd51189, 16'd61487, 16'd8340, 16'd61513, 16'd11138, 16'd3570, 16'd61716, 16'd63364, 16'd64895, 16'd2147, 16'd43226, 16'd30619, 16'd55139, 16'd34447, 16'd27688, 16'd2484, 16'd58945, 16'd55176, 16'd35287, 16'd54757});
	test_expansion(128'h0d9a08a79b150e9ce6318e4815c60311, {16'd47624, 16'd35046, 16'd31688, 16'd53743, 16'd55478, 16'd51977, 16'd57334, 16'd2036, 16'd62791, 16'd59753, 16'd6947, 16'd23340, 16'd9487, 16'd34933, 16'd40713, 16'd29356, 16'd46780, 16'd23793, 16'd37756, 16'd57290, 16'd46701, 16'd11427, 16'd7134, 16'd53390, 16'd48427, 16'd50129});
	test_expansion(128'ha1ae820d23b7251fa8329819d0b7d6ca, {16'd9726, 16'd34086, 16'd18723, 16'd14250, 16'd59120, 16'd8705, 16'd5512, 16'd61977, 16'd2901, 16'd35119, 16'd16088, 16'd32528, 16'd47900, 16'd34787, 16'd62805, 16'd57034, 16'd15700, 16'd54456, 16'd39039, 16'd43168, 16'd29654, 16'd8752, 16'd43833, 16'd52933, 16'd21660, 16'd47898});
	test_expansion(128'ha3305cfcd6d3d5ccf5b424c32564b338, {16'd20437, 16'd45079, 16'd50708, 16'd36366, 16'd7681, 16'd43848, 16'd37118, 16'd41539, 16'd35916, 16'd53889, 16'd36115, 16'd22100, 16'd47875, 16'd2845, 16'd32969, 16'd32351, 16'd62454, 16'd29582, 16'd15279, 16'd30955, 16'd34792, 16'd48995, 16'd40698, 16'd5456, 16'd61475, 16'd52285});
	test_expansion(128'h1ee1c4a644b9fedd8b3e22bbae3f93c2, {16'd21402, 16'd28974, 16'd50333, 16'd39480, 16'd17872, 16'd42460, 16'd7653, 16'd52109, 16'd22773, 16'd28194, 16'd30103, 16'd19478, 16'd54773, 16'd9495, 16'd7120, 16'd32260, 16'd28443, 16'd34467, 16'd11517, 16'd13452, 16'd32676, 16'd38649, 16'd63140, 16'd55705, 16'd23730, 16'd9694});
	test_expansion(128'he566882c048b17b81f5c918e8e2df584, {16'd46759, 16'd28823, 16'd26442, 16'd21961, 16'd27720, 16'd3685, 16'd26800, 16'd7891, 16'd14705, 16'd51760, 16'd47895, 16'd21613, 16'd22979, 16'd40121, 16'd20554, 16'd37615, 16'd55087, 16'd37875, 16'd2199, 16'd37445, 16'd40100, 16'd45657, 16'd62587, 16'd3458, 16'd31087, 16'd46465});
	test_expansion(128'h6c8470392e0106b4b689e3022e1c19ec, {16'd25074, 16'd30859, 16'd42862, 16'd25314, 16'd58732, 16'd56401, 16'd18844, 16'd56862, 16'd56116, 16'd57865, 16'd64374, 16'd38747, 16'd15659, 16'd37259, 16'd46090, 16'd35028, 16'd15886, 16'd9490, 16'd15773, 16'd52923, 16'd566, 16'd56820, 16'd14046, 16'd5231, 16'd41522, 16'd1565});
	test_expansion(128'h03c91a6050c5b4a6a08e817cb751e30a, {16'd48708, 16'd7313, 16'd39925, 16'd34278, 16'd4172, 16'd45299, 16'd21456, 16'd63524, 16'd6725, 16'd30612, 16'd26418, 16'd29162, 16'd59304, 16'd22342, 16'd29433, 16'd39318, 16'd26662, 16'd7492, 16'd3496, 16'd18678, 16'd12316, 16'd10770, 16'd29150, 16'd58354, 16'd41465, 16'd29027});
	test_expansion(128'h6903c49e21b32dfb2ed3ff1a72e71ea2, {16'd18031, 16'd59399, 16'd54874, 16'd34010, 16'd63451, 16'd6751, 16'd4874, 16'd59726, 16'd19638, 16'd35711, 16'd49002, 16'd15593, 16'd50350, 16'd58579, 16'd31788, 16'd21579, 16'd799, 16'd5187, 16'd58957, 16'd38437, 16'd9105, 16'd58760, 16'd40601, 16'd57499, 16'd21714, 16'd40674});
	test_expansion(128'hfd285bd6c9663f5e7bd1a948d115210f, {16'd21077, 16'd55173, 16'd21032, 16'd46309, 16'd44543, 16'd20984, 16'd41244, 16'd23076, 16'd56435, 16'd8965, 16'd60191, 16'd10588, 16'd31294, 16'd63110, 16'd5949, 16'd22168, 16'd25603, 16'd34337, 16'd6719, 16'd154, 16'd530, 16'd8979, 16'd47572, 16'd48507, 16'd19056, 16'd1670});
	test_expansion(128'h9a9a23ebb7e29323bc71d4eb10ecfee2, {16'd32991, 16'd3233, 16'd14251, 16'd17579, 16'd36862, 16'd26759, 16'd56687, 16'd32678, 16'd59983, 16'd47532, 16'd63159, 16'd57879, 16'd51874, 16'd8861, 16'd22638, 16'd37314, 16'd32305, 16'd38737, 16'd64340, 16'd51282, 16'd53041, 16'd30339, 16'd4986, 16'd52034, 16'd59597, 16'd2415});
	test_expansion(128'h7cef3714f1a0eb01fefa731e9aeb1873, {16'd55555, 16'd34446, 16'd11547, 16'd15249, 16'd11354, 16'd61846, 16'd5862, 16'd38723, 16'd16427, 16'd43303, 16'd58855, 16'd30749, 16'd59843, 16'd61172, 16'd10581, 16'd3835, 16'd52321, 16'd19803, 16'd39708, 16'd47828, 16'd35113, 16'd46845, 16'd49463, 16'd58599, 16'd57125, 16'd18801});
	test_expansion(128'h0ebc673aa292158ea6c6e13897ed99c1, {16'd41409, 16'd13063, 16'd23859, 16'd12086, 16'd3460, 16'd26357, 16'd13806, 16'd13673, 16'd49869, 16'd39780, 16'd46387, 16'd14073, 16'd9289, 16'd33511, 16'd41742, 16'd9916, 16'd11532, 16'd11692, 16'd62289, 16'd48692, 16'd56208, 16'd24463, 16'd15156, 16'd18542, 16'd29986, 16'd44983});
	test_expansion(128'hebbe779d5a230f5213e0341fbd893681, {16'd6225, 16'd57631, 16'd2293, 16'd56782, 16'd61400, 16'd57604, 16'd59519, 16'd58166, 16'd47582, 16'd10865, 16'd18015, 16'd42183, 16'd2490, 16'd1134, 16'd22459, 16'd21547, 16'd60230, 16'd47919, 16'd10492, 16'd6447, 16'd14825, 16'd359, 16'd37587, 16'd32823, 16'd33115, 16'd19983});
	test_expansion(128'h8b72a2e6df51947805d9d199a529afa6, {16'd36565, 16'd32912, 16'd6358, 16'd31034, 16'd4114, 16'd2959, 16'd13391, 16'd23472, 16'd13346, 16'd53346, 16'd27661, 16'd15535, 16'd40935, 16'd60539, 16'd51328, 16'd47549, 16'd18709, 16'd62297, 16'd29965, 16'd19788, 16'd18938, 16'd6685, 16'd80, 16'd57251, 16'd20078, 16'd32870});
	test_expansion(128'h8e77fc6ca1ab6627e6ff6bc2acba19c0, {16'd12751, 16'd34713, 16'd39327, 16'd42703, 16'd61391, 16'd52269, 16'd16956, 16'd37423, 16'd1429, 16'd39347, 16'd20388, 16'd9315, 16'd26847, 16'd553, 16'd32118, 16'd63327, 16'd13889, 16'd63132, 16'd51173, 16'd752, 16'd62298, 16'd31428, 16'd60423, 16'd54646, 16'd45600, 16'd29718});
	test_expansion(128'hff3124d01819409475da48f02d3542ff, {16'd21610, 16'd60055, 16'd48815, 16'd59883, 16'd50281, 16'd41253, 16'd45009, 16'd48109, 16'd15506, 16'd6974, 16'd12106, 16'd5710, 16'd11699, 16'd14058, 16'd9316, 16'd13187, 16'd25504, 16'd8674, 16'd38292, 16'd43109, 16'd15805, 16'd21250, 16'd65231, 16'd37833, 16'd46633, 16'd10824});
	test_expansion(128'hedaa8ad550e3a0f13feb9aaf5fa6e831, {16'd53911, 16'd9883, 16'd57211, 16'd4395, 16'd26014, 16'd41379, 16'd48544, 16'd53872, 16'd12507, 16'd5378, 16'd64194, 16'd58429, 16'd38327, 16'd39391, 16'd49601, 16'd14471, 16'd7360, 16'd19920, 16'd32736, 16'd45683, 16'd54103, 16'd11348, 16'd49684, 16'd17162, 16'd4981, 16'd20467});
	test_expansion(128'ha1190d01ee70ff5c59c96aa570679c23, {16'd25444, 16'd28439, 16'd7631, 16'd46949, 16'd53851, 16'd30368, 16'd42701, 16'd6869, 16'd5941, 16'd56248, 16'd12807, 16'd34105, 16'd57955, 16'd36310, 16'd20238, 16'd4814, 16'd13704, 16'd61608, 16'd1752, 16'd35979, 16'd4751, 16'd5584, 16'd54699, 16'd41650, 16'd7565, 16'd26484});
	test_expansion(128'h16f976f1398a3befe8559dbacd62d694, {16'd25358, 16'd27160, 16'd4391, 16'd4679, 16'd48280, 16'd7705, 16'd43794, 16'd34702, 16'd15071, 16'd36281, 16'd1719, 16'd48731, 16'd13116, 16'd42260, 16'd34721, 16'd16509, 16'd22168, 16'd625, 16'd53656, 16'd58888, 16'd51887, 16'd25576, 16'd26525, 16'd8225, 16'd16075, 16'd40665});
	test_expansion(128'hcf29f8417472f1d228188175582c801a, {16'd23359, 16'd22734, 16'd51410, 16'd4580, 16'd20439, 16'd22355, 16'd40870, 16'd33040, 16'd59917, 16'd43528, 16'd39931, 16'd63306, 16'd29775, 16'd49025, 16'd60869, 16'd24870, 16'd28428, 16'd25277, 16'd34812, 16'd10870, 16'd33982, 16'd32425, 16'd10632, 16'd27126, 16'd20326, 16'd43818});
	test_expansion(128'h6489162948d92de7544f2349cd896bb7, {16'd50993, 16'd10065, 16'd45216, 16'd54812, 16'd5579, 16'd18455, 16'd48150, 16'd36209, 16'd754, 16'd19359, 16'd4638, 16'd36987, 16'd22289, 16'd6221, 16'd48050, 16'd3566, 16'd15293, 16'd8869, 16'd13625, 16'd18477, 16'd2543, 16'd10254, 16'd63020, 16'd44861, 16'd3162, 16'd47866});
	test_expansion(128'h3ca658c6016fe96d9fa0af2165444535, {16'd42849, 16'd41904, 16'd7102, 16'd18263, 16'd33921, 16'd34212, 16'd26354, 16'd24533, 16'd44965, 16'd20680, 16'd63099, 16'd58528, 16'd17539, 16'd8839, 16'd65309, 16'd27219, 16'd50935, 16'd3775, 16'd698, 16'd30846, 16'd42877, 16'd16073, 16'd56712, 16'd21282, 16'd30653, 16'd8950});
	test_expansion(128'h704e42ffa4337ca156496da23759260e, {16'd21069, 16'd16109, 16'd22884, 16'd12256, 16'd19702, 16'd27782, 16'd29906, 16'd34050, 16'd31127, 16'd16983, 16'd48284, 16'd10887, 16'd60953, 16'd46885, 16'd16535, 16'd60680, 16'd63974, 16'd8030, 16'd24749, 16'd60532, 16'd41930, 16'd4901, 16'd34248, 16'd51430, 16'd46629, 16'd35202});
	test_expansion(128'hd5f322a0abe40ce4eb727e075127d120, {16'd17190, 16'd11014, 16'd64063, 16'd32664, 16'd51436, 16'd55781, 16'd13767, 16'd57170, 16'd26971, 16'd23847, 16'd36138, 16'd64410, 16'd29417, 16'd42944, 16'd32034, 16'd57284, 16'd56394, 16'd24044, 16'd49035, 16'd31531, 16'd41277, 16'd45686, 16'd62158, 16'd31251, 16'd19592, 16'd8511});
	test_expansion(128'he3001ff1bb890e312b22dc076829cea3, {16'd44731, 16'd34267, 16'd49202, 16'd18440, 16'd29618, 16'd46832, 16'd33716, 16'd15538, 16'd65480, 16'd9832, 16'd43752, 16'd63264, 16'd53526, 16'd44075, 16'd4089, 16'd36484, 16'd8547, 16'd17898, 16'd12409, 16'd2152, 16'd64668, 16'd5867, 16'd12529, 16'd30289, 16'd53462, 16'd65054});
	test_expansion(128'h9323c93567c6ff3eefd7e713c75e36e5, {16'd49109, 16'd21288, 16'd56634, 16'd51094, 16'd47216, 16'd14248, 16'd45808, 16'd60760, 16'd22894, 16'd27451, 16'd7324, 16'd9073, 16'd57351, 16'd41656, 16'd61756, 16'd52845, 16'd16082, 16'd14491, 16'd20350, 16'd53139, 16'd24720, 16'd42859, 16'd24107, 16'd23302, 16'd28452, 16'd48353});
	test_expansion(128'h8f63ebe3c23f5e2d832df0cd702686f2, {16'd19098, 16'd21252, 16'd16009, 16'd16615, 16'd31863, 16'd35312, 16'd37996, 16'd7485, 16'd47712, 16'd5741, 16'd1387, 16'd55716, 16'd29923, 16'd43354, 16'd1234, 16'd43018, 16'd32055, 16'd23363, 16'd40821, 16'd31191, 16'd23261, 16'd10575, 16'd2436, 16'd63192, 16'd47639, 16'd40770});
	test_expansion(128'h18237aaae58f8a5332478944bddc9fea, {16'd57208, 16'd43120, 16'd34960, 16'd25803, 16'd20635, 16'd35864, 16'd31444, 16'd45401, 16'd58988, 16'd17959, 16'd60207, 16'd9958, 16'd19034, 16'd41113, 16'd56519, 16'd43479, 16'd49315, 16'd2402, 16'd50661, 16'd21691, 16'd34336, 16'd40404, 16'd29030, 16'd46333, 16'd11522, 16'd55446});
	test_expansion(128'h9de5bc8aba630505ce5cd6fd6c8ee9ab, {16'd20989, 16'd55558, 16'd2338, 16'd32827, 16'd45780, 16'd5491, 16'd57999, 16'd41902, 16'd10241, 16'd20038, 16'd25335, 16'd12853, 16'd54933, 16'd34725, 16'd15666, 16'd47361, 16'd177, 16'd47921, 16'd46254, 16'd58430, 16'd13406, 16'd53405, 16'd60477, 16'd22233, 16'd65287, 16'd28986});
	test_expansion(128'hd031c9c45fef3e116904a3e34220f810, {16'd59805, 16'd49487, 16'd54844, 16'd57612, 16'd28953, 16'd64920, 16'd60792, 16'd30988, 16'd57797, 16'd20117, 16'd26991, 16'd62526, 16'd10343, 16'd15063, 16'd22474, 16'd58340, 16'd44932, 16'd62593, 16'd46354, 16'd18421, 16'd62718, 16'd64034, 16'd12634, 16'd61085, 16'd12511, 16'd20027});
	test_expansion(128'h3b71400106577e22e2b3c4c92f4cc63d, {16'd54486, 16'd7683, 16'd61035, 16'd58251, 16'd37957, 16'd2126, 16'd10054, 16'd62969, 16'd40261, 16'd59722, 16'd9520, 16'd4521, 16'd24415, 16'd6174, 16'd20308, 16'd33483, 16'd53758, 16'd47435, 16'd42742, 16'd20901, 16'd24216, 16'd43376, 16'd21459, 16'd24162, 16'd12319, 16'd51184});
	test_expansion(128'hbd6080fb99db1afb1792a9e4c90e25fb, {16'd8602, 16'd50134, 16'd36327, 16'd50132, 16'd10945, 16'd6193, 16'd5584, 16'd60626, 16'd13177, 16'd39772, 16'd55403, 16'd35577, 16'd45779, 16'd28093, 16'd8353, 16'd15545, 16'd29686, 16'd8418, 16'd52494, 16'd37428, 16'd22143, 16'd35126, 16'd44183, 16'd16750, 16'd12036, 16'd40825});
	test_expansion(128'h8744342c56d39dbc99aefcf76b1735c4, {16'd60742, 16'd60543, 16'd62764, 16'd7130, 16'd46437, 16'd63704, 16'd40565, 16'd38474, 16'd58991, 16'd50577, 16'd60875, 16'd28528, 16'd48091, 16'd38461, 16'd45481, 16'd29637, 16'd41574, 16'd63624, 16'd1100, 16'd42777, 16'd1492, 16'd24636, 16'd50620, 16'd24865, 16'd37574, 16'd42957});
	test_expansion(128'h3bec6e3bdb9140b0043112315e6893ee, {16'd8628, 16'd8951, 16'd9644, 16'd2211, 16'd256, 16'd18622, 16'd5310, 16'd52368, 16'd59282, 16'd62123, 16'd37234, 16'd38526, 16'd14198, 16'd33119, 16'd41146, 16'd54207, 16'd11066, 16'd47535, 16'd56385, 16'd25279, 16'd30755, 16'd24089, 16'd42203, 16'd26019, 16'd47102, 16'd28560});
	test_expansion(128'h548eac21096e2103b9b19cee7ae82e55, {16'd51850, 16'd15222, 16'd62740, 16'd35024, 16'd50355, 16'd5003, 16'd12294, 16'd40392, 16'd48916, 16'd45235, 16'd52311, 16'd22985, 16'd44220, 16'd61691, 16'd35880, 16'd49198, 16'd55573, 16'd43780, 16'd62408, 16'd44929, 16'd53395, 16'd36107, 16'd30133, 16'd62393, 16'd14055, 16'd21427});
	test_expansion(128'h513bd8fd670922de98eab416531a3ad4, {16'd14590, 16'd50881, 16'd60151, 16'd11202, 16'd7152, 16'd56772, 16'd50110, 16'd37092, 16'd57972, 16'd44197, 16'd49899, 16'd48455, 16'd46031, 16'd14818, 16'd46394, 16'd31771, 16'd12764, 16'd64537, 16'd6265, 16'd51086, 16'd34905, 16'd59577, 16'd36807, 16'd13659, 16'd20701, 16'd61025});
	test_expansion(128'h1aa66c5fbe25bc9f714fca792a48be86, {16'd32743, 16'd46460, 16'd29856, 16'd62577, 16'd37073, 16'd57668, 16'd1432, 16'd28882, 16'd13043, 16'd53009, 16'd49236, 16'd42022, 16'd40862, 16'd19085, 16'd44922, 16'd31197, 16'd27281, 16'd15969, 16'd31024, 16'd8666, 16'd62723, 16'd14424, 16'd12054, 16'd17131, 16'd60622, 16'd49806});
	test_expansion(128'h1b34f1926b13afb7769274c6ec90bf34, {16'd31398, 16'd51254, 16'd40728, 16'd14460, 16'd9010, 16'd1295, 16'd7805, 16'd53588, 16'd59457, 16'd55555, 16'd64682, 16'd35961, 16'd58579, 16'd2139, 16'd36051, 16'd11148, 16'd39519, 16'd49853, 16'd26216, 16'd50618, 16'd677, 16'd51838, 16'd11788, 16'd52104, 16'd52945, 16'd47677});
	test_expansion(128'h20cafa41f89da951d049ff3f1f99e3b6, {16'd64009, 16'd1812, 16'd21442, 16'd43972, 16'd12504, 16'd47088, 16'd44225, 16'd23546, 16'd57406, 16'd58487, 16'd44357, 16'd61073, 16'd60165, 16'd64243, 16'd6069, 16'd42219, 16'd21406, 16'd40208, 16'd18444, 16'd64840, 16'd55682, 16'd21417, 16'd2624, 16'd63939, 16'd28443, 16'd65174});
	test_expansion(128'hb38c550c2668f44c08937189e02f002d, {16'd17081, 16'd37309, 16'd64905, 16'd29877, 16'd4044, 16'd24667, 16'd19795, 16'd31720, 16'd1650, 16'd22418, 16'd39781, 16'd27580, 16'd11629, 16'd54084, 16'd18509, 16'd46355, 16'd5613, 16'd61061, 16'd26287, 16'd11004, 16'd64754, 16'd36879, 16'd19808, 16'd19282, 16'd57778, 16'd10948});
	test_expansion(128'hb9afbd5d9ad01062a646cdd69017ab35, {16'd22931, 16'd51129, 16'd15484, 16'd56275, 16'd50260, 16'd15435, 16'd17383, 16'd24542, 16'd37403, 16'd31913, 16'd40618, 16'd40209, 16'd60900, 16'd47301, 16'd56321, 16'd27925, 16'd5935, 16'd58924, 16'd24205, 16'd24099, 16'd16802, 16'd50256, 16'd49336, 16'd54436, 16'd23023, 16'd31717});
	test_expansion(128'h86e297239d6978d6d59743d5b401caa8, {16'd65249, 16'd18924, 16'd60238, 16'd49050, 16'd33354, 16'd56470, 16'd47662, 16'd45308, 16'd5712, 16'd39102, 16'd51117, 16'd24973, 16'd2103, 16'd17573, 16'd29756, 16'd2217, 16'd3036, 16'd28610, 16'd60451, 16'd61577, 16'd14226, 16'd31849, 16'd49827, 16'd1471, 16'd38792, 16'd6640});
	test_expansion(128'hfebe1ca3dfb941e3f9e35ecdbf7bcec3, {16'd19841, 16'd24566, 16'd1940, 16'd13481, 16'd58162, 16'd47715, 16'd12836, 16'd49343, 16'd61260, 16'd28547, 16'd6622, 16'd23734, 16'd24132, 16'd2351, 16'd54458, 16'd19997, 16'd36940, 16'd32539, 16'd56819, 16'd10533, 16'd10218, 16'd27373, 16'd40095, 16'd4575, 16'd28696, 16'd5575});
	test_expansion(128'haac0d179b0b8d4749ea401e3f3dc1a62, {16'd5391, 16'd10435, 16'd51095, 16'd31771, 16'd24494, 16'd49668, 16'd57531, 16'd52876, 16'd56512, 16'd28328, 16'd15345, 16'd26405, 16'd54823, 16'd27882, 16'd30637, 16'd35266, 16'd7321, 16'd42102, 16'd61116, 16'd3574, 16'd45479, 16'd58106, 16'd55757, 16'd545, 16'd58167, 16'd32618});
	test_expansion(128'h9b205f10d19b303546973077eb6f709f, {16'd60884, 16'd31164, 16'd60814, 16'd55953, 16'd14575, 16'd40952, 16'd17132, 16'd12184, 16'd29151, 16'd17964, 16'd34913, 16'd31317, 16'd2858, 16'd65077, 16'd57704, 16'd50522, 16'd33440, 16'd743, 16'd16330, 16'd34590, 16'd40689, 16'd12367, 16'd40346, 16'd8629, 16'd23482, 16'd27191});
	test_expansion(128'h2fab5d674f8d6fa0eae54e3aa8496ca4, {16'd20885, 16'd45628, 16'd15747, 16'd20732, 16'd36119, 16'd40965, 16'd29358, 16'd37301, 16'd27236, 16'd3017, 16'd899, 16'd30674, 16'd35158, 16'd65145, 16'd47744, 16'd32685, 16'd59246, 16'd41197, 16'd64087, 16'd63589, 16'd30470, 16'd41684, 16'd7882, 16'd43997, 16'd65411, 16'd55936});
	test_expansion(128'h810ec1eecbf85cd1aa4d3f6026a48f9b, {16'd22666, 16'd15332, 16'd10586, 16'd57428, 16'd23201, 16'd14147, 16'd28465, 16'd30072, 16'd22645, 16'd9639, 16'd12428, 16'd8274, 16'd31742, 16'd62516, 16'd13726, 16'd5844, 16'd57216, 16'd51619, 16'd44840, 16'd49543, 16'd55283, 16'd6393, 16'd30622, 16'd47557, 16'd7655, 16'd25567});
	test_expansion(128'hd3c3c13c88c77263ebc10e2f9164339d, {16'd22353, 16'd6091, 16'd52906, 16'd46750, 16'd15904, 16'd23894, 16'd35545, 16'd9907, 16'd52172, 16'd44481, 16'd28013, 16'd14698, 16'd26940, 16'd34376, 16'd30641, 16'd61870, 16'd27366, 16'd29147, 16'd62056, 16'd42988, 16'd62534, 16'd5950, 16'd7081, 16'd49307, 16'd56645, 16'd4857});
	test_expansion(128'h25200c2d91f0ac1f6c59aea4aaf3141c, {16'd38460, 16'd2536, 16'd34537, 16'd60100, 16'd40844, 16'd45466, 16'd54286, 16'd31556, 16'd26441, 16'd58586, 16'd58789, 16'd27342, 16'd63160, 16'd20134, 16'd43896, 16'd22113, 16'd51211, 16'd6739, 16'd7037, 16'd65271, 16'd22972, 16'd22483, 16'd43141, 16'd44313, 16'd17627, 16'd37605});
	test_expansion(128'h7e9bd98c52b8fe7450909764d8ddaf17, {16'd63834, 16'd5843, 16'd45684, 16'd8961, 16'd4442, 16'd29172, 16'd45336, 16'd44089, 16'd18307, 16'd18636, 16'd19255, 16'd35947, 16'd44396, 16'd58022, 16'd61037, 16'd43028, 16'd27108, 16'd51431, 16'd9369, 16'd1384, 16'd59747, 16'd7584, 16'd49498, 16'd9166, 16'd13067, 16'd36312});
	test_expansion(128'hbb142c67cceca8ecc8868213e822a9aa, {16'd38203, 16'd13617, 16'd57724, 16'd61598, 16'd41073, 16'd25130, 16'd41981, 16'd32317, 16'd34297, 16'd3819, 16'd19814, 16'd58893, 16'd3448, 16'd38090, 16'd48552, 16'd41101, 16'd30087, 16'd63396, 16'd154, 16'd49691, 16'd50724, 16'd55194, 16'd55052, 16'd37388, 16'd57652, 16'd41966});
	test_expansion(128'hb1ce7a7ffd4143067635fd3beb3f6283, {16'd63628, 16'd6570, 16'd36945, 16'd58728, 16'd46581, 16'd21564, 16'd7185, 16'd47157, 16'd40683, 16'd9752, 16'd21329, 16'd47801, 16'd15094, 16'd30089, 16'd17790, 16'd23322, 16'd13940, 16'd9094, 16'd27274, 16'd17350, 16'd36233, 16'd21989, 16'd6472, 16'd38699, 16'd43569, 16'd53637});
	test_expansion(128'hf6a480b39df1f6b31e0dd81ac7740fe9, {16'd54693, 16'd35848, 16'd37015, 16'd39106, 16'd25448, 16'd28358, 16'd23030, 16'd44743, 16'd19109, 16'd3717, 16'd26680, 16'd40090, 16'd29903, 16'd34397, 16'd38802, 16'd63859, 16'd38186, 16'd9005, 16'd54565, 16'd21951, 16'd50384, 16'd48223, 16'd23728, 16'd22615, 16'd62467, 16'd14639});
	test_expansion(128'h8d6ffb456f7222c446249ffb39eab0e2, {16'd55787, 16'd40409, 16'd15475, 16'd30528, 16'd5616, 16'd12213, 16'd34128, 16'd46937, 16'd16585, 16'd42815, 16'd7286, 16'd32927, 16'd4409, 16'd39284, 16'd17037, 16'd37453, 16'd20367, 16'd6272, 16'd48554, 16'd60182, 16'd28531, 16'd17386, 16'd6986, 16'd36294, 16'd6428, 16'd19209});
	test_expansion(128'h9a984d8c9f3ea7764632fcee8f2bbed6, {16'd5268, 16'd27124, 16'd16652, 16'd39937, 16'd42501, 16'd31110, 16'd47166, 16'd32971, 16'd3293, 16'd41387, 16'd36413, 16'd8417, 16'd45944, 16'd59178, 16'd37924, 16'd7357, 16'd41255, 16'd55448, 16'd3268, 16'd11923, 16'd57207, 16'd62282, 16'd64187, 16'd51012, 16'd22484, 16'd50924});
	test_expansion(128'h8b115bc0dc74c86c11364098f29a7ca4, {16'd46962, 16'd763, 16'd62393, 16'd9292, 16'd54816, 16'd4777, 16'd16971, 16'd11657, 16'd27933, 16'd6844, 16'd44365, 16'd33122, 16'd58495, 16'd3356, 16'd33135, 16'd15573, 16'd59462, 16'd15757, 16'd54426, 16'd22832, 16'd24107, 16'd18966, 16'd1356, 16'd35288, 16'd44718, 16'd29558});
	test_expansion(128'hfbc2b5c4c5ebec723e2556ab1e87efb2, {16'd2255, 16'd61360, 16'd24888, 16'd36852, 16'd11013, 16'd23662, 16'd40552, 16'd29597, 16'd16592, 16'd60650, 16'd57690, 16'd65102, 16'd60926, 16'd20806, 16'd3648, 16'd29052, 16'd29014, 16'd52949, 16'd13175, 16'd35373, 16'd58985, 16'd45998, 16'd47358, 16'd3487, 16'd62591, 16'd9372});
	test_expansion(128'haa50dc43ebe3aa98f28e1a9407ccd354, {16'd53671, 16'd55063, 16'd16716, 16'd655, 16'd5176, 16'd24310, 16'd45221, 16'd64452, 16'd53561, 16'd11833, 16'd42487, 16'd16107, 16'd60960, 16'd41462, 16'd9183, 16'd26676, 16'd46394, 16'd4638, 16'd7044, 16'd64575, 16'd47884, 16'd63122, 16'd25636, 16'd6915, 16'd40996, 16'd27644});
	test_expansion(128'hcbe799644750f039622a6a6e2c968abc, {16'd44257, 16'd36479, 16'd46025, 16'd20969, 16'd40290, 16'd31999, 16'd27379, 16'd43683, 16'd53316, 16'd54296, 16'd44858, 16'd18516, 16'd51216, 16'd42504, 16'd56471, 16'd22784, 16'd21065, 16'd44705, 16'd63050, 16'd8885, 16'd13006, 16'd63479, 16'd26252, 16'd51241, 16'd47724, 16'd57128});
	test_expansion(128'h5a6a00950c05958e26ebfc4982090f09, {16'd54820, 16'd12729, 16'd59766, 16'd36298, 16'd14216, 16'd54808, 16'd48483, 16'd1448, 16'd34766, 16'd16242, 16'd26166, 16'd20598, 16'd19313, 16'd13133, 16'd3662, 16'd3432, 16'd57245, 16'd50071, 16'd5213, 16'd2717, 16'd50785, 16'd26399, 16'd12553, 16'd40704, 16'd29072, 16'd44692});
	test_expansion(128'hf55d6a98a6b6eeb24932b0111c462af6, {16'd56922, 16'd50461, 16'd46610, 16'd53478, 16'd38481, 16'd7774, 16'd58400, 16'd8022, 16'd64912, 16'd7329, 16'd44554, 16'd30839, 16'd60587, 16'd16131, 16'd10008, 16'd22330, 16'd18782, 16'd14272, 16'd18860, 16'd54941, 16'd46476, 16'd24742, 16'd33255, 16'd40279, 16'd1878, 16'd58747});
	test_expansion(128'h7b62f68787d74505425f6a693bb7f077, {16'd16637, 16'd47319, 16'd38640, 16'd61724, 16'd18395, 16'd48799, 16'd4367, 16'd37953, 16'd51103, 16'd58997, 16'd10308, 16'd57572, 16'd13146, 16'd46756, 16'd56322, 16'd42258, 16'd29271, 16'd11824, 16'd33835, 16'd65328, 16'd17813, 16'd219, 16'd26888, 16'd55604, 16'd5945, 16'd5527});
	test_expansion(128'h2cc2f2df00642dd08b48e73b9e9459b2, {16'd16834, 16'd60700, 16'd22221, 16'd63085, 16'd43785, 16'd45242, 16'd5575, 16'd29303, 16'd22213, 16'd3602, 16'd17591, 16'd5086, 16'd34134, 16'd17030, 16'd59307, 16'd34310, 16'd59684, 16'd33542, 16'd54666, 16'd62857, 16'd50414, 16'd10782, 16'd43423, 16'd10457, 16'd38049, 16'd64367});
	test_expansion(128'h03a12367b8d0d3484ebb071a4905a119, {16'd19555, 16'd58352, 16'd63671, 16'd6381, 16'd59693, 16'd41260, 16'd2468, 16'd55259, 16'd16248, 16'd62866, 16'd62022, 16'd34407, 16'd35527, 16'd16460, 16'd50404, 16'd47027, 16'd41043, 16'd6725, 16'd55174, 16'd4933, 16'd16671, 16'd15231, 16'd1262, 16'd21779, 16'd64313, 16'd30338});
	test_expansion(128'h93bc757f87e3b967bcb46991186bcb42, {16'd38697, 16'd10685, 16'd41366, 16'd7977, 16'd61099, 16'd36798, 16'd38727, 16'd59750, 16'd25644, 16'd43339, 16'd3493, 16'd11747, 16'd40324, 16'd57081, 16'd57373, 16'd32939, 16'd2373, 16'd3025, 16'd46367, 16'd48133, 16'd48848, 16'd47303, 16'd56830, 16'd35695, 16'd46377, 16'd45405});
	test_expansion(128'h0169ded84ea68f004d8a93487cd000f6, {16'd38139, 16'd25997, 16'd21643, 16'd40306, 16'd50919, 16'd32426, 16'd56297, 16'd51143, 16'd54694, 16'd24632, 16'd6587, 16'd5788, 16'd35953, 16'd12785, 16'd15087, 16'd11263, 16'd3813, 16'd48212, 16'd21743, 16'd13960, 16'd51698, 16'd34666, 16'd21236, 16'd61796, 16'd85, 16'd5758});
	test_expansion(128'h169ccd57286a6f19749801acc9274751, {16'd1109, 16'd31302, 16'd54128, 16'd41302, 16'd12701, 16'd18733, 16'd34922, 16'd52996, 16'd27795, 16'd1864, 16'd44569, 16'd35661, 16'd49134, 16'd30627, 16'd14981, 16'd9757, 16'd328, 16'd49662, 16'd43594, 16'd60947, 16'd35434, 16'd55214, 16'd39420, 16'd43464, 16'd30143, 16'd45953});
	test_expansion(128'h2b345cf8d4d57756d1ab87b830126027, {16'd63217, 16'd14624, 16'd3347, 16'd9788, 16'd23982, 16'd37991, 16'd3426, 16'd42476, 16'd31042, 16'd26968, 16'd29999, 16'd64283, 16'd54163, 16'd53481, 16'd44898, 16'd63652, 16'd54477, 16'd35294, 16'd18167, 16'd20647, 16'd29725, 16'd53385, 16'd46680, 16'd38474, 16'd55943, 16'd55313});
	test_expansion(128'h83f8c5690e1475c81a4f6f393353c575, {16'd19560, 16'd6423, 16'd64624, 16'd36460, 16'd23213, 16'd2346, 16'd32473, 16'd14954, 16'd47145, 16'd16545, 16'd34830, 16'd32714, 16'd739, 16'd57774, 16'd24212, 16'd4859, 16'd22373, 16'd60659, 16'd65480, 16'd1250, 16'd9658, 16'd40645, 16'd47067, 16'd36637, 16'd36676, 16'd16270});
	test_expansion(128'hbe052c9c9dffa309cc2f2555ddf7ddd3, {16'd38398, 16'd9902, 16'd13803, 16'd5545, 16'd9069, 16'd54477, 16'd59483, 16'd19955, 16'd52474, 16'd31852, 16'd7540, 16'd23020, 16'd25091, 16'd11505, 16'd35929, 16'd62479, 16'd9378, 16'd55612, 16'd41613, 16'd15972, 16'd14058, 16'd30365, 16'd42782, 16'd27181, 16'd62671, 16'd56778});
	test_expansion(128'h5f86f3107fa661273d2d8257b9788eb8, {16'd8849, 16'd30270, 16'd3001, 16'd28567, 16'd36748, 16'd60666, 16'd59920, 16'd29759, 16'd56806, 16'd4513, 16'd46679, 16'd21003, 16'd6932, 16'd39105, 16'd27364, 16'd28275, 16'd30526, 16'd61109, 16'd27561, 16'd46886, 16'd58360, 16'd25545, 16'd64226, 16'd40797, 16'd44324, 16'd51803});
	test_expansion(128'h38331515e86cd1d92932515c60aa2599, {16'd9692, 16'd48092, 16'd37971, 16'd13510, 16'd14632, 16'd65247, 16'd18644, 16'd8274, 16'd12833, 16'd49828, 16'd29518, 16'd22159, 16'd47409, 16'd46212, 16'd7903, 16'd11265, 16'd15165, 16'd30550, 16'd25566, 16'd39290, 16'd39520, 16'd16002, 16'd46231, 16'd14816, 16'd2036, 16'd41179});
	test_expansion(128'h22e28c6f16993f7009a0f2986ce7904f, {16'd60116, 16'd52492, 16'd45389, 16'd61917, 16'd53320, 16'd53213, 16'd30292, 16'd28365, 16'd49763, 16'd62359, 16'd17456, 16'd30657, 16'd40735, 16'd53443, 16'd33903, 16'd22712, 16'd10910, 16'd40225, 16'd33186, 16'd58289, 16'd8201, 16'd40133, 16'd14962, 16'd12776, 16'd13728, 16'd30439});
	test_expansion(128'h5c64d14907043a7dd1c71f35851eb5a8, {16'd45890, 16'd11331, 16'd3352, 16'd57732, 16'd36403, 16'd1936, 16'd49691, 16'd7501, 16'd49826, 16'd16798, 16'd42882, 16'd65525, 16'd12986, 16'd9205, 16'd32737, 16'd190, 16'd52035, 16'd14576, 16'd2346, 16'd41753, 16'd58600, 16'd7214, 16'd50622, 16'd46931, 16'd6813, 16'd29573});
	test_expansion(128'he922e829c2c99b0955f93083beacd59e, {16'd5742, 16'd57423, 16'd44993, 16'd26891, 16'd15277, 16'd9395, 16'd31391, 16'd56188, 16'd43718, 16'd16871, 16'd39319, 16'd52661, 16'd56852, 16'd7809, 16'd41872, 16'd12047, 16'd47762, 16'd27151, 16'd31775, 16'd37762, 16'd11524, 16'd36776, 16'd8133, 16'd27497, 16'd53594, 16'd47990});
	test_expansion(128'h9f5aafbeb6572cfba63aa10cc50003b6, {16'd63689, 16'd22963, 16'd28555, 16'd50754, 16'd3471, 16'd39063, 16'd1301, 16'd31661, 16'd26283, 16'd30087, 16'd15929, 16'd54234, 16'd18389, 16'd974, 16'd58021, 16'd14946, 16'd22293, 16'd45294, 16'd9287, 16'd15945, 16'd51691, 16'd11247, 16'd32110, 16'd14022, 16'd12789, 16'd14844});
	test_expansion(128'hecff9f2553434b8fe0629a596c16b503, {16'd15560, 16'd5244, 16'd52145, 16'd15696, 16'd17754, 16'd37942, 16'd43805, 16'd63658, 16'd61819, 16'd50359, 16'd55824, 16'd17312, 16'd4296, 16'd34471, 16'd35090, 16'd36530, 16'd6908, 16'd9007, 16'd32962, 16'd48948, 16'd35884, 16'd30972, 16'd41748, 16'd38543, 16'd32034, 16'd26865});
	test_expansion(128'h9dcab53da207710fc44d71c8adbc163f, {16'd23409, 16'd28802, 16'd10682, 16'd19430, 16'd56873, 16'd41542, 16'd14849, 16'd55517, 16'd3069, 16'd17986, 16'd27172, 16'd53628, 16'd9437, 16'd54600, 16'd43115, 16'd38447, 16'd11012, 16'd14930, 16'd59327, 16'd13931, 16'd28130, 16'd59459, 16'd44757, 16'd19111, 16'd6317, 16'd57565});
	test_expansion(128'h8b4a586e38107360d72e6c46a7ef9a9a, {16'd59925, 16'd42465, 16'd25157, 16'd50403, 16'd53338, 16'd50245, 16'd45488, 16'd36515, 16'd53592, 16'd32577, 16'd33911, 16'd62509, 16'd39625, 16'd24089, 16'd20700, 16'd38420, 16'd200, 16'd44100, 16'd20191, 16'd25285, 16'd50562, 16'd52094, 16'd29079, 16'd17686, 16'd49210, 16'd16765});
	test_expansion(128'h882aaea4c55f65ece80e131e8cca49e0, {16'd3052, 16'd50381, 16'd10694, 16'd29928, 16'd23022, 16'd20239, 16'd35435, 16'd58233, 16'd48189, 16'd65108, 16'd6546, 16'd25997, 16'd15846, 16'd60336, 16'd47233, 16'd3504, 16'd41673, 16'd1460, 16'd22294, 16'd653, 16'd14715, 16'd25854, 16'd38324, 16'd28109, 16'd44362, 16'd55808});
	test_expansion(128'hdb8cded5b0f5afa3323f0329ed35d434, {16'd42539, 16'd3592, 16'd3104, 16'd35001, 16'd44190, 16'd5735, 16'd61175, 16'd5556, 16'd49544, 16'd10754, 16'd60422, 16'd10636, 16'd42514, 16'd48408, 16'd4035, 16'd42170, 16'd53744, 16'd27134, 16'd39163, 16'd6826, 16'd18404, 16'd34361, 16'd5820, 16'd46522, 16'd11897, 16'd39085});
	test_expansion(128'h4593c48a9478722b37bedc60f9956b5e, {16'd61560, 16'd3929, 16'd42977, 16'd16918, 16'd65431, 16'd63303, 16'd56924, 16'd34992, 16'd8696, 16'd60781, 16'd13862, 16'd14121, 16'd40307, 16'd36675, 16'd8210, 16'd187, 16'd20057, 16'd40443, 16'd27411, 16'd14756, 16'd36331, 16'd43546, 16'd57839, 16'd54594, 16'd58820, 16'd7483});
	test_expansion(128'hc7d939a172c2efef2a7b3ab2a54ca63a, {16'd7506, 16'd34084, 16'd63063, 16'd38941, 16'd8013, 16'd28003, 16'd59790, 16'd62309, 16'd58288, 16'd31688, 16'd37435, 16'd13807, 16'd49906, 16'd18978, 16'd56559, 16'd17716, 16'd54018, 16'd2052, 16'd10916, 16'd56092, 16'd59055, 16'd7085, 16'd27741, 16'd10128, 16'd13098, 16'd51561});
	test_expansion(128'h33b8e553bc5d5d7a04339e0f99a766c6, {16'd49487, 16'd19382, 16'd7356, 16'd21629, 16'd33019, 16'd27820, 16'd60523, 16'd23379, 16'd10239, 16'd31240, 16'd29766, 16'd30791, 16'd52129, 16'd36082, 16'd56075, 16'd33424, 16'd6829, 16'd3381, 16'd59078, 16'd17156, 16'd45183, 16'd56702, 16'd55994, 16'd31138, 16'd23748, 16'd22506});
	test_expansion(128'hfd815fdc38c77192c984df09ee7be043, {16'd20536, 16'd567, 16'd11701, 16'd61481, 16'd61389, 16'd14793, 16'd6150, 16'd51346, 16'd36346, 16'd54879, 16'd10913, 16'd40993, 16'd47499, 16'd4311, 16'd39437, 16'd41260, 16'd16206, 16'd5425, 16'd5661, 16'd2829, 16'd49722, 16'd51368, 16'd29041, 16'd15739, 16'd6973, 16'd47852});
	test_expansion(128'h11e75372358291735c2c46c42d410ea3, {16'd57979, 16'd15447, 16'd21118, 16'd41926, 16'd63677, 16'd15307, 16'd44122, 16'd37175, 16'd28936, 16'd30215, 16'd39309, 16'd24656, 16'd17688, 16'd40887, 16'd22466, 16'd47639, 16'd53155, 16'd61766, 16'd19753, 16'd17574, 16'd23416, 16'd53193, 16'd60348, 16'd61809, 16'd38144, 16'd60470});
	test_expansion(128'ha75aa81b301e986929cfce2087ed2157, {16'd3178, 16'd40870, 16'd46091, 16'd58706, 16'd8424, 16'd59754, 16'd36546, 16'd22149, 16'd44946, 16'd8154, 16'd9044, 16'd32770, 16'd55397, 16'd63560, 16'd45814, 16'd49483, 16'd65396, 16'd19448, 16'd49772, 16'd42272, 16'd11726, 16'd42297, 16'd1854, 16'd58480, 16'd61834, 16'd38472});
	test_expansion(128'h1364c1943c1ef1f5d76509353d30bb9f, {16'd24988, 16'd5796, 16'd61120, 16'd64108, 16'd14744, 16'd56463, 16'd19348, 16'd63402, 16'd50239, 16'd31443, 16'd10113, 16'd2141, 16'd54822, 16'd35977, 16'd51966, 16'd64360, 16'd4552, 16'd27903, 16'd12596, 16'd15232, 16'd40639, 16'd26352, 16'd27946, 16'd49203, 16'd62884, 16'd36825});
	test_expansion(128'h7039487c55b0d8f2e119e1c7c6397729, {16'd31116, 16'd28960, 16'd37950, 16'd57103, 16'd12688, 16'd22080, 16'd64630, 16'd32920, 16'd4907, 16'd45746, 16'd30484, 16'd11157, 16'd17647, 16'd31308, 16'd44282, 16'd20156, 16'd13539, 16'd63131, 16'd52685, 16'd41966, 16'd44435, 16'd32383, 16'd21978, 16'd11397, 16'd36187, 16'd11723});
	test_expansion(128'h0d5e079d86bd33ce563ce4353be54807, {16'd18843, 16'd14497, 16'd14864, 16'd16470, 16'd7923, 16'd59026, 16'd10340, 16'd35024, 16'd3803, 16'd55111, 16'd64153, 16'd26419, 16'd40681, 16'd47268, 16'd18204, 16'd1314, 16'd16293, 16'd46129, 16'd44454, 16'd25815, 16'd56121, 16'd30637, 16'd19496, 16'd6731, 16'd31282, 16'd43130});
	test_expansion(128'h5c56636b6b49b8daa14250fbf5dfe9d3, {16'd35763, 16'd2864, 16'd61416, 16'd10971, 16'd45974, 16'd28228, 16'd7819, 16'd16449, 16'd57062, 16'd52225, 16'd27810, 16'd52574, 16'd30631, 16'd17816, 16'd22172, 16'd62812, 16'd20140, 16'd62428, 16'd2799, 16'd52644, 16'd35186, 16'd7271, 16'd49779, 16'd39215, 16'd63813, 16'd55149});
	test_expansion(128'h1c110b47c05cd67152874ed46d7fca76, {16'd21457, 16'd16426, 16'd38818, 16'd62643, 16'd64437, 16'd12861, 16'd8672, 16'd25361, 16'd53682, 16'd15327, 16'd45076, 16'd8168, 16'd2483, 16'd9173, 16'd25743, 16'd17638, 16'd54462, 16'd27081, 16'd46697, 16'd19613, 16'd53348, 16'd23425, 16'd44395, 16'd63562, 16'd58522, 16'd47852});
	test_expansion(128'h3a75fd3bae363162ee3c65983f1214ef, {16'd12490, 16'd53660, 16'd8661, 16'd14405, 16'd52430, 16'd22220, 16'd62161, 16'd20367, 16'd20347, 16'd58606, 16'd25124, 16'd38178, 16'd19949, 16'd14306, 16'd17350, 16'd9284, 16'd19058, 16'd31401, 16'd9456, 16'd49144, 16'd18311, 16'd3696, 16'd40859, 16'd63119, 16'd16786, 16'd34277});
	test_expansion(128'he59d031b2dd44bb4fae3ca6ad03bbd86, {16'd12513, 16'd8026, 16'd1463, 16'd7312, 16'd20439, 16'd57126, 16'd23555, 16'd27991, 16'd13391, 16'd102, 16'd61988, 16'd43043, 16'd33021, 16'd35885, 16'd4910, 16'd40199, 16'd28449, 16'd46818, 16'd7312, 16'd12701, 16'd27177, 16'd41778, 16'd61824, 16'd37495, 16'd49772, 16'd64606});
	test_expansion(128'h65af145e4f7d5485b9a774b102e053cc, {16'd45863, 16'd950, 16'd20944, 16'd46283, 16'd19609, 16'd64235, 16'd40760, 16'd64921, 16'd45976, 16'd13675, 16'd34755, 16'd64954, 16'd2021, 16'd32903, 16'd33424, 16'd10827, 16'd49401, 16'd22676, 16'd60850, 16'd11280, 16'd22250, 16'd3805, 16'd40686, 16'd37002, 16'd48009, 16'd59746});
	test_expansion(128'h38fd32a4abd6214434d7d370929e994b, {16'd4230, 16'd59562, 16'd53079, 16'd57730, 16'd15108, 16'd42025, 16'd39449, 16'd10863, 16'd60050, 16'd25268, 16'd49046, 16'd17675, 16'd15161, 16'd56327, 16'd40591, 16'd29698, 16'd401, 16'd6166, 16'd58324, 16'd61026, 16'd58440, 16'd47725, 16'd10751, 16'd28384, 16'd24958, 16'd45804});
	test_expansion(128'ha943e03fda6ddd951d7d580f2b833a18, {16'd46115, 16'd16990, 16'd26784, 16'd34811, 16'd52310, 16'd29649, 16'd42851, 16'd31314, 16'd5132, 16'd56937, 16'd60448, 16'd42722, 16'd39136, 16'd44922, 16'd9604, 16'd40880, 16'd56817, 16'd6979, 16'd22189, 16'd14065, 16'd61170, 16'd32284, 16'd58423, 16'd56700, 16'd50541, 16'd15050});
	test_expansion(128'hf8c44b98d22d50117b06fb540a720aca, {16'd1774, 16'd15450, 16'd41827, 16'd38676, 16'd8043, 16'd50132, 16'd35683, 16'd54816, 16'd8421, 16'd51922, 16'd22366, 16'd24870, 16'd12454, 16'd54749, 16'd64786, 16'd16660, 16'd13543, 16'd21103, 16'd45052, 16'd9742, 16'd28911, 16'd6947, 16'd36211, 16'd49061, 16'd17866, 16'd48088});
	test_expansion(128'hf9f56c2fd6678a00160726e753cddb0f, {16'd33516, 16'd1585, 16'd12095, 16'd19539, 16'd21550, 16'd42999, 16'd49018, 16'd20037, 16'd19593, 16'd573, 16'd37904, 16'd36686, 16'd50832, 16'd1008, 16'd740, 16'd61894, 16'd12625, 16'd16578, 16'd41729, 16'd49790, 16'd25129, 16'd28475, 16'd43068, 16'd62728, 16'd24172, 16'd29866});
	test_expansion(128'h4a0edb9b6da5efc5ed95e95412099363, {16'd50608, 16'd55250, 16'd34045, 16'd53012, 16'd23082, 16'd25525, 16'd32287, 16'd51914, 16'd48839, 16'd11765, 16'd14809, 16'd47992, 16'd32437, 16'd20591, 16'd35475, 16'd23170, 16'd12744, 16'd14508, 16'd11670, 16'd45784, 16'd8351, 16'd7112, 16'd34766, 16'd26850, 16'd7584, 16'd62468});
	test_expansion(128'h7a2a540918b6f3a1461df435241766bf, {16'd43636, 16'd44479, 16'd9095, 16'd15709, 16'd14802, 16'd10699, 16'd12820, 16'd15916, 16'd35974, 16'd25012, 16'd52840, 16'd47739, 16'd24413, 16'd43844, 16'd18836, 16'd40328, 16'd33561, 16'd36243, 16'd36009, 16'd33449, 16'd45344, 16'd39680, 16'd36493, 16'd31868, 16'd33640, 16'd39073});
	test_expansion(128'h8ba02bc4ffc27bf642ed73b636a44349, {16'd60649, 16'd57279, 16'd57735, 16'd5796, 16'd3609, 16'd25830, 16'd3164, 16'd40492, 16'd7359, 16'd16579, 16'd13801, 16'd7892, 16'd24843, 16'd34771, 16'd40973, 16'd9798, 16'd15683, 16'd21961, 16'd38972, 16'd34538, 16'd30483, 16'd5523, 16'd61492, 16'd13153, 16'd432, 16'd5382});
	test_expansion(128'h38edff4eec8c85447ac243ae5b286dcf, {16'd29297, 16'd41464, 16'd46825, 16'd16673, 16'd8087, 16'd13952, 16'd3180, 16'd58775, 16'd13958, 16'd50392, 16'd5491, 16'd857, 16'd61877, 16'd21174, 16'd28366, 16'd63030, 16'd39866, 16'd46231, 16'd54079, 16'd8301, 16'd40608, 16'd4905, 16'd52769, 16'd10699, 16'd50098, 16'd59433});
	test_expansion(128'h288ce1e9ea8cc14f02760b5e63041cd9, {16'd41956, 16'd8504, 16'd26721, 16'd62085, 16'd29294, 16'd2232, 16'd20896, 16'd43083, 16'd20786, 16'd46559, 16'd27391, 16'd9358, 16'd50534, 16'd27155, 16'd61011, 16'd34477, 16'd33243, 16'd43978, 16'd53814, 16'd1173, 16'd43716, 16'd43392, 16'd56824, 16'd29396, 16'd61318, 16'd27881});
	test_expansion(128'h90a2845d457aac3898e7e0eb0bf16c21, {16'd13038, 16'd42102, 16'd33092, 16'd20507, 16'd40687, 16'd43727, 16'd111, 16'd48558, 16'd8589, 16'd520, 16'd48989, 16'd46657, 16'd38092, 16'd11679, 16'd2039, 16'd16685, 16'd37097, 16'd59358, 16'd12207, 16'd52260, 16'd64086, 16'd6185, 16'd25503, 16'd13598, 16'd58266, 16'd34308});
	test_expansion(128'h8c319d73e0aeaf9eb1e9bd0f8c744bb9, {16'd30084, 16'd61421, 16'd20953, 16'd29726, 16'd5279, 16'd920, 16'd2051, 16'd15312, 16'd49831, 16'd19684, 16'd34453, 16'd35047, 16'd47235, 16'd42748, 16'd43287, 16'd16360, 16'd6897, 16'd50763, 16'd37274, 16'd22334, 16'd24840, 16'd27702, 16'd42850, 16'd42839, 16'd36873, 16'd55606});
	test_expansion(128'h16cb70ae594af3d13acdcffca0363df2, {16'd46258, 16'd50331, 16'd9556, 16'd50958, 16'd23014, 16'd3818, 16'd60340, 16'd33841, 16'd57246, 16'd60698, 16'd32948, 16'd5905, 16'd46592, 16'd48994, 16'd53839, 16'd37776, 16'd34343, 16'd13715, 16'd1258, 16'd46123, 16'd5315, 16'd18160, 16'd6917, 16'd37812, 16'd2356, 16'd2710});
	test_expansion(128'hae48deb012a8d8e607d73f77cca0542c, {16'd43937, 16'd61600, 16'd54828, 16'd9657, 16'd36276, 16'd33498, 16'd50680, 16'd48459, 16'd12140, 16'd1135, 16'd64171, 16'd48687, 16'd1528, 16'd4957, 16'd58926, 16'd33014, 16'd46709, 16'd42588, 16'd14112, 16'd3635, 16'd15491, 16'd8422, 16'd29104, 16'd33805, 16'd42199, 16'd47906});
	test_expansion(128'h11129136573072876cb036e19ed308c9, {16'd3370, 16'd8898, 16'd28134, 16'd45747, 16'd40603, 16'd2350, 16'd50779, 16'd53479, 16'd48958, 16'd38073, 16'd20725, 16'd10021, 16'd19740, 16'd46292, 16'd18937, 16'd24014, 16'd2297, 16'd38844, 16'd1722, 16'd59974, 16'd23496, 16'd8613, 16'd40957, 16'd5631, 16'd12188, 16'd51405});
	test_expansion(128'h012aeca6430b9741e9b1741a62637c42, {16'd4548, 16'd27667, 16'd10423, 16'd360, 16'd30481, 16'd10319, 16'd4999, 16'd24873, 16'd33826, 16'd40069, 16'd24394, 16'd45257, 16'd21801, 16'd37371, 16'd27409, 16'd33863, 16'd34672, 16'd63902, 16'd45718, 16'd50536, 16'd23654, 16'd56493, 16'd31866, 16'd10500, 16'd6491, 16'd37801});
	test_expansion(128'hd95c5b19e9b2f225212b3c31616504b4, {16'd13651, 16'd17813, 16'd20051, 16'd37740, 16'd35944, 16'd35821, 16'd4884, 16'd58806, 16'd63464, 16'd53826, 16'd13033, 16'd40389, 16'd47868, 16'd30616, 16'd56726, 16'd63390, 16'd63129, 16'd64752, 16'd24490, 16'd5000, 16'd7416, 16'd35134, 16'd51941, 16'd51257, 16'd2254, 16'd16273});
	test_expansion(128'hf2427bfaef323f0749e683682804da55, {16'd52908, 16'd56921, 16'd30488, 16'd28351, 16'd22813, 16'd39521, 16'd45695, 16'd19309, 16'd49249, 16'd58540, 16'd22311, 16'd17626, 16'd9627, 16'd53044, 16'd17327, 16'd63428, 16'd8100, 16'd19126, 16'd17995, 16'd61227, 16'd21603, 16'd30401, 16'd8678, 16'd11099, 16'd33535, 16'd28871});
	test_expansion(128'hfc537ec0ab167e4298e2db1adce84cee, {16'd57605, 16'd63715, 16'd27729, 16'd8720, 16'd18096, 16'd11614, 16'd23023, 16'd24983, 16'd48515, 16'd44531, 16'd9152, 16'd31526, 16'd56369, 16'd45041, 16'd46721, 16'd28797, 16'd4395, 16'd46360, 16'd30913, 16'd50512, 16'd7938, 16'd55539, 16'd23220, 16'd1277, 16'd9098, 16'd48506});
	test_expansion(128'hdf6655080688d6672c1563bcde69950b, {16'd16873, 16'd1981, 16'd50117, 16'd9169, 16'd12617, 16'd36824, 16'd28782, 16'd16615, 16'd46747, 16'd55696, 16'd51698, 16'd54858, 16'd62195, 16'd60344, 16'd25544, 16'd62337, 16'd22908, 16'd28294, 16'd31653, 16'd21812, 16'd29498, 16'd54147, 16'd23844, 16'd24927, 16'd32573, 16'd1396});
	test_expansion(128'h4c55d4e791b020aad0ced3ebef8a62ce, {16'd29980, 16'd27820, 16'd44622, 16'd50680, 16'd24674, 16'd20575, 16'd4628, 16'd41290, 16'd31395, 16'd2164, 16'd52579, 16'd27531, 16'd65287, 16'd36060, 16'd51371, 16'd18011, 16'd59864, 16'd35771, 16'd13257, 16'd14720, 16'd28411, 16'd37164, 16'd31309, 16'd18955, 16'd3808, 16'd28570});
	test_expansion(128'h753ba536582e53c4b88abb97f544d1cd, {16'd55755, 16'd38037, 16'd54245, 16'd64267, 16'd27519, 16'd8557, 16'd35566, 16'd35671, 16'd63192, 16'd9519, 16'd6045, 16'd57521, 16'd22918, 16'd48724, 16'd16890, 16'd24993, 16'd12047, 16'd594, 16'd47553, 16'd43888, 16'd19943, 16'd54403, 16'd63405, 16'd43117, 16'd3345, 16'd24712});
	test_expansion(128'hd9d4202c2522049916951412fc855a32, {16'd16608, 16'd44851, 16'd53425, 16'd65535, 16'd15107, 16'd47910, 16'd2277, 16'd11675, 16'd38753, 16'd12101, 16'd64038, 16'd26596, 16'd54415, 16'd12208, 16'd15868, 16'd3102, 16'd46329, 16'd1147, 16'd58133, 16'd60223, 16'd48262, 16'd31942, 16'd5411, 16'd17468, 16'd35027, 16'd44059});
	test_expansion(128'h22cb0c35b5b3e0bca643716a4a4c77e6, {16'd11106, 16'd59295, 16'd29824, 16'd13932, 16'd19813, 16'd31068, 16'd4089, 16'd42898, 16'd64204, 16'd30642, 16'd33269, 16'd25860, 16'd35576, 16'd57287, 16'd60776, 16'd33441, 16'd9528, 16'd50316, 16'd25070, 16'd25346, 16'd26250, 16'd52784, 16'd10304, 16'd24038, 16'd2971, 16'd55473});
	test_expansion(128'ha8d4aa0b20d2da5f81c8474ad0181fc5, {16'd52253, 16'd37559, 16'd53494, 16'd33753, 16'd39560, 16'd3450, 16'd42534, 16'd15760, 16'd16747, 16'd29219, 16'd37534, 16'd57326, 16'd60724, 16'd8697, 16'd58767, 16'd22628, 16'd42190, 16'd37098, 16'd35272, 16'd41631, 16'd21011, 16'd28557, 16'd47335, 16'd10013, 16'd44898, 16'd25022});
	test_expansion(128'h2c7b1e8efc357fe496160521279be25d, {16'd13547, 16'd22721, 16'd55464, 16'd65442, 16'd32540, 16'd6415, 16'd2522, 16'd26504, 16'd5982, 16'd7683, 16'd28230, 16'd63922, 16'd13595, 16'd32929, 16'd24596, 16'd49030, 16'd17533, 16'd59536, 16'd2216, 16'd39181, 16'd41955, 16'd27686, 16'd54704, 16'd2704, 16'd26145, 16'd34077});
	test_expansion(128'h4d42999916efad95db61980ed69adb5e, {16'd36002, 16'd15331, 16'd27016, 16'd35168, 16'd46309, 16'd28935, 16'd7166, 16'd31881, 16'd16226, 16'd3133, 16'd20171, 16'd9608, 16'd38221, 16'd15540, 16'd55293, 16'd45565, 16'd29412, 16'd13974, 16'd21258, 16'd47450, 16'd53673, 16'd59328, 16'd55094, 16'd3472, 16'd2575, 16'd41417});
	test_expansion(128'hd11948bb0894e928e99a67fe8da9ffb4, {16'd31138, 16'd45379, 16'd49185, 16'd19137, 16'd15425, 16'd9253, 16'd41362, 16'd61710, 16'd55497, 16'd14280, 16'd28580, 16'd9276, 16'd29973, 16'd57708, 16'd52250, 16'd1614, 16'd58159, 16'd45822, 16'd4934, 16'd50556, 16'd49427, 16'd46577, 16'd54897, 16'd26195, 16'd17654, 16'd45159});
	test_expansion(128'h0f1fa510a9eb47bf16ee41adadb16255, {16'd61019, 16'd21295, 16'd53153, 16'd12753, 16'd50608, 16'd33395, 16'd11452, 16'd6151, 16'd30615, 16'd27237, 16'd15680, 16'd8459, 16'd52443, 16'd57002, 16'd48060, 16'd56045, 16'd12170, 16'd23426, 16'd57283, 16'd29699, 16'd24799, 16'd36098, 16'd222, 16'd16834, 16'd46700, 16'd50347});
	test_expansion(128'hfce6de6b5bba9cb2e226a3e87d8d7047, {16'd61550, 16'd26698, 16'd49381, 16'd21565, 16'd42684, 16'd48742, 16'd2881, 16'd27053, 16'd33360, 16'd30020, 16'd62042, 16'd42590, 16'd24085, 16'd24211, 16'd904, 16'd24746, 16'd53152, 16'd13052, 16'd33478, 16'd10870, 16'd53043, 16'd35779, 16'd75, 16'd30006, 16'd54025, 16'd11772});
	test_expansion(128'h196ca1ddaf063e2a402d5839c202156b, {16'd38130, 16'd41546, 16'd24981, 16'd56954, 16'd20097, 16'd58523, 16'd34233, 16'd53146, 16'd55415, 16'd65279, 16'd12996, 16'd9061, 16'd1431, 16'd16458, 16'd23556, 16'd24254, 16'd37231, 16'd6589, 16'd56281, 16'd12583, 16'd20747, 16'd7735, 16'd18156, 16'd30088, 16'd51150, 16'd43412});
	test_expansion(128'h71e8529cf67ab73b0301a2ac2993a03b, {16'd38595, 16'd63487, 16'd1888, 16'd4061, 16'd30548, 16'd25361, 16'd10519, 16'd64411, 16'd3446, 16'd48182, 16'd15315, 16'd26354, 16'd3885, 16'd25115, 16'd29520, 16'd54164, 16'd55952, 16'd53417, 16'd6664, 16'd64828, 16'd28408, 16'd36966, 16'd5670, 16'd58356, 16'd14252, 16'd17258});
	test_expansion(128'h21ec26e1983872e243aa849d2159b6f4, {16'd18853, 16'd63880, 16'd2608, 16'd3822, 16'd41811, 16'd62645, 16'd51792, 16'd44342, 16'd29226, 16'd27765, 16'd6359, 16'd14623, 16'd28628, 16'd12689, 16'd39860, 16'd59416, 16'd21503, 16'd38465, 16'd2884, 16'd54337, 16'd2511, 16'd38751, 16'd56942, 16'd45890, 16'd44232, 16'd20374});
	test_expansion(128'h764f3207ad87265ee30214d55812165e, {16'd55764, 16'd57248, 16'd44905, 16'd28417, 16'd53231, 16'd33669, 16'd823, 16'd63594, 16'd41575, 16'd21048, 16'd59365, 16'd27558, 16'd63966, 16'd42674, 16'd20253, 16'd62099, 16'd18361, 16'd35576, 16'd56647, 16'd39176, 16'd11445, 16'd11751, 16'd1319, 16'd40591, 16'd17935, 16'd47405});
	test_expansion(128'ha538981d9e62ea476db7cfb0e65d601c, {16'd24126, 16'd49501, 16'd26874, 16'd2804, 16'd37738, 16'd39434, 16'd49331, 16'd63850, 16'd37646, 16'd1607, 16'd23019, 16'd25336, 16'd4642, 16'd20936, 16'd25087, 16'd37194, 16'd3847, 16'd45285, 16'd2732, 16'd21783, 16'd65275, 16'd58425, 16'd5462, 16'd59075, 16'd54342, 16'd60541});
	test_expansion(128'h1a5f098b0731743c48f2bd7dc33d4687, {16'd55721, 16'd36668, 16'd20982, 16'd51657, 16'd1149, 16'd58027, 16'd49581, 16'd62224, 16'd30469, 16'd4806, 16'd2790, 16'd38852, 16'd54734, 16'd22552, 16'd14846, 16'd59602, 16'd22296, 16'd38873, 16'd5232, 16'd3484, 16'd37345, 16'd50262, 16'd6985, 16'd28691, 16'd22053, 16'd23768});
	test_expansion(128'he83c208b65204b6dff0e0611972d815c, {16'd37473, 16'd7115, 16'd48371, 16'd37345, 16'd37221, 16'd38011, 16'd38125, 16'd33334, 16'd48425, 16'd51623, 16'd58259, 16'd20991, 16'd19640, 16'd35680, 16'd63245, 16'd37035, 16'd56108, 16'd7804, 16'd59688, 16'd33962, 16'd22619, 16'd11477, 16'd2992, 16'd45957, 16'd24585, 16'd50166});
	test_expansion(128'h3c7970969c68e7bcf1a921d65150391e, {16'd32777, 16'd60846, 16'd21431, 16'd5068, 16'd61823, 16'd58657, 16'd22830, 16'd47467, 16'd34568, 16'd45606, 16'd13455, 16'd63461, 16'd29540, 16'd52560, 16'd32473, 16'd5817, 16'd43622, 16'd44410, 16'd35844, 16'd10838, 16'd43797, 16'd60123, 16'd3324, 16'd23257, 16'd25486, 16'd6451});
	test_expansion(128'hdb3beaa5578742e05f466db03420403b, {16'd19119, 16'd37296, 16'd5726, 16'd12714, 16'd5949, 16'd27109, 16'd25482, 16'd5014, 16'd35741, 16'd13755, 16'd47520, 16'd37038, 16'd39010, 16'd26121, 16'd63182, 16'd15988, 16'd8267, 16'd42240, 16'd39123, 16'd29418, 16'd2302, 16'd32380, 16'd61691, 16'd320, 16'd8349, 16'd36836});
	test_expansion(128'h0e25dd631bd9acc7330d5706311ae371, {16'd45763, 16'd23335, 16'd61429, 16'd29562, 16'd24210, 16'd2381, 16'd51666, 16'd47021, 16'd21786, 16'd5931, 16'd52521, 16'd55846, 16'd32033, 16'd19213, 16'd45325, 16'd38663, 16'd11633, 16'd49911, 16'd41494, 16'd37047, 16'd64656, 16'd32518, 16'd57201, 16'd27937, 16'd6932, 16'd50689});
	test_expansion(128'h1eb183f474834a34f6f4b43d7c0ad179, {16'd54423, 16'd805, 16'd4700, 16'd54914, 16'd59748, 16'd55704, 16'd3064, 16'd58432, 16'd34748, 16'd51598, 16'd9072, 16'd37147, 16'd8908, 16'd32912, 16'd26808, 16'd62688, 16'd18044, 16'd26182, 16'd6387, 16'd40464, 16'd52570, 16'd4180, 16'd30740, 16'd5960, 16'd28058, 16'd42361});
	test_expansion(128'hd3c0cb7b1131e1bd703cd786331d27d8, {16'd64284, 16'd55118, 16'd18668, 16'd18699, 16'd36944, 16'd25420, 16'd33740, 16'd57539, 16'd27482, 16'd34226, 16'd61426, 16'd9343, 16'd30136, 16'd40910, 16'd23365, 16'd52409, 16'd16356, 16'd21669, 16'd17064, 16'd54885, 16'd53430, 16'd63203, 16'd25900, 16'd64934, 16'd38303, 16'd32637});
	test_expansion(128'h4a440e5f24d2169a480229aa9e05e94a, {16'd57047, 16'd43236, 16'd69, 16'd14990, 16'd5708, 16'd37273, 16'd37795, 16'd4823, 16'd40826, 16'd39012, 16'd26230, 16'd20316, 16'd51191, 16'd48884, 16'd12903, 16'd33319, 16'd15274, 16'd10743, 16'd59226, 16'd12638, 16'd33793, 16'd25449, 16'd13475, 16'd56958, 16'd27848, 16'd34203});
	test_expansion(128'h281de745421ad3bbe02e128aa560f273, {16'd21469, 16'd40664, 16'd8512, 16'd32716, 16'd16892, 16'd64821, 16'd65149, 16'd2824, 16'd57646, 16'd9297, 16'd18197, 16'd53066, 16'd29400, 16'd17082, 16'd31890, 16'd22427, 16'd60391, 16'd55204, 16'd27553, 16'd45195, 16'd59227, 16'd21778, 16'd30572, 16'd56829, 16'd31519, 16'd4832});
	test_expansion(128'hc773aa20738ae443e97d5281cc8cd82c, {16'd54018, 16'd50274, 16'd35509, 16'd42916, 16'd38739, 16'd36051, 16'd28262, 16'd16231, 16'd47957, 16'd631, 16'd59394, 16'd32515, 16'd27131, 16'd49607, 16'd4226, 16'd59112, 16'd39878, 16'd51139, 16'd27521, 16'd44674, 16'd63396, 16'd29845, 16'd44264, 16'd10142, 16'd55713, 16'd41247});
	test_expansion(128'h11ccd9e5ec04d3b54ca23f93d709c7c6, {16'd44529, 16'd18604, 16'd65361, 16'd11082, 16'd57190, 16'd5215, 16'd63683, 16'd23643, 16'd55136, 16'd27760, 16'd15151, 16'd14382, 16'd52605, 16'd38199, 16'd24237, 16'd45968, 16'd54365, 16'd58304, 16'd50528, 16'd53318, 16'd46643, 16'd30252, 16'd25348, 16'd20390, 16'd27831, 16'd41871});
	test_expansion(128'hbe8dd61b0e053b3f35178544ad883965, {16'd62176, 16'd51533, 16'd56459, 16'd53104, 16'd29029, 16'd13013, 16'd9427, 16'd52574, 16'd33851, 16'd37270, 16'd9726, 16'd4977, 16'd2404, 16'd8956, 16'd5667, 16'd63268, 16'd64641, 16'd37895, 16'd40359, 16'd64039, 16'd51099, 16'd62615, 16'd60018, 16'd49788, 16'd39912, 16'd30400});
	test_expansion(128'hb6e149036c651752bc9cbae4cc394e52, {16'd4694, 16'd3801, 16'd7843, 16'd33996, 16'd4516, 16'd44127, 16'd17604, 16'd43186, 16'd50579, 16'd51586, 16'd5271, 16'd23588, 16'd65044, 16'd25729, 16'd7665, 16'd53680, 16'd61901, 16'd32933, 16'd9574, 16'd2523, 16'd53026, 16'd33456, 16'd48539, 16'd20171, 16'd37093, 16'd26520});
	test_expansion(128'he0874c7818d2b2e7e66c6ac724ef6f2d, {16'd59635, 16'd53639, 16'd14434, 16'd59519, 16'd27238, 16'd4242, 16'd4130, 16'd39648, 16'd22066, 16'd1392, 16'd42853, 16'd51891, 16'd7884, 16'd21811, 16'd44785, 16'd37039, 16'd34424, 16'd4473, 16'd47699, 16'd20750, 16'd48749, 16'd22834, 16'd48776, 16'd64140, 16'd30657, 16'd19714});
	test_expansion(128'h3b6bd4361e4161ab011a61f364c1dbac, {16'd36883, 16'd59226, 16'd62550, 16'd44109, 16'd63278, 16'd63157, 16'd50978, 16'd55480, 16'd40567, 16'd57117, 16'd58261, 16'd1570, 16'd26573, 16'd5091, 16'd60232, 16'd30243, 16'd30192, 16'd5335, 16'd32188, 16'd24774, 16'd16960, 16'd1126, 16'd1737, 16'd23433, 16'd46566, 16'd61837});
	test_expansion(128'h63e950c1b53ba0d2ebd7234f27cccdc5, {16'd21390, 16'd60649, 16'd50411, 16'd53317, 16'd15095, 16'd22573, 16'd47502, 16'd3401, 16'd61736, 16'd2949, 16'd11434, 16'd2381, 16'd23360, 16'd38258, 16'd13386, 16'd15724, 16'd64442, 16'd23214, 16'd35540, 16'd48879, 16'd32098, 16'd37830, 16'd49147, 16'd63905, 16'd23105, 16'd2244});
	test_expansion(128'h5a73abdebe1fa4d5ec62b61393d267ff, {16'd2296, 16'd32923, 16'd53110, 16'd37940, 16'd22183, 16'd3696, 16'd7065, 16'd19341, 16'd12880, 16'd33579, 16'd56572, 16'd4859, 16'd5637, 16'd57376, 16'd25456, 16'd8848, 16'd55196, 16'd5354, 16'd43726, 16'd45428, 16'd39140, 16'd23795, 16'd17703, 16'd45668, 16'd43429, 16'd18150});
	test_expansion(128'h1f3db53d25d4c908e3d355286bbe6688, {16'd3414, 16'd13639, 16'd52197, 16'd20104, 16'd39461, 16'd51538, 16'd41476, 16'd61426, 16'd50358, 16'd49338, 16'd42560, 16'd63284, 16'd61169, 16'd21395, 16'd53044, 16'd47503, 16'd51788, 16'd44591, 16'd36737, 16'd5814, 16'd52434, 16'd28403, 16'd58639, 16'd13859, 16'd13464, 16'd48527});
	test_expansion(128'h4d6863a19d5cd85900fe0af5b3797d8a, {16'd14185, 16'd7045, 16'd16721, 16'd41096, 16'd33605, 16'd60095, 16'd43764, 16'd17766, 16'd21919, 16'd13959, 16'd1905, 16'd4593, 16'd25763, 16'd26243, 16'd42539, 16'd61618, 16'd27690, 16'd17544, 16'd29468, 16'd23176, 16'd40034, 16'd62257, 16'd14082, 16'd25523, 16'd13421, 16'd55567});
	test_expansion(128'hb95c2bbc1661f910d44b2faedf39cd8f, {16'd58162, 16'd42894, 16'd15409, 16'd17299, 16'd58569, 16'd60891, 16'd10907, 16'd64725, 16'd47983, 16'd11886, 16'd25072, 16'd2193, 16'd57481, 16'd12801, 16'd8239, 16'd34175, 16'd8928, 16'd15039, 16'd38781, 16'd7268, 16'd34977, 16'd59656, 16'd9540, 16'd21987, 16'd40084, 16'd41477});
	test_expansion(128'h4aac8e89bcf7017c622a002391a2e75c, {16'd35032, 16'd45592, 16'd43796, 16'd770, 16'd4461, 16'd20942, 16'd51518, 16'd55616, 16'd29851, 16'd5550, 16'd49069, 16'd24167, 16'd15129, 16'd34714, 16'd15549, 16'd46274, 16'd5764, 16'd46629, 16'd43238, 16'd14054, 16'd23846, 16'd27950, 16'd43216, 16'd34680, 16'd12651, 16'd11042});
	test_expansion(128'he5e8aa680743c3d5de271868ab007f0a, {16'd57051, 16'd2965, 16'd62873, 16'd14610, 16'd4067, 16'd49978, 16'd17733, 16'd36460, 16'd13633, 16'd41464, 16'd21831, 16'd42249, 16'd4846, 16'd47336, 16'd24085, 16'd2891, 16'd49438, 16'd20125, 16'd10265, 16'd14302, 16'd2814, 16'd55666, 16'd62757, 16'd32822, 16'd32283, 16'd49655});
	test_expansion(128'hd88d8ac08b7bdfae68855681045b5b6c, {16'd28577, 16'd2921, 16'd34391, 16'd50047, 16'd56915, 16'd16227, 16'd45295, 16'd35383, 16'd20256, 16'd2805, 16'd20645, 16'd14497, 16'd39285, 16'd34644, 16'd8516, 16'd64914, 16'd53729, 16'd30130, 16'd34726, 16'd38309, 16'd30583, 16'd14624, 16'd2404, 16'd57217, 16'd47851, 16'd57194});
	test_expansion(128'h374393e8fb2a6dc6ddb0a8cd3c90326a, {16'd48476, 16'd28813, 16'd49201, 16'd20792, 16'd28644, 16'd8446, 16'd11552, 16'd48449, 16'd15806, 16'd24560, 16'd62184, 16'd13539, 16'd53241, 16'd52435, 16'd28279, 16'd2597, 16'd31360, 16'd45817, 16'd50792, 16'd30625, 16'd6804, 16'd64185, 16'd35849, 16'd65392, 16'd25519, 16'd3152});
	test_expansion(128'h660d952e22c8c703a1ba74547a6427e1, {16'd41105, 16'd3011, 16'd41745, 16'd4843, 16'd22613, 16'd62758, 16'd21118, 16'd56692, 16'd22071, 16'd55965, 16'd42070, 16'd34094, 16'd33605, 16'd49946, 16'd29215, 16'd36521, 16'd63332, 16'd3195, 16'd426, 16'd41450, 16'd15012, 16'd9500, 16'd37560, 16'd41164, 16'd18157, 16'd59178});
	test_expansion(128'hbe36cbbeb65d8446576dec5acb71b8f4, {16'd28357, 16'd26045, 16'd44749, 16'd34032, 16'd32403, 16'd48799, 16'd554, 16'd20446, 16'd47768, 16'd26757, 16'd41681, 16'd41004, 16'd34669, 16'd39589, 16'd55699, 16'd47436, 16'd2444, 16'd10401, 16'd60358, 16'd20480, 16'd11598, 16'd10385, 16'd26519, 16'd19554, 16'd12738, 16'd56478});
	test_expansion(128'h915abdd36b15932794def49ba1ef6215, {16'd54343, 16'd30582, 16'd21713, 16'd64803, 16'd39815, 16'd40980, 16'd8328, 16'd19983, 16'd12659, 16'd9085, 16'd10508, 16'd31247, 16'd24791, 16'd32200, 16'd29906, 16'd63234, 16'd61768, 16'd43933, 16'd14409, 16'd29276, 16'd39822, 16'd11549, 16'd29110, 16'd17392, 16'd9134, 16'd4073});
	test_expansion(128'h580234e680afb2a5462b5a133a2e5835, {16'd32608, 16'd18003, 16'd43597, 16'd10347, 16'd399, 16'd48, 16'd2552, 16'd47355, 16'd35582, 16'd51447, 16'd21686, 16'd35139, 16'd21434, 16'd45665, 16'd30484, 16'd58144, 16'd23754, 16'd9609, 16'd56490, 16'd63435, 16'd45723, 16'd40287, 16'd49847, 16'd13116, 16'd6058, 16'd54253});
	test_expansion(128'hee84a5806b61e3be7ee725747696d8a6, {16'd10139, 16'd19824, 16'd49603, 16'd54175, 16'd43201, 16'd29624, 16'd53994, 16'd36081, 16'd60602, 16'd55798, 16'd24947, 16'd10469, 16'd31514, 16'd35331, 16'd59305, 16'd43443, 16'd40343, 16'd62329, 16'd7823, 16'd31070, 16'd25469, 16'd51424, 16'd17348, 16'd26600, 16'd52211, 16'd14508});
	test_expansion(128'h292ac2c202f89503ce0b0adf25c4eb77, {16'd61714, 16'd8728, 16'd13750, 16'd60647, 16'd61501, 16'd21683, 16'd16730, 16'd26245, 16'd7105, 16'd19004, 16'd54153, 16'd31561, 16'd62621, 16'd7670, 16'd89, 16'd38981, 16'd28963, 16'd38199, 16'd9400, 16'd56661, 16'd52419, 16'd21080, 16'd43303, 16'd19760, 16'd52875, 16'd29959});
	test_expansion(128'h7ce37e4f5ea0a488e799f179339b4f13, {16'd51820, 16'd9424, 16'd270, 16'd63629, 16'd28816, 16'd23392, 16'd19712, 16'd22313, 16'd1480, 16'd43691, 16'd61139, 16'd60019, 16'd37613, 16'd9259, 16'd5381, 16'd40549, 16'd50534, 16'd4345, 16'd33393, 16'd2132, 16'd39328, 16'd44076, 16'd12421, 16'd24168, 16'd49456, 16'd56360});
	test_expansion(128'h848ea7c500edd1b38f29e16b08f9e458, {16'd19523, 16'd61384, 16'd50689, 16'd58168, 16'd63873, 16'd44450, 16'd54349, 16'd30129, 16'd4765, 16'd64800, 16'd30913, 16'd18674, 16'd56777, 16'd4225, 16'd22840, 16'd41655, 16'd15282, 16'd29677, 16'd6433, 16'd8849, 16'd43182, 16'd38803, 16'd58500, 16'd52124, 16'd62097, 16'd3481});
	test_expansion(128'hd66f53e0b8b0ae95052dace4b4f82ea0, {16'd60140, 16'd41791, 16'd13471, 16'd20126, 16'd58255, 16'd62734, 16'd41232, 16'd49865, 16'd59053, 16'd10578, 16'd43029, 16'd38089, 16'd31057, 16'd17205, 16'd64623, 16'd2477, 16'd8216, 16'd60142, 16'd51572, 16'd26131, 16'd45307, 16'd4136, 16'd10391, 16'd33769, 16'd43302, 16'd44043});
	test_expansion(128'h0272c4d882ac8df92d5934f42f880ac0, {16'd4106, 16'd48203, 16'd15917, 16'd57861, 16'd41167, 16'd25009, 16'd15291, 16'd12006, 16'd28109, 16'd47646, 16'd31263, 16'd59645, 16'd7109, 16'd2583, 16'd9663, 16'd31472, 16'd15840, 16'd33593, 16'd40970, 16'd27840, 16'd8093, 16'd32465, 16'd6754, 16'd23730, 16'd53038, 16'd702});
	test_expansion(128'hfd53b52941233776fd79611bfc9a95e4, {16'd56654, 16'd14405, 16'd450, 16'd63500, 16'd35860, 16'd8405, 16'd52367, 16'd52263, 16'd63104, 16'd19035, 16'd30572, 16'd48352, 16'd5922, 16'd34854, 16'd50058, 16'd33949, 16'd17261, 16'd20616, 16'd20323, 16'd30484, 16'd26547, 16'd35505, 16'd35034, 16'd30040, 16'd36202, 16'd59612});
	test_expansion(128'h33057f84c1ff659ceca931c46bbe50f7, {16'd5485, 16'd24950, 16'd33279, 16'd61122, 16'd44466, 16'd3637, 16'd57699, 16'd39610, 16'd27739, 16'd44711, 16'd53052, 16'd34906, 16'd58200, 16'd56055, 16'd10695, 16'd17337, 16'd310, 16'd16209, 16'd55496, 16'd30087, 16'd24973, 16'd20343, 16'd12229, 16'd40848, 16'd3525, 16'd47118});
	test_expansion(128'h77e8599ca110495edfb511fdd4cea3b9, {16'd23747, 16'd63812, 16'd26780, 16'd56198, 16'd54817, 16'd12161, 16'd52520, 16'd18456, 16'd2514, 16'd29187, 16'd19039, 16'd12657, 16'd27344, 16'd60567, 16'd62877, 16'd62418, 16'd8096, 16'd51768, 16'd31818, 16'd26546, 16'd3216, 16'd15930, 16'd53229, 16'd30382, 16'd57589, 16'd55425});
	test_expansion(128'h5de64d32761be3984cd7918c9fdd9fc0, {16'd9600, 16'd50896, 16'd3186, 16'd24662, 16'd2867, 16'd49119, 16'd16887, 16'd49078, 16'd35416, 16'd40890, 16'd63655, 16'd12178, 16'd6984, 16'd4559, 16'd63305, 16'd16538, 16'd6725, 16'd44841, 16'd26197, 16'd49041, 16'd50921, 16'd10760, 16'd17783, 16'd31849, 16'd44976, 16'd24166});
	test_expansion(128'h552626b24e026de48561413df98d3714, {16'd52662, 16'd41993, 16'd22686, 16'd16415, 16'd54087, 16'd7849, 16'd56012, 16'd61705, 16'd45871, 16'd38464, 16'd16864, 16'd45891, 16'd25848, 16'd56424, 16'd32851, 16'd29154, 16'd36863, 16'd49084, 16'd59023, 16'd1971, 16'd58400, 16'd12916, 16'd3680, 16'd35474, 16'd14035, 16'd33465});
	test_expansion(128'hbe43b0b70b23a817ecd8289c9f0e44ee, {16'd33197, 16'd22243, 16'd43086, 16'd14163, 16'd36994, 16'd4860, 16'd65290, 16'd18288, 16'd53036, 16'd2650, 16'd3738, 16'd16178, 16'd24402, 16'd19703, 16'd3682, 16'd15400, 16'd56552, 16'd41927, 16'd57580, 16'd22234, 16'd13958, 16'd7381, 16'd64101, 16'd62756, 16'd60551, 16'd42483});
	test_expansion(128'he990273132199a28dbc6b28a0f90ada9, {16'd17856, 16'd57696, 16'd22974, 16'd28381, 16'd37161, 16'd33530, 16'd3129, 16'd60892, 16'd16682, 16'd49273, 16'd27247, 16'd41158, 16'd25306, 16'd45578, 16'd65192, 16'd25801, 16'd2342, 16'd26295, 16'd21002, 16'd63127, 16'd4294, 16'd9400, 16'd33259, 16'd45166, 16'd43725, 16'd62054});
	test_expansion(128'h00ec6852e694f89685c7f903b8132a69, {16'd28227, 16'd39280, 16'd31925, 16'd9973, 16'd26185, 16'd16773, 16'd11553, 16'd43896, 16'd7129, 16'd15810, 16'd61530, 16'd56590, 16'd3721, 16'd29357, 16'd14463, 16'd41351, 16'd11292, 16'd25577, 16'd41635, 16'd29622, 16'd10231, 16'd46093, 16'd39759, 16'd29059, 16'd14067, 16'd56715});
	test_expansion(128'h215d73d226d9341f558f764dd0a07afd, {16'd44299, 16'd58376, 16'd47330, 16'd55124, 16'd41023, 16'd37105, 16'd15599, 16'd11996, 16'd26224, 16'd668, 16'd61853, 16'd43224, 16'd44317, 16'd36400, 16'd59659, 16'd21374, 16'd40315, 16'd1913, 16'd49957, 16'd47112, 16'd21634, 16'd7877, 16'd39259, 16'd53249, 16'd22769, 16'd15436});
	test_expansion(128'ha62fb57745100a5765248915ddabcaad, {16'd49487, 16'd8833, 16'd24463, 16'd53072, 16'd52700, 16'd34808, 16'd9117, 16'd47437, 16'd21123, 16'd40017, 16'd39385, 16'd22716, 16'd35641, 16'd19166, 16'd41835, 16'd15194, 16'd25580, 16'd42552, 16'd50970, 16'd24316, 16'd61445, 16'd24384, 16'd52101, 16'd62656, 16'd57643, 16'd51475});
	test_expansion(128'h5ba34c094b0793e4249be5767977e11f, {16'd39691, 16'd23343, 16'd13879, 16'd44661, 16'd445, 16'd57319, 16'd49905, 16'd1469, 16'd1967, 16'd62290, 16'd23445, 16'd63351, 16'd58841, 16'd10779, 16'd55279, 16'd27368, 16'd19227, 16'd46553, 16'd15136, 16'd20928, 16'd47333, 16'd17489, 16'd59729, 16'd1454, 16'd40987, 16'd47986});
	test_expansion(128'hab8769c88b5b02f1e1de96ba6e965dee, {16'd17186, 16'd28641, 16'd3794, 16'd49171, 16'd54127, 16'd54041, 16'd19378, 16'd57598, 16'd62633, 16'd59091, 16'd24864, 16'd56562, 16'd18715, 16'd42454, 16'd39351, 16'd35521, 16'd20924, 16'd922, 16'd201, 16'd7632, 16'd18804, 16'd27404, 16'd43828, 16'd51116, 16'd52066, 16'd47858});
	test_expansion(128'h683a16d737e9bafe191ca48e2466afe0, {16'd61981, 16'd31795, 16'd50959, 16'd28423, 16'd60723, 16'd26865, 16'd36323, 16'd55253, 16'd19885, 16'd61426, 16'd21818, 16'd18733, 16'd34438, 16'd20508, 16'd32910, 16'd23402, 16'd14772, 16'd39721, 16'd26806, 16'd10916, 16'd43534, 16'd14441, 16'd46145, 16'd1030, 16'd59796, 16'd53814});
	test_expansion(128'h9fbe4aa9bfa14f17af0ffdc9713d3491, {16'd44636, 16'd59403, 16'd42822, 16'd32824, 16'd49738, 16'd10788, 16'd11026, 16'd65357, 16'd63404, 16'd4674, 16'd45931, 16'd25255, 16'd29186, 16'd65404, 16'd46681, 16'd18762, 16'd13714, 16'd7739, 16'd5300, 16'd37597, 16'd61391, 16'd29149, 16'd12326, 16'd22134, 16'd49921, 16'd21971});
	test_expansion(128'hf7657a7e12edfc8dd3e98bdecc971365, {16'd38078, 16'd13690, 16'd51472, 16'd28374, 16'd21088, 16'd26115, 16'd60378, 16'd28270, 16'd60191, 16'd37067, 16'd28030, 16'd10634, 16'd27316, 16'd13136, 16'd64463, 16'd49752, 16'd34970, 16'd54192, 16'd49040, 16'd49001, 16'd9309, 16'd119, 16'd51308, 16'd20620, 16'd61690, 16'd59874});
	test_expansion(128'h41dc5eb5f84aeb2dbb3578d68a18540e, {16'd2057, 16'd12570, 16'd20437, 16'd49248, 16'd32803, 16'd36575, 16'd3986, 16'd39570, 16'd31501, 16'd58902, 16'd41042, 16'd61802, 16'd20573, 16'd6964, 16'd46610, 16'd29417, 16'd34039, 16'd7377, 16'd39224, 16'd2196, 16'd55491, 16'd20777, 16'd65059, 16'd21593, 16'd2769, 16'd46334});
	test_expansion(128'h07e52d674119cc3e994ea6e2cea30a54, {16'd21420, 16'd27403, 16'd53414, 16'd19335, 16'd10313, 16'd55611, 16'd33034, 16'd52512, 16'd65012, 16'd29437, 16'd48610, 16'd61582, 16'd18888, 16'd582, 16'd28288, 16'd13114, 16'd61296, 16'd41511, 16'd39163, 16'd16438, 16'd60646, 16'd12544, 16'd42782, 16'd56438, 16'd43298, 16'd48916});
	test_expansion(128'ha9d48de5ddaec35b21408328295c4acd, {16'd8506, 16'd39599, 16'd48554, 16'd55878, 16'd23443, 16'd45603, 16'd57689, 16'd43234, 16'd52330, 16'd41844, 16'd4836, 16'd31977, 16'd55286, 16'd30064, 16'd29353, 16'd12062, 16'd31283, 16'd4234, 16'd51825, 16'd36279, 16'd14020, 16'd16111, 16'd35685, 16'd53109, 16'd48513, 16'd30845});
	test_expansion(128'h79de8e59b5b64955b90f2fb60ea70ee8, {16'd16607, 16'd136, 16'd26021, 16'd62277, 16'd4337, 16'd51567, 16'd33500, 16'd42879, 16'd49963, 16'd7409, 16'd55187, 16'd16386, 16'd40059, 16'd49498, 16'd49343, 16'd28288, 16'd61014, 16'd6817, 16'd8140, 16'd35499, 16'd18961, 16'd6402, 16'd59599, 16'd41928, 16'd19075, 16'd60106});
	test_expansion(128'h903259aea5c9cd132cc561acd8e50680, {16'd64704, 16'd60416, 16'd39604, 16'd622, 16'd30596, 16'd7347, 16'd17663, 16'd21035, 16'd12345, 16'd21561, 16'd34322, 16'd44135, 16'd7070, 16'd32299, 16'd12123, 16'd61007, 16'd26994, 16'd30901, 16'd7475, 16'd4689, 16'd60910, 16'd27713, 16'd27038, 16'd39610, 16'd20243, 16'd17063});
	test_expansion(128'h3211c9202edfaaa71504daa3bd1ee318, {16'd61587, 16'd62612, 16'd31495, 16'd48152, 16'd47600, 16'd30915, 16'd48165, 16'd12094, 16'd45426, 16'd10131, 16'd27064, 16'd53432, 16'd55761, 16'd38077, 16'd12675, 16'd56978, 16'd2253, 16'd49521, 16'd29930, 16'd39563, 16'd31520, 16'd30936, 16'd46405, 16'd14919, 16'd17006, 16'd40192});
	test_expansion(128'h4a7ed52c9ba0a839b7f5ac1cb2735f81, {16'd56715, 16'd31250, 16'd35854, 16'd31680, 16'd22035, 16'd10784, 16'd17820, 16'd28352, 16'd47710, 16'd64465, 16'd28736, 16'd33407, 16'd4230, 16'd54151, 16'd12306, 16'd498, 16'd13834, 16'd60529, 16'd59746, 16'd37544, 16'd29877, 16'd19447, 16'd14087, 16'd36665, 16'd29676, 16'd117});
	test_expansion(128'he9bacce059a2b0397ece3bcffc3f7695, {16'd33470, 16'd57219, 16'd50957, 16'd60316, 16'd45376, 16'd1960, 16'd10690, 16'd1627, 16'd50000, 16'd57366, 16'd23101, 16'd13673, 16'd26151, 16'd36185, 16'd11570, 16'd59070, 16'd42989, 16'd21380, 16'd9193, 16'd41665, 16'd52864, 16'd22641, 16'd40867, 16'd26442, 16'd50148, 16'd19679});
	test_expansion(128'h2e0e017dd98d5f9aba26cf90c9e26d3a, {16'd14121, 16'd118, 16'd23548, 16'd17815, 16'd42315, 16'd27852, 16'd55488, 16'd18803, 16'd29094, 16'd32470, 16'd16589, 16'd64625, 16'd4889, 16'd22819, 16'd9268, 16'd24342, 16'd48744, 16'd39996, 16'd33624, 16'd21855, 16'd30893, 16'd36584, 16'd50645, 16'd25317, 16'd1118, 16'd26587});
	test_expansion(128'h93893de22339654bbc3e0a5f1079d801, {16'd29091, 16'd51791, 16'd43171, 16'd10065, 16'd4645, 16'd13374, 16'd19265, 16'd59324, 16'd64525, 16'd28488, 16'd65502, 16'd15537, 16'd59756, 16'd59859, 16'd17375, 16'd53171, 16'd10385, 16'd32838, 16'd46262, 16'd4293, 16'd25743, 16'd47257, 16'd21516, 16'd35374, 16'd12481, 16'd28155});
	test_expansion(128'hd4d807f9cc0812ab7874875539c10ffb, {16'd57424, 16'd16515, 16'd6701, 16'd55139, 16'd32959, 16'd31510, 16'd23302, 16'd55047, 16'd841, 16'd20291, 16'd58267, 16'd62370, 16'd64812, 16'd55299, 16'd8379, 16'd64079, 16'd39161, 16'd34122, 16'd25618, 16'd13645, 16'd22263, 16'd48469, 16'd12225, 16'd1056, 16'd35677, 16'd7674});
	test_expansion(128'h9b918e37df882c7395b9c9302ab301df, {16'd32488, 16'd48141, 16'd21456, 16'd25917, 16'd14996, 16'd2728, 16'd50152, 16'd15988, 16'd31742, 16'd33372, 16'd20195, 16'd37420, 16'd7342, 16'd50019, 16'd21592, 16'd41029, 16'd39613, 16'd60938, 16'd12265, 16'd52065, 16'd27055, 16'd60404, 16'd25760, 16'd30333, 16'd45375, 16'd38011});
	test_expansion(128'h90436ae1e7460d9faf01d74abb54dfc2, {16'd33616, 16'd25151, 16'd4860, 16'd41581, 16'd26555, 16'd43500, 16'd8201, 16'd25113, 16'd54145, 16'd53846, 16'd7067, 16'd14448, 16'd14890, 16'd34815, 16'd4616, 16'd44953, 16'd12174, 16'd6315, 16'd10994, 16'd43084, 16'd18582, 16'd3587, 16'd26296, 16'd22862, 16'd37147, 16'd45886});
	test_expansion(128'hb69658a4b4ec73155d7cfb04888b20fc, {16'd43043, 16'd4657, 16'd6277, 16'd27712, 16'd47135, 16'd2999, 16'd8970, 16'd48456, 16'd44814, 16'd33531, 16'd38400, 16'd37256, 16'd5008, 16'd49729, 16'd54721, 16'd49050, 16'd6169, 16'd26168, 16'd50472, 16'd32395, 16'd56814, 16'd8866, 16'd28866, 16'd2120, 16'd45720, 16'd42540});
	test_expansion(128'hef47fbd61c6b2f1b97f67722b4b2abd2, {16'd54034, 16'd53041, 16'd42544, 16'd3021, 16'd13780, 16'd49591, 16'd33186, 16'd31524, 16'd26302, 16'd38936, 16'd21640, 16'd13242, 16'd49766, 16'd43638, 16'd60904, 16'd51512, 16'd22815, 16'd2714, 16'd13064, 16'd32339, 16'd7375, 16'd22875, 16'd50344, 16'd42419, 16'd17278, 16'd16923});
	test_expansion(128'h59f8d5f712ceebeb03ccfaa685ba7ba8, {16'd27825, 16'd5683, 16'd28988, 16'd54846, 16'd19020, 16'd60774, 16'd10632, 16'd49974, 16'd39468, 16'd12674, 16'd13003, 16'd41800, 16'd33563, 16'd48190, 16'd29013, 16'd18347, 16'd38054, 16'd40309, 16'd28557, 16'd27961, 16'd51387, 16'd27696, 16'd5610, 16'd47186, 16'd63573, 16'd28754});
	test_expansion(128'hf8b9a53a3fe69bd82d5cdf568ab84661, {16'd64524, 16'd54039, 16'd12099, 16'd19673, 16'd58989, 16'd20434, 16'd22892, 16'd343, 16'd42697, 16'd23554, 16'd25622, 16'd52175, 16'd59442, 16'd65505, 16'd16902, 16'd49323, 16'd19049, 16'd33031, 16'd61307, 16'd49527, 16'd48446, 16'd45935, 16'd61830, 16'd58591, 16'd8040, 16'd40602});
	test_expansion(128'h4d5166b2f314a3385af771a0fce2589f, {16'd27905, 16'd36228, 16'd27914, 16'd18821, 16'd35744, 16'd43975, 16'd40945, 16'd1213, 16'd7563, 16'd29026, 16'd48606, 16'd11773, 16'd64500, 16'd27187, 16'd47839, 16'd36876, 16'd46687, 16'd58966, 16'd30409, 16'd33126, 16'd51980, 16'd50099, 16'd23608, 16'd2658, 16'd26984, 16'd36676});
	test_expansion(128'h3e9a34ad198ac6e85ac913f62520b15a, {16'd35346, 16'd3221, 16'd44700, 16'd20604, 16'd5004, 16'd1851, 16'd55733, 16'd15171, 16'd18662, 16'd56465, 16'd54201, 16'd55991, 16'd23536, 16'd6395, 16'd52062, 16'd5708, 16'd21228, 16'd40332, 16'd17821, 16'd33165, 16'd28139, 16'd13523, 16'd42002, 16'd60885, 16'd33364, 16'd44582});
	test_expansion(128'he4588274223a0abe76cee5dbc10b4f34, {16'd9742, 16'd34089, 16'd45913, 16'd37055, 16'd8612, 16'd24076, 16'd27069, 16'd64171, 16'd46770, 16'd63943, 16'd64638, 16'd14769, 16'd46398, 16'd49199, 16'd24398, 16'd35157, 16'd15656, 16'd58903, 16'd9779, 16'd45032, 16'd48830, 16'd5917, 16'd44379, 16'd59150, 16'd497, 16'd33367});
	test_expansion(128'h7baecf992adb0976ccd2950cdf676d93, {16'd21961, 16'd34031, 16'd23383, 16'd36985, 16'd56366, 16'd48399, 16'd39392, 16'd60999, 16'd29186, 16'd2566, 16'd38372, 16'd34733, 16'd12803, 16'd43561, 16'd27125, 16'd46095, 16'd64211, 16'd3929, 16'd47103, 16'd63253, 16'd65385, 16'd3851, 16'd27616, 16'd34187, 16'd12654, 16'd8884});
	test_expansion(128'hbbc47d1e0c313b159f6cb63fbb155b2d, {16'd22664, 16'd61741, 16'd22996, 16'd12107, 16'd32633, 16'd8687, 16'd61624, 16'd15578, 16'd51215, 16'd33523, 16'd45341, 16'd53337, 16'd21083, 16'd46615, 16'd45068, 16'd10414, 16'd55371, 16'd2612, 16'd38799, 16'd18288, 16'd42846, 16'd332, 16'd51970, 16'd34249, 16'd6005, 16'd29464});
	test_expansion(128'h19d2cb6e764946c9520067a324252849, {16'd27105, 16'd2038, 16'd53751, 16'd4222, 16'd14436, 16'd16170, 16'd55587, 16'd64197, 16'd9312, 16'd43136, 16'd11713, 16'd49309, 16'd23494, 16'd63607, 16'd57684, 16'd2726, 16'd41681, 16'd56143, 16'd40257, 16'd7515, 16'd29369, 16'd10255, 16'd25093, 16'd55580, 16'd60689, 16'd56357});
	test_expansion(128'hbce028cbd82c9fb264a49ac1e9d3e04a, {16'd18804, 16'd49021, 16'd11205, 16'd29743, 16'd13334, 16'd50924, 16'd4610, 16'd19853, 16'd52052, 16'd17702, 16'd10593, 16'd2642, 16'd35875, 16'd32221, 16'd58681, 16'd42457, 16'd15143, 16'd55841, 16'd24644, 16'd40597, 16'd5070, 16'd51597, 16'd44053, 16'd46544, 16'd54110, 16'd3415});
	test_expansion(128'hedbaf092b45b2c1f886917d772352c19, {16'd26937, 16'd2496, 16'd14452, 16'd9469, 16'd15924, 16'd59666, 16'd20864, 16'd30177, 16'd38609, 16'd53560, 16'd28830, 16'd61165, 16'd11968, 16'd22855, 16'd5775, 16'd11171, 16'd2796, 16'd46184, 16'd15914, 16'd61566, 16'd11791, 16'd63937, 16'd8364, 16'd13683, 16'd24961, 16'd25156});
	test_expansion(128'h9b474da12dbde78aa933cc8e8671106d, {16'd48208, 16'd20765, 16'd58350, 16'd58586, 16'd63355, 16'd15840, 16'd58572, 16'd38697, 16'd52626, 16'd22444, 16'd4151, 16'd35856, 16'd42016, 16'd31445, 16'd48190, 16'd36824, 16'd11172, 16'd56786, 16'd11400, 16'd37198, 16'd24262, 16'd51193, 16'd23330, 16'd64129, 16'd45915, 16'd20473});
	test_expansion(128'h62c194ccaea62566748d6ed0c4abecfd, {16'd53168, 16'd2649, 16'd64036, 16'd51138, 16'd64966, 16'd63777, 16'd45546, 16'd78, 16'd55857, 16'd8674, 16'd15434, 16'd5695, 16'd55323, 16'd32663, 16'd5022, 16'd39559, 16'd52932, 16'd50695, 16'd9562, 16'd60794, 16'd39520, 16'd12774, 16'd57745, 16'd25241, 16'd4432, 16'd39096});
	test_expansion(128'hd38f2a1c77b92fa09e669329dc6b3b33, {16'd26726, 16'd36372, 16'd25522, 16'd3469, 16'd33089, 16'd59446, 16'd41077, 16'd48515, 16'd2575, 16'd10794, 16'd7449, 16'd50592, 16'd17505, 16'd44766, 16'd43542, 16'd10666, 16'd17497, 16'd32403, 16'd32403, 16'd62300, 16'd32727, 16'd37006, 16'd32183, 16'd48504, 16'd44085, 16'd55882});
	test_expansion(128'hd84ffdb6dfbd573206e64c9f4ccd0cb4, {16'd29414, 16'd5599, 16'd64325, 16'd372, 16'd47680, 16'd48323, 16'd47417, 16'd51756, 16'd10379, 16'd57244, 16'd35140, 16'd19218, 16'd26028, 16'd18055, 16'd54105, 16'd42482, 16'd21420, 16'd3273, 16'd3491, 16'd22484, 16'd26109, 16'd57543, 16'd1905, 16'd25955, 16'd27719, 16'd36140});
	test_expansion(128'h9e07be9b737b82aad9fc15f9eee1321b, {16'd20169, 16'd61820, 16'd4375, 16'd5397, 16'd37932, 16'd44072, 16'd1712, 16'd19945, 16'd15962, 16'd4686, 16'd18810, 16'd15266, 16'd31409, 16'd53186, 16'd64404, 16'd44307, 16'd37773, 16'd17251, 16'd44426, 16'd51388, 16'd39959, 16'd64145, 16'd3297, 16'd9478, 16'd64799, 16'd4852});
	test_expansion(128'hee83e371d3ee0cdcc36fbcfddabfc3fb, {16'd62150, 16'd44344, 16'd28113, 16'd11315, 16'd56731, 16'd39117, 16'd52805, 16'd21274, 16'd4319, 16'd33094, 16'd3540, 16'd43167, 16'd38724, 16'd54002, 16'd50468, 16'd40836, 16'd55276, 16'd61396, 16'd28434, 16'd65449, 16'd61698, 16'd39971, 16'd58188, 16'd783, 16'd37267, 16'd27503});
	test_expansion(128'hba166bf1597416978070636348891b6c, {16'd2078, 16'd60625, 16'd54368, 16'd41907, 16'd11440, 16'd1102, 16'd51727, 16'd2216, 16'd23715, 16'd56649, 16'd42112, 16'd11119, 16'd48127, 16'd88, 16'd36320, 16'd30127, 16'd34087, 16'd48516, 16'd18564, 16'd10480, 16'd58407, 16'd53038, 16'd22534, 16'd16449, 16'd51021, 16'd38248});
	test_expansion(128'h2112250fc25ca460e836b0b699a4fd6f, {16'd64377, 16'd33816, 16'd54278, 16'd56398, 16'd2166, 16'd35457, 16'd35876, 16'd5531, 16'd25333, 16'd38948, 16'd59970, 16'd22391, 16'd51932, 16'd40185, 16'd10220, 16'd51376, 16'd10605, 16'd58826, 16'd44306, 16'd8528, 16'd17031, 16'd8878, 16'd44440, 16'd16280, 16'd47936, 16'd4963});
	test_expansion(128'h3a4661ff57ff082bac89c2cc32b3a394, {16'd19270, 16'd41398, 16'd53158, 16'd56384, 16'd25166, 16'd60552, 16'd17336, 16'd13122, 16'd33558, 16'd55290, 16'd1568, 16'd22287, 16'd46390, 16'd20325, 16'd19122, 16'd32131, 16'd26963, 16'd29557, 16'd37295, 16'd51452, 16'd57436, 16'd36033, 16'd13605, 16'd27051, 16'd40029, 16'd46450});
	test_expansion(128'h6d490853a1535acd962ed9089781f90c, {16'd30884, 16'd4294, 16'd57233, 16'd21538, 16'd20032, 16'd55160, 16'd57053, 16'd54147, 16'd21792, 16'd39108, 16'd24634, 16'd53506, 16'd6082, 16'd61327, 16'd3298, 16'd45564, 16'd33921, 16'd64789, 16'd31287, 16'd19924, 16'd30747, 16'd56949, 16'd20092, 16'd43608, 16'd42161, 16'd12682});
	test_expansion(128'hea456069b5c190969dc008f5ae32422f, {16'd738, 16'd21505, 16'd63526, 16'd17058, 16'd22820, 16'd57960, 16'd22237, 16'd61195, 16'd35955, 16'd54692, 16'd58364, 16'd6517, 16'd7386, 16'd57988, 16'd43735, 16'd22911, 16'd18507, 16'd48702, 16'd50319, 16'd19352, 16'd50162, 16'd4294, 16'd25440, 16'd41230, 16'd59650, 16'd2657});
	test_expansion(128'h8762b6c66eb92a1e9d4a0ad1e85a15bb, {16'd28484, 16'd36022, 16'd10796, 16'd43713, 16'd9922, 16'd50764, 16'd44806, 16'd36479, 16'd8631, 16'd27623, 16'd51489, 16'd40598, 16'd10281, 16'd57710, 16'd44751, 16'd32978, 16'd24522, 16'd44558, 16'd20151, 16'd21058, 16'd19842, 16'd29274, 16'd37946, 16'd20623, 16'd18006, 16'd23551});
	test_expansion(128'h5832f4fb54e3828f1838094175263d35, {16'd2279, 16'd5473, 16'd3015, 16'd10336, 16'd565, 16'd60337, 16'd50762, 16'd55898, 16'd49833, 16'd22917, 16'd31058, 16'd64459, 16'd49927, 16'd65159, 16'd59926, 16'd11007, 16'd21010, 16'd6452, 16'd44021, 16'd61814, 16'd26738, 16'd37325, 16'd43739, 16'd44811, 16'd7815, 16'd15511});
	test_expansion(128'h716834d6804f0d0fa4aefe7b78c08b7f, {16'd35867, 16'd28928, 16'd60706, 16'd50541, 16'd6974, 16'd35250, 16'd35809, 16'd4471, 16'd24708, 16'd9655, 16'd32478, 16'd57500, 16'd9152, 16'd37622, 16'd54919, 16'd2913, 16'd18418, 16'd34456, 16'd13225, 16'd5926, 16'd17132, 16'd39768, 16'd62411, 16'd9665, 16'd44883, 16'd8825});
	test_expansion(128'h5e5189072e32351fad86d177706533ff, {16'd31361, 16'd63929, 16'd31651, 16'd39421, 16'd18802, 16'd17597, 16'd42238, 16'd50093, 16'd22570, 16'd18109, 16'd17857, 16'd26671, 16'd13805, 16'd20478, 16'd21316, 16'd50126, 16'd9298, 16'd39689, 16'd54700, 16'd15704, 16'd61541, 16'd59171, 16'd34367, 16'd1575, 16'd289, 16'd27391});
	test_expansion(128'h9a7f84201b15db658331c442820cb580, {16'd65221, 16'd60465, 16'd4015, 16'd40127, 16'd20515, 16'd37682, 16'd38776, 16'd21955, 16'd56261, 16'd17348, 16'd56568, 16'd7865, 16'd65438, 16'd24515, 16'd35580, 16'd64163, 16'd50126, 16'd44405, 16'd43637, 16'd2978, 16'd1535, 16'd23264, 16'd12747, 16'd52332, 16'd1259, 16'd39756});
	test_expansion(128'hf15e853277d495c738d0ec59d63f3223, {16'd11065, 16'd62097, 16'd61541, 16'd9966, 16'd25555, 16'd144, 16'd22914, 16'd62146, 16'd58188, 16'd1625, 16'd5267, 16'd54750, 16'd40304, 16'd65204, 16'd328, 16'd11810, 16'd38675, 16'd10397, 16'd33234, 16'd8578, 16'd37312, 16'd60441, 16'd7841, 16'd17532, 16'd30183, 16'd17359});
	test_expansion(128'hb65676257badb44d52f1538905c1db77, {16'd19536, 16'd46209, 16'd53462, 16'd12891, 16'd26733, 16'd17559, 16'd23306, 16'd9341, 16'd6878, 16'd54011, 16'd11189, 16'd60704, 16'd18534, 16'd19959, 16'd15474, 16'd10349, 16'd12675, 16'd22883, 16'd25369, 16'd26324, 16'd18571, 16'd41878, 16'd51411, 16'd51178, 16'd46666, 16'd24583});
	test_expansion(128'h058fc01e6fac096f0728f4c5faf08f56, {16'd45434, 16'd32907, 16'd42085, 16'd11695, 16'd48029, 16'd10303, 16'd59984, 16'd27959, 16'd5971, 16'd34513, 16'd42900, 16'd43260, 16'd24666, 16'd61183, 16'd28058, 16'd59159, 16'd47077, 16'd58130, 16'd25667, 16'd52491, 16'd54247, 16'd39988, 16'd15209, 16'd48825, 16'd42995, 16'd1260});
	test_expansion(128'h89ccc5133907c87258fdbd71c30f4875, {16'd45977, 16'd5113, 16'd38484, 16'd984, 16'd33482, 16'd40251, 16'd27148, 16'd6112, 16'd6591, 16'd4475, 16'd49567, 16'd44986, 16'd29589, 16'd16463, 16'd31, 16'd61736, 16'd5543, 16'd15779, 16'd32555, 16'd20989, 16'd46250, 16'd32278, 16'd54945, 16'd17133, 16'd5488, 16'd5858});
	test_expansion(128'h5b3b1a29a35a36dfa7986f38b84f2311, {16'd14203, 16'd34209, 16'd57284, 16'd59483, 16'd37979, 16'd17718, 16'd20419, 16'd52397, 16'd62471, 16'd28750, 16'd9571, 16'd40166, 16'd14941, 16'd28131, 16'd57487, 16'd48727, 16'd13449, 16'd52513, 16'd17742, 16'd9745, 16'd21301, 16'd45980, 16'd30122, 16'd45222, 16'd51055, 16'd12895});
	test_expansion(128'hfbf784d2c14a1cc68a9343ff260c80ff, {16'd15321, 16'd30457, 16'd6507, 16'd34754, 16'd52821, 16'd22422, 16'd17742, 16'd36947, 16'd5158, 16'd61461, 16'd16506, 16'd19753, 16'd56749, 16'd50742, 16'd27373, 16'd14280, 16'd55066, 16'd15541, 16'd16675, 16'd10666, 16'd38754, 16'd51356, 16'd2385, 16'd6224, 16'd9460, 16'd62937});
	test_expansion(128'h7879ae5b6300e198e35f30b57e5c862c, {16'd31519, 16'd5869, 16'd57980, 16'd14752, 16'd6475, 16'd25698, 16'd16906, 16'd28729, 16'd32458, 16'd62876, 16'd13485, 16'd42539, 16'd50156, 16'd9328, 16'd20956, 16'd28284, 16'd15242, 16'd16730, 16'd41564, 16'd20763, 16'd20073, 16'd49429, 16'd18674, 16'd31705, 16'd45388, 16'd26214});
	test_expansion(128'h64fe0e0baf84e5af78cd83c3dd8c9e7b, {16'd64210, 16'd62959, 16'd6148, 16'd52293, 16'd47632, 16'd46585, 16'd14219, 16'd9587, 16'd34868, 16'd36517, 16'd37702, 16'd24765, 16'd20933, 16'd16203, 16'd13123, 16'd59275, 16'd64275, 16'd60896, 16'd1148, 16'd41587, 16'd46603, 16'd31076, 16'd37847, 16'd20789, 16'd30060, 16'd46777});
	test_expansion(128'ha3166f3ceb180f5506f32a18ecd2b19b, {16'd59988, 16'd15409, 16'd16500, 16'd24291, 16'd40840, 16'd60789, 16'd54853, 16'd64304, 16'd27077, 16'd40540, 16'd27715, 16'd7561, 16'd44964, 16'd3023, 16'd25823, 16'd5855, 16'd58260, 16'd53793, 16'd25070, 16'd33055, 16'd26896, 16'd42738, 16'd58786, 16'd37314, 16'd43750, 16'd3915});
	test_expansion(128'hebaedcc0ff79ae7c11b442775881d949, {16'd7978, 16'd44921, 16'd61927, 16'd11357, 16'd37000, 16'd31931, 16'd13233, 16'd29215, 16'd33649, 16'd50215, 16'd26567, 16'd44635, 16'd53046, 16'd47207, 16'd53511, 16'd49257, 16'd9941, 16'd52506, 16'd59995, 16'd44312, 16'd15104, 16'd64330, 16'd36248, 16'd41578, 16'd20385, 16'd13949});
	test_expansion(128'hf323b943ce0258466846505ed2678988, {16'd56201, 16'd29280, 16'd64705, 16'd61620, 16'd20777, 16'd32762, 16'd24691, 16'd21433, 16'd23285, 16'd24623, 16'd18756, 16'd58522, 16'd37954, 16'd64314, 16'd14520, 16'd27665, 16'd56373, 16'd51331, 16'd38848, 16'd7934, 16'd29732, 16'd56238, 16'd50283, 16'd17636, 16'd32347, 16'd31657});
	test_expansion(128'h58a3e37eb24a8f9a07963edc6506e951, {16'd47898, 16'd10304, 16'd52759, 16'd13756, 16'd44376, 16'd61298, 16'd47615, 16'd39649, 16'd56111, 16'd20008, 16'd9726, 16'd31704, 16'd258, 16'd22346, 16'd53581, 16'd12432, 16'd14552, 16'd48818, 16'd32666, 16'd13970, 16'd31324, 16'd42276, 16'd65510, 16'd61340, 16'd43227, 16'd31440});
	test_expansion(128'hc3b1c79765041b29123aa95dce95724d, {16'd47871, 16'd54995, 16'd57366, 16'd55931, 16'd35489, 16'd27733, 16'd36533, 16'd34600, 16'd35079, 16'd24656, 16'd36238, 16'd56491, 16'd22541, 16'd10116, 16'd8469, 16'd10356, 16'd40206, 16'd53048, 16'd4878, 16'd34885, 16'd57355, 16'd11507, 16'd60219, 16'd29239, 16'd16846, 16'd58578});
	test_expansion(128'h2c42c27529aa0b5e54a8c185eaeea4f4, {16'd9202, 16'd3519, 16'd24080, 16'd22903, 16'd2630, 16'd10368, 16'd18013, 16'd62840, 16'd55950, 16'd42871, 16'd8934, 16'd16520, 16'd42125, 16'd11815, 16'd10076, 16'd17732, 16'd9768, 16'd43022, 16'd33398, 16'd55052, 16'd51492, 16'd47629, 16'd2396, 16'd53865, 16'd49124, 16'd41818});
	test_expansion(128'h7a5961773a49e10d704fed002c246e86, {16'd55963, 16'd61894, 16'd12920, 16'd34093, 16'd55419, 16'd8699, 16'd41722, 16'd15555, 16'd12168, 16'd44976, 16'd54942, 16'd8875, 16'd54643, 16'd24983, 16'd41968, 16'd41389, 16'd34674, 16'd37840, 16'd58172, 16'd24877, 16'd21796, 16'd20685, 16'd26694, 16'd25837, 16'd40738, 16'd46018});
	test_expansion(128'hd8dde62b8ea63418d4bcaf0f8cdf0ef0, {16'd17964, 16'd22333, 16'd54704, 16'd53922, 16'd14404, 16'd38276, 16'd6644, 16'd5169, 16'd24368, 16'd6639, 16'd24153, 16'd8338, 16'd42969, 16'd35043, 16'd880, 16'd14287, 16'd12286, 16'd40306, 16'd12294, 16'd6370, 16'd37134, 16'd29935, 16'd47641, 16'd43660, 16'd12077, 16'd60973});
	test_expansion(128'he01eace780564f0483c26664e5d8e364, {16'd14591, 16'd59288, 16'd39448, 16'd61, 16'd3295, 16'd63353, 16'd7523, 16'd39904, 16'd38274, 16'd51077, 16'd16150, 16'd43534, 16'd44739, 16'd1774, 16'd49043, 16'd33219, 16'd25825, 16'd43523, 16'd21972, 16'd49252, 16'd47721, 16'd10868, 16'd24336, 16'd26826, 16'd18505, 16'd48748});
	test_expansion(128'h8324c2d0586042d7beb27025295883c9, {16'd48355, 16'd2931, 16'd1317, 16'd31170, 16'd29394, 16'd25660, 16'd33045, 16'd38451, 16'd45004, 16'd58021, 16'd5472, 16'd14779, 16'd46628, 16'd54039, 16'd15940, 16'd57844, 16'd2589, 16'd31845, 16'd1996, 16'd59776, 16'd31105, 16'd22000, 16'd16671, 16'd24315, 16'd17808, 16'd62915});
	test_expansion(128'hf364f8d09c434479770726e633d10bab, {16'd25638, 16'd36113, 16'd8881, 16'd59644, 16'd64996, 16'd33680, 16'd43209, 16'd21114, 16'd44128, 16'd22403, 16'd23606, 16'd61711, 16'd58460, 16'd24524, 16'd34733, 16'd28840, 16'd22861, 16'd24249, 16'd2956, 16'd25848, 16'd1132, 16'd64001, 16'd41142, 16'd31522, 16'd9182, 16'd13309});
	test_expansion(128'h54099b90de5876bab71af6a1a172b8ae, {16'd44991, 16'd43640, 16'd36732, 16'd54530, 16'd63152, 16'd28530, 16'd25792, 16'd25537, 16'd48493, 16'd22010, 16'd7201, 16'd55669, 16'd32035, 16'd48784, 16'd39223, 16'd10239, 16'd32090, 16'd49969, 16'd41531, 16'd6904, 16'd92, 16'd53995, 16'd49410, 16'd39395, 16'd62377, 16'd16967});
	test_expansion(128'hff327c6b7046d3272fa2e50bf72d34e0, {16'd14435, 16'd53449, 16'd48400, 16'd65226, 16'd29318, 16'd26692, 16'd7447, 16'd59956, 16'd27917, 16'd61083, 16'd18369, 16'd43514, 16'd31517, 16'd22782, 16'd44419, 16'd28799, 16'd14504, 16'd11240, 16'd38629, 16'd3626, 16'd47903, 16'd43141, 16'd47465, 16'd40757, 16'd3142, 16'd31990});
	test_expansion(128'h99f2aa4d0ec12b6011236fca10805de7, {16'd6762, 16'd52217, 16'd41816, 16'd52833, 16'd42516, 16'd43359, 16'd31500, 16'd4710, 16'd6446, 16'd34, 16'd3687, 16'd20895, 16'd1254, 16'd41132, 16'd18600, 16'd35368, 16'd13451, 16'd39612, 16'd49463, 16'd3351, 16'd22927, 16'd57873, 16'd56941, 16'd47394, 16'd8411, 16'd6891});
	test_expansion(128'h4d0f535b87350a3fbb16714b1ffaea2f, {16'd63832, 16'd29390, 16'd41073, 16'd31677, 16'd273, 16'd52871, 16'd1802, 16'd28967, 16'd23991, 16'd63373, 16'd26850, 16'd10979, 16'd55062, 16'd19083, 16'd1904, 16'd62563, 16'd24340, 16'd21451, 16'd26209, 16'd59572, 16'd9771, 16'd33969, 16'd45077, 16'd60849, 16'd16934, 16'd16422});
	test_expansion(128'h4b793008129c63356726873248252db8, {16'd51087, 16'd23199, 16'd61020, 16'd18178, 16'd7271, 16'd31634, 16'd61487, 16'd45723, 16'd50272, 16'd10260, 16'd61701, 16'd22140, 16'd45342, 16'd50084, 16'd58041, 16'd57145, 16'd23153, 16'd29659, 16'd46352, 16'd59079, 16'd52173, 16'd30097, 16'd9568, 16'd536, 16'd23910, 16'd28584});
	test_expansion(128'h403afede5d0ec629b365bb8c4204725e, {16'd27237, 16'd6417, 16'd23483, 16'd51151, 16'd41526, 16'd55672, 16'd44247, 16'd51506, 16'd2171, 16'd195, 16'd62571, 16'd52153, 16'd7963, 16'd10579, 16'd48260, 16'd40472, 16'd20280, 16'd7301, 16'd26012, 16'd17027, 16'd9382, 16'd64621, 16'd31740, 16'd43304, 16'd55319, 16'd16031});
	test_expansion(128'h5cf0dfa5d0099fa40b34043bb387bbf4, {16'd28004, 16'd28646, 16'd37086, 16'd33620, 16'd20200, 16'd32203, 16'd42222, 16'd38101, 16'd4461, 16'd8032, 16'd52769, 16'd60561, 16'd44332, 16'd26851, 16'd14902, 16'd63065, 16'd35775, 16'd57526, 16'd9376, 16'd30219, 16'd27090, 16'd28634, 16'd59431, 16'd27435, 16'd29949, 16'd5097});
	test_expansion(128'hf21b318038d9e34cd1fc36af047b4eb9, {16'd61768, 16'd8011, 16'd5302, 16'd27674, 16'd57611, 16'd28278, 16'd2970, 16'd56608, 16'd15110, 16'd25689, 16'd58794, 16'd10719, 16'd22919, 16'd17454, 16'd21162, 16'd59391, 16'd17583, 16'd59235, 16'd49797, 16'd45248, 16'd31696, 16'd62848, 16'd62038, 16'd60577, 16'd1984, 16'd21775});
	test_expansion(128'h78c451adaf6d9c28c10935cdbf398ace, {16'd32647, 16'd5695, 16'd36633, 16'd61241, 16'd52877, 16'd53383, 16'd22876, 16'd52634, 16'd42306, 16'd24725, 16'd60638, 16'd5508, 16'd17938, 16'd20683, 16'd50646, 16'd19604, 16'd32210, 16'd31360, 16'd44306, 16'd23764, 16'd55798, 16'd11184, 16'd55372, 16'd31592, 16'd15744, 16'd37097});
	test_expansion(128'heaac876db213b668685ee6c7e76c8ffb, {16'd27187, 16'd21236, 16'd28047, 16'd782, 16'd11876, 16'd40898, 16'd49346, 16'd11557, 16'd2213, 16'd41360, 16'd1561, 16'd37999, 16'd31273, 16'd25430, 16'd28937, 16'd11779, 16'd47823, 16'd16179, 16'd11704, 16'd11743, 16'd31085, 16'd5062, 16'd46614, 16'd26127, 16'd16207, 16'd16841});
	test_expansion(128'h7e652a680a9aa7896d9e6776d508b4e7, {16'd41366, 16'd8138, 16'd669, 16'd22219, 16'd50002, 16'd45208, 16'd24229, 16'd46806, 16'd58567, 16'd30053, 16'd50087, 16'd15598, 16'd37967, 16'd64557, 16'd29389, 16'd4230, 16'd24315, 16'd31230, 16'd55614, 16'd4071, 16'd23122, 16'd23026, 16'd50114, 16'd1281, 16'd55029, 16'd14407});
	test_expansion(128'h614c4fd3e0bca4403fbcea950f1700be, {16'd31277, 16'd20328, 16'd13212, 16'd19507, 16'd20569, 16'd453, 16'd3074, 16'd55980, 16'd17686, 16'd41550, 16'd56174, 16'd34510, 16'd18965, 16'd6030, 16'd36364, 16'd30198, 16'd23060, 16'd20308, 16'd24029, 16'd44865, 16'd13882, 16'd22766, 16'd58041, 16'd32045, 16'd33347, 16'd49263});
	test_expansion(128'hed76df7482b63c891e0de172efc219ae, {16'd9335, 16'd20066, 16'd60352, 16'd34539, 16'd24139, 16'd4227, 16'd59369, 16'd22871, 16'd33511, 16'd41689, 16'd3422, 16'd8467, 16'd51362, 16'd60794, 16'd11759, 16'd60975, 16'd1673, 16'd8794, 16'd7025, 16'd53372, 16'd32530, 16'd57194, 16'd64244, 16'd28461, 16'd25086, 16'd29025});
	test_expansion(128'h01391070b30c7ef010426204a8168fd4, {16'd8674, 16'd50220, 16'd17051, 16'd48339, 16'd49815, 16'd852, 16'd21371, 16'd50586, 16'd50720, 16'd47054, 16'd13411, 16'd47450, 16'd12663, 16'd65012, 16'd54069, 16'd36532, 16'd37575, 16'd22618, 16'd40607, 16'd3396, 16'd28147, 16'd42696, 16'd42561, 16'd23875, 16'd2031, 16'd56211});
	test_expansion(128'h6629c0d27bede89e6eed86d53cbb06bf, {16'd65064, 16'd59214, 16'd33452, 16'd15147, 16'd4756, 16'd25854, 16'd32941, 16'd8588, 16'd21602, 16'd22910, 16'd47096, 16'd9809, 16'd47238, 16'd42446, 16'd18306, 16'd3084, 16'd29874, 16'd30290, 16'd18057, 16'd15244, 16'd64069, 16'd60774, 16'd43755, 16'd13746, 16'd52698, 16'd954});
	test_expansion(128'hd698b3eb484360022c09699c48fdec17, {16'd1901, 16'd40296, 16'd10330, 16'd12543, 16'd31353, 16'd22161, 16'd7495, 16'd62659, 16'd4986, 16'd64631, 16'd56859, 16'd34673, 16'd25108, 16'd56502, 16'd63961, 16'd50420, 16'd51303, 16'd16121, 16'd60879, 16'd7141, 16'd21019, 16'd29046, 16'd13414, 16'd45, 16'd63540, 16'd57415});
	test_expansion(128'hc0fbca0d1a1576f13a7cb74bb8663c63, {16'd61858, 16'd12456, 16'd44188, 16'd45645, 16'd42699, 16'd28246, 16'd33138, 16'd29831, 16'd15162, 16'd60951, 16'd47318, 16'd24983, 16'd60641, 16'd10262, 16'd64060, 16'd15388, 16'd28856, 16'd65230, 16'd1335, 16'd52702, 16'd15341, 16'd56378, 16'd13627, 16'd46346, 16'd10954, 16'd7047});
	test_expansion(128'hcac93c6162f95f7c7a0662bf7661076f, {16'd50072, 16'd13910, 16'd7690, 16'd61567, 16'd11385, 16'd25892, 16'd53927, 16'd24066, 16'd64395, 16'd19038, 16'd37320, 16'd2475, 16'd47110, 16'd31048, 16'd59797, 16'd24669, 16'd35088, 16'd5468, 16'd2933, 16'd28198, 16'd44733, 16'd15358, 16'd55949, 16'd47152, 16'd57512, 16'd23074});
	test_expansion(128'h0c798c5c9bd8e4b603563db7ca535071, {16'd7703, 16'd63510, 16'd47435, 16'd5252, 16'd55788, 16'd38466, 16'd47725, 16'd41046, 16'd24865, 16'd10315, 16'd2069, 16'd4740, 16'd7013, 16'd42675, 16'd54709, 16'd16378, 16'd17920, 16'd54510, 16'd31413, 16'd22747, 16'd48426, 16'd18328, 16'd52640, 16'd22166, 16'd52721, 16'd47971});
	test_expansion(128'h6287dc3114a38aae7eee0d091062a7e8, {16'd60720, 16'd36334, 16'd3106, 16'd13888, 16'd40617, 16'd39277, 16'd909, 16'd26676, 16'd64981, 16'd23792, 16'd8908, 16'd45139, 16'd49541, 16'd22825, 16'd7680, 16'd44482, 16'd40970, 16'd41606, 16'd26400, 16'd31518, 16'd22895, 16'd39085, 16'd19536, 16'd3975, 16'd30039, 16'd29386});
	test_expansion(128'h1e530b2ba49d5a1583a2b96d49f00d89, {16'd5897, 16'd18483, 16'd32839, 16'd24824, 16'd61660, 16'd10223, 16'd42732, 16'd21327, 16'd11803, 16'd34018, 16'd29652, 16'd60550, 16'd52846, 16'd58100, 16'd8585, 16'd24805, 16'd26686, 16'd9493, 16'd21682, 16'd16802, 16'd43034, 16'd24049, 16'd15195, 16'd29845, 16'd8283, 16'd37767});
	test_expansion(128'hc7bd806dab96c7f1ae48afce5be39948, {16'd17609, 16'd49648, 16'd23825, 16'd39229, 16'd19053, 16'd16038, 16'd65407, 16'd62738, 16'd54203, 16'd7318, 16'd20775, 16'd33874, 16'd23611, 16'd13138, 16'd46035, 16'd39871, 16'd13810, 16'd29438, 16'd45714, 16'd15521, 16'd33252, 16'd63625, 16'd49990, 16'd37322, 16'd24799, 16'd2185});
	test_expansion(128'h195ad54e021a982a19ac4af1d7202716, {16'd30135, 16'd50425, 16'd43358, 16'd65464, 16'd26326, 16'd26012, 16'd9447, 16'd49684, 16'd13201, 16'd54819, 16'd34237, 16'd54759, 16'd3369, 16'd63216, 16'd39304, 16'd30628, 16'd38558, 16'd18539, 16'd42981, 16'd44260, 16'd22028, 16'd3683, 16'd4758, 16'd52820, 16'd58394, 16'd64533});
	test_expansion(128'hb7db694532f95da8a923fdcc4e1554d9, {16'd15330, 16'd2504, 16'd45221, 16'd55690, 16'd58990, 16'd52002, 16'd50685, 16'd4559, 16'd20917, 16'd44780, 16'd30307, 16'd5985, 16'd7018, 16'd23194, 16'd43389, 16'd49026, 16'd58959, 16'd5835, 16'd56667, 16'd54581, 16'd56811, 16'd60869, 16'd19992, 16'd33566, 16'd37309, 16'd33834});
	test_expansion(128'ha747e9b4895d8507eabffc37e9f18f1b, {16'd6116, 16'd61558, 16'd59912, 16'd55495, 16'd39445, 16'd52793, 16'd37357, 16'd46744, 16'd23479, 16'd61412, 16'd3792, 16'd8390, 16'd2282, 16'd34986, 16'd48924, 16'd64893, 16'd56905, 16'd42584, 16'd25704, 16'd28719, 16'd48022, 16'd22006, 16'd27746, 16'd12953, 16'd50348, 16'd32118});
	test_expansion(128'h8abe70c47ff30aa5834ae613e821bd34, {16'd10724, 16'd24500, 16'd15383, 16'd32011, 16'd2664, 16'd42090, 16'd21898, 16'd9929, 16'd33764, 16'd45547, 16'd50414, 16'd27454, 16'd29122, 16'd41990, 16'd16745, 16'd44383, 16'd48663, 16'd2458, 16'd47520, 16'd61464, 16'd35335, 16'd9685, 16'd473, 16'd60220, 16'd47764, 16'd34517});
	test_expansion(128'h05bec2bb4a87d615d9c08df5010aa573, {16'd21328, 16'd7473, 16'd10355, 16'd42315, 16'd62955, 16'd21926, 16'd21199, 16'd3818, 16'd6695, 16'd46496, 16'd63025, 16'd64534, 16'd33938, 16'd44150, 16'd32809, 16'd15419, 16'd60669, 16'd61798, 16'd2572, 16'd29488, 16'd63587, 16'd29690, 16'd4724, 16'd48367, 16'd56532, 16'd12610});
	test_expansion(128'he7497f8e5f90e9640e2d216c67131c5e, {16'd26220, 16'd58121, 16'd17164, 16'd21112, 16'd52149, 16'd36094, 16'd14925, 16'd44972, 16'd4529, 16'd28434, 16'd6991, 16'd59564, 16'd25008, 16'd62848, 16'd54294, 16'd55433, 16'd16793, 16'd2629, 16'd40536, 16'd12611, 16'd1392, 16'd486, 16'd29678, 16'd19264, 16'd30873, 16'd18566});
	test_expansion(128'hb4b3c2dcbe7eb5cc756aacc3c5c45c2b, {16'd46342, 16'd31556, 16'd21069, 16'd52039, 16'd41912, 16'd29490, 16'd33393, 16'd15774, 16'd45071, 16'd30397, 16'd50138, 16'd15677, 16'd6854, 16'd27786, 16'd34009, 16'd44075, 16'd44837, 16'd3975, 16'd18823, 16'd61754, 16'd60512, 16'd42061, 16'd28634, 16'd15468, 16'd50610, 16'd5597});
	test_expansion(128'h1d617f1c2ae34f189132c600fe1b14ef, {16'd54811, 16'd36862, 16'd40263, 16'd9163, 16'd40172, 16'd32699, 16'd56370, 16'd1905, 16'd21692, 16'd60434, 16'd62551, 16'd21878, 16'd38074, 16'd37087, 16'd29415, 16'd17748, 16'd50170, 16'd60604, 16'd50660, 16'd63714, 16'd53860, 16'd42319, 16'd54149, 16'd28531, 16'd23762, 16'd47576});
	test_expansion(128'hd953bbab8857be9e6ba6e4050a4af4d6, {16'd16667, 16'd13300, 16'd40986, 16'd16135, 16'd30763, 16'd13841, 16'd40442, 16'd22682, 16'd2267, 16'd64564, 16'd49588, 16'd5740, 16'd12547, 16'd24880, 16'd51835, 16'd27863, 16'd10142, 16'd30127, 16'd16251, 16'd43790, 16'd65096, 16'd3523, 16'd53349, 16'd65513, 16'd12286, 16'd3152});
	test_expansion(128'hce75150d547cc8d4ab46d54cee3a70e8, {16'd7513, 16'd27278, 16'd15714, 16'd7224, 16'd60971, 16'd58123, 16'd10456, 16'd31848, 16'd6269, 16'd50879, 16'd10285, 16'd17831, 16'd24960, 16'd6941, 16'd8612, 16'd8611, 16'd38265, 16'd15707, 16'd15353, 16'd23159, 16'd47835, 16'd2828, 16'd6656, 16'd26957, 16'd6624, 16'd42533});
	test_expansion(128'hb6ad99558be8b2f4201007bc3f022f35, {16'd58006, 16'd33317, 16'd35685, 16'd35385, 16'd23393, 16'd28131, 16'd62731, 16'd59784, 16'd10185, 16'd3852, 16'd29042, 16'd37628, 16'd55437, 16'd11068, 16'd35025, 16'd21647, 16'd51682, 16'd11601, 16'd10402, 16'd65120, 16'd7382, 16'd45029, 16'd65121, 16'd49265, 16'd51819, 16'd28447});
	test_expansion(128'h9ddf0562d5411a611fe66165c902887f, {16'd2291, 16'd4160, 16'd57157, 16'd60638, 16'd56171, 16'd25615, 16'd51598, 16'd802, 16'd12027, 16'd33698, 16'd47650, 16'd61492, 16'd63217, 16'd41455, 16'd16237, 16'd65445, 16'd22226, 16'd49503, 16'd26188, 16'd45969, 16'd40297, 16'd53231, 16'd4934, 16'd16952, 16'd50644, 16'd24736});
	test_expansion(128'hca4940c0a0528767f9fc15138953a9c6, {16'd5549, 16'd9056, 16'd4663, 16'd41182, 16'd11717, 16'd13660, 16'd18396, 16'd36210, 16'd896, 16'd22100, 16'd41113, 16'd32122, 16'd29423, 16'd56212, 16'd45307, 16'd37527, 16'd426, 16'd22155, 16'd13559, 16'd289, 16'd50968, 16'd48701, 16'd21279, 16'd63612, 16'd59136, 16'd6517});
	test_expansion(128'h026ed9fd59fc6e48965820db2190944f, {16'd15710, 16'd60128, 16'd17084, 16'd22522, 16'd5391, 16'd28834, 16'd17695, 16'd4019, 16'd52430, 16'd42021, 16'd56761, 16'd18740, 16'd62467, 16'd48406, 16'd50679, 16'd8186, 16'd15227, 16'd4853, 16'd41651, 16'd16218, 16'd32160, 16'd13909, 16'd18515, 16'd26584, 16'd35826, 16'd57360});
	test_expansion(128'hafccea7aaed4dc2158990137402a1a29, {16'd14668, 16'd13953, 16'd30863, 16'd5063, 16'd39560, 16'd60572, 16'd51391, 16'd27565, 16'd9007, 16'd855, 16'd55108, 16'd4447, 16'd28916, 16'd28423, 16'd60595, 16'd29576, 16'd21855, 16'd10315, 16'd64038, 16'd40376, 16'd11230, 16'd20030, 16'd43276, 16'd52021, 16'd2869, 16'd41952});
	test_expansion(128'h1d75c6891b5d2af7320c3d1ac6990102, {16'd32633, 16'd53782, 16'd33438, 16'd63753, 16'd8981, 16'd13017, 16'd21083, 16'd7470, 16'd33729, 16'd6810, 16'd65227, 16'd31299, 16'd26869, 16'd43139, 16'd22764, 16'd64341, 16'd10253, 16'd4618, 16'd13312, 16'd15954, 16'd55067, 16'd10994, 16'd51977, 16'd59915, 16'd32897, 16'd4027});
	test_expansion(128'h2a4cc5dd9eaa74563ca339af7b9e8730, {16'd27051, 16'd62968, 16'd5166, 16'd12290, 16'd32721, 16'd7580, 16'd50042, 16'd12457, 16'd14243, 16'd13201, 16'd18509, 16'd55182, 16'd31599, 16'd45445, 16'd16173, 16'd23547, 16'd58922, 16'd16866, 16'd53303, 16'd14260, 16'd53345, 16'd31284, 16'd35751, 16'd35416, 16'd39113, 16'd33738});
	test_expansion(128'h50c6664f68b909db6a5b1a3f472caeaa, {16'd63966, 16'd30506, 16'd10190, 16'd21682, 16'd29098, 16'd45109, 16'd2699, 16'd12915, 16'd24459, 16'd28986, 16'd48849, 16'd28367, 16'd48097, 16'd27945, 16'd27172, 16'd21056, 16'd20166, 16'd8417, 16'd64330, 16'd4909, 16'd19778, 16'd42443, 16'd28648, 16'd8354, 16'd2905, 16'd25484});
	test_expansion(128'h1567bee0e59bbaea789cc6cbd3bcf6fd, {16'd51948, 16'd18149, 16'd39078, 16'd37095, 16'd49480, 16'd34836, 16'd40649, 16'd29176, 16'd63192, 16'd18883, 16'd46701, 16'd45452, 16'd61414, 16'd57550, 16'd62480, 16'd20227, 16'd49984, 16'd57945, 16'd40730, 16'd35939, 16'd58565, 16'd39444, 16'd31071, 16'd18535, 16'd9956, 16'd40083});
	test_expansion(128'hc4f1f1b97944f0d316614d6ce2e531d8, {16'd14486, 16'd42581, 16'd53155, 16'd54528, 16'd1085, 16'd38925, 16'd58061, 16'd13545, 16'd44277, 16'd52545, 16'd52591, 16'd59524, 16'd3315, 16'd56361, 16'd20682, 16'd64697, 16'd37586, 16'd23178, 16'd52800, 16'd27900, 16'd48745, 16'd31030, 16'd55254, 16'd50959, 16'd27185, 16'd24236});
	test_expansion(128'hc8b583b5bc756c00bcaf9d46e02d03cb, {16'd16920, 16'd12016, 16'd28250, 16'd3946, 16'd16101, 16'd51055, 16'd45625, 16'd38599, 16'd58030, 16'd30418, 16'd44835, 16'd63512, 16'd27639, 16'd40885, 16'd46174, 16'd63550, 16'd64149, 16'd62520, 16'd39496, 16'd1668, 16'd22210, 16'd22119, 16'd42573, 16'd22837, 16'd28000, 16'd52265});
	test_expansion(128'h506b236528e96319210f28b774cbc77f, {16'd31242, 16'd20970, 16'd1698, 16'd59229, 16'd23155, 16'd23188, 16'd46445, 16'd21215, 16'd62750, 16'd22662, 16'd29056, 16'd28896, 16'd38083, 16'd14676, 16'd20353, 16'd34641, 16'd49918, 16'd8126, 16'd9990, 16'd28138, 16'd43194, 16'd897, 16'd12830, 16'd27366, 16'd57105, 16'd18864});
	test_expansion(128'h50e0c9e96bedbb44e8a1660bacaf198a, {16'd39722, 16'd41627, 16'd40321, 16'd5980, 16'd26183, 16'd23182, 16'd11712, 16'd49224, 16'd8227, 16'd49109, 16'd19190, 16'd39312, 16'd2878, 16'd131, 16'd55453, 16'd61677, 16'd11619, 16'd46670, 16'd20073, 16'd29886, 16'd53069, 16'd19758, 16'd52501, 16'd21688, 16'd55389, 16'd56790});
	test_expansion(128'h5d280d88a22bf1182300d685604ca9f2, {16'd2973, 16'd51938, 16'd48097, 16'd55068, 16'd4126, 16'd63600, 16'd30273, 16'd51907, 16'd43151, 16'd10603, 16'd31978, 16'd26218, 16'd41818, 16'd35792, 16'd29089, 16'd32208, 16'd11714, 16'd1323, 16'd8655, 16'd41365, 16'd46712, 16'd27580, 16'd17907, 16'd10997, 16'd5299, 16'd64618});
	test_expansion(128'h8480baa294e93df91217c7f017abe437, {16'd50248, 16'd49492, 16'd8980, 16'd14806, 16'd24858, 16'd27124, 16'd10179, 16'd1426, 16'd1509, 16'd61248, 16'd19123, 16'd24210, 16'd21503, 16'd34233, 16'd45603, 16'd39848, 16'd50351, 16'd15278, 16'd43579, 16'd33508, 16'd56263, 16'd46132, 16'd32144, 16'd14172, 16'd58703, 16'd10710});
	test_expansion(128'hd8c8b582cee9be5087e7927a1f0b4caa, {16'd5717, 16'd47198, 16'd7989, 16'd44349, 16'd46889, 16'd47063, 16'd39804, 16'd65316, 16'd37732, 16'd55948, 16'd24182, 16'd39333, 16'd18009, 16'd49076, 16'd45037, 16'd57450, 16'd61382, 16'd40286, 16'd14236, 16'd62276, 16'd32529, 16'd36633, 16'd37956, 16'd19390, 16'd26341, 16'd1343});
	test_expansion(128'h9dc1fed1be377a3fdbc32dc49e3b8045, {16'd38970, 16'd57896, 16'd1279, 16'd24243, 16'd23865, 16'd38358, 16'd5856, 16'd15423, 16'd16824, 16'd42891, 16'd51200, 16'd64812, 16'd48494, 16'd14899, 16'd46354, 16'd52120, 16'd35225, 16'd43785, 16'd33342, 16'd3614, 16'd4250, 16'd55672, 16'd64818, 16'd12049, 16'd8469, 16'd55864});
	test_expansion(128'h06b8d712bf187db3134481e4d61ab955, {16'd39174, 16'd41388, 16'd37417, 16'd16638, 16'd36840, 16'd59356, 16'd26166, 16'd33811, 16'd703, 16'd16906, 16'd29504, 16'd58673, 16'd53414, 16'd60798, 16'd39309, 16'd10448, 16'd65468, 16'd6477, 16'd24358, 16'd47238, 16'd22087, 16'd44366, 16'd47020, 16'd48645, 16'd10394, 16'd4842});
	test_expansion(128'h0e0b026b0f0ff1858fd2d81b2c848c59, {16'd5143, 16'd39180, 16'd55725, 16'd33413, 16'd20305, 16'd55628, 16'd64128, 16'd13202, 16'd48431, 16'd43087, 16'd34623, 16'd23414, 16'd61084, 16'd61996, 16'd61000, 16'd3520, 16'd40283, 16'd52832, 16'd51484, 16'd42116, 16'd2224, 16'd38238, 16'd21248, 16'd37263, 16'd26949, 16'd60868});
	test_expansion(128'hc56fbecb0749fdd3e92ae8dc0a793b42, {16'd52771, 16'd38882, 16'd55234, 16'd63045, 16'd52529, 16'd40329, 16'd17363, 16'd32341, 16'd46926, 16'd14049, 16'd59602, 16'd39008, 16'd37290, 16'd21088, 16'd8383, 16'd40142, 16'd59875, 16'd55570, 16'd1243, 16'd45351, 16'd43070, 16'd43793, 16'd25747, 16'd35593, 16'd46188, 16'd45182});
	test_expansion(128'ha6ef9e3aa2b16951edcf4598e49ddb4b, {16'd35678, 16'd23105, 16'd59774, 16'd23844, 16'd63383, 16'd11883, 16'd48213, 16'd12175, 16'd55007, 16'd38725, 16'd45982, 16'd16594, 16'd8972, 16'd43657, 16'd10755, 16'd47947, 16'd47478, 16'd40770, 16'd39612, 16'd37421, 16'd40213, 16'd11942, 16'd21515, 16'd37661, 16'd61171, 16'd12553});
	test_expansion(128'h17bb8380519d456439ac49be8804db65, {16'd32227, 16'd19171, 16'd56931, 16'd54806, 16'd21454, 16'd47202, 16'd57394, 16'd2035, 16'd13696, 16'd36454, 16'd43560, 16'd51467, 16'd54262, 16'd10613, 16'd18267, 16'd56856, 16'd27069, 16'd59484, 16'd7813, 16'd17960, 16'd23455, 16'd28087, 16'd51084, 16'd2388, 16'd26470, 16'd18602});
	test_expansion(128'hb61fa13a94f8cf94dfacceda271c94ce, {16'd17916, 16'd17542, 16'd46118, 16'd29363, 16'd61436, 16'd8854, 16'd64788, 16'd41694, 16'd10813, 16'd56822, 16'd64515, 16'd33155, 16'd1181, 16'd47903, 16'd64227, 16'd33703, 16'd26008, 16'd20978, 16'd4432, 16'd52828, 16'd5936, 16'd19718, 16'd22648, 16'd56935, 16'd54596, 16'd2729});
	test_expansion(128'hd623543b3658bac118ad4834b5f31181, {16'd41217, 16'd42709, 16'd54284, 16'd22902, 16'd64044, 16'd7774, 16'd62882, 16'd46148, 16'd14770, 16'd59719, 16'd49235, 16'd9967, 16'd31788, 16'd16497, 16'd19719, 16'd31334, 16'd43466, 16'd55378, 16'd34402, 16'd27017, 16'd61460, 16'd44097, 16'd6819, 16'd41434, 16'd25028, 16'd52375});
	test_expansion(128'haeedfe1957d738d16f57ddd4e4b62311, {16'd1064, 16'd37468, 16'd46434, 16'd32433, 16'd56844, 16'd22558, 16'd10046, 16'd29397, 16'd18511, 16'd33585, 16'd59319, 16'd35753, 16'd55395, 16'd24739, 16'd61734, 16'd43867, 16'd54654, 16'd26304, 16'd709, 16'd36042, 16'd35509, 16'd61788, 16'd64026, 16'd62039, 16'd46220, 16'd33710});
	test_expansion(128'hb8f91dc82e447ab302b5a93dc031647b, {16'd11611, 16'd39020, 16'd24289, 16'd9201, 16'd7320, 16'd3065, 16'd15544, 16'd64734, 16'd20019, 16'd743, 16'd17193, 16'd9907, 16'd2297, 16'd54905, 16'd14166, 16'd60688, 16'd56745, 16'd16427, 16'd27297, 16'd16169, 16'd50964, 16'd6081, 16'd6229, 16'd47850, 16'd5748, 16'd7037});
	test_expansion(128'h92bb0d29d465787631d698baa60eb5a7, {16'd47018, 16'd47092, 16'd59850, 16'd44436, 16'd52393, 16'd42792, 16'd25842, 16'd2391, 16'd25897, 16'd27613, 16'd51282, 16'd34145, 16'd52471, 16'd14897, 16'd47177, 16'd6773, 16'd47250, 16'd28833, 16'd4876, 16'd14372, 16'd58666, 16'd4610, 16'd9815, 16'd22196, 16'd31785, 16'd40131});
	test_expansion(128'h72bd058b740a3fdb8553b1f19b2df62c, {16'd26715, 16'd13033, 16'd6543, 16'd55860, 16'd55178, 16'd26316, 16'd65372, 16'd14874, 16'd43927, 16'd33389, 16'd19238, 16'd61669, 16'd26277, 16'd37553, 16'd7523, 16'd17905, 16'd55838, 16'd31498, 16'd40806, 16'd6370, 16'd55177, 16'd7926, 16'd12137, 16'd47443, 16'd8679, 16'd33096});
	test_expansion(128'hb5d158d4812b590fcdd147d33e572315, {16'd39806, 16'd26833, 16'd31755, 16'd18559, 16'd59282, 16'd37813, 16'd60371, 16'd50552, 16'd16325, 16'd42379, 16'd557, 16'd57373, 16'd42592, 16'd61027, 16'd47835, 16'd24234, 16'd645, 16'd58622, 16'd19276, 16'd39844, 16'd37665, 16'd60356, 16'd19355, 16'd51747, 16'd16561, 16'd54093});
	test_expansion(128'h7a57d34f2a20c6c02ded8f08c5b70999, {16'd11893, 16'd35095, 16'd55283, 16'd41226, 16'd57419, 16'd62986, 16'd58092, 16'd55665, 16'd48859, 16'd45889, 16'd56804, 16'd1940, 16'd65349, 16'd4684, 16'd64268, 16'd60709, 16'd50242, 16'd20818, 16'd63060, 16'd21890, 16'd4533, 16'd13362, 16'd63612, 16'd18697, 16'd46860, 16'd43497});
	test_expansion(128'h28fac6a850b80d8833e5756f8b4bd363, {16'd64626, 16'd63558, 16'd18445, 16'd52621, 16'd44268, 16'd2899, 16'd1818, 16'd62380, 16'd931, 16'd25723, 16'd50221, 16'd9688, 16'd13240, 16'd15984, 16'd61173, 16'd43445, 16'd32897, 16'd8581, 16'd6997, 16'd53439, 16'd29423, 16'd1412, 16'd57845, 16'd25548, 16'd2092, 16'd25539});
	test_expansion(128'ha4a897ffd4a32de1e89d0e877b3abecd, {16'd9605, 16'd46319, 16'd20263, 16'd30830, 16'd22740, 16'd28884, 16'd50566, 16'd18080, 16'd27629, 16'd51176, 16'd37233, 16'd32829, 16'd61168, 16'd8959, 16'd61378, 16'd6460, 16'd15105, 16'd33320, 16'd7937, 16'd30755, 16'd61727, 16'd60358, 16'd33876, 16'd43117, 16'd29770, 16'd770});
	test_expansion(128'h2b82a1cf190f205fde7c6a6f694abdad, {16'd25691, 16'd1759, 16'd32423, 16'd11524, 16'd34231, 16'd55227, 16'd16766, 16'd53557, 16'd1899, 16'd15665, 16'd27617, 16'd38168, 16'd2475, 16'd32562, 16'd62471, 16'd65428, 16'd58944, 16'd55495, 16'd56821, 16'd10956, 16'd40343, 16'd59831, 16'd49484, 16'd26495, 16'd17123, 16'd5196});
	test_expansion(128'h08ae4851b068af951259acadfb2aa4bc, {16'd36619, 16'd25183, 16'd45200, 16'd48846, 16'd783, 16'd61673, 16'd51483, 16'd31484, 16'd2071, 16'd909, 16'd12320, 16'd138, 16'd46053, 16'd14515, 16'd2848, 16'd47438, 16'd20426, 16'd20867, 16'd35469, 16'd63862, 16'd20213, 16'd38237, 16'd5735, 16'd46838, 16'd49024, 16'd7620});
	test_expansion(128'hd6876ae6abe457d6f9cbbc0ea9fbac7d, {16'd2996, 16'd24091, 16'd57305, 16'd38981, 16'd12719, 16'd29132, 16'd8821, 16'd42147, 16'd31756, 16'd24746, 16'd4904, 16'd35353, 16'd14070, 16'd10492, 16'd23456, 16'd29998, 16'd26098, 16'd31057, 16'd13815, 16'd32834, 16'd21024, 16'd38450, 16'd317, 16'd50214, 16'd8915, 16'd14518});
	test_expansion(128'hf6e034693834168d365a3f7a68bcbca6, {16'd55633, 16'd3057, 16'd2682, 16'd3419, 16'd44050, 16'd18415, 16'd19666, 16'd44365, 16'd63903, 16'd46989, 16'd36589, 16'd6582, 16'd715, 16'd39981, 16'd31739, 16'd35818, 16'd17231, 16'd21568, 16'd47250, 16'd37749, 16'd31260, 16'd36157, 16'd19859, 16'd31405, 16'd15697, 16'd46450});
	test_expansion(128'h585bb30d67e26cf76c537d2651b6f4c2, {16'd53910, 16'd34351, 16'd18151, 16'd8548, 16'd54320, 16'd64225, 16'd8073, 16'd45743, 16'd8571, 16'd32901, 16'd5899, 16'd28834, 16'd11599, 16'd31741, 16'd15920, 16'd21401, 16'd54296, 16'd41244, 16'd52975, 16'd345, 16'd44712, 16'd41199, 16'd48220, 16'd19431, 16'd9433, 16'd4574});
	test_expansion(128'h9c23808f9f8826ec371e2ec3e5a8b564, {16'd57143, 16'd39841, 16'd47786, 16'd59169, 16'd4348, 16'd8514, 16'd12699, 16'd41366, 16'd35592, 16'd34081, 16'd65511, 16'd44915, 16'd348, 16'd37819, 16'd17992, 16'd50470, 16'd305, 16'd56388, 16'd32597, 16'd45040, 16'd4808, 16'd23961, 16'd48727, 16'd26078, 16'd64415, 16'd50691});
	test_expansion(128'h645629731c8534ba1ed5639fcb43f116, {16'd50804, 16'd5071, 16'd37625, 16'd22214, 16'd65389, 16'd3049, 16'd45797, 16'd27010, 16'd60297, 16'd53700, 16'd41560, 16'd17358, 16'd23874, 16'd7277, 16'd38228, 16'd51524, 16'd48907, 16'd56689, 16'd15926, 16'd25377, 16'd16730, 16'd31867, 16'd53154, 16'd32448, 16'd44906, 16'd30042});
	test_expansion(128'h798877a0b20c2e3be345a58853ac855b, {16'd357, 16'd3908, 16'd65066, 16'd24402, 16'd56590, 16'd64201, 16'd1672, 16'd109, 16'd43247, 16'd38502, 16'd2390, 16'd24400, 16'd16334, 16'd2939, 16'd57101, 16'd45582, 16'd12576, 16'd13696, 16'd53863, 16'd37334, 16'd58723, 16'd59674, 16'd31071, 16'd19960, 16'd10024, 16'd1339});
	test_expansion(128'hc294012af5a35844866009e944a7ab08, {16'd50349, 16'd44291, 16'd22691, 16'd38386, 16'd16735, 16'd14838, 16'd52710, 16'd64710, 16'd14801, 16'd31086, 16'd30488, 16'd55770, 16'd16507, 16'd37971, 16'd21863, 16'd7083, 16'd33581, 16'd40440, 16'd48615, 16'd32362, 16'd6214, 16'd10150, 16'd45097, 16'd33318, 16'd46020, 16'd45254});
	test_expansion(128'h1fc559d087e2d23bd98c4c94096a4fd5, {16'd2929, 16'd19373, 16'd50927, 16'd62733, 16'd23650, 16'd56716, 16'd57177, 16'd9250, 16'd52334, 16'd59310, 16'd56606, 16'd46605, 16'd18224, 16'd26578, 16'd2930, 16'd16496, 16'd44452, 16'd33559, 16'd22814, 16'd27640, 16'd55932, 16'd25883, 16'd21649, 16'd53064, 16'd37894, 16'd31796});
	test_expansion(128'h4e43728625074aecfa5c99e0a1e48a01, {16'd26879, 16'd14129, 16'd53166, 16'd95, 16'd41075, 16'd51194, 16'd19417, 16'd5390, 16'd25044, 16'd34667, 16'd45874, 16'd31138, 16'd43675, 16'd62571, 16'd57731, 16'd8906, 16'd13389, 16'd22622, 16'd51840, 16'd19283, 16'd9042, 16'd42563, 16'd46763, 16'd32600, 16'd14303, 16'd354});
	test_expansion(128'hbe23a24928600f381de86e96bd055351, {16'd53377, 16'd45461, 16'd1331, 16'd19111, 16'd33879, 16'd50248, 16'd36606, 16'd71, 16'd65002, 16'd51501, 16'd44976, 16'd60803, 16'd11457, 16'd44503, 16'd57007, 16'd17819, 16'd55465, 16'd7683, 16'd19420, 16'd23717, 16'd12035, 16'd56484, 16'd17118, 16'd64365, 16'd13402, 16'd34736});
	test_expansion(128'h3ae5ccd62b1ffedb5a680ec28c9f11d0, {16'd50082, 16'd51945, 16'd29022, 16'd18670, 16'd23126, 16'd16323, 16'd6663, 16'd24148, 16'd53196, 16'd54124, 16'd50500, 16'd8179, 16'd34860, 16'd22037, 16'd32924, 16'd35928, 16'd50141, 16'd36732, 16'd42155, 16'd40829, 16'd63937, 16'd63545, 16'd3555, 16'd13493, 16'd61536, 16'd45420});
	test_expansion(128'h2f31157767e6d0e979e8f7996268c6fa, {16'd29708, 16'd47282, 16'd21994, 16'd20937, 16'd19893, 16'd21311, 16'd29513, 16'd55830, 16'd5337, 16'd32515, 16'd45742, 16'd15212, 16'd24109, 16'd18545, 16'd19436, 16'd20258, 16'd51567, 16'd48923, 16'd56899, 16'd49616, 16'd3012, 16'd51704, 16'd62912, 16'd56409, 16'd56015, 16'd58469});
	test_expansion(128'h2d78973468c2207e8d4de983f5c2d455, {16'd7516, 16'd30492, 16'd12333, 16'd21795, 16'd43967, 16'd52490, 16'd24235, 16'd61255, 16'd23104, 16'd14262, 16'd3316, 16'd56113, 16'd7424, 16'd48323, 16'd33902, 16'd58069, 16'd22425, 16'd9960, 16'd50847, 16'd45366, 16'd7874, 16'd42229, 16'd12341, 16'd48253, 16'd24960, 16'd46200});
	test_expansion(128'ha3b54d4f98dcbdb5bc38690e108a2b13, {16'd44802, 16'd6426, 16'd58682, 16'd61440, 16'd640, 16'd25257, 16'd43431, 16'd12304, 16'd38420, 16'd33256, 16'd37437, 16'd22836, 16'd23955, 16'd1690, 16'd33299, 16'd61334, 16'd11109, 16'd60321, 16'd43743, 16'd51836, 16'd58941, 16'd28074, 16'd29933, 16'd12227, 16'd19727, 16'd58765});
	test_expansion(128'haa6c413b9c9fb4cf5d2272d9253fbd41, {16'd40682, 16'd1532, 16'd16851, 16'd40458, 16'd12769, 16'd971, 16'd53066, 16'd21173, 16'd62697, 16'd49455, 16'd35771, 16'd59286, 16'd45223, 16'd3020, 16'd10194, 16'd42654, 16'd16988, 16'd63150, 16'd431, 16'd18199, 16'd28844, 16'd63365, 16'd52357, 16'd11002, 16'd9222, 16'd16143});
	test_expansion(128'h6a68638ca65b651044edecd1fd9fd032, {16'd17150, 16'd18675, 16'd31344, 16'd59567, 16'd1506, 16'd50631, 16'd45382, 16'd33812, 16'd27575, 16'd54248, 16'd11411, 16'd61227, 16'd24470, 16'd38865, 16'd41638, 16'd53329, 16'd56832, 16'd59961, 16'd32604, 16'd35136, 16'd30208, 16'd50931, 16'd5188, 16'd53885, 16'd63378, 16'd43687});
	test_expansion(128'h72914726d26451666bcf832a2f351869, {16'd44192, 16'd15681, 16'd52419, 16'd671, 16'd8949, 16'd12308, 16'd55656, 16'd56142, 16'd37021, 16'd62146, 16'd32372, 16'd27853, 16'd507, 16'd40306, 16'd30684, 16'd32089, 16'd63223, 16'd64893, 16'd18113, 16'd30537, 16'd59011, 16'd21244, 16'd403, 16'd29674, 16'd20127, 16'd48246});
	test_expansion(128'h5776c27a68269490ce26c8ee632afc8c, {16'd63529, 16'd58400, 16'd29387, 16'd40907, 16'd29871, 16'd5381, 16'd51355, 16'd61717, 16'd44964, 16'd57011, 16'd8070, 16'd59283, 16'd1738, 16'd63853, 16'd42333, 16'd63898, 16'd27988, 16'd17463, 16'd44884, 16'd3009, 16'd16841, 16'd29900, 16'd48354, 16'd45300, 16'd39093, 16'd27630});
	test_expansion(128'hc128bd5d47c3d7c8659c53599f5dc1bc, {16'd57617, 16'd28693, 16'd54460, 16'd41401, 16'd14418, 16'd31253, 16'd48113, 16'd61564, 16'd34638, 16'd62080, 16'd11984, 16'd38447, 16'd48228, 16'd63788, 16'd47542, 16'd61491, 16'd22252, 16'd15240, 16'd65365, 16'd44977, 16'd10306, 16'd8459, 16'd54904, 16'd15455, 16'd45133, 16'd17112});
	test_expansion(128'h9abf545d6b2d1979dbcf5c210ab59592, {16'd21497, 16'd21912, 16'd59514, 16'd60813, 16'd15955, 16'd3055, 16'd5965, 16'd22426, 16'd21202, 16'd60767, 16'd53739, 16'd37330, 16'd20249, 16'd6900, 16'd61536, 16'd39521, 16'd32932, 16'd4571, 16'd47948, 16'd58281, 16'd33420, 16'd34240, 16'd47098, 16'd37871, 16'd1046, 16'd35689});
	test_expansion(128'h104e323b749423554d692bc9ef7fcf5c, {16'd14750, 16'd11727, 16'd2316, 16'd23182, 16'd21883, 16'd44870, 16'd36620, 16'd56237, 16'd46216, 16'd11447, 16'd15621, 16'd30873, 16'd59883, 16'd56631, 16'd15587, 16'd64704, 16'd54619, 16'd27326, 16'd46047, 16'd35053, 16'd44977, 16'd42105, 16'd27960, 16'd42851, 16'd41973, 16'd16091});
	test_expansion(128'hf1bf3009f2deb1bbc1be6f96c5119994, {16'd44849, 16'd61864, 16'd56934, 16'd28759, 16'd34312, 16'd62976, 16'd47360, 16'd39982, 16'd2232, 16'd27221, 16'd31044, 16'd39835, 16'd63984, 16'd27028, 16'd27332, 16'd30669, 16'd43393, 16'd18448, 16'd6770, 16'd13300, 16'd63746, 16'd53654, 16'd62639, 16'd23273, 16'd61708, 16'd55851});
	test_expansion(128'hd8e809d9457204d94ad849396ee63570, {16'd36238, 16'd1151, 16'd54386, 16'd11267, 16'd45627, 16'd60400, 16'd60286, 16'd19477, 16'd33161, 16'd58293, 16'd49342, 16'd27166, 16'd63448, 16'd30297, 16'd26990, 16'd62628, 16'd7576, 16'd34840, 16'd41647, 16'd49652, 16'd33441, 16'd32390, 16'd32337, 16'd46587, 16'd39530, 16'd57489});
	test_expansion(128'h55ff90ac7b2fdab16409bb0bbe0f2d1f, {16'd63417, 16'd40687, 16'd16731, 16'd59796, 16'd28326, 16'd36141, 16'd46861, 16'd29162, 16'd9548, 16'd39571, 16'd59460, 16'd5602, 16'd3318, 16'd2661, 16'd5963, 16'd47392, 16'd25360, 16'd54356, 16'd5013, 16'd45081, 16'd41025, 16'd4326, 16'd19666, 16'd14368, 16'd49175, 16'd12773});
	test_expansion(128'hf6510a5f1d019a9428861969bca7fe44, {16'd42859, 16'd49121, 16'd60686, 16'd63511, 16'd22083, 16'd48272, 16'd21731, 16'd9652, 16'd62295, 16'd40843, 16'd20378, 16'd40765, 16'd9172, 16'd34067, 16'd43108, 16'd9532, 16'd22916, 16'd39165, 16'd13469, 16'd35560, 16'd8310, 16'd32249, 16'd62606, 16'd49970, 16'd5146, 16'd17780});
	test_expansion(128'h8a3add5403cb1ee9d30cdfabedbe37db, {16'd25995, 16'd64914, 16'd64143, 16'd43517, 16'd3663, 16'd45438, 16'd60038, 16'd45855, 16'd16319, 16'd28170, 16'd56533, 16'd17460, 16'd61135, 16'd19068, 16'd20623, 16'd6480, 16'd20144, 16'd13723, 16'd39911, 16'd63967, 16'd21513, 16'd22961, 16'd12284, 16'd22792, 16'd12165, 16'd11314});
	test_expansion(128'h2a553a0a1dc5ab3c90c448fa2b33c7bc, {16'd18365, 16'd52642, 16'd48072, 16'd43271, 16'd30879, 16'd29978, 16'd40990, 16'd62285, 16'd39571, 16'd30268, 16'd54658, 16'd42255, 16'd43270, 16'd42243, 16'd24645, 16'd36109, 16'd13394, 16'd32010, 16'd62730, 16'd15582, 16'd16208, 16'd38044, 16'd41579, 16'd10708, 16'd19787, 16'd25952});
	test_expansion(128'h1c6c49412c21cc92b3adb5d206cf3a47, {16'd5765, 16'd17103, 16'd30002, 16'd62015, 16'd55452, 16'd60772, 16'd12873, 16'd42399, 16'd56991, 16'd29761, 16'd45357, 16'd8282, 16'd10168, 16'd56260, 16'd58240, 16'd54980, 16'd53184, 16'd49466, 16'd42313, 16'd58946, 16'd17338, 16'd47816, 16'd45206, 16'd23668, 16'd56558, 16'd24182});
	test_expansion(128'h51f80ca4a82bc5f06061093f0fb88b96, {16'd10004, 16'd13867, 16'd26076, 16'd25261, 16'd6015, 16'd35908, 16'd52793, 16'd20844, 16'd13186, 16'd32189, 16'd16878, 16'd57139, 16'd43356, 16'd18985, 16'd23195, 16'd19992, 16'd40377, 16'd64432, 16'd64960, 16'd45433, 16'd26200, 16'd50761, 16'd46869, 16'd29677, 16'd54207, 16'd17481});
	test_expansion(128'h63883aa1fd58021c671c2f6b888d5eea, {16'd53042, 16'd32684, 16'd54318, 16'd13569, 16'd26029, 16'd21295, 16'd49478, 16'd60862, 16'd36780, 16'd53447, 16'd42961, 16'd43318, 16'd55232, 16'd18176, 16'd27979, 16'd59524, 16'd57208, 16'd20196, 16'd317, 16'd15986, 16'd54529, 16'd8616, 16'd24778, 16'd62922, 16'd22161, 16'd3503});
	test_expansion(128'h9bb9241123e617e82c4acc5252f4cab4, {16'd51586, 16'd41331, 16'd12031, 16'd46555, 16'd46238, 16'd22574, 16'd61536, 16'd28930, 16'd45874, 16'd51222, 16'd40632, 16'd48491, 16'd23612, 16'd52912, 16'd1134, 16'd62312, 16'd35180, 16'd10245, 16'd49643, 16'd10723, 16'd32788, 16'd30154, 16'd64784, 16'd41916, 16'd37106, 16'd13807});
	test_expansion(128'heb6d599429d09d6f97ff9e5c39820e6a, {16'd12625, 16'd31202, 16'd4690, 16'd49176, 16'd28476, 16'd15488, 16'd46170, 16'd451, 16'd49367, 16'd47409, 16'd558, 16'd38600, 16'd3661, 16'd26767, 16'd46543, 16'd42203, 16'd56583, 16'd21223, 16'd15094, 16'd29709, 16'd15802, 16'd45695, 16'd7670, 16'd30047, 16'd19252, 16'd43861});
	test_expansion(128'hb3944b5725d0467fa705c21b39f8e8c4, {16'd62137, 16'd17518, 16'd52546, 16'd32760, 16'd46569, 16'd23654, 16'd29270, 16'd60506, 16'd61310, 16'd20293, 16'd414, 16'd53408, 16'd3071, 16'd36420, 16'd51049, 16'd46719, 16'd8884, 16'd13932, 16'd10221, 16'd63507, 16'd23642, 16'd983, 16'd12714, 16'd2055, 16'd26470, 16'd49311});
	test_expansion(128'h947f061d6262f819ea421d05dd9d77a0, {16'd64294, 16'd64903, 16'd24671, 16'd42409, 16'd36156, 16'd30743, 16'd45830, 16'd60036, 16'd23514, 16'd43606, 16'd30948, 16'd57602, 16'd36606, 16'd15578, 16'd47304, 16'd46666, 16'd17658, 16'd62293, 16'd64911, 16'd33139, 16'd23317, 16'd48209, 16'd32123, 16'd63106, 16'd45970, 16'd49274});
	test_expansion(128'h941c8e0492ff42642957abe3b9bb9e92, {16'd41941, 16'd29044, 16'd10537, 16'd38442, 16'd41994, 16'd42056, 16'd3857, 16'd27925, 16'd31070, 16'd42065, 16'd61437, 16'd45938, 16'd51168, 16'd55604, 16'd21297, 16'd56986, 16'd19195, 16'd40136, 16'd47625, 16'd27649, 16'd28599, 16'd32304, 16'd8219, 16'd25789, 16'd57218, 16'd37815});
	test_expansion(128'hfc2cd4b5c7a4f4c64e174e58892456b1, {16'd40813, 16'd10715, 16'd24636, 16'd52888, 16'd58324, 16'd43677, 16'd60532, 16'd59359, 16'd50931, 16'd15365, 16'd64695, 16'd63879, 16'd28377, 16'd10730, 16'd7081, 16'd21894, 16'd19615, 16'd48079, 16'd38806, 16'd21487, 16'd50223, 16'd54705, 16'd64663, 16'd53129, 16'd62227, 16'd33128});
	test_expansion(128'h89e87bdcdb44d41781652969bf4fde9e, {16'd12471, 16'd36094, 16'd49647, 16'd9526, 16'd46176, 16'd9946, 16'd40697, 16'd43349, 16'd58342, 16'd6934, 16'd40930, 16'd22874, 16'd17452, 16'd18056, 16'd18185, 16'd17458, 16'd36229, 16'd6908, 16'd11809, 16'd15939, 16'd42305, 16'd48757, 16'd46492, 16'd55820, 16'd18784, 16'd30305});
	test_expansion(128'h60a123a90c112a15da953322973706bd, {16'd53183, 16'd19442, 16'd49342, 16'd46876, 16'd57951, 16'd38843, 16'd21191, 16'd33674, 16'd57941, 16'd17123, 16'd12503, 16'd47758, 16'd54520, 16'd2004, 16'd12834, 16'd34151, 16'd48609, 16'd3084, 16'd3761, 16'd63106, 16'd31676, 16'd4192, 16'd62652, 16'd47631, 16'd28129, 16'd61916});
	test_expansion(128'hf2e064d979379a2ad9a5217668b1e885, {16'd19550, 16'd8464, 16'd799, 16'd25970, 16'd10465, 16'd51402, 16'd53596, 16'd23209, 16'd52630, 16'd56479, 16'd60247, 16'd50383, 16'd25160, 16'd53270, 16'd35851, 16'd32087, 16'd61257, 16'd30438, 16'd4466, 16'd58352, 16'd55517, 16'd29802, 16'd24506, 16'd57185, 16'd22799, 16'd57734});
	test_expansion(128'h352e37f471c8488a7d4b5e5990a92020, {16'd7957, 16'd31432, 16'd17132, 16'd15227, 16'd41098, 16'd40165, 16'd17524, 16'd47934, 16'd57280, 16'd55363, 16'd24518, 16'd24065, 16'd62104, 16'd39784, 16'd1556, 16'd12142, 16'd14504, 16'd65436, 16'd16987, 16'd30674, 16'd20988, 16'd17511, 16'd45511, 16'd63283, 16'd46891, 16'd36776});
	test_expansion(128'h62a706ffedc888b3a5176cf5d72cdd7f, {16'd9949, 16'd13551, 16'd45273, 16'd48880, 16'd32498, 16'd7565, 16'd41275, 16'd51138, 16'd11557, 16'd10421, 16'd36234, 16'd4296, 16'd63379, 16'd47350, 16'd4181, 16'd9397, 16'd37890, 16'd726, 16'd31685, 16'd50225, 16'd48264, 16'd30730, 16'd55887, 16'd30901, 16'd15731, 16'd59311});
	test_expansion(128'hd1401c663822da1d7305407c2a461458, {16'd40958, 16'd41682, 16'd58944, 16'd42476, 16'd10067, 16'd7386, 16'd29218, 16'd38794, 16'd13165, 16'd1406, 16'd35297, 16'd58975, 16'd33081, 16'd45838, 16'd4026, 16'd34765, 16'd23469, 16'd57489, 16'd46922, 16'd22991, 16'd48603, 16'd50560, 16'd44201, 16'd50364, 16'd52616, 16'd36112});
	test_expansion(128'hba589bdf2ccc0542546706e5c5ebe4bc, {16'd49151, 16'd13934, 16'd64990, 16'd30896, 16'd61171, 16'd9617, 16'd7591, 16'd30704, 16'd7930, 16'd16996, 16'd49534, 16'd46318, 16'd21245, 16'd60450, 16'd14375, 16'd1643, 16'd60062, 16'd56259, 16'd0, 16'd18122, 16'd58827, 16'd14286, 16'd33036, 16'd11899, 16'd59620, 16'd13668});
	test_expansion(128'hf287448ddd6061bd1c5b5e60c987f98e, {16'd55205, 16'd42245, 16'd33154, 16'd38877, 16'd37310, 16'd28694, 16'd37110, 16'd16442, 16'd42510, 16'd51812, 16'd4960, 16'd61572, 16'd7467, 16'd47941, 16'd51817, 16'd29722, 16'd48898, 16'd9546, 16'd32779, 16'd62166, 16'd11544, 16'd54169, 16'd30508, 16'd37700, 16'd64027, 16'd44504});
	test_expansion(128'h391ebfa5dab91b2e8f7672b56f7d32c0, {16'd45202, 16'd13919, 16'd1308, 16'd60794, 16'd44813, 16'd37407, 16'd26777, 16'd53677, 16'd40735, 16'd40401, 16'd62592, 16'd46400, 16'd63373, 16'd20765, 16'd30055, 16'd58917, 16'd33078, 16'd4894, 16'd5648, 16'd7686, 16'd56899, 16'd42116, 16'd318, 16'd48455, 16'd17498, 16'd60152});
	test_expansion(128'h02c3dc194ebfd05a571a7a23b13e112a, {16'd47309, 16'd60317, 16'd47974, 16'd38595, 16'd700, 16'd50662, 16'd40564, 16'd26028, 16'd3373, 16'd54359, 16'd24194, 16'd54868, 16'd1902, 16'd43984, 16'd25582, 16'd55826, 16'd35936, 16'd58407, 16'd18965, 16'd41421, 16'd3416, 16'd27011, 16'd27757, 16'd23740, 16'd4278, 16'd44709});
	test_expansion(128'h8814e82535af278dcfc0ac9ff0c98b1f, {16'd9840, 16'd61223, 16'd51791, 16'd6423, 16'd16152, 16'd35335, 16'd6101, 16'd49413, 16'd38899, 16'd40814, 16'd25212, 16'd53608, 16'd27425, 16'd44710, 16'd42066, 16'd37295, 16'd67, 16'd62221, 16'd31202, 16'd20969, 16'd31774, 16'd27732, 16'd12494, 16'd39297, 16'd49640, 16'd2458});
	test_expansion(128'hc5230423246e48310c28f520d3d8ed39, {16'd13662, 16'd16749, 16'd16690, 16'd13274, 16'd23171, 16'd55511, 16'd41510, 16'd544, 16'd23446, 16'd19955, 16'd54599, 16'd44022, 16'd46431, 16'd12434, 16'd52719, 16'd58543, 16'd62435, 16'd26814, 16'd31310, 16'd11631, 16'd24643, 16'd18883, 16'd51707, 16'd61282, 16'd50699, 16'd37546});
	test_expansion(128'h676b0ad483613231e3ef9b7124833cbe, {16'd13804, 16'd32739, 16'd64712, 16'd29727, 16'd8422, 16'd58873, 16'd34375, 16'd41829, 16'd24582, 16'd58041, 16'd46391, 16'd62300, 16'd8247, 16'd27021, 16'd25036, 16'd15613, 16'd60504, 16'd8146, 16'd32110, 16'd33098, 16'd63436, 16'd3311, 16'd59532, 16'd12911, 16'd3117, 16'd50293});
	test_expansion(128'h5cdd88838a4bc478917a7744b4436e80, {16'd59320, 16'd26912, 16'd9226, 16'd14420, 16'd55888, 16'd6061, 16'd15468, 16'd64714, 16'd988, 16'd57802, 16'd23921, 16'd14658, 16'd23821, 16'd15106, 16'd60403, 16'd22529, 16'd6476, 16'd25310, 16'd59981, 16'd43424, 16'd46632, 16'd60107, 16'd50702, 16'd64281, 16'd28932, 16'd32100});
	test_expansion(128'h02617dc8262e5c785bd993b59d990f27, {16'd26523, 16'd61571, 16'd22096, 16'd58146, 16'd12496, 16'd51993, 16'd41467, 16'd15323, 16'd4712, 16'd34561, 16'd11508, 16'd16337, 16'd1050, 16'd34786, 16'd35123, 16'd51872, 16'd41266, 16'd59552, 16'd42431, 16'd37356, 16'd48082, 16'd57090, 16'd53066, 16'd61356, 16'd49696, 16'd3375});
	test_expansion(128'hea9f67ec4886a89bcf9f17bf80dd60c3, {16'd23612, 16'd42717, 16'd53448, 16'd19808, 16'd59327, 16'd3771, 16'd17012, 16'd40950, 16'd25239, 16'd47056, 16'd38780, 16'd61183, 16'd2097, 16'd47067, 16'd23278, 16'd49912, 16'd36668, 16'd55967, 16'd52999, 16'd24130, 16'd50731, 16'd43012, 16'd58496, 16'd30412, 16'd6540, 16'd33490});
	test_expansion(128'h33effd6e7a7d26523138e1bbbd3df3e0, {16'd31789, 16'd61728, 16'd55641, 16'd56959, 16'd23329, 16'd48073, 16'd20994, 16'd36289, 16'd46210, 16'd22046, 16'd26228, 16'd16354, 16'd63542, 16'd49601, 16'd22113, 16'd26557, 16'd25341, 16'd19128, 16'd60339, 16'd20560, 16'd11486, 16'd50937, 16'd62986, 16'd904, 16'd49578, 16'd21205});
	test_expansion(128'h7c71332be8e813b4180e031acbde267e, {16'd50101, 16'd18788, 16'd25639, 16'd32628, 16'd304, 16'd9341, 16'd29970, 16'd14698, 16'd61334, 16'd57391, 16'd793, 16'd57790, 16'd12790, 16'd32699, 16'd43042, 16'd55210, 16'd32746, 16'd4384, 16'd31898, 16'd54963, 16'd19821, 16'd15522, 16'd21154, 16'd64453, 16'd5105, 16'd40986});
	test_expansion(128'h61b07b37968cecb2d0520607100c2d56, {16'd30990, 16'd13477, 16'd6363, 16'd54366, 16'd22310, 16'd17879, 16'd48862, 16'd61952, 16'd36146, 16'd61906, 16'd59951, 16'd21965, 16'd26945, 16'd42939, 16'd64730, 16'd44895, 16'd57801, 16'd54672, 16'd7143, 16'd25563, 16'd19222, 16'd46900, 16'd27203, 16'd59143, 16'd45066, 16'd12801});
	test_expansion(128'h11a8e67e147ead4f86e6c6427b2949a8, {16'd37635, 16'd11857, 16'd47302, 16'd50838, 16'd58301, 16'd39259, 16'd48090, 16'd29705, 16'd36026, 16'd39709, 16'd25542, 16'd30654, 16'd11207, 16'd58508, 16'd19349, 16'd61336, 16'd29111, 16'd46675, 16'd33374, 16'd27566, 16'd30455, 16'd34635, 16'd7449, 16'd11616, 16'd37910, 16'd54906});
	test_expansion(128'h69cdca3c2f83538880c32d53eac3d66d, {16'd24823, 16'd42379, 16'd12684, 16'd60832, 16'd22412, 16'd52770, 16'd45542, 16'd10800, 16'd32824, 16'd62169, 16'd58545, 16'd29680, 16'd36487, 16'd41804, 16'd17593, 16'd22321, 16'd10250, 16'd20299, 16'd64802, 16'd31992, 16'd30798, 16'd35291, 16'd49822, 16'd54503, 16'd27511, 16'd54750});
	test_expansion(128'h60d9e8884a23006d88fd50af41d709ff, {16'd55228, 16'd20403, 16'd39845, 16'd39440, 16'd39488, 16'd3087, 16'd9189, 16'd52570, 16'd10770, 16'd5489, 16'd43741, 16'd7246, 16'd19810, 16'd52721, 16'd52678, 16'd9441, 16'd33756, 16'd50472, 16'd35000, 16'd32187, 16'd48066, 16'd2139, 16'd32251, 16'd40084, 16'd50602, 16'd20791});
	test_expansion(128'h2cb36d02e304be03fed3ce0f23defbbb, {16'd15641, 16'd2219, 16'd17759, 16'd17841, 16'd41572, 16'd12425, 16'd1530, 16'd25563, 16'd46203, 16'd50304, 16'd18167, 16'd38601, 16'd35884, 16'd39349, 16'd64446, 16'd33275, 16'd20062, 16'd44551, 16'd51186, 16'd42341, 16'd17436, 16'd7829, 16'd12963, 16'd40702, 16'd19655, 16'd1499});
	test_expansion(128'h0ee34dabbe4833e903ac9402142794ef, {16'd64520, 16'd9035, 16'd45438, 16'd1912, 16'd28400, 16'd62384, 16'd50563, 16'd46550, 16'd57880, 16'd44613, 16'd65135, 16'd7669, 16'd25478, 16'd32358, 16'd16033, 16'd62221, 16'd57672, 16'd22974, 16'd36381, 16'd8548, 16'd38106, 16'd46973, 16'd32634, 16'd52205, 16'd23174, 16'd37846});
	test_expansion(128'hc74e22bc3d39281487b66b3f7c0585e6, {16'd56083, 16'd27395, 16'd29085, 16'd58475, 16'd41346, 16'd17375, 16'd6284, 16'd24109, 16'd49678, 16'd24533, 16'd23188, 16'd29776, 16'd11518, 16'd24631, 16'd61296, 16'd57336, 16'd24444, 16'd12083, 16'd18888, 16'd42575, 16'd2733, 16'd13741, 16'd2745, 16'd29462, 16'd62289, 16'd43969});
	test_expansion(128'h2d48a090dfbe37730bdc600a97e0d558, {16'd21044, 16'd50745, 16'd25170, 16'd23355, 16'd38524, 16'd32105, 16'd52226, 16'd11718, 16'd6404, 16'd9316, 16'd60064, 16'd6190, 16'd488, 16'd33379, 16'd11069, 16'd20334, 16'd40642, 16'd29754, 16'd40853, 16'd37841, 16'd47688, 16'd5591, 16'd274, 16'd17470, 16'd36701, 16'd6613});
	test_expansion(128'ha2b327fdc27cda2b52567ce4b06c6123, {16'd22671, 16'd17205, 16'd28095, 16'd1545, 16'd52526, 16'd63944, 16'd42347, 16'd13054, 16'd31747, 16'd46079, 16'd3610, 16'd58664, 16'd43774, 16'd38720, 16'd4055, 16'd8527, 16'd26900, 16'd7986, 16'd34033, 16'd42342, 16'd40467, 16'd65218, 16'd32012, 16'd60592, 16'd18377, 16'd2959});
	test_expansion(128'h8d4679d87d7fb2ec2d1603cc2056239f, {16'd30479, 16'd2335, 16'd18642, 16'd27465, 16'd41891, 16'd57245, 16'd47196, 16'd54510, 16'd17373, 16'd48657, 16'd48457, 16'd29560, 16'd7666, 16'd59969, 16'd9214, 16'd35806, 16'd48267, 16'd15710, 16'd10718, 16'd3734, 16'd54305, 16'd5717, 16'd11227, 16'd4461, 16'd40453, 16'd2032});
	test_expansion(128'hfe6a4aad31a3e6385abdb209e381ec17, {16'd7493, 16'd59097, 16'd12050, 16'd60508, 16'd12576, 16'd12830, 16'd32107, 16'd21268, 16'd25000, 16'd6329, 16'd41274, 16'd7043, 16'd18467, 16'd32607, 16'd22447, 16'd6990, 16'd51318, 16'd1667, 16'd42776, 16'd19647, 16'd50011, 16'd21209, 16'd33866, 16'd55944, 16'd10486, 16'd30146});
	test_expansion(128'h87db4318e73934c798f5c072953a32c4, {16'd4347, 16'd23400, 16'd19647, 16'd34805, 16'd53721, 16'd14953, 16'd43038, 16'd57533, 16'd31752, 16'd62410, 16'd54464, 16'd65314, 16'd19790, 16'd45445, 16'd31338, 16'd18359, 16'd29632, 16'd45367, 16'd63354, 16'd32286, 16'd31620, 16'd41242, 16'd29068, 16'd43360, 16'd49426, 16'd5646});
	test_expansion(128'hfc981ebd7867ba367736e9202b0ad662, {16'd31330, 16'd29710, 16'd23902, 16'd47042, 16'd16684, 16'd12478, 16'd54808, 16'd60640, 16'd7723, 16'd17804, 16'd20930, 16'd35374, 16'd52803, 16'd20466, 16'd42755, 16'd5551, 16'd40507, 16'd420, 16'd36381, 16'd4155, 16'd5847, 16'd23278, 16'd22751, 16'd37105, 16'd15475, 16'd44518});
	test_expansion(128'hdbd377a03a81c561374c7a6bb9a30fa3, {16'd26303, 16'd34678, 16'd48856, 16'd40303, 16'd27401, 16'd8053, 16'd27103, 16'd49608, 16'd45580, 16'd62011, 16'd23263, 16'd31532, 16'd51652, 16'd28214, 16'd39717, 16'd28391, 16'd58077, 16'd43926, 16'd20622, 16'd5582, 16'd13272, 16'd13982, 16'd3829, 16'd17167, 16'd25906, 16'd17382});
	test_expansion(128'h6302a3cdb15e177eca9b43bd3dccadb9, {16'd14783, 16'd41509, 16'd29820, 16'd57547, 16'd44891, 16'd38303, 16'd62837, 16'd356, 16'd52083, 16'd57572, 16'd4371, 16'd26391, 16'd22052, 16'd14540, 16'd1861, 16'd19771, 16'd50652, 16'd39448, 16'd7897, 16'd34210, 16'd23963, 16'd41132, 16'd11395, 16'd18427, 16'd26833, 16'd1802});
	test_expansion(128'h7be24c6e0b06194a63b4fb37161a348c, {16'd6952, 16'd49420, 16'd60863, 16'd25260, 16'd52305, 16'd21798, 16'd46043, 16'd12655, 16'd3481, 16'd35259, 16'd44784, 16'd22004, 16'd15401, 16'd58727, 16'd57525, 16'd30105, 16'd13869, 16'd59001, 16'd37938, 16'd34385, 16'd56020, 16'd32334, 16'd63571, 16'd42294, 16'd12780, 16'd7875});
	test_expansion(128'hfd76378a1efada7ace01696bd4c0c421, {16'd26010, 16'd3679, 16'd45472, 16'd22813, 16'd11419, 16'd11422, 16'd33079, 16'd45903, 16'd52326, 16'd44798, 16'd34632, 16'd36649, 16'd52381, 16'd59539, 16'd7458, 16'd9146, 16'd55155, 16'd11405, 16'd59486, 16'd63067, 16'd46776, 16'd26049, 16'd44522, 16'd51301, 16'd61131, 16'd2034});
	test_expansion(128'h567e172d6008b597d2e0246b65cdefd2, {16'd31808, 16'd37766, 16'd40345, 16'd21888, 16'd13060, 16'd2916, 16'd58241, 16'd18031, 16'd35540, 16'd16991, 16'd31574, 16'd60455, 16'd21174, 16'd31595, 16'd27470, 16'd25331, 16'd63658, 16'd9358, 16'd18374, 16'd7185, 16'd39286, 16'd18818, 16'd44268, 16'd35708, 16'd22331, 16'd36674});
	test_expansion(128'h6d6a1b4a397000dc714c1e9bb7595d50, {16'd439, 16'd12460, 16'd33266, 16'd174, 16'd45660, 16'd54303, 16'd29248, 16'd53037, 16'd35130, 16'd44208, 16'd45292, 16'd28142, 16'd57885, 16'd52979, 16'd53890, 16'd30970, 16'd9345, 16'd5451, 16'd9433, 16'd42390, 16'd62368, 16'd59156, 16'd23915, 16'd64046, 16'd10366, 16'd52560});
	test_expansion(128'h3209155e87fb87911ba822a9b80201ca, {16'd19306, 16'd7730, 16'd45366, 16'd34368, 16'd7573, 16'd6703, 16'd21394, 16'd1531, 16'd2677, 16'd1043, 16'd1780, 16'd52422, 16'd30395, 16'd51216, 16'd64663, 16'd52228, 16'd54529, 16'd41601, 16'd15445, 16'd1370, 16'd13169, 16'd14047, 16'd37068, 16'd48845, 16'd53789, 16'd57349});
	test_expansion(128'ha2b46f112fbeda83c2e51051bbf7f2a1, {16'd55140, 16'd22857, 16'd48913, 16'd30295, 16'd47720, 16'd36500, 16'd43788, 16'd61669, 16'd18089, 16'd6340, 16'd55656, 16'd49215, 16'd35356, 16'd50393, 16'd44242, 16'd18158, 16'd47091, 16'd15194, 16'd23672, 16'd5350, 16'd11019, 16'd48719, 16'd29356, 16'd22510, 16'd47635, 16'd15291});
	test_expansion(128'hb555ee949b9552a3d7a0a4a754a9a607, {16'd31291, 16'd1728, 16'd3938, 16'd2006, 16'd63613, 16'd39698, 16'd11440, 16'd36225, 16'd13753, 16'd13434, 16'd12256, 16'd199, 16'd63249, 16'd17437, 16'd63363, 16'd64167, 16'd36100, 16'd49429, 16'd58825, 16'd24289, 16'd7071, 16'd2221, 16'd10106, 16'd49100, 16'd24268, 16'd51424});
	test_expansion(128'ha3207eeffac345b68ce7ea5a0958e301, {16'd24546, 16'd16302, 16'd51267, 16'd1653, 16'd59234, 16'd6297, 16'd57513, 16'd31003, 16'd47788, 16'd59867, 16'd39924, 16'd35337, 16'd57103, 16'd24271, 16'd61064, 16'd51845, 16'd51982, 16'd50297, 16'd18896, 16'd64154, 16'd61054, 16'd39815, 16'd2645, 16'd51650, 16'd62198, 16'd4837});
	test_expansion(128'hb940a0a1cf38469bc96e9b4c2554d188, {16'd36644, 16'd42159, 16'd32492, 16'd32468, 16'd27775, 16'd1084, 16'd38702, 16'd7640, 16'd51778, 16'd15606, 16'd50313, 16'd53128, 16'd65171, 16'd31797, 16'd58047, 16'd22281, 16'd24516, 16'd10664, 16'd60888, 16'd9061, 16'd25977, 16'd20589, 16'd5860, 16'd54448, 16'd63048, 16'd46662});
	test_expansion(128'h6648631e86b7d6b14cbc0a34416236d3, {16'd48385, 16'd42389, 16'd63101, 16'd24682, 16'd56552, 16'd32488, 16'd41946, 16'd14322, 16'd38658, 16'd54648, 16'd35123, 16'd42599, 16'd51857, 16'd61534, 16'd8453, 16'd2388, 16'd64885, 16'd24475, 16'd32803, 16'd38828, 16'd44637, 16'd35809, 16'd50035, 16'd33299, 16'd44932, 16'd46430});
	test_expansion(128'hf8752ed2b59b1eeb25e1b424cc69e147, {16'd45656, 16'd6540, 16'd37448, 16'd54532, 16'd8600, 16'd53041, 16'd19423, 16'd2207, 16'd30951, 16'd58941, 16'd34365, 16'd62160, 16'd35911, 16'd62419, 16'd60555, 16'd14883, 16'd27213, 16'd9348, 16'd64686, 16'd58332, 16'd60930, 16'd59919, 16'd23674, 16'd17803, 16'd45865, 16'd10807});
	test_expansion(128'h2cec00beef04253f98be4c7823bbd794, {16'd12064, 16'd39772, 16'd40353, 16'd59195, 16'd62632, 16'd58289, 16'd49998, 16'd56130, 16'd62405, 16'd37808, 16'd19332, 16'd6596, 16'd24948, 16'd58836, 16'd44929, 16'd18925, 16'd16255, 16'd36676, 16'd15906, 16'd2551, 16'd59599, 16'd61047, 16'd46146, 16'd7928, 16'd58969, 16'd51027});
	test_expansion(128'h241f4cc39aeb4f290da8aeec1bde4670, {16'd871, 16'd23189, 16'd10209, 16'd24191, 16'd36548, 16'd32660, 16'd4420, 16'd39912, 16'd54994, 16'd51390, 16'd25678, 16'd32969, 16'd21178, 16'd50800, 16'd35047, 16'd55877, 16'd52260, 16'd2520, 16'd53594, 16'd40725, 16'd46209, 16'd26929, 16'd53736, 16'd10333, 16'd5416, 16'd24894});
	test_expansion(128'hba35f516b55298d0751383c2a95c11f6, {16'd50847, 16'd43725, 16'd58695, 16'd31818, 16'd4448, 16'd41132, 16'd20764, 16'd51634, 16'd44880, 16'd49725, 16'd16012, 16'd1709, 16'd7674, 16'd42014, 16'd23100, 16'd34646, 16'd31402, 16'd30846, 16'd60978, 16'd37681, 16'd15330, 16'd40832, 16'd9672, 16'd56913, 16'd41599, 16'd34711});
	test_expansion(128'h1dad1c3471255d7b7de05be140f69156, {16'd5682, 16'd24856, 16'd56981, 16'd49936, 16'd25465, 16'd14792, 16'd26907, 16'd46314, 16'd13110, 16'd29306, 16'd42713, 16'd19008, 16'd39896, 16'd12467, 16'd2206, 16'd37418, 16'd61277, 16'd54683, 16'd55383, 16'd54271, 16'd61853, 16'd21573, 16'd32419, 16'd14139, 16'd35749, 16'd35764});
	test_expansion(128'ha6db8151aa0dea00599405d5ea9c6be3, {16'd55019, 16'd8407, 16'd28124, 16'd6241, 16'd49152, 16'd58863, 16'd15280, 16'd34437, 16'd281, 16'd34995, 16'd47654, 16'd13316, 16'd35604, 16'd11089, 16'd29714, 16'd37715, 16'd41371, 16'd18722, 16'd61220, 16'd39004, 16'd22168, 16'd37154, 16'd11137, 16'd49430, 16'd14453, 16'd42016});
	test_expansion(128'hd5fe526a98dcbb6857f6d0f8390091c5, {16'd20236, 16'd28108, 16'd57613, 16'd52618, 16'd47079, 16'd36030, 16'd23675, 16'd5198, 16'd1380, 16'd18172, 16'd64545, 16'd51998, 16'd7782, 16'd27326, 16'd53887, 16'd13790, 16'd41506, 16'd39027, 16'd11693, 16'd39483, 16'd8750, 16'd57879, 16'd30405, 16'd32398, 16'd30491, 16'd42644});
	test_expansion(128'hd7f7de833dbf775696bee797b6ba5f2d, {16'd6536, 16'd40660, 16'd51132, 16'd22441, 16'd45597, 16'd27780, 16'd7229, 16'd33092, 16'd44755, 16'd41667, 16'd48329, 16'd13316, 16'd134, 16'd27543, 16'd21906, 16'd50404, 16'd36422, 16'd31953, 16'd51308, 16'd11306, 16'd36960, 16'd60017, 16'd54526, 16'd13489, 16'd11071, 16'd34825});
	test_expansion(128'hbae18c91bf46ea63be7054b93c32e3fc, {16'd42693, 16'd42046, 16'd32235, 16'd34623, 16'd50230, 16'd33144, 16'd42169, 16'd35169, 16'd2743, 16'd49949, 16'd2935, 16'd5765, 16'd32158, 16'd1466, 16'd18659, 16'd16223, 16'd30805, 16'd63882, 16'd25179, 16'd57208, 16'd36601, 16'd26476, 16'd26686, 16'd65088, 16'd30883, 16'd9682});
	test_expansion(128'hcaadc66c0ab9853c70936300c85ced53, {16'd12254, 16'd18871, 16'd55484, 16'd23657, 16'd28622, 16'd5968, 16'd51813, 16'd63696, 16'd19147, 16'd21182, 16'd60671, 16'd5324, 16'd35712, 16'd40371, 16'd36379, 16'd27821, 16'd7906, 16'd53602, 16'd36570, 16'd62365, 16'd23028, 16'd61186, 16'd9036, 16'd23720, 16'd22325, 16'd21});
	test_expansion(128'h22d1a3b4169e20a79876d933a4f9cc76, {16'd16453, 16'd23642, 16'd62444, 16'd39799, 16'd61554, 16'd56952, 16'd46581, 16'd39834, 16'd9138, 16'd56254, 16'd47545, 16'd17036, 16'd51450, 16'd52077, 16'd55652, 16'd25692, 16'd50856, 16'd33905, 16'd1550, 16'd880, 16'd21771, 16'd4799, 16'd41065, 16'd30340, 16'd62294, 16'd59451});
	test_expansion(128'h852acb772d28121eae41e8b5dd18b25b, {16'd9701, 16'd19961, 16'd47954, 16'd34993, 16'd49762, 16'd1208, 16'd56846, 16'd8225, 16'd34993, 16'd41897, 16'd38432, 16'd44413, 16'd9910, 16'd30969, 16'd21698, 16'd52426, 16'd13666, 16'd22103, 16'd41130, 16'd17665, 16'd28721, 16'd61327, 16'd43591, 16'd25877, 16'd48986, 16'd47553});
	test_expansion(128'h54db1358a36a6812ff8b4c4d4da57329, {16'd32961, 16'd18092, 16'd23445, 16'd37516, 16'd36978, 16'd35827, 16'd5281, 16'd14309, 16'd55461, 16'd29001, 16'd35950, 16'd49632, 16'd3474, 16'd43974, 16'd30937, 16'd16855, 16'd51798, 16'd54111, 16'd17366, 16'd23316, 16'd25319, 16'd42740, 16'd48358, 16'd47446, 16'd26967, 16'd17223});
	test_expansion(128'h22160d9265bcd30fdeaf90858678da38, {16'd51534, 16'd29979, 16'd29724, 16'd39614, 16'd11417, 16'd12326, 16'd15509, 16'd16179, 16'd4064, 16'd3911, 16'd11670, 16'd28082, 16'd28707, 16'd292, 16'd41034, 16'd6581, 16'd45809, 16'd578, 16'd23953, 16'd63932, 16'd24611, 16'd38029, 16'd45008, 16'd48070, 16'd7595, 16'd4519});
	test_expansion(128'hbf922589ad410fb414a39a8be880ae3c, {16'd199, 16'd5878, 16'd17313, 16'd7238, 16'd36217, 16'd3418, 16'd3586, 16'd2673, 16'd32066, 16'd30878, 16'd32319, 16'd42396, 16'd18044, 16'd33280, 16'd43286, 16'd64969, 16'd57890, 16'd41855, 16'd15808, 16'd16621, 16'd34657, 16'd32661, 16'd29290, 16'd13434, 16'd30861, 16'd23219});
	test_expansion(128'h5ca1c63d426d0b63099d70b3784ed135, {16'd40668, 16'd7809, 16'd54372, 16'd65073, 16'd39176, 16'd56109, 16'd7118, 16'd43422, 16'd6786, 16'd22475, 16'd64266, 16'd63177, 16'd54161, 16'd55625, 16'd25853, 16'd14578, 16'd53595, 16'd46496, 16'd26738, 16'd15664, 16'd43417, 16'd27405, 16'd42238, 16'd22672, 16'd57733, 16'd23579});
	test_expansion(128'h9debff2f03671bb1385d3f07423b3b6f, {16'd51588, 16'd13917, 16'd63055, 16'd52548, 16'd1179, 16'd49132, 16'd44129, 16'd16939, 16'd38778, 16'd34220, 16'd25860, 16'd47981, 16'd29577, 16'd13076, 16'd41180, 16'd45914, 16'd38708, 16'd38704, 16'd30733, 16'd58676, 16'd57841, 16'd48361, 16'd23522, 16'd32787, 16'd9103, 16'd34181});
	test_expansion(128'hfe4bab4b8300162ed54b7f59d2f4c92c, {16'd20968, 16'd42015, 16'd31938, 16'd3061, 16'd13619, 16'd61534, 16'd17698, 16'd30205, 16'd4939, 16'd16554, 16'd59820, 16'd31046, 16'd17641, 16'd18857, 16'd296, 16'd37668, 16'd19847, 16'd24093, 16'd44353, 16'd1006, 16'd61527, 16'd38501, 16'd11589, 16'd10341, 16'd16874, 16'd18623});
	test_expansion(128'h60849f7dc8f2d2c0fd7636a19ee94909, {16'd20663, 16'd26831, 16'd9610, 16'd22462, 16'd13601, 16'd43385, 16'd24611, 16'd55031, 16'd42529, 16'd9840, 16'd26144, 16'd46168, 16'd24226, 16'd51080, 16'd1976, 16'd35635, 16'd53949, 16'd62226, 16'd4076, 16'd21175, 16'd24282, 16'd3048, 16'd9805, 16'd1725, 16'd53265, 16'd7576});
	test_expansion(128'h8c23eaccea6e0abe1136557d2dbb4fcc, {16'd47579, 16'd33869, 16'd10071, 16'd39373, 16'd13055, 16'd10731, 16'd47662, 16'd63354, 16'd8017, 16'd33814, 16'd61662, 16'd42626, 16'd25589, 16'd28621, 16'd53463, 16'd49554, 16'd42042, 16'd2626, 16'd61055, 16'd4843, 16'd37320, 16'd16268, 16'd41082, 16'd2056, 16'd26783, 16'd16242});
	test_expansion(128'hbe107efef73fa03e07d906419d132fd4, {16'd22134, 16'd8471, 16'd4212, 16'd52136, 16'd53568, 16'd30505, 16'd30569, 16'd30289, 16'd29433, 16'd46174, 16'd10656, 16'd1235, 16'd48369, 16'd26645, 16'd42944, 16'd18982, 16'd63747, 16'd48295, 16'd60599, 16'd12156, 16'd43184, 16'd62720, 16'd6592, 16'd38006, 16'd35726, 16'd37689});
	test_expansion(128'h8d751493324b37e6e6aaa6ec10fc5f87, {16'd29748, 16'd29380, 16'd60936, 16'd37614, 16'd60276, 16'd36373, 16'd5845, 16'd30656, 16'd45768, 16'd57735, 16'd27560, 16'd9353, 16'd21360, 16'd20349, 16'd29511, 16'd64343, 16'd60752, 16'd8607, 16'd17365, 16'd25357, 16'd36658, 16'd32956, 16'd28988, 16'd37806, 16'd44073, 16'd11516});
	test_expansion(128'h2294efcb6761c2c5d24916b44ce0d92b, {16'd25683, 16'd43380, 16'd32970, 16'd25750, 16'd58287, 16'd46452, 16'd64011, 16'd42739, 16'd19719, 16'd25908, 16'd9119, 16'd23275, 16'd23580, 16'd33348, 16'd1214, 16'd9049, 16'd46756, 16'd52115, 16'd62023, 16'd27732, 16'd61039, 16'd34101, 16'd47608, 16'd17123, 16'd6560, 16'd20772});
	test_expansion(128'h3953504cb3d24b6b7c7d2dfdae7ef913, {16'd55267, 16'd19292, 16'd63020, 16'd39398, 16'd14274, 16'd63543, 16'd9780, 16'd36257, 16'd44713, 16'd48884, 16'd38957, 16'd23487, 16'd12372, 16'd14459, 16'd42194, 16'd8353, 16'd57815, 16'd11404, 16'd22879, 16'd47614, 16'd35976, 16'd31562, 16'd38837, 16'd62455, 16'd44042, 16'd45697});
	test_expansion(128'h089e3420f03096986f7615416e119405, {16'd1650, 16'd25266, 16'd9089, 16'd62593, 16'd28227, 16'd20687, 16'd47747, 16'd29948, 16'd8823, 16'd59416, 16'd61830, 16'd53291, 16'd60042, 16'd55209, 16'd45603, 16'd34943, 16'd62436, 16'd20944, 16'd64451, 16'd33151, 16'd59708, 16'd64579, 16'd36994, 16'd28089, 16'd44992, 16'd14788});
	test_expansion(128'h94be024278e01e6e07bcfb8f46a73d6c, {16'd19861, 16'd14374, 16'd14878, 16'd34544, 16'd14021, 16'd50169, 16'd24004, 16'd29781, 16'd62006, 16'd19646, 16'd1293, 16'd17266, 16'd1589, 16'd47896, 16'd21777, 16'd59082, 16'd20867, 16'd51164, 16'd48737, 16'd31797, 16'd45071, 16'd56716, 16'd27763, 16'd60052, 16'd4084, 16'd15481});
	test_expansion(128'h4f40f0675a8251c7f0a156d584f4bfa9, {16'd48380, 16'd29726, 16'd62131, 16'd8649, 16'd3931, 16'd1785, 16'd7553, 16'd15776, 16'd29477, 16'd34213, 16'd31280, 16'd53978, 16'd57856, 16'd43890, 16'd39965, 16'd34020, 16'd37165, 16'd14378, 16'd4254, 16'd26164, 16'd15327, 16'd2041, 16'd1086, 16'd62080, 16'd1221, 16'd65125});
	test_expansion(128'h59a564e52d9f13638811abec649bfc23, {16'd3794, 16'd31325, 16'd52641, 16'd4239, 16'd30034, 16'd16630, 16'd11258, 16'd37350, 16'd36438, 16'd64781, 16'd17173, 16'd44030, 16'd31959, 16'd57122, 16'd55492, 16'd4032, 16'd19577, 16'd51172, 16'd45714, 16'd6913, 16'd8730, 16'd34728, 16'd3641, 16'd16730, 16'd36470, 16'd48389});
	test_expansion(128'h7aa81910398716c09b63029460cfa846, {16'd2609, 16'd23235, 16'd1700, 16'd29631, 16'd15068, 16'd49469, 16'd34809, 16'd41561, 16'd47692, 16'd58130, 16'd4646, 16'd20349, 16'd12223, 16'd18474, 16'd11715, 16'd28453, 16'd13326, 16'd28012, 16'd20900, 16'd18064, 16'd25993, 16'd62277, 16'd17085, 16'd26294, 16'd40537, 16'd14648});
	test_expansion(128'h37b391dbdfc555d33fab72c69b83d828, {16'd27660, 16'd16173, 16'd51234, 16'd37616, 16'd46229, 16'd12421, 16'd22672, 16'd51042, 16'd15695, 16'd19291, 16'd31839, 16'd30016, 16'd39026, 16'd49141, 16'd28876, 16'd11609, 16'd50381, 16'd57841, 16'd52272, 16'd52843, 16'd18886, 16'd50737, 16'd41283, 16'd56945, 16'd2852, 16'd59751});
	test_expansion(128'h5cfec92daf2a4f66e67d7606d80bc821, {16'd1201, 16'd11935, 16'd39229, 16'd20918, 16'd47389, 16'd41473, 16'd42670, 16'd23441, 16'd50508, 16'd28413, 16'd54673, 16'd23161, 16'd49683, 16'd49901, 16'd42186, 16'd8319, 16'd26050, 16'd59451, 16'd46839, 16'd38718, 16'd53532, 16'd14722, 16'd15562, 16'd22207, 16'd54633, 16'd55022});
	test_expansion(128'h9aaaf3fab3c73e8e74813fab212f29c2, {16'd60333, 16'd19967, 16'd32448, 16'd6794, 16'd5157, 16'd62385, 16'd14404, 16'd51626, 16'd36090, 16'd29564, 16'd6767, 16'd40422, 16'd16691, 16'd42105, 16'd56754, 16'd4634, 16'd54841, 16'd27376, 16'd17160, 16'd56601, 16'd18802, 16'd20592, 16'd29887, 16'd59309, 16'd18505, 16'd54822});
	test_expansion(128'h8529bcc6994de801758bb6e1b36ee81d, {16'd3167, 16'd23794, 16'd13917, 16'd65097, 16'd59407, 16'd25607, 16'd28802, 16'd41492, 16'd62450, 16'd5172, 16'd44048, 16'd45789, 16'd54791, 16'd34394, 16'd40162, 16'd63461, 16'd33526, 16'd62377, 16'd2871, 16'd61034, 16'd11958, 16'd16119, 16'd14048, 16'd4388, 16'd34360, 16'd34707});
	test_expansion(128'h69a58143f34600c97f7001e06dc5ebd6, {16'd26943, 16'd27461, 16'd47791, 16'd62963, 16'd13669, 16'd24806, 16'd51548, 16'd10870, 16'd799, 16'd20690, 16'd46421, 16'd25866, 16'd30866, 16'd39178, 16'd47131, 16'd59652, 16'd63228, 16'd30863, 16'd65275, 16'd23040, 16'd6116, 16'd6134, 16'd49806, 16'd8043, 16'd7249, 16'd31210});
	test_expansion(128'h5d66f8590f52e39208a64673848ff1e8, {16'd47259, 16'd51829, 16'd63379, 16'd10484, 16'd39999, 16'd11119, 16'd61702, 16'd39455, 16'd31861, 16'd28349, 16'd20408, 16'd13875, 16'd13991, 16'd17315, 16'd3021, 16'd26417, 16'd1176, 16'd43968, 16'd25896, 16'd34115, 16'd60107, 16'd43756, 16'd40441, 16'd13622, 16'd42548, 16'd65320});
	test_expansion(128'h3cab79eaa3f2b77dcfcf8af57bf8ab59, {16'd50547, 16'd32868, 16'd53449, 16'd58440, 16'd58514, 16'd37861, 16'd63471, 16'd41451, 16'd31422, 16'd57477, 16'd37241, 16'd17258, 16'd9211, 16'd43320, 16'd62206, 16'd18854, 16'd22490, 16'd32325, 16'd14735, 16'd18212, 16'd7674, 16'd21217, 16'd2427, 16'd456, 16'd60798, 16'd28527});
	test_expansion(128'h61f98d953b9536c160823d8164516364, {16'd4763, 16'd47923, 16'd50979, 16'd23067, 16'd27214, 16'd56324, 16'd1596, 16'd43341, 16'd39886, 16'd47405, 16'd16139, 16'd43328, 16'd64737, 16'd32131, 16'd7255, 16'd10656, 16'd54128, 16'd11990, 16'd15402, 16'd64570, 16'd35927, 16'd23711, 16'd5910, 16'd14954, 16'd38358, 16'd2586});
	test_expansion(128'h3a7ddd6f2f2624ab8fd15236edc74c1d, {16'd41475, 16'd36273, 16'd23896, 16'd22349, 16'd45117, 16'd34666, 16'd53685, 16'd1791, 16'd47033, 16'd63702, 16'd27608, 16'd18473, 16'd39904, 16'd17229, 16'd26723, 16'd9622, 16'd25065, 16'd13639, 16'd17982, 16'd47178, 16'd50096, 16'd4113, 16'd31945, 16'd36014, 16'd40921, 16'd48266});
	test_expansion(128'haee3bf70f460826666502d71a5b2d906, {16'd54960, 16'd29398, 16'd31936, 16'd19879, 16'd35278, 16'd8153, 16'd64005, 16'd54785, 16'd13930, 16'd26756, 16'd6935, 16'd21157, 16'd28702, 16'd27735, 16'd8659, 16'd21428, 16'd50397, 16'd32836, 16'd31335, 16'd23409, 16'd60847, 16'd28689, 16'd56427, 16'd19464, 16'd33563, 16'd26265});
	test_expansion(128'h3082e17f61c82f36f0a312c6458ebe82, {16'd6202, 16'd21083, 16'd34303, 16'd45518, 16'd62613, 16'd16885, 16'd52116, 16'd8234, 16'd23781, 16'd40142, 16'd58228, 16'd12314, 16'd20929, 16'd54534, 16'd1886, 16'd516, 16'd35724, 16'd63876, 16'd19936, 16'd63461, 16'd582, 16'd1010, 16'd44533, 16'd9515, 16'd37792, 16'd16278});
	test_expansion(128'h8dea4106ccfd421a2646b629400bd89e, {16'd38033, 16'd42079, 16'd544, 16'd34169, 16'd3983, 16'd50369, 16'd32065, 16'd47231, 16'd12127, 16'd2196, 16'd50972, 16'd52848, 16'd65096, 16'd7779, 16'd12344, 16'd25943, 16'd52372, 16'd8669, 16'd57820, 16'd62214, 16'd2067, 16'd51974, 16'd47431, 16'd23576, 16'd30626, 16'd28613});
	test_expansion(128'h0ff32770bbfe821209c329b21b6fa1e8, {16'd56894, 16'd2809, 16'd46947, 16'd53680, 16'd63186, 16'd37127, 16'd28518, 16'd18712, 16'd12514, 16'd20263, 16'd21447, 16'd26825, 16'd62262, 16'd2647, 16'd5262, 16'd6505, 16'd43326, 16'd47299, 16'd3662, 16'd42592, 16'd28519, 16'd43122, 16'd12610, 16'd45024, 16'd12091, 16'd23073});
	test_expansion(128'h627f1a5fde3b7762250668c4076cbba1, {16'd7776, 16'd54716, 16'd1720, 16'd28052, 16'd7297, 16'd28539, 16'd34630, 16'd26648, 16'd51195, 16'd30450, 16'd22701, 16'd17316, 16'd45887, 16'd49150, 16'd31490, 16'd47560, 16'd15948, 16'd62196, 16'd10429, 16'd43422, 16'd32907, 16'd65208, 16'd31343, 16'd1186, 16'd11783, 16'd45918});
	test_expansion(128'hb9f62fb33598465844575ee8968e59de, {16'd21046, 16'd55444, 16'd27165, 16'd24097, 16'd33256, 16'd14970, 16'd6360, 16'd21105, 16'd27911, 16'd30720, 16'd8194, 16'd26915, 16'd48551, 16'd34503, 16'd5328, 16'd45017, 16'd13136, 16'd1461, 16'd33784, 16'd16772, 16'd47428, 16'd6342, 16'd53658, 16'd18066, 16'd48304, 16'd8811});
	test_expansion(128'h75e5b8909a5956e43c89529b08074b34, {16'd35153, 16'd11992, 16'd63675, 16'd10488, 16'd56700, 16'd5883, 16'd17971, 16'd45966, 16'd18485, 16'd45014, 16'd28662, 16'd29570, 16'd48033, 16'd30922, 16'd59505, 16'd46381, 16'd56307, 16'd8978, 16'd63791, 16'd13530, 16'd21840, 16'd48843, 16'd26351, 16'd18947, 16'd52884, 16'd64623});
	test_expansion(128'hd7301c41899f6ab794bb62da5609fe88, {16'd30053, 16'd24408, 16'd54487, 16'd64933, 16'd14519, 16'd6664, 16'd48590, 16'd17243, 16'd64483, 16'd42879, 16'd50999, 16'd15306, 16'd22390, 16'd8335, 16'd59873, 16'd16439, 16'd44455, 16'd13858, 16'd6667, 16'd413, 16'd29569, 16'd2534, 16'd11214, 16'd39097, 16'd60509, 16'd48594});
	test_expansion(128'h7c97ed26d394a368370ed21a98479418, {16'd21792, 16'd24876, 16'd31765, 16'd35994, 16'd25163, 16'd17835, 16'd38034, 16'd38673, 16'd32148, 16'd61765, 16'd39984, 16'd31526, 16'd354, 16'd53805, 16'd17730, 16'd6267, 16'd63699, 16'd65400, 16'd61255, 16'd52507, 16'd8809, 16'd61988, 16'd19390, 16'd8244, 16'd31386, 16'd18760});
	test_expansion(128'h8b1744c5a5a9b91d6fa189a6d2c519db, {16'd34029, 16'd39777, 16'd63518, 16'd8848, 16'd60434, 16'd29435, 16'd40547, 16'd54513, 16'd17683, 16'd55095, 16'd579, 16'd47326, 16'd11801, 16'd23507, 16'd18097, 16'd43873, 16'd38779, 16'd57767, 16'd21842, 16'd28499, 16'd57369, 16'd32083, 16'd45996, 16'd18642, 16'd32470, 16'd63985});
	test_expansion(128'h044783cdaaee018e537903d9a08432cd, {16'd22277, 16'd15700, 16'd55643, 16'd1218, 16'd16602, 16'd43449, 16'd17664, 16'd51628, 16'd47878, 16'd33578, 16'd3210, 16'd39312, 16'd39295, 16'd17834, 16'd38541, 16'd57967, 16'd49873, 16'd62649, 16'd35391, 16'd63792, 16'd11631, 16'd15813, 16'd44557, 16'd18533, 16'd65106, 16'd40622});
	test_expansion(128'h08c3d1b2c6627c82fa73f382519584e4, {16'd185, 16'd48557, 16'd13609, 16'd13306, 16'd2725, 16'd14226, 16'd54168, 16'd27611, 16'd40078, 16'd21745, 16'd63131, 16'd15913, 16'd4035, 16'd22212, 16'd21596, 16'd40191, 16'd10971, 16'd50648, 16'd40974, 16'd60384, 16'd34539, 16'd40909, 16'd30856, 16'd58263, 16'd18409, 16'd57492});
	test_expansion(128'h2dc56e3501c6103a9ba811fd08c2c198, {16'd16468, 16'd62225, 16'd36120, 16'd40828, 16'd48242, 16'd61887, 16'd51618, 16'd4388, 16'd20023, 16'd15328, 16'd38233, 16'd25717, 16'd15197, 16'd4939, 16'd56893, 16'd17562, 16'd63842, 16'd61124, 16'd47334, 16'd44596, 16'd34402, 16'd28974, 16'd36015, 16'd53978, 16'd23087, 16'd25521});
	test_expansion(128'h1e94f95f3f7ce0cd2d10af6590baec81, {16'd12347, 16'd54052, 16'd55585, 16'd47361, 16'd49544, 16'd44957, 16'd45168, 16'd58807, 16'd46991, 16'd26701, 16'd4963, 16'd62355, 16'd4496, 16'd59330, 16'd10774, 16'd48092, 16'd29223, 16'd28628, 16'd45027, 16'd45139, 16'd23927, 16'd57515, 16'd51344, 16'd22824, 16'd65407, 16'd7015});
	test_expansion(128'hc0c6d8bf0d16998902e824e130f7b3f3, {16'd47325, 16'd46720, 16'd24448, 16'd21519, 16'd3001, 16'd25263, 16'd29972, 16'd18772, 16'd52163, 16'd72, 16'd57347, 16'd6263, 16'd63987, 16'd61533, 16'd36664, 16'd37233, 16'd4937, 16'd17689, 16'd9579, 16'd12070, 16'd41586, 16'd9515, 16'd42997, 16'd982, 16'd44659, 16'd56071});
	test_expansion(128'hcc260b3de92f6cd199b8a81766e7a0d2, {16'd45376, 16'd16279, 16'd19631, 16'd57708, 16'd51153, 16'd9836, 16'd15551, 16'd54123, 16'd55550, 16'd19135, 16'd55410, 16'd42970, 16'd64029, 16'd17933, 16'd2539, 16'd21757, 16'd15840, 16'd57542, 16'd18582, 16'd22219, 16'd43327, 16'd60374, 16'd20238, 16'd35636, 16'd32886, 16'd55822});
	test_expansion(128'h240f7f371db0a11e67a91c85f3b2b706, {16'd34652, 16'd3988, 16'd17933, 16'd28553, 16'd20612, 16'd63136, 16'd7571, 16'd27889, 16'd14137, 16'd64391, 16'd7580, 16'd52992, 16'd64874, 16'd7560, 16'd40483, 16'd52707, 16'd53769, 16'd35979, 16'd28276, 16'd41089, 16'd14530, 16'd23879, 16'd56764, 16'd58321, 16'd19215, 16'd46368});
	test_expansion(128'h21534483aae067d68bab48da037e9cf3, {16'd24282, 16'd58482, 16'd16846, 16'd58461, 16'd7221, 16'd58033, 16'd56569, 16'd61200, 16'd30447, 16'd27775, 16'd54635, 16'd14498, 16'd12808, 16'd23528, 16'd46774, 16'd24401, 16'd48438, 16'd27058, 16'd39309, 16'd33338, 16'd11600, 16'd43775, 16'd40163, 16'd10372, 16'd7857, 16'd12032});
	test_expansion(128'h575830e7ec76421032457a160a7faa18, {16'd29744, 16'd18031, 16'd7016, 16'd48721, 16'd44942, 16'd50134, 16'd11600, 16'd38228, 16'd36324, 16'd6159, 16'd7262, 16'd32826, 16'd42584, 16'd57879, 16'd45, 16'd20137, 16'd57112, 16'd4146, 16'd16304, 16'd45388, 16'd24183, 16'd38717, 16'd56100, 16'd40173, 16'd15303, 16'd29897});
	test_expansion(128'he44ac8d76434272c8fc71caceb920e9c, {16'd16051, 16'd36575, 16'd38744, 16'd61823, 16'd6605, 16'd7627, 16'd44473, 16'd44846, 16'd29766, 16'd13838, 16'd63478, 16'd30806, 16'd45067, 16'd3691, 16'd49345, 16'd36602, 16'd13666, 16'd62283, 16'd61721, 16'd63591, 16'd56293, 16'd55460, 16'd8669, 16'd15615, 16'd14627, 16'd32967});
	test_expansion(128'h420389542905fcaf4334e7464157e968, {16'd27668, 16'd7620, 16'd14198, 16'd48571, 16'd28294, 16'd26585, 16'd51735, 16'd50576, 16'd1772, 16'd44303, 16'd38568, 16'd1335, 16'd15268, 16'd4464, 16'd1388, 16'd32360, 16'd53333, 16'd6075, 16'd52884, 16'd9690, 16'd29347, 16'd44843, 16'd4867, 16'd32675, 16'd15296, 16'd20542});
	test_expansion(128'h3db312e37d31cb667df92104e7a1d3d4, {16'd20599, 16'd11403, 16'd32519, 16'd25782, 16'd8168, 16'd52843, 16'd57300, 16'd24963, 16'd25011, 16'd59200, 16'd733, 16'd64095, 16'd10702, 16'd42932, 16'd63810, 16'd29404, 16'd37905, 16'd4341, 16'd12838, 16'd20702, 16'd36393, 16'd1643, 16'd51336, 16'd40995, 16'd48135, 16'd30766});
	test_expansion(128'hed59c26a27c65d1a199abd97c860e9f0, {16'd17377, 16'd50828, 16'd63913, 16'd58778, 16'd30388, 16'd10966, 16'd3458, 16'd10705, 16'd21198, 16'd5519, 16'd40412, 16'd43561, 16'd23659, 16'd38444, 16'd6653, 16'd13458, 16'd31864, 16'd23588, 16'd12940, 16'd1932, 16'd794, 16'd56956, 16'd63331, 16'd10304, 16'd33121, 16'd23611});
	test_expansion(128'h01c7c87c85dc53b99e0b582ce824d525, {16'd47584, 16'd41769, 16'd29323, 16'd58079, 16'd58971, 16'd54526, 16'd49514, 16'd20078, 16'd38608, 16'd19607, 16'd24318, 16'd42123, 16'd17464, 16'd36145, 16'd2885, 16'd21773, 16'd56839, 16'd45363, 16'd9567, 16'd24336, 16'd53546, 16'd37280, 16'd65261, 16'd7259, 16'd40702, 16'd59353});
	test_expansion(128'ha99fd8f90cbb05c44111b7c0784e0052, {16'd39376, 16'd50810, 16'd55938, 16'd45434, 16'd54116, 16'd64198, 16'd60197, 16'd17093, 16'd47704, 16'd10533, 16'd27572, 16'd53968, 16'd10561, 16'd63914, 16'd41058, 16'd39612, 16'd23908, 16'd55312, 16'd51251, 16'd8621, 16'd21578, 16'd29734, 16'd29078, 16'd16701, 16'd48097, 16'd2772});
	test_expansion(128'h84763592fb275e606c9a90375d8cf781, {16'd42912, 16'd61328, 16'd64319, 16'd22578, 16'd50994, 16'd12063, 16'd19938, 16'd49911, 16'd39126, 16'd45104, 16'd61408, 16'd37257, 16'd51838, 16'd9772, 16'd24982, 16'd47047, 16'd60291, 16'd52599, 16'd21444, 16'd16098, 16'd41040, 16'd60292, 16'd4977, 16'd10945, 16'd40157, 16'd21357});
	test_expansion(128'he8756de13b713078bb486d0ba049a02c, {16'd2642, 16'd49155, 16'd54573, 16'd36147, 16'd12916, 16'd64013, 16'd15930, 16'd6647, 16'd5703, 16'd18017, 16'd23698, 16'd6064, 16'd29800, 16'd2375, 16'd25819, 16'd33881, 16'd62434, 16'd65434, 16'd24092, 16'd17709, 16'd48264, 16'd52125, 16'd64771, 16'd25133, 16'd52199, 16'd48984});
	test_expansion(128'h197d22e09676a712a3e8362d1e97041c, {16'd60592, 16'd42532, 16'd20371, 16'd8305, 16'd648, 16'd18860, 16'd4563, 16'd14111, 16'd62686, 16'd40436, 16'd17827, 16'd24164, 16'd48384, 16'd13252, 16'd5392, 16'd20126, 16'd58063, 16'd7921, 16'd24795, 16'd3027, 16'd2193, 16'd58498, 16'd22003, 16'd45096, 16'd61751, 16'd54157});
	test_expansion(128'h19b11075bea435fca61bed7ebc3e988d, {16'd63307, 16'd44423, 16'd54323, 16'd5657, 16'd53471, 16'd29657, 16'd54719, 16'd49063, 16'd60965, 16'd61542, 16'd29419, 16'd54500, 16'd42149, 16'd36909, 16'd12242, 16'd60406, 16'd8059, 16'd18229, 16'd16249, 16'd63222, 16'd43476, 16'd13054, 16'd15133, 16'd6488, 16'd61222, 16'd14036});
	test_expansion(128'he8196ed08317f49a01d9bb4805df52d3, {16'd33772, 16'd48530, 16'd51783, 16'd17803, 16'd18613, 16'd46662, 16'd16854, 16'd25693, 16'd14228, 16'd15717, 16'd23610, 16'd25806, 16'd26907, 16'd50904, 16'd2009, 16'd63874, 16'd33113, 16'd47066, 16'd26737, 16'd40041, 16'd53075, 16'd37169, 16'd14130, 16'd8639, 16'd1559, 16'd45484});
	test_expansion(128'hdf879cf8f8256f817fb97d7db8d5338f, {16'd12880, 16'd2037, 16'd62632, 16'd17028, 16'd39424, 16'd15768, 16'd32182, 16'd51796, 16'd34993, 16'd15628, 16'd60054, 16'd25176, 16'd42347, 16'd20210, 16'd18652, 16'd58030, 16'd47791, 16'd104, 16'd47063, 16'd34233, 16'd55913, 16'd55201, 16'd16000, 16'd48814, 16'd23585, 16'd47942});
	test_expansion(128'h88ab065f6a8e47d355a9768dc6c35198, {16'd54881, 16'd3366, 16'd9969, 16'd46387, 16'd9737, 16'd43356, 16'd17517, 16'd36094, 16'd4229, 16'd60513, 16'd62845, 16'd32301, 16'd21907, 16'd6976, 16'd19394, 16'd2262, 16'd51359, 16'd34048, 16'd57664, 16'd7977, 16'd52983, 16'd4876, 16'd714, 16'd53712, 16'd12442, 16'd25555});
	test_expansion(128'h122f280aeb391a316cb0d98d551d0bab, {16'd14461, 16'd5210, 16'd11420, 16'd1923, 16'd47065, 16'd39904, 16'd17234, 16'd18387, 16'd4029, 16'd28556, 16'd12491, 16'd33929, 16'd54170, 16'd54237, 16'd49206, 16'd32290, 16'd6194, 16'd24069, 16'd38080, 16'd5066, 16'd32142, 16'd61640, 16'd6797, 16'd45622, 16'd2171, 16'd27006});
	test_expansion(128'h65ad73064085ea0629c111b585f6e46a, {16'd33812, 16'd57381, 16'd15247, 16'd64729, 16'd7043, 16'd25224, 16'd21950, 16'd17441, 16'd34511, 16'd41975, 16'd52850, 16'd29725, 16'd64602, 16'd25868, 16'd52368, 16'd4222, 16'd42206, 16'd43057, 16'd65313, 16'd19162, 16'd21360, 16'd1143, 16'd2999, 16'd24110, 16'd56311, 16'd46135});
	test_expansion(128'h468b57230e7468ed68ea10fa873955f7, {16'd59231, 16'd6591, 16'd13386, 16'd35024, 16'd23249, 16'd56277, 16'd27834, 16'd42961, 16'd23778, 16'd60817, 16'd31471, 16'd39684, 16'd9528, 16'd33504, 16'd17696, 16'd53430, 16'd63185, 16'd56193, 16'd52685, 16'd10919, 16'd18583, 16'd4169, 16'd3178, 16'd12802, 16'd25501, 16'd35454});
	test_expansion(128'hdc483ec6e41826c0951396ecc496fcd6, {16'd26170, 16'd31577, 16'd12748, 16'd48154, 16'd17945, 16'd20449, 16'd57665, 16'd31224, 16'd23107, 16'd58575, 16'd12077, 16'd64026, 16'd63307, 16'd3299, 16'd60172, 16'd51606, 16'd17867, 16'd5720, 16'd27614, 16'd1359, 16'd3044, 16'd19611, 16'd52373, 16'd39015, 16'd13846, 16'd49561});
	test_expansion(128'hfcc5bcf9b4c5ce05f954cbd7f9139c2b, {16'd27960, 16'd5299, 16'd53224, 16'd41104, 16'd9000, 16'd5786, 16'd65490, 16'd54953, 16'd48784, 16'd49351, 16'd39645, 16'd51430, 16'd35993, 16'd13571, 16'd23121, 16'd53872, 16'd46461, 16'd45082, 16'd19062, 16'd45163, 16'd21265, 16'd59003, 16'd32642, 16'd36170, 16'd27421, 16'd55838});
	test_expansion(128'h97621cf24eed7451d50c24832f08e775, {16'd26768, 16'd34038, 16'd23912, 16'd29163, 16'd57309, 16'd31323, 16'd8406, 16'd9977, 16'd15412, 16'd41591, 16'd59176, 16'd32739, 16'd26769, 16'd52100, 16'd57748, 16'd47869, 16'd35959, 16'd32170, 16'd9642, 16'd32022, 16'd7970, 16'd32924, 16'd45063, 16'd32199, 16'd38265, 16'd21341});
	test_expansion(128'hd549617a9281054e498371f1a01a0d79, {16'd62721, 16'd21569, 16'd33555, 16'd2407, 16'd17767, 16'd62589, 16'd5983, 16'd23815, 16'd61227, 16'd27152, 16'd23574, 16'd11493, 16'd22189, 16'd23556, 16'd15555, 16'd56793, 16'd6153, 16'd32533, 16'd48499, 16'd51914, 16'd51367, 16'd15019, 16'd9959, 16'd22495, 16'd45056, 16'd7033});
	test_expansion(128'h1ff9fce38cdf132c15b503d0311ad8dd, {16'd16302, 16'd1587, 16'd21664, 16'd28479, 16'd19819, 16'd55603, 16'd21585, 16'd19510, 16'd28126, 16'd16722, 16'd40035, 16'd52501, 16'd43260, 16'd41576, 16'd44855, 16'd20600, 16'd30158, 16'd8026, 16'd32486, 16'd55856, 16'd54450, 16'd47560, 16'd16561, 16'd27067, 16'd38268, 16'd24172});
	test_expansion(128'h4ddf5c8748de95ab4ec918acb03cba97, {16'd60522, 16'd9440, 16'd37918, 16'd32308, 16'd54117, 16'd9028, 16'd12810, 16'd13462, 16'd5154, 16'd7969, 16'd7715, 16'd9017, 16'd10142, 16'd10424, 16'd29806, 16'd7444, 16'd40400, 16'd47757, 16'd61563, 16'd16275, 16'd62673, 16'd30777, 16'd63421, 16'd61710, 16'd15763, 16'd25230});
	test_expansion(128'h678c0767f6a6ff39233706adf30b67d6, {16'd28283, 16'd53126, 16'd27529, 16'd38505, 16'd32210, 16'd14366, 16'd48546, 16'd46323, 16'd36259, 16'd16584, 16'd13986, 16'd45453, 16'd38148, 16'd29070, 16'd1372, 16'd45409, 16'd42590, 16'd25559, 16'd56229, 16'd1436, 16'd59716, 16'd63451, 16'd28238, 16'd12394, 16'd52273, 16'd20912});
	test_expansion(128'h476188190b0d3bfeb4b474e69561d289, {16'd39647, 16'd7694, 16'd3650, 16'd47973, 16'd28447, 16'd30022, 16'd19641, 16'd51480, 16'd26024, 16'd978, 16'd48404, 16'd476, 16'd54392, 16'd51790, 16'd44290, 16'd7010, 16'd32631, 16'd1810, 16'd46953, 16'd30808, 16'd39331, 16'd14702, 16'd13086, 16'd36624, 16'd14184, 16'd19273});
	test_expansion(128'hbaf3aa988621e9f1e50a3df1fb337b2a, {16'd41969, 16'd34296, 16'd27757, 16'd47266, 16'd98, 16'd63455, 16'd712, 16'd47876, 16'd54344, 16'd18165, 16'd7573, 16'd706, 16'd57326, 16'd2988, 16'd61597, 16'd11401, 16'd27579, 16'd15578, 16'd28327, 16'd5220, 16'd14447, 16'd25788, 16'd25479, 16'd7687, 16'd64305, 16'd25506});
	test_expansion(128'h9b6df4dba754ff2bb38e6e673919cce3, {16'd10644, 16'd21781, 16'd21260, 16'd60748, 16'd48471, 16'd28063, 16'd57343, 16'd50576, 16'd15430, 16'd2741, 16'd39850, 16'd11663, 16'd1667, 16'd32606, 16'd36338, 16'd31916, 16'd2729, 16'd168, 16'd8146, 16'd4490, 16'd19052, 16'd6098, 16'd53512, 16'd33751, 16'd8481, 16'd34998});
	test_expansion(128'h537ca78648291dead4ccac28944e2119, {16'd12157, 16'd40792, 16'd2304, 16'd42035, 16'd3269, 16'd16058, 16'd53176, 16'd9431, 16'd11881, 16'd29221, 16'd8484, 16'd4472, 16'd5257, 16'd4218, 16'd49454, 16'd18038, 16'd26637, 16'd41352, 16'd23607, 16'd40818, 16'd55621, 16'd34995, 16'd10452, 16'd45466, 16'd64923, 16'd4489});
	test_expansion(128'hc9e86faf0b88f020ee4330d7a003597a, {16'd32227, 16'd48142, 16'd57703, 16'd13163, 16'd64261, 16'd31155, 16'd44708, 16'd37688, 16'd59465, 16'd28823, 16'd32907, 16'd35226, 16'd57351, 16'd15923, 16'd48781, 16'd38482, 16'd57733, 16'd27498, 16'd33220, 16'd22514, 16'd50848, 16'd48857, 16'd62165, 16'd60372, 16'd11523, 16'd779});
	test_expansion(128'h87ca0e24bfede9a0bcf474249e28344a, {16'd57275, 16'd930, 16'd33285, 16'd49518, 16'd50489, 16'd32400, 16'd28844, 16'd18238, 16'd7273, 16'd64353, 16'd5868, 16'd33798, 16'd8735, 16'd30400, 16'd50757, 16'd33691, 16'd40606, 16'd8737, 16'd5547, 16'd31879, 16'd4013, 16'd11777, 16'd29838, 16'd39189, 16'd22737, 16'd14082});
	test_expansion(128'h4b6c0da7acf32efbdcf66ab4c32953d5, {16'd10407, 16'd29713, 16'd14556, 16'd13002, 16'd24199, 16'd51908, 16'd6698, 16'd16416, 16'd40172, 16'd35613, 16'd25512, 16'd49588, 16'd54508, 16'd45641, 16'd42415, 16'd5662, 16'd50417, 16'd12248, 16'd52945, 16'd30434, 16'd48359, 16'd37844, 16'd38125, 16'd17723, 16'd12130, 16'd49693});
	test_expansion(128'h480be66265bac3b0e6a0c385a355f84c, {16'd51378, 16'd19392, 16'd41404, 16'd23891, 16'd64107, 16'd8825, 16'd16393, 16'd51704, 16'd64128, 16'd49691, 16'd10859, 16'd2878, 16'd29022, 16'd16391, 16'd14503, 16'd10969, 16'd39749, 16'd20508, 16'd52986, 16'd7681, 16'd33768, 16'd19409, 16'd14765, 16'd30106, 16'd7010, 16'd26413});
	test_expansion(128'hc385e5cbc1360143de083b3c4e9d6d91, {16'd11047, 16'd19238, 16'd61651, 16'd27649, 16'd20427, 16'd64186, 16'd41146, 16'd55372, 16'd40470, 16'd44304, 16'd13396, 16'd48594, 16'd62384, 16'd53116, 16'd59750, 16'd44484, 16'd38006, 16'd59911, 16'd41452, 16'd30479, 16'd6588, 16'd33325, 16'd61604, 16'd11554, 16'd6211, 16'd40523});
	test_expansion(128'ha01724c16357ac77af812fe459bb372c, {16'd41106, 16'd65136, 16'd32475, 16'd2315, 16'd64007, 16'd7587, 16'd63333, 16'd49120, 16'd60481, 16'd60500, 16'd57060, 16'd63239, 16'd26149, 16'd41093, 16'd16708, 16'd9483, 16'd33864, 16'd8216, 16'd61740, 16'd59840, 16'd35186, 16'd62921, 16'd47830, 16'd30257, 16'd64864, 16'd24539});
	test_expansion(128'h369ce1148a4d7f7b0d4aac9ec1777f55, {16'd53612, 16'd56948, 16'd45071, 16'd46103, 16'd15028, 16'd48193, 16'd63924, 16'd1803, 16'd4068, 16'd42667, 16'd182, 16'd17219, 16'd41097, 16'd13088, 16'd12713, 16'd8328, 16'd34542, 16'd13999, 16'd62338, 16'd8171, 16'd55930, 16'd6481, 16'd8525, 16'd57125, 16'd26988, 16'd15334});
	test_expansion(128'h6c96b9854f12dad256fa99a5bce0a597, {16'd55898, 16'd4653, 16'd50881, 16'd35144, 16'd42454, 16'd16692, 16'd7801, 16'd63518, 16'd41610, 16'd59162, 16'd38054, 16'd46160, 16'd14011, 16'd13232, 16'd7977, 16'd38413, 16'd57677, 16'd34600, 16'd30689, 16'd58143, 16'd21884, 16'd18276, 16'd42856, 16'd34554, 16'd14778, 16'd37156});
	test_expansion(128'h47f108f94418af569e4ca41785fcd70b, {16'd48380, 16'd49619, 16'd9220, 16'd23932, 16'd22623, 16'd37706, 16'd53465, 16'd43170, 16'd7954, 16'd45626, 16'd4847, 16'd16759, 16'd56029, 16'd41844, 16'd20326, 16'd14651, 16'd30803, 16'd8282, 16'd31909, 16'd28659, 16'd21333, 16'd9715, 16'd51727, 16'd30195, 16'd58007, 16'd42657});
	test_expansion(128'h41f121ef83b78e373e5345aaba552f97, {16'd10563, 16'd4386, 16'd6484, 16'd15628, 16'd5101, 16'd60380, 16'd57109, 16'd11311, 16'd55103, 16'd34034, 16'd38431, 16'd42717, 16'd47630, 16'd52360, 16'd43174, 16'd52576, 16'd6841, 16'd1942, 16'd62096, 16'd24888, 16'd48852, 16'd38858, 16'd34125, 16'd25689, 16'd54781, 16'd22355});
	test_expansion(128'h103f99cf8622fd4e171ee46dbbf78d7b, {16'd31154, 16'd35033, 16'd42224, 16'd53179, 16'd26156, 16'd11148, 16'd61812, 16'd37409, 16'd6609, 16'd50535, 16'd48016, 16'd17873, 16'd3370, 16'd28650, 16'd43289, 16'd15861, 16'd62229, 16'd2347, 16'd26614, 16'd50325, 16'd55439, 16'd23371, 16'd27539, 16'd15623, 16'd6703, 16'd17309});
	test_expansion(128'hf5d547b5a3b6ff4f57d38c83f3d9662d, {16'd13722, 16'd47247, 16'd51507, 16'd56234, 16'd9728, 16'd19990, 16'd37909, 16'd20306, 16'd23565, 16'd5039, 16'd4702, 16'd3816, 16'd65445, 16'd30556, 16'd49263, 16'd61300, 16'd19922, 16'd49641, 16'd37292, 16'd18340, 16'd55670, 16'd31384, 16'd37798, 16'd12945, 16'd40221, 16'd51899});
	test_expansion(128'h6ef7a825c46231386d85feff3050c92e, {16'd6117, 16'd57073, 16'd11037, 16'd49655, 16'd64002, 16'd184, 16'd62221, 16'd65197, 16'd15185, 16'd12552, 16'd15963, 16'd4209, 16'd10448, 16'd33666, 16'd58082, 16'd3196, 16'd58349, 16'd34119, 16'd47669, 16'd5987, 16'd50264, 16'd30667, 16'd8933, 16'd30577, 16'd45819, 16'd39261});
	test_expansion(128'h306b9f8a1377fc67f8f73bfe8787e1fa, {16'd28683, 16'd58533, 16'd17676, 16'd17343, 16'd13349, 16'd6124, 16'd52490, 16'd38061, 16'd60701, 16'd7205, 16'd19365, 16'd63724, 16'd61581, 16'd37847, 16'd54466, 16'd28355, 16'd54735, 16'd23498, 16'd28630, 16'd34405, 16'd32164, 16'd899, 16'd60898, 16'd14001, 16'd14013, 16'd47673});
	test_expansion(128'hc6ae8298336bc3ccb657e2fe14190c13, {16'd33841, 16'd34761, 16'd17063, 16'd17055, 16'd52431, 16'd5366, 16'd45980, 16'd57067, 16'd43089, 16'd11167, 16'd17957, 16'd3876, 16'd27803, 16'd60295, 16'd61664, 16'd9161, 16'd64265, 16'd38630, 16'd36328, 16'd60598, 16'd51720, 16'd49500, 16'd49229, 16'd21347, 16'd54901, 16'd33245});
	test_expansion(128'h310efeabe74afeed65202ad8c59e8aab, {16'd46094, 16'd31043, 16'd8692, 16'd27002, 16'd55853, 16'd9217, 16'd55330, 16'd11324, 16'd25965, 16'd3262, 16'd32063, 16'd37745, 16'd42922, 16'd64603, 16'd25307, 16'd47002, 16'd19702, 16'd61157, 16'd12535, 16'd22870, 16'd27285, 16'd23141, 16'd24240, 16'd17398, 16'd19867, 16'd20761});
	test_expansion(128'h0a8382a1e22df87e2d66d304a8cd1821, {16'd8742, 16'd38834, 16'd49421, 16'd49549, 16'd36325, 16'd59988, 16'd47876, 16'd16484, 16'd58041, 16'd63025, 16'd47526, 16'd21196, 16'd44127, 16'd44149, 16'd45980, 16'd9383, 16'd33188, 16'd45622, 16'd48539, 16'd15145, 16'd21802, 16'd51097, 16'd10948, 16'd36596, 16'd42058, 16'd54685});
	test_expansion(128'h382df6617ff9269657de14330c1cbee8, {16'd60983, 16'd49538, 16'd3808, 16'd56, 16'd25331, 16'd30114, 16'd50734, 16'd49109, 16'd21953, 16'd33827, 16'd35240, 16'd31216, 16'd9672, 16'd50222, 16'd16773, 16'd61840, 16'd35234, 16'd13514, 16'd27496, 16'd60153, 16'd4136, 16'd39643, 16'd59471, 16'd43611, 16'd2710, 16'd60006});
	test_expansion(128'h6895bb2b2dcad30741de3a2167bf1b57, {16'd2543, 16'd60424, 16'd19253, 16'd46752, 16'd31277, 16'd27013, 16'd11990, 16'd11574, 16'd5592, 16'd11341, 16'd8407, 16'd55609, 16'd24402, 16'd54824, 16'd21350, 16'd27108, 16'd38547, 16'd47874, 16'd37962, 16'd60774, 16'd9865, 16'd37781, 16'd42023, 16'd41455, 16'd505, 16'd16140});
	test_expansion(128'ha8cedaab13a8b0deaf51bcd0c9361b16, {16'd50257, 16'd25523, 16'd7156, 16'd42402, 16'd24510, 16'd46871, 16'd21960, 16'd18104, 16'd31647, 16'd35429, 16'd26309, 16'd49975, 16'd55238, 16'd35055, 16'd38720, 16'd61913, 16'd16197, 16'd56130, 16'd29649, 16'd37405, 16'd51592, 16'd1548, 16'd47129, 16'd3816, 16'd19465, 16'd43553});
	test_expansion(128'h812644747a04c9bb0dd0fe7f42f62096, {16'd43206, 16'd21427, 16'd44904, 16'd50252, 16'd16720, 16'd64858, 16'd49319, 16'd51502, 16'd1839, 16'd3637, 16'd61623, 16'd52662, 16'd27565, 16'd53381, 16'd55883, 16'd6162, 16'd32308, 16'd59732, 16'd18739, 16'd29088, 16'd10434, 16'd5112, 16'd1219, 16'd50563, 16'd18976, 16'd25147});
	test_expansion(128'hb4202126c753e557760d571bcaf41e1a, {16'd10445, 16'd35011, 16'd62407, 16'd2084, 16'd38569, 16'd37004, 16'd35179, 16'd51563, 16'd59539, 16'd47387, 16'd29728, 16'd53608, 16'd23331, 16'd27443, 16'd20892, 16'd22881, 16'd43672, 16'd10959, 16'd49208, 16'd54017, 16'd3325, 16'd51993, 16'd20312, 16'd32185, 16'd7376, 16'd36684});
	test_expansion(128'h704f503a021c3f05f23caf5ea7fe9111, {16'd5245, 16'd39146, 16'd6495, 16'd45429, 16'd4765, 16'd64707, 16'd1507, 16'd19848, 16'd26593, 16'd60020, 16'd57255, 16'd10710, 16'd53826, 16'd46132, 16'd27482, 16'd11376, 16'd58557, 16'd44836, 16'd40238, 16'd62754, 16'd60328, 16'd64190, 16'd28770, 16'd1747, 16'd5805, 16'd11354});
	test_expansion(128'hfb83dc694aaa8c79f952b7472e444cc4, {16'd37192, 16'd32707, 16'd60686, 16'd4936, 16'd63291, 16'd16738, 16'd50836, 16'd10409, 16'd58982, 16'd9875, 16'd17545, 16'd36242, 16'd33513, 16'd25236, 16'd18607, 16'd26849, 16'd49480, 16'd55128, 16'd55808, 16'd22681, 16'd50521, 16'd15479, 16'd34470, 16'd30937, 16'd26556, 16'd12282});
	test_expansion(128'hdb8bf1a087413d5869e35283dd4be691, {16'd1592, 16'd1039, 16'd16990, 16'd40540, 16'd8383, 16'd38208, 16'd48848, 16'd30459, 16'd47653, 16'd48010, 16'd3876, 16'd15740, 16'd42225, 16'd45480, 16'd11880, 16'd12687, 16'd32190, 16'd16872, 16'd23001, 16'd16078, 16'd64159, 16'd60248, 16'd188, 16'd23857, 16'd64578, 16'd61257});
	test_expansion(128'h41332e4f5cd8510ea395d5af6f9e4c78, {16'd8931, 16'd50232, 16'd56578, 16'd44404, 16'd12947, 16'd12941, 16'd31746, 16'd49280, 16'd48527, 16'd10091, 16'd36838, 16'd4137, 16'd60505, 16'd36508, 16'd60290, 16'd27126, 16'd4099, 16'd13808, 16'd16689, 16'd27157, 16'd20310, 16'd59924, 16'd5207, 16'd44862, 16'd52615, 16'd13289});
	test_expansion(128'h21950f2f82e6739efeb7fd724bba26d8, {16'd6899, 16'd26398, 16'd14482, 16'd47761, 16'd59509, 16'd30654, 16'd56707, 16'd64355, 16'd20336, 16'd1468, 16'd47625, 16'd15743, 16'd18623, 16'd20167, 16'd61645, 16'd51648, 16'd51821, 16'd50994, 16'd48169, 16'd59769, 16'd3920, 16'd26227, 16'd32480, 16'd1041, 16'd29113, 16'd50270});
	test_expansion(128'h94acdfc5f4d83f913576e9768b4bb511, {16'd3157, 16'd12978, 16'd31647, 16'd16161, 16'd36914, 16'd35875, 16'd11908, 16'd14477, 16'd48482, 16'd34325, 16'd39419, 16'd3459, 16'd20879, 16'd25231, 16'd1912, 16'd65121, 16'd35149, 16'd49263, 16'd2122, 16'd64597, 16'd173, 16'd22990, 16'd46420, 16'd39663, 16'd23012, 16'd14377});
	test_expansion(128'h238f160dd91f1731bf34fbb5d38f8dc7, {16'd65464, 16'd49182, 16'd40062, 16'd1157, 16'd54241, 16'd55586, 16'd57766, 16'd58326, 16'd2031, 16'd48646, 16'd51056, 16'd55683, 16'd11583, 16'd56661, 16'd50599, 16'd4861, 16'd52375, 16'd38858, 16'd49910, 16'd28694, 16'd16066, 16'd3210, 16'd2551, 16'd53752, 16'd36895, 16'd10011});
	test_expansion(128'hfb8cf300de47318a3f80dc2c48cc74f7, {16'd41264, 16'd39105, 16'd62103, 16'd39022, 16'd33949, 16'd45252, 16'd2405, 16'd25259, 16'd46711, 16'd29032, 16'd26168, 16'd4096, 16'd14557, 16'd11197, 16'd1022, 16'd20640, 16'd9970, 16'd8178, 16'd22588, 16'd14312, 16'd47071, 16'd22178, 16'd3443, 16'd65082, 16'd51710, 16'd2459});
	test_expansion(128'h176b2d684d458f18ca2706e19514d521, {16'd4984, 16'd28937, 16'd60437, 16'd51551, 16'd61479, 16'd1771, 16'd42798, 16'd61497, 16'd1583, 16'd55873, 16'd49089, 16'd6587, 16'd46721, 16'd7585, 16'd36427, 16'd58100, 16'd770, 16'd5507, 16'd41906, 16'd14334, 16'd12838, 16'd1921, 16'd29921, 16'd10565, 16'd25417, 16'd25873});
	test_expansion(128'h5953eb34fbbf0b742b52733e4580a5d3, {16'd38693, 16'd20037, 16'd35554, 16'd62783, 16'd36827, 16'd15092, 16'd36722, 16'd5885, 16'd27742, 16'd59350, 16'd59530, 16'd33096, 16'd31134, 16'd21168, 16'd49007, 16'd2027, 16'd44641, 16'd12277, 16'd23391, 16'd27646, 16'd11192, 16'd50315, 16'd1926, 16'd8277, 16'd42836, 16'd52438});
	test_expansion(128'h22fc06557f29afdaca13e0c8b35dbc87, {16'd49958, 16'd43870, 16'd25490, 16'd63739, 16'd43464, 16'd45418, 16'd17772, 16'd28703, 16'd59376, 16'd11005, 16'd48531, 16'd17086, 16'd5031, 16'd16496, 16'd54177, 16'd26524, 16'd55478, 16'd34149, 16'd46256, 16'd15073, 16'd3879, 16'd42023, 16'd36784, 16'd11488, 16'd46324, 16'd38974});
	test_expansion(128'h76cccf5f3ea38aa753a55a28ee9136b4, {16'd31324, 16'd12861, 16'd56412, 16'd50003, 16'd44353, 16'd29183, 16'd59113, 16'd29695, 16'd63288, 16'd6032, 16'd38655, 16'd53888, 16'd4411, 16'd37405, 16'd19874, 16'd45034, 16'd16407, 16'd21509, 16'd14857, 16'd8925, 16'd50990, 16'd37155, 16'd33553, 16'd9629, 16'd17939, 16'd7344});
	test_expansion(128'hcb1435ea6f177f22c74997f9c768bdf7, {16'd62739, 16'd17970, 16'd62295, 16'd20758, 16'd47891, 16'd37839, 16'd10802, 16'd8857, 16'd18024, 16'd61815, 16'd10890, 16'd47411, 16'd12743, 16'd32608, 16'd53957, 16'd19439, 16'd6633, 16'd21051, 16'd49411, 16'd12568, 16'd10947, 16'd23762, 16'd32343, 16'd60664, 16'd12459, 16'd64838});
	test_expansion(128'h97220cd693b1cf16a1aeb9c3e4982bd1, {16'd65101, 16'd9420, 16'd41227, 16'd39174, 16'd1200, 16'd37745, 16'd56960, 16'd28852, 16'd170, 16'd62481, 16'd60158, 16'd7139, 16'd34713, 16'd13097, 16'd6766, 16'd41477, 16'd55880, 16'd44623, 16'd22402, 16'd65204, 16'd35483, 16'd22596, 16'd17691, 16'd11254, 16'd17095, 16'd53056});
	test_expansion(128'h618bec7a0e84787482fcaa17b7070864, {16'd42532, 16'd21825, 16'd46342, 16'd41562, 16'd34783, 16'd43644, 16'd56274, 16'd42037, 16'd5461, 16'd63101, 16'd9923, 16'd36105, 16'd8312, 16'd23736, 16'd43637, 16'd37932, 16'd27915, 16'd26622, 16'd61795, 16'd40946, 16'd22417, 16'd35481, 16'd5828, 16'd47691, 16'd50716, 16'd53358});
	test_expansion(128'h2ecb9890ca838abc832cbe5d4e37cf90, {16'd57939, 16'd30218, 16'd3965, 16'd32713, 16'd41000, 16'd38157, 16'd48429, 16'd28045, 16'd34540, 16'd55622, 16'd22594, 16'd55278, 16'd21889, 16'd19835, 16'd56310, 16'd35552, 16'd21853, 16'd32579, 16'd15987, 16'd1546, 16'd41420, 16'd52561, 16'd1787, 16'd64271, 16'd14112, 16'd57777});
	test_expansion(128'h75a6652a861c023bfd007e3020b970b9, {16'd44770, 16'd41789, 16'd58624, 16'd60722, 16'd39787, 16'd60540, 16'd19557, 16'd46892, 16'd47696, 16'd22829, 16'd21811, 16'd26961, 16'd48269, 16'd39092, 16'd3356, 16'd14031, 16'd35725, 16'd64738, 16'd59863, 16'd4161, 16'd27223, 16'd59790, 16'd19624, 16'd47215, 16'd64582, 16'd46307});
	test_expansion(128'h647f8946fc372c0f3b035cccf118fa75, {16'd60854, 16'd54936, 16'd43187, 16'd57078, 16'd36056, 16'd48306, 16'd48323, 16'd46438, 16'd12156, 16'd4583, 16'd30047, 16'd39481, 16'd4734, 16'd42350, 16'd3560, 16'd46124, 16'd44960, 16'd32401, 16'd46688, 16'd14736, 16'd49492, 16'd56557, 16'd1292, 16'd58605, 16'd4063, 16'd43764});
	test_expansion(128'hc55ace7871d9ac251224d641953e7f5f, {16'd23468, 16'd49372, 16'd8845, 16'd53519, 16'd44968, 16'd3923, 16'd35218, 16'd29999, 16'd44099, 16'd1877, 16'd14848, 16'd12160, 16'd51206, 16'd62076, 16'd16205, 16'd47316, 16'd11060, 16'd12274, 16'd5259, 16'd45734, 16'd7159, 16'd55065, 16'd31831, 16'd22814, 16'd35657, 16'd20222});
	test_expansion(128'hd9bf922709fb472cec403619c179401c, {16'd5903, 16'd36644, 16'd7992, 16'd46389, 16'd31925, 16'd51664, 16'd23213, 16'd32817, 16'd45469, 16'd6650, 16'd57269, 16'd15113, 16'd40377, 16'd34991, 16'd10282, 16'd62834, 16'd55681, 16'd33655, 16'd15690, 16'd34131, 16'd36337, 16'd18819, 16'd60014, 16'd33991, 16'd34675, 16'd35432});
	test_expansion(128'h467e0a66b31561e66fbeaabfcbe419f3, {16'd47865, 16'd20788, 16'd62829, 16'd39020, 16'd14972, 16'd11237, 16'd43265, 16'd12273, 16'd37912, 16'd11698, 16'd3692, 16'd62825, 16'd11469, 16'd34951, 16'd46464, 16'd48458, 16'd57642, 16'd47414, 16'd21613, 16'd39904, 16'd12431, 16'd13093, 16'd13, 16'd46222, 16'd5796, 16'd30757});
	test_expansion(128'h4c0f27cdec3492aca094a97d02505cfd, {16'd50366, 16'd30133, 16'd20046, 16'd23546, 16'd32066, 16'd35773, 16'd43604, 16'd64442, 16'd50615, 16'd30702, 16'd38837, 16'd30736, 16'd21380, 16'd37521, 16'd7281, 16'd57589, 16'd24648, 16'd7444, 16'd27405, 16'd23977, 16'd52619, 16'd23710, 16'd48693, 16'd8016, 16'd62082, 16'd57015});
	test_expansion(128'h3b351a9934886f0d08e524cb48abd814, {16'd24172, 16'd9890, 16'd54998, 16'd25120, 16'd32879, 16'd27972, 16'd36224, 16'd64270, 16'd64492, 16'd59323, 16'd40690, 16'd30689, 16'd24624, 16'd38424, 16'd10115, 16'd42033, 16'd8638, 16'd51591, 16'd25369, 16'd44763, 16'd25932, 16'd59241, 16'd30301, 16'd27516, 16'd23135, 16'd41146});
	test_expansion(128'h2b7599318730bc1e942e856b00183d55, {16'd21982, 16'd5488, 16'd47696, 16'd143, 16'd65505, 16'd59524, 16'd22524, 16'd19121, 16'd25945, 16'd65496, 16'd48480, 16'd1002, 16'd60258, 16'd30631, 16'd25378, 16'd38198, 16'd45543, 16'd8692, 16'd21497, 16'd6595, 16'd45076, 16'd52697, 16'd61205, 16'd20614, 16'd56568, 16'd55405});
	test_expansion(128'hc653260bf56a24fc37665d90feb28a9e, {16'd45824, 16'd14661, 16'd2398, 16'd970, 16'd34908, 16'd34024, 16'd24517, 16'd30016, 16'd54369, 16'd6104, 16'd36724, 16'd41481, 16'd9148, 16'd54957, 16'd45885, 16'd2637, 16'd52845, 16'd47094, 16'd37503, 16'd4858, 16'd59172, 16'd48949, 16'd14318, 16'd57611, 16'd58449, 16'd27502});
	test_expansion(128'h2e874e2d187db5bcc9fbf710c91d08c9, {16'd27551, 16'd11532, 16'd59793, 16'd51365, 16'd4775, 16'd29729, 16'd12746, 16'd65092, 16'd8, 16'd17418, 16'd52611, 16'd13641, 16'd46714, 16'd16212, 16'd58115, 16'd41200, 16'd13403, 16'd49798, 16'd17421, 16'd12032, 16'd25051, 16'd64989, 16'd56691, 16'd47293, 16'd44992, 16'd31343});
	test_expansion(128'hf976db111ca87c1b1dd0e1a06206020e, {16'd64569, 16'd23498, 16'd35282, 16'd27902, 16'd8912, 16'd1990, 16'd30731, 16'd44459, 16'd39301, 16'd48697, 16'd5295, 16'd15804, 16'd9752, 16'd61598, 16'd4299, 16'd29600, 16'd54939, 16'd64685, 16'd34239, 16'd30725, 16'd8770, 16'd5317, 16'd30129, 16'd20616, 16'd61874, 16'd5631});
	test_expansion(128'h84de8dbe1ff575f90f81249c8fbde37d, {16'd62341, 16'd854, 16'd30086, 16'd35838, 16'd18109, 16'd58466, 16'd59506, 16'd52877, 16'd14579, 16'd19857, 16'd16738, 16'd33720, 16'd48162, 16'd63636, 16'd35189, 16'd52117, 16'd21222, 16'd59258, 16'd34578, 16'd17762, 16'd14928, 16'd61707, 16'd45773, 16'd24962, 16'd55860, 16'd62806});
	test_expansion(128'h30fa9ac1c71525ade4671b42fedca9c4, {16'd25562, 16'd1006, 16'd37742, 16'd36379, 16'd42521, 16'd63853, 16'd943, 16'd35011, 16'd22617, 16'd64026, 16'd40797, 16'd60497, 16'd50200, 16'd41325, 16'd21130, 16'd52303, 16'd20452, 16'd41062, 16'd23696, 16'd27598, 16'd44820, 16'd33712, 16'd25429, 16'd58265, 16'd45546, 16'd58986});
	test_expansion(128'h3def4afba3897eb154c4231a75759d04, {16'd34583, 16'd53181, 16'd57786, 16'd2234, 16'd383, 16'd10093, 16'd37263, 16'd52295, 16'd2826, 16'd47797, 16'd17218, 16'd58624, 16'd18837, 16'd43274, 16'd10896, 16'd46152, 16'd61933, 16'd58994, 16'd33827, 16'd21263, 16'd18258, 16'd19913, 16'd28817, 16'd64958, 16'd34241, 16'd20843});
	test_expansion(128'hc581e358b5ef50ed47cae0d0d2f53592, {16'd20054, 16'd35967, 16'd10236, 16'd25768, 16'd9570, 16'd47923, 16'd37249, 16'd37881, 16'd43708, 16'd62339, 16'd4891, 16'd39225, 16'd57562, 16'd31511, 16'd10343, 16'd61153, 16'd25002, 16'd58222, 16'd48574, 16'd46355, 16'd11521, 16'd10819, 16'd61549, 16'd44747, 16'd1753, 16'd53845});
	test_expansion(128'h2908a95b22bc58eac2fabd0769275f7f, {16'd10154, 16'd59702, 16'd14525, 16'd63478, 16'd5248, 16'd9293, 16'd55168, 16'd45878, 16'd42522, 16'd52666, 16'd60333, 16'd64374, 16'd15419, 16'd62439, 16'd35895, 16'd12025, 16'd31792, 16'd14137, 16'd62244, 16'd51084, 16'd12192, 16'd10915, 16'd23136, 16'd44079, 16'd33664, 16'd43632});
	test_expansion(128'hd7ded8b1888cde7cbc17fa574ec16498, {16'd614, 16'd21458, 16'd53670, 16'd33770, 16'd51052, 16'd61684, 16'd39339, 16'd25272, 16'd18851, 16'd61827, 16'd21460, 16'd62945, 16'd16889, 16'd39915, 16'd25400, 16'd56517, 16'd31969, 16'd974, 16'd5833, 16'd8787, 16'd6760, 16'd1784, 16'd34161, 16'd42705, 16'd11044, 16'd13188});
	test_expansion(128'h48fca29d109ce84dededf062f6ceeb67, {16'd32733, 16'd9077, 16'd58432, 16'd41482, 16'd28024, 16'd49000, 16'd6286, 16'd25513, 16'd2499, 16'd33502, 16'd59849, 16'd14443, 16'd18101, 16'd36210, 16'd9844, 16'd11438, 16'd63709, 16'd28815, 16'd61431, 16'd8277, 16'd37498, 16'd31690, 16'd42285, 16'd64154, 16'd803, 16'd31269});
	test_expansion(128'h201de9749a07a78b1dd4321e42dc0194, {16'd60938, 16'd2754, 16'd41063, 16'd28270, 16'd3926, 16'd47169, 16'd26100, 16'd33057, 16'd60329, 16'd35677, 16'd1858, 16'd63394, 16'd31060, 16'd29814, 16'd1568, 16'd14863, 16'd1653, 16'd61838, 16'd7469, 16'd52054, 16'd16911, 16'd32633, 16'd46182, 16'd23002, 16'd20462, 16'd4387});
	test_expansion(128'h9471ef564210df56e90ba231f7a5fe7b, {16'd20865, 16'd25118, 16'd13427, 16'd18831, 16'd38072, 16'd8419, 16'd24309, 16'd60865, 16'd40820, 16'd61228, 16'd7532, 16'd32608, 16'd47030, 16'd37128, 16'd6527, 16'd30068, 16'd9941, 16'd16828, 16'd39924, 16'd16735, 16'd43499, 16'd59761, 16'd34637, 16'd31180, 16'd16141, 16'd9351});
	test_expansion(128'h868dfb7ac87f344665ed25b5fbef2d19, {16'd9583, 16'd17024, 16'd7977, 16'd15756, 16'd52872, 16'd54150, 16'd4078, 16'd17133, 16'd23679, 16'd53434, 16'd65319, 16'd43953, 16'd7351, 16'd16783, 16'd62681, 16'd28004, 16'd39987, 16'd837, 16'd22056, 16'd35508, 16'd26299, 16'd25750, 16'd46333, 16'd28620, 16'd23182, 16'd40556});
	test_expansion(128'h8ce774c2475ac54c7b48047137bc217d, {16'd7213, 16'd24399, 16'd25514, 16'd8286, 16'd50451, 16'd42500, 16'd26949, 16'd16296, 16'd9377, 16'd748, 16'd17865, 16'd14713, 16'd37267, 16'd62700, 16'd60653, 16'd49759, 16'd54676, 16'd25091, 16'd16011, 16'd54637, 16'd55330, 16'd47566, 16'd16206, 16'd23523, 16'd41649, 16'd2637});
	test_expansion(128'hf7ed91f6793b2c1fbe45009f4891a938, {16'd31655, 16'd30118, 16'd9559, 16'd3617, 16'd20082, 16'd12628, 16'd16593, 16'd64218, 16'd63263, 16'd4911, 16'd29384, 16'd34723, 16'd7612, 16'd53765, 16'd59189, 16'd24938, 16'd41195, 16'd11307, 16'd38407, 16'd9242, 16'd34462, 16'd27270, 16'd37288, 16'd50985, 16'd37647, 16'd3991});
	test_expansion(128'h852c62eab45ccc8aa735c92c1243fdfc, {16'd54782, 16'd32898, 16'd54684, 16'd38909, 16'd60257, 16'd58146, 16'd11786, 16'd63930, 16'd58824, 16'd43249, 16'd45549, 16'd47152, 16'd10791, 16'd31196, 16'd42528, 16'd47384, 16'd44066, 16'd45148, 16'd20979, 16'd43517, 16'd957, 16'd50692, 16'd40365, 16'd62166, 16'd42433, 16'd54964});
	test_expansion(128'hf49530876e0e213f977686c2c4462f71, {16'd54887, 16'd64073, 16'd2225, 16'd12674, 16'd10584, 16'd22069, 16'd28153, 16'd26774, 16'd28036, 16'd44431, 16'd36691, 16'd36931, 16'd31221, 16'd8689, 16'd16790, 16'd38341, 16'd32902, 16'd21782, 16'd18377, 16'd31205, 16'd19547, 16'd14383, 16'd48386, 16'd14565, 16'd33814, 16'd47215});
	test_expansion(128'h90cb54cf0eef74f98faed1659c3f7335, {16'd64001, 16'd21628, 16'd31554, 16'd11626, 16'd48970, 16'd11383, 16'd42289, 16'd11919, 16'd13215, 16'd34463, 16'd43325, 16'd30373, 16'd59229, 16'd55678, 16'd19239, 16'd62738, 16'd53731, 16'd61055, 16'd4556, 16'd1066, 16'd14603, 16'd37481, 16'd51656, 16'd6536, 16'd65395, 16'd27561});
	test_expansion(128'h3f24d38e5d89472ab53303d55fd4200c, {16'd23873, 16'd50179, 16'd32085, 16'd40593, 16'd62531, 16'd15141, 16'd48507, 16'd30754, 16'd1694, 16'd22930, 16'd393, 16'd31375, 16'd22138, 16'd6452, 16'd43482, 16'd886, 16'd2299, 16'd42262, 16'd21375, 16'd10414, 16'd45472, 16'd16016, 16'd59793, 16'd19341, 16'd47446, 16'd28571});
	test_expansion(128'h49fa31bda5d901990384df7f35dbf94e, {16'd30262, 16'd19881, 16'd30703, 16'd23134, 16'd37658, 16'd47871, 16'd24536, 16'd21337, 16'd16669, 16'd62260, 16'd20689, 16'd5715, 16'd23094, 16'd61100, 16'd22777, 16'd51069, 16'd13207, 16'd46859, 16'd56391, 16'd25736, 16'd27618, 16'd50765, 16'd6217, 16'd32034, 16'd37796, 16'd50941});
	test_expansion(128'hcc1ee99e0702c6c8dba05dc6cad8e39b, {16'd5163, 16'd5303, 16'd62300, 16'd20156, 16'd14967, 16'd59906, 16'd19061, 16'd52753, 16'd51540, 16'd50958, 16'd34016, 16'd38408, 16'd25968, 16'd59683, 16'd53287, 16'd33911, 16'd41600, 16'd22881, 16'd47052, 16'd40014, 16'd41576, 16'd55617, 16'd18643, 16'd9933, 16'd38182, 16'd19254});
	test_expansion(128'h2c3db765d409c6748330df0621385744, {16'd54685, 16'd60984, 16'd27203, 16'd18517, 16'd25705, 16'd32436, 16'd47478, 16'd48147, 16'd57643, 16'd20417, 16'd13374, 16'd12560, 16'd54105, 16'd16373, 16'd15018, 16'd12986, 16'd33860, 16'd31924, 16'd11789, 16'd30770, 16'd50766, 16'd61569, 16'd43571, 16'd53943, 16'd46572, 16'd48146});
	test_expansion(128'h8f9f58e485ef4029f79746a4db2c55b5, {16'd27013, 16'd47165, 16'd29840, 16'd59948, 16'd18250, 16'd46749, 16'd59296, 16'd14756, 16'd2175, 16'd38548, 16'd19664, 16'd26425, 16'd24605, 16'd50882, 16'd18424, 16'd38883, 16'd44253, 16'd24795, 16'd64573, 16'd8926, 16'd28085, 16'd30848, 16'd48335, 16'd40279, 16'd14920, 16'd58444});
	test_expansion(128'h8e9cd7d051ed24d47beb95d992aa1f11, {16'd41471, 16'd40412, 16'd25124, 16'd37926, 16'd59483, 16'd5872, 16'd28192, 16'd30539, 16'd41168, 16'd49007, 16'd31196, 16'd24710, 16'd48964, 16'd21835, 16'd62196, 16'd24142, 16'd14938, 16'd38683, 16'd34599, 16'd9083, 16'd54447, 16'd29726, 16'd15911, 16'd22034, 16'd39871, 16'd51708});
	test_expansion(128'h6b86e0e21f8088fc0ead6a1070b802ec, {16'd58099, 16'd3001, 16'd50367, 16'd32400, 16'd26341, 16'd26375, 16'd27997, 16'd18352, 16'd24047, 16'd40647, 16'd23999, 16'd25398, 16'd57436, 16'd59325, 16'd27852, 16'd2853, 16'd49714, 16'd6046, 16'd25365, 16'd42199, 16'd28611, 16'd22592, 16'd18157, 16'd23306, 16'd24416, 16'd9176});
	test_expansion(128'haa0d765c76bd8fa2a04ac3cb8ee2c526, {16'd13929, 16'd19797, 16'd54924, 16'd65192, 16'd43546, 16'd25625, 16'd44259, 16'd14618, 16'd51717, 16'd50116, 16'd1462, 16'd31557, 16'd28182, 16'd48510, 16'd13719, 16'd49265, 16'd26722, 16'd32113, 16'd35550, 16'd20050, 16'd14531, 16'd12529, 16'd14538, 16'd26659, 16'd26597, 16'd34196});
	test_expansion(128'he3cae460858ef20843cfcbf47418f275, {16'd39062, 16'd51861, 16'd41246, 16'd51379, 16'd36219, 16'd10074, 16'd62495, 16'd61482, 16'd21692, 16'd50335, 16'd21735, 16'd22794, 16'd17288, 16'd33743, 16'd44699, 16'd56943, 16'd49785, 16'd18968, 16'd2633, 16'd62664, 16'd20911, 16'd24990, 16'd49855, 16'd7779, 16'd31803, 16'd19959});
	test_expansion(128'hb122ffa07e25c0d12a27531a82ebaba2, {16'd5418, 16'd49984, 16'd22178, 16'd22661, 16'd58937, 16'd53742, 16'd10309, 16'd30342, 16'd53632, 16'd45673, 16'd38927, 16'd57050, 16'd38867, 16'd2860, 16'd26809, 16'd58094, 16'd46993, 16'd42786, 16'd15858, 16'd50004, 16'd61359, 16'd24062, 16'd40509, 16'd33337, 16'd36764, 16'd60193});
	test_expansion(128'ha9301e66da3967092616eb1c2d304a92, {16'd18503, 16'd57679, 16'd36663, 16'd43948, 16'd22132, 16'd59130, 16'd44737, 16'd22691, 16'd33392, 16'd4469, 16'd40327, 16'd31372, 16'd140, 16'd35899, 16'd64249, 16'd50486, 16'd36723, 16'd27185, 16'd60037, 16'd7121, 16'd8050, 16'd54508, 16'd1761, 16'd30197, 16'd18036, 16'd8520});
	test_expansion(128'h0eec2c727af674e41b7818a3cc55c74f, {16'd35297, 16'd53050, 16'd3413, 16'd12279, 16'd58148, 16'd15498, 16'd56633, 16'd50127, 16'd55047, 16'd34672, 16'd32613, 16'd13345, 16'd57997, 16'd62071, 16'd45196, 16'd5708, 16'd46115, 16'd31051, 16'd17157, 16'd50030, 16'd50875, 16'd12146, 16'd47855, 16'd8062, 16'd63921, 16'd11643});
	test_expansion(128'hf02d47fb63058d833cfbf087dbe637da, {16'd9308, 16'd64462, 16'd34346, 16'd38555, 16'd15301, 16'd45207, 16'd41748, 16'd13477, 16'd63556, 16'd41237, 16'd56878, 16'd48691, 16'd21207, 16'd35958, 16'd58987, 16'd13995, 16'd33208, 16'd27778, 16'd5850, 16'd12720, 16'd6896, 16'd49959, 16'd19381, 16'd14835, 16'd54737, 16'd16539});
	test_expansion(128'hc62d1dbaea158278f1fed39876d16983, {16'd1886, 16'd35936, 16'd32583, 16'd53097, 16'd10811, 16'd31907, 16'd62470, 16'd56946, 16'd12530, 16'd52744, 16'd1966, 16'd12483, 16'd45959, 16'd28450, 16'd50232, 16'd28315, 16'd14584, 16'd6275, 16'd41061, 16'd24469, 16'd57232, 16'd38591, 16'd60417, 16'd9387, 16'd47279, 16'd57168});
	test_expansion(128'hb7483696a67c0e38abb6cc21ba8854b1, {16'd36825, 16'd30978, 16'd18122, 16'd31003, 16'd14567, 16'd9254, 16'd51712, 16'd17661, 16'd18226, 16'd54273, 16'd35960, 16'd30368, 16'd9535, 16'd10539, 16'd38140, 16'd61693, 16'd61145, 16'd58405, 16'd6143, 16'd11804, 16'd11393, 16'd37603, 16'd28465, 16'd50939, 16'd276, 16'd41474});
	test_expansion(128'h6d803935065668059c01cb1e96a12f7e, {16'd742, 16'd920, 16'd61700, 16'd60819, 16'd22187, 16'd3519, 16'd36015, 16'd62686, 16'd28223, 16'd4738, 16'd36425, 16'd38378, 16'd63078, 16'd37993, 16'd29522, 16'd53120, 16'd28236, 16'd25369, 16'd22307, 16'd51860, 16'd40230, 16'd24430, 16'd20739, 16'd44567, 16'd14833, 16'd9541});
	test_expansion(128'heba36eb4985e48dd8a13f019490b9f22, {16'd36506, 16'd49812, 16'd27205, 16'd18231, 16'd11914, 16'd46959, 16'd18687, 16'd9010, 16'd3406, 16'd64514, 16'd41815, 16'd26560, 16'd64416, 16'd10740, 16'd42721, 16'd33064, 16'd39768, 16'd58525, 16'd13958, 16'd29302, 16'd40747, 16'd9040, 16'd37924, 16'd64761, 16'd45149, 16'd33714});
	test_expansion(128'hb7e1823f8bfb35eb7dec3849c641ade8, {16'd9604, 16'd39704, 16'd40522, 16'd20508, 16'd15222, 16'd49452, 16'd37035, 16'd14260, 16'd23234, 16'd44424, 16'd4065, 16'd30643, 16'd7807, 16'd59074, 16'd11389, 16'd11893, 16'd26663, 16'd27296, 16'd32185, 16'd27626, 16'd60410, 16'd23577, 16'd18793, 16'd48806, 16'd64320, 16'd15563});
	test_expansion(128'h23c7fd07eb9d9413d2a77951f010f08c, {16'd30219, 16'd15914, 16'd34673, 16'd38345, 16'd55623, 16'd46970, 16'd10869, 16'd54264, 16'd43013, 16'd53303, 16'd51167, 16'd16659, 16'd1352, 16'd12934, 16'd39288, 16'd10545, 16'd59366, 16'd46739, 16'd32747, 16'd41557, 16'd42633, 16'd1902, 16'd38919, 16'd20050, 16'd10048, 16'd44172});
	test_expansion(128'h9779634e3a2bd8da8df59982b6f6c38c, {16'd12685, 16'd42659, 16'd43015, 16'd23262, 16'd24639, 16'd19058, 16'd55710, 16'd19757, 16'd4620, 16'd44311, 16'd23840, 16'd28505, 16'd47006, 16'd27371, 16'd58774, 16'd4127, 16'd53574, 16'd2886, 16'd50763, 16'd34212, 16'd36135, 16'd27569, 16'd25193, 16'd53709, 16'd63146, 16'd47164});
	test_expansion(128'h2c44b975d1f6448a62b307ef1692619b, {16'd19342, 16'd5974, 16'd59536, 16'd48750, 16'd50162, 16'd32024, 16'd35448, 16'd44818, 16'd5730, 16'd42717, 16'd32678, 16'd17559, 16'd34041, 16'd27254, 16'd37980, 16'd55258, 16'd58353, 16'd55594, 16'd58841, 16'd53974, 16'd60272, 16'd22567, 16'd20967, 16'd48003, 16'd10632, 16'd21671});
	test_expansion(128'he1d4279bffbf81de030dc18bc9eff4b4, {16'd2048, 16'd12736, 16'd47242, 16'd7212, 16'd60863, 16'd11202, 16'd39494, 16'd9390, 16'd1141, 16'd52813, 16'd273, 16'd56415, 16'd34011, 16'd58565, 16'd22706, 16'd14070, 16'd8040, 16'd37600, 16'd51586, 16'd55392, 16'd16489, 16'd23370, 16'd26714, 16'd26553, 16'd44541, 16'd7732});
	test_expansion(128'h22d9a2e79e960727a9538466c7995479, {16'd55306, 16'd9717, 16'd16029, 16'd19113, 16'd17506, 16'd50343, 16'd26744, 16'd46722, 16'd28604, 16'd1437, 16'd1448, 16'd41821, 16'd63738, 16'd9136, 16'd34000, 16'd16284, 16'd47968, 16'd61424, 16'd5182, 16'd47281, 16'd21901, 16'd4956, 16'd6452, 16'd54241, 16'd58947, 16'd27162});
	test_expansion(128'hc0aa2fe10d520c3690b0a7a17e2e6574, {16'd58570, 16'd49602, 16'd16491, 16'd60660, 16'd2514, 16'd40221, 16'd25665, 16'd5179, 16'd47811, 16'd40033, 16'd29642, 16'd19456, 16'd48094, 16'd50570, 16'd7768, 16'd3250, 16'd3298, 16'd26009, 16'd60761, 16'd38691, 16'd6026, 16'd36643, 16'd28967, 16'd2092, 16'd11663, 16'd59061});
	test_expansion(128'h4f3bfcea62eff9b4dfe9beca02b6f8ea, {16'd4248, 16'd26958, 16'd42482, 16'd12654, 16'd37858, 16'd53114, 16'd472, 16'd14146, 16'd15821, 16'd37514, 16'd50896, 16'd32295, 16'd47914, 16'd8247, 16'd57972, 16'd42378, 16'd22751, 16'd8697, 16'd57316, 16'd37405, 16'd17838, 16'd24184, 16'd1923, 16'd26357, 16'd21623, 16'd9804});
	test_expansion(128'hc5166e90ef51c3583b52147c2d6cc875, {16'd5539, 16'd46951, 16'd33373, 16'd43885, 16'd48265, 16'd53299, 16'd48918, 16'd53979, 16'd5387, 16'd65163, 16'd8686, 16'd22222, 16'd59817, 16'd51789, 16'd5687, 16'd18022, 16'd38593, 16'd23603, 16'd62338, 16'd23135, 16'd55787, 16'd27907, 16'd733, 16'd40533, 16'd60998, 16'd48396});
	test_expansion(128'h9f9b5cc8617bf6f8e904c7a25989f69d, {16'd24839, 16'd50857, 16'd26471, 16'd10742, 16'd8720, 16'd19946, 16'd38201, 16'd55826, 16'd20857, 16'd65422, 16'd59746, 16'd48638, 16'd35846, 16'd40950, 16'd34553, 16'd31052, 16'd26387, 16'd40594, 16'd18389, 16'd56925, 16'd49982, 16'd23186, 16'd19247, 16'd50874, 16'd1933, 16'd49998});
	test_expansion(128'hfb85f25e83cb963538b888a496fc4ed1, {16'd28798, 16'd19350, 16'd24224, 16'd24943, 16'd31410, 16'd60821, 16'd52394, 16'd5190, 16'd36692, 16'd7262, 16'd61390, 16'd32566, 16'd3799, 16'd58277, 16'd17579, 16'd24963, 16'd57233, 16'd16954, 16'd19527, 16'd14938, 16'd10527, 16'd51260, 16'd1895, 16'd3213, 16'd33575, 16'd51487});
	test_expansion(128'h89f1e305e924e7e622b6eeca0195dae5, {16'd7445, 16'd43256, 16'd10001, 16'd8902, 16'd11747, 16'd31110, 16'd24690, 16'd58400, 16'd12377, 16'd44723, 16'd40598, 16'd23155, 16'd31458, 16'd15541, 16'd64531, 16'd63484, 16'd27180, 16'd48871, 16'd9412, 16'd31561, 16'd15403, 16'd42223, 16'd14829, 16'd58602, 16'd58310, 16'd31825});
	test_expansion(128'hc977cc6e30037ed0ef995c2e420a6052, {16'd58966, 16'd403, 16'd3115, 16'd33939, 16'd13478, 16'd32217, 16'd39649, 16'd35106, 16'd45756, 16'd22753, 16'd65416, 16'd46000, 16'd33710, 16'd63212, 16'd54123, 16'd1373, 16'd15152, 16'd21295, 16'd17290, 16'd59862, 16'd63558, 16'd34291, 16'd4211, 16'd55896, 16'd55385, 16'd59537});
	test_expansion(128'h9ce19079080910f537d495d918b77bc3, {16'd39525, 16'd49596, 16'd26647, 16'd45731, 16'd12430, 16'd22430, 16'd21190, 16'd31938, 16'd38639, 16'd31814, 16'd64786, 16'd4080, 16'd3718, 16'd54577, 16'd17656, 16'd44977, 16'd30051, 16'd25651, 16'd25588, 16'd51981, 16'd57145, 16'd10944, 16'd8116, 16'd21426, 16'd27224, 16'd34727});
	test_expansion(128'hee5cb0cd5e9c99363f92bfa9b20cc35d, {16'd54411, 16'd19811, 16'd57612, 16'd32322, 16'd13321, 16'd27265, 16'd24957, 16'd17884, 16'd65194, 16'd47220, 16'd52822, 16'd39764, 16'd21983, 16'd52413, 16'd60660, 16'd29705, 16'd60578, 16'd48832, 16'd50310, 16'd10541, 16'd59321, 16'd64975, 16'd9884, 16'd55510, 16'd4211, 16'd58572});
	test_expansion(128'h301ed8bd5686b607419e889a09a87c1a, {16'd26820, 16'd15309, 16'd53245, 16'd60473, 16'd21909, 16'd50958, 16'd41583, 16'd481, 16'd52480, 16'd62088, 16'd45915, 16'd853, 16'd27390, 16'd56243, 16'd41344, 16'd6225, 16'd19713, 16'd8685, 16'd49559, 16'd24936, 16'd19544, 16'd6290, 16'd18260, 16'd47723, 16'd41637, 16'd58600});
	test_expansion(128'h7709611d1a8d6507c85f17facbcda630, {16'd32199, 16'd15141, 16'd4300, 16'd60653, 16'd35399, 16'd5196, 16'd59758, 16'd56966, 16'd44853, 16'd39511, 16'd65016, 16'd23007, 16'd62146, 16'd37976, 16'd21529, 16'd23759, 16'd13041, 16'd33114, 16'd2711, 16'd61246, 16'd18002, 16'd47550, 16'd44303, 16'd9481, 16'd9302, 16'd23707});
	test_expansion(128'h1cf59356bb37bd5fb399b383eebb6026, {16'd5162, 16'd52212, 16'd1746, 16'd31588, 16'd56589, 16'd40722, 16'd60972, 16'd573, 16'd45565, 16'd46563, 16'd24752, 16'd36501, 16'd29525, 16'd7104, 16'd19670, 16'd7553, 16'd30040, 16'd22181, 16'd42985, 16'd45473, 16'd47120, 16'd31739, 16'd61793, 16'd59654, 16'd64453, 16'd45917});
	test_expansion(128'h29dd078508a3077327177aaee6faedca, {16'd14810, 16'd52889, 16'd7489, 16'd43507, 16'd56693, 16'd11686, 16'd43434, 16'd46400, 16'd49731, 16'd44588, 16'd41306, 16'd24582, 16'd60128, 16'd56942, 16'd49903, 16'd47120, 16'd30486, 16'd57802, 16'd27015, 16'd31053, 16'd27437, 16'd31913, 16'd59283, 16'd37086, 16'd55410, 16'd40044});
	test_expansion(128'h3e7a1820754a9735ca8f0976016f7925, {16'd48401, 16'd34440, 16'd57106, 16'd30881, 16'd18987, 16'd40826, 16'd23297, 16'd4834, 16'd54849, 16'd13210, 16'd27522, 16'd28127, 16'd5918, 16'd3799, 16'd25424, 16'd63629, 16'd65393, 16'd2581, 16'd6221, 16'd11495, 16'd50870, 16'd8521, 16'd28444, 16'd12420, 16'd29789, 16'd23061});
	test_expansion(128'h9f4cee659eeff14693a11a69d7e80692, {16'd51500, 16'd36429, 16'd43378, 16'd26396, 16'd40739, 16'd52135, 16'd64889, 16'd19533, 16'd25805, 16'd17409, 16'd5457, 16'd15929, 16'd42676, 16'd37530, 16'd63522, 16'd27976, 16'd19844, 16'd35056, 16'd36740, 16'd54663, 16'd50447, 16'd10208, 16'd49060, 16'd18754, 16'd42289, 16'd6187});
	test_expansion(128'ha490c49201fefc5a2cd71a2ef4d9db7a, {16'd64856, 16'd57411, 16'd7375, 16'd51804, 16'd9978, 16'd41699, 16'd19237, 16'd58059, 16'd13513, 16'd39866, 16'd39710, 16'd3045, 16'd1639, 16'd64303, 16'd64675, 16'd32694, 16'd57090, 16'd5957, 16'd4470, 16'd36441, 16'd60344, 16'd10080, 16'd15507, 16'd56498, 16'd23672, 16'd44615});
	test_expansion(128'h7eed68d8ddb140968c7bc0ff98bafce1, {16'd45519, 16'd6194, 16'd30739, 16'd8987, 16'd58368, 16'd46214, 16'd40200, 16'd30178, 16'd24331, 16'd64981, 16'd45616, 16'd35199, 16'd54794, 16'd31714, 16'd30808, 16'd50434, 16'd60398, 16'd53041, 16'd3216, 16'd18296, 16'd57077, 16'd49240, 16'd23725, 16'd17341, 16'd60816, 16'd5023});
	test_expansion(128'hec4bccd7ae0a27e7645588178aa8d344, {16'd43395, 16'd7776, 16'd49406, 16'd62325, 16'd57814, 16'd33993, 16'd59360, 16'd17251, 16'd27329, 16'd36566, 16'd11827, 16'd33866, 16'd22421, 16'd37955, 16'd62317, 16'd8268, 16'd46415, 16'd3026, 16'd5335, 16'd2480, 16'd168, 16'd15468, 16'd61894, 16'd22304, 16'd22956, 16'd18335});
	test_expansion(128'h386103a7bd95c7c39c6f5619d3083d03, {16'd26118, 16'd56311, 16'd52153, 16'd21005, 16'd36813, 16'd62896, 16'd440, 16'd17440, 16'd25137, 16'd32239, 16'd51147, 16'd52390, 16'd36445, 16'd39621, 16'd31495, 16'd23820, 16'd43752, 16'd31231, 16'd14888, 16'd63133, 16'd39206, 16'd6804, 16'd59358, 16'd27747, 16'd60175, 16'd58590});
	test_expansion(128'h1fe719bc9dfb8102ae99c456fd40ac21, {16'd50391, 16'd12253, 16'd12512, 16'd48463, 16'd35309, 16'd20470, 16'd11587, 16'd7317, 16'd59886, 16'd3688, 16'd39968, 16'd54141, 16'd13256, 16'd50876, 16'd17083, 16'd49247, 16'd55276, 16'd59552, 16'd52183, 16'd54972, 16'd61938, 16'd41877, 16'd33329, 16'd63049, 16'd56358, 16'd62356});
	test_expansion(128'hce541eb16a375d2feb618d1bfb85a9f1, {16'd14316, 16'd60780, 16'd37520, 16'd118, 16'd29037, 16'd1040, 16'd54521, 16'd19292, 16'd10083, 16'd17031, 16'd64270, 16'd36799, 16'd41143, 16'd37725, 16'd57099, 16'd19356, 16'd21620, 16'd53120, 16'd40925, 16'd12862, 16'd58792, 16'd27657, 16'd47770, 16'd50521, 16'd38748, 16'd65455});
	test_expansion(128'hd2eb8e243f95baa896281a5f1a821ac6, {16'd3010, 16'd60869, 16'd21589, 16'd52772, 16'd35552, 16'd23904, 16'd34679, 16'd39839, 16'd40754, 16'd26749, 16'd26631, 16'd61730, 16'd39250, 16'd63507, 16'd47686, 16'd24024, 16'd53245, 16'd63436, 16'd20742, 16'd2939, 16'd43817, 16'd11447, 16'd1289, 16'd27865, 16'd45335, 16'd44920});
	test_expansion(128'h8f1d79ed78c3013d9606724fade7b4cf, {16'd14720, 16'd15623, 16'd57643, 16'd29454, 16'd18465, 16'd42966, 16'd25484, 16'd48471, 16'd12878, 16'd5874, 16'd41022, 16'd5605, 16'd20017, 16'd14999, 16'd64882, 16'd31794, 16'd44095, 16'd29362, 16'd41145, 16'd14062, 16'd51275, 16'd37349, 16'd59994, 16'd63417, 16'd14273, 16'd50470});
	test_expansion(128'h7cad94946d5fc4936fd6b5298549abf1, {16'd2919, 16'd29744, 16'd15630, 16'd14862, 16'd12584, 16'd59025, 16'd43926, 16'd29699, 16'd16235, 16'd30673, 16'd16088, 16'd58480, 16'd24686, 16'd12041, 16'd57975, 16'd10776, 16'd13887, 16'd4880, 16'd51521, 16'd29609, 16'd63651, 16'd4625, 16'd56163, 16'd53988, 16'd39589, 16'd12978});
	test_expansion(128'h7deb6ab8188682bee52c487884827010, {16'd39608, 16'd38980, 16'd65050, 16'd7113, 16'd54548, 16'd23001, 16'd48244, 16'd64601, 16'd27552, 16'd51675, 16'd43469, 16'd28889, 16'd48481, 16'd53730, 16'd38110, 16'd18226, 16'd24966, 16'd5529, 16'd36287, 16'd27129, 16'd28083, 16'd9183, 16'd55668, 16'd45391, 16'd42760, 16'd31150});
	test_expansion(128'hae8cfec1ab745d257b0b9a0c2eed9f69, {16'd4165, 16'd64392, 16'd18966, 16'd5889, 16'd1712, 16'd8393, 16'd55257, 16'd49786, 16'd16718, 16'd16000, 16'd19026, 16'd36699, 16'd6588, 16'd47685, 16'd47600, 16'd6196, 16'd42788, 16'd9869, 16'd62420, 16'd28697, 16'd28878, 16'd58030, 16'd62372, 16'd22106, 16'd53792, 16'd13389});
	test_expansion(128'he5e0758e7b4634d3cc97b5a4b7cd69ce, {16'd52668, 16'd24195, 16'd12369, 16'd33041, 16'd36568, 16'd39461, 16'd19867, 16'd61405, 16'd13358, 16'd37528, 16'd16182, 16'd6619, 16'd45207, 16'd8517, 16'd9523, 16'd63705, 16'd31151, 16'd25965, 16'd26568, 16'd47268, 16'd59995, 16'd52344, 16'd51963, 16'd40543, 16'd29013, 16'd41688});
	test_expansion(128'h0e64f6dc0db284455471e44229597782, {16'd26135, 16'd12915, 16'd31611, 16'd7573, 16'd7159, 16'd56352, 16'd23884, 16'd4190, 16'd50698, 16'd58188, 16'd12964, 16'd32452, 16'd30011, 16'd60093, 16'd63239, 16'd54118, 16'd511, 16'd56041, 16'd27528, 16'd36375, 16'd50244, 16'd29809, 16'd23382, 16'd2807, 16'd51276, 16'd44038});
	test_expansion(128'h8e361ac8f651f38cf9fe780c88031e70, {16'd12664, 16'd42675, 16'd41070, 16'd47773, 16'd16367, 16'd42469, 16'd1697, 16'd51585, 16'd17113, 16'd64970, 16'd51348, 16'd53874, 16'd5490, 16'd43856, 16'd10249, 16'd46802, 16'd25045, 16'd60081, 16'd53867, 16'd9038, 16'd7125, 16'd47694, 16'd44743, 16'd50603, 16'd47279, 16'd41157});
	test_expansion(128'h7f85086e0bb7bd9f5d47b30e3790f987, {16'd31559, 16'd48708, 16'd59660, 16'd22824, 16'd2683, 16'd9753, 16'd42963, 16'd64070, 16'd33711, 16'd59616, 16'd62654, 16'd52971, 16'd16826, 16'd6390, 16'd33004, 16'd29717, 16'd25085, 16'd43799, 16'd39803, 16'd1344, 16'd48896, 16'd60510, 16'd39876, 16'd58189, 16'd5995, 16'd21344});
	test_expansion(128'h4fb592e9549374368025a20ddca1fb37, {16'd3390, 16'd36764, 16'd21113, 16'd23005, 16'd10800, 16'd60517, 16'd8569, 16'd3506, 16'd26448, 16'd62689, 16'd56890, 16'd48681, 16'd1331, 16'd41230, 16'd34018, 16'd41824, 16'd38948, 16'd51320, 16'd9443, 16'd52791, 16'd7183, 16'd56292, 16'd6146, 16'd52456, 16'd17986, 16'd21015});
	test_expansion(128'h798a9c63f9b3f84574fd4dcc3c501baf, {16'd16235, 16'd5245, 16'd7262, 16'd10607, 16'd11810, 16'd25808, 16'd45957, 16'd58881, 16'd47817, 16'd23382, 16'd31753, 16'd6983, 16'd38593, 16'd19567, 16'd30422, 16'd3163, 16'd60032, 16'd791, 16'd678, 16'd3754, 16'd1320, 16'd18563, 16'd21473, 16'd59852, 16'd11112, 16'd60924});
	test_expansion(128'h1894d792dfeb46875fbe5c368aac442b, {16'd28657, 16'd14715, 16'd20728, 16'd13275, 16'd34171, 16'd9754, 16'd48567, 16'd41403, 16'd2942, 16'd34949, 16'd10552, 16'd15172, 16'd38688, 16'd10936, 16'd26076, 16'd1820, 16'd24464, 16'd1359, 16'd34028, 16'd39150, 16'd11245, 16'd49941, 16'd15888, 16'd59838, 16'd4097, 16'd17234});
	test_expansion(128'h428711ee9bd8b2df90ee5acf7ac21d5e, {16'd16192, 16'd34060, 16'd23760, 16'd63173, 16'd7568, 16'd65022, 16'd58184, 16'd17872, 16'd4352, 16'd45535, 16'd1416, 16'd8965, 16'd61611, 16'd32540, 16'd9170, 16'd13775, 16'd55062, 16'd96, 16'd7663, 16'd37506, 16'd48281, 16'd6179, 16'd46903, 16'd23745, 16'd27078, 16'd23276});
	test_expansion(128'h2ffa4067e20ffd4a1c6090ee735615d8, {16'd51827, 16'd39713, 16'd40145, 16'd17878, 16'd17968, 16'd14416, 16'd37069, 16'd21975, 16'd60006, 16'd61934, 16'd13961, 16'd64860, 16'd57449, 16'd7994, 16'd22325, 16'd10369, 16'd39431, 16'd9644, 16'd5727, 16'd62033, 16'd17901, 16'd51275, 16'd37099, 16'd6157, 16'd37419, 16'd16327});
	test_expansion(128'h6908141b92edce18570a7d2e01720270, {16'd32562, 16'd21389, 16'd62366, 16'd21256, 16'd49375, 16'd30497, 16'd56277, 16'd30832, 16'd57804, 16'd45055, 16'd25878, 16'd38575, 16'd3202, 16'd17656, 16'd46740, 16'd15226, 16'd64225, 16'd26707, 16'd739, 16'd31018, 16'd27476, 16'd31885, 16'd41115, 16'd37608, 16'd10957, 16'd18642});
	test_expansion(128'h2a69706c3f89f8381ed06f4685fc4a6d, {16'd16994, 16'd62128, 16'd23560, 16'd15252, 16'd58599, 16'd25703, 16'd51936, 16'd27272, 16'd27378, 16'd61854, 16'd45755, 16'd30617, 16'd48964, 16'd40188, 16'd36387, 16'd1212, 16'd32372, 16'd13939, 16'd12568, 16'd49639, 16'd55398, 16'd16734, 16'd43427, 16'd58609, 16'd28423, 16'd59220});
	test_expansion(128'h0bd4e7a6cf1ee1aa581106c69ddd11de, {16'd51714, 16'd5532, 16'd34861, 16'd49098, 16'd56925, 16'd22605, 16'd38235, 16'd20155, 16'd47648, 16'd55248, 16'd51840, 16'd4689, 16'd43947, 16'd9263, 16'd25084, 16'd26068, 16'd23780, 16'd21409, 16'd58094, 16'd44821, 16'd21291, 16'd1729, 16'd8473, 16'd45200, 16'd4921, 16'd28356});
	test_expansion(128'h55882ff468a604b306be5c0039ca8e90, {16'd25472, 16'd4094, 16'd28175, 16'd63399, 16'd11494, 16'd16537, 16'd11701, 16'd9288, 16'd31160, 16'd47557, 16'd5415, 16'd74, 16'd30124, 16'd12067, 16'd58958, 16'd55490, 16'd46800, 16'd26870, 16'd38468, 16'd56092, 16'd36376, 16'd10858, 16'd9218, 16'd63575, 16'd59684, 16'd51720});
	test_expansion(128'h7a7f92e4a65ce4147be3db30c56a5629, {16'd26786, 16'd51232, 16'd61958, 16'd47617, 16'd53579, 16'd58079, 16'd9307, 16'd61556, 16'd22553, 16'd36116, 16'd14639, 16'd49422, 16'd52911, 16'd43209, 16'd52455, 16'd51232, 16'd40333, 16'd42836, 16'd46982, 16'd45085, 16'd14635, 16'd49038, 16'd5183, 16'd1205, 16'd29143, 16'd55471});
	test_expansion(128'hc2b03cb52d0da7d70286d1e6d80e39a3, {16'd18660, 16'd18768, 16'd39626, 16'd10272, 16'd24621, 16'd33560, 16'd13652, 16'd65071, 16'd12086, 16'd33693, 16'd29539, 16'd4690, 16'd39964, 16'd31242, 16'd53001, 16'd63623, 16'd64977, 16'd54135, 16'd53403, 16'd30936, 16'd32107, 16'd21412, 16'd44947, 16'd36738, 16'd6529, 16'd18172});
	test_expansion(128'h22e7eb8a91e5655dc18b799c0a4f0d3a, {16'd19347, 16'd19297, 16'd61900, 16'd7545, 16'd47722, 16'd57643, 16'd59337, 16'd39515, 16'd7275, 16'd18294, 16'd40180, 16'd27075, 16'd10180, 16'd26783, 16'd9564, 16'd27338, 16'd2904, 16'd52208, 16'd12257, 16'd36631, 16'd50407, 16'd18158, 16'd27213, 16'd803, 16'd7426, 16'd5131});
	test_expansion(128'hefd5ed0139eac17dfb8a71ac63159136, {16'd24986, 16'd33478, 16'd41409, 16'd25107, 16'd1469, 16'd61897, 16'd20756, 16'd59136, 16'd42899, 16'd31674, 16'd33736, 16'd9329, 16'd19828, 16'd1919, 16'd17689, 16'd13517, 16'd41166, 16'd32152, 16'd62156, 16'd36970, 16'd57848, 16'd19630, 16'd6980, 16'd14292, 16'd33427, 16'd20230});
	test_expansion(128'h85eb5a4d87b9cf683cf97664727b6a57, {16'd38919, 16'd34023, 16'd16108, 16'd40359, 16'd20935, 16'd19654, 16'd60369, 16'd18947, 16'd1452, 16'd1742, 16'd32443, 16'd20839, 16'd29377, 16'd526, 16'd30465, 16'd45715, 16'd23386, 16'd8119, 16'd28513, 16'd21506, 16'd63470, 16'd34749, 16'd26024, 16'd46380, 16'd60908, 16'd29202});
	test_expansion(128'h0ade7d6b9f8d0ea5aa439c6b30294241, {16'd17312, 16'd945, 16'd29302, 16'd34496, 16'd48505, 16'd2597, 16'd1394, 16'd11073, 16'd32797, 16'd2823, 16'd55118, 16'd11284, 16'd38511, 16'd9833, 16'd19427, 16'd57560, 16'd59899, 16'd12939, 16'd8392, 16'd17714, 16'd4605, 16'd64708, 16'd27603, 16'd21534, 16'd26845, 16'd45421});
	test_expansion(128'h6238590c80b1013014d8269d67b58ff8, {16'd29097, 16'd61817, 16'd58425, 16'd7176, 16'd27191, 16'd43768, 16'd3083, 16'd28379, 16'd21954, 16'd31439, 16'd5102, 16'd55426, 16'd63261, 16'd35417, 16'd8229, 16'd3412, 16'd27892, 16'd9484, 16'd15822, 16'd29346, 16'd46117, 16'd15117, 16'd27164, 16'd1886, 16'd19451, 16'd46300});
	test_expansion(128'h216cb3f2160a90ed1fefff58d29c90d9, {16'd48163, 16'd28992, 16'd26554, 16'd28326, 16'd12674, 16'd34122, 16'd56034, 16'd34741, 16'd23249, 16'd62975, 16'd14880, 16'd41786, 16'd37656, 16'd33145, 16'd62290, 16'd45245, 16'd23126, 16'd28701, 16'd30217, 16'd57405, 16'd35585, 16'd3660, 16'd40537, 16'd13341, 16'd41576, 16'd21194});
	test_expansion(128'he0936dac119c68fce0d24c7cc322e563, {16'd50060, 16'd54072, 16'd47615, 16'd31318, 16'd23384, 16'd1382, 16'd32902, 16'd39439, 16'd4032, 16'd22851, 16'd1330, 16'd37592, 16'd44032, 16'd59391, 16'd44117, 16'd36847, 16'd31773, 16'd54769, 16'd41845, 16'd38689, 16'd9177, 16'd33603, 16'd25643, 16'd62962, 16'd23615, 16'd61286});
	test_expansion(128'h9686ad4ae86c3b6f5b69a2c0f9ab049c, {16'd3240, 16'd57893, 16'd27481, 16'd15271, 16'd63858, 16'd11733, 16'd21024, 16'd52499, 16'd16914, 16'd44153, 16'd32057, 16'd39548, 16'd35784, 16'd4830, 16'd13131, 16'd1207, 16'd23271, 16'd64477, 16'd12240, 16'd45851, 16'd65120, 16'd4257, 16'd12791, 16'd2040, 16'd14366, 16'd16745});
	test_expansion(128'h0386dd6f83a1b7337b237d77f3f548ab, {16'd25014, 16'd59636, 16'd20501, 16'd2563, 16'd29144, 16'd41244, 16'd9713, 16'd47737, 16'd33534, 16'd53579, 16'd30063, 16'd4173, 16'd23581, 16'd49301, 16'd51681, 16'd19107, 16'd9210, 16'd17353, 16'd33886, 16'd59380, 16'd53706, 16'd16706, 16'd45899, 16'd55462, 16'd11870, 16'd53928});
	test_expansion(128'hc3f1b6b1fcd419b10d1f3dac35dc9ee8, {16'd42278, 16'd48885, 16'd16215, 16'd51875, 16'd57126, 16'd63734, 16'd48913, 16'd31214, 16'd39787, 16'd39295, 16'd25526, 16'd6258, 16'd19767, 16'd16659, 16'd57522, 16'd15144, 16'd16096, 16'd14554, 16'd45649, 16'd41618, 16'd17855, 16'd16992, 16'd34450, 16'd13550, 16'd4987, 16'd52120});
	test_expansion(128'h571e9770a74eea96e24408b0a1939a5a, {16'd55853, 16'd26717, 16'd12532, 16'd46611, 16'd58598, 16'd55977, 16'd55969, 16'd50787, 16'd5881, 16'd46253, 16'd16007, 16'd42773, 16'd28601, 16'd55084, 16'd32263, 16'd17796, 16'd40539, 16'd10595, 16'd27383, 16'd35993, 16'd62755, 16'd36373, 16'd43079, 16'd63382, 16'd10020, 16'd49686});
	test_expansion(128'h3f3d88d276dee74b4499f9cec4d89fbe, {16'd36945, 16'd50241, 16'd10135, 16'd47762, 16'd52070, 16'd34406, 16'd17997, 16'd11218, 16'd58888, 16'd61136, 16'd15007, 16'd34547, 16'd42390, 16'd17543, 16'd64463, 16'd37391, 16'd4381, 16'd53024, 16'd60820, 16'd33556, 16'd13614, 16'd37907, 16'd5307, 16'd23303, 16'd18687, 16'd51363});
	test_expansion(128'h33bb67089583cad3b70b242a0adcfff9, {16'd7995, 16'd16920, 16'd45055, 16'd43265, 16'd28725, 16'd24333, 16'd41957, 16'd39342, 16'd22485, 16'd9725, 16'd61940, 16'd64769, 16'd18202, 16'd62915, 16'd46792, 16'd59220, 16'd64315, 16'd5651, 16'd11549, 16'd26585, 16'd21544, 16'd23154, 16'd64598, 16'd50311, 16'd62017, 16'd59879});
	test_expansion(128'h09205a056fbf0653364a5a3360e501da, {16'd4278, 16'd31651, 16'd32530, 16'd20032, 16'd33224, 16'd65085, 16'd35033, 16'd37336, 16'd60856, 16'd622, 16'd590, 16'd21934, 16'd768, 16'd37869, 16'd36062, 16'd42427, 16'd44857, 16'd2297, 16'd56580, 16'd43887, 16'd20299, 16'd20633, 16'd9206, 16'd61461, 16'd11647, 16'd44906});
	test_expansion(128'h6a5136ae798a8eb76669ae99bdacf77d, {16'd41522, 16'd19394, 16'd56257, 16'd6423, 16'd36613, 16'd44133, 16'd24340, 16'd64426, 16'd37928, 16'd23191, 16'd17439, 16'd23015, 16'd39291, 16'd25479, 16'd16069, 16'd43929, 16'd48727, 16'd19316, 16'd11581, 16'd4008, 16'd26781, 16'd60101, 16'd6785, 16'd57453, 16'd28850, 16'd36132});
	test_expansion(128'h21fbe08d391075c23496bacee3ded775, {16'd51866, 16'd64280, 16'd64943, 16'd58685, 16'd1444, 16'd41082, 16'd27952, 16'd25786, 16'd1642, 16'd14095, 16'd16359, 16'd21418, 16'd40709, 16'd44426, 16'd2817, 16'd54737, 16'd61885, 16'd18077, 16'd41156, 16'd19262, 16'd13012, 16'd54349, 16'd26221, 16'd23578, 16'd57964, 16'd61521});
	test_expansion(128'h724c3716dabc310a4e9951515230266f, {16'd56831, 16'd52437, 16'd38694, 16'd51682, 16'd22665, 16'd37330, 16'd5597, 16'd63046, 16'd7492, 16'd10183, 16'd53337, 16'd5961, 16'd55458, 16'd9798, 16'd49360, 16'd1951, 16'd1966, 16'd16287, 16'd10945, 16'd35821, 16'd13748, 16'd29170, 16'd30217, 16'd17385, 16'd12753, 16'd34187});
	test_expansion(128'h2a8b2686dc61b2566b4c868e6caa68b5, {16'd53604, 16'd22112, 16'd61191, 16'd34094, 16'd14649, 16'd1938, 16'd31546, 16'd24782, 16'd43581, 16'd17824, 16'd1733, 16'd18334, 16'd43972, 16'd36560, 16'd63798, 16'd7553, 16'd9442, 16'd35415, 16'd1228, 16'd36869, 16'd59087, 16'd49757, 16'd39431, 16'd63469, 16'd11402, 16'd7175});
	test_expansion(128'hb2e76e5bd69e22682b9030f3b03bc336, {16'd8249, 16'd10030, 16'd13550, 16'd12748, 16'd57321, 16'd47962, 16'd49895, 16'd31664, 16'd8943, 16'd53566, 16'd62602, 16'd56470, 16'd39618, 16'd21544, 16'd7042, 16'd51536, 16'd44904, 16'd13786, 16'd52012, 16'd57906, 16'd24329, 16'd64008, 16'd44733, 16'd13474, 16'd24886, 16'd57517});
	test_expansion(128'h3f6c3201e3e56739cdf14236121cf5aa, {16'd25683, 16'd36700, 16'd62615, 16'd12027, 16'd46528, 16'd32818, 16'd5887, 16'd58240, 16'd26701, 16'd4739, 16'd30934, 16'd26792, 16'd48566, 16'd33256, 16'd37721, 16'd2487, 16'd58652, 16'd12311, 16'd45755, 16'd45100, 16'd5611, 16'd26185, 16'd51046, 16'd38716, 16'd12975, 16'd49530});
	test_expansion(128'hd335ec1a866db1d0cd10913cd55da281, {16'd60368, 16'd776, 16'd54283, 16'd7975, 16'd33713, 16'd3054, 16'd62155, 16'd45715, 16'd9624, 16'd9756, 16'd18431, 16'd45723, 16'd3974, 16'd28560, 16'd10531, 16'd52405, 16'd19705, 16'd15476, 16'd33489, 16'd10555, 16'd53470, 16'd49677, 16'd8278, 16'd23212, 16'd7520, 16'd65455});
	test_expansion(128'hadab5ec07ff5d27df0688ba4fb3a311e, {16'd46544, 16'd64570, 16'd60543, 16'd45319, 16'd11272, 16'd48372, 16'd20012, 16'd26548, 16'd64139, 16'd25848, 16'd40299, 16'd39751, 16'd18228, 16'd22791, 16'd33830, 16'd1379, 16'd3989, 16'd37970, 16'd202, 16'd51142, 16'd23464, 16'd56356, 16'd29886, 16'd50813, 16'd51913, 16'd32179});
	test_expansion(128'hd9c3427f568d3dbe73e8c951172c4c95, {16'd31559, 16'd10355, 16'd54389, 16'd43320, 16'd36881, 16'd6990, 16'd26502, 16'd33189, 16'd49628, 16'd25593, 16'd54864, 16'd267, 16'd7845, 16'd62334, 16'd5549, 16'd58422, 16'd26336, 16'd41870, 16'd53052, 16'd7613, 16'd56676, 16'd10731, 16'd921, 16'd55900, 16'd36882, 16'd8534});
	test_expansion(128'h86a04a37543074fe0c348eed33328505, {16'd62019, 16'd39084, 16'd51160, 16'd10873, 16'd43610, 16'd53896, 16'd46593, 16'd3120, 16'd56450, 16'd9444, 16'd51067, 16'd21365, 16'd5685, 16'd63155, 16'd23070, 16'd34851, 16'd37438, 16'd53963, 16'd27522, 16'd35435, 16'd27100, 16'd39477, 16'd38520, 16'd16186, 16'd8301, 16'd37275});
	test_expansion(128'h595b6af4be967230d3f2f31ec09c185b, {16'd55904, 16'd56103, 16'd38114, 16'd19435, 16'd8374, 16'd3253, 16'd58052, 16'd18336, 16'd56901, 16'd36328, 16'd17510, 16'd9069, 16'd26886, 16'd44701, 16'd28721, 16'd49158, 16'd18121, 16'd41190, 16'd15956, 16'd4250, 16'd51966, 16'd42875, 16'd5826, 16'd27502, 16'd53187, 16'd28062});
	test_expansion(128'h5fe4ce3d71aeeebc144c4f9534e7bc4d, {16'd19474, 16'd57910, 16'd56500, 16'd11552, 16'd26442, 16'd51170, 16'd9278, 16'd37583, 16'd3550, 16'd47856, 16'd16642, 16'd26644, 16'd38129, 16'd19448, 16'd21213, 16'd55069, 16'd23237, 16'd63564, 16'd26153, 16'd49051, 16'd13651, 16'd19705, 16'd11902, 16'd35540, 16'd16909, 16'd24600});
	test_expansion(128'h6bfb8daf09844750549a403d2e590507, {16'd30912, 16'd16240, 16'd43443, 16'd58988, 16'd10354, 16'd26819, 16'd1647, 16'd28724, 16'd47272, 16'd44404, 16'd49221, 16'd9983, 16'd8772, 16'd10560, 16'd11656, 16'd5316, 16'd15370, 16'd13237, 16'd20243, 16'd19777, 16'd43977, 16'd6076, 16'd6940, 16'd57760, 16'd16294, 16'd41574});
	test_expansion(128'h8ee7238c08b1282727049f2c8c2b081c, {16'd32214, 16'd53342, 16'd15403, 16'd21044, 16'd39737, 16'd64675, 16'd34921, 16'd1954, 16'd56076, 16'd33169, 16'd57709, 16'd10386, 16'd51548, 16'd62740, 16'd17365, 16'd7916, 16'd7475, 16'd64722, 16'd56270, 16'd1621, 16'd16956, 16'd40689, 16'd8732, 16'd58504, 16'd12243, 16'd22657});
	test_expansion(128'h22648ead8fe0456aab73da9226cd67c2, {16'd61319, 16'd17765, 16'd12757, 16'd59951, 16'd21312, 16'd56379, 16'd11333, 16'd18543, 16'd45941, 16'd3130, 16'd31786, 16'd16830, 16'd391, 16'd59371, 16'd50617, 16'd24944, 16'd32905, 16'd61755, 16'd16382, 16'd51420, 16'd49369, 16'd9450, 16'd5329, 16'd14919, 16'd40908, 16'd48245});
	test_expansion(128'h1de012abcd0c13d2faba98c06af8e5d9, {16'd38435, 16'd14068, 16'd44191, 16'd55590, 16'd23039, 16'd9785, 16'd30988, 16'd1938, 16'd44303, 16'd42731, 16'd44971, 16'd26487, 16'd6115, 16'd7085, 16'd13277, 16'd25283, 16'd4755, 16'd25135, 16'd41240, 16'd11901, 16'd4624, 16'd26958, 16'd44434, 16'd9653, 16'd36430, 16'd11547});
	test_expansion(128'heedb093faff8c735a188b4df71649368, {16'd28141, 16'd41762, 16'd38404, 16'd64649, 16'd55236, 16'd7269, 16'd46494, 16'd48937, 16'd48710, 16'd4882, 16'd65136, 16'd62763, 16'd18201, 16'd23190, 16'd1672, 16'd49126, 16'd33395, 16'd10250, 16'd56266, 16'd33350, 16'd13908, 16'd51723, 16'd47405, 16'd3494, 16'd43055, 16'd25872});
	test_expansion(128'h0bdf34fb21ca32ddee17939f75b29671, {16'd30644, 16'd59170, 16'd48988, 16'd59659, 16'd24979, 16'd30348, 16'd15797, 16'd4658, 16'd47375, 16'd23777, 16'd1381, 16'd30765, 16'd61284, 16'd14218, 16'd50682, 16'd17571, 16'd17793, 16'd52566, 16'd20044, 16'd17252, 16'd30964, 16'd38773, 16'd53891, 16'd30906, 16'd36354, 16'd18994});
	test_expansion(128'hae056f52fab8dccc516f45e132c5d83d, {16'd52635, 16'd21392, 16'd50494, 16'd47045, 16'd63717, 16'd60759, 16'd52516, 16'd33064, 16'd32011, 16'd5789, 16'd31326, 16'd53630, 16'd5863, 16'd59529, 16'd28953, 16'd23152, 16'd16493, 16'd21214, 16'd21217, 16'd58569, 16'd36934, 16'd52461, 16'd8689, 16'd23812, 16'd27423, 16'd61802});
	test_expansion(128'hb74882509a98269f73212f021e879272, {16'd12765, 16'd57448, 16'd64652, 16'd39171, 16'd50211, 16'd59210, 16'd2876, 16'd29385, 16'd61146, 16'd39498, 16'd25913, 16'd4319, 16'd55888, 16'd42390, 16'd58687, 16'd2213, 16'd49247, 16'd21411, 16'd3058, 16'd56872, 16'd24916, 16'd1466, 16'd776, 16'd3851, 16'd51914, 16'd50885});
	test_expansion(128'h8ae0e0dcfe0da975edf9fbf923baecea, {16'd61396, 16'd58889, 16'd43744, 16'd44852, 16'd58237, 16'd10929, 16'd22043, 16'd47388, 16'd8720, 16'd49657, 16'd19636, 16'd36125, 16'd20793, 16'd33397, 16'd51503, 16'd7332, 16'd58322, 16'd49109, 16'd30170, 16'd15399, 16'd64296, 16'd36568, 16'd44006, 16'd7072, 16'd18164, 16'd7941});
	test_expansion(128'h76fc99eb8b1ba9a97b818d792ed4d936, {16'd27377, 16'd30320, 16'd42735, 16'd42433, 16'd1079, 16'd37154, 16'd59362, 16'd45948, 16'd48620, 16'd6345, 16'd47399, 16'd47136, 16'd25707, 16'd56967, 16'd47461, 16'd28876, 16'd1330, 16'd9412, 16'd10488, 16'd1252, 16'd56845, 16'd25356, 16'd30494, 16'd20011, 16'd9214, 16'd14687});
	test_expansion(128'h9a45088da1abb5130b8e515ae34cc823, {16'd62049, 16'd48320, 16'd37140, 16'd11903, 16'd24156, 16'd62134, 16'd22272, 16'd62052, 16'd4878, 16'd12512, 16'd29808, 16'd59331, 16'd40283, 16'd5701, 16'd10552, 16'd10730, 16'd45230, 16'd50467, 16'd17595, 16'd20824, 16'd61146, 16'd53074, 16'd26184, 16'd36277, 16'd58237, 16'd14897});
	test_expansion(128'hea337fa15a23c91f0decbb88636437ca, {16'd21066, 16'd54611, 16'd53899, 16'd57159, 16'd19193, 16'd6925, 16'd58207, 16'd4092, 16'd57187, 16'd8481, 16'd45082, 16'd12261, 16'd61026, 16'd60319, 16'd25839, 16'd30225, 16'd65372, 16'd11358, 16'd13930, 16'd12421, 16'd16483, 16'd60573, 16'd64833, 16'd59646, 16'd46623, 16'd19045});
	test_expansion(128'ha739f3f8250de74a82cde8fb6cec3595, {16'd52831, 16'd22740, 16'd19084, 16'd2853, 16'd14719, 16'd35290, 16'd30893, 16'd30737, 16'd56285, 16'd34154, 16'd63124, 16'd12832, 16'd7032, 16'd5700, 16'd24185, 16'd36030, 16'd9950, 16'd33265, 16'd3301, 16'd23789, 16'd20637, 16'd13550, 16'd56772, 16'd51588, 16'd52741, 16'd27560});
	test_expansion(128'hc9cf7a53ead63fdcdd3e3a9fa480b411, {16'd3339, 16'd49213, 16'd63902, 16'd50448, 16'd498, 16'd9342, 16'd53883, 16'd49669, 16'd36847, 16'd32982, 16'd6272, 16'd10827, 16'd54018, 16'd53463, 16'd30062, 16'd1618, 16'd25999, 16'd49853, 16'd4809, 16'd29743, 16'd53486, 16'd32486, 16'd61982, 16'd35516, 16'd61706, 16'd37799});
	test_expansion(128'h67c87bc4a2e42584392761a010db58e7, {16'd47767, 16'd19004, 16'd61041, 16'd43271, 16'd44225, 16'd30228, 16'd61054, 16'd65062, 16'd18689, 16'd7907, 16'd60457, 16'd55615, 16'd54143, 16'd12021, 16'd36546, 16'd55726, 16'd29804, 16'd20792, 16'd34383, 16'd11478, 16'd23863, 16'd5150, 16'd48499, 16'd25607, 16'd28937, 16'd11047});
	test_expansion(128'h10298b470baf11633482a532684abfe2, {16'd33467, 16'd38910, 16'd5232, 16'd23938, 16'd312, 16'd58208, 16'd45132, 16'd21551, 16'd30893, 16'd15062, 16'd65206, 16'd62674, 16'd36669, 16'd30750, 16'd46173, 16'd2141, 16'd39144, 16'd9209, 16'd37897, 16'd36176, 16'd47418, 16'd61114, 16'd7730, 16'd8979, 16'd62016, 16'd14015});
	test_expansion(128'h33940059688dde6d6b8d0280d1367af5, {16'd39204, 16'd37277, 16'd23357, 16'd30670, 16'd25364, 16'd61999, 16'd35133, 16'd18964, 16'd20698, 16'd44253, 16'd10468, 16'd32282, 16'd20088, 16'd48646, 16'd63552, 16'd25678, 16'd55872, 16'd28244, 16'd17721, 16'd11587, 16'd7068, 16'd56851, 16'd61361, 16'd41500, 16'd4103, 16'd18770});
	test_expansion(128'hff37d60585b3c8931866b80d9e701af4, {16'd54109, 16'd9608, 16'd6780, 16'd89, 16'd48472, 16'd6834, 16'd7828, 16'd332, 16'd46475, 16'd30603, 16'd37301, 16'd22280, 16'd37917, 16'd28514, 16'd30791, 16'd52006, 16'd30565, 16'd9757, 16'd42255, 16'd53858, 16'd34075, 16'd50702, 16'd24171, 16'd16852, 16'd41390, 16'd21849});
	test_expansion(128'hf01dd229d4f389876455c7e973ae4ce2, {16'd31259, 16'd64124, 16'd9810, 16'd9827, 16'd10027, 16'd29718, 16'd5143, 16'd8015, 16'd56149, 16'd45185, 16'd41932, 16'd18367, 16'd26973, 16'd21468, 16'd7675, 16'd13394, 16'd7171, 16'd14652, 16'd42678, 16'd29068, 16'd11569, 16'd22847, 16'd472, 16'd20716, 16'd9827, 16'd50227});
	test_expansion(128'h9a1ea7dfe2880712c07622cc2a08bb4b, {16'd25951, 16'd17073, 16'd30698, 16'd1247, 16'd62285, 16'd4603, 16'd21397, 16'd29008, 16'd58528, 16'd24096, 16'd23656, 16'd16056, 16'd57676, 16'd33028, 16'd39213, 16'd62525, 16'd37242, 16'd35139, 16'd12282, 16'd5477, 16'd53213, 16'd9403, 16'd25270, 16'd10676, 16'd12300, 16'd59005});
	test_expansion(128'hbbb7fc3d26328c2f0a39216928e8b45e, {16'd11148, 16'd19809, 16'd56874, 16'd53736, 16'd56054, 16'd41610, 16'd9374, 16'd33997, 16'd28310, 16'd37069, 16'd35965, 16'd48922, 16'd64325, 16'd21065, 16'd40751, 16'd49959, 16'd45078, 16'd5627, 16'd15343, 16'd19124, 16'd16508, 16'd29986, 16'd60556, 16'd53057, 16'd60492, 16'd54629});
	test_expansion(128'h521cf5e3d923fd760e3e9353ca139a5e, {16'd27480, 16'd55498, 16'd13778, 16'd40555, 16'd6276, 16'd22977, 16'd61957, 16'd19546, 16'd15034, 16'd8568, 16'd25312, 16'd33492, 16'd14241, 16'd20410, 16'd11365, 16'd62010, 16'd23140, 16'd60782, 16'd21995, 16'd22128, 16'd46013, 16'd55946, 16'd33429, 16'd50945, 16'd56287, 16'd24759});
	test_expansion(128'h291174c2458d70492fe1fdc02404c8b9, {16'd24809, 16'd17164, 16'd54671, 16'd17409, 16'd40518, 16'd30493, 16'd54052, 16'd10092, 16'd44887, 16'd1090, 16'd18421, 16'd34732, 16'd16960, 16'd27066, 16'd42802, 16'd52358, 16'd44557, 16'd20569, 16'd135, 16'd4650, 16'd52309, 16'd15335, 16'd54765, 16'd4152, 16'd64000, 16'd22339});
	test_expansion(128'hce2cb17a883f23c47fd57808b2f8d9cd, {16'd795, 16'd29604, 16'd59840, 16'd53736, 16'd20465, 16'd16649, 16'd26720, 16'd25655, 16'd17035, 16'd33292, 16'd4673, 16'd51949, 16'd50032, 16'd2366, 16'd30573, 16'd23165, 16'd18445, 16'd50163, 16'd49373, 16'd7635, 16'd15269, 16'd15944, 16'd26432, 16'd34241, 16'd55367, 16'd24897});
	test_expansion(128'h925b004da93e07fa050afd4d40465c80, {16'd21477, 16'd16500, 16'd8111, 16'd8182, 16'd38805, 16'd1059, 16'd4759, 16'd54618, 16'd23173, 16'd12033, 16'd32103, 16'd41694, 16'd56980, 16'd11177, 16'd10679, 16'd3894, 16'd61689, 16'd62352, 16'd13069, 16'd8772, 16'd65106, 16'd17533, 16'd30080, 16'd58051, 16'd64536, 16'd64563});
	test_expansion(128'h4ea1a4a233f7168ee375b6f91293744b, {16'd51656, 16'd34080, 16'd13709, 16'd19331, 16'd43261, 16'd41699, 16'd58775, 16'd7091, 16'd15985, 16'd56103, 16'd11028, 16'd51124, 16'd43113, 16'd43363, 16'd10396, 16'd11935, 16'd33315, 16'd40841, 16'd24147, 16'd64213, 16'd55268, 16'd6064, 16'd1335, 16'd4628, 16'd63888, 16'd60860});
	test_expansion(128'h8f03cbf1c381b2a05b4f433a8b17605d, {16'd25834, 16'd62984, 16'd34503, 16'd21375, 16'd54078, 16'd20432, 16'd20743, 16'd3239, 16'd25742, 16'd4727, 16'd17902, 16'd5502, 16'd14781, 16'd31597, 16'd10493, 16'd16842, 16'd61506, 16'd15516, 16'd46640, 16'd11907, 16'd3682, 16'd37393, 16'd29962, 16'd8530, 16'd31498, 16'd15279});
	test_expansion(128'hced548fde37188bc628d4d4f793f95a0, {16'd3848, 16'd44365, 16'd39288, 16'd5475, 16'd22937, 16'd30253, 16'd24087, 16'd56689, 16'd17350, 16'd48631, 16'd31057, 16'd35503, 16'd52602, 16'd2681, 16'd50647, 16'd64349, 16'd907, 16'd27600, 16'd35194, 16'd61601, 16'd61346, 16'd45330, 16'd10706, 16'd25120, 16'd10215, 16'd10910});
	test_expansion(128'h0ff000f73fc691002f6699067b734d19, {16'd50477, 16'd14730, 16'd38751, 16'd39133, 16'd41364, 16'd28793, 16'd8759, 16'd30686, 16'd7766, 16'd48054, 16'd38933, 16'd64754, 16'd10489, 16'd34237, 16'd37582, 16'd64606, 16'd29896, 16'd2375, 16'd60292, 16'd7175, 16'd6964, 16'd15185, 16'd13378, 16'd35116, 16'd18836, 16'd5266});
	test_expansion(128'h525e6792201f055b223cdfe0d9522b4b, {16'd1085, 16'd15107, 16'd3928, 16'd39026, 16'd38637, 16'd15703, 16'd55673, 16'd38770, 16'd62155, 16'd21997, 16'd5096, 16'd28866, 16'd9106, 16'd9179, 16'd56943, 16'd15504, 16'd28611, 16'd48584, 16'd8772, 16'd3620, 16'd9942, 16'd20436, 16'd14818, 16'd60460, 16'd43615, 16'd22609});
	test_expansion(128'h7323b526a33b36c73d2e1e02c37a3589, {16'd49148, 16'd497, 16'd18493, 16'd17783, 16'd45754, 16'd16169, 16'd34679, 16'd18867, 16'd45258, 16'd59873, 16'd11046, 16'd11969, 16'd27668, 16'd32147, 16'd32310, 16'd61048, 16'd62749, 16'd20287, 16'd30524, 16'd12612, 16'd60126, 16'd16069, 16'd48195, 16'd43663, 16'd25729, 16'd8433});
	test_expansion(128'hbb17d134a3884a300099ff8a88b42ae9, {16'd62280, 16'd42251, 16'd7426, 16'd11465, 16'd24742, 16'd28040, 16'd55225, 16'd33427, 16'd20260, 16'd40349, 16'd25364, 16'd38691, 16'd48223, 16'd16380, 16'd3336, 16'd61581, 16'd53860, 16'd43729, 16'd25099, 16'd57136, 16'd49565, 16'd33444, 16'd15635, 16'd18513, 16'd18136, 16'd6145});
	test_expansion(128'h8509af111d4ae0fac5080e26df205e76, {16'd55174, 16'd5790, 16'd31548, 16'd1827, 16'd38966, 16'd60775, 16'd52363, 16'd40919, 16'd11676, 16'd16566, 16'd37539, 16'd63742, 16'd39840, 16'd29941, 16'd6456, 16'd23936, 16'd12058, 16'd23859, 16'd28228, 16'd64575, 16'd61107, 16'd24791, 16'd4360, 16'd26158, 16'd56802, 16'd36892});
	test_expansion(128'h5ed2c3de4b79b119c78b521d478f8791, {16'd28382, 16'd29773, 16'd31204, 16'd1817, 16'd15462, 16'd10653, 16'd13041, 16'd4701, 16'd2495, 16'd20750, 16'd4261, 16'd26694, 16'd27247, 16'd64453, 16'd43031, 16'd65291, 16'd12066, 16'd44507, 16'd9246, 16'd27042, 16'd16932, 16'd27404, 16'd34258, 16'd61285, 16'd31987, 16'd9383});
	test_expansion(128'h4df97b7a12bde0f6ccb46b96d0bd5fa9, {16'd34574, 16'd11408, 16'd39931, 16'd38957, 16'd52045, 16'd22398, 16'd1237, 16'd16546, 16'd15771, 16'd21536, 16'd54922, 16'd48301, 16'd36313, 16'd3380, 16'd22251, 16'd16535, 16'd46725, 16'd13093, 16'd33682, 16'd806, 16'd24530, 16'd45969, 16'd47470, 16'd48871, 16'd32778, 16'd4729});
	test_expansion(128'h7aa9371a2072067bdd076313aa418e66, {16'd10628, 16'd55714, 16'd57053, 16'd33268, 16'd28179, 16'd51633, 16'd63968, 16'd13297, 16'd57177, 16'd35623, 16'd20925, 16'd10215, 16'd35496, 16'd11757, 16'd42992, 16'd43151, 16'd50317, 16'd29629, 16'd47881, 16'd9740, 16'd20586, 16'd65509, 16'd48989, 16'd40629, 16'd19427, 16'd19659});
	test_expansion(128'h77536e3e9c912efec0e32e82c9f36191, {16'd30135, 16'd51135, 16'd23247, 16'd47442, 16'd45672, 16'd11285, 16'd41078, 16'd6763, 16'd38035, 16'd6029, 16'd2121, 16'd63227, 16'd706, 16'd33825, 16'd56018, 16'd30596, 16'd45092, 16'd23900, 16'd22915, 16'd8936, 16'd40503, 16'd11125, 16'd48594, 16'd50232, 16'd22339, 16'd15162});
	test_expansion(128'h60542ad9aaf12a371e22bea2a376a542, {16'd11222, 16'd32726, 16'd6600, 16'd9427, 16'd55162, 16'd65478, 16'd27964, 16'd20866, 16'd36099, 16'd28789, 16'd65002, 16'd24822, 16'd26413, 16'd58256, 16'd50829, 16'd36279, 16'd28520, 16'd3159, 16'd24418, 16'd10199, 16'd61750, 16'd32719, 16'd21773, 16'd32904, 16'd61719, 16'd7415});
	test_expansion(128'hd9b1999a3a6ae442dc273825910695a4, {16'd10497, 16'd46166, 16'd22837, 16'd49738, 16'd53472, 16'd5944, 16'd3633, 16'd14490, 16'd22571, 16'd37683, 16'd51182, 16'd35552, 16'd39219, 16'd6983, 16'd62752, 16'd63985, 16'd6891, 16'd28965, 16'd16245, 16'd58344, 16'd64498, 16'd22810, 16'd14815, 16'd46759, 16'd10733, 16'd30267});
	test_expansion(128'ha39384c8a81a21c63af24c5dd53bedbd, {16'd57364, 16'd10026, 16'd24059, 16'd9273, 16'd9637, 16'd1557, 16'd43785, 16'd49852, 16'd24322, 16'd17000, 16'd25971, 16'd61660, 16'd52578, 16'd4143, 16'd32951, 16'd47653, 16'd24938, 16'd43996, 16'd44520, 16'd32319, 16'd24150, 16'd39378, 16'd20537, 16'd64945, 16'd47758, 16'd26318});
	test_expansion(128'h6cc446c9a2fe003a08d08768d8a30624, {16'd34915, 16'd46856, 16'd47040, 16'd35725, 16'd63877, 16'd22841, 16'd6812, 16'd62717, 16'd24782, 16'd29087, 16'd32242, 16'd44974, 16'd50734, 16'd41192, 16'd53262, 16'd36055, 16'd12305, 16'd54594, 16'd50072, 16'd48238, 16'd18782, 16'd63221, 16'd51792, 16'd50874, 16'd12311, 16'd43417});
	test_expansion(128'h8ac07f08699e26a828d6b5da29f47cb1, {16'd54864, 16'd38031, 16'd9378, 16'd53927, 16'd50046, 16'd27322, 16'd364, 16'd36791, 16'd33524, 16'd11132, 16'd5952, 16'd12058, 16'd28049, 16'd16820, 16'd57758, 16'd39712, 16'd36538, 16'd590, 16'd33047, 16'd31724, 16'd28451, 16'd17338, 16'd39038, 16'd35759, 16'd1990, 16'd5458});
	test_expansion(128'hab0b7cd9326b563021251434de91c917, {16'd55720, 16'd29758, 16'd59017, 16'd57289, 16'd3371, 16'd61598, 16'd64294, 16'd2568, 16'd46290, 16'd13333, 16'd30369, 16'd20168, 16'd45939, 16'd5619, 16'd36190, 16'd45829, 16'd53214, 16'd39082, 16'd10864, 16'd22653, 16'd7372, 16'd56228, 16'd51151, 16'd17087, 16'd45670, 16'd2591});
	test_expansion(128'h1519ea005133836f5112d9a41e59924e, {16'd64860, 16'd59333, 16'd44680, 16'd1785, 16'd43376, 16'd3686, 16'd16976, 16'd39818, 16'd35837, 16'd35051, 16'd10032, 16'd19787, 16'd26457, 16'd53288, 16'd37385, 16'd34970, 16'd37091, 16'd7588, 16'd63061, 16'd32732, 16'd2755, 16'd33891, 16'd54123, 16'd50844, 16'd38657, 16'd26179});
	test_expansion(128'h8ed687263266cd1b4fed9fa41d9892b6, {16'd63265, 16'd17020, 16'd26892, 16'd10294, 16'd28768, 16'd58097, 16'd43935, 16'd4016, 16'd10253, 16'd57173, 16'd41437, 16'd34660, 16'd39675, 16'd54453, 16'd15382, 16'd33945, 16'd55287, 16'd27755, 16'd6421, 16'd19668, 16'd24796, 16'd61034, 16'd5573, 16'd62448, 16'd55528, 16'd65250});
	test_expansion(128'h85109fac0966b3a3b43f6a0783b1adeb, {16'd29787, 16'd39480, 16'd16741, 16'd4205, 16'd25059, 16'd48402, 16'd32726, 16'd62082, 16'd53447, 16'd62483, 16'd5098, 16'd56257, 16'd20928, 16'd33114, 16'd1994, 16'd51128, 16'd39599, 16'd28353, 16'd18216, 16'd4316, 16'd11657, 16'd296, 16'd27643, 16'd24609, 16'd53916, 16'd44916});
	test_expansion(128'h05d3d0f8821763397dcd3a9b6e2d07e3, {16'd6746, 16'd16863, 16'd65525, 16'd13618, 16'd30128, 16'd39150, 16'd60215, 16'd48990, 16'd29873, 16'd47200, 16'd17011, 16'd10960, 16'd11244, 16'd33796, 16'd35346, 16'd31546, 16'd59390, 16'd7565, 16'd52260, 16'd19687, 16'd2863, 16'd2544, 16'd8694, 16'd35995, 16'd54411, 16'd65292});
	test_expansion(128'h87b1042851b711cf0a17f33d7f889056, {16'd22499, 16'd55248, 16'd39491, 16'd10888, 16'd32646, 16'd50663, 16'd13191, 16'd698, 16'd22921, 16'd41859, 16'd17652, 16'd18418, 16'd2390, 16'd7170, 16'd9326, 16'd59526, 16'd39021, 16'd10354, 16'd43086, 16'd4511, 16'd35652, 16'd35910, 16'd60359, 16'd25001, 16'd11015, 16'd63991});
	test_expansion(128'hfe0346ce4686e3a31e06dcf192a83097, {16'd25088, 16'd5942, 16'd20634, 16'd46270, 16'd791, 16'd10944, 16'd34649, 16'd6906, 16'd30933, 16'd41940, 16'd31789, 16'd53836, 16'd28836, 16'd55567, 16'd64188, 16'd18863, 16'd58155, 16'd54800, 16'd53145, 16'd58406, 16'd10379, 16'd58733, 16'd17397, 16'd19731, 16'd30240, 16'd31718});
	test_expansion(128'hd586a791538d54ab32cc86a479d9f2a1, {16'd23854, 16'd64987, 16'd58922, 16'd38540, 16'd37492, 16'd48014, 16'd17091, 16'd52121, 16'd43363, 16'd64171, 16'd17339, 16'd16969, 16'd30034, 16'd31091, 16'd26899, 16'd5068, 16'd60167, 16'd45962, 16'd50417, 16'd62935, 16'd45986, 16'd42615, 16'd30911, 16'd32291, 16'd29519, 16'd44782});
	test_expansion(128'h6f3ecc818a54ca05c59d2872fc56f26a, {16'd29692, 16'd63114, 16'd36332, 16'd16211, 16'd60132, 16'd630, 16'd50097, 16'd57687, 16'd13832, 16'd51682, 16'd3798, 16'd50499, 16'd39374, 16'd21164, 16'd7894, 16'd61574, 16'd28529, 16'd29583, 16'd51127, 16'd20840, 16'd34261, 16'd2092, 16'd49936, 16'd7668, 16'd24726, 16'd54238});
	test_expansion(128'hd9910fd0c2f434dd7c88b30f85e6c0e2, {16'd64061, 16'd22370, 16'd37245, 16'd54374, 16'd43767, 16'd35694, 16'd16366, 16'd28850, 16'd47285, 16'd62268, 16'd47140, 16'd42932, 16'd31826, 16'd51772, 16'd8854, 16'd16039, 16'd45002, 16'd12679, 16'd15413, 16'd39567, 16'd44280, 16'd46300, 16'd23684, 16'd672, 16'd27606, 16'd46828});
	test_expansion(128'hc526af426b608a6159d355f6a347c4c0, {16'd60236, 16'd43418, 16'd57332, 16'd16514, 16'd75, 16'd3428, 16'd38729, 16'd21238, 16'd43451, 16'd12722, 16'd56451, 16'd41337, 16'd60265, 16'd13413, 16'd11806, 16'd8236, 16'd11642, 16'd38476, 16'd31047, 16'd44021, 16'd55468, 16'd34829, 16'd55726, 16'd49469, 16'd33542, 16'd40428});
	test_expansion(128'h467c3478b88518dc4829b0e1e406f8e0, {16'd12038, 16'd52542, 16'd57747, 16'd54519, 16'd25885, 16'd24947, 16'd26149, 16'd64577, 16'd6024, 16'd27389, 16'd41945, 16'd19318, 16'd42200, 16'd61027, 16'd27812, 16'd19689, 16'd57255, 16'd52433, 16'd36205, 16'd53864, 16'd62428, 16'd29865, 16'd29607, 16'd61270, 16'd34934, 16'd12364});
	test_expansion(128'ha36b82bb3dcc4ea2e6d7abda3b155810, {16'd50603, 16'd55929, 16'd37517, 16'd35634, 16'd15181, 16'd62742, 16'd55518, 16'd2487, 16'd54489, 16'd32805, 16'd39117, 16'd10181, 16'd29699, 16'd59897, 16'd28648, 16'd42171, 16'd54990, 16'd17152, 16'd17060, 16'd41401, 16'd27, 16'd15195, 16'd49147, 16'd64371, 16'd10724, 16'd20033});
	test_expansion(128'hea5ca1b454de391ef8fb6b024653f3ca, {16'd17597, 16'd45393, 16'd22472, 16'd22151, 16'd35908, 16'd21351, 16'd21137, 16'd47952, 16'd21093, 16'd58505, 16'd18736, 16'd22031, 16'd16619, 16'd42105, 16'd41909, 16'd16711, 16'd8127, 16'd56418, 16'd8847, 16'd33847, 16'd49223, 16'd5444, 16'd123, 16'd23891, 16'd63961, 16'd50971});
	test_expansion(128'hc7ff8117e69c3935f1ac875fe6e2eb85, {16'd12415, 16'd38005, 16'd47136, 16'd63987, 16'd4033, 16'd12437, 16'd28301, 16'd44575, 16'd44422, 16'd25919, 16'd11105, 16'd53268, 16'd8301, 16'd33033, 16'd21099, 16'd14835, 16'd43497, 16'd25745, 16'd43865, 16'd1449, 16'd17514, 16'd50686, 16'd39175, 16'd19945, 16'd33691, 16'd4551});
	test_expansion(128'h202f7aa172b63e6b5675eaf327014638, {16'd11323, 16'd33443, 16'd13792, 16'd49978, 16'd24042, 16'd29060, 16'd59735, 16'd50384, 16'd9148, 16'd22696, 16'd46884, 16'd16903, 16'd32950, 16'd20856, 16'd49827, 16'd52229, 16'd22193, 16'd46764, 16'd22545, 16'd6760, 16'd13498, 16'd41607, 16'd35812, 16'd62255, 16'd10538, 16'd52572});
	test_expansion(128'hf631ddaebb65519cfe48c776e83ba692, {16'd17008, 16'd16697, 16'd44745, 16'd8073, 16'd38945, 16'd40242, 16'd13033, 16'd62700, 16'd42404, 16'd41790, 16'd49283, 16'd40080, 16'd44801, 16'd32016, 16'd64186, 16'd13252, 16'd38414, 16'd41735, 16'd8458, 16'd34587, 16'd331, 16'd58702, 16'd59062, 16'd15570, 16'd47371, 16'd17994});
	test_expansion(128'h4024ce9528e936f097b0ea540961f7b2, {16'd59289, 16'd47589, 16'd55729, 16'd27089, 16'd57861, 16'd22762, 16'd21522, 16'd9134, 16'd32487, 16'd15502, 16'd24851, 16'd53661, 16'd52471, 16'd14609, 16'd13597, 16'd61107, 16'd17548, 16'd17558, 16'd13920, 16'd4432, 16'd26223, 16'd14400, 16'd21907, 16'd46942, 16'd29580, 16'd61959});
	test_expansion(128'hcbbf3a7fb803029a178535f49a742911, {16'd42344, 16'd35969, 16'd9910, 16'd19697, 16'd13130, 16'd57210, 16'd51029, 16'd36668, 16'd3114, 16'd28691, 16'd34477, 16'd25685, 16'd49527, 16'd27821, 16'd47162, 16'd60170, 16'd9281, 16'd2351, 16'd15182, 16'd53832, 16'd20818, 16'd19096, 16'd24047, 16'd35454, 16'd42830, 16'd33262});
	test_expansion(128'he58edad27cc2878403741883a7ceb28d, {16'd10220, 16'd33159, 16'd20951, 16'd31693, 16'd6296, 16'd38223, 16'd53620, 16'd60106, 16'd35282, 16'd33601, 16'd7831, 16'd33681, 16'd20737, 16'd215, 16'd35817, 16'd5871, 16'd13373, 16'd49650, 16'd44639, 16'd35070, 16'd4593, 16'd52192, 16'd17170, 16'd63825, 16'd54981, 16'd8396});
	test_expansion(128'h1c595684ba4bf6a86f120fbc62203de2, {16'd2858, 16'd5936, 16'd48374, 16'd6520, 16'd4385, 16'd54661, 16'd32101, 16'd56923, 16'd56876, 16'd26896, 16'd51760, 16'd31417, 16'd21401, 16'd12121, 16'd26042, 16'd34768, 16'd18953, 16'd989, 16'd41266, 16'd47573, 16'd11297, 16'd18887, 16'd64282, 16'd38818, 16'd27869, 16'd56621});
	test_expansion(128'hb4383754a1286499c8583ea6fbe29d7c, {16'd40293, 16'd49177, 16'd43115, 16'd27517, 16'd1602, 16'd40613, 16'd12961, 16'd56940, 16'd30196, 16'd8822, 16'd11099, 16'd61289, 16'd161, 16'd14492, 16'd52906, 16'd46360, 16'd50083, 16'd48067, 16'd56189, 16'd49128, 16'd18818, 16'd49261, 16'd18083, 16'd16446, 16'd2679, 16'd18430});
	test_expansion(128'he88024dbf278eb6cad69a610c9165bdb, {16'd55879, 16'd44471, 16'd54428, 16'd62506, 16'd2957, 16'd56285, 16'd64530, 16'd4856, 16'd57363, 16'd27032, 16'd63458, 16'd12017, 16'd49815, 16'd20461, 16'd2147, 16'd48695, 16'd28628, 16'd48348, 16'd11959, 16'd15559, 16'd60335, 16'd65478, 16'd43816, 16'd52021, 16'd43896, 16'd23399});
	test_expansion(128'hb7933673a7559e781121f4294d273be3, {16'd45874, 16'd14529, 16'd12950, 16'd6741, 16'd62367, 16'd61260, 16'd51012, 16'd30444, 16'd8547, 16'd7045, 16'd38870, 16'd32207, 16'd53834, 16'd46470, 16'd29936, 16'd22900, 16'd19518, 16'd36475, 16'd52823, 16'd9422, 16'd13471, 16'd49831, 16'd52366, 16'd21801, 16'd32307, 16'd55796});
	test_expansion(128'h536fe5694fe09271fb08fc31c96a7292, {16'd6726, 16'd60686, 16'd29415, 16'd28123, 16'd56061, 16'd14292, 16'd19333, 16'd55528, 16'd27898, 16'd19844, 16'd19082, 16'd50627, 16'd21686, 16'd37741, 16'd17857, 16'd22557, 16'd32162, 16'd25007, 16'd39131, 16'd25824, 16'd61072, 16'd6103, 16'd28091, 16'd29270, 16'd20195, 16'd6878});
	test_expansion(128'h65accb0d86bc31ca37d6993d009e93ae, {16'd54020, 16'd41349, 16'd42002, 16'd61422, 16'd36541, 16'd37145, 16'd46660, 16'd4727, 16'd44720, 16'd48091, 16'd64944, 16'd62921, 16'd44958, 16'd4222, 16'd38157, 16'd3535, 16'd45011, 16'd31241, 16'd10182, 16'd19482, 16'd14858, 16'd47912, 16'd3681, 16'd42340, 16'd44503, 16'd32112});
	test_expansion(128'hfead37404e77448406031112c3837a87, {16'd62571, 16'd20622, 16'd53047, 16'd51454, 16'd19960, 16'd51026, 16'd19333, 16'd11655, 16'd44235, 16'd42131, 16'd45919, 16'd54138, 16'd40240, 16'd10921, 16'd10015, 16'd61927, 16'd8151, 16'd4400, 16'd41941, 16'd13543, 16'd48864, 16'd9629, 16'd46030, 16'd57008, 16'd39337, 16'd8530});
	test_expansion(128'h7f144e75c4c7677493be5c60c2d38ec7, {16'd38137, 16'd29706, 16'd51415, 16'd7024, 16'd20686, 16'd49310, 16'd26386, 16'd3476, 16'd33538, 16'd44555, 16'd48891, 16'd16512, 16'd59891, 16'd56308, 16'd23341, 16'd42444, 16'd18782, 16'd209, 16'd56433, 16'd44764, 16'd14804, 16'd63515, 16'd1691, 16'd5324, 16'd46660, 16'd50317});
	test_expansion(128'h1ceae82958281b4315241095b31422aa, {16'd40806, 16'd7885, 16'd34157, 16'd53331, 16'd37361, 16'd25971, 16'd50926, 16'd31387, 16'd15254, 16'd16518, 16'd6119, 16'd5703, 16'd33895, 16'd14761, 16'd14720, 16'd13142, 16'd58445, 16'd42059, 16'd2875, 16'd5070, 16'd37591, 16'd40973, 16'd17524, 16'd35020, 16'd44650, 16'd46201});
	test_expansion(128'ha5cb7cc6f1e49b35594a9fce84aca7e8, {16'd7214, 16'd59802, 16'd30020, 16'd54926, 16'd59214, 16'd48833, 16'd6325, 16'd31348, 16'd2558, 16'd19464, 16'd26765, 16'd405, 16'd58326, 16'd24327, 16'd6957, 16'd65263, 16'd45151, 16'd59366, 16'd51732, 16'd2773, 16'd30541, 16'd52584, 16'd37078, 16'd13468, 16'd33283, 16'd18697});
	test_expansion(128'h30cc13062948b447768e8e35f81e9fcc, {16'd47655, 16'd5804, 16'd65534, 16'd4473, 16'd39829, 16'd20498, 16'd35434, 16'd63037, 16'd60953, 16'd24714, 16'd14014, 16'd64702, 16'd25806, 16'd11524, 16'd27656, 16'd35379, 16'd57855, 16'd52392, 16'd64891, 16'd38552, 16'd15340, 16'd60630, 16'd6695, 16'd50749, 16'd27499, 16'd17251});
	test_expansion(128'h9636d0497c89ea3315f378e9de988396, {16'd40843, 16'd56968, 16'd9116, 16'd14895, 16'd56271, 16'd3025, 16'd46627, 16'd6378, 16'd3318, 16'd36290, 16'd11249, 16'd51265, 16'd2582, 16'd39525, 16'd9503, 16'd42720, 16'd35551, 16'd8502, 16'd31221, 16'd34643, 16'd5797, 16'd22856, 16'd21136, 16'd58474, 16'd39616, 16'd33979});
	test_expansion(128'h996ea255af90257ec253aab7ab85671e, {16'd62052, 16'd42, 16'd33299, 16'd43179, 16'd65306, 16'd29316, 16'd19454, 16'd25555, 16'd41807, 16'd31443, 16'd25981, 16'd1918, 16'd44970, 16'd3382, 16'd46141, 16'd15306, 16'd55184, 16'd30919, 16'd6829, 16'd21234, 16'd42920, 16'd18355, 16'd24465, 16'd61191, 16'd59083, 16'd50097});
	test_expansion(128'hc78c2f8fbc9733816e42eff0d693b636, {16'd3985, 16'd46713, 16'd60992, 16'd35599, 16'd18412, 16'd31912, 16'd53701, 16'd45256, 16'd9115, 16'd58583, 16'd57828, 16'd37470, 16'd64269, 16'd57157, 16'd41314, 16'd25232, 16'd43203, 16'd26132, 16'd9191, 16'd1836, 16'd52942, 16'd43140, 16'd17899, 16'd22926, 16'd20293, 16'd30349});
	test_expansion(128'h0d47cf15e74f8be69381e8b18f6a42cb, {16'd46937, 16'd22073, 16'd32013, 16'd26732, 16'd46121, 16'd23347, 16'd55231, 16'd64388, 16'd54437, 16'd53411, 16'd35694, 16'd65406, 16'd30223, 16'd9985, 16'd49558, 16'd16708, 16'd52483, 16'd38347, 16'd16012, 16'd6553, 16'd58748, 16'd18648, 16'd6022, 16'd35513, 16'd43537, 16'd61237});
	test_expansion(128'h9222ff45d4cdc26681d7393096c02b9b, {16'd62195, 16'd12238, 16'd42833, 16'd43157, 16'd55003, 16'd50870, 16'd62454, 16'd44059, 16'd40635, 16'd6515, 16'd63789, 16'd23686, 16'd39838, 16'd82, 16'd44973, 16'd51182, 16'd5888, 16'd14776, 16'd48565, 16'd4857, 16'd64482, 16'd55335, 16'd48974, 16'd51538, 16'd37568, 16'd18623});
	test_expansion(128'hb770055f56dd405ef6a79ebb7e2a9fa9, {16'd61497, 16'd49515, 16'd5292, 16'd4044, 16'd39631, 16'd60765, 16'd36842, 16'd19419, 16'd37915, 16'd36096, 16'd31115, 16'd30365, 16'd44340, 16'd42370, 16'd12684, 16'd29318, 16'd17630, 16'd50809, 16'd27570, 16'd36705, 16'd38443, 16'd7137, 16'd9592, 16'd26234, 16'd40339, 16'd57132});
	test_expansion(128'h2982ef9c6adf5f0bcaf7c556c4512bb8, {16'd62137, 16'd23865, 16'd53316, 16'd60506, 16'd44359, 16'd10837, 16'd39920, 16'd38207, 16'd5495, 16'd47725, 16'd54151, 16'd16642, 16'd48545, 16'd26579, 16'd13955, 16'd34116, 16'd20199, 16'd24435, 16'd33133, 16'd56527, 16'd29546, 16'd55527, 16'd37223, 16'd62322, 16'd30532, 16'd59639});
	test_expansion(128'h86638e352b96572ec4e291d2e21e8ef7, {16'd63329, 16'd23575, 16'd28625, 16'd9801, 16'd6960, 16'd49634, 16'd12858, 16'd4185, 16'd42648, 16'd20238, 16'd44763, 16'd35070, 16'd45211, 16'd27635, 16'd30644, 16'd63385, 16'd57425, 16'd43449, 16'd64456, 16'd3764, 16'd43102, 16'd60713, 16'd46763, 16'd35707, 16'd4694, 16'd41207});
	test_expansion(128'h645bbbb554feec01ee87a715ad7027e5, {16'd55579, 16'd27692, 16'd57828, 16'd12772, 16'd38738, 16'd4709, 16'd24063, 16'd54207, 16'd23765, 16'd34915, 16'd16619, 16'd28012, 16'd21693, 16'd56607, 16'd20629, 16'd50715, 16'd4428, 16'd62258, 16'd8422, 16'd62828, 16'd18558, 16'd5993, 16'd58715, 16'd1082, 16'd39156, 16'd9972});
	test_expansion(128'h8342f660521f53200f519ddd48589dc7, {16'd13297, 16'd6705, 16'd38342, 16'd13099, 16'd11822, 16'd58675, 16'd61813, 16'd45085, 16'd294, 16'd61647, 16'd37841, 16'd57600, 16'd12496, 16'd60915, 16'd53617, 16'd31021, 16'd46329, 16'd4749, 16'd14150, 16'd49839, 16'd14425, 16'd57580, 16'd44437, 16'd17717, 16'd6496, 16'd8666});
	test_expansion(128'hde9862b6c36b806abe3cbb3ca0552548, {16'd49612, 16'd53015, 16'd26212, 16'd47563, 16'd63121, 16'd7137, 16'd9415, 16'd23293, 16'd9313, 16'd17896, 16'd23829, 16'd40469, 16'd15269, 16'd1188, 16'd31238, 16'd60954, 16'd23504, 16'd16797, 16'd14777, 16'd54717, 16'd10228, 16'd39363, 16'd32386, 16'd46835, 16'd22428, 16'd25126});
	test_expansion(128'h20e1fd072fbdcd28eafbc9205c595af9, {16'd35135, 16'd10110, 16'd64994, 16'd56459, 16'd10234, 16'd57918, 16'd34890, 16'd61342, 16'd44345, 16'd29404, 16'd26253, 16'd38878, 16'd1708, 16'd32053, 16'd40606, 16'd14416, 16'd48336, 16'd12416, 16'd35545, 16'd56304, 16'd19713, 16'd37172, 16'd581, 16'd40626, 16'd46225, 16'd12390});
	test_expansion(128'hb8ef214d59fc7058f8df2ba47d4c118b, {16'd41429, 16'd65324, 16'd33114, 16'd14963, 16'd60783, 16'd10417, 16'd36276, 16'd15786, 16'd52483, 16'd20008, 16'd34380, 16'd4248, 16'd19842, 16'd54167, 16'd51528, 16'd437, 16'd29160, 16'd46837, 16'd52357, 16'd53255, 16'd3643, 16'd50560, 16'd45156, 16'd7453, 16'd62435, 16'd48843});
	test_expansion(128'hdef2c830875ab3e8bccb14f792dceba7, {16'd62029, 16'd172, 16'd37073, 16'd40755, 16'd1599, 16'd11547, 16'd58112, 16'd1439, 16'd24597, 16'd52584, 16'd47227, 16'd34344, 16'd53908, 16'd14364, 16'd30339, 16'd17133, 16'd51995, 16'd19399, 16'd39777, 16'd10526, 16'd46797, 16'd64663, 16'd42198, 16'd38566, 16'd65100, 16'd6820});
	test_expansion(128'ha6a8a19d4077e9a4803d9cf5723fc321, {16'd19829, 16'd665, 16'd17592, 16'd30890, 16'd1406, 16'd8041, 16'd48118, 16'd18031, 16'd20651, 16'd28582, 16'd38711, 16'd26258, 16'd248, 16'd25475, 16'd44040, 16'd35131, 16'd1389, 16'd35410, 16'd24640, 16'd28644, 16'd42973, 16'd123, 16'd31923, 16'd52383, 16'd51807, 16'd12919});
	test_expansion(128'h062acaf8bc50c023dd6b39d82f0bf776, {16'd5404, 16'd19618, 16'd3250, 16'd18186, 16'd29339, 16'd34638, 16'd55116, 16'd24233, 16'd36718, 16'd43662, 16'd27817, 16'd23540, 16'd24369, 16'd50033, 16'd49370, 16'd50735, 16'd46161, 16'd17450, 16'd36297, 16'd65461, 16'd2767, 16'd21993, 16'd33970, 16'd38505, 16'd31982, 16'd38030});
	test_expansion(128'h683846d19c6b60e670176bde8605ef74, {16'd44529, 16'd22007, 16'd57376, 16'd42854, 16'd3584, 16'd28397, 16'd11, 16'd2919, 16'd18046, 16'd55626, 16'd50930, 16'd58824, 16'd44214, 16'd13452, 16'd61016, 16'd56200, 16'd47734, 16'd9691, 16'd27723, 16'd16435, 16'd18553, 16'd64886, 16'd53836, 16'd51804, 16'd49416, 16'd64435});
	test_expansion(128'h7fa2729e240489eeb17ebb5e91182a1c, {16'd51628, 16'd50217, 16'd47173, 16'd17057, 16'd42142, 16'd62399, 16'd864, 16'd6494, 16'd29058, 16'd5263, 16'd2081, 16'd724, 16'd50231, 16'd31903, 16'd33223, 16'd55752, 16'd9741, 16'd8756, 16'd56904, 16'd17043, 16'd53448, 16'd40336, 16'd36901, 16'd64300, 16'd38572, 16'd54012});
	test_expansion(128'h286f82fa1d4a68506fbf9808dfce1278, {16'd59507, 16'd28678, 16'd57062, 16'd20875, 16'd41547, 16'd61444, 16'd21106, 16'd18154, 16'd10145, 16'd46567, 16'd28058, 16'd50848, 16'd41277, 16'd58336, 16'd23440, 16'd57287, 16'd1943, 16'd15109, 16'd572, 16'd2474, 16'd34598, 16'd19425, 16'd58275, 16'd61041, 16'd41551, 16'd7582});
	test_expansion(128'h545e2e2a7cc6f5c86176dbab452848e1, {16'd26467, 16'd41137, 16'd36137, 16'd43338, 16'd5590, 16'd53608, 16'd17209, 16'd54295, 16'd40657, 16'd29240, 16'd5425, 16'd30605, 16'd9654, 16'd20575, 16'd12130, 16'd64721, 16'd47639, 16'd856, 16'd41078, 16'd43224, 16'd1576, 16'd60998, 16'd52607, 16'd14142, 16'd44210, 16'd64618});
	test_expansion(128'h5609ef211972a9df8c622ebb5d7b9e28, {16'd42271, 16'd55747, 16'd1634, 16'd50791, 16'd31525, 16'd23662, 16'd27883, 16'd17304, 16'd32119, 16'd12220, 16'd50612, 16'd1616, 16'd46505, 16'd12018, 16'd59857, 16'd23363, 16'd54559, 16'd1279, 16'd42051, 16'd21186, 16'd65000, 16'd57230, 16'd15421, 16'd35675, 16'd49945, 16'd51220});
	test_expansion(128'h91922c3f59453210f8b4ffce2be8e291, {16'd25712, 16'd35710, 16'd59627, 16'd61606, 16'd46897, 16'd15203, 16'd14240, 16'd4941, 16'd34627, 16'd1477, 16'd1721, 16'd13436, 16'd19625, 16'd58773, 16'd7344, 16'd44960, 16'd58720, 16'd14984, 16'd13587, 16'd46245, 16'd56957, 16'd18442, 16'd13487, 16'd723, 16'd24250, 16'd3410});
	test_expansion(128'hf08e8f35b619f9751d350fcef7f0f804, {16'd15838, 16'd39913, 16'd58438, 16'd21257, 16'd32204, 16'd20433, 16'd23562, 16'd14990, 16'd61214, 16'd34766, 16'd16206, 16'd2229, 16'd40228, 16'd52471, 16'd15243, 16'd34766, 16'd18797, 16'd56365, 16'd57137, 16'd4696, 16'd39547, 16'd8567, 16'd22654, 16'd6254, 16'd45841, 16'd61551});
	test_expansion(128'h407aed8089da58393df480eccf835d2e, {16'd40738, 16'd53, 16'd28598, 16'd4547, 16'd4329, 16'd60877, 16'd5295, 16'd38802, 16'd53073, 16'd2401, 16'd18247, 16'd53399, 16'd19254, 16'd28295, 16'd15105, 16'd12458, 16'd4043, 16'd15542, 16'd44671, 16'd59293, 16'd44418, 16'd3069, 16'd26275, 16'd64875, 16'd34934, 16'd2684});
	test_expansion(128'h0e9c8548dad5b967fb152536eab72365, {16'd14555, 16'd37268, 16'd64301, 16'd29438, 16'd61525, 16'd51496, 16'd65275, 16'd2848, 16'd17375, 16'd32690, 16'd41132, 16'd36149, 16'd11105, 16'd1917, 16'd29198, 16'd52532, 16'd29054, 16'd49045, 16'd9181, 16'd55784, 16'd36223, 16'd48895, 16'd19861, 16'd40348, 16'd25277, 16'd32769});
	test_expansion(128'hdd86b3c72c6bb85f1de045d670b26a47, {16'd64374, 16'd26940, 16'd53799, 16'd20414, 16'd32868, 16'd33810, 16'd22001, 16'd5957, 16'd10912, 16'd19506, 16'd48887, 16'd62480, 16'd17089, 16'd31807, 16'd33165, 16'd4779, 16'd62060, 16'd31315, 16'd34755, 16'd46196, 16'd7215, 16'd52434, 16'd19331, 16'd51566, 16'd19117, 16'd17284});
	test_expansion(128'h2ac40fca3287f432fbcdde7639b25d03, {16'd40410, 16'd8255, 16'd54728, 16'd46664, 16'd4648, 16'd14561, 16'd60298, 16'd3081, 16'd59574, 16'd63333, 16'd23613, 16'd20041, 16'd22644, 16'd40194, 16'd27470, 16'd30248, 16'd10912, 16'd30258, 16'd61811, 16'd14759, 16'd47827, 16'd51498, 16'd60059, 16'd10775, 16'd4238, 16'd10856});
	test_expansion(128'h8b2cb2088db96b36bef74fe2aa9759d1, {16'd47209, 16'd62896, 16'd58147, 16'd33202, 16'd8814, 16'd62648, 16'd1924, 16'd23994, 16'd37640, 16'd47281, 16'd44738, 16'd28087, 16'd41695, 16'd28288, 16'd19107, 16'd8056, 16'd53276, 16'd17031, 16'd36327, 16'd8702, 16'd28678, 16'd62577, 16'd14129, 16'd24066, 16'd7410, 16'd65069});
	test_expansion(128'h6371f3459b8ac68f20b0656c9ccafa2b, {16'd27541, 16'd50341, 16'd28270, 16'd48595, 16'd56460, 16'd28886, 16'd27272, 16'd51550, 16'd59566, 16'd1033, 16'd22319, 16'd21897, 16'd11432, 16'd24559, 16'd41255, 16'd16473, 16'd14495, 16'd64259, 16'd27066, 16'd17738, 16'd39302, 16'd55171, 16'd23143, 16'd60975, 16'd4181, 16'd28256});
	test_expansion(128'h7aec816ba5fd1ed79e886a7700819b31, {16'd13651, 16'd53486, 16'd62872, 16'd49641, 16'd13440, 16'd27388, 16'd64, 16'd47982, 16'd62333, 16'd44646, 16'd25857, 16'd35647, 16'd61881, 16'd2245, 16'd36717, 16'd29371, 16'd30549, 16'd33948, 16'd62992, 16'd30033, 16'd55771, 16'd17661, 16'd40139, 16'd30108, 16'd52224, 16'd26464});
	test_expansion(128'h6e1ca2a2a27124477e14a8b0828110f9, {16'd17271, 16'd20967, 16'd62355, 16'd51048, 16'd7638, 16'd47023, 16'd27707, 16'd60801, 16'd1096, 16'd40080, 16'd12955, 16'd35267, 16'd28588, 16'd35179, 16'd22437, 16'd59753, 16'd22115, 16'd41700, 16'd8349, 16'd26925, 16'd16276, 16'd29871, 16'd58832, 16'd45482, 16'd13283, 16'd14896});
	test_expansion(128'h392a09874f67038c471111361ac65e5e, {16'd48229, 16'd59254, 16'd35551, 16'd62553, 16'd52072, 16'd18501, 16'd25186, 16'd31560, 16'd59133, 16'd7819, 16'd14898, 16'd29548, 16'd6019, 16'd22550, 16'd26220, 16'd13288, 16'd51629, 16'd16525, 16'd31161, 16'd57797, 16'd63764, 16'd33550, 16'd16883, 16'd35345, 16'd56552, 16'd29056});
	test_expansion(128'hfd2bc639096e667c31567bdb5ea3574d, {16'd65086, 16'd63115, 16'd50833, 16'd52054, 16'd50551, 16'd53122, 16'd46457, 16'd18148, 16'd63610, 16'd50195, 16'd53519, 16'd57410, 16'd63493, 16'd1273, 16'd281, 16'd34526, 16'd19504, 16'd3343, 16'd32894, 16'd35603, 16'd15547, 16'd13781, 16'd53502, 16'd1782, 16'd30366, 16'd48200});
	test_expansion(128'he52cb96b438c8ece9653fa542b4874a6, {16'd19354, 16'd28187, 16'd29789, 16'd57739, 16'd25669, 16'd11508, 16'd44040, 16'd23580, 16'd36283, 16'd54991, 16'd20174, 16'd59547, 16'd45976, 16'd31934, 16'd27426, 16'd15170, 16'd24204, 16'd19235, 16'd11901, 16'd15111, 16'd46383, 16'd39822, 16'd51214, 16'd28587, 16'd48954, 16'd60075});
	test_expansion(128'hfd8bb7e6f5ede45616ebccf160143dce, {16'd55921, 16'd17868, 16'd7554, 16'd9746, 16'd14747, 16'd16155, 16'd4413, 16'd12039, 16'd47623, 16'd39902, 16'd30080, 16'd22519, 16'd36547, 16'd9144, 16'd1583, 16'd1921, 16'd4315, 16'd30975, 16'd24524, 16'd28045, 16'd39540, 16'd5057, 16'd20352, 16'd45181, 16'd42844, 16'd2598});
	test_expansion(128'hd87d083c174b699db69bd935097594ec, {16'd30929, 16'd16870, 16'd27627, 16'd55259, 16'd5670, 16'd38792, 16'd406, 16'd41637, 16'd31833, 16'd32345, 16'd4686, 16'd52890, 16'd23334, 16'd55261, 16'd42077, 16'd47783, 16'd18881, 16'd61321, 16'd55964, 16'd22132, 16'd7765, 16'd11270, 16'd37460, 16'd20457, 16'd63036, 16'd10685});
	test_expansion(128'hbf160b5997838fb6feb79a00c69ffde5, {16'd36897, 16'd4880, 16'd33502, 16'd27453, 16'd30274, 16'd41584, 16'd6243, 16'd59008, 16'd4764, 16'd24505, 16'd21151, 16'd10477, 16'd56721, 16'd46701, 16'd19006, 16'd34710, 16'd53166, 16'd6400, 16'd6776, 16'd35803, 16'd54699, 16'd4593, 16'd10645, 16'd28473, 16'd47936, 16'd18499});
	test_expansion(128'hdd5e169ab96f1ff5de79d127558d2e81, {16'd55269, 16'd57182, 16'd58242, 16'd56465, 16'd11877, 16'd12700, 16'd4823, 16'd29723, 16'd23358, 16'd60880, 16'd54103, 16'd52870, 16'd64424, 16'd3124, 16'd64948, 16'd35915, 16'd6797, 16'd2261, 16'd59577, 16'd52562, 16'd39740, 16'd50199, 16'd34187, 16'd65273, 16'd22435, 16'd33046});
	test_expansion(128'h50575c37359f2308b405f204a3f26a02, {16'd28496, 16'd58325, 16'd16194, 16'd27630, 16'd62277, 16'd17373, 16'd2187, 16'd65336, 16'd56105, 16'd30500, 16'd63468, 16'd44797, 16'd41359, 16'd36473, 16'd12731, 16'd58034, 16'd13333, 16'd15037, 16'd55244, 16'd13064, 16'd24844, 16'd34898, 16'd6640, 16'd33519, 16'd54742, 16'd50628});
	test_expansion(128'hdd92ce49afd83ad1410f90a9eb2ab2df, {16'd52992, 16'd42568, 16'd61810, 16'd2513, 16'd57025, 16'd15502, 16'd63465, 16'd47465, 16'd7534, 16'd23502, 16'd3827, 16'd20087, 16'd6285, 16'd11641, 16'd36420, 16'd50503, 16'd37479, 16'd16220, 16'd194, 16'd42039, 16'd45792, 16'd51529, 16'd29583, 16'd4376, 16'd37796, 16'd19237});
	test_expansion(128'h16d91025e7fa00f139d2aa91855aea93, {16'd23819, 16'd62022, 16'd15422, 16'd50235, 16'd33202, 16'd36071, 16'd33505, 16'd24186, 16'd509, 16'd4364, 16'd58334, 16'd3961, 16'd30523, 16'd51389, 16'd44818, 16'd10653, 16'd53554, 16'd2503, 16'd60047, 16'd35693, 16'd16583, 16'd27501, 16'd13833, 16'd14537, 16'd4356, 16'd55577});
	test_expansion(128'hfaa790b595dcd8def7afd422815abe9f, {16'd14872, 16'd55724, 16'd31435, 16'd47049, 16'd56987, 16'd34543, 16'd41127, 16'd48846, 16'd23150, 16'd7808, 16'd28927, 16'd30622, 16'd6080, 16'd27371, 16'd38962, 16'd29514, 16'd42234, 16'd53308, 16'd49685, 16'd42032, 16'd51900, 16'd41112, 16'd45786, 16'd3152, 16'd18465, 16'd36422});
	test_expansion(128'h6e4787ae8d20fcf23df6db09fe3a5799, {16'd41758, 16'd12163, 16'd4291, 16'd17713, 16'd7862, 16'd29264, 16'd38954, 16'd534, 16'd45363, 16'd65088, 16'd23859, 16'd61962, 16'd38927, 16'd16088, 16'd9686, 16'd37134, 16'd4827, 16'd47013, 16'd2846, 16'd42649, 16'd61594, 16'd59595, 16'd5363, 16'd65043, 16'd21504, 16'd54057});
	test_expansion(128'h54d52220b56a6b93782e58ae31d592c0, {16'd52484, 16'd41871, 16'd5652, 16'd48671, 16'd60145, 16'd59536, 16'd686, 16'd10746, 16'd6358, 16'd31903, 16'd1374, 16'd21982, 16'd4696, 16'd22689, 16'd18574, 16'd7159, 16'd34993, 16'd39533, 16'd38655, 16'd3563, 16'd59469, 16'd62584, 16'd29336, 16'd41395, 16'd4371, 16'd30045});
	test_expansion(128'hae5b750d3b81892d70ce9f047a5588d7, {16'd41993, 16'd6161, 16'd38071, 16'd349, 16'd31991, 16'd10071, 16'd11297, 16'd60294, 16'd22615, 16'd7391, 16'd22637, 16'd39194, 16'd15976, 16'd273, 16'd13817, 16'd34860, 16'd13652, 16'd4955, 16'd6270, 16'd35535, 16'd49463, 16'd24525, 16'd16233, 16'd35461, 16'd62452, 16'd16392});
	test_expansion(128'h706f2e0b3d920c108d4237594a88f0f9, {16'd5481, 16'd59542, 16'd2772, 16'd62865, 16'd9349, 16'd50488, 16'd33617, 16'd31404, 16'd41003, 16'd61536, 16'd64941, 16'd8719, 16'd18217, 16'd53376, 16'd14936, 16'd34143, 16'd40894, 16'd19209, 16'd11688, 16'd60747, 16'd30727, 16'd64861, 16'd45126, 16'd11797, 16'd57755, 16'd6415});
	test_expansion(128'h45c4a5279d9a968c97c9960ed418962f, {16'd25659, 16'd61766, 16'd25709, 16'd53448, 16'd37682, 16'd15399, 16'd63923, 16'd46647, 16'd42448, 16'd18532, 16'd58268, 16'd65123, 16'd27970, 16'd10993, 16'd46324, 16'd27530, 16'd4921, 16'd22446, 16'd805, 16'd49393, 16'd23663, 16'd7770, 16'd38034, 16'd48955, 16'd13308, 16'd54494});
	test_expansion(128'h09350d59b685635066b2891fc6323a4c, {16'd1298, 16'd47159, 16'd26780, 16'd59, 16'd41847, 16'd53105, 16'd7313, 16'd44264, 16'd26944, 16'd20359, 16'd59743, 16'd64805, 16'd39, 16'd25071, 16'd62387, 16'd18624, 16'd51228, 16'd40814, 16'd61510, 16'd39789, 16'd53045, 16'd8680, 16'd21412, 16'd63256, 16'd23198, 16'd46411});
	test_expansion(128'hc038088e3ba885a3523f0057b4c7207a, {16'd52771, 16'd13402, 16'd53609, 16'd36411, 16'd33274, 16'd5457, 16'd12132, 16'd46686, 16'd36245, 16'd24901, 16'd57328, 16'd56581, 16'd17246, 16'd41912, 16'd17386, 16'd17198, 16'd11035, 16'd4067, 16'd3443, 16'd25408, 16'd22841, 16'd20640, 16'd10175, 16'd23934, 16'd44289, 16'd30920});
	test_expansion(128'hab5afe00fba75fde3ef675f4e1b45159, {16'd62329, 16'd38665, 16'd11517, 16'd4863, 16'd29604, 16'd19342, 16'd12049, 16'd42905, 16'd58736, 16'd47052, 16'd64369, 16'd723, 16'd28915, 16'd45425, 16'd1601, 16'd14453, 16'd51678, 16'd35074, 16'd27386, 16'd33920, 16'd29518, 16'd52197, 16'd17204, 16'd45848, 16'd38588, 16'd28546});
	test_expansion(128'h4438ac42e2dfb82acffd2258b86db526, {16'd43395, 16'd8696, 16'd22732, 16'd63802, 16'd52910, 16'd22778, 16'd60430, 16'd60985, 16'd12657, 16'd21172, 16'd27277, 16'd63246, 16'd41281, 16'd64023, 16'd23472, 16'd46883, 16'd24658, 16'd55572, 16'd42355, 16'd10114, 16'd4256, 16'd3724, 16'd3012, 16'd46595, 16'd12985, 16'd54847});
	test_expansion(128'hf2875bdb2d08e34b11fec85795a63acc, {16'd53650, 16'd45658, 16'd36971, 16'd33228, 16'd50745, 16'd28442, 16'd32264, 16'd59650, 16'd691, 16'd16027, 16'd43096, 16'd41100, 16'd21310, 16'd22612, 16'd20949, 16'd60061, 16'd51583, 16'd35822, 16'd57299, 16'd62506, 16'd11244, 16'd59152, 16'd29175, 16'd52540, 16'd57471, 16'd56773});
	test_expansion(128'hb1757808a4a10d47dab3113548fa31ad, {16'd38012, 16'd26074, 16'd28975, 16'd44673, 16'd14187, 16'd29075, 16'd52686, 16'd58524, 16'd44116, 16'd27372, 16'd46898, 16'd58018, 16'd2959, 16'd58798, 16'd28980, 16'd46895, 16'd53534, 16'd55010, 16'd38603, 16'd1594, 16'd44902, 16'd11583, 16'd10484, 16'd55376, 16'd52144, 16'd26622});
	test_expansion(128'he616c2b945ab8016389c58dd94aba7e7, {16'd22602, 16'd12747, 16'd33985, 16'd57629, 16'd10873, 16'd43401, 16'd17121, 16'd11033, 16'd8114, 16'd38399, 16'd63866, 16'd8403, 16'd52976, 16'd30254, 16'd3230, 16'd2832, 16'd272, 16'd37826, 16'd57715, 16'd3, 16'd51821, 16'd44423, 16'd48440, 16'd56491, 16'd6363, 16'd59888});
	test_expansion(128'h0cb7f8312fe7e6704aa40e89bacf5092, {16'd33865, 16'd55716, 16'd7182, 16'd56494, 16'd23574, 16'd58226, 16'd62522, 16'd32368, 16'd1879, 16'd26667, 16'd42154, 16'd539, 16'd19331, 16'd18633, 16'd30366, 16'd65095, 16'd24946, 16'd24932, 16'd64207, 16'd3701, 16'd46311, 16'd51875, 16'd30122, 16'd13945, 16'd15291, 16'd43338});
	test_expansion(128'h9650250c19aabca000682666faf12d2e, {16'd25435, 16'd8082, 16'd38885, 16'd13173, 16'd54408, 16'd30671, 16'd31375, 16'd53726, 16'd18456, 16'd49658, 16'd12714, 16'd47866, 16'd13707, 16'd34693, 16'd48221, 16'd15250, 16'd4256, 16'd15286, 16'd14263, 16'd51921, 16'd31646, 16'd37036, 16'd7781, 16'd7927, 16'd52485, 16'd65295});
	test_expansion(128'hd77bc9ed8ba92a87091517a27269bb24, {16'd6117, 16'd18817, 16'd3119, 16'd56252, 16'd20787, 16'd58395, 16'd24941, 16'd25196, 16'd52086, 16'd2884, 16'd30612, 16'd58377, 16'd29734, 16'd49772, 16'd4673, 16'd19159, 16'd2344, 16'd46498, 16'd9755, 16'd21904, 16'd6936, 16'd44273, 16'd27410, 16'd34294, 16'd35287, 16'd34931});
	test_expansion(128'h03fbf5b26de03723074ddd05a622e13c, {16'd45735, 16'd50415, 16'd8332, 16'd60071, 16'd13878, 16'd41950, 16'd8320, 16'd17479, 16'd36533, 16'd48888, 16'd39142, 16'd18374, 16'd48079, 16'd2474, 16'd38697, 16'd28638, 16'd19018, 16'd55321, 16'd60772, 16'd46991, 16'd32956, 16'd2174, 16'd18886, 16'd38011, 16'd17516, 16'd30486});
	test_expansion(128'h1ab55362cbc676392b324c6838b07b4b, {16'd42059, 16'd31936, 16'd2908, 16'd38019, 16'd49356, 16'd52760, 16'd11799, 16'd35519, 16'd10285, 16'd26245, 16'd37145, 16'd61971, 16'd50253, 16'd6149, 16'd15206, 16'd26094, 16'd52410, 16'd13118, 16'd25012, 16'd37894, 16'd6835, 16'd527, 16'd35577, 16'd56100, 16'd23891, 16'd32463});
	test_expansion(128'h2c5b44ab81e52f955836cc6ec23ac1bd, {16'd11589, 16'd6696, 16'd2574, 16'd39197, 16'd60531, 16'd12957, 16'd48122, 16'd62734, 16'd18148, 16'd39706, 16'd42743, 16'd3722, 16'd20960, 16'd26210, 16'd40346, 16'd40268, 16'd29192, 16'd28229, 16'd38508, 16'd6017, 16'd52888, 16'd64810, 16'd13163, 16'd4960, 16'd59402, 16'd16675});
	test_expansion(128'hc69786a26d54f503ab096526ee3725cd, {16'd46873, 16'd60447, 16'd65139, 16'd41355, 16'd18681, 16'd16679, 16'd43621, 16'd24795, 16'd1277, 16'd62175, 16'd49088, 16'd20028, 16'd47179, 16'd28426, 16'd54148, 16'd52116, 16'd15838, 16'd16586, 16'd49790, 16'd31184, 16'd40524, 16'd21998, 16'd2195, 16'd49932, 16'd26103, 16'd14563});
	test_expansion(128'hdc6ce9a28bb2e63d72193171bc82a157, {16'd1605, 16'd4136, 16'd42522, 16'd38216, 16'd28747, 16'd9140, 16'd22631, 16'd41625, 16'd36119, 16'd48805, 16'd58636, 16'd45155, 16'd22328, 16'd21897, 16'd62703, 16'd59340, 16'd15890, 16'd30643, 16'd35489, 16'd12666, 16'd26410, 16'd12464, 16'd57582, 16'd12985, 16'd38626, 16'd64342});
	test_expansion(128'h73fd296cc5746f64bf21fce8d3b5aa57, {16'd28593, 16'd30900, 16'd2209, 16'd9919, 16'd15615, 16'd10936, 16'd52985, 16'd38078, 16'd9124, 16'd32492, 16'd50258, 16'd4393, 16'd7372, 16'd6715, 16'd54371, 16'd32916, 16'd61105, 16'd25405, 16'd23396, 16'd57877, 16'd45701, 16'd62127, 16'd1612, 16'd63843, 16'd15576, 16'd62397});
	test_expansion(128'ha4b887671a40e54d2d2138c759b38338, {16'd11299, 16'd56567, 16'd19674, 16'd1901, 16'd51344, 16'd44006, 16'd50609, 16'd13976, 16'd45075, 16'd54110, 16'd65189, 16'd44824, 16'd24216, 16'd32525, 16'd1663, 16'd15004, 16'd55278, 16'd46280, 16'd18666, 16'd47253, 16'd23873, 16'd18300, 16'd55096, 16'd63121, 16'd48748, 16'd10293});
	test_expansion(128'h9080cb2cde2524dd3ef6551a20550495, {16'd21276, 16'd13310, 16'd44613, 16'd60901, 16'd20843, 16'd20744, 16'd18960, 16'd25635, 16'd4854, 16'd49322, 16'd6282, 16'd59041, 16'd46990, 16'd5888, 16'd10368, 16'd58428, 16'd45355, 16'd62035, 16'd57537, 16'd5038, 16'd6830, 16'd64258, 16'd5597, 16'd37858, 16'd51048, 16'd5073});
	test_expansion(128'h8f4f7933a35a67b28e93e98403bafb12, {16'd46421, 16'd50611, 16'd34653, 16'd28667, 16'd47863, 16'd7498, 16'd812, 16'd16772, 16'd60381, 16'd27105, 16'd38471, 16'd40638, 16'd31514, 16'd44090, 16'd47047, 16'd31650, 16'd29649, 16'd6145, 16'd60840, 16'd21696, 16'd45376, 16'd47432, 16'd38243, 16'd9796, 16'd58994, 16'd37560});
	test_expansion(128'h87ff0b799e2ae6138eb9cfe372b3777b, {16'd46424, 16'd42271, 16'd65320, 16'd2370, 16'd12003, 16'd17539, 16'd65174, 16'd23315, 16'd6461, 16'd25012, 16'd39984, 16'd49924, 16'd62345, 16'd4116, 16'd10538, 16'd62802, 16'd33300, 16'd2930, 16'd49475, 16'd7657, 16'd1162, 16'd16356, 16'd50025, 16'd19141, 16'd56424, 16'd10243});
	test_expansion(128'h2b6e49e949200022a56715c0d44cade5, {16'd54616, 16'd47704, 16'd14797, 16'd6442, 16'd14661, 16'd16825, 16'd17898, 16'd44234, 16'd30365, 16'd59116, 16'd36822, 16'd11857, 16'd12249, 16'd56119, 16'd36069, 16'd46814, 16'd34679, 16'd28573, 16'd28713, 16'd51124, 16'd9902, 16'd30683, 16'd33742, 16'd19290, 16'd31982, 16'd39719});
	test_expansion(128'hafe703011f924858d2a02a31f02b9a2a, {16'd16002, 16'd50617, 16'd21708, 16'd19748, 16'd63485, 16'd4829, 16'd3171, 16'd45355, 16'd29474, 16'd49783, 16'd1886, 16'd4712, 16'd49091, 16'd56054, 16'd54178, 16'd36132, 16'd14840, 16'd60485, 16'd413, 16'd18900, 16'd9307, 16'd5815, 16'd17195, 16'd35259, 16'd36911, 16'd61685});
	test_expansion(128'h013f1bbc737e6c09c3878c65a9010b48, {16'd45476, 16'd45416, 16'd60301, 16'd61233, 16'd27729, 16'd16993, 16'd9609, 16'd38168, 16'd63406, 16'd62290, 16'd44477, 16'd44929, 16'd28842, 16'd2365, 16'd21286, 16'd26161, 16'd47062, 16'd38249, 16'd45487, 16'd41404, 16'd58150, 16'd9731, 16'd4296, 16'd18960, 16'd41518, 16'd53354});
	test_expansion(128'h5a9b35d789a7c4f04526ed8bbb05ce29, {16'd27848, 16'd40171, 16'd35121, 16'd35968, 16'd5783, 16'd34557, 16'd2346, 16'd41139, 16'd24577, 16'd55345, 16'd37097, 16'd29626, 16'd38978, 16'd63283, 16'd14858, 16'd61709, 16'd22357, 16'd4870, 16'd39838, 16'd33627, 16'd12165, 16'd24543, 16'd41308, 16'd20436, 16'd34374, 16'd42022});
	test_expansion(128'hdba2d93a9353752499d5627d1cd8b927, {16'd51897, 16'd61896, 16'd34543, 16'd31690, 16'd7926, 16'd45753, 16'd12302, 16'd31118, 16'd1087, 16'd62645, 16'd29384, 16'd47438, 16'd38195, 16'd12895, 16'd17019, 16'd45389, 16'd32516, 16'd9303, 16'd37934, 16'd31970, 16'd30617, 16'd18589, 16'd58465, 16'd47885, 16'd47753, 16'd62220});
	test_expansion(128'h008196122bf7ad373e0acc149de5f1de, {16'd38325, 16'd18030, 16'd54929, 16'd12368, 16'd48895, 16'd7376, 16'd59417, 16'd43405, 16'd41968, 16'd42804, 16'd29521, 16'd9527, 16'd19157, 16'd17357, 16'd46269, 16'd27480, 16'd34009, 16'd57355, 16'd26460, 16'd22801, 16'd53793, 16'd12585, 16'd61516, 16'd31981, 16'd6029, 16'd35054});
	test_expansion(128'he44290f770d1f433b4edc578471338aa, {16'd19752, 16'd45874, 16'd57149, 16'd45100, 16'd6392, 16'd56768, 16'd20231, 16'd15619, 16'd43182, 16'd3062, 16'd9939, 16'd705, 16'd18173, 16'd52088, 16'd5091, 16'd60450, 16'd62418, 16'd19169, 16'd55484, 16'd63260, 16'd29798, 16'd41676, 16'd23385, 16'd61868, 16'd37608, 16'd53129});
	test_expansion(128'h3d52288ec11a2873e533e011f2a77206, {16'd22679, 16'd25074, 16'd15550, 16'd46716, 16'd18417, 16'd51325, 16'd62732, 16'd54812, 16'd31489, 16'd13525, 16'd59989, 16'd27096, 16'd24036, 16'd1861, 16'd18213, 16'd47532, 16'd5858, 16'd7713, 16'd7232, 16'd45701, 16'd28109, 16'd12455, 16'd26911, 16'd41688, 16'd50286, 16'd39517});
	test_expansion(128'hfb30d86298f30423368b2e79c4b39dde, {16'd7783, 16'd50967, 16'd54396, 16'd56916, 16'd38590, 16'd14645, 16'd6899, 16'd41870, 16'd60142, 16'd36743, 16'd23649, 16'd40222, 16'd6350, 16'd60329, 16'd46171, 16'd61983, 16'd37440, 16'd18870, 16'd11308, 16'd12469, 16'd49694, 16'd38726, 16'd24628, 16'd29956, 16'd54468, 16'd23969});
	test_expansion(128'hc69944bdee23e13ee9d5328adb7a1fc8, {16'd63354, 16'd53460, 16'd264, 16'd44528, 16'd2008, 16'd12466, 16'd20574, 16'd44847, 16'd48806, 16'd1331, 16'd51440, 16'd23808, 16'd6225, 16'd13088, 16'd23158, 16'd1550, 16'd245, 16'd61773, 16'd6459, 16'd5732, 16'd24588, 16'd23121, 16'd50468, 16'd5705, 16'd28835, 16'd9031});
	test_expansion(128'h8417c8280844035a6cd7be45f2d4dd63, {16'd48135, 16'd5947, 16'd59697, 16'd24706, 16'd47268, 16'd48783, 16'd34993, 16'd16456, 16'd29891, 16'd61632, 16'd42793, 16'd22253, 16'd13259, 16'd26949, 16'd3570, 16'd513, 16'd52613, 16'd63578, 16'd3066, 16'd19680, 16'd17043, 16'd19704, 16'd64394, 16'd56025, 16'd20443, 16'd31073});
	test_expansion(128'hd15fda2094a7b566cff253612812bbb6, {16'd30899, 16'd22652, 16'd25487, 16'd9760, 16'd60565, 16'd30716, 16'd21093, 16'd48589, 16'd43517, 16'd57846, 16'd30166, 16'd7149, 16'd37082, 16'd36180, 16'd15405, 16'd35460, 16'd43913, 16'd6481, 16'd12020, 16'd15702, 16'd18483, 16'd64436, 16'd48817, 16'd19485, 16'd60484, 16'd26716});
	test_expansion(128'hdcb687273f357e8097a698ff38064b9e, {16'd21731, 16'd1746, 16'd45060, 16'd25976, 16'd37215, 16'd20389, 16'd14474, 16'd41321, 16'd8843, 16'd16489, 16'd55418, 16'd15348, 16'd9889, 16'd36670, 16'd28419, 16'd49355, 16'd44077, 16'd38434, 16'd14300, 16'd21066, 16'd47995, 16'd17647, 16'd47613, 16'd46012, 16'd44511, 16'd55113});
	test_expansion(128'hd9948422c21b5cab1b4bc82f3bdcfcdb, {16'd37496, 16'd42797, 16'd52632, 16'd3571, 16'd22012, 16'd55344, 16'd2640, 16'd29198, 16'd15681, 16'd45292, 16'd60068, 16'd23085, 16'd52871, 16'd47538, 16'd29976, 16'd6553, 16'd1883, 16'd31870, 16'd49513, 16'd2234, 16'd61214, 16'd10832, 16'd33892, 16'd50795, 16'd17165, 16'd4289});
	test_expansion(128'hc6b816e5a4c24eec1b477c4c2d9919d0, {16'd18167, 16'd22660, 16'd27207, 16'd48501, 16'd1066, 16'd47710, 16'd40445, 16'd51016, 16'd65228, 16'd61886, 16'd6731, 16'd29920, 16'd17702, 16'd10983, 16'd19914, 16'd2101, 16'd61697, 16'd49551, 16'd43962, 16'd8050, 16'd52731, 16'd43432, 16'd2088, 16'd18632, 16'd39438, 16'd27288});
	test_expansion(128'hd86c41da8fe8bd5f516c85cd473b2948, {16'd2608, 16'd38019, 16'd51397, 16'd32394, 16'd14237, 16'd42833, 16'd7658, 16'd64947, 16'd38329, 16'd38877, 16'd9910, 16'd59237, 16'd37815, 16'd62646, 16'd6662, 16'd2991, 16'd736, 16'd7753, 16'd6892, 16'd16375, 16'd25136, 16'd53296, 16'd35436, 16'd12247, 16'd37494, 16'd40928});
	test_expansion(128'h04bd3c62fe8d4a53899936ed018865ee, {16'd59706, 16'd32389, 16'd55329, 16'd63366, 16'd22795, 16'd32421, 16'd13757, 16'd41689, 16'd3159, 16'd59698, 16'd57442, 16'd27356, 16'd54202, 16'd3740, 16'd26960, 16'd59368, 16'd3927, 16'd56680, 16'd24004, 16'd47116, 16'd58476, 16'd6377, 16'd19979, 16'd24347, 16'd43500, 16'd40681});
	test_expansion(128'ha045535aab124a0b023ef2f23f4c7c1c, {16'd26704, 16'd60489, 16'd27549, 16'd294, 16'd32503, 16'd31786, 16'd2849, 16'd16021, 16'd51796, 16'd26987, 16'd19549, 16'd16987, 16'd60373, 16'd22153, 16'd17524, 16'd14538, 16'd7400, 16'd33978, 16'd59201, 16'd61033, 16'd60770, 16'd6252, 16'd15279, 16'd9442, 16'd21846, 16'd36841});
	test_expansion(128'hdb06a539dfdb2ae70e1401af497be1b4, {16'd8242, 16'd50990, 16'd59633, 16'd43799, 16'd62890, 16'd9726, 16'd1297, 16'd25986, 16'd17303, 16'd39097, 16'd62407, 16'd2316, 16'd11297, 16'd56080, 16'd2262, 16'd28927, 16'd32286, 16'd49237, 16'd63974, 16'd52559, 16'd24869, 16'd36675, 16'd28218, 16'd19140, 16'd55690, 16'd42506});
	test_expansion(128'h765c6d39acdafc9d5fbf85f45dd45a59, {16'd17887, 16'd28994, 16'd11014, 16'd31838, 16'd22997, 16'd49183, 16'd62311, 16'd37656, 16'd37976, 16'd33873, 16'd18184, 16'd20466, 16'd28478, 16'd27348, 16'd15230, 16'd21444, 16'd17415, 16'd17741, 16'd31232, 16'd17418, 16'd38446, 16'd54039, 16'd23431, 16'd5527, 16'd25792, 16'd2330});
	test_expansion(128'h9fb4d4a1034ccdbec570bd0659854b16, {16'd22909, 16'd16653, 16'd35843, 16'd30212, 16'd60620, 16'd37142, 16'd40608, 16'd56769, 16'd3094, 16'd7037, 16'd36669, 16'd44096, 16'd46824, 16'd62619, 16'd20312, 16'd34917, 16'd6235, 16'd48941, 16'd26485, 16'd58082, 16'd2016, 16'd22000, 16'd45784, 16'd233, 16'd57697, 16'd36307});
	test_expansion(128'h0a91c7dfe9e34509cb07b2c1913df9da, {16'd2921, 16'd52529, 16'd39283, 16'd65008, 16'd24919, 16'd40524, 16'd12101, 16'd27701, 16'd14831, 16'd36058, 16'd34993, 16'd26996, 16'd28601, 16'd19563, 16'd25762, 16'd62512, 16'd13560, 16'd35136, 16'd39469, 16'd5172, 16'd30726, 16'd63218, 16'd2373, 16'd56020, 16'd62044, 16'd10332});
	test_expansion(128'h672db02c061160ad1c50543d8960cdf7, {16'd7852, 16'd22906, 16'd23016, 16'd56964, 16'd32618, 16'd4708, 16'd56584, 16'd54594, 16'd40332, 16'd24449, 16'd3802, 16'd39018, 16'd53251, 16'd18390, 16'd51540, 16'd1284, 16'd34662, 16'd18019, 16'd30438, 16'd47312, 16'd3246, 16'd11227, 16'd44766, 16'd2980, 16'd18711, 16'd47596});
	test_expansion(128'h855b68dead0b7242a60b0f496cf86a61, {16'd8669, 16'd10159, 16'd26188, 16'd62388, 16'd29169, 16'd54559, 16'd6886, 16'd5909, 16'd45795, 16'd62275, 16'd46047, 16'd46913, 16'd59093, 16'd50615, 16'd24463, 16'd6836, 16'd29475, 16'd5228, 16'd13810, 16'd12583, 16'd64894, 16'd49571, 16'd63373, 16'd1156, 16'd27222, 16'd17697});
	test_expansion(128'hd3e4f0f680cffed85b333ba074ba44d7, {16'd21212, 16'd49252, 16'd29351, 16'd20940, 16'd53465, 16'd18378, 16'd10933, 16'd39288, 16'd14710, 16'd33677, 16'd35340, 16'd39007, 16'd31252, 16'd43196, 16'd40014, 16'd35003, 16'd12508, 16'd51438, 16'd51581, 16'd43371, 16'd36459, 16'd9700, 16'd48230, 16'd6509, 16'd23345, 16'd62170});
	test_expansion(128'h08dbaf644e298c1d59455cfb18b3f257, {16'd43119, 16'd59537, 16'd46246, 16'd45996, 16'd23910, 16'd51442, 16'd237, 16'd58118, 16'd9669, 16'd14155, 16'd62637, 16'd48844, 16'd10186, 16'd2191, 16'd49021, 16'd22376, 16'd25789, 16'd33941, 16'd45004, 16'd8574, 16'd35540, 16'd60569, 16'd5628, 16'd20061, 16'd8106, 16'd25416});
	test_expansion(128'he97f28f8f4796965fe858db758605901, {16'd47530, 16'd65314, 16'd4825, 16'd24320, 16'd54237, 16'd25988, 16'd44647, 16'd63497, 16'd59345, 16'd7717, 16'd32004, 16'd31972, 16'd8203, 16'd61801, 16'd34616, 16'd47730, 16'd3142, 16'd37258, 16'd14122, 16'd15270, 16'd55642, 16'd1927, 16'd29133, 16'd62615, 16'd56495, 16'd6593});
	test_expansion(128'hda341074013edf5dc4d6053cd065972f, {16'd31743, 16'd28599, 16'd13840, 16'd42816, 16'd43117, 16'd42779, 16'd10028, 16'd49829, 16'd33425, 16'd55952, 16'd24363, 16'd63605, 16'd30210, 16'd40586, 16'd49308, 16'd42052, 16'd49051, 16'd25511, 16'd57013, 16'd21897, 16'd29305, 16'd47328, 16'd1411, 16'd19112, 16'd33801, 16'd44035});
	test_expansion(128'h9695872d8146a8ccf428bea6a15ccde4, {16'd40083, 16'd56651, 16'd42039, 16'd52814, 16'd17739, 16'd36923, 16'd12192, 16'd36113, 16'd38518, 16'd6602, 16'd37693, 16'd65317, 16'd45301, 16'd25568, 16'd3272, 16'd63132, 16'd46228, 16'd11956, 16'd34926, 16'd51290, 16'd33748, 16'd27218, 16'd37097, 16'd34945, 16'd3130, 16'd60383});
	test_expansion(128'hf0080ca400a9b9689b719cbfa4be421f, {16'd25165, 16'd34658, 16'd273, 16'd24636, 16'd24838, 16'd32906, 16'd4619, 16'd33143, 16'd34366, 16'd63561, 16'd62726, 16'd24954, 16'd14606, 16'd33568, 16'd2464, 16'd41455, 16'd58018, 16'd22941, 16'd27174, 16'd36588, 16'd20969, 16'd28785, 16'd31152, 16'd13395, 16'd39627, 16'd7388});
	test_expansion(128'h15afc3cfbac69570683c52831146456d, {16'd20909, 16'd6954, 16'd45345, 16'd40095, 16'd32043, 16'd27028, 16'd12857, 16'd26680, 16'd32189, 16'd32155, 16'd20158, 16'd55286, 16'd35302, 16'd5431, 16'd11777, 16'd32154, 16'd51642, 16'd35523, 16'd6361, 16'd18723, 16'd20091, 16'd63378, 16'd48760, 16'd47815, 16'd7082, 16'd24620});
	test_expansion(128'h46a431bb0b0d66a452ab0c2adfc34a57, {16'd6063, 16'd49383, 16'd27037, 16'd15177, 16'd18395, 16'd25101, 16'd38884, 16'd23332, 16'd2609, 16'd27778, 16'd36599, 16'd639, 16'd36125, 16'd30533, 16'd14820, 16'd33154, 16'd44063, 16'd20812, 16'd43780, 16'd25239, 16'd61827, 16'd27010, 16'd45543, 16'd45604, 16'd17862, 16'd885});
	test_expansion(128'h34141c2004f64ba97cd05afcc6c3ab31, {16'd40526, 16'd59667, 16'd44388, 16'd19532, 16'd38998, 16'd15660, 16'd16384, 16'd40289, 16'd40494, 16'd15678, 16'd29214, 16'd20102, 16'd42150, 16'd8312, 16'd59392, 16'd51350, 16'd34548, 16'd44668, 16'd40230, 16'd38851, 16'd27112, 16'd5070, 16'd54493, 16'd9248, 16'd56580, 16'd20202});
	test_expansion(128'h28f637af461ec47de5206be351ed4e84, {16'd8980, 16'd36529, 16'd37069, 16'd29741, 16'd9424, 16'd33740, 16'd24708, 16'd64705, 16'd55765, 16'd41268, 16'd6651, 16'd15143, 16'd37298, 16'd16677, 16'd10873, 16'd7137, 16'd8239, 16'd38878, 16'd8618, 16'd4629, 16'd64948, 16'd62796, 16'd13587, 16'd29135, 16'd30157, 16'd62747});
	test_expansion(128'hb1e7d20bc1fb1ac4ee415ea69990aa72, {16'd3208, 16'd26385, 16'd55859, 16'd31847, 16'd38725, 16'd47934, 16'd48780, 16'd55853, 16'd48450, 16'd15539, 16'd31266, 16'd37805, 16'd9056, 16'd51747, 16'd49253, 16'd24515, 16'd11857, 16'd40214, 16'd1862, 16'd28996, 16'd34737, 16'd27352, 16'd10560, 16'd33437, 16'd32069, 16'd62615});
	test_expansion(128'ha7f242e34a65a0b34e3b1e05ae598f74, {16'd44334, 16'd20237, 16'd35817, 16'd42549, 16'd48683, 16'd55617, 16'd41246, 16'd63727, 16'd50771, 16'd43481, 16'd49582, 16'd64088, 16'd5027, 16'd29642, 16'd35896, 16'd40861, 16'd17567, 16'd41522, 16'd26345, 16'd4862, 16'd20545, 16'd28416, 16'd31962, 16'd17277, 16'd58559, 16'd27659});
	test_expansion(128'h9b122cb9017343af38f8300b89ab9af4, {16'd52272, 16'd4889, 16'd46921, 16'd51371, 16'd20009, 16'd28657, 16'd7493, 16'd25056, 16'd22286, 16'd36803, 16'd56116, 16'd51975, 16'd57299, 16'd42067, 16'd59117, 16'd9910, 16'd29991, 16'd50016, 16'd3207, 16'd35644, 16'd42675, 16'd33607, 16'd14928, 16'd37508, 16'd4400, 16'd7784});
	test_expansion(128'h2ed8cf11533dd6cef414e23729dd06bc, {16'd56748, 16'd61599, 16'd2505, 16'd48120, 16'd47504, 16'd33047, 16'd51940, 16'd2786, 16'd50573, 16'd24824, 16'd43778, 16'd65228, 16'd15546, 16'd15303, 16'd28334, 16'd39038, 16'd16998, 16'd22492, 16'd36993, 16'd30624, 16'd26885, 16'd27579, 16'd14443, 16'd35300, 16'd23159, 16'd22489});
	test_expansion(128'h0fae209b7725161adc72d96fb31243f3, {16'd22438, 16'd7861, 16'd49035, 16'd51667, 16'd51988, 16'd29976, 16'd50644, 16'd45684, 16'd24141, 16'd4693, 16'd60807, 16'd58074, 16'd29475, 16'd34691, 16'd32625, 16'd52902, 16'd14509, 16'd17919, 16'd22149, 16'd8562, 16'd47600, 16'd4157, 16'd46859, 16'd17671, 16'd55046, 16'd6212});
	test_expansion(128'h82c40e23a83062ca6bd551c7e6e3572f, {16'd17424, 16'd8259, 16'd40066, 16'd10707, 16'd19083, 16'd57965, 16'd21135, 16'd13450, 16'd55719, 16'd47212, 16'd27800, 16'd59780, 16'd30330, 16'd3490, 16'd2636, 16'd47549, 16'd59740, 16'd41333, 16'd61442, 16'd23172, 16'd43967, 16'd64818, 16'd62222, 16'd62572, 16'd31003, 16'd28350});
	test_expansion(128'h263f69f7e10e409c693976eea6321b5c, {16'd4065, 16'd17438, 16'd5732, 16'd32784, 16'd18206, 16'd18335, 16'd49111, 16'd29933, 16'd39159, 16'd54009, 16'd20654, 16'd56937, 16'd25517, 16'd27597, 16'd58492, 16'd58347, 16'd63651, 16'd47430, 16'd36183, 16'd42821, 16'd32288, 16'd63032, 16'd10556, 16'd31371, 16'd40618, 16'd34122});
	test_expansion(128'h04ca068dcfd98f1a53fabcf036d9501b, {16'd43165, 16'd28958, 16'd40691, 16'd60943, 16'd34525, 16'd24649, 16'd60410, 16'd50648, 16'd38443, 16'd58822, 16'd20289, 16'd54345, 16'd12176, 16'd16126, 16'd73, 16'd9215, 16'd43757, 16'd34362, 16'd52255, 16'd43385, 16'd24019, 16'd26829, 16'd29487, 16'd64423, 16'd9130, 16'd1083});
	test_expansion(128'h193033c859cb9aa6c394d7c5b7140ffc, {16'd37022, 16'd5702, 16'd34183, 16'd18116, 16'd50741, 16'd61285, 16'd1986, 16'd53333, 16'd13870, 16'd3877, 16'd45936, 16'd4661, 16'd21573, 16'd49930, 16'd39786, 16'd24087, 16'd18248, 16'd37954, 16'd38172, 16'd35598, 16'd57531, 16'd34340, 16'd64255, 16'd5562, 16'd34489, 16'd51797});
	test_expansion(128'h6b77c63ee52b976ed1fb3db640a6b260, {16'd51753, 16'd41523, 16'd65448, 16'd8188, 16'd21165, 16'd11035, 16'd32109, 16'd45339, 16'd54333, 16'd26789, 16'd19545, 16'd53353, 16'd5348, 16'd20397, 16'd31249, 16'd9830, 16'd16269, 16'd59216, 16'd39574, 16'd29749, 16'd24590, 16'd5286, 16'd20050, 16'd63738, 16'd23438, 16'd47191});
	test_expansion(128'h8e420cc91bbabd78363a0829b92cdc4e, {16'd8954, 16'd57404, 16'd11169, 16'd53768, 16'd33471, 16'd54558, 16'd19193, 16'd50610, 16'd21189, 16'd39610, 16'd49782, 16'd7790, 16'd39048, 16'd16059, 16'd55452, 16'd4045, 16'd45547, 16'd59327, 16'd17640, 16'd130, 16'd25506, 16'd21655, 16'd62909, 16'd47670, 16'd7779, 16'd17145});
	test_expansion(128'h0ae964beef7c14f1866a522161d5606a, {16'd35129, 16'd3251, 16'd8383, 16'd33285, 16'd3109, 16'd14095, 16'd64319, 16'd37631, 16'd12120, 16'd31257, 16'd8253, 16'd58997, 16'd4410, 16'd50033, 16'd4149, 16'd41657, 16'd58235, 16'd12603, 16'd65432, 16'd63792, 16'd29854, 16'd54574, 16'd31966, 16'd43238, 16'd31454, 16'd33222});
	test_expansion(128'hb10f1913299861feab086113850654eb, {16'd16917, 16'd16017, 16'd51318, 16'd44870, 16'd21902, 16'd52039, 16'd12119, 16'd42534, 16'd598, 16'd65171, 16'd62242, 16'd21762, 16'd63452, 16'd24146, 16'd52456, 16'd9522, 16'd16784, 16'd33922, 16'd3251, 16'd25622, 16'd34867, 16'd51250, 16'd31, 16'd22151, 16'd28834, 16'd2868});
	test_expansion(128'h57e42c55dad948deb9b27eac7ac4a3d0, {16'd38739, 16'd65425, 16'd54079, 16'd8414, 16'd32877, 16'd61586, 16'd49148, 16'd32932, 16'd5491, 16'd61139, 16'd40816, 16'd33399, 16'd14332, 16'd28043, 16'd57984, 16'd61739, 16'd24146, 16'd8901, 16'd42165, 16'd52922, 16'd25764, 16'd25790, 16'd61475, 16'd22334, 16'd50414, 16'd13485});
	test_expansion(128'h3e065cfac866269da6a9b2c361e77a8e, {16'd11399, 16'd65341, 16'd20101, 16'd29845, 16'd35039, 16'd33429, 16'd64581, 16'd32523, 16'd45665, 16'd36901, 16'd25857, 16'd21800, 16'd54716, 16'd9228, 16'd800, 16'd16546, 16'd59315, 16'd35581, 16'd45394, 16'd42990, 16'd27160, 16'd58993, 16'd2706, 16'd30395, 16'd39265, 16'd14137});
	test_expansion(128'h612c214272d7f197411659c055b58d4f, {16'd62694, 16'd16318, 16'd5010, 16'd3309, 16'd17271, 16'd52604, 16'd63977, 16'd30380, 16'd44254, 16'd49936, 16'd20358, 16'd58612, 16'd2968, 16'd56105, 16'd58340, 16'd40445, 16'd56569, 16'd2265, 16'd59632, 16'd30487, 16'd58399, 16'd17835, 16'd64214, 16'd51433, 16'd17165, 16'd53239});
	test_expansion(128'hf3269bdc4b74471e29582ae4079df541, {16'd6414, 16'd48798, 16'd61451, 16'd17359, 16'd47376, 16'd49691, 16'd3942, 16'd56842, 16'd17680, 16'd62267, 16'd5273, 16'd6266, 16'd26641, 16'd63106, 16'd22302, 16'd30155, 16'd11731, 16'd41811, 16'd19570, 16'd19959, 16'd6165, 16'd19094, 16'd56865, 16'd2701, 16'd29961, 16'd55175});
	test_expansion(128'hbbf71493c045599889896c577f86177d, {16'd41705, 16'd41917, 16'd14142, 16'd57715, 16'd48759, 16'd48170, 16'd12533, 16'd32890, 16'd944, 16'd43216, 16'd60616, 16'd11684, 16'd60508, 16'd37277, 16'd21100, 16'd56380, 16'd11911, 16'd17230, 16'd11417, 16'd65200, 16'd38677, 16'd19615, 16'd11826, 16'd15876, 16'd4576, 16'd7488});
	test_expansion(128'h771e9026090b1a1c5d840fef0d5a391a, {16'd35163, 16'd52671, 16'd26601, 16'd38798, 16'd48682, 16'd27993, 16'd37399, 16'd39408, 16'd4894, 16'd12380, 16'd9743, 16'd48448, 16'd43007, 16'd36186, 16'd48567, 16'd457, 16'd3631, 16'd28101, 16'd50495, 16'd6911, 16'd55719, 16'd56403, 16'd64434, 16'd59812, 16'd36655, 16'd8482});
	test_expansion(128'h147ec9855806fe01d023894fa6e3292a, {16'd43046, 16'd10988, 16'd6603, 16'd32727, 16'd1344, 16'd37185, 16'd55719, 16'd39627, 16'd1069, 16'd16458, 16'd5960, 16'd32738, 16'd3764, 16'd51995, 16'd10041, 16'd51295, 16'd13899, 16'd3932, 16'd19604, 16'd25254, 16'd36749, 16'd51905, 16'd55022, 16'd32667, 16'd47495, 16'd56751});
	test_expansion(128'hd7418a1db68eca2d0f976bf9574c3065, {16'd10420, 16'd13872, 16'd57474, 16'd60030, 16'd5664, 16'd38357, 16'd16292, 16'd26006, 16'd17818, 16'd22812, 16'd4625, 16'd10325, 16'd47929, 16'd4074, 16'd5627, 16'd46245, 16'd37153, 16'd12924, 16'd39712, 16'd65357, 16'd28679, 16'd24052, 16'd47916, 16'd17751, 16'd52788, 16'd62602});
	test_expansion(128'h3157e58fdde051e0ffee4814f68530d9, {16'd31121, 16'd2816, 16'd26974, 16'd4698, 16'd48936, 16'd43309, 16'd64973, 16'd2941, 16'd16482, 16'd14724, 16'd48244, 16'd33016, 16'd53919, 16'd40902, 16'd27383, 16'd47013, 16'd9001, 16'd4284, 16'd29205, 16'd62476, 16'd41429, 16'd50977, 16'd61692, 16'd41147, 16'd38896, 16'd46851});
	test_expansion(128'h0addf8c961681c9e5c46f0072a4f7c70, {16'd13476, 16'd28904, 16'd27142, 16'd5076, 16'd38019, 16'd20864, 16'd51376, 16'd227, 16'd35687, 16'd42661, 16'd19176, 16'd47846, 16'd49652, 16'd6017, 16'd18617, 16'd5371, 16'd4828, 16'd60535, 16'd10388, 16'd38377, 16'd53999, 16'd9436, 16'd18663, 16'd202, 16'd30745, 16'd20035});
	test_expansion(128'h5ce34a9edb4939694901e5000c76eead, {16'd63657, 16'd43939, 16'd27270, 16'd47210, 16'd34832, 16'd2652, 16'd33109, 16'd15106, 16'd7417, 16'd56267, 16'd60907, 16'd27042, 16'd62566, 16'd40955, 16'd34083, 16'd21448, 16'd27329, 16'd64150, 16'd31536, 16'd52793, 16'd35023, 16'd45469, 16'd10812, 16'd33521, 16'd55114, 16'd27774});
	test_expansion(128'hb99d58cce19a6ce7b5a2d7bd3b4e2a51, {16'd35261, 16'd53443, 16'd62382, 16'd53081, 16'd7906, 16'd51502, 16'd3663, 16'd31944, 16'd36627, 16'd31170, 16'd42407, 16'd31449, 16'd42311, 16'd34000, 16'd58725, 16'd1937, 16'd41823, 16'd61738, 16'd39157, 16'd4647, 16'd30867, 16'd15515, 16'd38843, 16'd12092, 16'd8890, 16'd46573});
	test_expansion(128'hd2572117fae41eb916554b640452497a, {16'd9732, 16'd45002, 16'd61650, 16'd4861, 16'd35848, 16'd40163, 16'd36953, 16'd1180, 16'd22770, 16'd34143, 16'd21945, 16'd15065, 16'd48246, 16'd58922, 16'd46331, 16'd12196, 16'd22729, 16'd54293, 16'd25638, 16'd16223, 16'd10490, 16'd25650, 16'd21890, 16'd10883, 16'd59895, 16'd823});
	test_expansion(128'hf3eea997e1f18f9322f7c8e82843ff56, {16'd29705, 16'd56349, 16'd30753, 16'd5707, 16'd60801, 16'd9213, 16'd18566, 16'd60322, 16'd20882, 16'd62886, 16'd18221, 16'd45860, 16'd35269, 16'd2390, 16'd33042, 16'd15611, 16'd49881, 16'd62174, 16'd45023, 16'd46764, 16'd29801, 16'd9323, 16'd23488, 16'd53085, 16'd9921, 16'd33327});
	test_expansion(128'he358a00c5bec28b28e459361e822a667, {16'd65515, 16'd13605, 16'd30845, 16'd16695, 16'd40978, 16'd44701, 16'd41510, 16'd12025, 16'd59984, 16'd29691, 16'd37735, 16'd42600, 16'd47942, 16'd50770, 16'd19636, 16'd60841, 16'd55790, 16'd14178, 16'd47407, 16'd28565, 16'd56737, 16'd32073, 16'd58905, 16'd56822, 16'd2409, 16'd31810});
	test_expansion(128'h06526f883d7df0d456593fabb9e69796, {16'd7072, 16'd26394, 16'd42345, 16'd48190, 16'd23093, 16'd46146, 16'd48980, 16'd23693, 16'd49090, 16'd33942, 16'd10813, 16'd54532, 16'd64777, 16'd47044, 16'd1700, 16'd7868, 16'd37807, 16'd34082, 16'd54657, 16'd9246, 16'd64717, 16'd21695, 16'd62265, 16'd15484, 16'd10751, 16'd18430});
	test_expansion(128'h0b37d5a4f64f753eb998d3c9be5618c2, {16'd26871, 16'd42977, 16'd21007, 16'd37162, 16'd62851, 16'd46762, 16'd64947, 16'd24122, 16'd35716, 16'd187, 16'd43672, 16'd34189, 16'd17588, 16'd25214, 16'd30412, 16'd37922, 16'd2821, 16'd62133, 16'd56186, 16'd58372, 16'd47600, 16'd6105, 16'd8902, 16'd14280, 16'd17313, 16'd26818});
	test_expansion(128'h7afeb5bbd01ee7f6ef85d8e2327ceee1, {16'd8496, 16'd57733, 16'd8568, 16'd21555, 16'd7707, 16'd32199, 16'd34034, 16'd48757, 16'd37174, 16'd16317, 16'd51435, 16'd45437, 16'd38206, 16'd39661, 16'd7462, 16'd58128, 16'd47952, 16'd36481, 16'd48785, 16'd7511, 16'd3915, 16'd38611, 16'd21441, 16'd48673, 16'd31663, 16'd11017});
	test_expansion(128'h55f29780218f7233fd657f3997c4ddbf, {16'd64126, 16'd36346, 16'd63791, 16'd51445, 16'd41365, 16'd59430, 16'd6869, 16'd8149, 16'd16986, 16'd37665, 16'd20205, 16'd1456, 16'd44044, 16'd40115, 16'd23159, 16'd42155, 16'd53335, 16'd59364, 16'd50830, 16'd61310, 16'd53899, 16'd47956, 16'd62429, 16'd45850, 16'd44385, 16'd12217});
	test_expansion(128'hcd077dc56d56d427969018972c4a3dfd, {16'd28141, 16'd5428, 16'd39987, 16'd59133, 16'd26446, 16'd54405, 16'd18580, 16'd30326, 16'd42727, 16'd4372, 16'd13393, 16'd36177, 16'd27110, 16'd55338, 16'd57855, 16'd33822, 16'd12087, 16'd54855, 16'd3339, 16'd30422, 16'd29518, 16'd2434, 16'd19344, 16'd36447, 16'd204, 16'd14255});
	test_expansion(128'hdb9d5c7efdfa2af4169d101c4d52ff66, {16'd30895, 16'd38386, 16'd64983, 16'd59292, 16'd11587, 16'd7657, 16'd8431, 16'd10993, 16'd6625, 16'd38808, 16'd15788, 16'd60291, 16'd11052, 16'd64152, 16'd41022, 16'd6090, 16'd58974, 16'd30118, 16'd17660, 16'd32084, 16'd22741, 16'd45164, 16'd21838, 16'd17923, 16'd31647, 16'd14321});
	test_expansion(128'h28dfc9ee8374f4fe81aaef0b30bb1365, {16'd9066, 16'd33401, 16'd42641, 16'd5341, 16'd10334, 16'd51465, 16'd61943, 16'd33207, 16'd16407, 16'd43084, 16'd27230, 16'd55041, 16'd24333, 16'd37018, 16'd6027, 16'd32519, 16'd16971, 16'd32636, 16'd45142, 16'd41348, 16'd49952, 16'd11007, 16'd55152, 16'd46125, 16'd10296, 16'd59944});
	test_expansion(128'h5c39af213700930894f2ac042f749644, {16'd34607, 16'd46230, 16'd14136, 16'd26329, 16'd7512, 16'd40749, 16'd44825, 16'd548, 16'd38837, 16'd1550, 16'd56075, 16'd62689, 16'd2818, 16'd63662, 16'd38940, 16'd47156, 16'd11429, 16'd49066, 16'd30341, 16'd54662, 16'd50188, 16'd2895, 16'd39843, 16'd34822, 16'd49823, 16'd62147});
	test_expansion(128'had8eadf87de28fe17bd59912842e9cd6, {16'd11218, 16'd23734, 16'd33190, 16'd2891, 16'd7269, 16'd6631, 16'd60717, 16'd54274, 16'd1862, 16'd63705, 16'd23684, 16'd17645, 16'd45011, 16'd35062, 16'd47817, 16'd48201, 16'd61142, 16'd53077, 16'd11787, 16'd41280, 16'd55987, 16'd10747, 16'd28614, 16'd15459, 16'd14357, 16'd55595});
	test_expansion(128'h5c55efa9844dabe5fad50694208961bf, {16'd36133, 16'd36414, 16'd7474, 16'd51236, 16'd56906, 16'd47026, 16'd9942, 16'd44163, 16'd40642, 16'd17029, 16'd58897, 16'd31295, 16'd49721, 16'd21957, 16'd5927, 16'd17366, 16'd51370, 16'd10016, 16'd15114, 16'd25079, 16'd46104, 16'd58229, 16'd36196, 16'd63295, 16'd34241, 16'd8908});
	test_expansion(128'h26797f6bbdc8ec80d2ee6505edeeb2b0, {16'd63650, 16'd63722, 16'd25356, 16'd65394, 16'd61411, 16'd7228, 16'd32008, 16'd2344, 16'd63134, 16'd65071, 16'd8325, 16'd36369, 16'd40426, 16'd2754, 16'd58801, 16'd22447, 16'd9716, 16'd64901, 16'd49930, 16'd21812, 16'd60988, 16'd54644, 16'd25849, 16'd28365, 16'd20410, 16'd29715});
	test_expansion(128'h44a0056728af22f094a86e782d35caee, {16'd32931, 16'd47525, 16'd33042, 16'd24022, 16'd65351, 16'd60476, 16'd40638, 16'd26934, 16'd2272, 16'd61392, 16'd11277, 16'd13047, 16'd29533, 16'd23726, 16'd19406, 16'd47421, 16'd35412, 16'd11090, 16'd37891, 16'd36876, 16'd40249, 16'd61557, 16'd24532, 16'd15642, 16'd19379, 16'd57734});
	test_expansion(128'h3a89afa42dbc612d469121ba31ac75de, {16'd48622, 16'd8504, 16'd3842, 16'd14963, 16'd6814, 16'd60351, 16'd62015, 16'd9569, 16'd23207, 16'd51234, 16'd24194, 16'd26966, 16'd35794, 16'd23636, 16'd14255, 16'd24175, 16'd20379, 16'd45083, 16'd1951, 16'd12944, 16'd40206, 16'd16701, 16'd60208, 16'd29975, 16'd48196, 16'd48388});
	test_expansion(128'he5bf705965b1765d857c2af1edbce4d7, {16'd27129, 16'd50244, 16'd65445, 16'd38332, 16'd20923, 16'd20044, 16'd51118, 16'd20356, 16'd58091, 16'd19274, 16'd25773, 16'd47098, 16'd48257, 16'd38532, 16'd45813, 16'd51193, 16'd62424, 16'd2013, 16'd34908, 16'd33934, 16'd52845, 16'd58753, 16'd36840, 16'd20954, 16'd21783, 16'd21307});
	test_expansion(128'h21a0c6c8b2cb966212fc6e312ad228c5, {16'd58946, 16'd40242, 16'd53779, 16'd35803, 16'd65404, 16'd51298, 16'd46098, 16'd54810, 16'd42513, 16'd37000, 16'd14755, 16'd42274, 16'd26561, 16'd3992, 16'd17282, 16'd14032, 16'd52097, 16'd32305, 16'd62928, 16'd9630, 16'd15920, 16'd15825, 16'd22033, 16'd49392, 16'd56331, 16'd53065});
	test_expansion(128'he6d1a521efc07d9cdb782d997b1fa33e, {16'd11896, 16'd43978, 16'd22660, 16'd25915, 16'd9137, 16'd4263, 16'd3317, 16'd58622, 16'd31254, 16'd54263, 16'd30879, 16'd43988, 16'd26783, 16'd10999, 16'd5331, 16'd165, 16'd665, 16'd57102, 16'd35441, 16'd28822, 16'd1557, 16'd10537, 16'd36214, 16'd17184, 16'd13435, 16'd55330});
	test_expansion(128'h700fe0090a7216edcecc94729f39eb10, {16'd18910, 16'd50072, 16'd30868, 16'd46678, 16'd54923, 16'd15362, 16'd52431, 16'd59831, 16'd4923, 16'd2452, 16'd40604, 16'd24739, 16'd34503, 16'd35649, 16'd55796, 16'd56337, 16'd3210, 16'd1855, 16'd50859, 16'd26976, 16'd45761, 16'd63725, 16'd58906, 16'd62695, 16'd13272, 16'd60964});
	test_expansion(128'h1854da363f65e178e83a923927444f6e, {16'd26850, 16'd56100, 16'd61755, 16'd44791, 16'd36862, 16'd57078, 16'd57620, 16'd46268, 16'd6576, 16'd62021, 16'd9963, 16'd46051, 16'd13438, 16'd12336, 16'd35835, 16'd33127, 16'd28337, 16'd48918, 16'd40798, 16'd33885, 16'd26815, 16'd27764, 16'd3898, 16'd16105, 16'd49799, 16'd43859});
	test_expansion(128'h447e6d8552ed56b0bf5bc86aa2fa78cc, {16'd18296, 16'd62003, 16'd57673, 16'd15883, 16'd35874, 16'd54845, 16'd65150, 16'd28846, 16'd26394, 16'd55749, 16'd48594, 16'd41360, 16'd15078, 16'd22228, 16'd64964, 16'd13138, 16'd5768, 16'd24242, 16'd36200, 16'd56069, 16'd40507, 16'd22429, 16'd48178, 16'd26032, 16'd47888, 16'd18750});
	test_expansion(128'hda2a3bbcdc8693b7a2efb2e09de5297f, {16'd20795, 16'd21082, 16'd37766, 16'd58675, 16'd53585, 16'd17511, 16'd57805, 16'd35374, 16'd36542, 16'd35566, 16'd51458, 16'd30912, 16'd33381, 16'd10926, 16'd23089, 16'd46216, 16'd43737, 16'd8980, 16'd39665, 16'd24452, 16'd40232, 16'd21493, 16'd62760, 16'd24738, 16'd27715, 16'd53614});
	test_expansion(128'hff63190a2fa3036cd9f65661cfd8cffe, {16'd19694, 16'd5155, 16'd39010, 16'd57958, 16'd60913, 16'd59571, 16'd65127, 16'd33261, 16'd49892, 16'd52713, 16'd40969, 16'd64158, 16'd253, 16'd48932, 16'd5880, 16'd33344, 16'd4978, 16'd25570, 16'd57415, 16'd44633, 16'd4674, 16'd15957, 16'd64670, 16'd58738, 16'd36185, 16'd12604});
	test_expansion(128'h4207c930e7ce44016ac412dfdcbc05cf, {16'd64763, 16'd8407, 16'd38151, 16'd56713, 16'd58184, 16'd11091, 16'd42247, 16'd4022, 16'd20564, 16'd2841, 16'd49836, 16'd31053, 16'd58978, 16'd56612, 16'd3562, 16'd58179, 16'd4253, 16'd56665, 16'd32125, 16'd61382, 16'd41685, 16'd49579, 16'd50623, 16'd46321, 16'd48759, 16'd47606});
	test_expansion(128'hb58974cacd46996d67e4ae67dcc675ab, {16'd40530, 16'd57221, 16'd36449, 16'd30813, 16'd57463, 16'd27593, 16'd59087, 16'd58565, 16'd19718, 16'd9670, 16'd17444, 16'd7082, 16'd47473, 16'd23114, 16'd640, 16'd50890, 16'd53236, 16'd61503, 16'd40506, 16'd6544, 16'd56448, 16'd20874, 16'd22769, 16'd27063, 16'd38904, 16'd59742});
	test_expansion(128'h60496bfade0feb0e57609e81b282bedc, {16'd48879, 16'd35995, 16'd12762, 16'd55547, 16'd63377, 16'd43780, 16'd21307, 16'd62005, 16'd33200, 16'd39145, 16'd20559, 16'd3156, 16'd8386, 16'd19167, 16'd37177, 16'd37023, 16'd806, 16'd58262, 16'd60896, 16'd38336, 16'd49772, 16'd7952, 16'd42703, 16'd57507, 16'd56865, 16'd55441});
	test_expansion(128'h14deac421124bfeedc55aebb95104012, {16'd8750, 16'd45784, 16'd58262, 16'd49132, 16'd26006, 16'd63398, 16'd28485, 16'd49459, 16'd5600, 16'd52612, 16'd8482, 16'd19731, 16'd22405, 16'd39083, 16'd16374, 16'd39551, 16'd13026, 16'd37075, 16'd5008, 16'd33549, 16'd28490, 16'd24804, 16'd16743, 16'd26721, 16'd34359, 16'd53050});
	test_expansion(128'he02d77884c45114f1543d358a714fd1e, {16'd21525, 16'd14388, 16'd30606, 16'd52076, 16'd29485, 16'd1327, 16'd59005, 16'd27696, 16'd13671, 16'd63697, 16'd57845, 16'd8414, 16'd41091, 16'd11989, 16'd51075, 16'd42144, 16'd29170, 16'd21854, 16'd14557, 16'd32242, 16'd21506, 16'd900, 16'd17703, 16'd61540, 16'd57677, 16'd16013});
	test_expansion(128'h25eb8e5b3c27cd58ba40e477d2fe3da0, {16'd16799, 16'd9821, 16'd35096, 16'd9861, 16'd20809, 16'd40884, 16'd26377, 16'd62070, 16'd20285, 16'd38123, 16'd33699, 16'd5259, 16'd58724, 16'd3899, 16'd42528, 16'd56245, 16'd56327, 16'd873, 16'd3325, 16'd11476, 16'd20115, 16'd14907, 16'd10729, 16'd51956, 16'd40617, 16'd47968});
	test_expansion(128'he412294edc34c23b9526973659f92106, {16'd48195, 16'd40783, 16'd58749, 16'd46394, 16'd1746, 16'd188, 16'd14198, 16'd21410, 16'd37502, 16'd60585, 16'd55736, 16'd3924, 16'd46846, 16'd19928, 16'd62862, 16'd63170, 16'd56126, 16'd7318, 16'd25389, 16'd40198, 16'd40394, 16'd51718, 16'd51124, 16'd42897, 16'd38611, 16'd27183});
	test_expansion(128'h64bb2ea5812496349a3a87cdfbdf21f0, {16'd3096, 16'd52203, 16'd12603, 16'd23772, 16'd7888, 16'd58862, 16'd3472, 16'd32489, 16'd10364, 16'd34152, 16'd30895, 16'd44113, 16'd39144, 16'd7893, 16'd16386, 16'd22492, 16'd1952, 16'd61279, 16'd5713, 16'd4797, 16'd47450, 16'd53828, 16'd30218, 16'd55423, 16'd8568, 16'd19414});
	test_expansion(128'hc1f04ca2768d1ab5cbb25e98a06255e8, {16'd54821, 16'd47863, 16'd46313, 16'd44082, 16'd9184, 16'd50106, 16'd47308, 16'd16085, 16'd63268, 16'd25099, 16'd6445, 16'd9879, 16'd39240, 16'd24701, 16'd8395, 16'd14946, 16'd34939, 16'd33647, 16'd18239, 16'd11442, 16'd24326, 16'd36096, 16'd36606, 16'd37702, 16'd49898, 16'd46289});
	test_expansion(128'h2d594e3f27a0299b0abd9f876f9daac8, {16'd43269, 16'd40190, 16'd54290, 16'd42897, 16'd22790, 16'd8359, 16'd44865, 16'd34286, 16'd4576, 16'd61982, 16'd50616, 16'd55048, 16'd27353, 16'd28202, 16'd46688, 16'd60041, 16'd31504, 16'd645, 16'd55413, 16'd58300, 16'd37179, 16'd61199, 16'd10720, 16'd57594, 16'd8429, 16'd65438});
	test_expansion(128'h9a73294625f67ab13fe24259932559ad, {16'd32294, 16'd63268, 16'd47159, 16'd37685, 16'd7778, 16'd2131, 16'd53995, 16'd32180, 16'd26366, 16'd28674, 16'd49882, 16'd33337, 16'd40340, 16'd50953, 16'd21087, 16'd53495, 16'd54565, 16'd707, 16'd55634, 16'd28314, 16'd22685, 16'd31382, 16'd63075, 16'd47008, 16'd35487, 16'd19990});
	test_expansion(128'h0851730521ea6d0dd7a6c8b8df51098b, {16'd60215, 16'd1790, 16'd9873, 16'd54504, 16'd34940, 16'd21262, 16'd24420, 16'd29138, 16'd28948, 16'd47853, 16'd45644, 16'd65320, 16'd45963, 16'd17560, 16'd49515, 16'd42753, 16'd40339, 16'd50281, 16'd63463, 16'd46905, 16'd45715, 16'd60176, 16'd31936, 16'd27524, 16'd27526, 16'd21693});
	test_expansion(128'h135e656c6e7d8f36c6638d117d69359d, {16'd56148, 16'd4422, 16'd24407, 16'd35009, 16'd6169, 16'd16892, 16'd5747, 16'd45994, 16'd58015, 16'd54710, 16'd1734, 16'd2031, 16'd55066, 16'd47606, 16'd63794, 16'd39111, 16'd22117, 16'd61162, 16'd55100, 16'd19562, 16'd34877, 16'd42586, 16'd24066, 16'd394, 16'd17851, 16'd58303});
	test_expansion(128'h8d283f0f8b29c5f857afe74455df8de6, {16'd18307, 16'd35120, 16'd55379, 16'd43194, 16'd3070, 16'd61397, 16'd11909, 16'd30820, 16'd39387, 16'd30368, 16'd48237, 16'd21564, 16'd40178, 16'd5369, 16'd23641, 16'd47180, 16'd33927, 16'd62961, 16'd36734, 16'd22014, 16'd11027, 16'd62565, 16'd43078, 16'd20437, 16'd60058, 16'd20128});
	test_expansion(128'ha16b9e5a268f3a3bea6db7a04261b2e8, {16'd27320, 16'd19280, 16'd42293, 16'd21169, 16'd64589, 16'd54464, 16'd8456, 16'd41667, 16'd26778, 16'd17096, 16'd5149, 16'd11960, 16'd13865, 16'd43334, 16'd38622, 16'd13279, 16'd60502, 16'd25597, 16'd530, 16'd31101, 16'd40566, 16'd56666, 16'd64864, 16'd6246, 16'd43770, 16'd21643});
	test_expansion(128'hea875092525f9b6d4c5540c5d827669b, {16'd18333, 16'd17816, 16'd21800, 16'd30225, 16'd19342, 16'd54419, 16'd33260, 16'd39462, 16'd45061, 16'd47971, 16'd53405, 16'd63681, 16'd20177, 16'd17305, 16'd44630, 16'd51647, 16'd50868, 16'd11241, 16'd56418, 16'd59178, 16'd53661, 16'd30667, 16'd37530, 16'd60941, 16'd1821, 16'd34470});
	test_expansion(128'h79d0b44add2a6caa7df796b1a63ac436, {16'd23279, 16'd25150, 16'd42260, 16'd19105, 16'd61389, 16'd43565, 16'd21782, 16'd12899, 16'd46894, 16'd25340, 16'd65014, 16'd28609, 16'd11583, 16'd43034, 16'd28370, 16'd53065, 16'd39999, 16'd37336, 16'd10664, 16'd32735, 16'd24709, 16'd20393, 16'd42898, 16'd46171, 16'd22878, 16'd53561});
	test_expansion(128'hf6de6b5ba42b746e540614af80dbfe7f, {16'd48366, 16'd34647, 16'd32535, 16'd4319, 16'd45469, 16'd64032, 16'd33409, 16'd32144, 16'd422, 16'd7642, 16'd46769, 16'd65274, 16'd29391, 16'd5996, 16'd59886, 16'd30132, 16'd21291, 16'd13851, 16'd57783, 16'd25135, 16'd7747, 16'd41003, 16'd58249, 16'd32899, 16'd40132, 16'd40242});
	test_expansion(128'hb3a01bd9fac69d937ae94b6670297efb, {16'd22009, 16'd21350, 16'd53555, 16'd39431, 16'd42048, 16'd28878, 16'd18505, 16'd52058, 16'd39297, 16'd26698, 16'd26525, 16'd61717, 16'd13980, 16'd9617, 16'd5919, 16'd3409, 16'd55621, 16'd1725, 16'd24800, 16'd6444, 16'd43126, 16'd12065, 16'd56340, 16'd9086, 16'd35237, 16'd28347});
	test_expansion(128'he11e3566b352e22786f4c0b743945eb8, {16'd58447, 16'd17732, 16'd25082, 16'd59977, 16'd46188, 16'd16520, 16'd41821, 16'd45388, 16'd17314, 16'd61104, 16'd4996, 16'd38308, 16'd10613, 16'd3043, 16'd52987, 16'd23132, 16'd26185, 16'd5919, 16'd47173, 16'd24457, 16'd25688, 16'd55176, 16'd38615, 16'd3596, 16'd60914, 16'd43483});
	test_expansion(128'h5ea2a4bfa8e01c845f0ad7e635f481f8, {16'd20638, 16'd47223, 16'd49204, 16'd17076, 16'd58903, 16'd45974, 16'd59577, 16'd16593, 16'd36686, 16'd38604, 16'd64909, 16'd36589, 16'd11767, 16'd51551, 16'd58812, 16'd31531, 16'd9827, 16'd63603, 16'd47873, 16'd4673, 16'd42070, 16'd4619, 16'd59847, 16'd7532, 16'd60259, 16'd53537});
	test_expansion(128'h391b72d1c2cfb983a5766f49260b2d92, {16'd22406, 16'd37875, 16'd52083, 16'd59883, 16'd52519, 16'd53320, 16'd49746, 16'd3448, 16'd41361, 16'd23761, 16'd20912, 16'd51070, 16'd54962, 16'd31926, 16'd7066, 16'd30860, 16'd17731, 16'd63019, 16'd37427, 16'd35793, 16'd44197, 16'd59044, 16'd17153, 16'd40950, 16'd16121, 16'd3797});
	test_expansion(128'h5621994827217280eb2e8259b39aa884, {16'd53858, 16'd46161, 16'd28750, 16'd47506, 16'd53429, 16'd63364, 16'd62497, 16'd13840, 16'd59648, 16'd31733, 16'd62597, 16'd52994, 16'd21987, 16'd54152, 16'd25, 16'd43063, 16'd42065, 16'd60536, 16'd35300, 16'd52645, 16'd37207, 16'd59431, 16'd27399, 16'd6208, 16'd937, 16'd3802});
	test_expansion(128'h033535e1ce7e8174595afebdd600e1fe, {16'd27704, 16'd19039, 16'd38600, 16'd46968, 16'd50432, 16'd59506, 16'd23853, 16'd25372, 16'd29404, 16'd51171, 16'd1051, 16'd64544, 16'd50511, 16'd12346, 16'd23646, 16'd17657, 16'd50297, 16'd18450, 16'd53894, 16'd44124, 16'd15416, 16'd2474, 16'd29283, 16'd46778, 16'd45873, 16'd14301});
	test_expansion(128'h87b98ccdd3ab9d398606c332dec9cd26, {16'd35279, 16'd65426, 16'd45067, 16'd30815, 16'd4081, 16'd4872, 16'd26472, 16'd33583, 16'd45809, 16'd50351, 16'd7652, 16'd60458, 16'd64213, 16'd34019, 16'd55594, 16'd40463, 16'd6914, 16'd53136, 16'd4085, 16'd6313, 16'd40407, 16'd28515, 16'd46876, 16'd14832, 16'd21601, 16'd46041});
	test_expansion(128'h1b5b1d52c66a518e0d0fccda87f65591, {16'd47079, 16'd19786, 16'd8708, 16'd56604, 16'd64613, 16'd17653, 16'd59492, 16'd38762, 16'd25508, 16'd4236, 16'd62443, 16'd24696, 16'd12655, 16'd44273, 16'd54944, 16'd63890, 16'd32358, 16'd12419, 16'd65345, 16'd2323, 16'd31138, 16'd13973, 16'd16604, 16'd27683, 16'd52524, 16'd31541});
	test_expansion(128'h0abe213568e4752a015a2cf682ee3664, {16'd33475, 16'd20725, 16'd26358, 16'd7621, 16'd61550, 16'd24635, 16'd38944, 16'd53676, 16'd31494, 16'd16149, 16'd30620, 16'd10581, 16'd5031, 16'd54591, 16'd6850, 16'd8159, 16'd12748, 16'd20202, 16'd42169, 16'd6864, 16'd52066, 16'd21546, 16'd7080, 16'd19646, 16'd59121, 16'd22751});
	test_expansion(128'h372ecc8bfd447cbdba4f81d0fa6c15d9, {16'd23640, 16'd59031, 16'd10442, 16'd27575, 16'd54129, 16'd3016, 16'd46492, 16'd9366, 16'd60295, 16'd27931, 16'd6193, 16'd24920, 16'd25804, 16'd39528, 16'd47420, 16'd16743, 16'd53468, 16'd51501, 16'd49755, 16'd9519, 16'd9387, 16'd47665, 16'd29714, 16'd57154, 16'd24116, 16'd41124});
	test_expansion(128'h7cb8f10fb730bebe01f89ea5c4a49886, {16'd28686, 16'd18090, 16'd47918, 16'd41462, 16'd25556, 16'd35269, 16'd8218, 16'd18516, 16'd7694, 16'd5722, 16'd4877, 16'd14170, 16'd29289, 16'd49588, 16'd47489, 16'd49723, 16'd10214, 16'd54703, 16'd39572, 16'd37895, 16'd34007, 16'd53681, 16'd7798, 16'd13009, 16'd64956, 16'd34207});
	test_expansion(128'ha84dfb9d34b3cb0d3a011f7ad3b308a1, {16'd13020, 16'd15108, 16'd57986, 16'd43283, 16'd5637, 16'd53379, 16'd44293, 16'd28946, 16'd27856, 16'd41197, 16'd32543, 16'd7763, 16'd28750, 16'd30323, 16'd31275, 16'd38579, 16'd57533, 16'd19649, 16'd44747, 16'd34516, 16'd47536, 16'd18342, 16'd19555, 16'd37990, 16'd46146, 16'd58759});
	test_expansion(128'h2664f156a1fce8094c13f31b9a0c72e4, {16'd10632, 16'd56055, 16'd24309, 16'd23432, 16'd25322, 16'd64447, 16'd51016, 16'd39744, 16'd34737, 16'd36865, 16'd47008, 16'd22543, 16'd15215, 16'd35713, 16'd21303, 16'd31118, 16'd60908, 16'd46114, 16'd35323, 16'd17914, 16'd44333, 16'd3435, 16'd52630, 16'd18500, 16'd64152, 16'd20432});
	test_expansion(128'h8a8ff9aba4b73b0c1a54cfef4492008a, {16'd28859, 16'd35807, 16'd35354, 16'd52125, 16'd24480, 16'd51773, 16'd429, 16'd18241, 16'd31595, 16'd57977, 16'd56197, 16'd19066, 16'd35674, 16'd50020, 16'd60686, 16'd21245, 16'd57529, 16'd10542, 16'd20730, 16'd32482, 16'd54885, 16'd28426, 16'd1744, 16'd35471, 16'd8532, 16'd33638});
	test_expansion(128'h5abc9cdcf48e76be818c1450745e62db, {16'd24267, 16'd40302, 16'd33071, 16'd18350, 16'd44048, 16'd25764, 16'd49581, 16'd64609, 16'd11676, 16'd2700, 16'd63796, 16'd10300, 16'd14388, 16'd16795, 16'd51673, 16'd16967, 16'd24021, 16'd49840, 16'd2088, 16'd23388, 16'd43362, 16'd36763, 16'd42355, 16'd31155, 16'd19030, 16'd14475});
	test_expansion(128'h47147492eca965cd8d6cb0a4aa316bc8, {16'd6442, 16'd35872, 16'd26902, 16'd65185, 16'd25450, 16'd51596, 16'd15765, 16'd59805, 16'd62500, 16'd37348, 16'd61839, 16'd25576, 16'd50455, 16'd61386, 16'd40243, 16'd55059, 16'd8658, 16'd18264, 16'd27734, 16'd43296, 16'd11721, 16'd30097, 16'd13786, 16'd26388, 16'd9083, 16'd18653});
	test_expansion(128'hccea312f0aebcd51b9672bc8f6989943, {16'd14012, 16'd1140, 16'd4902, 16'd13738, 16'd53240, 16'd9013, 16'd41995, 16'd25317, 16'd10534, 16'd33673, 16'd5564, 16'd13931, 16'd10732, 16'd10542, 16'd2933, 16'd2836, 16'd12070, 16'd40844, 16'd57824, 16'd9494, 16'd50981, 16'd52341, 16'd10307, 16'd46263, 16'd34736, 16'd37912});
	test_expansion(128'h572ee9176e802db23ffb084a289c9f00, {16'd17793, 16'd22955, 16'd37368, 16'd37617, 16'd42082, 16'd22529, 16'd20709, 16'd14647, 16'd15676, 16'd33142, 16'd62681, 16'd41256, 16'd30554, 16'd47217, 16'd39659, 16'd41912, 16'd22432, 16'd40240, 16'd57287, 16'd38984, 16'd48017, 16'd44062, 16'd48166, 16'd17918, 16'd50270, 16'd2929});
	test_expansion(128'hc96624d06dc858f4a58d18b36ff21b4b, {16'd31743, 16'd21919, 16'd24476, 16'd55970, 16'd30777, 16'd51779, 16'd4649, 16'd23802, 16'd63501, 16'd61737, 16'd64615, 16'd35078, 16'd35283, 16'd27592, 16'd30148, 16'd48687, 16'd576, 16'd16622, 16'd11264, 16'd7136, 16'd39050, 16'd60855, 16'd28774, 16'd4274, 16'd38664, 16'd50950});
	test_expansion(128'h6ac1d0e371afda9352c7238f145d11b7, {16'd55762, 16'd40028, 16'd63881, 16'd59275, 16'd47050, 16'd52418, 16'd57747, 16'd37566, 16'd10748, 16'd62355, 16'd35072, 16'd62999, 16'd15603, 16'd58962, 16'd17677, 16'd27048, 16'd45082, 16'd59782, 16'd8005, 16'd3520, 16'd65374, 16'd55040, 16'd38590, 16'd25323, 16'd24659, 16'd14609});
	test_expansion(128'hebf35f6e6f1c144cd630e167637308e7, {16'd18585, 16'd52502, 16'd56646, 16'd7851, 16'd31131, 16'd36151, 16'd14016, 16'd23669, 16'd35758, 16'd57399, 16'd47597, 16'd62005, 16'd1826, 16'd54323, 16'd769, 16'd65287, 16'd40884, 16'd42576, 16'd60544, 16'd3787, 16'd33977, 16'd54001, 16'd55901, 16'd53094, 16'd15600, 16'd24369});
	test_expansion(128'h454bc8a56325f668a6eab5c64e537398, {16'd61772, 16'd16724, 16'd30736, 16'd34803, 16'd24841, 16'd4634, 16'd19336, 16'd7019, 16'd21466, 16'd56493, 16'd50572, 16'd49797, 16'd11144, 16'd10273, 16'd8925, 16'd32942, 16'd60242, 16'd25392, 16'd25100, 16'd119, 16'd9121, 16'd47655, 16'd4101, 16'd33169, 16'd4778, 16'd53370});
	test_expansion(128'h5746339abb8e49447b60c0fcf632cec3, {16'd45590, 16'd18386, 16'd47560, 16'd4543, 16'd27541, 16'd48497, 16'd29476, 16'd49245, 16'd12050, 16'd37699, 16'd3382, 16'd18921, 16'd61483, 16'd20202, 16'd18919, 16'd4645, 16'd19884, 16'd43500, 16'd42778, 16'd38812, 16'd56915, 16'd34900, 16'd37452, 16'd27184, 16'd44357, 16'd34776});
	test_expansion(128'h85f1f9d830ece2d3c2f225751bb29f23, {16'd63491, 16'd60973, 16'd39592, 16'd18216, 16'd31906, 16'd45608, 16'd35724, 16'd63736, 16'd26965, 16'd57585, 16'd34792, 16'd36607, 16'd32997, 16'd13556, 16'd19418, 16'd101, 16'd28152, 16'd60016, 16'd42375, 16'd48130, 16'd45274, 16'd16790, 16'd33532, 16'd27570, 16'd16771, 16'd5911});
	test_expansion(128'hb49a5e52b3a7f01b235ba4f82931b1d0, {16'd51181, 16'd10819, 16'd19566, 16'd48744, 16'd60274, 16'd23128, 16'd16925, 16'd33733, 16'd10658, 16'd9681, 16'd33948, 16'd28199, 16'd56232, 16'd10805, 16'd35162, 16'd17973, 16'd29504, 16'd8075, 16'd27416, 16'd48646, 16'd30300, 16'd39363, 16'd17392, 16'd32183, 16'd61665, 16'd38891});
	test_expansion(128'hdd3c1884c82dd8c4610075d26e211276, {16'd4868, 16'd53515, 16'd28434, 16'd9186, 16'd39500, 16'd18604, 16'd25350, 16'd1525, 16'd1868, 16'd22507, 16'd12755, 16'd4671, 16'd23020, 16'd17670, 16'd17570, 16'd63255, 16'd52655, 16'd51949, 16'd51585, 16'd54883, 16'd25810, 16'd58253, 16'd32520, 16'd55958, 16'd64023, 16'd64407});
	test_expansion(128'h4673a6cf7e4f2637938f632b6309c449, {16'd7537, 16'd36292, 16'd41859, 16'd27981, 16'd36472, 16'd59213, 16'd64060, 16'd44163, 16'd27227, 16'd15072, 16'd58549, 16'd20934, 16'd11193, 16'd15601, 16'd39787, 16'd30700, 16'd37715, 16'd18852, 16'd17165, 16'd32848, 16'd59483, 16'd60145, 16'd63147, 16'd63514, 16'd23240, 16'd49529});
	test_expansion(128'h8dfb6e2f617ddfa4517ceab9516e6705, {16'd8376, 16'd11127, 16'd10154, 16'd4445, 16'd58269, 16'd21459, 16'd12983, 16'd43807, 16'd48749, 16'd4754, 16'd56334, 16'd60252, 16'd3561, 16'd10736, 16'd554, 16'd54852, 16'd46931, 16'd8757, 16'd42984, 16'd24984, 16'd61825, 16'd29026, 16'd7511, 16'd61113, 16'd39484, 16'd48756});
	test_expansion(128'he56a6aefba351e8f039ca80a148c2904, {16'd60070, 16'd32454, 16'd49655, 16'd62215, 16'd56141, 16'd4848, 16'd54620, 16'd24603, 16'd59439, 16'd3254, 16'd11194, 16'd31140, 16'd8141, 16'd59708, 16'd33510, 16'd12975, 16'd38358, 16'd61377, 16'd9163, 16'd2223, 16'd12235, 16'd24141, 16'd5448, 16'd13294, 16'd1006, 16'd48998});
	test_expansion(128'h263cdb073944b07ba6df7530b2677e81, {16'd52387, 16'd17492, 16'd44001, 16'd63207, 16'd32485, 16'd40986, 16'd22622, 16'd54772, 16'd828, 16'd2657, 16'd32267, 16'd24302, 16'd58575, 16'd19430, 16'd21408, 16'd15595, 16'd6742, 16'd35398, 16'd39513, 16'd16593, 16'd44044, 16'd16495, 16'd15986, 16'd27031, 16'd21787, 16'd28265});
	test_expansion(128'h4463a832ed159cb9bc0c07935470ada9, {16'd62761, 16'd36098, 16'd64287, 16'd18712, 16'd1964, 16'd24600, 16'd30724, 16'd49508, 16'd42496, 16'd41470, 16'd18242, 16'd19602, 16'd34341, 16'd16856, 16'd44018, 16'd14804, 16'd42860, 16'd16080, 16'd3867, 16'd61843, 16'd30228, 16'd4579, 16'd7273, 16'd11872, 16'd38206, 16'd7136});
	test_expansion(128'h6b0d6df3238d185da6bf15c6bd584c11, {16'd14307, 16'd6931, 16'd59305, 16'd56490, 16'd52685, 16'd14079, 16'd40591, 16'd62500, 16'd56784, 16'd34685, 16'd5154, 16'd16702, 16'd18533, 16'd28548, 16'd11627, 16'd56557, 16'd1714, 16'd4139, 16'd41442, 16'd12443, 16'd63015, 16'd57870, 16'd19893, 16'd55874, 16'd35551, 16'd63765});
	test_expansion(128'hf1be19a924aeb768d1f8c444efac250a, {16'd2762, 16'd40236, 16'd25121, 16'd35584, 16'd45385, 16'd7718, 16'd40797, 16'd22538, 16'd43995, 16'd49795, 16'd22279, 16'd56605, 16'd20301, 16'd2948, 16'd24095, 16'd30985, 16'd63744, 16'd933, 16'd56195, 16'd14954, 16'd33327, 16'd40523, 16'd46804, 16'd12009, 16'd33349, 16'd23853});
	test_expansion(128'h1562126ebf95e06cf2dc9584dc926034, {16'd17008, 16'd56794, 16'd52005, 16'd14188, 16'd62844, 16'd29399, 16'd32098, 16'd62630, 16'd2764, 16'd16235, 16'd20344, 16'd37240, 16'd6725, 16'd18440, 16'd21939, 16'd30643, 16'd21472, 16'd40842, 16'd53761, 16'd23579, 16'd12325, 16'd16402, 16'd32575, 16'd31719, 16'd30971, 16'd38755});
	test_expansion(128'h8f12ef2f93c1649f1c289f05c55f2baf, {16'd32670, 16'd49990, 16'd54621, 16'd162, 16'd48859, 16'd50658, 16'd31130, 16'd23575, 16'd49549, 16'd25057, 16'd21879, 16'd49237, 16'd37259, 16'd14871, 16'd59036, 16'd47950, 16'd16189, 16'd28798, 16'd39323, 16'd54204, 16'd3513, 16'd45560, 16'd15176, 16'd65325, 16'd31666, 16'd42215});
	test_expansion(128'h60cbc5b68796a17771fe95896f2618c5, {16'd51533, 16'd32624, 16'd50243, 16'd51079, 16'd61379, 16'd32236, 16'd15502, 16'd64058, 16'd63269, 16'd5966, 16'd21962, 16'd4719, 16'd12661, 16'd60533, 16'd62432, 16'd60545, 16'd58699, 16'd14989, 16'd21864, 16'd9158, 16'd14115, 16'd3202, 16'd5485, 16'd5872, 16'd37155, 16'd57007});
	test_expansion(128'h38a469decf06faceeaae20aae410de9a, {16'd55137, 16'd9528, 16'd37510, 16'd20659, 16'd7139, 16'd26361, 16'd25215, 16'd47529, 16'd23782, 16'd1768, 16'd237, 16'd32515, 16'd30726, 16'd42268, 16'd5422, 16'd55710, 16'd40882, 16'd53571, 16'd30451, 16'd8687, 16'd61678, 16'd22736, 16'd60573, 16'd19796, 16'd12514, 16'd2945});
	test_expansion(128'hec2e8b7b130122a565428485b553d852, {16'd43805, 16'd21357, 16'd53993, 16'd48975, 16'd6263, 16'd49457, 16'd36121, 16'd64304, 16'd14084, 16'd4599, 16'd3111, 16'd32481, 16'd39114, 16'd55535, 16'd63608, 16'd2286, 16'd13227, 16'd53296, 16'd43191, 16'd4699, 16'd57430, 16'd27237, 16'd5332, 16'd58635, 16'd35367, 16'd46363});
	test_expansion(128'haaef1a55a5be192f5c80011dad72174a, {16'd53365, 16'd48774, 16'd48474, 16'd10152, 16'd15503, 16'd60331, 16'd35575, 16'd41179, 16'd7189, 16'd53227, 16'd59065, 16'd6430, 16'd33093, 16'd60025, 16'd18927, 16'd34954, 16'd1521, 16'd14866, 16'd44145, 16'd2966, 16'd14191, 16'd7228, 16'd4930, 16'd29004, 16'd62121, 16'd55213});
	test_expansion(128'h9fdc4dd27006070a4f880d76b0f11b27, {16'd23936, 16'd40863, 16'd34785, 16'd37772, 16'd7743, 16'd8867, 16'd35642, 16'd16199, 16'd6090, 16'd54957, 16'd45684, 16'd42830, 16'd54501, 16'd1530, 16'd43369, 16'd58533, 16'd23927, 16'd6092, 16'd23873, 16'd4264, 16'd3284, 16'd27433, 16'd43036, 16'd12396, 16'd20545, 16'd10619});
	test_expansion(128'h99207d0392efde6941a8a9232665704f, {16'd48925, 16'd41073, 16'd25976, 16'd44196, 16'd39830, 16'd21724, 16'd38289, 16'd32235, 16'd20951, 16'd49172, 16'd54227, 16'd30103, 16'd47820, 16'd20163, 16'd53018, 16'd57737, 16'd14981, 16'd52933, 16'd3854, 16'd17982, 16'd60151, 16'd22018, 16'd51755, 16'd35734, 16'd48996, 16'd28809});
	test_expansion(128'h7389e71887309242ba9f62ba5cfa5bbf, {16'd50144, 16'd894, 16'd41701, 16'd1417, 16'd26644, 16'd23787, 16'd58135, 16'd37948, 16'd37945, 16'd530, 16'd4076, 16'd50532, 16'd52245, 16'd29741, 16'd8433, 16'd59059, 16'd33325, 16'd48109, 16'd16893, 16'd55381, 16'd2441, 16'd59822, 16'd40048, 16'd26299, 16'd20691, 16'd55447});
	test_expansion(128'h29bf80f8deb1d66a72b44e410ee82b2a, {16'd9065, 16'd1680, 16'd47910, 16'd3163, 16'd43009, 16'd2148, 16'd40946, 16'd5562, 16'd5854, 16'd36026, 16'd27549, 16'd52417, 16'd2875, 16'd38490, 16'd41361, 16'd63513, 16'd14753, 16'd16089, 16'd37031, 16'd18106, 16'd2019, 16'd16049, 16'd36240, 16'd38640, 16'd50398, 16'd10216});
	test_expansion(128'hb3d1e87166a3cbda14a67068ea58c6cd, {16'd6039, 16'd24836, 16'd59510, 16'd36642, 16'd55212, 16'd65057, 16'd43780, 16'd13767, 16'd49714, 16'd13551, 16'd26939, 16'd46573, 16'd7687, 16'd61527, 16'd61074, 16'd54086, 16'd33509, 16'd17645, 16'd58980, 16'd23192, 16'd42850, 16'd6527, 16'd24930, 16'd41292, 16'd2454, 16'd51059});
	test_expansion(128'h8992a3e0ddfeb75be62b1b38113985c7, {16'd50987, 16'd64286, 16'd44408, 16'd10956, 16'd37833, 16'd32971, 16'd15496, 16'd56272, 16'd23072, 16'd25619, 16'd23444, 16'd52001, 16'd5369, 16'd33005, 16'd38939, 16'd18379, 16'd25750, 16'd39263, 16'd60009, 16'd7961, 16'd34612, 16'd43453, 16'd37476, 16'd10512, 16'd7589, 16'd64381});
	test_expansion(128'h076f4f44624625c7bec6f66e2d2444f2, {16'd4478, 16'd12650, 16'd25552, 16'd41033, 16'd34731, 16'd38932, 16'd19157, 16'd26831, 16'd19965, 16'd27382, 16'd31189, 16'd28715, 16'd33952, 16'd44014, 16'd18143, 16'd49468, 16'd30553, 16'd773, 16'd10706, 16'd47735, 16'd6393, 16'd14333, 16'd5720, 16'd17244, 16'd12802, 16'd54824});
	test_expansion(128'h0e2044639f7b4c101f7de31a51e57ed4, {16'd44526, 16'd57575, 16'd48347, 16'd36366, 16'd52660, 16'd27518, 16'd52141, 16'd48273, 16'd11809, 16'd45924, 16'd17321, 16'd50078, 16'd61152, 16'd54978, 16'd33599, 16'd13245, 16'd46718, 16'd29576, 16'd39806, 16'd32948, 16'd51709, 16'd45894, 16'd37902, 16'd7601, 16'd34329, 16'd36019});
	test_expansion(128'h71c05811c148b2cfa792a196c195d212, {16'd19909, 16'd46667, 16'd35605, 16'd17195, 16'd48645, 16'd11834, 16'd49874, 16'd41723, 16'd2817, 16'd53839, 16'd43909, 16'd24850, 16'd57568, 16'd26455, 16'd16739, 16'd60383, 16'd54070, 16'd23633, 16'd58865, 16'd46911, 16'd63530, 16'd59521, 16'd28851, 16'd53497, 16'd16997, 16'd51735});
	test_expansion(128'h8a9ea8c98e2a9e90da3d7219675268e1, {16'd53698, 16'd21462, 16'd8325, 16'd54062, 16'd49897, 16'd10085, 16'd53527, 16'd30557, 16'd46835, 16'd41382, 16'd60852, 16'd17221, 16'd38923, 16'd2356, 16'd20739, 16'd16028, 16'd61135, 16'd3201, 16'd54412, 16'd26852, 16'd15536, 16'd43659, 16'd1011, 16'd30385, 16'd40461, 16'd56579});
	test_expansion(128'hfd825c89d097b9dc05931fb2c8fb7b62, {16'd18189, 16'd26020, 16'd13106, 16'd18796, 16'd13348, 16'd34497, 16'd16564, 16'd36956, 16'd44215, 16'd38915, 16'd64904, 16'd33026, 16'd1778, 16'd5478, 16'd52863, 16'd58074, 16'd21295, 16'd23540, 16'd62118, 16'd36957, 16'd45953, 16'd33799, 16'd13860, 16'd1320, 16'd60686, 16'd44404});
	test_expansion(128'h2a4c280f966d4eacb84b9f02387797b5, {16'd5057, 16'd59052, 16'd11526, 16'd44134, 16'd5321, 16'd54451, 16'd62600, 16'd6517, 16'd19820, 16'd21477, 16'd55179, 16'd16934, 16'd8868, 16'd16114, 16'd7420, 16'd65085, 16'd44783, 16'd59733, 16'd4916, 16'd64997, 16'd3105, 16'd26415, 16'd51128, 16'd32822, 16'd45222, 16'd24388});
	test_expansion(128'h6ce607561a71b1b2490619c5542877c6, {16'd62540, 16'd51535, 16'd12483, 16'd5156, 16'd42052, 16'd61133, 16'd1063, 16'd44829, 16'd23630, 16'd38730, 16'd50805, 16'd3248, 16'd60264, 16'd54783, 16'd25222, 16'd46283, 16'd61093, 16'd58522, 16'd63655, 16'd25140, 16'd35516, 16'd57015, 16'd11411, 16'd62492, 16'd24737, 16'd54729});
	test_expansion(128'hb8b368ecf60b3c6b7a7114896f321089, {16'd51444, 16'd13246, 16'd65418, 16'd31699, 16'd38995, 16'd52710, 16'd60035, 16'd6155, 16'd5500, 16'd38316, 16'd42679, 16'd19099, 16'd37681, 16'd60267, 16'd44660, 16'd22837, 16'd36374, 16'd27032, 16'd55091, 16'd49100, 16'd43909, 16'd18301, 16'd48435, 16'd27617, 16'd14057, 16'd58121});
	test_expansion(128'h21ce6c08780ad42344b303651b9f6aea, {16'd46527, 16'd33669, 16'd58325, 16'd51555, 16'd13312, 16'd54600, 16'd19448, 16'd20710, 16'd12018, 16'd36191, 16'd39574, 16'd29942, 16'd34568, 16'd1214, 16'd46959, 16'd18710, 16'd25618, 16'd33816, 16'd57440, 16'd996, 16'd29553, 16'd52945, 16'd37512, 16'd18437, 16'd31225, 16'd31802});
	test_expansion(128'h4a1e0923084fb6331ddda15cc48615ba, {16'd63652, 16'd57619, 16'd32972, 16'd10124, 16'd40810, 16'd338, 16'd11791, 16'd51342, 16'd30281, 16'd42533, 16'd52897, 16'd61794, 16'd38050, 16'd45426, 16'd14213, 16'd9277, 16'd45713, 16'd52911, 16'd18893, 16'd28497, 16'd60143, 16'd63057, 16'd8905, 16'd36214, 16'd51938, 16'd25196});
	test_expansion(128'h723abf344bc2095da0a7063116129efa, {16'd19078, 16'd31540, 16'd3271, 16'd38874, 16'd23085, 16'd46531, 16'd35744, 16'd30732, 16'd36030, 16'd27283, 16'd31779, 16'd55053, 16'd54919, 16'd14441, 16'd41174, 16'd45251, 16'd64869, 16'd57516, 16'd39352, 16'd64481, 16'd23673, 16'd55369, 16'd17329, 16'd31238, 16'd57642, 16'd22451});
	test_expansion(128'h76d0bd221bb744548d0babab1feb9b07, {16'd41782, 16'd40207, 16'd47697, 16'd2096, 16'd62134, 16'd815, 16'd53123, 16'd52178, 16'd7441, 16'd50893, 16'd33119, 16'd53666, 16'd31686, 16'd9937, 16'd39419, 16'd33712, 16'd63465, 16'd29490, 16'd34942, 16'd3952, 16'd23898, 16'd35844, 16'd1848, 16'd12159, 16'd16709, 16'd48419});
	test_expansion(128'h8ab11f32586335c343a4d898344c2943, {16'd42174, 16'd12921, 16'd49181, 16'd17333, 16'd47209, 16'd54252, 16'd14888, 16'd35459, 16'd38252, 16'd9230, 16'd33063, 16'd24526, 16'd32657, 16'd39221, 16'd47680, 16'd60099, 16'd49900, 16'd20028, 16'd56170, 16'd61287, 16'd15391, 16'd52095, 16'd51511, 16'd9665, 16'd31163, 16'd2326});
	test_expansion(128'h3dcd59dbcda974590f3af265c47f07ab, {16'd26320, 16'd1694, 16'd51600, 16'd23701, 16'd3833, 16'd34822, 16'd20686, 16'd4171, 16'd56599, 16'd1277, 16'd6836, 16'd49740, 16'd22572, 16'd56823, 16'd32776, 16'd62535, 16'd39147, 16'd47271, 16'd45287, 16'd39618, 16'd54404, 16'd11121, 16'd32703, 16'd57016, 16'd53793, 16'd50240});
	test_expansion(128'hf98b39fc221bc40ece1e4262db447c17, {16'd48619, 16'd58473, 16'd6268, 16'd29865, 16'd19118, 16'd14252, 16'd26378, 16'd32104, 16'd22102, 16'd15556, 16'd16603, 16'd5961, 16'd26636, 16'd54934, 16'd16431, 16'd65132, 16'd48916, 16'd2622, 16'd55609, 16'd34094, 16'd48564, 16'd13973, 16'd40741, 16'd34731, 16'd52516, 16'd6665});
	test_expansion(128'h4c739ca9ce7505bda51e293a5f635c0e, {16'd6983, 16'd44001, 16'd41330, 16'd55747, 16'd52138, 16'd13859, 16'd56451, 16'd58517, 16'd7294, 16'd41507, 16'd31265, 16'd51354, 16'd44084, 16'd51793, 16'd16076, 16'd61974, 16'd6536, 16'd20421, 16'd22660, 16'd23003, 16'd22661, 16'd10617, 16'd57861, 16'd51821, 16'd22421, 16'd39563});
	test_expansion(128'h4f7d6cc89f7216efdd0777eb308db2a4, {16'd9696, 16'd55421, 16'd24357, 16'd49162, 16'd63628, 16'd1551, 16'd48845, 16'd23462, 16'd4610, 16'd57131, 16'd7237, 16'd53877, 16'd265, 16'd49867, 16'd25044, 16'd8126, 16'd25178, 16'd24209, 16'd35598, 16'd31957, 16'd62514, 16'd62739, 16'd65227, 16'd28733, 16'd37783, 16'd39483});
	test_expansion(128'h03fa2c75925c941480943cf440e76a91, {16'd31954, 16'd63814, 16'd3849, 16'd33296, 16'd17714, 16'd11728, 16'd25, 16'd43685, 16'd22085, 16'd28498, 16'd27237, 16'd32294, 16'd65026, 16'd55057, 16'd59514, 16'd1493, 16'd18555, 16'd3349, 16'd53673, 16'd7159, 16'd7140, 16'd23676, 16'd22294, 16'd41236, 16'd42423, 16'd2704});
	test_expansion(128'h8f7315afab2a1529f99b40d8f2b2db54, {16'd63087, 16'd42109, 16'd59876, 16'd53331, 16'd22440, 16'd47327, 16'd10486, 16'd44356, 16'd8098, 16'd56684, 16'd12577, 16'd32111, 16'd1511, 16'd14145, 16'd39576, 16'd37416, 16'd24774, 16'd25626, 16'd57036, 16'd39164, 16'd11662, 16'd7502, 16'd14924, 16'd50844, 16'd14224, 16'd19986});
	test_expansion(128'hd4cba44c510dd9112cbf1d96f72ebfa7, {16'd31504, 16'd5462, 16'd33277, 16'd21810, 16'd48691, 16'd35934, 16'd42000, 16'd50950, 16'd20995, 16'd409, 16'd34648, 16'd251, 16'd36313, 16'd47093, 16'd2317, 16'd55397, 16'd26207, 16'd46324, 16'd61055, 16'd36805, 16'd47622, 16'd34931, 16'd54941, 16'd15697, 16'd52849, 16'd2412});
	test_expansion(128'h8b94a56a4cd18a28f0ac8ac6cd34c0d0, {16'd42972, 16'd12369, 16'd41950, 16'd26643, 16'd25859, 16'd27939, 16'd9994, 16'd50237, 16'd60870, 16'd39390, 16'd23653, 16'd27303, 16'd47882, 16'd5926, 16'd37726, 16'd27704, 16'd63736, 16'd20690, 16'd56321, 16'd47017, 16'd6509, 16'd9680, 16'd22499, 16'd62235, 16'd21815, 16'd25378});
	test_expansion(128'hc8d87a209a6bc51f313a69d9a3f95001, {16'd13528, 16'd54589, 16'd6543, 16'd46122, 16'd29632, 16'd4118, 16'd21301, 16'd34599, 16'd6072, 16'd51060, 16'd31588, 16'd31294, 16'd25570, 16'd62351, 16'd49254, 16'd41229, 16'd59061, 16'd1676, 16'd53836, 16'd37218, 16'd41683, 16'd9428, 16'd2039, 16'd52447, 16'd35637, 16'd64479});
	test_expansion(128'h0639b7656a1da353cf822b7bff459bd9, {16'd61614, 16'd5227, 16'd52555, 16'd49331, 16'd43296, 16'd42061, 16'd8593, 16'd1638, 16'd21150, 16'd30172, 16'd25494, 16'd61787, 16'd44273, 16'd52482, 16'd558, 16'd54927, 16'd36806, 16'd57861, 16'd18761, 16'd56223, 16'd38397, 16'd61792, 16'd50632, 16'd35640, 16'd45816, 16'd47350});
	test_expansion(128'h48bf2e1819ded879340bb17e8450aac8, {16'd3918, 16'd4896, 16'd60528, 16'd57578, 16'd25633, 16'd36513, 16'd49014, 16'd7164, 16'd33457, 16'd32114, 16'd10140, 16'd10792, 16'd62383, 16'd1532, 16'd45063, 16'd57405, 16'd30864, 16'd18455, 16'd20389, 16'd23287, 16'd47334, 16'd19869, 16'd35847, 16'd58462, 16'd7231, 16'd63313});
	test_expansion(128'h01bf732ff598c915a97c314120fb6a39, {16'd23449, 16'd39065, 16'd19528, 16'd39594, 16'd4351, 16'd55593, 16'd33480, 16'd15269, 16'd22348, 16'd24558, 16'd38372, 16'd58551, 16'd10105, 16'd11376, 16'd50742, 16'd37375, 16'd5285, 16'd39743, 16'd42589, 16'd29707, 16'd13174, 16'd60237, 16'd21903, 16'd20709, 16'd52383, 16'd43874});
	test_expansion(128'h373a3d53ccbd289358a545dc67b1192e, {16'd7376, 16'd61903, 16'd16901, 16'd57298, 16'd47664, 16'd808, 16'd5029, 16'd10720, 16'd50042, 16'd36595, 16'd27689, 16'd5312, 16'd55478, 16'd53584, 16'd64448, 16'd14000, 16'd48233, 16'd49578, 16'd4550, 16'd16650, 16'd26620, 16'd54449, 16'd42335, 16'd13847, 16'd45762, 16'd56731});
	test_expansion(128'h827344b35eb436974216b1c05de34858, {16'd28298, 16'd64479, 16'd27201, 16'd43977, 16'd30221, 16'd24198, 16'd43945, 16'd44610, 16'd16030, 16'd30304, 16'd17030, 16'd16252, 16'd32482, 16'd13150, 16'd27870, 16'd57031, 16'd3974, 16'd56739, 16'd29133, 16'd54314, 16'd42030, 16'd44918, 16'd54838, 16'd50942, 16'd42975, 16'd7121});
	test_expansion(128'hcb878c1b1f8a5629610e25996dc8913b, {16'd36332, 16'd56481, 16'd62861, 16'd33459, 16'd45544, 16'd55192, 16'd24736, 16'd24649, 16'd26587, 16'd56003, 16'd5011, 16'd59311, 16'd16830, 16'd44263, 16'd3464, 16'd11259, 16'd46555, 16'd30002, 16'd49209, 16'd138, 16'd51738, 16'd62020, 16'd25525, 16'd58163, 16'd31456, 16'd23363});
	test_expansion(128'heedbd726de9f8c974bf0513584000573, {16'd33671, 16'd16214, 16'd59203, 16'd32836, 16'd31334, 16'd22850, 16'd49057, 16'd9388, 16'd22834, 16'd47727, 16'd24507, 16'd41693, 16'd40097, 16'd15061, 16'd41351, 16'd47923, 16'd42572, 16'd32795, 16'd12342, 16'd50690, 16'd39154, 16'd13495, 16'd63605, 16'd57677, 16'd27199, 16'd40049});
	test_expansion(128'ha779fedf44d242d918cd4bcefa6d3330, {16'd39624, 16'd61701, 16'd20626, 16'd32189, 16'd39388, 16'd24456, 16'd42176, 16'd56931, 16'd29514, 16'd58633, 16'd39647, 16'd41085, 16'd8687, 16'd14451, 16'd55917, 16'd5272, 16'd28194, 16'd48749, 16'd38585, 16'd62857, 16'd52008, 16'd57946, 16'd57624, 16'd14333, 16'd57106, 16'd50285});
	test_expansion(128'hde398442f53b86c60f345f8c31631e53, {16'd50807, 16'd40922, 16'd39396, 16'd60932, 16'd23561, 16'd38297, 16'd61600, 16'd52310, 16'd51787, 16'd1496, 16'd4892, 16'd40021, 16'd6448, 16'd45701, 16'd45264, 16'd56019, 16'd22061, 16'd19807, 16'd33848, 16'd10168, 16'd17067, 16'd32356, 16'd46912, 16'd36317, 16'd55838, 16'd65332});
	test_expansion(128'h863df21a94076322f1ae4659af6469d2, {16'd49793, 16'd44790, 16'd10213, 16'd34204, 16'd8923, 16'd23178, 16'd38373, 16'd15146, 16'd64415, 16'd56406, 16'd51441, 16'd40010, 16'd6978, 16'd13010, 16'd10645, 16'd26651, 16'd8783, 16'd55500, 16'd53069, 16'd41239, 16'd1887, 16'd60094, 16'd42715, 16'd13856, 16'd24961, 16'd9386});
	test_expansion(128'hc99685aaa350e909bcec8e41064cc21d, {16'd54188, 16'd49676, 16'd36557, 16'd10170, 16'd57951, 16'd23957, 16'd22392, 16'd41687, 16'd490, 16'd28165, 16'd45398, 16'd49450, 16'd23311, 16'd32854, 16'd29684, 16'd27396, 16'd6007, 16'd7652, 16'd15003, 16'd54845, 16'd58499, 16'd29798, 16'd55769, 16'd30417, 16'd15032, 16'd65081});
	test_expansion(128'he5067c54289649b35d7e26c694eb9714, {16'd50537, 16'd1974, 16'd46728, 16'd6847, 16'd33152, 16'd45917, 16'd49809, 16'd60359, 16'd23073, 16'd23821, 16'd52189, 16'd43917, 16'd10142, 16'd27953, 16'd13681, 16'd1014, 16'd53194, 16'd6396, 16'd26413, 16'd25689, 16'd5483, 16'd60703, 16'd1888, 16'd47627, 16'd49348, 16'd41722});
	test_expansion(128'hbc81086c5e84c0c9736ee6713c645a6d, {16'd27140, 16'd27976, 16'd26555, 16'd28124, 16'd21426, 16'd17497, 16'd36894, 16'd25490, 16'd15955, 16'd24893, 16'd15607, 16'd18693, 16'd23012, 16'd4578, 16'd42051, 16'd38124, 16'd23787, 16'd17479, 16'd35063, 16'd12723, 16'd4120, 16'd27376, 16'd57095, 16'd63934, 16'd38348, 16'd50777});
	test_expansion(128'h2f3e0f080088f2f6523d9dbc24b64607, {16'd45583, 16'd31492, 16'd46592, 16'd25162, 16'd42402, 16'd43628, 16'd43711, 16'd40889, 16'd12452, 16'd52140, 16'd11520, 16'd28061, 16'd14245, 16'd51506, 16'd3503, 16'd20797, 16'd11058, 16'd7016, 16'd25130, 16'd19181, 16'd43273, 16'd50620, 16'd61452, 16'd4373, 16'd30861, 16'd5642});
	test_expansion(128'hfab94661b8befc8731a8860b86220261, {16'd56838, 16'd18670, 16'd24889, 16'd46784, 16'd61174, 16'd31890, 16'd11563, 16'd19815, 16'd3572, 16'd7558, 16'd49785, 16'd46253, 16'd21194, 16'd37498, 16'd19457, 16'd53969, 16'd41619, 16'd37065, 16'd38352, 16'd41949, 16'd39252, 16'd60525, 16'd36339, 16'd64575, 16'd22779, 16'd41217});
	test_expansion(128'h1220f9f2362a6300ada3cfd36fb5e02b, {16'd19845, 16'd60203, 16'd64004, 16'd37247, 16'd23319, 16'd45666, 16'd37097, 16'd5752, 16'd13667, 16'd27688, 16'd62982, 16'd11556, 16'd37, 16'd35031, 16'd4241, 16'd32987, 16'd58094, 16'd37101, 16'd17813, 16'd15125, 16'd3576, 16'd38447, 16'd63423, 16'd19092, 16'd13824, 16'd40226});
	test_expansion(128'h180b3a8793c30ce3160cc6ee908f5b77, {16'd60772, 16'd43324, 16'd42332, 16'd36071, 16'd37848, 16'd15361, 16'd6809, 16'd22709, 16'd11799, 16'd13314, 16'd34621, 16'd909, 16'd22214, 16'd15486, 16'd9616, 16'd37531, 16'd5808, 16'd56281, 16'd9438, 16'd7377, 16'd24823, 16'd14951, 16'd24712, 16'd33574, 16'd31646, 16'd23447});
	test_expansion(128'h943cda25ddcd50160d1946b104756274, {16'd5664, 16'd49908, 16'd30724, 16'd47959, 16'd9891, 16'd22182, 16'd56739, 16'd61753, 16'd56977, 16'd13713, 16'd39173, 16'd20393, 16'd51353, 16'd27456, 16'd18884, 16'd38683, 16'd4841, 16'd53626, 16'd63650, 16'd4593, 16'd3853, 16'd9808, 16'd45329, 16'd65079, 16'd22869, 16'd52645});
	test_expansion(128'hff9a44e8393da872f499a834d1c9ed4e, {16'd9627, 16'd26674, 16'd59259, 16'd15425, 16'd60288, 16'd32368, 16'd30168, 16'd18671, 16'd27855, 16'd62733, 16'd65344, 16'd44065, 16'd43769, 16'd12675, 16'd52297, 16'd64744, 16'd64871, 16'd42267, 16'd4710, 16'd30315, 16'd36238, 16'd7611, 16'd14249, 16'd14199, 16'd38426, 16'd29384});
	test_expansion(128'h525782193dbfaebc723bb3a16d31bf99, {16'd13775, 16'd25013, 16'd37866, 16'd47861, 16'd22012, 16'd27117, 16'd32165, 16'd39208, 16'd37154, 16'd21917, 16'd42666, 16'd47126, 16'd19343, 16'd53813, 16'd44223, 16'd17312, 16'd16268, 16'd41980, 16'd11016, 16'd7636, 16'd7074, 16'd10560, 16'd17993, 16'd29062, 16'd40027, 16'd48068});
	test_expansion(128'h595d96aa02b5c330c7e883b9dabd50a9, {16'd64536, 16'd24480, 16'd13208, 16'd2366, 16'd60880, 16'd43821, 16'd56994, 16'd1322, 16'd842, 16'd61462, 16'd16656, 16'd169, 16'd16680, 16'd19808, 16'd34788, 16'd58432, 16'd46443, 16'd53877, 16'd24871, 16'd12701, 16'd37443, 16'd51789, 16'd49232, 16'd29064, 16'd4538, 16'd23606});
	test_expansion(128'h46f7f56e2d6668828cbe921939899a17, {16'd29489, 16'd48750, 16'd27405, 16'd16517, 16'd42934, 16'd17101, 16'd26189, 16'd12416, 16'd37688, 16'd46242, 16'd64992, 16'd19707, 16'd16537, 16'd30641, 16'd47853, 16'd45245, 16'd54558, 16'd38321, 16'd21700, 16'd35185, 16'd49086, 16'd18883, 16'd10705, 16'd33748, 16'd20233, 16'd18000});
	test_expansion(128'hde7d670351c1b9b12eb846e6a3d4dc43, {16'd33586, 16'd57587, 16'd19434, 16'd54064, 16'd8097, 16'd45319, 16'd29982, 16'd23742, 16'd55462, 16'd48227, 16'd31889, 16'd54714, 16'd9267, 16'd47428, 16'd26789, 16'd58353, 16'd59077, 16'd22460, 16'd4845, 16'd60916, 16'd30005, 16'd3064, 16'd8780, 16'd56479, 16'd3116, 16'd48081});
	test_expansion(128'h959fe430e36b491323a4f1208301c56d, {16'd11159, 16'd54474, 16'd44664, 16'd17922, 16'd52022, 16'd9530, 16'd15879, 16'd41887, 16'd46889, 16'd58408, 16'd55714, 16'd41446, 16'd38848, 16'd1435, 16'd35724, 16'd56796, 16'd21631, 16'd45969, 16'd5190, 16'd10947, 16'd13962, 16'd50295, 16'd18765, 16'd20488, 16'd31854, 16'd62375});
	test_expansion(128'hefac81e553b3e7511e6416fdf50a61df, {16'd3561, 16'd60479, 16'd62945, 16'd12388, 16'd57982, 16'd34408, 16'd28471, 16'd26974, 16'd34729, 16'd48118, 16'd28020, 16'd56546, 16'd35923, 16'd33982, 16'd37732, 16'd28377, 16'd6307, 16'd7431, 16'd41686, 16'd23216, 16'd28395, 16'd29811, 16'd47735, 16'd31268, 16'd33376, 16'd13172});
	test_expansion(128'hd6057b171250c2fd7c7312da03eebfc3, {16'd49932, 16'd58201, 16'd52886, 16'd10256, 16'd44629, 16'd49491, 16'd63844, 16'd23606, 16'd33343, 16'd25398, 16'd28460, 16'd42700, 16'd2686, 16'd34157, 16'd2941, 16'd36307, 16'd16941, 16'd26337, 16'd34037, 16'd51160, 16'd54691, 16'd26045, 16'd50147, 16'd27736, 16'd23573, 16'd65535});
	test_expansion(128'h6614a901036388bfeb083545dab6deec, {16'd26146, 16'd42070, 16'd46829, 16'd6292, 16'd21728, 16'd53944, 16'd53264, 16'd47428, 16'd39405, 16'd20169, 16'd54239, 16'd54728, 16'd3561, 16'd2877, 16'd2632, 16'd22036, 16'd36187, 16'd18965, 16'd55163, 16'd61049, 16'd26829, 16'd29898, 16'd32822, 16'd50292, 16'd23420, 16'd37508});
	test_expansion(128'h15f8b10c512af489e9733d151c34ac27, {16'd53990, 16'd22566, 16'd26853, 16'd24506, 16'd54522, 16'd29352, 16'd1478, 16'd53385, 16'd62641, 16'd19964, 16'd1801, 16'd36849, 16'd31368, 16'd36230, 16'd12889, 16'd52460, 16'd27017, 16'd63011, 16'd29406, 16'd4134, 16'd61593, 16'd39515, 16'd12104, 16'd18003, 16'd41931, 16'd7545});
	test_expansion(128'h151832e0ad69d56dca4cd75958d80d5b, {16'd47321, 16'd47796, 16'd24332, 16'd36975, 16'd45464, 16'd65231, 16'd51711, 16'd55763, 16'd20177, 16'd60543, 16'd26196, 16'd28651, 16'd21932, 16'd36678, 16'd59683, 16'd51049, 16'd2527, 16'd2334, 16'd41536, 16'd37873, 16'd24227, 16'd3980, 16'd51300, 16'd43811, 16'd9105, 16'd48857});
	test_expansion(128'h3eb80795b8dbdb39b4af0d1db1fb03b2, {16'd8352, 16'd6651, 16'd44780, 16'd55598, 16'd30974, 16'd13214, 16'd29177, 16'd25671, 16'd10893, 16'd27395, 16'd7835, 16'd22900, 16'd5772, 16'd28446, 16'd16914, 16'd62639, 16'd20737, 16'd27518, 16'd14838, 16'd8616, 16'd18901, 16'd35233, 16'd15040, 16'd10144, 16'd16731, 16'd61913});
	test_expansion(128'h4e581a07401891fea3606d908c374316, {16'd57828, 16'd42472, 16'd48885, 16'd17209, 16'd56806, 16'd45415, 16'd11772, 16'd35357, 16'd27042, 16'd54112, 16'd65529, 16'd53488, 16'd6794, 16'd14729, 16'd6503, 16'd61748, 16'd17560, 16'd26604, 16'd36127, 16'd18660, 16'd49037, 16'd46178, 16'd24064, 16'd58441, 16'd11686, 16'd65298});
	test_expansion(128'h0478d058ba64a732fd1e0d595d4465b0, {16'd49375, 16'd31591, 16'd17926, 16'd1769, 16'd50850, 16'd64566, 16'd48735, 16'd46647, 16'd3338, 16'd24008, 16'd40693, 16'd24047, 16'd31357, 16'd48888, 16'd63757, 16'd62801, 16'd19583, 16'd34088, 16'd35249, 16'd59271, 16'd12256, 16'd61486, 16'd23481, 16'd24808, 16'd38719, 16'd46410});
	test_expansion(128'hc0868b2526f99e40a68eea7fd63f8dcf, {16'd42094, 16'd28569, 16'd49563, 16'd61969, 16'd47406, 16'd29293, 16'd36892, 16'd43009, 16'd38907, 16'd52982, 16'd31648, 16'd26411, 16'd37682, 16'd36333, 16'd1379, 16'd22392, 16'd8690, 16'd32979, 16'd49057, 16'd34889, 16'd33177, 16'd63195, 16'd40885, 16'd62150, 16'd54798, 16'd61170});
	test_expansion(128'h55e3e8549218908ad119c5b8520e4327, {16'd2916, 16'd20157, 16'd53392, 16'd59986, 16'd28251, 16'd31879, 16'd63874, 16'd36175, 16'd36917, 16'd50480, 16'd42934, 16'd17424, 16'd47043, 16'd48107, 16'd50268, 16'd53051, 16'd54210, 16'd8966, 16'd10827, 16'd21448, 16'd53159, 16'd49252, 16'd32252, 16'd30630, 16'd2569, 16'd11531});
	test_expansion(128'h615930282a48a535ea60640fc2e3b0ae, {16'd60880, 16'd41341, 16'd28464, 16'd61190, 16'd26286, 16'd33181, 16'd3713, 16'd21074, 16'd51258, 16'd44806, 16'd22897, 16'd25095, 16'd63902, 16'd13675, 16'd49304, 16'd54508, 16'd58505, 16'd58745, 16'd52814, 16'd27405, 16'd26274, 16'd34690, 16'd53348, 16'd18712, 16'd54852, 16'd2366});
	test_expansion(128'h3092381eafff620571eb9ebe75c5887a, {16'd51986, 16'd54691, 16'd32684, 16'd7363, 16'd64295, 16'd17692, 16'd39235, 16'd30704, 16'd58082, 16'd8657, 16'd5599, 16'd59503, 16'd46403, 16'd54589, 16'd61839, 16'd2099, 16'd11561, 16'd14147, 16'd62066, 16'd45991, 16'd25684, 16'd41519, 16'd53245, 16'd27847, 16'd60479, 16'd35987});
	test_expansion(128'ha4ae7e22b64f7195e2b576197aa145c1, {16'd61558, 16'd32569, 16'd49854, 16'd55173, 16'd32905, 16'd19999, 16'd27842, 16'd21747, 16'd56497, 16'd22336, 16'd55820, 16'd39075, 16'd15537, 16'd19808, 16'd34433, 16'd54931, 16'd51142, 16'd18701, 16'd41980, 16'd50343, 16'd19002, 16'd56798, 16'd62235, 16'd5845, 16'd41785, 16'd6322});
	test_expansion(128'h78db9ec5ab3f2a0ad82bd701e978a4f2, {16'd37669, 16'd7876, 16'd17379, 16'd40141, 16'd115, 16'd3986, 16'd60214, 16'd37430, 16'd26748, 16'd50909, 16'd3149, 16'd44421, 16'd27813, 16'd24091, 16'd54882, 16'd59253, 16'd34832, 16'd57831, 16'd29414, 16'd62681, 16'd9354, 16'd10166, 16'd35040, 16'd14866, 16'd28750, 16'd6821});
	test_expansion(128'h50f96effe7f967380f45aaaffb9f3e2c, {16'd44082, 16'd16960, 16'd46932, 16'd49810, 16'd41545, 16'd52027, 16'd49234, 16'd7952, 16'd8535, 16'd25587, 16'd37401, 16'd24037, 16'd45702, 16'd49605, 16'd59086, 16'd32895, 16'd18445, 16'd62474, 16'd55098, 16'd16135, 16'd45258, 16'd9889, 16'd42239, 16'd39679, 16'd63897, 16'd53341});
	test_expansion(128'h47500b8b5920a9efbc85ea94cfc1932f, {16'd57354, 16'd1648, 16'd40713, 16'd32701, 16'd21973, 16'd12258, 16'd44041, 16'd12934, 16'd17231, 16'd57631, 16'd62348, 16'd23096, 16'd10356, 16'd57100, 16'd39160, 16'd47004, 16'd61548, 16'd24327, 16'd44288, 16'd49667, 16'd52224, 16'd15385, 16'd49062, 16'd39740, 16'd30473, 16'd47233});
	test_expansion(128'ha139ed6be85394151bd39719a68021fb, {16'd49808, 16'd28734, 16'd31050, 16'd35772, 16'd19197, 16'd48305, 16'd64763, 16'd11126, 16'd13852, 16'd14685, 16'd49267, 16'd34962, 16'd22508, 16'd12444, 16'd27256, 16'd58832, 16'd5937, 16'd56089, 16'd32314, 16'd57264, 16'd49725, 16'd24204, 16'd52589, 16'd37911, 16'd21977, 16'd12474});
	test_expansion(128'h247c0eda7ece4f4e77ee5c31c8327b59, {16'd868, 16'd56946, 16'd60216, 16'd56545, 16'd28966, 16'd2207, 16'd20765, 16'd13398, 16'd53920, 16'd42859, 16'd8764, 16'd44595, 16'd25000, 16'd64405, 16'd2836, 16'd19652, 16'd6176, 16'd39794, 16'd46324, 16'd62786, 16'd51837, 16'd50700, 16'd40574, 16'd35991, 16'd39547, 16'd40784});
	test_expansion(128'ha0d7d3a6bd2966fccc4a26922a3b36f2, {16'd5905, 16'd4684, 16'd26121, 16'd28038, 16'd50079, 16'd12365, 16'd52905, 16'd59294, 16'd51900, 16'd13537, 16'd30931, 16'd2308, 16'd49781, 16'd10779, 16'd19441, 16'd26032, 16'd62397, 16'd60952, 16'd30812, 16'd27048, 16'd37485, 16'd33304, 16'd30882, 16'd50302, 16'd63503, 16'd14715});
	test_expansion(128'h6be2127fa13ad8d918feec4647d2a225, {16'd17616, 16'd4266, 16'd53265, 16'd6563, 16'd60584, 16'd36413, 16'd49980, 16'd37931, 16'd3450, 16'd33179, 16'd29067, 16'd50895, 16'd63008, 16'd37890, 16'd24657, 16'd45215, 16'd57573, 16'd25980, 16'd18896, 16'd53070, 16'd2686, 16'd6595, 16'd40743, 16'd51319, 16'd54602, 16'd13834});
	test_expansion(128'hde09f25c158484233583b907191820ab, {16'd51222, 16'd61807, 16'd26109, 16'd46794, 16'd52392, 16'd50127, 16'd27421, 16'd60214, 16'd15500, 16'd24158, 16'd33090, 16'd45807, 16'd10125, 16'd45006, 16'd39315, 16'd62311, 16'd43065, 16'd49380, 16'd50215, 16'd26918, 16'd26767, 16'd37744, 16'd23982, 16'd7535, 16'd9657, 16'd29311});
	test_expansion(128'h128cfc3b3ea30239dca61385a0750cc5, {16'd55857, 16'd44696, 16'd39826, 16'd52335, 16'd60215, 16'd37199, 16'd50760, 16'd60238, 16'd59841, 16'd26964, 16'd17784, 16'd7180, 16'd55202, 16'd37080, 16'd53073, 16'd12051, 16'd22760, 16'd54833, 16'd28163, 16'd51963, 16'd9241, 16'd38869, 16'd30963, 16'd22086, 16'd4924, 16'd41202});
	test_expansion(128'h61e9dec3f51d88d8bf125cbd895fe94b, {16'd55860, 16'd45813, 16'd61719, 16'd9957, 16'd61161, 16'd35563, 16'd16583, 16'd1600, 16'd58995, 16'd64854, 16'd40295, 16'd28995, 16'd21398, 16'd30259, 16'd38834, 16'd30465, 16'd43425, 16'd41071, 16'd28985, 16'd7397, 16'd15924, 16'd4527, 16'd49471, 16'd29808, 16'd1088, 16'd20046});
	test_expansion(128'h7eb339d5a38db4400de3faadc63e8735, {16'd9524, 16'd10490, 16'd56791, 16'd49794, 16'd16886, 16'd17012, 16'd8489, 16'd16724, 16'd7906, 16'd53634, 16'd40549, 16'd52931, 16'd6276, 16'd6934, 16'd38783, 16'd62285, 16'd1505, 16'd10840, 16'd64334, 16'd38054, 16'd32972, 16'd18235, 16'd20601, 16'd33480, 16'd8198, 16'd34761});
	test_expansion(128'h08a3515bd04c26ca51744927353e50d8, {16'd22740, 16'd22262, 16'd42948, 16'd32292, 16'd10191, 16'd1285, 16'd35695, 16'd33578, 16'd2494, 16'd1523, 16'd45208, 16'd63508, 16'd1191, 16'd7862, 16'd51838, 16'd24811, 16'd46237, 16'd35162, 16'd21049, 16'd28243, 16'd23275, 16'd58069, 16'd15209, 16'd53264, 16'd64272, 16'd8686});
	test_expansion(128'h95a7b52e91f73903bfa089baeda02be6, {16'd62765, 16'd21508, 16'd20181, 16'd50493, 16'd24089, 16'd37264, 16'd48174, 16'd25201, 16'd39336, 16'd26331, 16'd58509, 16'd54160, 16'd3717, 16'd41256, 16'd45739, 16'd60928, 16'd41179, 16'd30912, 16'd1385, 16'd24790, 16'd21576, 16'd15515, 16'd50760, 16'd62655, 16'd38481, 16'd7250});
	test_expansion(128'h0d63404a95bc29e358582846de69ee9b, {16'd52771, 16'd57366, 16'd10676, 16'd53765, 16'd50672, 16'd21263, 16'd32202, 16'd19908, 16'd7027, 16'd43933, 16'd9506, 16'd64669, 16'd10311, 16'd41661, 16'd32144, 16'd2157, 16'd42826, 16'd39753, 16'd6337, 16'd18469, 16'd746, 16'd34185, 16'd9857, 16'd11908, 16'd42932, 16'd13483});
	test_expansion(128'hb2e0ac6d7c216d5ada842cef9f6c4150, {16'd28914, 16'd21086, 16'd5907, 16'd45233, 16'd31694, 16'd3870, 16'd10069, 16'd63212, 16'd1066, 16'd51769, 16'd11833, 16'd36002, 16'd51088, 16'd4672, 16'd8487, 16'd47400, 16'd5679, 16'd48015, 16'd2014, 16'd1576, 16'd47883, 16'd1662, 16'd41738, 16'd29674, 16'd12497, 16'd28203});
	test_expansion(128'h8dea2887761ecb9654b4c11776c72bb8, {16'd54488, 16'd27282, 16'd33129, 16'd33747, 16'd52372, 16'd64987, 16'd47259, 16'd50480, 16'd30659, 16'd16625, 16'd10942, 16'd28216, 16'd37993, 16'd3800, 16'd10593, 16'd50166, 16'd56704, 16'd32150, 16'd13608, 16'd33667, 16'd2110, 16'd57898, 16'd13738, 16'd33434, 16'd10546, 16'd26469});
	test_expansion(128'h203aea9521d0d94a9faa8b214b082f70, {16'd35448, 16'd15298, 16'd22236, 16'd55376, 16'd21771, 16'd59156, 16'd39251, 16'd4975, 16'd42683, 16'd25374, 16'd16225, 16'd20044, 16'd54543, 16'd765, 16'd7642, 16'd19091, 16'd7669, 16'd51037, 16'd19651, 16'd6966, 16'd10946, 16'd51082, 16'd64247, 16'd24058, 16'd7317, 16'd60583});
	test_expansion(128'h878dbcb55355afaf6d17892d12ddca28, {16'd51020, 16'd17666, 16'd54658, 16'd38494, 16'd7445, 16'd3652, 16'd61255, 16'd57792, 16'd6288, 16'd7956, 16'd19839, 16'd56778, 16'd17886, 16'd43870, 16'd29590, 16'd25903, 16'd38398, 16'd27732, 16'd46657, 16'd45245, 16'd166, 16'd5239, 16'd40717, 16'd38392, 16'd8073, 16'd39077});
	test_expansion(128'h94c59a526dc178159ea7b31a40621903, {16'd25082, 16'd51307, 16'd7364, 16'd14254, 16'd62798, 16'd59976, 16'd57129, 16'd63613, 16'd49937, 16'd23731, 16'd10636, 16'd21668, 16'd14495, 16'd20386, 16'd141, 16'd41054, 16'd25443, 16'd61953, 16'd56373, 16'd35496, 16'd60302, 16'd32291, 16'd20856, 16'd11251, 16'd34961, 16'd44116});
	test_expansion(128'h2e369e53eb62020c3e4725ae6b2449a6, {16'd19148, 16'd17928, 16'd12301, 16'd61899, 16'd64812, 16'd52910, 16'd9742, 16'd18649, 16'd49671, 16'd62445, 16'd10825, 16'd50481, 16'd32496, 16'd22227, 16'd48572, 16'd52233, 16'd56760, 16'd17806, 16'd50278, 16'd44439, 16'd5167, 16'd51980, 16'd45317, 16'd27479, 16'd42587, 16'd38809});
	test_expansion(128'h72146f2dec0ed3ed039616a8f225619d, {16'd26779, 16'd65043, 16'd28243, 16'd39958, 16'd47733, 16'd8794, 16'd62995, 16'd8481, 16'd61375, 16'd29323, 16'd39480, 16'd21848, 16'd35127, 16'd2964, 16'd765, 16'd31193, 16'd43339, 16'd48641, 16'd30744, 16'd46415, 16'd5634, 16'd484, 16'd52123, 16'd18179, 16'd56376, 16'd18882});
	test_expansion(128'h8e3ef09fa01e05e8a6074ed716fb2240, {16'd19938, 16'd1689, 16'd56687, 16'd7033, 16'd51715, 16'd41100, 16'd10996, 16'd27575, 16'd14403, 16'd43346, 16'd1778, 16'd48750, 16'd41279, 16'd62167, 16'd23036, 16'd26466, 16'd42083, 16'd1688, 16'd44278, 16'd54329, 16'd33179, 16'd56840, 16'd5467, 16'd16520, 16'd14583, 16'd38051});
	test_expansion(128'h35103dd4c38f297eaa530d2f6fe85629, {16'd31082, 16'd1035, 16'd7433, 16'd10015, 16'd8148, 16'd9220, 16'd34956, 16'd39137, 16'd32229, 16'd37612, 16'd15183, 16'd44433, 16'd60568, 16'd5268, 16'd57137, 16'd24335, 16'd21997, 16'd52901, 16'd65532, 16'd43611, 16'd11894, 16'd23127, 16'd24493, 16'd33291, 16'd65079, 16'd44487});
	test_expansion(128'h6c091c623b9f0effa9cf8b7034d12788, {16'd44241, 16'd63556, 16'd47290, 16'd58697, 16'd62042, 16'd23135, 16'd31731, 16'd31178, 16'd29121, 16'd32630, 16'd48062, 16'd7937, 16'd41083, 16'd38333, 16'd17946, 16'd52961, 16'd1050, 16'd8864, 16'd45500, 16'd39413, 16'd30587, 16'd65167, 16'd61080, 16'd25459, 16'd44435, 16'd65292});
	test_expansion(128'h1c26751d20fc74ef77657a1874993b24, {16'd56675, 16'd16048, 16'd20164, 16'd2159, 16'd27790, 16'd45341, 16'd10614, 16'd58561, 16'd34203, 16'd57114, 16'd35700, 16'd52744, 16'd29518, 16'd19185, 16'd52250, 16'd44357, 16'd65076, 16'd36165, 16'd7319, 16'd18617, 16'd22769, 16'd65076, 16'd55988, 16'd40684, 16'd38521, 16'd33501});
	test_expansion(128'h376e66d05cd43fd2b804450a67b8e3ab, {16'd51136, 16'd64692, 16'd7250, 16'd57568, 16'd41020, 16'd62793, 16'd62665, 16'd51787, 16'd60970, 16'd38790, 16'd55792, 16'd10153, 16'd27434, 16'd37688, 16'd46265, 16'd12940, 16'd11339, 16'd53253, 16'd36564, 16'd50192, 16'd23994, 16'd43507, 16'd43902, 16'd14621, 16'd57472, 16'd22037});
	test_expansion(128'hf97c5b7bdbf9ef250a63795b7679895f, {16'd19137, 16'd61717, 16'd46885, 16'd59222, 16'd32814, 16'd54265, 16'd8300, 16'd28289, 16'd55593, 16'd47968, 16'd17361, 16'd1124, 16'd11839, 16'd36400, 16'd40767, 16'd45913, 16'd29514, 16'd20725, 16'd4335, 16'd19615, 16'd237, 16'd41390, 16'd1237, 16'd5911, 16'd45212, 16'd20998});
	test_expansion(128'h816aab2abba9fcaa46c0f35e1e755882, {16'd48398, 16'd22038, 16'd4340, 16'd19148, 16'd62573, 16'd25221, 16'd35566, 16'd40861, 16'd15473, 16'd30032, 16'd34516, 16'd62242, 16'd30447, 16'd60879, 16'd25046, 16'd46899, 16'd30395, 16'd17357, 16'd6460, 16'd31556, 16'd14915, 16'd32651, 16'd39553, 16'd30327, 16'd47055, 16'd59409});
	test_expansion(128'hb7874219c8b63d8c3f5ba87db600fa1a, {16'd44290, 16'd24752, 16'd32983, 16'd64319, 16'd65503, 16'd7578, 16'd14449, 16'd17357, 16'd47742, 16'd14935, 16'd52234, 16'd30500, 16'd56162, 16'd59012, 16'd28459, 16'd20495, 16'd44732, 16'd63334, 16'd38309, 16'd64811, 16'd47796, 16'd21079, 16'd54103, 16'd20557, 16'd7208, 16'd62088});
	test_expansion(128'h8b4b64102c1ae15f056f339e5717303d, {16'd13604, 16'd52630, 16'd12277, 16'd47335, 16'd7530, 16'd36656, 16'd543, 16'd168, 16'd45739, 16'd55755, 16'd957, 16'd47804, 16'd31280, 16'd29011, 16'd35393, 16'd7215, 16'd53611, 16'd63853, 16'd48816, 16'd44720, 16'd4228, 16'd65024, 16'd18276, 16'd16415, 16'd49373, 16'd19145});
	test_expansion(128'h9436dd506b1f36e966f99f2b8992a322, {16'd31671, 16'd31788, 16'd57650, 16'd23961, 16'd59451, 16'd28457, 16'd56578, 16'd8578, 16'd39576, 16'd51749, 16'd60071, 16'd57912, 16'd35899, 16'd1607, 16'd59983, 16'd45025, 16'd11878, 16'd21660, 16'd25571, 16'd17731, 16'd8018, 16'd25606, 16'd63613, 16'd22709, 16'd30163, 16'd63115});
	test_expansion(128'ha641903bded435d36a7f71f9fa8fe18f, {16'd26977, 16'd63021, 16'd1352, 16'd39162, 16'd62810, 16'd19800, 16'd25821, 16'd36229, 16'd314, 16'd55974, 16'd53934, 16'd17647, 16'd46571, 16'd49793, 16'd45867, 16'd51111, 16'd45468, 16'd45914, 16'd17959, 16'd48617, 16'd56313, 16'd48505, 16'd30312, 16'd53649, 16'd13767, 16'd26898});
	test_expansion(128'hf89db11b60b51cead475f741af1d3b0c, {16'd58402, 16'd18593, 16'd16291, 16'd29738, 16'd53837, 16'd46739, 16'd9747, 16'd5747, 16'd17252, 16'd11058, 16'd62740, 16'd49986, 16'd27704, 16'd4945, 16'd46683, 16'd25233, 16'd41172, 16'd9588, 16'd60272, 16'd11745, 16'd11881, 16'd60192, 16'd1096, 16'd32266, 16'd27372, 16'd56204});
	test_expansion(128'h5b5341be567e2bef204c5ae6060da138, {16'd611, 16'd51999, 16'd48078, 16'd31880, 16'd10487, 16'd10307, 16'd49704, 16'd62990, 16'd48922, 16'd36101, 16'd16198, 16'd51812, 16'd58604, 16'd7729, 16'd18350, 16'd23300, 16'd32864, 16'd40842, 16'd64080, 16'd28657, 16'd17299, 16'd16990, 16'd61148, 16'd5050, 16'd27629, 16'd53606});
	test_expansion(128'hfa949ef945a53f3b9cd22d3b3afe30a4, {16'd12320, 16'd32141, 16'd40203, 16'd34379, 16'd47074, 16'd40451, 16'd14588, 16'd4927, 16'd57996, 16'd59185, 16'd41719, 16'd5407, 16'd49010, 16'd59589, 16'd30566, 16'd52983, 16'd56021, 16'd51636, 16'd6624, 16'd22001, 16'd6603, 16'd60947, 16'd30969, 16'd49869, 16'd58819, 16'd14913});
	test_expansion(128'hac4e9209dab67c585ff03371fda6523e, {16'd48411, 16'd25915, 16'd34313, 16'd41606, 16'd29904, 16'd35987, 16'd41934, 16'd41897, 16'd18415, 16'd56009, 16'd65200, 16'd10890, 16'd5733, 16'd32573, 16'd23946, 16'd48183, 16'd12086, 16'd19521, 16'd52052, 16'd58702, 16'd11410, 16'd41501, 16'd21505, 16'd44306, 16'd62831, 16'd3187});
	test_expansion(128'hc0834bc6314c3bc5ad136923af48e3d2, {16'd16592, 16'd57264, 16'd44566, 16'd25012, 16'd16568, 16'd51366, 16'd13468, 16'd30444, 16'd39677, 16'd43894, 16'd16168, 16'd43187, 16'd54984, 16'd16056, 16'd63802, 16'd53281, 16'd5867, 16'd19371, 16'd19523, 16'd49261, 16'd13280, 16'd32631, 16'd3646, 16'd46503, 16'd29899, 16'd43279});
	test_expansion(128'h43d661d825c6fbe26f719d26ba079f1f, {16'd20800, 16'd19496, 16'd56492, 16'd64290, 16'd59514, 16'd3813, 16'd1596, 16'd52346, 16'd876, 16'd61997, 16'd35110, 16'd3836, 16'd4653, 16'd28017, 16'd58916, 16'd3861, 16'd23871, 16'd47222, 16'd18184, 16'd29854, 16'd45793, 16'd54896, 16'd9969, 16'd7950, 16'd27026, 16'd13444});
	test_expansion(128'h4db179dd0fc354074ef16cc15d646696, {16'd9749, 16'd55964, 16'd61946, 16'd13271, 16'd32397, 16'd49617, 16'd11405, 16'd34298, 16'd53792, 16'd17005, 16'd31231, 16'd11353, 16'd26273, 16'd6592, 16'd15895, 16'd2381, 16'd7623, 16'd57654, 16'd57621, 16'd61015, 16'd48299, 16'd59690, 16'd3807, 16'd58946, 16'd48141, 16'd27745});
	test_expansion(128'hb849f86222dba8d8147e111895914e9a, {16'd51813, 16'd14146, 16'd15283, 16'd48849, 16'd17102, 16'd19929, 16'd50192, 16'd19184, 16'd23694, 16'd64962, 16'd9816, 16'd49828, 16'd61344, 16'd31552, 16'd61331, 16'd27147, 16'd30862, 16'd14243, 16'd41868, 16'd34278, 16'd59486, 16'd29081, 16'd7257, 16'd9821, 16'd15215, 16'd37173});
	test_expansion(128'h06d8282c65107081270b1e9f49a468d9, {16'd13438, 16'd39766, 16'd24653, 16'd65466, 16'd24840, 16'd43027, 16'd35354, 16'd40895, 16'd20161, 16'd11176, 16'd20978, 16'd28007, 16'd44873, 16'd51094, 16'd17114, 16'd48555, 16'd32018, 16'd16013, 16'd10758, 16'd55082, 16'd17331, 16'd20323, 16'd28772, 16'd34379, 16'd30327, 16'd26275});
	test_expansion(128'h0e419443098cc0fc00402fae87e7d0c1, {16'd10035, 16'd43718, 16'd23872, 16'd32841, 16'd57240, 16'd64716, 16'd6383, 16'd9140, 16'd29699, 16'd9358, 16'd15018, 16'd12662, 16'd6784, 16'd7885, 16'd15970, 16'd60260, 16'd12368, 16'd38268, 16'd32191, 16'd15459, 16'd25892, 16'd56628, 16'd57971, 16'd24772, 16'd44379, 16'd54727});
	test_expansion(128'h44abf029e964a52df7ddfc7e4a3c0abb, {16'd4064, 16'd33051, 16'd10, 16'd49461, 16'd13632, 16'd59462, 16'd27623, 16'd7179, 16'd40583, 16'd45609, 16'd38447, 16'd26561, 16'd2271, 16'd52683, 16'd49699, 16'd40976, 16'd36460, 16'd11492, 16'd59120, 16'd54211, 16'd39615, 16'd11290, 16'd19305, 16'd61430, 16'd50938, 16'd38143});
	test_expansion(128'hac4646641c45a55b395730cd111d0b2e, {16'd25973, 16'd60848, 16'd16798, 16'd26507, 16'd14897, 16'd51112, 16'd24136, 16'd16953, 16'd6319, 16'd56288, 16'd35571, 16'd37953, 16'd15691, 16'd38774, 16'd11581, 16'd34618, 16'd48368, 16'd54963, 16'd53984, 16'd48140, 16'd55454, 16'd10980, 16'd15801, 16'd43614, 16'd43605, 16'd35548});
	test_expansion(128'hce5c7e6035d4475a9f98532519853db7, {16'd41344, 16'd20435, 16'd13979, 16'd60854, 16'd8546, 16'd49293, 16'd7365, 16'd61660, 16'd50436, 16'd56266, 16'd11216, 16'd51328, 16'd56437, 16'd36266, 16'd40274, 16'd42881, 16'd20792, 16'd24935, 16'd56732, 16'd13219, 16'd35313, 16'd49782, 16'd11879, 16'd18428, 16'd458, 16'd49701});
	test_expansion(128'h222f37fe7df1034f208e2bf801b70b29, {16'd34448, 16'd27213, 16'd49643, 16'd26893, 16'd7754, 16'd43560, 16'd48379, 16'd60484, 16'd62468, 16'd7667, 16'd17159, 16'd62413, 16'd32936, 16'd28763, 16'd12649, 16'd37751, 16'd41432, 16'd25551, 16'd4764, 16'd15257, 16'd41759, 16'd54814, 16'd53786, 16'd56818, 16'd57574, 16'd9568});
	test_expansion(128'hf07c2dfc80f71a3b88b63136339970f1, {16'd45327, 16'd45236, 16'd48175, 16'd18490, 16'd64557, 16'd24809, 16'd27823, 16'd3052, 16'd24685, 16'd12598, 16'd61632, 16'd49408, 16'd12211, 16'd46994, 16'd54877, 16'd64287, 16'd10125, 16'd33060, 16'd43667, 16'd55251, 16'd30910, 16'd34564, 16'd57620, 16'd47578, 16'd6889, 16'd62361});
	test_expansion(128'h1a3360c5cd1a6930db727715d3d3e28c, {16'd62180, 16'd35879, 16'd7737, 16'd14075, 16'd32962, 16'd41748, 16'd14184, 16'd25660, 16'd42078, 16'd24463, 16'd17387, 16'd34619, 16'd16382, 16'd33667, 16'd45410, 16'd58916, 16'd47833, 16'd51203, 16'd44624, 16'd25268, 16'd58959, 16'd34341, 16'd39267, 16'd33836, 16'd55488, 16'd22564});
	test_expansion(128'hf9b72e430e62415343352c6ac218f53e, {16'd27427, 16'd22773, 16'd27611, 16'd17539, 16'd56221, 16'd35078, 16'd54216, 16'd55057, 16'd14703, 16'd75, 16'd14631, 16'd28704, 16'd59917, 16'd11273, 16'd42579, 16'd33444, 16'd38118, 16'd39987, 16'd39596, 16'd3048, 16'd4126, 16'd60422, 16'd44124, 16'd34007, 16'd52528, 16'd53392});
	test_expansion(128'h0db73ebed67d2e863b702b7444948b34, {16'd45323, 16'd60828, 16'd60933, 16'd48383, 16'd54776, 16'd29138, 16'd64894, 16'd19817, 16'd37784, 16'd29153, 16'd40090, 16'd28177, 16'd29266, 16'd15323, 16'd34117, 16'd46652, 16'd12267, 16'd40530, 16'd65464, 16'd45610, 16'd30662, 16'd12189, 16'd50903, 16'd20356, 16'd32030, 16'd22009});
	test_expansion(128'h6515d5b9f4e28f2fab42e353bd31c184, {16'd12895, 16'd19152, 16'd764, 16'd33602, 16'd18753, 16'd9490, 16'd60291, 16'd236, 16'd16696, 16'd12540, 16'd1259, 16'd27282, 16'd55520, 16'd48744, 16'd36407, 16'd27633, 16'd16930, 16'd21343, 16'd48993, 16'd11317, 16'd30102, 16'd8784, 16'd42421, 16'd7151, 16'd2465, 16'd37354});
	test_expansion(128'hefe65c356c70d4b3a63eeaa2df56f2cd, {16'd57076, 16'd45569, 16'd14544, 16'd51393, 16'd7381, 16'd44286, 16'd56175, 16'd36258, 16'd59286, 16'd22982, 16'd55639, 16'd30286, 16'd63693, 16'd9149, 16'd3988, 16'd24219, 16'd24890, 16'd44741, 16'd64937, 16'd58318, 16'd1188, 16'd39800, 16'd1883, 16'd55245, 16'd43212, 16'd37473});
	test_expansion(128'hc5ccf8dd60b1695f9f6c4db7bdf5163a, {16'd47911, 16'd44012, 16'd33330, 16'd13364, 16'd64747, 16'd52537, 16'd50139, 16'd38883, 16'd29108, 16'd46506, 16'd3154, 16'd6653, 16'd1572, 16'd12187, 16'd9989, 16'd9284, 16'd15082, 16'd32633, 16'd18716, 16'd59334, 16'd49863, 16'd63755, 16'd46804, 16'd57172, 16'd15177, 16'd31032});
	test_expansion(128'he3e67c30c183d34120eb36abd3c8c975, {16'd670, 16'd30424, 16'd25621, 16'd5166, 16'd27262, 16'd51010, 16'd41976, 16'd46577, 16'd25696, 16'd13531, 16'd41662, 16'd25765, 16'd19616, 16'd51967, 16'd59596, 16'd65315, 16'd24305, 16'd7195, 16'd51281, 16'd38295, 16'd46913, 16'd62817, 16'd41892, 16'd14778, 16'd35311, 16'd34054});
	test_expansion(128'h8a02d3cf3fe5d25484568fd8e7958796, {16'd49485, 16'd58214, 16'd14407, 16'd5055, 16'd61180, 16'd8326, 16'd53222, 16'd25444, 16'd14938, 16'd1569, 16'd10442, 16'd52439, 16'd35367, 16'd48486, 16'd16138, 16'd47535, 16'd48400, 16'd29343, 16'd37594, 16'd28594, 16'd14335, 16'd2483, 16'd41552, 16'd3825, 16'd40968, 16'd40649});
	test_expansion(128'h58718b4b04a0bf6aa18514faccae1207, {16'd65310, 16'd21890, 16'd49491, 16'd39030, 16'd28368, 16'd58244, 16'd39802, 16'd63079, 16'd59864, 16'd33020, 16'd9300, 16'd32399, 16'd15205, 16'd31345, 16'd6728, 16'd51599, 16'd10242, 16'd34193, 16'd62407, 16'd53511, 16'd8472, 16'd48224, 16'd64013, 16'd37256, 16'd26617, 16'd22626});
	test_expansion(128'h3968c9aaa01acb0e30cfc1c8721534cb, {16'd18964, 16'd44827, 16'd673, 16'd27182, 16'd12523, 16'd31618, 16'd1352, 16'd56020, 16'd9689, 16'd54371, 16'd54605, 16'd41178, 16'd25347, 16'd42738, 16'd27329, 16'd62568, 16'd42865, 16'd18425, 16'd57459, 16'd16734, 16'd5500, 16'd44780, 16'd62848, 16'd13792, 16'd63993, 16'd34021});
	test_expansion(128'hbbc09699b5bf03710bdb6c81e0b4901a, {16'd60251, 16'd51107, 16'd26447, 16'd42711, 16'd56328, 16'd29551, 16'd10122, 16'd2191, 16'd27462, 16'd57837, 16'd62125, 16'd46711, 16'd41842, 16'd8648, 16'd14230, 16'd56842, 16'd1814, 16'd46263, 16'd29750, 16'd61672, 16'd30971, 16'd48520, 16'd3913, 16'd52516, 16'd40393, 16'd32385});
	test_expansion(128'h9da81d827f631b5f0ec9932477a19dbc, {16'd28219, 16'd33639, 16'd4488, 16'd63313, 16'd58268, 16'd26273, 16'd40281, 16'd32721, 16'd57640, 16'd63612, 16'd31928, 16'd30051, 16'd23201, 16'd1583, 16'd26508, 16'd46371, 16'd23914, 16'd50880, 16'd62174, 16'd56409, 16'd12836, 16'd40177, 16'd56360, 16'd38791, 16'd14431, 16'd51333});
	test_expansion(128'h1bf1aaa3b10f0587ba3d7d6a02f94e44, {16'd43240, 16'd2000, 16'd53893, 16'd51814, 16'd45054, 16'd21532, 16'd20664, 16'd16645, 16'd46685, 16'd54135, 16'd41887, 16'd41233, 16'd60565, 16'd43120, 16'd18385, 16'd53482, 16'd29165, 16'd31774, 16'd1361, 16'd30442, 16'd16491, 16'd24446, 16'd46719, 16'd59621, 16'd35498, 16'd28877});
	test_expansion(128'hc779bcc0e90728d87b25b3ac466a5b62, {16'd37007, 16'd48386, 16'd25482, 16'd45898, 16'd53461, 16'd46551, 16'd37017, 16'd13862, 16'd21368, 16'd25828, 16'd31668, 16'd43648, 16'd21339, 16'd50886, 16'd42892, 16'd8058, 16'd10577, 16'd26892, 16'd21676, 16'd60974, 16'd33603, 16'd43960, 16'd4928, 16'd46754, 16'd47837, 16'd5193});
	test_expansion(128'h3d73c2e772d8ef0e43ec90be127d89b6, {16'd61462, 16'd52272, 16'd27287, 16'd37416, 16'd37435, 16'd36606, 16'd7151, 16'd25872, 16'd48115, 16'd49554, 16'd22438, 16'd446, 16'd43990, 16'd13988, 16'd49654, 16'd3253, 16'd48459, 16'd57808, 16'd48372, 16'd7510, 16'd63308, 16'd29580, 16'd44980, 16'd24073, 16'd26878, 16'd1949});
	test_expansion(128'hcbc16bd885732fdbec801b71effe8ede, {16'd53666, 16'd21545, 16'd41522, 16'd28456, 16'd60793, 16'd32301, 16'd8867, 16'd25036, 16'd2344, 16'd48991, 16'd15036, 16'd39475, 16'd8796, 16'd5164, 16'd40701, 16'd41618, 16'd29971, 16'd16242, 16'd32896, 16'd10217, 16'd42719, 16'd44371, 16'd8657, 16'd30759, 16'd20840, 16'd24151});
	test_expansion(128'hd12d7cb69351ca03e02dd6796578883d, {16'd34916, 16'd6473, 16'd55129, 16'd56427, 16'd44308, 16'd65267, 16'd16607, 16'd12027, 16'd6789, 16'd40336, 16'd15812, 16'd42301, 16'd37599, 16'd37194, 16'd25838, 16'd61877, 16'd52056, 16'd36615, 16'd61913, 16'd38019, 16'd25486, 16'd52000, 16'd1918, 16'd43398, 16'd7571, 16'd63022});
	test_expansion(128'h55634de8674db51643b763e07823ba12, {16'd65054, 16'd27269, 16'd41602, 16'd19321, 16'd7258, 16'd9710, 16'd56245, 16'd61348, 16'd44311, 16'd7370, 16'd16418, 16'd57151, 16'd8943, 16'd48197, 16'd61381, 16'd56845, 16'd10176, 16'd28314, 16'd26193, 16'd27521, 16'd26995, 16'd11193, 16'd65167, 16'd46660, 16'd63910, 16'd10087});
	test_expansion(128'he8e59c59bd207d119f7c3581e5eaad80, {16'd64576, 16'd35696, 16'd37112, 16'd6444, 16'd16981, 16'd51033, 16'd994, 16'd2241, 16'd16802, 16'd10921, 16'd61758, 16'd60683, 16'd37666, 16'd38969, 16'd30683, 16'd59165, 16'd16064, 16'd5009, 16'd35499, 16'd51470, 16'd40830, 16'd63706, 16'd29138, 16'd6716, 16'd61688, 16'd38835});
	test_expansion(128'h1e02a59c9ee76ea2d73b6e141d0a479d, {16'd12443, 16'd6658, 16'd5328, 16'd28178, 16'd36270, 16'd52980, 16'd29015, 16'd50945, 16'd30235, 16'd63785, 16'd62587, 16'd41509, 16'd12396, 16'd56011, 16'd43925, 16'd1233, 16'd1313, 16'd9249, 16'd37227, 16'd9600, 16'd62790, 16'd1908, 16'd44222, 16'd49355, 16'd53969, 16'd7999});
	test_expansion(128'h18a258c6f8b314c6955ddabb5380a93a, {16'd58651, 16'd4190, 16'd47459, 16'd10598, 16'd56638, 16'd41278, 16'd30481, 16'd40154, 16'd61246, 16'd44013, 16'd10073, 16'd6311, 16'd25245, 16'd201, 16'd37661, 16'd10285, 16'd23864, 16'd20847, 16'd60410, 16'd62404, 16'd32308, 16'd55727, 16'd2061, 16'd34867, 16'd42118, 16'd64371});
	test_expansion(128'h1ace80d856544677a6395b272c19a72e, {16'd2642, 16'd15703, 16'd21933, 16'd13311, 16'd26787, 16'd45770, 16'd47617, 16'd3918, 16'd33504, 16'd19355, 16'd51793, 16'd30703, 16'd22466, 16'd34489, 16'd39403, 16'd13899, 16'd3389, 16'd5924, 16'd23608, 16'd2227, 16'd58958, 16'd46399, 16'd51487, 16'd57156, 16'd29059, 16'd57363});
	test_expansion(128'h5d0f06fab1d9aad04ce7bdb4ce7920dd, {16'd51205, 16'd29703, 16'd15646, 16'd65337, 16'd25420, 16'd47087, 16'd51249, 16'd46218, 16'd43719, 16'd56021, 16'd38208, 16'd9451, 16'd33541, 16'd17142, 16'd13469, 16'd20378, 16'd2215, 16'd8007, 16'd56630, 16'd21888, 16'd22458, 16'd4440, 16'd32592, 16'd41773, 16'd23057, 16'd33325});
	test_expansion(128'h99e38d23d09f215b50e8284a2d0f5413, {16'd16767, 16'd62121, 16'd60204, 16'd61375, 16'd11865, 16'd9109, 16'd56132, 16'd53784, 16'd33689, 16'd35416, 16'd14035, 16'd24689, 16'd16670, 16'd64696, 16'd35822, 16'd20232, 16'd39341, 16'd28923, 16'd40257, 16'd10490, 16'd1516, 16'd40835, 16'd55248, 16'd50718, 16'd54139, 16'd8511});
	test_expansion(128'hc26b5d4b053cc90b5b5203ec054406f4, {16'd23896, 16'd56359, 16'd53777, 16'd37750, 16'd47942, 16'd38564, 16'd3131, 16'd46375, 16'd8441, 16'd26464, 16'd33270, 16'd7843, 16'd55535, 16'd18287, 16'd16563, 16'd44857, 16'd5779, 16'd47903, 16'd34973, 16'd43370, 16'd59638, 16'd19515, 16'd39452, 16'd36947, 16'd11365, 16'd38512});
	test_expansion(128'hc35598e4dbaf6b6076743e5482f0505e, {16'd6205, 16'd6294, 16'd54404, 16'd32933, 16'd18847, 16'd18178, 16'd65172, 16'd11527, 16'd35228, 16'd19348, 16'd10534, 16'd53922, 16'd20122, 16'd20960, 16'd6746, 16'd48015, 16'd60195, 16'd9766, 16'd5544, 16'd50719, 16'd38325, 16'd44243, 16'd52111, 16'd23357, 16'd65042, 16'd8640});
	test_expansion(128'hbbd7b8e9deca6ebc89193bbb0f6d811e, {16'd12434, 16'd27946, 16'd12795, 16'd6228, 16'd49751, 16'd42445, 16'd27667, 16'd1387, 16'd11949, 16'd57780, 16'd11152, 16'd58827, 16'd37904, 16'd8049, 16'd62205, 16'd56062, 16'd7001, 16'd62983, 16'd47098, 16'd24658, 16'd41857, 16'd43006, 16'd56377, 16'd19003, 16'd15239, 16'd30588});
	test_expansion(128'h2a02292ed9de2c61a9a9d861357b23c0, {16'd2658, 16'd23346, 16'd29847, 16'd49798, 16'd30486, 16'd37368, 16'd1153, 16'd32506, 16'd978, 16'd62271, 16'd31514, 16'd26070, 16'd58476, 16'd55767, 16'd45490, 16'd19162, 16'd17407, 16'd37574, 16'd4078, 16'd35598, 16'd45465, 16'd34932, 16'd43628, 16'd25216, 16'd11775, 16'd65508});
	test_expansion(128'h3972cd09fb0708be603585c3c3248a60, {16'd29402, 16'd58662, 16'd62377, 16'd6658, 16'd47633, 16'd48949, 16'd32189, 16'd33875, 16'd19587, 16'd16781, 16'd22880, 16'd43927, 16'd14070, 16'd8234, 16'd37411, 16'd45306, 16'd40991, 16'd805, 16'd15781, 16'd59061, 16'd18719, 16'd2799, 16'd8556, 16'd44436, 16'd59375, 16'd4322});
	test_expansion(128'h99beda141de502761df26d4a6daad115, {16'd28026, 16'd46807, 16'd12973, 16'd25923, 16'd22120, 16'd4029, 16'd65526, 16'd8261, 16'd446, 16'd59481, 16'd9766, 16'd61734, 16'd2242, 16'd55965, 16'd20968, 16'd23909, 16'd49913, 16'd24978, 16'd50185, 16'd20308, 16'd23833, 16'd14099, 16'd4643, 16'd32823, 16'd54863, 16'd45006});
	test_expansion(128'h5f3f49f2d3488af6ae28897493b79a61, {16'd18912, 16'd3221, 16'd22513, 16'd62993, 16'd54579, 16'd45921, 16'd18366, 16'd41575, 16'd29648, 16'd55881, 16'd16881, 16'd5258, 16'd11915, 16'd6628, 16'd22016, 16'd18639, 16'd54207, 16'd13399, 16'd54606, 16'd50170, 16'd12213, 16'd11497, 16'd5966, 16'd55932, 16'd16434, 16'd58375});
	test_expansion(128'hf5affb6e8999c68c551b35a714f78631, {16'd45661, 16'd62653, 16'd34035, 16'd29828, 16'd36167, 16'd53817, 16'd55343, 16'd21411, 16'd20465, 16'd3420, 16'd19258, 16'd2063, 16'd814, 16'd13401, 16'd32346, 16'd5307, 16'd15554, 16'd13050, 16'd20440, 16'd9554, 16'd31071, 16'd17511, 16'd23077, 16'd9781, 16'd53212, 16'd4952});
	test_expansion(128'h3eca8ce17123edd4ea2ba51eaf754f73, {16'd30668, 16'd32421, 16'd62832, 16'd16981, 16'd47462, 16'd32915, 16'd59710, 16'd21131, 16'd25743, 16'd46945, 16'd2977, 16'd21001, 16'd21568, 16'd3791, 16'd23359, 16'd27586, 16'd19662, 16'd43040, 16'd42682, 16'd41742, 16'd5031, 16'd50835, 16'd54547, 16'd61577, 16'd61241, 16'd10358});
	test_expansion(128'h3192b908ef8f6ec37a69bc33224e3e38, {16'd23850, 16'd8925, 16'd37432, 16'd58040, 16'd1581, 16'd63103, 16'd31001, 16'd16408, 16'd16446, 16'd182, 16'd40303, 16'd55500, 16'd25550, 16'd47020, 16'd28775, 16'd16764, 16'd25088, 16'd12364, 16'd25824, 16'd17130, 16'd1815, 16'd23164, 16'd6529, 16'd60539, 16'd20159, 16'd9568});
	test_expansion(128'h0b0e2f5c99d513a02ee4da9747b2a5c4, {16'd6479, 16'd43972, 16'd22118, 16'd24966, 16'd1757, 16'd52639, 16'd42520, 16'd2732, 16'd52495, 16'd20201, 16'd17435, 16'd59664, 16'd46341, 16'd41807, 16'd18295, 16'd11137, 16'd31731, 16'd48878, 16'd51703, 16'd54507, 16'd49971, 16'd22386, 16'd7755, 16'd50226, 16'd9687, 16'd9778});
	test_expansion(128'h9ae216c85ccb778f9396b76e0cf89f4e, {16'd29253, 16'd56381, 16'd38929, 16'd62875, 16'd14377, 16'd49483, 16'd63140, 16'd21779, 16'd18325, 16'd38824, 16'd6007, 16'd35279, 16'd53253, 16'd646, 16'd57008, 16'd36152, 16'd42925, 16'd49687, 16'd39412, 16'd14863, 16'd37550, 16'd4895, 16'd20921, 16'd63825, 16'd46005, 16'd46840});
	test_expansion(128'h5aa6ac15503fa107f6038a99d5035297, {16'd60643, 16'd8775, 16'd20670, 16'd12962, 16'd19179, 16'd25537, 16'd36231, 16'd63259, 16'd40636, 16'd15733, 16'd42198, 16'd39128, 16'd63809, 16'd35734, 16'd27014, 16'd60970, 16'd30264, 16'd4602, 16'd16924, 16'd40014, 16'd45130, 16'd19093, 16'd21422, 16'd5724, 16'd3283, 16'd1394});
	test_expansion(128'h7c7ca6c11bcfd1a52f7d857572f79a79, {16'd22564, 16'd15893, 16'd62380, 16'd14814, 16'd38057, 16'd5221, 16'd57300, 16'd56742, 16'd9364, 16'd51202, 16'd7930, 16'd10700, 16'd39642, 16'd59057, 16'd14659, 16'd26675, 16'd51907, 16'd41801, 16'd10938, 16'd48606, 16'd60368, 16'd15981, 16'd27154, 16'd6523, 16'd33558, 16'd40877});
	test_expansion(128'ha888362f7511671028d34a773fb4a74f, {16'd8619, 16'd10315, 16'd9733, 16'd41855, 16'd65524, 16'd15290, 16'd52779, 16'd40485, 16'd22393, 16'd58705, 16'd7501, 16'd3707, 16'd11759, 16'd48062, 16'd55371, 16'd5671, 16'd39946, 16'd18656, 16'd13914, 16'd41881, 16'd32589, 16'd53368, 16'd33067, 16'd58186, 16'd14966, 16'd16268});
	test_expansion(128'h362ef7aa3ca30ef43b4bf1107347ddcc, {16'd45460, 16'd38535, 16'd65111, 16'd34605, 16'd33756, 16'd28685, 16'd4403, 16'd34174, 16'd48359, 16'd32912, 16'd62478, 16'd37739, 16'd13271, 16'd40579, 16'd30662, 16'd11018, 16'd2740, 16'd34765, 16'd22493, 16'd60492, 16'd19949, 16'd25460, 16'd20730, 16'd55688, 16'd37324, 16'd20442});
	test_expansion(128'h7838562a7a29ccc05a572cd54e22bd41, {16'd26751, 16'd8123, 16'd28837, 16'd436, 16'd2651, 16'd46372, 16'd25545, 16'd16212, 16'd3629, 16'd50271, 16'd14906, 16'd60688, 16'd48654, 16'd53991, 16'd59298, 16'd27204, 16'd4773, 16'd41574, 16'd8619, 16'd28550, 16'd33425, 16'd37681, 16'd27841, 16'd18932, 16'd35097, 16'd2280});
	test_expansion(128'h9fbb970a1ab4d260575652d0083e8c77, {16'd20896, 16'd36797, 16'd42896, 16'd36786, 16'd56200, 16'd43816, 16'd34049, 16'd20633, 16'd54136, 16'd24460, 16'd41465, 16'd41867, 16'd11261, 16'd33382, 16'd14747, 16'd52633, 16'd16285, 16'd8867, 16'd5103, 16'd52878, 16'd55723, 16'd26879, 16'd2490, 16'd53622, 16'd11070, 16'd61738});
	test_expansion(128'h795c3e8182103026ffc0708d81eee4c2, {16'd7120, 16'd53436, 16'd35084, 16'd52798, 16'd9053, 16'd35825, 16'd40295, 16'd43012, 16'd23123, 16'd12887, 16'd11336, 16'd11288, 16'd47978, 16'd21377, 16'd36422, 16'd19200, 16'd31565, 16'd52805, 16'd20628, 16'd55079, 16'd20130, 16'd16226, 16'd26156, 16'd19947, 16'd10854, 16'd64593});
	test_expansion(128'h4d079267c72cbac200ebcef40be46eec, {16'd38814, 16'd2057, 16'd60269, 16'd29082, 16'd36961, 16'd41224, 16'd39748, 16'd3178, 16'd6802, 16'd5664, 16'd38628, 16'd29414, 16'd55923, 16'd29878, 16'd45095, 16'd57431, 16'd42228, 16'd12577, 16'd53597, 16'd17153, 16'd65219, 16'd37471, 16'd22150, 16'd43845, 16'd23422, 16'd51228});
	test_expansion(128'hdb198131df9ef5bd25ab07d18e6bfa0d, {16'd63254, 16'd59791, 16'd30350, 16'd18137, 16'd15997, 16'd53561, 16'd8146, 16'd8366, 16'd30527, 16'd10596, 16'd32906, 16'd32402, 16'd8253, 16'd3336, 16'd58713, 16'd23665, 16'd23697, 16'd53672, 16'd48316, 16'd15508, 16'd45027, 16'd33039, 16'd3712, 16'd29554, 16'd18989, 16'd57938});
	test_expansion(128'h1286e5dd057739eabfa011b9e426e37b, {16'd41003, 16'd24096, 16'd37408, 16'd34096, 16'd24792, 16'd35514, 16'd63523, 16'd43240, 16'd10084, 16'd28880, 16'd3989, 16'd47893, 16'd4244, 16'd56131, 16'd31143, 16'd20469, 16'd24750, 16'd19244, 16'd36062, 16'd9134, 16'd13586, 16'd22894, 16'd28736, 16'd54908, 16'd45293, 16'd31988});
	test_expansion(128'hb745d65c65597727dd50058793b0dc9e, {16'd19960, 16'd35172, 16'd43908, 16'd22242, 16'd56852, 16'd41855, 16'd31604, 16'd53265, 16'd8795, 16'd32220, 16'd35283, 16'd57230, 16'd24998, 16'd63316, 16'd11465, 16'd31082, 16'd30381, 16'd6830, 16'd65113, 16'd24921, 16'd20412, 16'd27295, 16'd47282, 16'd56673, 16'd10025, 16'd63073});
	test_expansion(128'h01ce196447d3fede9871a7092b77c9ef, {16'd45949, 16'd4524, 16'd40364, 16'd5506, 16'd40265, 16'd62952, 16'd63698, 16'd48248, 16'd55885, 16'd28222, 16'd20594, 16'd11958, 16'd15969, 16'd1190, 16'd56823, 16'd10474, 16'd27886, 16'd27598, 16'd47926, 16'd24997, 16'd33254, 16'd49790, 16'd4912, 16'd7184, 16'd44357, 16'd63077});
	test_expansion(128'h2f4deb46f8b7be72ec86f314b581ba77, {16'd38982, 16'd56549, 16'd28503, 16'd62204, 16'd8950, 16'd54041, 16'd43127, 16'd51468, 16'd8159, 16'd57913, 16'd33023, 16'd4688, 16'd20627, 16'd19261, 16'd45492, 16'd5962, 16'd14387, 16'd12934, 16'd32477, 16'd20334, 16'd44274, 16'd15045, 16'd45844, 16'd52931, 16'd48845, 16'd56555});
	test_expansion(128'h42384c7dd419c98a36b32fe236457714, {16'd60614, 16'd63323, 16'd35387, 16'd16624, 16'd36342, 16'd21539, 16'd5917, 16'd40371, 16'd3251, 16'd34841, 16'd21569, 16'd37247, 16'd57031, 16'd17546, 16'd22255, 16'd31321, 16'd34536, 16'd5295, 16'd63930, 16'd60195, 16'd74, 16'd24392, 16'd62014, 16'd63084, 16'd8464, 16'd26101});
	test_expansion(128'he9d29667349c0f04318151b87bc47e59, {16'd3825, 16'd10648, 16'd20740, 16'd23059, 16'd4872, 16'd55377, 16'd39368, 16'd15053, 16'd41718, 16'd6334, 16'd24384, 16'd57252, 16'd29134, 16'd34310, 16'd43320, 16'd41872, 16'd36468, 16'd58776, 16'd39664, 16'd41102, 16'd47775, 16'd29844, 16'd55957, 16'd33242, 16'd61405, 16'd59059});
	test_expansion(128'hadb259bdcdd5ce4146f34b3a5e71169c, {16'd35400, 16'd56056, 16'd61044, 16'd30155, 16'd29924, 16'd22227, 16'd14998, 16'd23628, 16'd9121, 16'd36527, 16'd8959, 16'd32001, 16'd58197, 16'd22574, 16'd33651, 16'd38963, 16'd53529, 16'd34221, 16'd29742, 16'd58904, 16'd47170, 16'd45126, 16'd6771, 16'd3703, 16'd43036, 16'd28170});
	test_expansion(128'h006d75270800e23c43ea791b62f9fa94, {16'd17109, 16'd44393, 16'd30469, 16'd36524, 16'd40309, 16'd47855, 16'd30722, 16'd50244, 16'd23512, 16'd13979, 16'd17739, 16'd54508, 16'd12795, 16'd24849, 16'd59984, 16'd9805, 16'd14335, 16'd61768, 16'd1360, 16'd29350, 16'd48684, 16'd20724, 16'd51280, 16'd51404, 16'd27954, 16'd19305});
	test_expansion(128'h6cbcabd34932387f4eafbe8ec7e606af, {16'd11853, 16'd28555, 16'd26864, 16'd62437, 16'd44655, 16'd8208, 16'd29524, 16'd4981, 16'd5314, 16'd33955, 16'd8383, 16'd48411, 16'd54153, 16'd50691, 16'd29861, 16'd32274, 16'd42749, 16'd13859, 16'd59435, 16'd58787, 16'd34001, 16'd53437, 16'd46134, 16'd62787, 16'd9974, 16'd8370});
	test_expansion(128'hceec8f188b136418db4926c5e33e3d87, {16'd15752, 16'd23537, 16'd18522, 16'd30389, 16'd6856, 16'd23966, 16'd36081, 16'd64306, 16'd64090, 16'd36031, 16'd59975, 16'd63305, 16'd27768, 16'd17836, 16'd58558, 16'd5019, 16'd17866, 16'd4221, 16'd49696, 16'd23811, 16'd25354, 16'd30057, 16'd61807, 16'd7921, 16'd25471, 16'd23744});
	test_expansion(128'hc3b2df93d643a607fa54fbd7f55bb38b, {16'd6646, 16'd61438, 16'd47080, 16'd53248, 16'd49998, 16'd4467, 16'd5733, 16'd1763, 16'd37823, 16'd29353, 16'd12846, 16'd17748, 16'd35859, 16'd16059, 16'd17195, 16'd14992, 16'd65227, 16'd549, 16'd50110, 16'd60519, 16'd56726, 16'd64486, 16'd55777, 16'd13088, 16'd52863, 16'd5120});
	test_expansion(128'hc408af76b3ca13688d68626f9c67feca, {16'd55053, 16'd59579, 16'd9009, 16'd18999, 16'd61797, 16'd20786, 16'd53893, 16'd65083, 16'd23770, 16'd26654, 16'd9601, 16'd50612, 16'd28266, 16'd52364, 16'd34451, 16'd32604, 16'd12548, 16'd44774, 16'd27820, 16'd5338, 16'd57872, 16'd44808, 16'd52818, 16'd40882, 16'd37993, 16'd63836});
	test_expansion(128'h0d9f6a512a51e0b795d9195bf0582f1e, {16'd2101, 16'd12539, 16'd21548, 16'd32910, 16'd42229, 16'd11492, 16'd47083, 16'd27214, 16'd37742, 16'd9656, 16'd3727, 16'd36263, 16'd32056, 16'd14083, 16'd18136, 16'd37151, 16'd22878, 16'd18856, 16'd10671, 16'd14274, 16'd34844, 16'd42468, 16'd2763, 16'd46275, 16'd56701, 16'd30597});
	test_expansion(128'hb6f932b73b983cd6db341f384f25cc2e, {16'd29115, 16'd19565, 16'd34703, 16'd48771, 16'd19121, 16'd20758, 16'd36781, 16'd44416, 16'd48853, 16'd18044, 16'd37640, 16'd51454, 16'd18064, 16'd39894, 16'd29328, 16'd64835, 16'd32799, 16'd47634, 16'd58168, 16'd47823, 16'd23475, 16'd8081, 16'd56141, 16'd45508, 16'd31163, 16'd10788});
	test_expansion(128'h246b78e10568dbc0c8f2fca96f11e135, {16'd15264, 16'd2690, 16'd54186, 16'd41202, 16'd56778, 16'd34410, 16'd55018, 16'd25653, 16'd50207, 16'd22025, 16'd28297, 16'd62205, 16'd6264, 16'd28274, 16'd51495, 16'd55756, 16'd18023, 16'd57600, 16'd38181, 16'd56468, 16'd11350, 16'd16489, 16'd46567, 16'd35191, 16'd13109, 16'd9302});
	test_expansion(128'h79a89b531c0869399b3ff921df5671b1, {16'd1102, 16'd34021, 16'd39043, 16'd44342, 16'd47871, 16'd58465, 16'd628, 16'd20965, 16'd47002, 16'd23464, 16'd239, 16'd10778, 16'd5287, 16'd8952, 16'd56564, 16'd9662, 16'd45822, 16'd56648, 16'd35826, 16'd53785, 16'd59762, 16'd8668, 16'd17400, 16'd44561, 16'd49489, 16'd32364});
	test_expansion(128'ha9f0d3461b67b722eb1be30f61a2bc72, {16'd12806, 16'd22567, 16'd29794, 16'd48130, 16'd57488, 16'd43908, 16'd4936, 16'd54694, 16'd20037, 16'd57207, 16'd5365, 16'd44477, 16'd17880, 16'd57194, 16'd28683, 16'd36740, 16'd59490, 16'd51640, 16'd31142, 16'd63199, 16'd63361, 16'd53002, 16'd35520, 16'd5400, 16'd15168, 16'd61754});
	test_expansion(128'h81d2c58855cda5393345dc99864bb8da, {16'd47458, 16'd50251, 16'd42070, 16'd17856, 16'd5285, 16'd39099, 16'd36249, 16'd61975, 16'd29421, 16'd30908, 16'd60632, 16'd60825, 16'd60670, 16'd29454, 16'd10905, 16'd56953, 16'd35548, 16'd44785, 16'd32709, 16'd20024, 16'd43598, 16'd25039, 16'd63845, 16'd53716, 16'd2405, 16'd29385});
	test_expansion(128'hd7eedff972e030e5474778c8b47571d1, {16'd58983, 16'd28657, 16'd23767, 16'd2500, 16'd23508, 16'd59396, 16'd363, 16'd774, 16'd49072, 16'd21927, 16'd44308, 16'd18159, 16'd41607, 16'd44869, 16'd53928, 16'd57079, 16'd31193, 16'd37503, 16'd29041, 16'd58962, 16'd32508, 16'd5766, 16'd62066, 16'd14714, 16'd57667, 16'd7383});
	test_expansion(128'h7095445dc7f0e7c2dd79a3e7f3e2b52c, {16'd42404, 16'd49823, 16'd42467, 16'd56189, 16'd12668, 16'd11796, 16'd45673, 16'd846, 16'd20990, 16'd55337, 16'd31655, 16'd17260, 16'd63257, 16'd56084, 16'd17303, 16'd26210, 16'd33086, 16'd8222, 16'd15750, 16'd43793, 16'd63183, 16'd17879, 16'd13929, 16'd48403, 16'd10495, 16'd65388});
	test_expansion(128'hefdb9f85ed3962e0ee426626d5c68c30, {16'd40908, 16'd300, 16'd11813, 16'd53600, 16'd12111, 16'd16176, 16'd46787, 16'd23279, 16'd26089, 16'd39806, 16'd21507, 16'd20164, 16'd15149, 16'd33791, 16'd3713, 16'd59680, 16'd10340, 16'd5125, 16'd59698, 16'd31391, 16'd58894, 16'd50786, 16'd27272, 16'd57602, 16'd38910, 16'd53556});
	test_expansion(128'h7617c22c94065897fb23858ea0b529a6, {16'd31424, 16'd55919, 16'd53931, 16'd60073, 16'd56032, 16'd24747, 16'd20593, 16'd38108, 16'd64221, 16'd40560, 16'd61390, 16'd23555, 16'd23148, 16'd23639, 16'd62091, 16'd24482, 16'd39520, 16'd12027, 16'd377, 16'd57145, 16'd1017, 16'd42027, 16'd18917, 16'd41419, 16'd43095, 16'd57912});
	test_expansion(128'h936c0d38ca01e2889a5abcd6057d8045, {16'd18297, 16'd34947, 16'd10114, 16'd18511, 16'd55807, 16'd10864, 16'd7826, 16'd56149, 16'd39627, 16'd30140, 16'd32778, 16'd11349, 16'd14545, 16'd37487, 16'd59563, 16'd54282, 16'd52885, 16'd15752, 16'd55563, 16'd52060, 16'd30927, 16'd29836, 16'd5043, 16'd21320, 16'd35807, 16'd59603});
	test_expansion(128'h547ea1b7b0f2d19cf071d8713a29d2d0, {16'd44042, 16'd11959, 16'd62294, 16'd16019, 16'd47856, 16'd9697, 16'd45537, 16'd37763, 16'd54739, 16'd53214, 16'd5882, 16'd59094, 16'd65292, 16'd40447, 16'd55869, 16'd60787, 16'd51102, 16'd29354, 16'd5015, 16'd3512, 16'd48101, 16'd1082, 16'd24989, 16'd61619, 16'd45966, 16'd31369});
	test_expansion(128'he80f3afbaedf7f0061cfed6fd71a717b, {16'd48424, 16'd59119, 16'd10571, 16'd33671, 16'd13916, 16'd39621, 16'd53824, 16'd51042, 16'd11579, 16'd7016, 16'd39942, 16'd49555, 16'd24662, 16'd34167, 16'd28370, 16'd43825, 16'd53295, 16'd16549, 16'd41979, 16'd64200, 16'd2740, 16'd11090, 16'd38607, 16'd54233, 16'd6939, 16'd39219});
	test_expansion(128'hbdf9acf0d96797accbfb514be4fd1598, {16'd50074, 16'd45845, 16'd58312, 16'd3946, 16'd24701, 16'd53662, 16'd56034, 16'd40288, 16'd6330, 16'd21286, 16'd21723, 16'd42929, 16'd17195, 16'd42949, 16'd65381, 16'd3304, 16'd13658, 16'd31489, 16'd22019, 16'd42501, 16'd57967, 16'd29733, 16'd55974, 16'd1395, 16'd6104, 16'd13516});
	test_expansion(128'ha4f9c1f15c12638742b43a473406e8f6, {16'd27881, 16'd36887, 16'd49201, 16'd630, 16'd14038, 16'd61373, 16'd38632, 16'd22214, 16'd28317, 16'd53607, 16'd45609, 16'd46782, 16'd56288, 16'd58357, 16'd42904, 16'd33142, 16'd28219, 16'd44721, 16'd27521, 16'd62217, 16'd44241, 16'd9164, 16'd60360, 16'd29296, 16'd3821, 16'd22505});
	test_expansion(128'h2cfeb17b4d8d2eed39554d191ec3b5f5, {16'd8222, 16'd44627, 16'd8676, 16'd10410, 16'd37977, 16'd15862, 16'd31870, 16'd24065, 16'd3279, 16'd62180, 16'd52205, 16'd63307, 16'd27912, 16'd19008, 16'd52640, 16'd14877, 16'd42356, 16'd53748, 16'd30297, 16'd2718, 16'd11976, 16'd21852, 16'd59126, 16'd49530, 16'd50714, 16'd47147});
	test_expansion(128'hd88c1e793a18b02d7d1f211212b1ca19, {16'd55042, 16'd10795, 16'd31049, 16'd4578, 16'd37159, 16'd48881, 16'd55188, 16'd28046, 16'd6875, 16'd41060, 16'd21970, 16'd44040, 16'd62086, 16'd37460, 16'd12436, 16'd21430, 16'd15838, 16'd33048, 16'd26066, 16'd10064, 16'd32214, 16'd44353, 16'd7954, 16'd31666, 16'd56824, 16'd41902});
	test_expansion(128'h00e270e49b7f67795ff8650ffc02f628, {16'd46527, 16'd46830, 16'd8487, 16'd38758, 16'd55378, 16'd2308, 16'd6784, 16'd5537, 16'd21568, 16'd1052, 16'd25916, 16'd22618, 16'd38787, 16'd28171, 16'd46668, 16'd45627, 16'd58139, 16'd4464, 16'd9516, 16'd22742, 16'd14083, 16'd37156, 16'd45539, 16'd56968, 16'd58861, 16'd44242});
	test_expansion(128'h361d5d5b2ccc982f8febc9f155ea7148, {16'd47590, 16'd4392, 16'd50415, 16'd18195, 16'd8039, 16'd62640, 16'd36391, 16'd24286, 16'd3652, 16'd55321, 16'd53221, 16'd15961, 16'd24573, 16'd31984, 16'd30852, 16'd47324, 16'd5111, 16'd37183, 16'd23510, 16'd35737, 16'd24571, 16'd18319, 16'd58918, 16'd44411, 16'd2497, 16'd57295});
	test_expansion(128'h2f20ddc8c17e2f167d05b5b25e2a8536, {16'd9053, 16'd26151, 16'd16004, 16'd40778, 16'd7682, 16'd17801, 16'd23420, 16'd25720, 16'd44615, 16'd52209, 16'd27897, 16'd12403, 16'd16117, 16'd41169, 16'd11001, 16'd42650, 16'd46311, 16'd56434, 16'd31680, 16'd17109, 16'd48346, 16'd47248, 16'd36240, 16'd10707, 16'd39055, 16'd42428});
	test_expansion(128'h3c10f0196e4177183cd12ca96bbfd725, {16'd47596, 16'd13158, 16'd21168, 16'd12262, 16'd6373, 16'd35965, 16'd5368, 16'd16861, 16'd58492, 16'd30358, 16'd45457, 16'd17782, 16'd65336, 16'd29823, 16'd23574, 16'd32896, 16'd49592, 16'd28398, 16'd49664, 16'd62955, 16'd55849, 16'd50948, 16'd41557, 16'd25647, 16'd37338, 16'd40086});
	test_expansion(128'h930dcd8770a82124b5243c5f02496757, {16'd337, 16'd58298, 16'd58888, 16'd27565, 16'd13647, 16'd13683, 16'd62168, 16'd150, 16'd38483, 16'd41488, 16'd21918, 16'd47681, 16'd10385, 16'd15809, 16'd38588, 16'd6870, 16'd36349, 16'd27784, 16'd61192, 16'd8396, 16'd41618, 16'd17669, 16'd7859, 16'd31312, 16'd14292, 16'd63972});
	test_expansion(128'h7a8fcf02bca1475b1b1621b40639b613, {16'd20105, 16'd41792, 16'd43634, 16'd10970, 16'd28076, 16'd64218, 16'd37608, 16'd45265, 16'd1921, 16'd19030, 16'd5583, 16'd25546, 16'd61692, 16'd10740, 16'd2500, 16'd54428, 16'd56881, 16'd57155, 16'd13673, 16'd23249, 16'd33004, 16'd42104, 16'd11793, 16'd57262, 16'd30611, 16'd33893});
	test_expansion(128'h35a3438db7bdf6f61f4830a6d22e7169, {16'd41590, 16'd52375, 16'd23881, 16'd49196, 16'd28293, 16'd11836, 16'd54073, 16'd3669, 16'd19311, 16'd4732, 16'd43611, 16'd26462, 16'd46627, 16'd62131, 16'd63925, 16'd22455, 16'd19201, 16'd44732, 16'd22208, 16'd42248, 16'd43885, 16'd63453, 16'd43300, 16'd53494, 16'd65047, 16'd43928});
	test_expansion(128'h7f75b46c34e589001142fef6c96bf475, {16'd7427, 16'd44978, 16'd4178, 16'd4705, 16'd7318, 16'd64601, 16'd33770, 16'd21241, 16'd38198, 16'd11727, 16'd50917, 16'd44661, 16'd52230, 16'd60912, 16'd52869, 16'd49257, 16'd3253, 16'd62501, 16'd9403, 16'd60029, 16'd59206, 16'd25527, 16'd22923, 16'd38252, 16'd15458, 16'd20143});
	test_expansion(128'hefa678c50873669a7e0ff3724fa93124, {16'd280, 16'd30170, 16'd47657, 16'd33163, 16'd46180, 16'd47278, 16'd52768, 16'd51126, 16'd33712, 16'd16279, 16'd36260, 16'd57499, 16'd19569, 16'd20012, 16'd32544, 16'd21243, 16'd63347, 16'd17777, 16'd60788, 16'd27621, 16'd48585, 16'd42768, 16'd32953, 16'd12311, 16'd771, 16'd61278});
	test_expansion(128'hb3072fe3dbdcc474cad73dde7bb24136, {16'd40658, 16'd50402, 16'd5447, 16'd18002, 16'd23823, 16'd18088, 16'd51039, 16'd4369, 16'd53990, 16'd16657, 16'd15789, 16'd24229, 16'd12802, 16'd64518, 16'd61045, 16'd12770, 16'd14286, 16'd58194, 16'd17722, 16'd5658, 16'd43171, 16'd40425, 16'd60859, 16'd2422, 16'd26966, 16'd54951});
	test_expansion(128'h349e3729b5db6254d2a01fae0d5d9a99, {16'd39672, 16'd33424, 16'd5668, 16'd44230, 16'd36449, 16'd36558, 16'd44339, 16'd12524, 16'd6406, 16'd15056, 16'd20007, 16'd8936, 16'd3935, 16'd26992, 16'd21347, 16'd25555, 16'd18431, 16'd32377, 16'd20344, 16'd19679, 16'd36120, 16'd11220, 16'd30825, 16'd6478, 16'd50671, 16'd19420});
	test_expansion(128'h2f0ee5bb4e8143f1a34340766917cede, {16'd40934, 16'd30523, 16'd31159, 16'd30992, 16'd61840, 16'd64717, 16'd27932, 16'd45561, 16'd52188, 16'd48824, 16'd27248, 16'd10554, 16'd33236, 16'd21976, 16'd53979, 16'd55207, 16'd60553, 16'd60786, 16'd33540, 16'd62885, 16'd35936, 16'd30764, 16'd8334, 16'd15350, 16'd28591, 16'd59670});
	test_expansion(128'h8dc051c5bd5139872e8df4cad85f20ae, {16'd15595, 16'd38000, 16'd46713, 16'd49078, 16'd6559, 16'd49654, 16'd42077, 16'd52741, 16'd48312, 16'd3393, 16'd43540, 16'd57492, 16'd35866, 16'd27166, 16'd31695, 16'd23121, 16'd61400, 16'd59783, 16'd48938, 16'd41432, 16'd28771, 16'd26039, 16'd25343, 16'd40874, 16'd32365, 16'd36908});
	test_expansion(128'hed3197f865a0b56562d0a607628b5a52, {16'd52658, 16'd49669, 16'd22690, 16'd20151, 16'd24164, 16'd28445, 16'd65237, 16'd17027, 16'd23017, 16'd5462, 16'd43342, 16'd5921, 16'd13263, 16'd30460, 16'd1301, 16'd5391, 16'd27067, 16'd60190, 16'd56471, 16'd23392, 16'd24725, 16'd11004, 16'd771, 16'd16693, 16'd7786, 16'd609});
	test_expansion(128'h865513329bcb284740d1c18dd0ca305e, {16'd23639, 16'd45463, 16'd63106, 16'd40467, 16'd6251, 16'd33235, 16'd15220, 16'd37859, 16'd8182, 16'd11695, 16'd28847, 16'd9495, 16'd57913, 16'd42947, 16'd23722, 16'd56712, 16'd47513, 16'd48129, 16'd41890, 16'd47044, 16'd10245, 16'd23042, 16'd50853, 16'd28295, 16'd7721, 16'd42153});
	test_expansion(128'hd71e50db286979a51535425ae60b3db7, {16'd1244, 16'd50819, 16'd62106, 16'd60492, 16'd3662, 16'd30620, 16'd58036, 16'd65476, 16'd4247, 16'd20803, 16'd22547, 16'd42227, 16'd12322, 16'd15705, 16'd45375, 16'd63539, 16'd58976, 16'd17724, 16'd21698, 16'd24408, 16'd61304, 16'd19733, 16'd231, 16'd5138, 16'd53630, 16'd5822});
	test_expansion(128'h0ae4dab11b72402f19dca2629f1596ed, {16'd16144, 16'd15240, 16'd10107, 16'd30998, 16'd5537, 16'd26990, 16'd9505, 16'd60718, 16'd49234, 16'd51440, 16'd43848, 16'd53809, 16'd44707, 16'd44094, 16'd5959, 16'd80, 16'd30769, 16'd11465, 16'd1827, 16'd13768, 16'd10805, 16'd26747, 16'd45085, 16'd57397, 16'd11155, 16'd13278});
	test_expansion(128'h370b77a69d782face336c2147b6c6f9b, {16'd14068, 16'd26599, 16'd42886, 16'd16128, 16'd25177, 16'd55465, 16'd3165, 16'd38879, 16'd46747, 16'd19164, 16'd4253, 16'd57907, 16'd49407, 16'd46397, 16'd20735, 16'd40948, 16'd7447, 16'd52973, 16'd50540, 16'd11623, 16'd33769, 16'd56728, 16'd21139, 16'd25291, 16'd9062, 16'd36713});
	test_expansion(128'h77c7f6d479b07d3f39176376eb191892, {16'd4488, 16'd18070, 16'd10553, 16'd19174, 16'd54130, 16'd55929, 16'd31343, 16'd6091, 16'd43430, 16'd13386, 16'd39867, 16'd54067, 16'd55711, 16'd38974, 16'd57705, 16'd26005, 16'd40724, 16'd65396, 16'd15083, 16'd32496, 16'd65307, 16'd19726, 16'd34471, 16'd37878, 16'd1543, 16'd13796});
	test_expansion(128'h6a31cb616f5af55a2471287ed0f691f6, {16'd12519, 16'd6351, 16'd12467, 16'd29738, 16'd43000, 16'd1781, 16'd39451, 16'd3922, 16'd59047, 16'd1505, 16'd30697, 16'd62385, 16'd9857, 16'd63969, 16'd11761, 16'd15917, 16'd14836, 16'd9995, 16'd26383, 16'd33058, 16'd16200, 16'd34877, 16'd19497, 16'd21331, 16'd35645, 16'd16147});
	test_expansion(128'hbca02250df761005b23f3b7e08729205, {16'd15622, 16'd55185, 16'd63017, 16'd16874, 16'd12941, 16'd47671, 16'd14224, 16'd56096, 16'd40967, 16'd26411, 16'd59023, 16'd52291, 16'd39972, 16'd59951, 16'd48224, 16'd56802, 16'd24216, 16'd36251, 16'd27067, 16'd28903, 16'd17637, 16'd52793, 16'd63492, 16'd22614, 16'd51638, 16'd52755});
	test_expansion(128'h253fb2031aa5e7ae96aecf6774246e76, {16'd39121, 16'd33607, 16'd3959, 16'd53477, 16'd43781, 16'd1427, 16'd23727, 16'd62625, 16'd17361, 16'd18622, 16'd48665, 16'd29180, 16'd17658, 16'd3506, 16'd60506, 16'd4722, 16'd28678, 16'd33738, 16'd54099, 16'd22478, 16'd2921, 16'd21474, 16'd7725, 16'd44587, 16'd64033, 16'd48601});
	test_expansion(128'hf8fe06627c11d9adf644eb92d341b3f7, {16'd49699, 16'd12356, 16'd61556, 16'd23731, 16'd28238, 16'd46774, 16'd39678, 16'd6870, 16'd24952, 16'd56321, 16'd61589, 16'd27289, 16'd54603, 16'd17805, 16'd10262, 16'd14840, 16'd3924, 16'd18318, 16'd10771, 16'd27035, 16'd14762, 16'd13361, 16'd27496, 16'd55873, 16'd40242, 16'd57208});
	test_expansion(128'ha4e91385909c774c62d6076e219cf746, {16'd1247, 16'd65351, 16'd31167, 16'd40579, 16'd23264, 16'd14719, 16'd48921, 16'd24465, 16'd55020, 16'd9241, 16'd62739, 16'd64160, 16'd35626, 16'd59395, 16'd10608, 16'd29212, 16'd2980, 16'd20620, 16'd48256, 16'd9563, 16'd39932, 16'd300, 16'd30663, 16'd15557, 16'd49282, 16'd9683});
	test_expansion(128'hadca113c7a5f7cb5c66787ac16fd7d23, {16'd44390, 16'd35739, 16'd16711, 16'd33416, 16'd35300, 16'd38193, 16'd30028, 16'd41124, 16'd34844, 16'd64343, 16'd29687, 16'd6515, 16'd3875, 16'd64199, 16'd7773, 16'd58019, 16'd37732, 16'd59642, 16'd8109, 16'd53464, 16'd10084, 16'd25636, 16'd46183, 16'd13893, 16'd45671, 16'd51650});
	test_expansion(128'hbebf072dfd329554a7bc071acb99fa67, {16'd36360, 16'd59065, 16'd32214, 16'd61138, 16'd30659, 16'd11502, 16'd64726, 16'd38338, 16'd21863, 16'd64725, 16'd5060, 16'd4562, 16'd63031, 16'd60951, 16'd20821, 16'd51338, 16'd1762, 16'd63561, 16'd16855, 16'd10347, 16'd13345, 16'd57769, 16'd46781, 16'd25112, 16'd41682, 16'd21300});
	test_expansion(128'h9ecf4a628ecbfa40b84d64b431d3f215, {16'd34054, 16'd62843, 16'd18339, 16'd50223, 16'd2705, 16'd58907, 16'd43166, 16'd28727, 16'd15371, 16'd24296, 16'd7502, 16'd10135, 16'd51989, 16'd379, 16'd42804, 16'd22554, 16'd49851, 16'd15078, 16'd544, 16'd64800, 16'd53643, 16'd54148, 16'd26704, 16'd36011, 16'd45440, 16'd52256});
	test_expansion(128'hd475459aca3eee85955000c683c48fed, {16'd4773, 16'd24979, 16'd8274, 16'd2530, 16'd64114, 16'd58085, 16'd20747, 16'd7355, 16'd12751, 16'd674, 16'd33480, 16'd8689, 16'd43919, 16'd6798, 16'd8513, 16'd25722, 16'd63282, 16'd59118, 16'd15736, 16'd3924, 16'd48232, 16'd61163, 16'd44532, 16'd48089, 16'd18379, 16'd2175});
	test_expansion(128'h762ba122e5defe1d9554d6b6fc38a931, {16'd16898, 16'd27016, 16'd15517, 16'd1433, 16'd53640, 16'd53058, 16'd42692, 16'd41079, 16'd62292, 16'd63766, 16'd17505, 16'd15736, 16'd32045, 16'd11625, 16'd17294, 16'd25517, 16'd10748, 16'd5402, 16'd61372, 16'd1918, 16'd41216, 16'd8263, 16'd20932, 16'd4575, 16'd16668, 16'd47041});
	test_expansion(128'hd11f2b4f7732910742b95055576cba58, {16'd40700, 16'd17013, 16'd13569, 16'd65065, 16'd4031, 16'd39380, 16'd64407, 16'd63160, 16'd16268, 16'd60065, 16'd46994, 16'd40871, 16'd59609, 16'd4895, 16'd65386, 16'd3293, 16'd1261, 16'd41813, 16'd8952, 16'd57007, 16'd37063, 16'd52107, 16'd2220, 16'd52895, 16'd33507, 16'd9534});
	test_expansion(128'h41b015b63e7320d58ba52b18ee4a5ad1, {16'd58504, 16'd25379, 16'd10518, 16'd9753, 16'd57234, 16'd58535, 16'd16500, 16'd9095, 16'd1254, 16'd24599, 16'd55118, 16'd40608, 16'd38939, 16'd57411, 16'd25452, 16'd780, 16'd16735, 16'd22075, 16'd17916, 16'd44197, 16'd11213, 16'd25084, 16'd22664, 16'd3997, 16'd44076, 16'd58774});
	test_expansion(128'h7ab6f28b42946283542f07c03a48063d, {16'd517, 16'd28586, 16'd59476, 16'd63806, 16'd51586, 16'd2871, 16'd25072, 16'd8432, 16'd35181, 16'd46893, 16'd47695, 16'd53059, 16'd26439, 16'd50499, 16'd18254, 16'd32233, 16'd12327, 16'd46906, 16'd50476, 16'd3562, 16'd39640, 16'd51802, 16'd5216, 16'd28296, 16'd53441, 16'd34268});
	test_expansion(128'he0ecffe4cbf4a6fa5ae6ffab05b834cd, {16'd30652, 16'd27066, 16'd53037, 16'd57999, 16'd49358, 16'd10813, 16'd4039, 16'd18031, 16'd58566, 16'd11457, 16'd62331, 16'd7830, 16'd58080, 16'd40200, 16'd15297, 16'd42094, 16'd38236, 16'd22630, 16'd12288, 16'd33567, 16'd11193, 16'd56882, 16'd43822, 16'd36418, 16'd58611, 16'd26879});
	test_expansion(128'h9efe986f07a5c996aa77de8e8d88db29, {16'd57990, 16'd59436, 16'd57392, 16'd62330, 16'd49218, 16'd21762, 16'd8824, 16'd12840, 16'd27565, 16'd28428, 16'd48512, 16'd19177, 16'd14880, 16'd37362, 16'd30175, 16'd45463, 16'd49414, 16'd30361, 16'd32614, 16'd54062, 16'd11425, 16'd15127, 16'd25830, 16'd27737, 16'd42884, 16'd35439});
	test_expansion(128'h09f45bee1927dc1a26878f65cd91f92f, {16'd4003, 16'd44403, 16'd52184, 16'd35019, 16'd55214, 16'd55314, 16'd5673, 16'd40703, 16'd57510, 16'd41936, 16'd35680, 16'd2913, 16'd15514, 16'd28480, 16'd48104, 16'd55561, 16'd17985, 16'd23918, 16'd4117, 16'd59726, 16'd19866, 16'd26976, 16'd42235, 16'd63224, 16'd44274, 16'd57157});
	test_expansion(128'h02462e3f611caac335dfcdbef859120c, {16'd17707, 16'd12947, 16'd37488, 16'd35535, 16'd56635, 16'd2664, 16'd13775, 16'd57283, 16'd27720, 16'd62116, 16'd16287, 16'd31963, 16'd63618, 16'd55707, 16'd40722, 16'd1524, 16'd10110, 16'd13356, 16'd49084, 16'd60559, 16'd48332, 16'd32903, 16'd62216, 16'd49368, 16'd60811, 16'd12714});
	test_expansion(128'h4df835f52a31fab00b7197100cfc04aa, {16'd49881, 16'd53249, 16'd20953, 16'd19096, 16'd44257, 16'd47442, 16'd30156, 16'd14173, 16'd2042, 16'd64475, 16'd7737, 16'd52475, 16'd25267, 16'd65269, 16'd20780, 16'd49650, 16'd60166, 16'd41591, 16'd64785, 16'd9221, 16'd39411, 16'd41941, 16'd44182, 16'd24667, 16'd40005, 16'd42499});
	test_expansion(128'h2473593c0fe11db2a4f9233b16ab9a46, {16'd62106, 16'd46547, 16'd10083, 16'd10381, 16'd28855, 16'd38869, 16'd46092, 16'd65384, 16'd57590, 16'd61763, 16'd40397, 16'd14261, 16'd60372, 16'd55270, 16'd22032, 16'd26149, 16'd42704, 16'd14895, 16'd60347, 16'd11702, 16'd24961, 16'd15326, 16'd9007, 16'd43674, 16'd59660, 16'd32453});
	test_expansion(128'h4d243a3638b76f36d10fed2f73ac2932, {16'd56248, 16'd45848, 16'd52872, 16'd43940, 16'd58652, 16'd29195, 16'd33473, 16'd16775, 16'd38095, 16'd11837, 16'd59720, 16'd20693, 16'd65134, 16'd46205, 16'd49596, 16'd40763, 16'd39508, 16'd59689, 16'd11396, 16'd12927, 16'd35625, 16'd5534, 16'd61005, 16'd61986, 16'd52265, 16'd32978});
	test_expansion(128'h8d43a8f86ae47924d18399f835e3680d, {16'd5517, 16'd23948, 16'd43516, 16'd9648, 16'd44252, 16'd31132, 16'd58641, 16'd45615, 16'd57070, 16'd17985, 16'd4925, 16'd39610, 16'd26442, 16'd29975, 16'd52666, 16'd26894, 16'd38456, 16'd36658, 16'd38357, 16'd61207, 16'd28168, 16'd54912, 16'd21443, 16'd60653, 16'd22588, 16'd19149});
	test_expansion(128'h3c9dd94b61a323c1ffa4e737409c57df, {16'd17481, 16'd15211, 16'd9022, 16'd25532, 16'd7104, 16'd63454, 16'd55486, 16'd16969, 16'd12530, 16'd58536, 16'd61270, 16'd27746, 16'd43018, 16'd51617, 16'd26522, 16'd29927, 16'd8969, 16'd21907, 16'd62802, 16'd6291, 16'd61374, 16'd41442, 16'd17828, 16'd11578, 16'd54633, 16'd20894});
	test_expansion(128'hef99dbc494fb0b9f1e4808f1caaa293e, {16'd44518, 16'd44439, 16'd30458, 16'd27206, 16'd48640, 16'd45352, 16'd52225, 16'd25239, 16'd43980, 16'd39150, 16'd3861, 16'd21409, 16'd8790, 16'd28771, 16'd13157, 16'd505, 16'd29545, 16'd7362, 16'd60493, 16'd2390, 16'd53233, 16'd47338, 16'd13004, 16'd59222, 16'd458, 16'd4708});
	test_expansion(128'hc92260a982568fbd0fe938bddd8d69ca, {16'd43341, 16'd43133, 16'd29391, 16'd46994, 16'd9574, 16'd6448, 16'd41073, 16'd45231, 16'd18882, 16'd18000, 16'd5467, 16'd44899, 16'd37251, 16'd23313, 16'd64394, 16'd3052, 16'd63015, 16'd58472, 16'd64149, 16'd30152, 16'd48050, 16'd55552, 16'd41238, 16'd34757, 16'd43508, 16'd56996});
	test_expansion(128'h1e75b8fcdf90cbee5c100b0a551fc5fd, {16'd11169, 16'd22458, 16'd32556, 16'd16225, 16'd23670, 16'd10033, 16'd17828, 16'd65081, 16'd42231, 16'd12253, 16'd5005, 16'd34874, 16'd42501, 16'd29121, 16'd18492, 16'd954, 16'd7142, 16'd17422, 16'd41413, 16'd12008, 16'd34802, 16'd28012, 16'd62268, 16'd27733, 16'd55958, 16'd15887});
	test_expansion(128'hb5db847bc319643997d5f4277f732d23, {16'd24524, 16'd65499, 16'd64930, 16'd8552, 16'd16849, 16'd47735, 16'd13860, 16'd36460, 16'd32267, 16'd61487, 16'd28108, 16'd49661, 16'd28080, 16'd45683, 16'd7330, 16'd51797, 16'd12245, 16'd5525, 16'd51957, 16'd34156, 16'd25418, 16'd14032, 16'd45583, 16'd23202, 16'd33982, 16'd33955});
	test_expansion(128'h6aa51dd3fcd5af8b85a939cc7a735ae0, {16'd51930, 16'd64190, 16'd36518, 16'd30352, 16'd13108, 16'd16311, 16'd60587, 16'd60188, 16'd919, 16'd24388, 16'd42069, 16'd15713, 16'd35470, 16'd33822, 16'd21047, 16'd60263, 16'd20468, 16'd46867, 16'd206, 16'd29219, 16'd63306, 16'd36477, 16'd19924, 16'd35738, 16'd32598, 16'd3391});
	test_expansion(128'hcb08a03d0f3245e2a6db1cf52af2d699, {16'd49445, 16'd60056, 16'd61652, 16'd22016, 16'd62464, 16'd64327, 16'd65522, 16'd28885, 16'd4172, 16'd54740, 16'd24711, 16'd5016, 16'd22212, 16'd26054, 16'd57118, 16'd18962, 16'd6348, 16'd29405, 16'd33853, 16'd40730, 16'd55241, 16'd48481, 16'd30382, 16'd6141, 16'd40713, 16'd26238});
	test_expansion(128'hd91980e9e131f8c78d650ec0f9b0689d, {16'd20872, 16'd39860, 16'd51531, 16'd31214, 16'd49834, 16'd1838, 16'd38095, 16'd45463, 16'd31508, 16'd35047, 16'd37554, 16'd29058, 16'd54128, 16'd43551, 16'd14989, 16'd60357, 16'd12490, 16'd29836, 16'd11044, 16'd15551, 16'd57165, 16'd8123, 16'd64094, 16'd12098, 16'd55764, 16'd12341});
	test_expansion(128'hc014aab8b9748da3d8409d33435c26d7, {16'd4755, 16'd61014, 16'd11314, 16'd57522, 16'd20386, 16'd29414, 16'd41110, 16'd23414, 16'd7914, 16'd27133, 16'd51239, 16'd27493, 16'd1108, 16'd21128, 16'd576, 16'd21989, 16'd3424, 16'd6006, 16'd12235, 16'd37859, 16'd12363, 16'd8026, 16'd47183, 16'd53698, 16'd49971, 16'd5956});
	test_expansion(128'h349ae0b3976f32e7641e43c971b924f3, {16'd8887, 16'd15487, 16'd55652, 16'd12465, 16'd45548, 16'd24145, 16'd23631, 16'd60881, 16'd45789, 16'd9907, 16'd32135, 16'd23736, 16'd50875, 16'd41058, 16'd15675, 16'd36646, 16'd42056, 16'd7167, 16'd13726, 16'd44133, 16'd38933, 16'd11981, 16'd4835, 16'd26826, 16'd58281, 16'd21445});
	test_expansion(128'h7ef91514a288644bbaa5cadaf8657e02, {16'd1048, 16'd7366, 16'd8049, 16'd50341, 16'd1002, 16'd49556, 16'd49218, 16'd40949, 16'd34150, 16'd26430, 16'd37049, 16'd39962, 16'd25460, 16'd4084, 16'd39423, 16'd59633, 16'd12103, 16'd5960, 16'd28231, 16'd1707, 16'd12765, 16'd57164, 16'd32008, 16'd52879, 16'd5815, 16'd38480});
	test_expansion(128'h49bc65c1397d8a24969a3bc9624423ee, {16'd36453, 16'd28720, 16'd41157, 16'd59137, 16'd34731, 16'd23418, 16'd4444, 16'd8885, 16'd19523, 16'd56413, 16'd38543, 16'd26264, 16'd58658, 16'd36582, 16'd53266, 16'd31132, 16'd58826, 16'd62778, 16'd53081, 16'd5954, 16'd9087, 16'd22798, 16'd41885, 16'd17398, 16'd51339, 16'd51072});
	test_expansion(128'h3b1a96fef746d5dd9510dfef899766bb, {16'd6231, 16'd1719, 16'd20658, 16'd30361, 16'd35345, 16'd21367, 16'd19581, 16'd64891, 16'd51335, 16'd54254, 16'd54182, 16'd46630, 16'd27674, 16'd13185, 16'd3478, 16'd54132, 16'd20071, 16'd15348, 16'd62542, 16'd50789, 16'd2986, 16'd36477, 16'd4611, 16'd36581, 16'd39431, 16'd26199});
	test_expansion(128'h70341fc1116431fafea72fbbc6f0f46b, {16'd39005, 16'd62248, 16'd43481, 16'd60252, 16'd36506, 16'd46445, 16'd20672, 16'd25248, 16'd63992, 16'd26446, 16'd2985, 16'd32955, 16'd722, 16'd10925, 16'd42297, 16'd51856, 16'd12968, 16'd27916, 16'd23033, 16'd2885, 16'd63617, 16'd7508, 16'd10881, 16'd47443, 16'd20319, 16'd61313});
	test_expansion(128'h5d1e6e3021a0be0e2d370d679563367c, {16'd9987, 16'd62889, 16'd14997, 16'd55120, 16'd8258, 16'd33673, 16'd16860, 16'd26329, 16'd8711, 16'd10161, 16'd58926, 16'd52141, 16'd30587, 16'd16993, 16'd43418, 16'd43940, 16'd36222, 16'd22251, 16'd43194, 16'd55441, 16'd32966, 16'd11986, 16'd10231, 16'd18443, 16'd52091, 16'd43791});
	test_expansion(128'hf16d1503f91cae3e0168e536f9b97b62, {16'd63620, 16'd28628, 16'd31317, 16'd15062, 16'd2691, 16'd10834, 16'd52911, 16'd15626, 16'd9128, 16'd31220, 16'd13049, 16'd187, 16'd65156, 16'd47227, 16'd1597, 16'd21248, 16'd36173, 16'd40587, 16'd36087, 16'd26258, 16'd53057, 16'd58703, 16'd42423, 16'd4877, 16'd3971, 16'd59868});
	test_expansion(128'h0be80b4d8c744bc8261186b3dc66c116, {16'd33291, 16'd57729, 16'd39913, 16'd28490, 16'd61981, 16'd22923, 16'd55930, 16'd35862, 16'd49851, 16'd22058, 16'd51545, 16'd22158, 16'd37957, 16'd1707, 16'd35565, 16'd21761, 16'd4771, 16'd5590, 16'd60440, 16'd28567, 16'd373, 16'd17879, 16'd63915, 16'd33047, 16'd48581, 16'd29541});
	test_expansion(128'h2446ad885e542857edae190189312d36, {16'd11413, 16'd958, 16'd7572, 16'd8697, 16'd2316, 16'd3971, 16'd24489, 16'd48343, 16'd45910, 16'd54209, 16'd51667, 16'd36055, 16'd47403, 16'd18131, 16'd13923, 16'd797, 16'd20966, 16'd22697, 16'd54107, 16'd26854, 16'd50324, 16'd42201, 16'd35955, 16'd13853, 16'd13980, 16'd19825});
	test_expansion(128'h2e429fafa777da7bf1b8db617021047b, {16'd685, 16'd42328, 16'd30225, 16'd18750, 16'd36255, 16'd22763, 16'd43116, 16'd61132, 16'd54529, 16'd28571, 16'd30423, 16'd39422, 16'd18732, 16'd45401, 16'd5138, 16'd14282, 16'd43650, 16'd60503, 16'd25521, 16'd55777, 16'd27277, 16'd51761, 16'd32956, 16'd22655, 16'd39506, 16'd52593});
	test_expansion(128'h12d8ef7f2ec15e277d7d6f733dc1ccf5, {16'd61928, 16'd48849, 16'd59587, 16'd65516, 16'd38608, 16'd26757, 16'd26938, 16'd21271, 16'd56040, 16'd33366, 16'd53504, 16'd7941, 16'd17541, 16'd46753, 16'd3358, 16'd59386, 16'd58178, 16'd12786, 16'd40024, 16'd41283, 16'd38293, 16'd43098, 16'd44580, 16'd5886, 16'd62913, 16'd15272});
	test_expansion(128'h07d738261518b65397bf9c478d864db9, {16'd40987, 16'd37955, 16'd18550, 16'd26067, 16'd58971, 16'd37959, 16'd6251, 16'd51344, 16'd63257, 16'd29360, 16'd63659, 16'd51894, 16'd3136, 16'd8427, 16'd55238, 16'd22441, 16'd19718, 16'd14028, 16'd59928, 16'd48538, 16'd61586, 16'd49285, 16'd37904, 16'd5271, 16'd56050, 16'd53843});
	test_expansion(128'h4c237525a1fe472bbf334077a6db9f77, {16'd27253, 16'd65378, 16'd8852, 16'd15049, 16'd62848, 16'd57729, 16'd3968, 16'd49849, 16'd62312, 16'd46444, 16'd26566, 16'd4189, 16'd24475, 16'd62770, 16'd54823, 16'd60704, 16'd839, 16'd2044, 16'd58271, 16'd53656, 16'd31463, 16'd25320, 16'd16223, 16'd17945, 16'd2711, 16'd19892});
	test_expansion(128'hb08a9906de70bc305ac3f70c48b66ed6, {16'd17683, 16'd9673, 16'd8739, 16'd30617, 16'd3021, 16'd18626, 16'd39386, 16'd47730, 16'd27528, 16'd39909, 16'd27170, 16'd39254, 16'd8561, 16'd26863, 16'd62387, 16'd23923, 16'd57641, 16'd19595, 16'd35294, 16'd23762, 16'd62489, 16'd51076, 16'd49346, 16'd36932, 16'd33179, 16'd27263});
	test_expansion(128'h34337f7fcf8bfa84961f5b4c8764f603, {16'd61678, 16'd56310, 16'd4263, 16'd29780, 16'd16763, 16'd28584, 16'd15100, 16'd52674, 16'd58319, 16'd45652, 16'd13355, 16'd34942, 16'd65296, 16'd39232, 16'd41374, 16'd11551, 16'd63275, 16'd22854, 16'd52092, 16'd4233, 16'd1879, 16'd46460, 16'd58166, 16'd31848, 16'd17556, 16'd5991});
	test_expansion(128'h4ab66611704625acbd0fecdd0edffa02, {16'd30423, 16'd58021, 16'd21088, 16'd33775, 16'd29125, 16'd24417, 16'd54491, 16'd46925, 16'd18493, 16'd29046, 16'd48312, 16'd22372, 16'd3938, 16'd54666, 16'd60910, 16'd63526, 16'd33217, 16'd45389, 16'd7223, 16'd19978, 16'd50475, 16'd30751, 16'd43267, 16'd37007, 16'd33291, 16'd40170});
	test_expansion(128'h8e377e9bf0c920042e259f8465c21464, {16'd59031, 16'd43093, 16'd21340, 16'd3182, 16'd33365, 16'd42327, 16'd22029, 16'd24108, 16'd53985, 16'd61907, 16'd49152, 16'd48770, 16'd64314, 16'd22924, 16'd19888, 16'd33869, 16'd32034, 16'd50518, 16'd8150, 16'd32094, 16'd44017, 16'd62075, 16'd24470, 16'd48489, 16'd45487, 16'd37249});
	test_expansion(128'h147318e95aa61b0d4bcc7164956ba80c, {16'd10467, 16'd10486, 16'd8997, 16'd60378, 16'd3057, 16'd21519, 16'd38457, 16'd32732, 16'd61663, 16'd9924, 16'd4354, 16'd49598, 16'd41534, 16'd58140, 16'd51099, 16'd44001, 16'd2330, 16'd1080, 16'd11496, 16'd24846, 16'd36765, 16'd63433, 16'd26556, 16'd30576, 16'd643, 16'd62955});
	test_expansion(128'h21aebcf99994407a68276d6b8e5b94e8, {16'd38746, 16'd64204, 16'd10194, 16'd16138, 16'd54607, 16'd55660, 16'd52376, 16'd6538, 16'd22669, 16'd12572, 16'd34482, 16'd59299, 16'd64598, 16'd30216, 16'd40050, 16'd25257, 16'd48228, 16'd47148, 16'd63498, 16'd19491, 16'd44231, 16'd42088, 16'd61062, 16'd42568, 16'd18207, 16'd61882});
	test_expansion(128'h8632be83c76af365ee311e00609a9a60, {16'd16221, 16'd30970, 16'd22501, 16'd34025, 16'd30609, 16'd36721, 16'd2523, 16'd46015, 16'd44335, 16'd10319, 16'd39719, 16'd22980, 16'd2670, 16'd46826, 16'd32589, 16'd20840, 16'd43355, 16'd49348, 16'd64989, 16'd20783, 16'd54208, 16'd893, 16'd48317, 16'd5669, 16'd50994, 16'd45489});
	test_expansion(128'h9b97ba13f0dea8c68e8b1846d9409a5b, {16'd51811, 16'd4682, 16'd51911, 16'd61581, 16'd27851, 16'd17499, 16'd59671, 16'd15480, 16'd54395, 16'd1957, 16'd43349, 16'd17464, 16'd8175, 16'd37074, 16'd11729, 16'd51031, 16'd8900, 16'd15152, 16'd32332, 16'd49288, 16'd13783, 16'd43110, 16'd58695, 16'd30915, 16'd58000, 16'd21125});
	test_expansion(128'hb5e011b8906fce6f3a6f699629016ff6, {16'd58225, 16'd296, 16'd45439, 16'd12003, 16'd29866, 16'd53762, 16'd18734, 16'd64098, 16'd16613, 16'd11511, 16'd63309, 16'd63266, 16'd34356, 16'd43651, 16'd26629, 16'd7394, 16'd31461, 16'd16355, 16'd28187, 16'd12042, 16'd64637, 16'd7548, 16'd30125, 16'd6837, 16'd35580, 16'd63533});
	test_expansion(128'h55b454b4be4f53a2d02d91b3308e3794, {16'd21104, 16'd20534, 16'd7320, 16'd41071, 16'd14278, 16'd29618, 16'd52459, 16'd53600, 16'd48983, 16'd37190, 16'd34657, 16'd62384, 16'd65533, 16'd56581, 16'd13972, 16'd61098, 16'd15425, 16'd61161, 16'd22113, 16'd35235, 16'd5117, 16'd38986, 16'd14435, 16'd28030, 16'd47984, 16'd15450});
	test_expansion(128'h632dcb8206160fc10dd6a07e6335b9e1, {16'd63533, 16'd55883, 16'd24700, 16'd64626, 16'd26102, 16'd31909, 16'd26366, 16'd58196, 16'd29713, 16'd9663, 16'd46130, 16'd53456, 16'd26928, 16'd24790, 16'd12169, 16'd55366, 16'd58769, 16'd13549, 16'd4690, 16'd12913, 16'd30243, 16'd25361, 16'd33922, 16'd41253, 16'd42023, 16'd2872});
	test_expansion(128'hc0633b329e8e2662448155f771b867f2, {16'd29589, 16'd20742, 16'd15641, 16'd53960, 16'd1542, 16'd57409, 16'd63397, 16'd43766, 16'd61364, 16'd8875, 16'd24995, 16'd39281, 16'd5636, 16'd25132, 16'd615, 16'd4029, 16'd43228, 16'd45163, 16'd42922, 16'd44092, 16'd1911, 16'd18752, 16'd35121, 16'd20521, 16'd41333, 16'd14161});
	test_expansion(128'h754b5e9d0ffcc55b592c3f6535406396, {16'd42627, 16'd29160, 16'd28289, 16'd36580, 16'd19800, 16'd14361, 16'd35887, 16'd53530, 16'd9172, 16'd44637, 16'd1001, 16'd50533, 16'd32177, 16'd58470, 16'd15197, 16'd1782, 16'd20698, 16'd30532, 16'd61543, 16'd54444, 16'd60213, 16'd17017, 16'd49262, 16'd62954, 16'd14223, 16'd57410});
	test_expansion(128'hd7c23355d59a0f7735a79551ec818f1a, {16'd61420, 16'd10194, 16'd50121, 16'd43079, 16'd19289, 16'd8692, 16'd6623, 16'd11719, 16'd1498, 16'd45496, 16'd2384, 16'd30569, 16'd12017, 16'd461, 16'd10250, 16'd57071, 16'd27919, 16'd30418, 16'd62658, 16'd2019, 16'd1470, 16'd7941, 16'd49114, 16'd21059, 16'd62825, 16'd14536});
	test_expansion(128'h84f9cc35f49da029920bf7e6900d01e4, {16'd12583, 16'd44887, 16'd41974, 16'd8165, 16'd65174, 16'd54471, 16'd49722, 16'd25806, 16'd53660, 16'd11131, 16'd1057, 16'd44100, 16'd1196, 16'd39451, 16'd23551, 16'd20156, 16'd32631, 16'd46314, 16'd23801, 16'd14415, 16'd27016, 16'd24481, 16'd63214, 16'd36911, 16'd1964, 16'd25369});
	test_expansion(128'h028c15b0fc2325233285769ca4169f5f, {16'd54133, 16'd34304, 16'd34586, 16'd28166, 16'd24515, 16'd33980, 16'd19591, 16'd16396, 16'd59606, 16'd21015, 16'd3842, 16'd13043, 16'd61095, 16'd27770, 16'd12506, 16'd28953, 16'd18078, 16'd61020, 16'd31518, 16'd3477, 16'd37530, 16'd5200, 16'd63910, 16'd26357, 16'd20249, 16'd10874});
	test_expansion(128'hc60223c7e9e4c451bb306c4085be2063, {16'd1719, 16'd63285, 16'd60499, 16'd33852, 16'd41772, 16'd27094, 16'd53206, 16'd39259, 16'd42992, 16'd13053, 16'd3140, 16'd49245, 16'd31353, 16'd2583, 16'd18934, 16'd39139, 16'd535, 16'd12070, 16'd15916, 16'd1644, 16'd56657, 16'd24177, 16'd19425, 16'd31249, 16'd58042, 16'd31839});
	test_expansion(128'hce931a2f753f11fface5626025d0d36f, {16'd20981, 16'd17751, 16'd21827, 16'd46487, 16'd43345, 16'd31285, 16'd44442, 16'd29653, 16'd15875, 16'd1754, 16'd22254, 16'd53062, 16'd18711, 16'd30952, 16'd25350, 16'd50949, 16'd32482, 16'd19627, 16'd19026, 16'd24939, 16'd29631, 16'd47247, 16'd30268, 16'd22471, 16'd43730, 16'd7943});
	test_expansion(128'haf6a57361102f3215c8e484724f1fa77, {16'd44339, 16'd36537, 16'd50609, 16'd27616, 16'd47210, 16'd51333, 16'd16541, 16'd7746, 16'd63670, 16'd54390, 16'd30482, 16'd63290, 16'd59987, 16'd24585, 16'd54755, 16'd38053, 16'd19421, 16'd6250, 16'd17670, 16'd4690, 16'd34376, 16'd36211, 16'd62449, 16'd19640, 16'd37670, 16'd6718});
	test_expansion(128'h170566f0a576f15f4091fd41684753a4, {16'd18121, 16'd36831, 16'd37371, 16'd5453, 16'd9400, 16'd54862, 16'd28604, 16'd6839, 16'd35634, 16'd56094, 16'd25523, 16'd19812, 16'd27507, 16'd25321, 16'd8711, 16'd5994, 16'd16141, 16'd18263, 16'd42875, 16'd5212, 16'd32546, 16'd43810, 16'd15420, 16'd29388, 16'd63517, 16'd13083});
	test_expansion(128'ha4840b1fe60b43ee2a96cbd85b248015, {16'd11639, 16'd15567, 16'd15368, 16'd51426, 16'd9561, 16'd24116, 16'd16012, 16'd16636, 16'd29916, 16'd57197, 16'd43757, 16'd13757, 16'd21003, 16'd47432, 16'd35598, 16'd65279, 16'd44112, 16'd53680, 16'd16316, 16'd5430, 16'd53397, 16'd42221, 16'd28011, 16'd25311, 16'd16948, 16'd45174});
	test_expansion(128'h45aff0b7cde5db4f72b022ad6a5d6975, {16'd1415, 16'd45921, 16'd37736, 16'd64948, 16'd14938, 16'd14138, 16'd48878, 16'd17910, 16'd50513, 16'd1953, 16'd9460, 16'd27652, 16'd33009, 16'd16100, 16'd52584, 16'd38888, 16'd61691, 16'd55369, 16'd1870, 16'd3866, 16'd13043, 16'd33870, 16'd50889, 16'd26625, 16'd61230, 16'd18600});
	test_expansion(128'h0d30d5c7c95fe24eea37bf4b3a6bc1a6, {16'd50707, 16'd45883, 16'd12981, 16'd36311, 16'd40244, 16'd29772, 16'd64445, 16'd46800, 16'd2368, 16'd9368, 16'd39904, 16'd9095, 16'd45664, 16'd4848, 16'd47813, 16'd30973, 16'd874, 16'd30138, 16'd24582, 16'd32012, 16'd20405, 16'd40037, 16'd18292, 16'd42114, 16'd18763, 16'd52271});
	test_expansion(128'h89a5eb79bb79afc4c8fefef0fb507267, {16'd51892, 16'd8860, 16'd474, 16'd14164, 16'd62371, 16'd62627, 16'd14181, 16'd52397, 16'd60720, 16'd20285, 16'd60490, 16'd27539, 16'd54998, 16'd40410, 16'd50674, 16'd31647, 16'd53555, 16'd17600, 16'd52733, 16'd51585, 16'd37475, 16'd50983, 16'd65262, 16'd28167, 16'd23814, 16'd6009});
	test_expansion(128'h84eb73858c5ae874e8896d05880e2647, {16'd51064, 16'd58233, 16'd3696, 16'd15686, 16'd560, 16'd57085, 16'd40930, 16'd57598, 16'd57703, 16'd42516, 16'd28290, 16'd50813, 16'd38129, 16'd48225, 16'd9447, 16'd43035, 16'd49954, 16'd19813, 16'd20547, 16'd48271, 16'd17195, 16'd22967, 16'd11903, 16'd51935, 16'd63662, 16'd10268});
	test_expansion(128'h528b6fba2454318fcad8dad255093251, {16'd64794, 16'd16274, 16'd13110, 16'd61875, 16'd57997, 16'd31270, 16'd2539, 16'd33981, 16'd3396, 16'd8324, 16'd5681, 16'd6781, 16'd28825, 16'd12411, 16'd55153, 16'd52428, 16'd30598, 16'd34034, 16'd29674, 16'd18944, 16'd11780, 16'd42038, 16'd42142, 16'd30111, 16'd51766, 16'd12492});
	test_expansion(128'h8c18aa6e87852d794bfaa43bfd4b151a, {16'd23840, 16'd5344, 16'd16096, 16'd13633, 16'd46186, 16'd59330, 16'd22013, 16'd11583, 16'd32208, 16'd1531, 16'd36635, 16'd62992, 16'd33107, 16'd28174, 16'd335, 16'd52780, 16'd13400, 16'd30281, 16'd35820, 16'd63349, 16'd56631, 16'd40204, 16'd50327, 16'd24349, 16'd51981, 16'd11908});
	test_expansion(128'hae178ccaed6614e42c83c022e037dd41, {16'd36310, 16'd37554, 16'd51108, 16'd4781, 16'd50896, 16'd8776, 16'd56466, 16'd8799, 16'd24162, 16'd31134, 16'd23765, 16'd51196, 16'd14959, 16'd50980, 16'd34606, 16'd18605, 16'd48697, 16'd16270, 16'd36192, 16'd8872, 16'd61876, 16'd47364, 16'd65117, 16'd36991, 16'd25585, 16'd7344});
	test_expansion(128'hbca4575e9f011a68700256428660f04e, {16'd4377, 16'd8130, 16'd17642, 16'd13271, 16'd61164, 16'd32971, 16'd2500, 16'd32321, 16'd31240, 16'd13911, 16'd41589, 16'd59380, 16'd57489, 16'd65098, 16'd13345, 16'd16831, 16'd17121, 16'd17192, 16'd65072, 16'd23717, 16'd3119, 16'd26659, 16'd32115, 16'd18675, 16'd20119, 16'd8300});
	test_expansion(128'ha5ae1e618d034c0bab4e33e77ca2d9da, {16'd49398, 16'd27489, 16'd40110, 16'd4852, 16'd18844, 16'd29816, 16'd14687, 16'd62023, 16'd33812, 16'd4666, 16'd64152, 16'd22496, 16'd29353, 16'd17125, 16'd4875, 16'd11541, 16'd43986, 16'd3560, 16'd61244, 16'd24552, 16'd4082, 16'd60931, 16'd668, 16'd37891, 16'd18615, 16'd59978});
	test_expansion(128'heb2774e8dfa83193b9252ad9f42a818f, {16'd15077, 16'd22143, 16'd45296, 16'd64067, 16'd48197, 16'd2206, 16'd62498, 16'd45566, 16'd1274, 16'd7457, 16'd17495, 16'd56451, 16'd21477, 16'd42500, 16'd26499, 16'd46035, 16'd17430, 16'd16432, 16'd28118, 16'd60100, 16'd31298, 16'd36139, 16'd59261, 16'd33141, 16'd46622, 16'd1021});
	test_expansion(128'h386d17810b6d9c1df193659e9c4f5ab2, {16'd9566, 16'd7030, 16'd60415, 16'd30124, 16'd64158, 16'd62375, 16'd45568, 16'd28588, 16'd35829, 16'd16447, 16'd33086, 16'd19780, 16'd6017, 16'd35689, 16'd9038, 16'd14780, 16'd29958, 16'd26588, 16'd60585, 16'd10981, 16'd52342, 16'd32641, 16'd58996, 16'd20629, 16'd21069, 16'd55816});
	test_expansion(128'h588a173f2c63b75d2a5b8054afff98d1, {16'd55119, 16'd56379, 16'd56525, 16'd58919, 16'd36414, 16'd33993, 16'd868, 16'd69, 16'd54705, 16'd21031, 16'd56358, 16'd34301, 16'd44771, 16'd9943, 16'd24470, 16'd20242, 16'd7747, 16'd49614, 16'd18915, 16'd57912, 16'd28482, 16'd53798, 16'd38774, 16'd14079, 16'd36879, 16'd58899});
	test_expansion(128'h857b65fef20f2b623459cea83617f6be, {16'd41974, 16'd64282, 16'd9058, 16'd13143, 16'd32617, 16'd32120, 16'd63364, 16'd62717, 16'd16186, 16'd30524, 16'd29296, 16'd62407, 16'd657, 16'd50245, 16'd27082, 16'd35918, 16'd42928, 16'd31126, 16'd14071, 16'd13150, 16'd55041, 16'd9689, 16'd42155, 16'd5867, 16'd21098, 16'd35240});
	test_expansion(128'hfbf4e0419452859045c7e78c1b14fbeb, {16'd38378, 16'd10023, 16'd36480, 16'd53694, 16'd11020, 16'd61133, 16'd44913, 16'd41937, 16'd35579, 16'd7696, 16'd18037, 16'd18956, 16'd39703, 16'd46701, 16'd19083, 16'd36796, 16'd17781, 16'd50072, 16'd26190, 16'd40881, 16'd9001, 16'd54242, 16'd15072, 16'd44555, 16'd31077, 16'd8852});
	test_expansion(128'h92b72907cef5b2d9abceb2916277aa7d, {16'd18523, 16'd60358, 16'd41902, 16'd23060, 16'd26113, 16'd63121, 16'd39410, 16'd20448, 16'd36833, 16'd39134, 16'd61970, 16'd19987, 16'd44456, 16'd41404, 16'd13174, 16'd15231, 16'd34582, 16'd41980, 16'd3142, 16'd22806, 16'd2127, 16'd16280, 16'd18207, 16'd19405, 16'd15027, 16'd60447});
	test_expansion(128'h4332c514335b9b6b9f891429c5244b62, {16'd13473, 16'd56945, 16'd6626, 16'd21574, 16'd8091, 16'd18514, 16'd35566, 16'd33957, 16'd4944, 16'd18899, 16'd61327, 16'd20290, 16'd26674, 16'd3213, 16'd43593, 16'd7463, 16'd35239, 16'd30890, 16'd33883, 16'd56743, 16'd34720, 16'd58241, 16'd58958, 16'd55353, 16'd22288, 16'd45639});
	test_expansion(128'he5a717767745237561d8a368a2add0ab, {16'd1168, 16'd56132, 16'd15268, 16'd3318, 16'd6308, 16'd16165, 16'd55412, 16'd54464, 16'd50523, 16'd847, 16'd48030, 16'd36500, 16'd59947, 16'd32780, 16'd14642, 16'd15287, 16'd16481, 16'd52927, 16'd56243, 16'd8725, 16'd20884, 16'd26971, 16'd59524, 16'd26564, 16'd48000, 16'd43146});
	test_expansion(128'h6e48616525fe13204a8bbd7f77933da7, {16'd4903, 16'd23506, 16'd56982, 16'd60977, 16'd31912, 16'd25761, 16'd55658, 16'd30484, 16'd40724, 16'd39977, 16'd35262, 16'd32807, 16'd54697, 16'd27269, 16'd61371, 16'd4947, 16'd13195, 16'd46157, 16'd38969, 16'd45904, 16'd44454, 16'd64379, 16'd6732, 16'd60467, 16'd41340, 16'd25022});
	test_expansion(128'hbf07605a7cab73f1d0671b8d5465696c, {16'd60792, 16'd37236, 16'd11780, 16'd15936, 16'd12626, 16'd51877, 16'd56227, 16'd37254, 16'd139, 16'd51566, 16'd38833, 16'd17563, 16'd31933, 16'd44979, 16'd42721, 16'd46516, 16'd20847, 16'd10847, 16'd23662, 16'd11896, 16'd5683, 16'd56278, 16'd62697, 16'd40116, 16'd8892, 16'd19024});
	test_expansion(128'h9984aca1a5ed62f79c78e3c90f539e50, {16'd13916, 16'd51152, 16'd53025, 16'd64387, 16'd12042, 16'd60154, 16'd47560, 16'd12692, 16'd16532, 16'd65084, 16'd20356, 16'd49226, 16'd10209, 16'd22852, 16'd18641, 16'd59426, 16'd28233, 16'd31446, 16'd35677, 16'd12174, 16'd45809, 16'd47455, 16'd3453, 16'd9266, 16'd30595, 16'd56597});
	test_expansion(128'hd5b84800f979421f8f5357d6f370d2c0, {16'd55794, 16'd5672, 16'd43010, 16'd1516, 16'd36943, 16'd61365, 16'd21352, 16'd45659, 16'd23779, 16'd52017, 16'd20444, 16'd44414, 16'd51299, 16'd50161, 16'd47786, 16'd20978, 16'd51062, 16'd28761, 16'd52205, 16'd44304, 16'd60389, 16'd14982, 16'd1392, 16'd29496, 16'd54393, 16'd39530});
	test_expansion(128'h1537a749988b5786872ba23ffe801585, {16'd6023, 16'd36675, 16'd60311, 16'd16888, 16'd21172, 16'd11437, 16'd31766, 16'd24706, 16'd873, 16'd51834, 16'd9875, 16'd23173, 16'd16611, 16'd35753, 16'd47763, 16'd26190, 16'd23898, 16'd44912, 16'd18968, 16'd65312, 16'd47178, 16'd39669, 16'd34187, 16'd63840, 16'd49607, 16'd53591});
	test_expansion(128'h2d97dfb8dfda3e4d81731fcbb96f7621, {16'd36795, 16'd32860, 16'd52403, 16'd49363, 16'd59037, 16'd7197, 16'd32224, 16'd18282, 16'd16188, 16'd26979, 16'd28637, 16'd60037, 16'd12457, 16'd486, 16'd17423, 16'd39851, 16'd11837, 16'd38798, 16'd64590, 16'd38658, 16'd26778, 16'd18016, 16'd32656, 16'd65348, 16'd39676, 16'd10760});
	test_expansion(128'he8edac96f91e0cee30c3be8f06304dfe, {16'd2691, 16'd39585, 16'd34273, 16'd54472, 16'd58637, 16'd2815, 16'd28320, 16'd60189, 16'd52881, 16'd46646, 16'd20539, 16'd12508, 16'd62482, 16'd55895, 16'd21460, 16'd11390, 16'd7169, 16'd37865, 16'd26085, 16'd40266, 16'd53303, 16'd18624, 16'd56770, 16'd24187, 16'd35346, 16'd24701});
	test_expansion(128'ha636fe5e78580cc8de7726fb885f8733, {16'd54138, 16'd40986, 16'd44353, 16'd42492, 16'd38047, 16'd47899, 16'd50570, 16'd26806, 16'd30115, 16'd9718, 16'd15250, 16'd26532, 16'd18902, 16'd21743, 16'd44951, 16'd43037, 16'd65139, 16'd38085, 16'd58473, 16'd65192, 16'd11982, 16'd34298, 16'd45703, 16'd22226, 16'd31460, 16'd26880});
	test_expansion(128'h34ffba270ac0af21621f1e93cad6da3f, {16'd51537, 16'd41886, 16'd26009, 16'd56590, 16'd49116, 16'd34497, 16'd3449, 16'd27595, 16'd47752, 16'd15084, 16'd24339, 16'd4757, 16'd64869, 16'd43121, 16'd3102, 16'd5722, 16'd52280, 16'd2540, 16'd15694, 16'd46741, 16'd15797, 16'd28013, 16'd48382, 16'd42420, 16'd46853, 16'd10180});
	test_expansion(128'h68b5ef8ca7b023325b5f6535db8698b2, {16'd32762, 16'd61755, 16'd10386, 16'd57587, 16'd39301, 16'd41140, 16'd10695, 16'd59026, 16'd50384, 16'd33398, 16'd38163, 16'd38870, 16'd3202, 16'd10361, 16'd43193, 16'd9759, 16'd49488, 16'd51680, 16'd41266, 16'd30454, 16'd65101, 16'd27525, 16'd23532, 16'd48564, 16'd27446, 16'd64920});
	test_expansion(128'h679f424c8e93d804c2a3dcafe610eeeb, {16'd34383, 16'd31436, 16'd25104, 16'd62871, 16'd56183, 16'd44446, 16'd36885, 16'd16330, 16'd24323, 16'd12810, 16'd39413, 16'd37856, 16'd35174, 16'd6970, 16'd62891, 16'd53646, 16'd35862, 16'd25965, 16'd4962, 16'd23125, 16'd3002, 16'd43044, 16'd48436, 16'd15722, 16'd3427, 16'd27229});
	test_expansion(128'ha4aad9cbc1ca56e9fb58c0bde66ffc15, {16'd15798, 16'd9504, 16'd38975, 16'd4760, 16'd34268, 16'd924, 16'd49127, 16'd59808, 16'd25388, 16'd20027, 16'd34657, 16'd2817, 16'd54091, 16'd24429, 16'd11964, 16'd5557, 16'd19817, 16'd22678, 16'd12103, 16'd23656, 16'd1888, 16'd34502, 16'd33834, 16'd432, 16'd42780, 16'd28423});
	test_expansion(128'hf21bd26b8718d2ad71be64d48530271f, {16'd52783, 16'd51266, 16'd28107, 16'd3837, 16'd10038, 16'd52821, 16'd27212, 16'd42935, 16'd62058, 16'd10661, 16'd38640, 16'd57208, 16'd52786, 16'd32632, 16'd4037, 16'd40240, 16'd7871, 16'd5292, 16'd43118, 16'd54181, 16'd51481, 16'd18506, 16'd3295, 16'd46527, 16'd18447, 16'd38781});
	test_expansion(128'had6a5a8a95719d293fe3e5bcba4bd891, {16'd42466, 16'd22281, 16'd50367, 16'd33357, 16'd9754, 16'd398, 16'd58569, 16'd57527, 16'd20851, 16'd998, 16'd41987, 16'd4748, 16'd29468, 16'd51077, 16'd23898, 16'd13154, 16'd7409, 16'd53042, 16'd32933, 16'd18900, 16'd36104, 16'd47843, 16'd60949, 16'd6225, 16'd7508, 16'd8448});
	test_expansion(128'hf0d180dbac46c50a87737e4d51f82c20, {16'd18607, 16'd32933, 16'd14954, 16'd19122, 16'd11914, 16'd51966, 16'd18966, 16'd25706, 16'd5537, 16'd51961, 16'd50072, 16'd35628, 16'd33338, 16'd16375, 16'd49564, 16'd34756, 16'd46404, 16'd18592, 16'd9487, 16'd44895, 16'd56035, 16'd43908, 16'd4215, 16'd18404, 16'd6670, 16'd24487});
	test_expansion(128'hf2ee893834d7ac532b741f2212d7f98b, {16'd28842, 16'd6511, 16'd13402, 16'd31554, 16'd63939, 16'd15122, 16'd17775, 16'd39681, 16'd3934, 16'd5550, 16'd59356, 16'd48493, 16'd57400, 16'd1610, 16'd46822, 16'd50316, 16'd56485, 16'd37722, 16'd10112, 16'd22384, 16'd28473, 16'd11431, 16'd13288, 16'd54359, 16'd26945, 16'd25896});
	test_expansion(128'hea2e030ab01e57798b92643e2e231541, {16'd12, 16'd56169, 16'd53549, 16'd39455, 16'd42002, 16'd10164, 16'd12973, 16'd25948, 16'd64594, 16'd5348, 16'd8039, 16'd34656, 16'd4085, 16'd42852, 16'd63154, 16'd32454, 16'd15781, 16'd60070, 16'd46901, 16'd47492, 16'd23996, 16'd37047, 16'd45892, 16'd55458, 16'd3803, 16'd45784});
	test_expansion(128'h75eb838484961feea71f6014ae87c826, {16'd30423, 16'd49012, 16'd63838, 16'd17734, 16'd43417, 16'd1226, 16'd29936, 16'd16937, 16'd29088, 16'd34351, 16'd10438, 16'd32935, 16'd51942, 16'd20831, 16'd22248, 16'd31880, 16'd54543, 16'd24038, 16'd18973, 16'd40921, 16'd44668, 16'd61705, 16'd56818, 16'd49345, 16'd65122, 16'd8494});
	test_expansion(128'h498d35fe396bc7fb2c974236bdce9147, {16'd38730, 16'd57005, 16'd33667, 16'd49454, 16'd42842, 16'd58373, 16'd18363, 16'd28782, 16'd17909, 16'd6261, 16'd25134, 16'd21696, 16'd46143, 16'd19851, 16'd53653, 16'd33003, 16'd30362, 16'd13414, 16'd10838, 16'd53573, 16'd32433, 16'd48653, 16'd11819, 16'd11418, 16'd41448, 16'd8078});
	test_expansion(128'h9b69bd73b07e0bcce60a639066d1a072, {16'd48483, 16'd28066, 16'd30661, 16'd42913, 16'd47719, 16'd25409, 16'd10927, 16'd32788, 16'd21526, 16'd12985, 16'd32366, 16'd12350, 16'd39763, 16'd56666, 16'd13882, 16'd455, 16'd64436, 16'd42599, 16'd997, 16'd2582, 16'd29450, 16'd483, 16'd30490, 16'd36871, 16'd40804, 16'd32561});
	test_expansion(128'h3b1d775bf942a84cd3e8fc283f804cf0, {16'd47605, 16'd44837, 16'd49173, 16'd15671, 16'd12300, 16'd13317, 16'd34974, 16'd38320, 16'd27692, 16'd27573, 16'd41127, 16'd44310, 16'd12629, 16'd604, 16'd60429, 16'd5028, 16'd7552, 16'd14277, 16'd10284, 16'd58082, 16'd54047, 16'd45328, 16'd24090, 16'd54362, 16'd35074, 16'd33763});
	test_expansion(128'h9201d368d03a7eaa399ba5004a76145d, {16'd59200, 16'd38471, 16'd54970, 16'd49831, 16'd18980, 16'd27974, 16'd25679, 16'd41122, 16'd51486, 16'd46579, 16'd33310, 16'd15210, 16'd41409, 16'd65486, 16'd13294, 16'd25661, 16'd40352, 16'd5883, 16'd19376, 16'd22521, 16'd2185, 16'd48330, 16'd53861, 16'd28837, 16'd31638, 16'd6512});
	test_expansion(128'hae28bbbe78d1019239c69897f166b111, {16'd42420, 16'd12750, 16'd51930, 16'd4190, 16'd29728, 16'd64261, 16'd35071, 16'd9252, 16'd26342, 16'd55638, 16'd41204, 16'd10369, 16'd37698, 16'd14206, 16'd60711, 16'd6426, 16'd34639, 16'd51581, 16'd31362, 16'd46379, 16'd38979, 16'd63111, 16'd5514, 16'd28812, 16'd32490, 16'd44889});
	test_expansion(128'hf4cab8e7b75bbef6ee84c924c80291d6, {16'd43652, 16'd49521, 16'd11811, 16'd5713, 16'd233, 16'd54902, 16'd28592, 16'd10899, 16'd36717, 16'd48330, 16'd55530, 16'd46709, 16'd62531, 16'd6789, 16'd48807, 16'd47573, 16'd53377, 16'd51316, 16'd9299, 16'd27686, 16'd33923, 16'd49055, 16'd59749, 16'd49958, 16'd49008, 16'd23776});
	test_expansion(128'hbe573f0f55452f8e0cb5d735fe499ada, {16'd5990, 16'd47387, 16'd28628, 16'd19494, 16'd29974, 16'd30539, 16'd1008, 16'd57327, 16'd19423, 16'd54322, 16'd1002, 16'd45055, 16'd64135, 16'd26641, 16'd30309, 16'd17921, 16'd384, 16'd28940, 16'd40164, 16'd34685, 16'd37488, 16'd29351, 16'd37969, 16'd10639, 16'd22498, 16'd23704});
	test_expansion(128'h4da64a685360afeae39947814f186f8b, {16'd16917, 16'd30862, 16'd44912, 16'd63892, 16'd60108, 16'd7241, 16'd7722, 16'd61184, 16'd8886, 16'd23226, 16'd60598, 16'd52327, 16'd31073, 16'd5923, 16'd7518, 16'd11906, 16'd23031, 16'd9505, 16'd41751, 16'd39277, 16'd53890, 16'd51841, 16'd58101, 16'd64652, 16'd28053, 16'd20384});
	test_expansion(128'hf1940bd9fb7f8c3169edb96b2f880f78, {16'd6079, 16'd1485, 16'd31175, 16'd20774, 16'd58342, 16'd15632, 16'd49859, 16'd36811, 16'd13683, 16'd33222, 16'd63315, 16'd62516, 16'd34204, 16'd49265, 16'd8273, 16'd56527, 16'd42451, 16'd24581, 16'd28697, 16'd52217, 16'd4371, 16'd49741, 16'd47296, 16'd30059, 16'd31845, 16'd47444});
	test_expansion(128'h221c97654afa71e297a46e9339cd0cba, {16'd3236, 16'd38364, 16'd59175, 16'd158, 16'd35289, 16'd29987, 16'd21314, 16'd32292, 16'd4774, 16'd48111, 16'd9834, 16'd51874, 16'd60059, 16'd1016, 16'd3805, 16'd49066, 16'd34082, 16'd35980, 16'd27305, 16'd65352, 16'd12516, 16'd55156, 16'd62002, 16'd11706, 16'd2421, 16'd25642});
	test_expansion(128'haf2d869d01f7867737a787dd7a981737, {16'd52871, 16'd35121, 16'd50230, 16'd61478, 16'd25598, 16'd62165, 16'd63532, 16'd55059, 16'd19757, 16'd29188, 16'd27036, 16'd41507, 16'd39903, 16'd31792, 16'd51417, 16'd30637, 16'd1723, 16'd9329, 16'd24894, 16'd9866, 16'd53275, 16'd26068, 16'd54147, 16'd10775, 16'd9574, 16'd43903});
	test_expansion(128'h760c23d96cfd23ec5a97c9b16beeff6f, {16'd2625, 16'd37370, 16'd56177, 16'd9859, 16'd39386, 16'd9210, 16'd45896, 16'd28850, 16'd45683, 16'd17237, 16'd52636, 16'd65013, 16'd52726, 16'd61629, 16'd64218, 16'd50513, 16'd60097, 16'd45532, 16'd10599, 16'd1450, 16'd31013, 16'd41093, 16'd3484, 16'd5153, 16'd52277, 16'd53800});
	test_expansion(128'hecb8c46b1082640f800dc93d48b6f33d, {16'd46933, 16'd60609, 16'd42000, 16'd55147, 16'd26372, 16'd3252, 16'd23838, 16'd50739, 16'd16572, 16'd47337, 16'd39136, 16'd9099, 16'd12067, 16'd19804, 16'd34854, 16'd40675, 16'd8609, 16'd59953, 16'd64770, 16'd31688, 16'd62922, 16'd41767, 16'd23106, 16'd56023, 16'd45769, 16'd6247});
	test_expansion(128'hd998a6b6a71feaf34c866224d37b1d6f, {16'd29429, 16'd39485, 16'd45021, 16'd26032, 16'd9300, 16'd34419, 16'd49273, 16'd58997, 16'd10312, 16'd50183, 16'd10991, 16'd59430, 16'd27696, 16'd17782, 16'd34125, 16'd396, 16'd13442, 16'd25741, 16'd1209, 16'd22084, 16'd57383, 16'd24219, 16'd22443, 16'd12588, 16'd6843, 16'd24651});
	test_expansion(128'h1a18fced2edd9e92156cd99d27f40014, {16'd42681, 16'd26294, 16'd64676, 16'd34658, 16'd37698, 16'd50361, 16'd19405, 16'd4251, 16'd29577, 16'd16257, 16'd55211, 16'd41234, 16'd39817, 16'd9152, 16'd24300, 16'd36342, 16'd55765, 16'd13557, 16'd24669, 16'd63126, 16'd52755, 16'd48161, 16'd53461, 16'd21011, 16'd62545, 16'd65497});
	test_expansion(128'h43d536054cd7397db8b427fad65e0163, {16'd46687, 16'd58095, 16'd10545, 16'd8631, 16'd50708, 16'd23307, 16'd45839, 16'd57955, 16'd1340, 16'd60203, 16'd19238, 16'd45670, 16'd17561, 16'd14013, 16'd63676, 16'd28841, 16'd58849, 16'd45685, 16'd13240, 16'd64656, 16'd30774, 16'd15986, 16'd39544, 16'd37769, 16'd8850, 16'd8762});
	test_expansion(128'h3dd10ea92b6712732b385d0a07f6fccc, {16'd19223, 16'd32305, 16'd34838, 16'd51487, 16'd39380, 16'd39667, 16'd18397, 16'd59784, 16'd19317, 16'd15042, 16'd19974, 16'd36758, 16'd36748, 16'd2360, 16'd16835, 16'd37845, 16'd38068, 16'd59283, 16'd48234, 16'd62737, 16'd57537, 16'd10343, 16'd17597, 16'd47089, 16'd10463, 16'd65487});
	test_expansion(128'hb00955bf94a7ead2bc0d94990c8e09d7, {16'd19224, 16'd54138, 16'd50490, 16'd32293, 16'd38388, 16'd21982, 16'd47307, 16'd30455, 16'd56704, 16'd3201, 16'd49887, 16'd51749, 16'd49818, 16'd38461, 16'd59350, 16'd16321, 16'd9254, 16'd33873, 16'd59538, 16'd9202, 16'd47173, 16'd45295, 16'd49758, 16'd1327, 16'd29664, 16'd63587});
	test_expansion(128'h4ee317d6436853aade4cc69133f1e045, {16'd42252, 16'd24297, 16'd14527, 16'd7244, 16'd15421, 16'd18299, 16'd65286, 16'd34907, 16'd53590, 16'd35541, 16'd21421, 16'd5244, 16'd24039, 16'd38767, 16'd50469, 16'd24605, 16'd65301, 16'd2640, 16'd63166, 16'd52564, 16'd33406, 16'd15272, 16'd40406, 16'd7020, 16'd48392, 16'd36386});
	test_expansion(128'h43e9ec796c3b3034d7ab450a1c412485, {16'd13549, 16'd13138, 16'd8159, 16'd20047, 16'd26545, 16'd41996, 16'd48312, 16'd26047, 16'd21484, 16'd3501, 16'd44346, 16'd2284, 16'd44819, 16'd13187, 16'd7153, 16'd1735, 16'd4697, 16'd32918, 16'd46084, 16'd6155, 16'd24628, 16'd10814, 16'd34267, 16'd55201, 16'd50134, 16'd26181});
	test_expansion(128'hfa0606ae5b2d45d606a5f251a5e05092, {16'd34116, 16'd56664, 16'd11616, 16'd49199, 16'd49770, 16'd36685, 16'd18632, 16'd50467, 16'd27055, 16'd55915, 16'd34608, 16'd31830, 16'd63280, 16'd21990, 16'd58055, 16'd37690, 16'd27353, 16'd61298, 16'd24657, 16'd63352, 16'd35617, 16'd15858, 16'd52002, 16'd22351, 16'd4008, 16'd29170});
	test_expansion(128'h3b95c7ff25464c8f3e89dea79f2d2750, {16'd58342, 16'd23919, 16'd61616, 16'd48185, 16'd49340, 16'd26919, 16'd30811, 16'd64503, 16'd50803, 16'd24306, 16'd47329, 16'd16881, 16'd20418, 16'd17621, 16'd6807, 16'd29937, 16'd2851, 16'd56576, 16'd44716, 16'd17423, 16'd22299, 16'd31785, 16'd59356, 16'd52602, 16'd29175, 16'd52611});
	test_expansion(128'h85fa48fd95dfc9ddf43b23e069e68f62, {16'd46027, 16'd8141, 16'd13648, 16'd44516, 16'd27007, 16'd11320, 16'd31541, 16'd41942, 16'd5121, 16'd37888, 16'd32260, 16'd47211, 16'd7300, 16'd15322, 16'd48127, 16'd589, 16'd55536, 16'd15483, 16'd17417, 16'd18791, 16'd37944, 16'd23615, 16'd52191, 16'd28185, 16'd53578, 16'd16654});
	test_expansion(128'hb14f962a258c6fc9c7f9170e1b89ff0b, {16'd16898, 16'd307, 16'd28170, 16'd38496, 16'd40525, 16'd42776, 16'd30673, 16'd23079, 16'd8807, 16'd27276, 16'd59767, 16'd42812, 16'd63685, 16'd31482, 16'd12748, 16'd16155, 16'd57980, 16'd15039, 16'd10119, 16'd62958, 16'd52706, 16'd55624, 16'd14087, 16'd36617, 16'd57255, 16'd36915});
	test_expansion(128'h09e12db4dbcd9ea5f385055dcf049c61, {16'd6981, 16'd59256, 16'd29267, 16'd39814, 16'd54383, 16'd31959, 16'd21774, 16'd52262, 16'd51403, 16'd61242, 16'd30446, 16'd46090, 16'd36486, 16'd10843, 16'd15389, 16'd55090, 16'd54537, 16'd25864, 16'd62439, 16'd50659, 16'd52315, 16'd56474, 16'd45501, 16'd58975, 16'd27459, 16'd23964});
	test_expansion(128'h02edc1db83b8c5d1139fa824f1d22348, {16'd45481, 16'd12048, 16'd42524, 16'd15604, 16'd39592, 16'd19067, 16'd36159, 16'd30493, 16'd15007, 16'd7029, 16'd46401, 16'd54267, 16'd36939, 16'd62211, 16'd3275, 16'd38501, 16'd19290, 16'd43033, 16'd18792, 16'd23900, 16'd2050, 16'd64597, 16'd17658, 16'd41, 16'd40874, 16'd3890});
	test_expansion(128'h7f7f474deabe4e8f34e19c3a3674141b, {16'd38682, 16'd60605, 16'd47448, 16'd4858, 16'd58965, 16'd12208, 16'd35269, 16'd29086, 16'd8690, 16'd33048, 16'd16475, 16'd64584, 16'd62863, 16'd28214, 16'd9858, 16'd40568, 16'd51697, 16'd43450, 16'd8840, 16'd55356, 16'd15859, 16'd31204, 16'd41644, 16'd2733, 16'd60579, 16'd48601});
	test_expansion(128'hf7ff5887eae1b0262c14839868947677, {16'd31195, 16'd35191, 16'd48772, 16'd54599, 16'd59159, 16'd25853, 16'd13269, 16'd48237, 16'd24579, 16'd58837, 16'd21462, 16'd6011, 16'd9634, 16'd6150, 16'd47523, 16'd5766, 16'd64935, 16'd14777, 16'd17499, 16'd16788, 16'd7887, 16'd30745, 16'd26723, 16'd10326, 16'd16830, 16'd34108});
	test_expansion(128'hc3e143e5fabae198001e4b2ba219cceb, {16'd3805, 16'd18878, 16'd35403, 16'd4841, 16'd7032, 16'd64618, 16'd45640, 16'd7184, 16'd42171, 16'd53187, 16'd59914, 16'd12210, 16'd54102, 16'd4803, 16'd54728, 16'd33298, 16'd47084, 16'd24091, 16'd26505, 16'd8254, 16'd41013, 16'd14648, 16'd40578, 16'd55547, 16'd29402, 16'd4738});
	test_expansion(128'h36cadaae31743f3a29f4ce4f76ddfa8f, {16'd15872, 16'd62803, 16'd27558, 16'd14033, 16'd8864, 16'd57850, 16'd64985, 16'd42793, 16'd18700, 16'd52849, 16'd39399, 16'd43188, 16'd15935, 16'd55879, 16'd45951, 16'd22622, 16'd48783, 16'd57802, 16'd32782, 16'd29540, 16'd14351, 16'd26027, 16'd29962, 16'd54391, 16'd23071, 16'd48363});
	test_expansion(128'hcda25c56d451952b096f3627665a6c31, {16'd41205, 16'd58311, 16'd34901, 16'd32193, 16'd45730, 16'd55603, 16'd43796, 16'd52088, 16'd5630, 16'd42298, 16'd62638, 16'd29545, 16'd37541, 16'd57938, 16'd52071, 16'd2675, 16'd53991, 16'd60372, 16'd57030, 16'd7482, 16'd5644, 16'd63236, 16'd60313, 16'd41373, 16'd8488, 16'd43085});
	test_expansion(128'h165b74756ce0d4ee71b9ba1048bf6c0d, {16'd57644, 16'd17409, 16'd15182, 16'd48740, 16'd20773, 16'd34337, 16'd21783, 16'd24205, 16'd26365, 16'd15809, 16'd471, 16'd34615, 16'd29040, 16'd30935, 16'd28776, 16'd23626, 16'd32517, 16'd37693, 16'd64165, 16'd8965, 16'd30453, 16'd50059, 16'd36558, 16'd8632, 16'd50246, 16'd42984});
	test_expansion(128'h7c9658fef7942b5c8e61e3f433b3d22c, {16'd56896, 16'd39748, 16'd31887, 16'd41735, 16'd28008, 16'd19239, 16'd65228, 16'd60420, 16'd46843, 16'd23358, 16'd41501, 16'd64601, 16'd57973, 16'd4011, 16'd15897, 16'd8483, 16'd7186, 16'd31413, 16'd18952, 16'd37367, 16'd59646, 16'd34214, 16'd65202, 16'd44996, 16'd56271, 16'd45229});
	test_expansion(128'h5dc61a07211122051bd593119f890b4b, {16'd36668, 16'd18888, 16'd15182, 16'd17753, 16'd1962, 16'd62595, 16'd20437, 16'd59987, 16'd60799, 16'd14047, 16'd63716, 16'd34197, 16'd46706, 16'd15446, 16'd55971, 16'd53964, 16'd11954, 16'd55413, 16'd23401, 16'd38563, 16'd45887, 16'd63322, 16'd23440, 16'd36290, 16'd33528, 16'd36606});
	test_expansion(128'h73de34862e2b3a659cf33df18a008456, {16'd25027, 16'd17773, 16'd15147, 16'd2711, 16'd54483, 16'd37281, 16'd13850, 16'd17142, 16'd30346, 16'd39203, 16'd45489, 16'd52383, 16'd52060, 16'd9764, 16'd55894, 16'd19255, 16'd62659, 16'd6540, 16'd9595, 16'd58370, 16'd22089, 16'd9709, 16'd53945, 16'd34115, 16'd9320, 16'd11661});
	test_expansion(128'h81399db4f5bbf20be23bcff2c0ba4ca5, {16'd50321, 16'd37864, 16'd36760, 16'd29526, 16'd47414, 16'd55226, 16'd16044, 16'd43875, 16'd38409, 16'd4330, 16'd49595, 16'd63023, 16'd14570, 16'd13014, 16'd40126, 16'd45855, 16'd18771, 16'd21031, 16'd6442, 16'd47635, 16'd64426, 16'd36515, 16'd60364, 16'd1986, 16'd8782, 16'd12110});
	test_expansion(128'h382092d452d5bf2911b0f5fb728c9c8a, {16'd29067, 16'd54514, 16'd2900, 16'd53193, 16'd11955, 16'd1160, 16'd17411, 16'd25607, 16'd29373, 16'd30922, 16'd34971, 16'd41960, 16'd45228, 16'd5157, 16'd49749, 16'd53888, 16'd38253, 16'd52660, 16'd21908, 16'd4540, 16'd11941, 16'd57479, 16'd21183, 16'd43397, 16'd23944, 16'd37504});
	test_expansion(128'h6ffca4c4d1b2abcdd4c6287f9a3e545b, {16'd57422, 16'd60215, 16'd30633, 16'd35619, 16'd19292, 16'd21190, 16'd37909, 16'd51882, 16'd14255, 16'd46789, 16'd44090, 16'd46664, 16'd3087, 16'd13958, 16'd21644, 16'd30376, 16'd5907, 16'd53217, 16'd51772, 16'd2829, 16'd33466, 16'd11283, 16'd15966, 16'd59310, 16'd33004, 16'd47178});
	test_expansion(128'h9ae1c033b4b4b48b6bb5b3a3b6b5129e, {16'd47113, 16'd21347, 16'd22690, 16'd778, 16'd36656, 16'd28282, 16'd21811, 16'd32104, 16'd50478, 16'd53168, 16'd31390, 16'd15200, 16'd11089, 16'd6383, 16'd16121, 16'd53333, 16'd32657, 16'd39827, 16'd25176, 16'd1010, 16'd55550, 16'd41151, 16'd62819, 16'd60830, 16'd41367, 16'd38024});
	test_expansion(128'hb711a22ec14924e6aa27d98d44c4daca, {16'd35444, 16'd57831, 16'd51251, 16'd25187, 16'd11273, 16'd10183, 16'd47602, 16'd49974, 16'd42519, 16'd32878, 16'd56760, 16'd51574, 16'd33550, 16'd5753, 16'd23325, 16'd4643, 16'd47543, 16'd39579, 16'd4706, 16'd35867, 16'd20365, 16'd3713, 16'd5530, 16'd38817, 16'd3602, 16'd7027});
	test_expansion(128'h53e1c8b896dad5af98481fc245c856e2, {16'd39492, 16'd24799, 16'd59577, 16'd12194, 16'd37231, 16'd3401, 16'd64012, 16'd19165, 16'd57536, 16'd1422, 16'd31793, 16'd2140, 16'd15564, 16'd33657, 16'd27404, 16'd18822, 16'd44869, 16'd9442, 16'd27554, 16'd6638, 16'd46739, 16'd22235, 16'd26664, 16'd9958, 16'd42110, 16'd42174});
	test_expansion(128'h98b773d6a908c548e4ac21301abffb20, {16'd41354, 16'd47154, 16'd9532, 16'd47157, 16'd23788, 16'd26344, 16'd35460, 16'd45009, 16'd23440, 16'd33986, 16'd62845, 16'd32840, 16'd42860, 16'd5350, 16'd28448, 16'd36544, 16'd47396, 16'd9038, 16'd21508, 16'd28377, 16'd12723, 16'd9930, 16'd50486, 16'd9608, 16'd39334, 16'd53828});
	test_expansion(128'h18ba1bcc1c38c438fa3f6aa96c7e8b80, {16'd10685, 16'd6604, 16'd30849, 16'd40492, 16'd6524, 16'd22777, 16'd63729, 16'd47219, 16'd6610, 16'd24577, 16'd62018, 16'd7989, 16'd28610, 16'd15426, 16'd16765, 16'd18362, 16'd2743, 16'd65130, 16'd10592, 16'd62040, 16'd8330, 16'd27640, 16'd10581, 16'd36983, 16'd41758, 16'd5389});
	test_expansion(128'h25d90283a2470149347d602e2262c519, {16'd14161, 16'd62027, 16'd3346, 16'd23286, 16'd58024, 16'd16432, 16'd27606, 16'd8967, 16'd60158, 16'd59722, 16'd18785, 16'd25631, 16'd1254, 16'd43691, 16'd50833, 16'd11747, 16'd37401, 16'd43107, 16'd32888, 16'd27575, 16'd17376, 16'd37550, 16'd2596, 16'd23714, 16'd39365, 16'd8099});
	test_expansion(128'h1e43d1a128b9df929132a93eca37b0de, {16'd31484, 16'd46980, 16'd52648, 16'd59640, 16'd15316, 16'd17658, 16'd56643, 16'd20081, 16'd7992, 16'd48728, 16'd45442, 16'd24678, 16'd57200, 16'd56596, 16'd50767, 16'd64957, 16'd13013, 16'd43525, 16'd49541, 16'd32979, 16'd15298, 16'd63573, 16'd44689, 16'd42933, 16'd61800, 16'd22412});
	test_expansion(128'h913bc87faff2cec684de1e555657a802, {16'd57149, 16'd16490, 16'd44371, 16'd3142, 16'd16768, 16'd11932, 16'd48522, 16'd52597, 16'd48361, 16'd33376, 16'd5890, 16'd14274, 16'd24795, 16'd39005, 16'd54154, 16'd28019, 16'd7893, 16'd52190, 16'd58521, 16'd20209, 16'd6415, 16'd34670, 16'd12907, 16'd53965, 16'd21414, 16'd36544});
	test_expansion(128'h9e455597dac911e2585ec49aadb2864f, {16'd60594, 16'd32744, 16'd26009, 16'd29154, 16'd38251, 16'd18156, 16'd3245, 16'd18325, 16'd16815, 16'd18924, 16'd29907, 16'd61707, 16'd54417, 16'd28264, 16'd56498, 16'd22128, 16'd10198, 16'd40779, 16'd29476, 16'd26405, 16'd56215, 16'd6645, 16'd64091, 16'd30395, 16'd52777, 16'd51424});
	test_expansion(128'hedb1df1b6c24402e3371f16c2c138ee2, {16'd62116, 16'd14917, 16'd27428, 16'd54960, 16'd50811, 16'd15466, 16'd9299, 16'd38171, 16'd56583, 16'd18555, 16'd44165, 16'd47411, 16'd49154, 16'd28014, 16'd9403, 16'd39382, 16'd56773, 16'd33165, 16'd65381, 16'd51702, 16'd5491, 16'd340, 16'd61728, 16'd5852, 16'd54293, 16'd13411});
	test_expansion(128'hbaca85fc95f010a1d3c4e34d2f2ff64c, {16'd56826, 16'd36303, 16'd42248, 16'd48148, 16'd30835, 16'd386, 16'd11357, 16'd19386, 16'd61332, 16'd54267, 16'd964, 16'd47999, 16'd34648, 16'd39486, 16'd24683, 16'd32116, 16'd40702, 16'd62483, 16'd8200, 16'd4066, 16'd23840, 16'd50756, 16'd1463, 16'd45391, 16'd59717, 16'd31823});
	test_expansion(128'hb3a67478c20abb77b2d027cf399d7484, {16'd64297, 16'd49876, 16'd22434, 16'd2387, 16'd51151, 16'd50057, 16'd65198, 16'd9511, 16'd58810, 16'd8794, 16'd65406, 16'd342, 16'd10137, 16'd316, 16'd51510, 16'd33608, 16'd46925, 16'd27232, 16'd7681, 16'd5254, 16'd23702, 16'd59125, 16'd17309, 16'd18943, 16'd56246, 16'd45845});
	test_expansion(128'hf8b0d139e3ece305436209440df20040, {16'd34405, 16'd39555, 16'd9731, 16'd22557, 16'd4030, 16'd8597, 16'd57712, 16'd8896, 16'd10177, 16'd59990, 16'd20593, 16'd19858, 16'd48131, 16'd55036, 16'd25336, 16'd4213, 16'd46207, 16'd615, 16'd23559, 16'd36589, 16'd44766, 16'd38932, 16'd9756, 16'd44933, 16'd13930, 16'd1446});
	test_expansion(128'ha33f657dc75aff8b8ee442698d4329ca, {16'd64371, 16'd62190, 16'd14013, 16'd57292, 16'd5670, 16'd4681, 16'd9116, 16'd30820, 16'd15525, 16'd3336, 16'd57892, 16'd17487, 16'd9604, 16'd25141, 16'd57116, 16'd6959, 16'd46135, 16'd49698, 16'd36280, 16'd22363, 16'd50895, 16'd34023, 16'd57172, 16'd29568, 16'd20857, 16'd263});
	test_expansion(128'h997c60b29c5674fc8fa029f18d45019a, {16'd52600, 16'd35577, 16'd15627, 16'd33979, 16'd56167, 16'd4071, 16'd20617, 16'd22417, 16'd43395, 16'd46696, 16'd60627, 16'd55562, 16'd48135, 16'd18246, 16'd18848, 16'd5274, 16'd55063, 16'd7742, 16'd22504, 16'd129, 16'd18017, 16'd25336, 16'd1117, 16'd35316, 16'd46651, 16'd11877});
	test_expansion(128'hc02d88920ed7f65709b788617b652596, {16'd2804, 16'd19926, 16'd14526, 16'd56922, 16'd49685, 16'd12039, 16'd22551, 16'd12423, 16'd52811, 16'd4197, 16'd63959, 16'd48464, 16'd1790, 16'd50297, 16'd4744, 16'd3766, 16'd47759, 16'd14410, 16'd57281, 16'd28623, 16'd63135, 16'd12650, 16'd8911, 16'd47094, 16'd21707, 16'd6635});
	test_expansion(128'hc777b4009342ed41e4bdccd0f4be5d32, {16'd65107, 16'd39865, 16'd9842, 16'd34596, 16'd23844, 16'd10796, 16'd46999, 16'd17080, 16'd51268, 16'd49140, 16'd26756, 16'd56789, 16'd31803, 16'd9048, 16'd32463, 16'd28863, 16'd27587, 16'd52326, 16'd4521, 16'd18728, 16'd16975, 16'd19047, 16'd61460, 16'd22724, 16'd11733, 16'd2878});
	test_expansion(128'h37d57c00673da880d4609bc3a49c7780, {16'd39310, 16'd62401, 16'd5666, 16'd31986, 16'd29030, 16'd9657, 16'd20733, 16'd60730, 16'd34194, 16'd64087, 16'd57612, 16'd47381, 16'd6982, 16'd11211, 16'd14729, 16'd20581, 16'd47690, 16'd11942, 16'd32632, 16'd60703, 16'd35687, 16'd5659, 16'd2960, 16'd41157, 16'd34792, 16'd14377});
	test_expansion(128'hf193e86fd087a84b152febab2a93a43b, {16'd11018, 16'd54971, 16'd30861, 16'd41179, 16'd21052, 16'd16996, 16'd43520, 16'd54815, 16'd54582, 16'd47687, 16'd38498, 16'd52500, 16'd58825, 16'd32809, 16'd12823, 16'd21958, 16'd58017, 16'd12037, 16'd62815, 16'd12123, 16'd32138, 16'd3667, 16'd18476, 16'd60833, 16'd4978, 16'd35949});
	test_expansion(128'ha46a540481cfba1f224f6322e2fd31b1, {16'd10984, 16'd59976, 16'd29386, 16'd50087, 16'd9038, 16'd25756, 16'd9701, 16'd20212, 16'd50331, 16'd12872, 16'd23283, 16'd18377, 16'd54103, 16'd45225, 16'd30818, 16'd5872, 16'd38033, 16'd21937, 16'd61428, 16'd18820, 16'd1751, 16'd49296, 16'd50482, 16'd5009, 16'd29797, 16'd32970});
	test_expansion(128'h58b3fa1f9247677502118f819c316190, {16'd49519, 16'd3977, 16'd19218, 16'd41799, 16'd26601, 16'd36554, 16'd22095, 16'd4479, 16'd2107, 16'd24941, 16'd47311, 16'd62034, 16'd37790, 16'd45218, 16'd23290, 16'd30711, 16'd17957, 16'd37682, 16'd44669, 16'd31472, 16'd116, 16'd63885, 16'd56707, 16'd31141, 16'd23919, 16'd8525});
	test_expansion(128'h3756928dcb632675166a8f669f66671d, {16'd14952, 16'd38108, 16'd62272, 16'd50329, 16'd61689, 16'd54226, 16'd6913, 16'd24416, 16'd62538, 16'd36180, 16'd31123, 16'd56740, 16'd44639, 16'd54298, 16'd3834, 16'd13577, 16'd45741, 16'd39101, 16'd37447, 16'd15033, 16'd12224, 16'd17566, 16'd40802, 16'd52049, 16'd7965, 16'd13677});
	test_expansion(128'h5f9fa36e50fe342005716bed5cb095ee, {16'd23713, 16'd50936, 16'd6871, 16'd47035, 16'd1175, 16'd19534, 16'd41119, 16'd29063, 16'd6330, 16'd28431, 16'd45461, 16'd15560, 16'd64489, 16'd29418, 16'd20255, 16'd26813, 16'd11057, 16'd5686, 16'd62729, 16'd17550, 16'd22823, 16'd6737, 16'd1193, 16'd42940, 16'd30204, 16'd52052});
	test_expansion(128'h8796faa4ce7bfc8a2a23de96054db717, {16'd45340, 16'd28852, 16'd57023, 16'd19496, 16'd49444, 16'd61797, 16'd27242, 16'd61429, 16'd23867, 16'd58669, 16'd49945, 16'd55952, 16'd28591, 16'd15255, 16'd45540, 16'd64827, 16'd13487, 16'd36126, 16'd59960, 16'd59682, 16'd1816, 16'd53767, 16'd6188, 16'd4597, 16'd29675, 16'd13716});
	test_expansion(128'h1bc3fea70f2ddfebf04af6a987d074a1, {16'd46506, 16'd63882, 16'd42620, 16'd4546, 16'd27060, 16'd62134, 16'd49910, 16'd27361, 16'd4665, 16'd43526, 16'd16415, 16'd51423, 16'd22431, 16'd63770, 16'd18790, 16'd39265, 16'd3998, 16'd48939, 16'd46116, 16'd51473, 16'd2264, 16'd38318, 16'd42933, 16'd38112, 16'd57021, 16'd59059});
	test_expansion(128'h6c7eeafdcc0dad7e235a14f4b586843e, {16'd23966, 16'd21191, 16'd43407, 16'd37595, 16'd41201, 16'd43760, 16'd14920, 16'd12231, 16'd10513, 16'd7549, 16'd41283, 16'd32815, 16'd50424, 16'd13237, 16'd55807, 16'd20015, 16'd47912, 16'd43365, 16'd22509, 16'd51256, 16'd25730, 16'd48694, 16'd1928, 16'd12843, 16'd450, 16'd49201});
	test_expansion(128'h3b35c44a52329cff9969940f3a38d507, {16'd9481, 16'd32831, 16'd54802, 16'd64283, 16'd28209, 16'd16969, 16'd19421, 16'd27349, 16'd30066, 16'd45183, 16'd6225, 16'd65289, 16'd38527, 16'd24057, 16'd16751, 16'd31286, 16'd62810, 16'd1055, 16'd22524, 16'd26301, 16'd22139, 16'd34128, 16'd49676, 16'd2623, 16'd5480, 16'd16438});
	test_expansion(128'hd989c66e0a36c23aa5fed756a8d3f039, {16'd47917, 16'd4572, 16'd34488, 16'd25874, 16'd9731, 16'd55280, 16'd61428, 16'd9798, 16'd61759, 16'd53056, 16'd6562, 16'd12655, 16'd16976, 16'd36790, 16'd37772, 16'd40447, 16'd58276, 16'd13909, 16'd62876, 16'd48674, 16'd33244, 16'd1085, 16'd25226, 16'd57021, 16'd27498, 16'd16987});
	test_expansion(128'h13c1b5eac0512ca493fe065cc228881a, {16'd61643, 16'd22700, 16'd32865, 16'd36198, 16'd57919, 16'd4943, 16'd48113, 16'd50674, 16'd15241, 16'd14526, 16'd62265, 16'd24814, 16'd49733, 16'd58768, 16'd12803, 16'd52524, 16'd28505, 16'd43498, 16'd44337, 16'd16714, 16'd57383, 16'd16188, 16'd45010, 16'd39900, 16'd62313, 16'd1171});
	test_expansion(128'h89d0124096d0aeaf5214dc9793777207, {16'd19701, 16'd35889, 16'd57616, 16'd8471, 16'd4131, 16'd62527, 16'd44324, 16'd6977, 16'd65398, 16'd9700, 16'd10840, 16'd3636, 16'd16196, 16'd48429, 16'd35296, 16'd31868, 16'd56360, 16'd29016, 16'd9485, 16'd33990, 16'd12366, 16'd64711, 16'd42979, 16'd59728, 16'd33349, 16'd45500});
	test_expansion(128'h48c1e99ac380bd9b915f820d88524a28, {16'd32291, 16'd23952, 16'd31408, 16'd59369, 16'd51284, 16'd29764, 16'd96, 16'd36310, 16'd19602, 16'd12197, 16'd27979, 16'd3249, 16'd65459, 16'd24627, 16'd45402, 16'd22797, 16'd7811, 16'd44676, 16'd15533, 16'd17198, 16'd33334, 16'd20059, 16'd54805, 16'd16923, 16'd6800, 16'd26333});
	test_expansion(128'h08566755cd9ad76f93a9a181ceceb070, {16'd43365, 16'd51911, 16'd50566, 16'd38896, 16'd30220, 16'd202, 16'd50519, 16'd19555, 16'd65226, 16'd52950, 16'd424, 16'd28879, 16'd39057, 16'd27677, 16'd20031, 16'd63457, 16'd36723, 16'd21462, 16'd5959, 16'd46565, 16'd36986, 16'd43758, 16'd58954, 16'd47786, 16'd54720, 16'd2702});
	test_expansion(128'h080fa6ce1f28dc7bbcf630637752a69f, {16'd14840, 16'd24062, 16'd31483, 16'd48263, 16'd39194, 16'd31062, 16'd39315, 16'd18586, 16'd12093, 16'd7787, 16'd41512, 16'd8412, 16'd47000, 16'd60911, 16'd13264, 16'd48140, 16'd42413, 16'd27895, 16'd64075, 16'd32097, 16'd15021, 16'd19834, 16'd15754, 16'd40831, 16'd60581, 16'd24302});
	test_expansion(128'h8da52e843268e6491b25a78c875ccde4, {16'd5410, 16'd49331, 16'd26063, 16'd6089, 16'd18397, 16'd2173, 16'd21896, 16'd5700, 16'd10540, 16'd65263, 16'd58942, 16'd13465, 16'd20872, 16'd3149, 16'd51009, 16'd1416, 16'd62757, 16'd44742, 16'd55960, 16'd25491, 16'd2787, 16'd20536, 16'd29718, 16'd12271, 16'd53870, 16'd38456});
	test_expansion(128'h2efd1108ac49584b32090002d7749882, {16'd44113, 16'd40345, 16'd33041, 16'd659, 16'd54379, 16'd18939, 16'd12106, 16'd55688, 16'd42101, 16'd6802, 16'd15431, 16'd23129, 16'd37334, 16'd33427, 16'd34442, 16'd16416, 16'd30844, 16'd58844, 16'd12583, 16'd27320, 16'd62673, 16'd60085, 16'd2201, 16'd47372, 16'd4448, 16'd16449});
	test_expansion(128'hc648a2b6d8a70be5271b86a4bc7d9aec, {16'd11031, 16'd46375, 16'd5186, 16'd35239, 16'd9663, 16'd53915, 16'd53481, 16'd14323, 16'd30554, 16'd46788, 16'd55796, 16'd4564, 16'd62275, 16'd21380, 16'd63462, 16'd61669, 16'd35956, 16'd27282, 16'd24327, 16'd73, 16'd40450, 16'd33239, 16'd26084, 16'd36556, 16'd8909, 16'd2705});
	test_expansion(128'h77c9662166db82637b2dd23631ad38c2, {16'd57180, 16'd11273, 16'd43954, 16'd4670, 16'd35154, 16'd37765, 16'd12621, 16'd11912, 16'd49235, 16'd9280, 16'd51455, 16'd47833, 16'd11199, 16'd22695, 16'd53133, 16'd55895, 16'd11180, 16'd27108, 16'd64170, 16'd37738, 16'd23497, 16'd2081, 16'd27153, 16'd15110, 16'd23966, 16'd55166});
	test_expansion(128'he9388b5003bca82235dcd196b514dfd3, {16'd61675, 16'd30871, 16'd10527, 16'd24566, 16'd48659, 16'd45486, 16'd40386, 16'd51496, 16'd40569, 16'd53685, 16'd34986, 16'd3583, 16'd10326, 16'd645, 16'd20456, 16'd29149, 16'd14552, 16'd13909, 16'd28461, 16'd34564, 16'd14273, 16'd44492, 16'd58162, 16'd36013, 16'd38861, 16'd14193});
	test_expansion(128'h1f14807e014f5eb466b9aab2af5f7678, {16'd23183, 16'd47080, 16'd30948, 16'd14682, 16'd47709, 16'd64866, 16'd49804, 16'd6776, 16'd47449, 16'd16529, 16'd19381, 16'd36094, 16'd19650, 16'd26075, 16'd58622, 16'd14928, 16'd17501, 16'd39010, 16'd48619, 16'd19341, 16'd46852, 16'd40570, 16'd63465, 16'd5393, 16'd55230, 16'd35489});
	test_expansion(128'h699caac0c61e6c864950bcaf4ede5923, {16'd10453, 16'd29029, 16'd25950, 16'd18706, 16'd47017, 16'd33917, 16'd29201, 16'd57663, 16'd62674, 16'd22998, 16'd36440, 16'd15495, 16'd49400, 16'd41837, 16'd65137, 16'd49757, 16'd32244, 16'd41123, 16'd22685, 16'd12546, 16'd21586, 16'd43435, 16'd35675, 16'd47383, 16'd51962, 16'd44199});
	test_expansion(128'hc194130202c70f1f530053741f16539e, {16'd27977, 16'd2454, 16'd21688, 16'd53348, 16'd5337, 16'd11201, 16'd27501, 16'd46051, 16'd17048, 16'd7172, 16'd57032, 16'd51580, 16'd52958, 16'd38096, 16'd45139, 16'd35607, 16'd46532, 16'd30026, 16'd41241, 16'd18617, 16'd52012, 16'd15338, 16'd7302, 16'd52243, 16'd25263, 16'd53710});
	test_expansion(128'h72318e272688ce65a3260e4fef28e1b0, {16'd62066, 16'd30023, 16'd26241, 16'd25158, 16'd45931, 16'd22036, 16'd28547, 16'd336, 16'd28845, 16'd43948, 16'd33816, 16'd34226, 16'd35039, 16'd22978, 16'd42323, 16'd29811, 16'd461, 16'd23990, 16'd60329, 16'd28736, 16'd56217, 16'd53125, 16'd16699, 16'd29883, 16'd63816, 16'd52665});
	test_expansion(128'h338ecc75710f1e825d777ae2b0a7a4fe, {16'd29745, 16'd1292, 16'd14398, 16'd43500, 16'd42618, 16'd48190, 16'd48558, 16'd51203, 16'd6295, 16'd43090, 16'd44610, 16'd6064, 16'd42581, 16'd2272, 16'd41090, 16'd48121, 16'd65055, 16'd64327, 16'd55152, 16'd7298, 16'd35448, 16'd28340, 16'd53934, 16'd15094, 16'd43447, 16'd12013});
	test_expansion(128'hea1d33d0e4ef43b340835b26df8d1327, {16'd61665, 16'd58695, 16'd50449, 16'd1827, 16'd42675, 16'd2735, 16'd418, 16'd9013, 16'd9573, 16'd19429, 16'd51423, 16'd55377, 16'd38420, 16'd24449, 16'd1379, 16'd15945, 16'd13320, 16'd39030, 16'd54650, 16'd19015, 16'd13325, 16'd14744, 16'd64647, 16'd19224, 16'd60716, 16'd53418});
	test_expansion(128'h15a88d311562b4200abd038f3a291331, {16'd33930, 16'd55394, 16'd44101, 16'd39702, 16'd1689, 16'd47476, 16'd59720, 16'd39518, 16'd23479, 16'd256, 16'd40043, 16'd6771, 16'd9448, 16'd19259, 16'd2201, 16'd44990, 16'd28341, 16'd33605, 16'd50154, 16'd27649, 16'd17734, 16'd10636, 16'd60866, 16'd63864, 16'd6908, 16'd12918});
	test_expansion(128'h0bfa8abc135954920734583470538f9a, {16'd53502, 16'd53531, 16'd45841, 16'd19000, 16'd57673, 16'd16418, 16'd24461, 16'd3458, 16'd49895, 16'd39187, 16'd51642, 16'd43520, 16'd21362, 16'd36896, 16'd55219, 16'd43870, 16'd12241, 16'd10779, 16'd50497, 16'd35830, 16'd16613, 16'd49647, 16'd64108, 16'd4694, 16'd27054, 16'd405});
	test_expansion(128'h40178842b3dea0ef74421690077d463c, {16'd33476, 16'd50886, 16'd20168, 16'd19748, 16'd8098, 16'd54518, 16'd41395, 16'd63142, 16'd63083, 16'd9306, 16'd60254, 16'd5868, 16'd54446, 16'd50024, 16'd49645, 16'd33059, 16'd30254, 16'd42162, 16'd11950, 16'd23824, 16'd39610, 16'd30296, 16'd37658, 16'd892, 16'd50219, 16'd7022});
	test_expansion(128'h74040ac65339863e516b82e8ee3a3ced, {16'd33977, 16'd30121, 16'd63018, 16'd8073, 16'd25688, 16'd43579, 16'd41286, 16'd5760, 16'd41904, 16'd54308, 16'd46452, 16'd57087, 16'd54243, 16'd31753, 16'd18468, 16'd33162, 16'd36155, 16'd59022, 16'd22579, 16'd19844, 16'd63249, 16'd17610, 16'd45964, 16'd42341, 16'd21183, 16'd62357});
	test_expansion(128'h6279e8839404f4d4bf4dc0df39037568, {16'd41271, 16'd3015, 16'd8674, 16'd40252, 16'd62940, 16'd34853, 16'd15314, 16'd7884, 16'd33478, 16'd20427, 16'd61739, 16'd50505, 16'd50156, 16'd22618, 16'd40321, 16'd1369, 16'd18314, 16'd39776, 16'd11465, 16'd6219, 16'd23942, 16'd2089, 16'd15920, 16'd43957, 16'd18568, 16'd1266});
	test_expansion(128'h86c141efd76277291d329a5a371b1be2, {16'd56768, 16'd54594, 16'd19909, 16'd49926, 16'd63742, 16'd58483, 16'd18952, 16'd13036, 16'd9431, 16'd64721, 16'd59092, 16'd10547, 16'd12798, 16'd14659, 16'd14394, 16'd7877, 16'd32369, 16'd10458, 16'd21347, 16'd30754, 16'd31323, 16'd52362, 16'd41572, 16'd35953, 16'd3785, 16'd23711});
	test_expansion(128'hffc8ae5550ac7067ec403a12cb1e1cc9, {16'd30950, 16'd12562, 16'd28563, 16'd27509, 16'd10869, 16'd46862, 16'd25509, 16'd26105, 16'd22443, 16'd42271, 16'd65399, 16'd51851, 16'd5114, 16'd23233, 16'd4894, 16'd63415, 16'd51447, 16'd51887, 16'd22713, 16'd26792, 16'd50620, 16'd1104, 16'd11548, 16'd24059, 16'd11995, 16'd866});
	test_expansion(128'h7ac4db20375a9ea3d09ec5ec652c454e, {16'd11433, 16'd7987, 16'd54073, 16'd50641, 16'd4043, 16'd52350, 16'd13246, 16'd31221, 16'd25529, 16'd54437, 16'd50604, 16'd38917, 16'd63973, 16'd50612, 16'd45774, 16'd4140, 16'd34399, 16'd6789, 16'd44572, 16'd5343, 16'd30894, 16'd2257, 16'd44857, 16'd15943, 16'd40140, 16'd43284});
	test_expansion(128'h13aca48337d3eec2da59a33765bdc2e4, {16'd54684, 16'd40411, 16'd6737, 16'd51651, 16'd11493, 16'd36585, 16'd2047, 16'd9295, 16'd11349, 16'd6535, 16'd43289, 16'd39116, 16'd20108, 16'd4004, 16'd14430, 16'd16451, 16'd13449, 16'd3309, 16'd32197, 16'd4068, 16'd24549, 16'd10975, 16'd16742, 16'd8286, 16'd44084, 16'd9848});
	test_expansion(128'h8ed5420570bbba9d398f42aa0069f283, {16'd42990, 16'd60859, 16'd19142, 16'd36821, 16'd29861, 16'd28644, 16'd11941, 16'd8985, 16'd48447, 16'd63633, 16'd17183, 16'd35088, 16'd15685, 16'd52928, 16'd30633, 16'd7527, 16'd13350, 16'd36311, 16'd1802, 16'd22211, 16'd55662, 16'd15513, 16'd14840, 16'd27098, 16'd61327, 16'd28644});
	test_expansion(128'hcaabe40d54b27758fc5262c2cff1293e, {16'd45489, 16'd17260, 16'd13025, 16'd6459, 16'd61168, 16'd23930, 16'd15154, 16'd4379, 16'd37041, 16'd15003, 16'd7168, 16'd62807, 16'd41140, 16'd58832, 16'd34977, 16'd27689, 16'd18065, 16'd42844, 16'd45554, 16'd55552, 16'd2805, 16'd46234, 16'd30771, 16'd41009, 16'd7311, 16'd27085});
	test_expansion(128'h30f716b58843e52e362881bba1bcba87, {16'd15401, 16'd26311, 16'd55839, 16'd4354, 16'd56008, 16'd36030, 16'd54313, 16'd63654, 16'd18489, 16'd9327, 16'd50050, 16'd59268, 16'd43579, 16'd32744, 16'd54973, 16'd21664, 16'd57860, 16'd65430, 16'd36073, 16'd2505, 16'd41647, 16'd56273, 16'd3327, 16'd2109, 16'd52761, 16'd7693});
	test_expansion(128'h04d506ea6523231632992a5920bca074, {16'd2287, 16'd18722, 16'd16849, 16'd54103, 16'd14358, 16'd38078, 16'd10662, 16'd63148, 16'd44091, 16'd46813, 16'd41624, 16'd47710, 16'd5304, 16'd64229, 16'd22202, 16'd47481, 16'd20367, 16'd41877, 16'd28145, 16'd23875, 16'd10567, 16'd23984, 16'd31449, 16'd34151, 16'd60498, 16'd37983});
	test_expansion(128'h9f5dccde532d8e41a01b0a53fd1b19c5, {16'd27154, 16'd28540, 16'd33275, 16'd33369, 16'd29401, 16'd4999, 16'd54392, 16'd25558, 16'd61241, 16'd17501, 16'd20034, 16'd32556, 16'd4584, 16'd4616, 16'd46823, 16'd47014, 16'd20869, 16'd6048, 16'd28302, 16'd43122, 16'd26981, 16'd18762, 16'd28317, 16'd28252, 16'd14569, 16'd6696});
	test_expansion(128'h8a24778a2c5d5916eab45527079b676f, {16'd22982, 16'd14106, 16'd51342, 16'd7288, 16'd25193, 16'd45318, 16'd54985, 16'd58621, 16'd62688, 16'd57723, 16'd37436, 16'd40746, 16'd13140, 16'd47369, 16'd30899, 16'd2661, 16'd41892, 16'd53013, 16'd47608, 16'd46460, 16'd11277, 16'd63770, 16'd59386, 16'd18089, 16'd1319, 16'd7314});
	test_expansion(128'hb7a7d034e3ebe21e6974ae10233453ff, {16'd37694, 16'd17195, 16'd13223, 16'd12680, 16'd58616, 16'd5220, 16'd14011, 16'd64843, 16'd58294, 16'd39165, 16'd52211, 16'd13383, 16'd19238, 16'd5275, 16'd52796, 16'd43374, 16'd24402, 16'd32013, 16'd25435, 16'd18840, 16'd49803, 16'd21011, 16'd18303, 16'd64902, 16'd57132, 16'd40719});
	test_expansion(128'h33d895a96d4a59cb5cfe5a691ff081f8, {16'd21116, 16'd58400, 16'd27858, 16'd11725, 16'd54117, 16'd24699, 16'd40805, 16'd24568, 16'd38676, 16'd22493, 16'd29101, 16'd11604, 16'd57983, 16'd43198, 16'd26526, 16'd60395, 16'd30230, 16'd55904, 16'd34745, 16'd22945, 16'd23886, 16'd18581, 16'd19229, 16'd63594, 16'd1951, 16'd12947});
	test_expansion(128'hc3f43553a7efa1265ba49be549e582d5, {16'd4116, 16'd18615, 16'd30059, 16'd34450, 16'd47948, 16'd36950, 16'd64641, 16'd52002, 16'd5930, 16'd36375, 16'd17030, 16'd2573, 16'd2224, 16'd27934, 16'd42383, 16'd11855, 16'd53235, 16'd28465, 16'd5804, 16'd8600, 16'd43120, 16'd36410, 16'd1974, 16'd40289, 16'd12498, 16'd8722});
	test_expansion(128'hf03a968200b183eb71ac9719e6039563, {16'd45705, 16'd20704, 16'd31147, 16'd54994, 16'd21148, 16'd21763, 16'd15322, 16'd26744, 16'd20365, 16'd53678, 16'd17018, 16'd770, 16'd59554, 16'd25686, 16'd54632, 16'd1043, 16'd50651, 16'd45075, 16'd40925, 16'd25496, 16'd44529, 16'd49297, 16'd53348, 16'd49006, 16'd25985, 16'd29});
	test_expansion(128'h2c2ca45331773081882af07fc34eb9fd, {16'd51557, 16'd16385, 16'd5789, 16'd4692, 16'd63884, 16'd8656, 16'd925, 16'd32366, 16'd33787, 16'd20501, 16'd31487, 16'd7786, 16'd33195, 16'd17237, 16'd9921, 16'd62150, 16'd24560, 16'd10608, 16'd11115, 16'd1778, 16'd24660, 16'd53880, 16'd9220, 16'd865, 16'd55055, 16'd58002});
	test_expansion(128'hf97c4b2b77067ff3896448d6b18a33dd, {16'd23767, 16'd64607, 16'd55594, 16'd29477, 16'd16329, 16'd65429, 16'd21180, 16'd42296, 16'd3550, 16'd4744, 16'd56671, 16'd21916, 16'd22024, 16'd22113, 16'd21349, 16'd51684, 16'd60195, 16'd5691, 16'd18, 16'd12425, 16'd9403, 16'd37171, 16'd52866, 16'd16888, 16'd5531, 16'd64855});
	test_expansion(128'hbc9663d87d0cc08cde5360ccd221fb77, {16'd35421, 16'd4320, 16'd14197, 16'd11024, 16'd19679, 16'd21415, 16'd27789, 16'd53549, 16'd37101, 16'd10043, 16'd44061, 16'd44097, 16'd37942, 16'd41434, 16'd51823, 16'd52725, 16'd5263, 16'd50483, 16'd10925, 16'd11371, 16'd64755, 16'd36428, 16'd27144, 16'd34344, 16'd27537, 16'd30039});
	test_expansion(128'h3f288085087b856331d44d641ca4ded3, {16'd39246, 16'd3518, 16'd51908, 16'd13673, 16'd27628, 16'd25464, 16'd1339, 16'd61412, 16'd64303, 16'd8976, 16'd23650, 16'd34093, 16'd40001, 16'd10137, 16'd21471, 16'd51193, 16'd51361, 16'd23572, 16'd38047, 16'd53658, 16'd24645, 16'd40021, 16'd57029, 16'd59155, 16'd47106, 16'd1831});
	test_expansion(128'h4674f713119c232b723da66bb63df94e, {16'd50755, 16'd6703, 16'd20497, 16'd29859, 16'd32030, 16'd9080, 16'd36978, 16'd57964, 16'd38734, 16'd27835, 16'd47176, 16'd42975, 16'd20335, 16'd3114, 16'd32037, 16'd58608, 16'd15252, 16'd14557, 16'd23558, 16'd41201, 16'd56614, 16'd7877, 16'd17041, 16'd14852, 16'd29189, 16'd23858});
	test_expansion(128'h4dd328a9b3a807b8e4737c0d43a1a676, {16'd6209, 16'd12743, 16'd21109, 16'd29385, 16'd17921, 16'd58584, 16'd63050, 16'd19444, 16'd24383, 16'd17920, 16'd24805, 16'd6790, 16'd28490, 16'd4352, 16'd58320, 16'd25613, 16'd49165, 16'd26072, 16'd10136, 16'd57469, 16'd52940, 16'd45441, 16'd32730, 16'd41738, 16'd29023, 16'd8178});
	test_expansion(128'h8698f43dfd3c608d67b5d07aab020df2, {16'd16979, 16'd11226, 16'd41390, 16'd32474, 16'd50172, 16'd1265, 16'd58811, 16'd39445, 16'd58181, 16'd61162, 16'd31062, 16'd39973, 16'd21550, 16'd64283, 16'd52882, 16'd55717, 16'd40639, 16'd56467, 16'd29048, 16'd17760, 16'd3558, 16'd24824, 16'd14394, 16'd8253, 16'd54184, 16'd31635});
	test_expansion(128'h0a217ebcf70fa81e91db8b6add2bc444, {16'd44785, 16'd63743, 16'd28864, 16'd5262, 16'd20886, 16'd35416, 16'd2597, 16'd23520, 16'd25985, 16'd1820, 16'd63392, 16'd18249, 16'd9123, 16'd51531, 16'd56662, 16'd8273, 16'd52451, 16'd60613, 16'd42998, 16'd39097, 16'd52951, 16'd929, 16'd16070, 16'd3860, 16'd4945, 16'd62770});
	test_expansion(128'h927e982b373dd5eca51191e2a7fe575e, {16'd62108, 16'd19539, 16'd5388, 16'd15168, 16'd22546, 16'd63831, 16'd27887, 16'd24011, 16'd51067, 16'd59005, 16'd14807, 16'd61817, 16'd27413, 16'd9333, 16'd61304, 16'd34210, 16'd22016, 16'd16518, 16'd30008, 16'd4986, 16'd3311, 16'd19346, 16'd34578, 16'd46065, 16'd60341, 16'd11972});
	test_expansion(128'h4d4d6eabfb1244f3d0859d74a6d931dc, {16'd13371, 16'd8100, 16'd16491, 16'd20134, 16'd48521, 16'd42691, 16'd4715, 16'd51102, 16'd31163, 16'd1648, 16'd56639, 16'd49685, 16'd12594, 16'd18599, 16'd43148, 16'd64043, 16'd277, 16'd51397, 16'd38223, 16'd59290, 16'd39775, 16'd11786, 16'd36367, 16'd61536, 16'd22761, 16'd60386});
	test_expansion(128'he5e76323d1a0113a2e3bb5b09ea80bd4, {16'd33932, 16'd38758, 16'd59936, 16'd50375, 16'd39895, 16'd22023, 16'd18110, 16'd41537, 16'd49103, 16'd44417, 16'd22768, 16'd33791, 16'd48027, 16'd47158, 16'd37726, 16'd12926, 16'd39143, 16'd8794, 16'd12303, 16'd64869, 16'd64536, 16'd10383, 16'd52558, 16'd26551, 16'd3450, 16'd35450});
	test_expansion(128'h419d798ba4d74b187ebec82fc57dd852, {16'd21291, 16'd19915, 16'd20216, 16'd30035, 16'd13798, 16'd16406, 16'd1478, 16'd5170, 16'd56403, 16'd59783, 16'd59600, 16'd8779, 16'd61067, 16'd11028, 16'd32955, 16'd57449, 16'd15626, 16'd45908, 16'd54041, 16'd57587, 16'd53681, 16'd16060, 16'd27319, 16'd35431, 16'd12583, 16'd41174});
	test_expansion(128'h976f3f3f1825b701069df899c797bdb6, {16'd31433, 16'd36028, 16'd38243, 16'd13788, 16'd55235, 16'd48998, 16'd44298, 16'd7518, 16'd27881, 16'd60009, 16'd9673, 16'd42406, 16'd11465, 16'd37087, 16'd28627, 16'd51781, 16'd52979, 16'd3085, 16'd30089, 16'd39142, 16'd27908, 16'd4362, 16'd18458, 16'd48888, 16'd5265, 16'd57603});
	test_expansion(128'ha841780df8a2d70d9a931a5da5f10f0f, {16'd43940, 16'd59214, 16'd45844, 16'd31274, 16'd41457, 16'd59640, 16'd30763, 16'd58738, 16'd9771, 16'd9282, 16'd64954, 16'd24465, 16'd9477, 16'd8038, 16'd44584, 16'd19286, 16'd44615, 16'd65100, 16'd29113, 16'd64401, 16'd49999, 16'd9167, 16'd47022, 16'd34409, 16'd2325, 16'd20901});
	test_expansion(128'h5899bb72d8d834c3eee8e3ccba940c1c, {16'd35261, 16'd35963, 16'd2114, 16'd10151, 16'd65496, 16'd53867, 16'd59749, 16'd7431, 16'd16406, 16'd61908, 16'd32904, 16'd45660, 16'd9525, 16'd18631, 16'd35928, 16'd52636, 16'd58120, 16'd39758, 16'd34978, 16'd58255, 16'd30842, 16'd37790, 16'd59177, 16'd1628, 16'd61734, 16'd27274});
	test_expansion(128'h385ac947c436950aa68356db7e8b7d37, {16'd58322, 16'd47155, 16'd58714, 16'd35154, 16'd32864, 16'd39449, 16'd25924, 16'd15054, 16'd32250, 16'd45060, 16'd27598, 16'd16348, 16'd46718, 16'd43149, 16'd32683, 16'd25225, 16'd38539, 16'd14928, 16'd2286, 16'd61179, 16'd27658, 16'd25315, 16'd29050, 16'd8876, 16'd44976, 16'd13226});
	test_expansion(128'h413d41d2c1744a783997df52308d248b, {16'd13064, 16'd18397, 16'd13019, 16'd28211, 16'd54692, 16'd31071, 16'd34326, 16'd37559, 16'd27236, 16'd18860, 16'd36069, 16'd59135, 16'd543, 16'd60055, 16'd17778, 16'd56943, 16'd54426, 16'd63262, 16'd5275, 16'd1485, 16'd16648, 16'd22713, 16'd26845, 16'd56615, 16'd6270, 16'd33728});
	test_expansion(128'hc33fc6fd5c94ed118ed443802b0f8c45, {16'd9056, 16'd12958, 16'd12375, 16'd908, 16'd11685, 16'd54796, 16'd14619, 16'd53051, 16'd44514, 16'd21828, 16'd60435, 16'd15096, 16'd1025, 16'd18205, 16'd15962, 16'd7914, 16'd59417, 16'd29543, 16'd25851, 16'd41533, 16'd26069, 16'd57040, 16'd1176, 16'd50220, 16'd27753, 16'd64690});
	test_expansion(128'h99a7ce47f789916e1117102b2ca2d472, {16'd18447, 16'd29317, 16'd53941, 16'd63060, 16'd12770, 16'd62887, 16'd50809, 16'd55188, 16'd28390, 16'd42086, 16'd11293, 16'd22125, 16'd41144, 16'd4815, 16'd50463, 16'd45522, 16'd37931, 16'd20766, 16'd30445, 16'd22922, 16'd55624, 16'd25425, 16'd50219, 16'd62672, 16'd19732, 16'd50591});
	test_expansion(128'h4bcbffb73ea7f474d674fb1bfb314272, {16'd59153, 16'd28395, 16'd51320, 16'd58714, 16'd33465, 16'd23266, 16'd36565, 16'd7901, 16'd11179, 16'd34288, 16'd635, 16'd64006, 16'd44199, 16'd32990, 16'd64213, 16'd55591, 16'd53916, 16'd28610, 16'd1204, 16'd844, 16'd24473, 16'd15208, 16'd63460, 16'd22547, 16'd10629, 16'd26782});
	test_expansion(128'h285e77303da5de2a112b0e5e06aca887, {16'd33138, 16'd54384, 16'd19735, 16'd64000, 16'd16826, 16'd32300, 16'd31010, 16'd13940, 16'd42497, 16'd30264, 16'd53852, 16'd9409, 16'd43933, 16'd35085, 16'd7834, 16'd46454, 16'd43571, 16'd32372, 16'd51600, 16'd18210, 16'd64225, 16'd54056, 16'd14255, 16'd34517, 16'd55611, 16'd55269});
	test_expansion(128'h4fcdc4ce2c703e9f434aa923464edd2d, {16'd1544, 16'd59702, 16'd47385, 16'd31887, 16'd27643, 16'd33226, 16'd11211, 16'd28732, 16'd43057, 16'd35337, 16'd8316, 16'd5155, 16'd58667, 16'd35215, 16'd56484, 16'd47581, 16'd3260, 16'd24442, 16'd4931, 16'd35702, 16'd26835, 16'd4714, 16'd42416, 16'd35473, 16'd924, 16'd53397});
	test_expansion(128'h0a0aaf2359ef43aaa2a5b10c37642bb5, {16'd11452, 16'd49870, 16'd49962, 16'd30779, 16'd24176, 16'd27582, 16'd65401, 16'd13315, 16'd62671, 16'd5494, 16'd38280, 16'd27436, 16'd55002, 16'd25585, 16'd45039, 16'd10115, 16'd23199, 16'd37351, 16'd47541, 16'd32505, 16'd21139, 16'd41596, 16'd29063, 16'd7885, 16'd32764, 16'd5671});
	test_expansion(128'h5a7ade906990fb67ab0fb8a2da5f2d42, {16'd62285, 16'd6170, 16'd9820, 16'd20156, 16'd49182, 16'd55530, 16'd9622, 16'd2897, 16'd33048, 16'd10018, 16'd59044, 16'd60013, 16'd7090, 16'd20964, 16'd39651, 16'd6194, 16'd64287, 16'd13631, 16'd6318, 16'd54953, 16'd59291, 16'd46375, 16'd37613, 16'd57314, 16'd32659, 16'd17555});
	test_expansion(128'h68eeab0b5a7e0898b1c2a1eb14f577c4, {16'd55469, 16'd46220, 16'd1993, 16'd47629, 16'd7920, 16'd65462, 16'd512, 16'd4712, 16'd12417, 16'd3976, 16'd9666, 16'd26977, 16'd47923, 16'd20162, 16'd62798, 16'd21670, 16'd29741, 16'd65502, 16'd38093, 16'd64555, 16'd34330, 16'd54802, 16'd19031, 16'd61512, 16'd18400, 16'd52564});
	test_expansion(128'h4b533bd705b6fc040fa0b6440dfa6739, {16'd62877, 16'd50072, 16'd32604, 16'd30171, 16'd54204, 16'd590, 16'd46260, 16'd55531, 16'd51781, 16'd28927, 16'd10668, 16'd49223, 16'd32120, 16'd39711, 16'd41904, 16'd33575, 16'd17817, 16'd57254, 16'd5932, 16'd13533, 16'd25497, 16'd15296, 16'd58409, 16'd17385, 16'd34640, 16'd7841});
	test_expansion(128'ha327fb069be6e60b19c08b3b19bdd2e1, {16'd53395, 16'd47980, 16'd8799, 16'd33803, 16'd5407, 16'd18657, 16'd12107, 16'd48482, 16'd4705, 16'd23005, 16'd24136, 16'd16621, 16'd12868, 16'd1737, 16'd37255, 16'd6272, 16'd46145, 16'd22482, 16'd25881, 16'd4749, 16'd732, 16'd63162, 16'd34804, 16'd54665, 16'd41344, 16'd14871});
	test_expansion(128'ha103a4a77386a71472a3540b54d182ae, {16'd7120, 16'd51722, 16'd42908, 16'd65014, 16'd8141, 16'd12308, 16'd20253, 16'd50745, 16'd60959, 16'd21332, 16'd28415, 16'd55085, 16'd11564, 16'd26482, 16'd41836, 16'd7436, 16'd41314, 16'd30512, 16'd3062, 16'd63736, 16'd36346, 16'd52731, 16'd53786, 16'd4350, 16'd63412, 16'd1322});
	test_expansion(128'h150305f68bed0ba348f96382356ccc55, {16'd38415, 16'd26117, 16'd59401, 16'd61057, 16'd39841, 16'd55438, 16'd63937, 16'd48348, 16'd26085, 16'd59523, 16'd25624, 16'd6066, 16'd9814, 16'd53130, 16'd60164, 16'd51032, 16'd24664, 16'd30699, 16'd64664, 16'd21794, 16'd16411, 16'd56560, 16'd45841, 16'd35651, 16'd57880, 16'd37724});
	test_expansion(128'ha80086db4dc0faa74da1f907dfe7589f, {16'd31442, 16'd32023, 16'd14906, 16'd24479, 16'd42171, 16'd25434, 16'd34252, 16'd56362, 16'd49034, 16'd46222, 16'd63398, 16'd57600, 16'd18584, 16'd65270, 16'd45791, 16'd7417, 16'd16428, 16'd2392, 16'd4705, 16'd55478, 16'd7577, 16'd20195, 16'd20007, 16'd31392, 16'd58696, 16'd18629});
	test_expansion(128'h6cf965e782af66a383e283c85f1b4725, {16'd60525, 16'd6133, 16'd60771, 16'd46861, 16'd32923, 16'd62001, 16'd44513, 16'd25578, 16'd45469, 16'd28154, 16'd34263, 16'd31501, 16'd19256, 16'd4524, 16'd28666, 16'd15674, 16'd58816, 16'd10059, 16'd22362, 16'd15704, 16'd48397, 16'd27870, 16'd64599, 16'd37102, 16'd35955, 16'd25027});
	test_expansion(128'h8ed1e15f5713931ba57f0f62375bc97d, {16'd5402, 16'd56456, 16'd20846, 16'd41379, 16'd22002, 16'd24713, 16'd35217, 16'd21465, 16'd4200, 16'd59455, 16'd17016, 16'd10947, 16'd6790, 16'd16486, 16'd38335, 16'd61361, 16'd31680, 16'd2737, 16'd18160, 16'd60079, 16'd27145, 16'd41676, 16'd21729, 16'd61329, 16'd63386, 16'd50785});
	test_expansion(128'h188e38d4738809a08a60816b01e7eb73, {16'd65113, 16'd45362, 16'd38575, 16'd20461, 16'd19019, 16'd48563, 16'd64676, 16'd46125, 16'd4338, 16'd18835, 16'd49058, 16'd36210, 16'd32928, 16'd19872, 16'd30899, 16'd26359, 16'd5820, 16'd15839, 16'd53279, 16'd65032, 16'd38995, 16'd54122, 16'd18834, 16'd46516, 16'd14566, 16'd56027});
	test_expansion(128'h3d5f922f5ae8257211383f5de8ab5014, {16'd63132, 16'd11363, 16'd48058, 16'd64377, 16'd26114, 16'd64309, 16'd39406, 16'd29139, 16'd21750, 16'd56039, 16'd50485, 16'd26280, 16'd10390, 16'd7468, 16'd16869, 16'd5547, 16'd4648, 16'd41770, 16'd37224, 16'd10511, 16'd25842, 16'd60435, 16'd8975, 16'd22484, 16'd30113, 16'd58673});
	test_expansion(128'ha9e387c8d850631feb5d64ce5d41aa0c, {16'd33809, 16'd48275, 16'd10022, 16'd40798, 16'd28128, 16'd27045, 16'd5895, 16'd62866, 16'd38048, 16'd38282, 16'd64363, 16'd19732, 16'd50356, 16'd63256, 16'd48074, 16'd7577, 16'd2886, 16'd64678, 16'd45567, 16'd34062, 16'd23445, 16'd37189, 16'd913, 16'd54012, 16'd17368, 16'd48483});
	test_expansion(128'h76b4f7b291c29bd865a9bc88acd9ccc4, {16'd56099, 16'd5629, 16'd43355, 16'd45248, 16'd12669, 16'd60827, 16'd17452, 16'd34657, 16'd54548, 16'd28856, 16'd46032, 16'd14988, 16'd13322, 16'd52171, 16'd25441, 16'd57547, 16'd41876, 16'd19973, 16'd10375, 16'd41613, 16'd9628, 16'd17393, 16'd32876, 16'd35252, 16'd7354, 16'd59031});
	test_expansion(128'h9452d5dc208ce95d8720f8469dbb7797, {16'd5585, 16'd5287, 16'd13514, 16'd18967, 16'd49611, 16'd38589, 16'd40936, 16'd57015, 16'd42318, 16'd48495, 16'd55324, 16'd40584, 16'd416, 16'd29992, 16'd15281, 16'd18598, 16'd53760, 16'd15867, 16'd36286, 16'd16812, 16'd27171, 16'd42940, 16'd4186, 16'd22014, 16'd37547, 16'd19120});
	test_expansion(128'h9129b89ecd2097b305a35645550bac85, {16'd59083, 16'd49278, 16'd20240, 16'd52057, 16'd42902, 16'd36135, 16'd473, 16'd25653, 16'd18212, 16'd47180, 16'd45686, 16'd57654, 16'd38823, 16'd57003, 16'd59296, 16'd50002, 16'd17805, 16'd64413, 16'd49477, 16'd41548, 16'd60530, 16'd11412, 16'd19257, 16'd36877, 16'd51112, 16'd45467});
	test_expansion(128'hfdcdc91e0e8e3ff12c3885b0b9950f54, {16'd54482, 16'd47198, 16'd50287, 16'd56666, 16'd12670, 16'd39944, 16'd27321, 16'd31822, 16'd63557, 16'd825, 16'd20384, 16'd59805, 16'd15952, 16'd51607, 16'd6537, 16'd60628, 16'd46291, 16'd36355, 16'd9707, 16'd31283, 16'd15771, 16'd59781, 16'd17047, 16'd36787, 16'd40928, 16'd4615});
	test_expansion(128'h72fdcd336fa3041c8a95751e072b213d, {16'd24959, 16'd59445, 16'd13104, 16'd28268, 16'd60315, 16'd4949, 16'd16826, 16'd20511, 16'd65029, 16'd44041, 16'd5821, 16'd52519, 16'd33805, 16'd8697, 16'd46704, 16'd63027, 16'd48512, 16'd11302, 16'd36493, 16'd16099, 16'd46481, 16'd9175, 16'd9971, 16'd63605, 16'd62972, 16'd27879});
	test_expansion(128'hf2e9e78963aee96953bbbaf597044ec7, {16'd15007, 16'd9913, 16'd35267, 16'd18918, 16'd7850, 16'd19536, 16'd57234, 16'd41756, 16'd34919, 16'd12381, 16'd35296, 16'd26043, 16'd7344, 16'd56786, 16'd35701, 16'd650, 16'd41049, 16'd47949, 16'd19168, 16'd19593, 16'd33362, 16'd24086, 16'd49831, 16'd61759, 16'd6815, 16'd19651});
	test_expansion(128'hd20c758c5dda77b198d7157d619b3942, {16'd15690, 16'd61519, 16'd45082, 16'd33054, 16'd64585, 16'd23623, 16'd62242, 16'd4676, 16'd56632, 16'd28032, 16'd14983, 16'd56571, 16'd62480, 16'd23984, 16'd62533, 16'd62614, 16'd63199, 16'd23454, 16'd18892, 16'd2863, 16'd37743, 16'd12300, 16'd11893, 16'd10963, 16'd61528, 16'd53514});
	test_expansion(128'h18558271fc146403964ddd688e3d3d5b, {16'd48968, 16'd16604, 16'd47951, 16'd1291, 16'd55189, 16'd19396, 16'd14866, 16'd63299, 16'd51198, 16'd27546, 16'd42919, 16'd1860, 16'd6120, 16'd4101, 16'd38139, 16'd60330, 16'd59450, 16'd49898, 16'd34839, 16'd54360, 16'd12863, 16'd58089, 16'd56431, 16'd30925, 16'd49109, 16'd34480});
	test_expansion(128'h7d5560f9f8d054658db881bef5cd9dec, {16'd50232, 16'd51314, 16'd58899, 16'd25773, 16'd22821, 16'd44301, 16'd40262, 16'd64548, 16'd19584, 16'd18625, 16'd32868, 16'd873, 16'd23608, 16'd33900, 16'd32549, 16'd38979, 16'd29866, 16'd29082, 16'd34080, 16'd20535, 16'd27370, 16'd56929, 16'd10875, 16'd48124, 16'd31241, 16'd16202});
	test_expansion(128'h8b28a1261493c553ef60e5935ddbbe05, {16'd61160, 16'd52561, 16'd12089, 16'd43611, 16'd63051, 16'd48676, 16'd50119, 16'd5778, 16'd40649, 16'd979, 16'd17506, 16'd15485, 16'd28469, 16'd36299, 16'd46520, 16'd40885, 16'd14984, 16'd12624, 16'd43087, 16'd20659, 16'd29301, 16'd58523, 16'd25640, 16'd23777, 16'd59511, 16'd29500});
	test_expansion(128'h20ffceb48afc995a84a23d426949e089, {16'd52260, 16'd16461, 16'd55186, 16'd45603, 16'd10503, 16'd21828, 16'd32847, 16'd11551, 16'd65462, 16'd15443, 16'd10781, 16'd77, 16'd50075, 16'd25536, 16'd25862, 16'd65408, 16'd55130, 16'd38866, 16'd7255, 16'd23331, 16'd12466, 16'd38003, 16'd43569, 16'd1702, 16'd53480, 16'd64603});
	test_expansion(128'h4d4f4062b962ea1a1bd8bc10784bb918, {16'd50453, 16'd19236, 16'd29346, 16'd31423, 16'd7885, 16'd39596, 16'd54587, 16'd36761, 16'd39650, 16'd46962, 16'd41494, 16'd35136, 16'd29307, 16'd48472, 16'd17360, 16'd50210, 16'd17409, 16'd18985, 16'd63103, 16'd25039, 16'd52436, 16'd2001, 16'd16877, 16'd35361, 16'd63368, 16'd21681});
	test_expansion(128'hec952c037e3f18a7e70733660bb07005, {16'd55065, 16'd61913, 16'd58864, 16'd35839, 16'd46146, 16'd30853, 16'd65067, 16'd11082, 16'd53141, 16'd55199, 16'd38476, 16'd37049, 16'd52944, 16'd15917, 16'd51275, 16'd16563, 16'd25814, 16'd54622, 16'd11615, 16'd28756, 16'd28683, 16'd39715, 16'd10648, 16'd34538, 16'd37214, 16'd34018});
	test_expansion(128'h708ac88037430ab890c86320730a7483, {16'd48451, 16'd33508, 16'd40038, 16'd1327, 16'd50513, 16'd36164, 16'd27447, 16'd25350, 16'd1579, 16'd13579, 16'd20799, 16'd60725, 16'd50161, 16'd34818, 16'd53211, 16'd22056, 16'd20151, 16'd34174, 16'd10839, 16'd34852, 16'd52190, 16'd51257, 16'd42588, 16'd56438, 16'd47012, 16'd23628});
	test_expansion(128'haf78a8052f13eef8c173dc4e13b32bcb, {16'd3099, 16'd18354, 16'd32172, 16'd31350, 16'd22917, 16'd48402, 16'd33706, 16'd41455, 16'd53260, 16'd17252, 16'd15176, 16'd185, 16'd52040, 16'd44872, 16'd26197, 16'd10270, 16'd39875, 16'd4374, 16'd12896, 16'd42289, 16'd61340, 16'd62083, 16'd62133, 16'd34476, 16'd61179, 16'd30390});
	test_expansion(128'ha5c7750df0c4ebf808d42670297a6625, {16'd59862, 16'd51796, 16'd37282, 16'd29290, 16'd4282, 16'd38041, 16'd19387, 16'd32442, 16'd6623, 16'd19555, 16'd22923, 16'd30, 16'd13989, 16'd16622, 16'd8812, 16'd28830, 16'd50821, 16'd61187, 16'd55148, 16'd12102, 16'd3274, 16'd57485, 16'd10555, 16'd17141, 16'd37677, 16'd18707});
	test_expansion(128'hf7022da7eca774f7d3249d96aa46c6fa, {16'd6130, 16'd38220, 16'd58458, 16'd1143, 16'd32498, 16'd33252, 16'd52557, 16'd48220, 16'd3591, 16'd65065, 16'd57004, 16'd20361, 16'd63775, 16'd39954, 16'd26245, 16'd41327, 16'd61044, 16'd45301, 16'd27920, 16'd35563, 16'd51387, 16'd34702, 16'd53071, 16'd7005, 16'd63196, 16'd40816});
	test_expansion(128'hf7b5a352ddcf7b61cdf99ffbd94d8376, {16'd19132, 16'd9439, 16'd45305, 16'd17485, 16'd32246, 16'd4246, 16'd15427, 16'd55216, 16'd39595, 16'd36870, 16'd26549, 16'd43081, 16'd8247, 16'd58235, 16'd47297, 16'd36117, 16'd32716, 16'd4115, 16'd2313, 16'd50376, 16'd10459, 16'd45811, 16'd54606, 16'd6277, 16'd44097, 16'd5438});
	test_expansion(128'h5cf87e6b70de1ff1ffe5c42b833b7483, {16'd58063, 16'd11391, 16'd20541, 16'd10143, 16'd45290, 16'd48164, 16'd27378, 16'd22844, 16'd41476, 16'd31018, 16'd11914, 16'd24034, 16'd3648, 16'd34732, 16'd47995, 16'd46112, 16'd28921, 16'd22426, 16'd64982, 16'd33158, 16'd33340, 16'd11399, 16'd43367, 16'd36676, 16'd49284, 16'd34168});
	test_expansion(128'h5d66558b60fcc4b8870bc7267f1ca6b5, {16'd18109, 16'd64008, 16'd34895, 16'd30399, 16'd43431, 16'd25972, 16'd43596, 16'd5510, 16'd49378, 16'd49905, 16'd35556, 16'd35866, 16'd65394, 16'd61160, 16'd42513, 16'd61842, 16'd25975, 16'd65212, 16'd37517, 16'd64374, 16'd15744, 16'd23621, 16'd36359, 16'd65525, 16'd21152, 16'd59406});
	test_expansion(128'h830272f4444caeefe473f243ad747a5e, {16'd4589, 16'd50183, 16'd56910, 16'd37709, 16'd21620, 16'd37598, 16'd34529, 16'd47671, 16'd11689, 16'd41576, 16'd58592, 16'd33727, 16'd50233, 16'd60274, 16'd8162, 16'd55863, 16'd54233, 16'd8588, 16'd24019, 16'd56332, 16'd65070, 16'd41180, 16'd38579, 16'd39289, 16'd3723, 16'd12819});
	test_expansion(128'h129685b22b41708be09225a39be67faa, {16'd24795, 16'd45587, 16'd54262, 16'd12356, 16'd45944, 16'd54715, 16'd40656, 16'd15400, 16'd55978, 16'd44197, 16'd48372, 16'd50299, 16'd44286, 16'd48739, 16'd62128, 16'd3503, 16'd44750, 16'd16766, 16'd21315, 16'd418, 16'd9887, 16'd7442, 16'd16808, 16'd42590, 16'd56705, 16'd22176});
	test_expansion(128'hc62097adc059ad7000d59f5e7f4fd143, {16'd12201, 16'd2118, 16'd45147, 16'd7969, 16'd63710, 16'd52427, 16'd42829, 16'd13284, 16'd15478, 16'd52790, 16'd7613, 16'd12482, 16'd28700, 16'd4964, 16'd62743, 16'd59195, 16'd10978, 16'd60079, 16'd28925, 16'd20965, 16'd62888, 16'd28827, 16'd59766, 16'd41847, 16'd46504, 16'd62077});
	test_expansion(128'h354385e2f8136d15127c6c0f53b0e38b, {16'd6915, 16'd25888, 16'd36620, 16'd64128, 16'd4280, 16'd52977, 16'd20295, 16'd21893, 16'd12083, 16'd64806, 16'd62632, 16'd52811, 16'd52127, 16'd54145, 16'd16557, 16'd2091, 16'd48132, 16'd56703, 16'd12046, 16'd6814, 16'd33123, 16'd30763, 16'd65320, 16'd20192, 16'd48869, 16'd60148});
	test_expansion(128'hf24885a3a6ee291d8b5f9ec2bca13910, {16'd47581, 16'd48152, 16'd47478, 16'd49702, 16'd51818, 16'd14791, 16'd52991, 16'd60262, 16'd22888, 16'd1677, 16'd25265, 16'd6733, 16'd4660, 16'd11920, 16'd5341, 16'd17531, 16'd46752, 16'd15245, 16'd17084, 16'd36367, 16'd13565, 16'd61897, 16'd4642, 16'd26894, 16'd18883, 16'd52131});
	test_expansion(128'h2bb9902f2e9ab71ddc6de4b96634837b, {16'd54045, 16'd15383, 16'd22181, 16'd54227, 16'd41465, 16'd36386, 16'd52906, 16'd49245, 16'd57672, 16'd14537, 16'd11286, 16'd28835, 16'd48862, 16'd64238, 16'd41024, 16'd62783, 16'd56040, 16'd4862, 16'd2514, 16'd9099, 16'd34644, 16'd19884, 16'd13110, 16'd38136, 16'd44268, 16'd54612});
	test_expansion(128'h9978c339eb5c09094288fa57591cc73b, {16'd35336, 16'd28023, 16'd34720, 16'd32290, 16'd59262, 16'd24352, 16'd27355, 16'd29832, 16'd63728, 16'd36907, 16'd23776, 16'd33515, 16'd9450, 16'd54198, 16'd35706, 16'd41908, 16'd2436, 16'd1262, 16'd18485, 16'd18619, 16'd9293, 16'd15759, 16'd37409, 16'd39112, 16'd20430, 16'd30925});
	test_expansion(128'h01bba90332b6d0e76edd698031e34ae7, {16'd35560, 16'd22742, 16'd60655, 16'd10362, 16'd16680, 16'd41320, 16'd156, 16'd11777, 16'd27226, 16'd51166, 16'd44458, 16'd24777, 16'd48711, 16'd1877, 16'd40491, 16'd38334, 16'd30511, 16'd63998, 16'd27840, 16'd14748, 16'd18416, 16'd3470, 16'd34563, 16'd28226, 16'd26352, 16'd31368});
	test_expansion(128'h9889061c5070dcc3fa61bc67ff2a2dd2, {16'd4893, 16'd28592, 16'd18436, 16'd37120, 16'd39734, 16'd25408, 16'd43359, 16'd19448, 16'd1701, 16'd10112, 16'd59716, 16'd47945, 16'd26822, 16'd53972, 16'd51730, 16'd32114, 16'd23204, 16'd46559, 16'd28917, 16'd25881, 16'd38200, 16'd5726, 16'd27038, 16'd61942, 16'd36258, 16'd28990});
	test_expansion(128'hd30df877829feb7b5ac3fce8fa2d27bf, {16'd51168, 16'd15504, 16'd21828, 16'd21075, 16'd21490, 16'd43581, 16'd50375, 16'd2591, 16'd13513, 16'd13595, 16'd12414, 16'd1959, 16'd40382, 16'd49023, 16'd16182, 16'd33057, 16'd5020, 16'd31570, 16'd4950, 16'd6350, 16'd5129, 16'd9521, 16'd43476, 16'd11667, 16'd19073, 16'd3557});
	test_expansion(128'hcd462bc4cb77eff48704d5d9dea15af6, {16'd20212, 16'd2712, 16'd17881, 16'd64520, 16'd11143, 16'd22189, 16'd52977, 16'd31397, 16'd36420, 16'd52611, 16'd41848, 16'd21178, 16'd49851, 16'd54719, 16'd50929, 16'd33154, 16'd26303, 16'd22601, 16'd36505, 16'd15975, 16'd65207, 16'd49864, 16'd53463, 16'd52031, 16'd27900, 16'd22179});
	test_expansion(128'hb51f189e6214b37b79ef3c1bb32ba40a, {16'd49984, 16'd8217, 16'd28818, 16'd15019, 16'd31885, 16'd2920, 16'd16020, 16'd44019, 16'd41716, 16'd33208, 16'd40810, 16'd33371, 16'd65332, 16'd37213, 16'd16891, 16'd24638, 16'd25781, 16'd62458, 16'd22790, 16'd28468, 16'd61801, 16'd61973, 16'd28955, 16'd57020, 16'd8291, 16'd44168});
	test_expansion(128'hc62d3223662bf81386ab019e3109d588, {16'd45018, 16'd12730, 16'd53108, 16'd2072, 16'd24833, 16'd57521, 16'd39878, 16'd61961, 16'd32626, 16'd4435, 16'd52302, 16'd28713, 16'd2019, 16'd30624, 16'd29368, 16'd46556, 16'd23893, 16'd51483, 16'd4846, 16'd4889, 16'd18546, 16'd62477, 16'd20006, 16'd22282, 16'd55526, 16'd38740});
	test_expansion(128'h1f53016e788eab040c4079c440456362, {16'd14095, 16'd22284, 16'd62838, 16'd61443, 16'd17505, 16'd20950, 16'd57987, 16'd26039, 16'd331, 16'd40346, 16'd51857, 16'd17197, 16'd51636, 16'd4726, 16'd61820, 16'd8640, 16'd32626, 16'd51546, 16'd57945, 16'd44347, 16'd12174, 16'd15696, 16'd54100, 16'd45425, 16'd11366, 16'd15172});
	test_expansion(128'hcb65aefeeb1cd66a97d2338e2c889488, {16'd63863, 16'd19311, 16'd25066, 16'd18266, 16'd40563, 16'd11694, 16'd61405, 16'd11300, 16'd57503, 16'd5259, 16'd46413, 16'd34352, 16'd11343, 16'd38465, 16'd49242, 16'd18057, 16'd39112, 16'd12414, 16'd57628, 16'd35667, 16'd13936, 16'd48361, 16'd49132, 16'd8704, 16'd44415, 16'd15639});
	test_expansion(128'h1eda1bc6a0933f4e1712f66e88bb01a2, {16'd13818, 16'd54154, 16'd64711, 16'd28039, 16'd28111, 16'd21350, 16'd53220, 16'd42371, 16'd36769, 16'd46884, 16'd16292, 16'd22222, 16'd48774, 16'd8737, 16'd39514, 16'd14428, 16'd28863, 16'd38238, 16'd8000, 16'd23021, 16'd27127, 16'd51424, 16'd63102, 16'd27770, 16'd43343, 16'd22756});
	test_expansion(128'h9b69462aca96affffe37f6324355d56f, {16'd13694, 16'd45004, 16'd54834, 16'd9151, 16'd34639, 16'd45255, 16'd907, 16'd25185, 16'd7387, 16'd28846, 16'd60205, 16'd21710, 16'd56787, 16'd29918, 16'd60779, 16'd47398, 16'd44348, 16'd29698, 16'd17627, 16'd65230, 16'd25832, 16'd20775, 16'd12530, 16'd7785, 16'd29645, 16'd63051});
	test_expansion(128'hc925c67863d9746894e7ae5c81b6f391, {16'd45728, 16'd53990, 16'd40257, 16'd48878, 16'd24985, 16'd56954, 16'd12900, 16'd46252, 16'd58005, 16'd28702, 16'd41872, 16'd50854, 16'd40319, 16'd40957, 16'd523, 16'd30200, 16'd41292, 16'd59109, 16'd42430, 16'd64568, 16'd38639, 16'd57165, 16'd27201, 16'd3137, 16'd22005, 16'd44775});
	test_expansion(128'ha3ab5a734d2b07bce899e0ad6013a475, {16'd29839, 16'd36479, 16'd63456, 16'd56231, 16'd60479, 16'd33099, 16'd35280, 16'd63752, 16'd63539, 16'd39242, 16'd36495, 16'd25905, 16'd18272, 16'd30746, 16'd62768, 16'd14890, 16'd33546, 16'd22778, 16'd60127, 16'd58162, 16'd21400, 16'd40883, 16'd39287, 16'd3236, 16'd10337, 16'd45523});
	test_expansion(128'hbff711a7f186dae645e6f49685e86b37, {16'd32637, 16'd44785, 16'd22454, 16'd18565, 16'd41174, 16'd29953, 16'd23401, 16'd38976, 16'd19446, 16'd52113, 16'd47958, 16'd27052, 16'd41222, 16'd16997, 16'd34938, 16'd35786, 16'd49922, 16'd3890, 16'd31490, 16'd61887, 16'd8898, 16'd24269, 16'd38795, 16'd42902, 16'd5282, 16'd51342});
	test_expansion(128'h0e53dffadcd3991a736a31dcf28d4491, {16'd55772, 16'd40357, 16'd5684, 16'd33383, 16'd4415, 16'd31165, 16'd44339, 16'd22090, 16'd8405, 16'd7460, 16'd42364, 16'd63227, 16'd26460, 16'd33650, 16'd41346, 16'd39476, 16'd61604, 16'd4786, 16'd45650, 16'd7249, 16'd61365, 16'd35117, 16'd18705, 16'd46234, 16'd27702, 16'd51219});
	test_expansion(128'hd47df56e45c41e61840a317acf128643, {16'd38737, 16'd2443, 16'd17820, 16'd32677, 16'd45025, 16'd19079, 16'd39465, 16'd28091, 16'd56709, 16'd20884, 16'd20263, 16'd53835, 16'd34228, 16'd6193, 16'd38432, 16'd65054, 16'd63980, 16'd38591, 16'd48109, 16'd57792, 16'd299, 16'd39923, 16'd48299, 16'd51381, 16'd19376, 16'd48139});
	test_expansion(128'h31df58de3d78211ea6c4cc4c57e007bd, {16'd53482, 16'd43940, 16'd62435, 16'd44710, 16'd26582, 16'd40535, 16'd37740, 16'd25360, 16'd50939, 16'd49974, 16'd60435, 16'd21179, 16'd5673, 16'd21841, 16'd6636, 16'd36934, 16'd48499, 16'd4109, 16'd29042, 16'd60975, 16'd12301, 16'd51660, 16'd57669, 16'd47097, 16'd6740, 16'd50119});
	test_expansion(128'ha46962f8770d777fb719770e0bb72fc8, {16'd43844, 16'd19259, 16'd37891, 16'd39394, 16'd39619, 16'd43273, 16'd35537, 16'd64460, 16'd11176, 16'd1904, 16'd49069, 16'd42996, 16'd11119, 16'd28622, 16'd38580, 16'd57881, 16'd53793, 16'd37702, 16'd33149, 16'd36756, 16'd13381, 16'd49777, 16'd50542, 16'd14841, 16'd39484, 16'd37025});
	test_expansion(128'hddf219c2f9e162c5e93e89c684f3d6a9, {16'd1415, 16'd20998, 16'd7928, 16'd216, 16'd31354, 16'd55003, 16'd29484, 16'd47966, 16'd59633, 16'd47925, 16'd52436, 16'd58908, 16'd33027, 16'd16641, 16'd59553, 16'd13986, 16'd11911, 16'd39478, 16'd64032, 16'd54282, 16'd61899, 16'd24443, 16'd4044, 16'd13088, 16'd43064, 16'd33907});
	test_expansion(128'hcf7d40e7219a9bcae9dfee0102632236, {16'd32754, 16'd4260, 16'd2977, 16'd38255, 16'd29978, 16'd5857, 16'd40669, 16'd35430, 16'd22545, 16'd46468, 16'd31263, 16'd33573, 16'd16142, 16'd58569, 16'd18116, 16'd6116, 16'd11237, 16'd17201, 16'd15925, 16'd55480, 16'd62701, 16'd60307, 16'd36707, 16'd14615, 16'd19911, 16'd51653});
	test_expansion(128'hf5d1ebe2632d8de51db0c73a4df1e479, {16'd43950, 16'd53074, 16'd2225, 16'd47917, 16'd8924, 16'd41106, 16'd57893, 16'd57430, 16'd6631, 16'd5188, 16'd3187, 16'd59291, 16'd45406, 16'd17207, 16'd62555, 16'd1356, 16'd29528, 16'd48689, 16'd65466, 16'd13543, 16'd53049, 16'd1436, 16'd57245, 16'd12208, 16'd52724, 16'd6657});
	test_expansion(128'hb3776554f9f8b94d41328a6b42044f76, {16'd7098, 16'd40520, 16'd23404, 16'd38474, 16'd56385, 16'd9291, 16'd41794, 16'd18414, 16'd20657, 16'd35267, 16'd47008, 16'd22845, 16'd40426, 16'd6280, 16'd32069, 16'd53131, 16'd37135, 16'd6513, 16'd55670, 16'd19695, 16'd9065, 16'd32572, 16'd3159, 16'd24445, 16'd15079, 16'd4839});
	test_expansion(128'hb15b53d97d596ce2fe5d8da865816f69, {16'd33126, 16'd44747, 16'd4482, 16'd20941, 16'd1374, 16'd30095, 16'd5088, 16'd26306, 16'd34967, 16'd33852, 16'd54191, 16'd9389, 16'd39107, 16'd38598, 16'd24703, 16'd28599, 16'd32422, 16'd39814, 16'd46374, 16'd7678, 16'd36739, 16'd39975, 16'd19721, 16'd38835, 16'd29761, 16'd27141});
	test_expansion(128'h0064c48a33a55ce5b738da6677b84f93, {16'd53214, 16'd24536, 16'd17567, 16'd58399, 16'd9889, 16'd33342, 16'd48595, 16'd42116, 16'd64518, 16'd38913, 16'd38917, 16'd239, 16'd10726, 16'd64373, 16'd31862, 16'd62956, 16'd30496, 16'd37608, 16'd1386, 16'd36511, 16'd28387, 16'd51174, 16'd62518, 16'd28289, 16'd15780, 16'd51507});
	test_expansion(128'h34e94d82daa889d5911f109a3c73c2f8, {16'd11673, 16'd5581, 16'd38494, 16'd31071, 16'd34767, 16'd31593, 16'd52877, 16'd43051, 16'd16618, 16'd38852, 16'd26475, 16'd29265, 16'd16363, 16'd53630, 16'd30057, 16'd54570, 16'd43060, 16'd8192, 16'd45312, 16'd58643, 16'd55422, 16'd33292, 16'd63432, 16'd3027, 16'd53087, 16'd17957});
	test_expansion(128'hb4fae3b85b1d364b481b3eae725db6ac, {16'd35498, 16'd7942, 16'd26265, 16'd10477, 16'd45132, 16'd49699, 16'd56959, 16'd64155, 16'd28262, 16'd58066, 16'd8531, 16'd3661, 16'd51212, 16'd36932, 16'd41390, 16'd12414, 16'd24523, 16'd48484, 16'd4261, 16'd58134, 16'd33455, 16'd1637, 16'd34981, 16'd41892, 16'd7551, 16'd46915});
	test_expansion(128'ha0b621248cb53f4232cddbce3636d5de, {16'd13506, 16'd44093, 16'd19165, 16'd45041, 16'd6104, 16'd38575, 16'd41902, 16'd54664, 16'd11001, 16'd16378, 16'd50963, 16'd21299, 16'd28031, 16'd14765, 16'd11641, 16'd20670, 16'd12951, 16'd25475, 16'd9655, 16'd14999, 16'd43229, 16'd33392, 16'd62357, 16'd52250, 16'd41549, 16'd24530});
	test_expansion(128'h73d196a44b8e486bd5c33e200af7751c, {16'd43027, 16'd55315, 16'd38986, 16'd41330, 16'd13783, 16'd32890, 16'd41803, 16'd52189, 16'd27403, 16'd19283, 16'd183, 16'd40070, 16'd42357, 16'd59918, 16'd18823, 16'd58229, 16'd31291, 16'd2100, 16'd14921, 16'd58090, 16'd33784, 16'd49334, 16'd38491, 16'd28434, 16'd15237, 16'd37252});
	test_expansion(128'h831e60b531600181f5f89590b469ef21, {16'd57496, 16'd11440, 16'd48496, 16'd2906, 16'd48010, 16'd2096, 16'd52754, 16'd30641, 16'd64802, 16'd16027, 16'd9850, 16'd42788, 16'd64516, 16'd56092, 16'd20604, 16'd44433, 16'd63267, 16'd46569, 16'd62765, 16'd59572, 16'd51469, 16'd2515, 16'd19987, 16'd27959, 16'd37141, 16'd40033});
	test_expansion(128'h7a8abaee243d880955acaaf2eb5251e1, {16'd13331, 16'd10250, 16'd2223, 16'd21921, 16'd16667, 16'd41909, 16'd3363, 16'd62279, 16'd46744, 16'd19565, 16'd30250, 16'd51249, 16'd17551, 16'd10217, 16'd19913, 16'd17643, 16'd64942, 16'd43498, 16'd42981, 16'd10157, 16'd53678, 16'd45412, 16'd13792, 16'd61515, 16'd40290, 16'd42421});
	test_expansion(128'hf2b989525376e82b38e5aa322c56a9b4, {16'd23818, 16'd13833, 16'd22094, 16'd57090, 16'd65280, 16'd22793, 16'd55546, 16'd42666, 16'd22203, 16'd16839, 16'd12799, 16'd24551, 16'd51412, 16'd7407, 16'd9744, 16'd16105, 16'd7814, 16'd6320, 16'd22569, 16'd57933, 16'd61519, 16'd31748, 16'd59897, 16'd16508, 16'd42796, 16'd14706});
	test_expansion(128'hea182fa1335d6a20d15495bff17c69ad, {16'd3699, 16'd38601, 16'd39907, 16'd10698, 16'd37481, 16'd667, 16'd55453, 16'd29133, 16'd4943, 16'd26711, 16'd33153, 16'd20543, 16'd23825, 16'd22438, 16'd63671, 16'd10577, 16'd2728, 16'd3911, 16'd442, 16'd11470, 16'd1764, 16'd57587, 16'd18237, 16'd41828, 16'd41265, 16'd55105});
	test_expansion(128'he000c962190082a573056e029507d58b, {16'd23590, 16'd48484, 16'd2309, 16'd53503, 16'd12030, 16'd7587, 16'd61616, 16'd13190, 16'd49248, 16'd35060, 16'd22739, 16'd52099, 16'd50775, 16'd19984, 16'd59502, 16'd37162, 16'd3600, 16'd53618, 16'd22454, 16'd31848, 16'd26095, 16'd29423, 16'd47263, 16'd11520, 16'd40435, 16'd46913});
	test_expansion(128'h6d8023faeea68d7072459179b39a38e1, {16'd62302, 16'd41298, 16'd42756, 16'd17000, 16'd49859, 16'd18207, 16'd59906, 16'd15656, 16'd32294, 16'd27438, 16'd50678, 16'd56981, 16'd12231, 16'd909, 16'd12116, 16'd9647, 16'd20428, 16'd62871, 16'd54174, 16'd1605, 16'd1814, 16'd10928, 16'd13770, 16'd61456, 16'd34741, 16'd4935});
	test_expansion(128'h2c4c5ba518d7066aada1d28ea3dfc12c, {16'd44925, 16'd634, 16'd28559, 16'd36856, 16'd47291, 16'd48734, 16'd32768, 16'd46699, 16'd62297, 16'd46768, 16'd57843, 16'd14977, 16'd45940, 16'd38731, 16'd24623, 16'd12247, 16'd51700, 16'd41206, 16'd54519, 16'd5573, 16'd65533, 16'd36914, 16'd64930, 16'd55665, 16'd16362, 16'd57961});
	test_expansion(128'hc992c72a11874ada0077b459ca5562c3, {16'd8052, 16'd32133, 16'd24893, 16'd2634, 16'd42826, 16'd7987, 16'd1829, 16'd47119, 16'd39505, 16'd57490, 16'd8450, 16'd17573, 16'd264, 16'd41068, 16'd6362, 16'd25192, 16'd33523, 16'd26379, 16'd40712, 16'd14671, 16'd52645, 16'd3662, 16'd47034, 16'd45526, 16'd44899, 16'd51336});
	test_expansion(128'h5bab352a30cc2645b80638300971c6e4, {16'd15129, 16'd19111, 16'd52399, 16'd47151, 16'd35784, 16'd3354, 16'd51012, 16'd25925, 16'd62534, 16'd49077, 16'd62311, 16'd52827, 16'd42522, 16'd37646, 16'd8814, 16'd1007, 16'd64668, 16'd26258, 16'd60678, 16'd33327, 16'd34233, 16'd14362, 16'd26759, 16'd7982, 16'd8790, 16'd55259});
	test_expansion(128'hc9a39e1e2c3189e04e0ce2572be4075c, {16'd9709, 16'd26388, 16'd46200, 16'd14397, 16'd803, 16'd39436, 16'd49140, 16'd26421, 16'd46917, 16'd9790, 16'd1264, 16'd54346, 16'd58375, 16'd48489, 16'd45975, 16'd64409, 16'd18512, 16'd53132, 16'd12980, 16'd50309, 16'd59853, 16'd30332, 16'd62332, 16'd9302, 16'd34605, 16'd59904});
	test_expansion(128'he604f59cb17f51f351394f0543176ea3, {16'd54840, 16'd31045, 16'd17926, 16'd25182, 16'd29201, 16'd23576, 16'd31860, 16'd5832, 16'd11611, 16'd40790, 16'd53708, 16'd21761, 16'd6222, 16'd34887, 16'd13317, 16'd21658, 16'd48828, 16'd31633, 16'd14263, 16'd54238, 16'd35159, 16'd63132, 16'd46867, 16'd52932, 16'd6566, 16'd46583});
	test_expansion(128'h9edfc87fafad192a437a4785e47bc95e, {16'd54493, 16'd57398, 16'd31000, 16'd36478, 16'd62255, 16'd31119, 16'd62500, 16'd22766, 16'd25276, 16'd33858, 16'd44614, 16'd8119, 16'd7536, 16'd48329, 16'd10598, 16'd40119, 16'd60705, 16'd10293, 16'd38580, 16'd45263, 16'd33406, 16'd15973, 16'd53892, 16'd39725, 16'd585, 16'd17957});
	test_expansion(128'hb73a844a98a2556c7c966972a3cd9085, {16'd42965, 16'd42190, 16'd5448, 16'd59833, 16'd65501, 16'd64663, 16'd26274, 16'd40141, 16'd22153, 16'd30085, 16'd49171, 16'd21429, 16'd28917, 16'd24378, 16'd7662, 16'd22013, 16'd31959, 16'd50785, 16'd43243, 16'd15662, 16'd53908, 16'd58886, 16'd44534, 16'd49197, 16'd50951, 16'd56767});
	test_expansion(128'hb00f0ea537805b4306ef9a3fd60b3474, {16'd46247, 16'd32511, 16'd12958, 16'd39495, 16'd16861, 16'd64394, 16'd19747, 16'd29841, 16'd50223, 16'd44941, 16'd39870, 16'd51070, 16'd20008, 16'd59736, 16'd536, 16'd54397, 16'd62941, 16'd24117, 16'd29550, 16'd43562, 16'd15026, 16'd34450, 16'd49525, 16'd64205, 16'd30615, 16'd61812});
	test_expansion(128'hcff3fe9e3b78303655569e40c32cdb09, {16'd65314, 16'd39016, 16'd35766, 16'd42956, 16'd29747, 16'd34491, 16'd8539, 16'd48753, 16'd6163, 16'd41171, 16'd27820, 16'd52317, 16'd55118, 16'd10029, 16'd33865, 16'd23494, 16'd30110, 16'd53411, 16'd21309, 16'd50285, 16'd14992, 16'd34882, 16'd13431, 16'd37881, 16'd38779, 16'd4114});
	test_expansion(128'hbe550145e0800b734d3348df29cf4b4d, {16'd53827, 16'd63091, 16'd37744, 16'd33269, 16'd43314, 16'd50965, 16'd29500, 16'd7739, 16'd35361, 16'd45060, 16'd46714, 16'd31955, 16'd10971, 16'd50404, 16'd2063, 16'd7377, 16'd7557, 16'd23572, 16'd27234, 16'd1577, 16'd52764, 16'd45538, 16'd21810, 16'd9215, 16'd17928, 16'd39234});
	test_expansion(128'hfdc0826314827f63ce45309f94e89332, {16'd30122, 16'd19103, 16'd28040, 16'd21410, 16'd57201, 16'd32359, 16'd33636, 16'd17089, 16'd11932, 16'd34254, 16'd41468, 16'd15190, 16'd19431, 16'd4654, 16'd57787, 16'd15929, 16'd13975, 16'd51957, 16'd10062, 16'd64120, 16'd12383, 16'd49277, 16'd40352, 16'd32042, 16'd9405, 16'd26838});
	test_expansion(128'h9aba644271094f80d98d247f2d1d70f7, {16'd57025, 16'd50901, 16'd49240, 16'd51462, 16'd3194, 16'd22708, 16'd61485, 16'd17714, 16'd1221, 16'd43091, 16'd63492, 16'd38183, 16'd62854, 16'd42791, 16'd46320, 16'd43997, 16'd549, 16'd2989, 16'd37925, 16'd19635, 16'd52903, 16'd49927, 16'd12842, 16'd7924, 16'd15977, 16'd40844});
	test_expansion(128'h8d114da7b7471115468cbec819bd32f4, {16'd4088, 16'd62543, 16'd61728, 16'd60418, 16'd42784, 16'd4215, 16'd17365, 16'd7924, 16'd48643, 16'd10375, 16'd45191, 16'd36646, 16'd10849, 16'd59224, 16'd48797, 16'd37724, 16'd4870, 16'd12321, 16'd1341, 16'd51524, 16'd13090, 16'd39640, 16'd35686, 16'd40601, 16'd22168, 16'd21169});
	test_expansion(128'h6251e93585981a7561246a696d66bf09, {16'd50784, 16'd30943, 16'd5771, 16'd42896, 16'd30623, 16'd45705, 16'd6317, 16'd11966, 16'd33156, 16'd27990, 16'd317, 16'd36658, 16'd26932, 16'd41970, 16'd48204, 16'd35368, 16'd2253, 16'd7834, 16'd30881, 16'd4596, 16'd30987, 16'd16739, 16'd21022, 16'd19284, 16'd29105, 16'd44100});
	test_expansion(128'h53062dfbadec034a266f1f19f1ed3d9b, {16'd18175, 16'd48642, 16'd27645, 16'd2000, 16'd18791, 16'd16540, 16'd63388, 16'd30467, 16'd42402, 16'd3151, 16'd49567, 16'd29932, 16'd17186, 16'd12955, 16'd35798, 16'd9527, 16'd59319, 16'd48209, 16'd29382, 16'd19087, 16'd63129, 16'd35768, 16'd27314, 16'd21813, 16'd39640, 16'd42766});
	test_expansion(128'h289f4d8ecd2e1e3ecd8626aae91c04f7, {16'd4313, 16'd8788, 16'd11329, 16'd17467, 16'd40122, 16'd20855, 16'd47528, 16'd52943, 16'd52293, 16'd54297, 16'd41698, 16'd14247, 16'd16146, 16'd61528, 16'd24369, 16'd38539, 16'd38149, 16'd51267, 16'd46908, 16'd42707, 16'd55924, 16'd32224, 16'd33776, 16'd62058, 16'd46518, 16'd12460});
	test_expansion(128'h96ea6932b0366c741b16193b1980acd2, {16'd10420, 16'd4522, 16'd28718, 16'd30666, 16'd15162, 16'd39284, 16'd60149, 16'd58998, 16'd56128, 16'd56532, 16'd3233, 16'd59215, 16'd39558, 16'd36857, 16'd48170, 16'd30045, 16'd49809, 16'd3120, 16'd7469, 16'd42777, 16'd51748, 16'd58266, 16'd49880, 16'd37352, 16'd34037, 16'd53667});
	test_expansion(128'h21adcc5a3e458d942c80b4bfed02d910, {16'd33007, 16'd27898, 16'd35681, 16'd2940, 16'd9650, 16'd27081, 16'd31679, 16'd48078, 16'd42360, 16'd21161, 16'd65281, 16'd44975, 16'd42732, 16'd23539, 16'd47805, 16'd56344, 16'd28734, 16'd48090, 16'd30216, 16'd17000, 16'd670, 16'd41679, 16'd37415, 16'd41212, 16'd3772, 16'd14706});
	test_expansion(128'h8b78c0b2b6d5a0e736b4677765549154, {16'd7145, 16'd19912, 16'd21527, 16'd52707, 16'd20193, 16'd48453, 16'd3716, 16'd3538, 16'd890, 16'd43628, 16'd56470, 16'd43146, 16'd20041, 16'd34900, 16'd45172, 16'd14407, 16'd48029, 16'd40070, 16'd53345, 16'd9163, 16'd64487, 16'd421, 16'd51631, 16'd36449, 16'd59938, 16'd28821});
	test_expansion(128'h650c7c712943dd073a8e68922fe078b7, {16'd23824, 16'd63952, 16'd61247, 16'd2199, 16'd45550, 16'd26238, 16'd38399, 16'd42338, 16'd14296, 16'd23287, 16'd31589, 16'd61980, 16'd12470, 16'd59924, 16'd32557, 16'd64822, 16'd53223, 16'd32447, 16'd38748, 16'd14895, 16'd31397, 16'd12957, 16'd7594, 16'd53559, 16'd58830, 16'd41727});
	test_expansion(128'h7542129423aa97b22c3e6c31887f7165, {16'd1389, 16'd17606, 16'd31086, 16'd30118, 16'd63606, 16'd15534, 16'd11493, 16'd44386, 16'd20163, 16'd54816, 16'd56199, 16'd50083, 16'd46339, 16'd3320, 16'd58306, 16'd23398, 16'd11888, 16'd31841, 16'd3695, 16'd51437, 16'd19854, 16'd7614, 16'd19902, 16'd51333, 16'd36055, 16'd10605});
	test_expansion(128'h1a00159ce331806e8a7e579ad997f861, {16'd51957, 16'd3995, 16'd55476, 16'd58112, 16'd43844, 16'd2206, 16'd34464, 16'd63652, 16'd40112, 16'd16858, 16'd62040, 16'd3558, 16'd39507, 16'd43684, 16'd18375, 16'd52416, 16'd44083, 16'd3424, 16'd43069, 16'd60996, 16'd53657, 16'd18486, 16'd18320, 16'd49479, 16'd2013, 16'd39293});
	test_expansion(128'h023131b67ab2533b26ce41e99237f0f3, {16'd65420, 16'd43846, 16'd30787, 16'd49151, 16'd22385, 16'd4989, 16'd23274, 16'd21462, 16'd39868, 16'd39610, 16'd39471, 16'd50158, 16'd13677, 16'd14086, 16'd6181, 16'd21418, 16'd64680, 16'd29360, 16'd47664, 16'd40749, 16'd62118, 16'd51432, 16'd4217, 16'd40014, 16'd30124, 16'd43519});
	test_expansion(128'hc63672f4184cf513af224949ce7e84c7, {16'd14832, 16'd62932, 16'd30357, 16'd63590, 16'd60094, 16'd52851, 16'd8511, 16'd4326, 16'd7182, 16'd52963, 16'd40067, 16'd48150, 16'd44258, 16'd64791, 16'd9823, 16'd11361, 16'd3801, 16'd28311, 16'd51241, 16'd11462, 16'd11678, 16'd15697, 16'd59159, 16'd23084, 16'd46340, 16'd33847});
	test_expansion(128'h3f7b4678107a2a919f0eac22a4acf2c1, {16'd53938, 16'd36685, 16'd55821, 16'd49100, 16'd28072, 16'd27802, 16'd8271, 16'd7225, 16'd44883, 16'd61917, 16'd32761, 16'd45613, 16'd64168, 16'd62266, 16'd5624, 16'd29966, 16'd14145, 16'd18093, 16'd17439, 16'd60368, 16'd38330, 16'd26879, 16'd64087, 16'd64208, 16'd47227, 16'd14129});
	test_expansion(128'hbcca9b0a31896f2150f426bd849fab9d, {16'd41479, 16'd58683, 16'd49512, 16'd46581, 16'd55702, 16'd49484, 16'd7905, 16'd6373, 16'd2341, 16'd57331, 16'd41568, 16'd49782, 16'd22168, 16'd55410, 16'd39082, 16'd4585, 16'd27856, 16'd9288, 16'd51647, 16'd43747, 16'd62237, 16'd17862, 16'd1029, 16'd44741, 16'd63797, 16'd46683});
	test_expansion(128'h18f772e0b3b142a6f40b954aa6087724, {16'd51868, 16'd53058, 16'd46054, 16'd57719, 16'd40709, 16'd26471, 16'd43567, 16'd62232, 16'd24348, 16'd19847, 16'd2226, 16'd57019, 16'd11448, 16'd63456, 16'd36304, 16'd25694, 16'd38336, 16'd42253, 16'd57368, 16'd59719, 16'd36244, 16'd9344, 16'd15761, 16'd3858, 16'd28493, 16'd7749});
	test_expansion(128'h8dcc6182388b7864d3b11fdf20af6355, {16'd8252, 16'd10698, 16'd14976, 16'd59156, 16'd32371, 16'd23053, 16'd30834, 16'd9494, 16'd36644, 16'd22446, 16'd29482, 16'd52318, 16'd7756, 16'd59325, 16'd1327, 16'd34303, 16'd907, 16'd43040, 16'd27127, 16'd13069, 16'd9812, 16'd53663, 16'd38978, 16'd50489, 16'd5379, 16'd39021});
	test_expansion(128'h4de5b2574d940c0cec6e6c62936e0d95, {16'd15255, 16'd44718, 16'd61265, 16'd36279, 16'd45630, 16'd8101, 16'd21301, 16'd1555, 16'd35495, 16'd11466, 16'd45402, 16'd58385, 16'd20427, 16'd18971, 16'd30564, 16'd52258, 16'd9214, 16'd33735, 16'd15518, 16'd47988, 16'd53895, 16'd23079, 16'd38838, 16'd372, 16'd65359, 16'd18217});
	test_expansion(128'hc488bdecdcf526673db898df0b5e29d0, {16'd36951, 16'd47409, 16'd14369, 16'd34788, 16'd40944, 16'd52590, 16'd48481, 16'd55132, 16'd58535, 16'd65509, 16'd41428, 16'd44544, 16'd21872, 16'd38828, 16'd51841, 16'd48222, 16'd34921, 16'd55291, 16'd3415, 16'd47100, 16'd42884, 16'd33828, 16'd45550, 16'd33934, 16'd59810, 16'd10211});
	test_expansion(128'h8114a482f29253023389b676aecff0ec, {16'd60905, 16'd16538, 16'd28830, 16'd10153, 16'd23166, 16'd38321, 16'd6167, 16'd9858, 16'd4937, 16'd36381, 16'd16487, 16'd29812, 16'd46720, 16'd49718, 16'd23553, 16'd22157, 16'd40936, 16'd10028, 16'd7327, 16'd56084, 16'd34138, 16'd57712, 16'd14821, 16'd40624, 16'd7875, 16'd35034});
	test_expansion(128'h0d97fad0983935427941ccea84383ea8, {16'd37534, 16'd44884, 16'd55108, 16'd41530, 16'd15474, 16'd32896, 16'd27702, 16'd40807, 16'd34356, 16'd3535, 16'd52349, 16'd57311, 16'd10878, 16'd16430, 16'd39747, 16'd18617, 16'd26747, 16'd30406, 16'd24051, 16'd15799, 16'd30782, 16'd39674, 16'd34628, 16'd23383, 16'd48959, 16'd16475});
	test_expansion(128'h0a7c944e1edd70701ff48eff7c1dda3b, {16'd27161, 16'd24138, 16'd5421, 16'd33501, 16'd46027, 16'd24229, 16'd62580, 16'd14165, 16'd18086, 16'd60251, 16'd39075, 16'd54510, 16'd24177, 16'd62845, 16'd64574, 16'd33695, 16'd36879, 16'd30280, 16'd61492, 16'd53703, 16'd56500, 16'd54892, 16'd36751, 16'd31943, 16'd29218, 16'd50774});
	test_expansion(128'h609bfc6871e7549905182472826605cb, {16'd536, 16'd42256, 16'd34301, 16'd41570, 16'd10740, 16'd24605, 16'd59921, 16'd10075, 16'd31986, 16'd33747, 16'd33791, 16'd41549, 16'd12353, 16'd4610, 16'd55885, 16'd27053, 16'd34251, 16'd40168, 16'd41588, 16'd53238, 16'd45330, 16'd101, 16'd32007, 16'd43870, 16'd13145, 16'd41079});
	test_expansion(128'hbb6d82bfb01d08b86616482dbd332e03, {16'd18092, 16'd64626, 16'd46694, 16'd24219, 16'd10630, 16'd55069, 16'd24681, 16'd13608, 16'd41074, 16'd60235, 16'd49927, 16'd28644, 16'd35425, 16'd53399, 16'd23374, 16'd23779, 16'd8146, 16'd28454, 16'd9808, 16'd57212, 16'd7343, 16'd20572, 16'd35086, 16'd31301, 16'd58454, 16'd59276});
	test_expansion(128'hfa7c7823178f621c980feb05ce7d6c8a, {16'd37448, 16'd58018, 16'd1753, 16'd37922, 16'd18381, 16'd13153, 16'd51932, 16'd41217, 16'd788, 16'd61921, 16'd58854, 16'd26837, 16'd3065, 16'd54214, 16'd27391, 16'd6465, 16'd53387, 16'd65483, 16'd5025, 16'd50224, 16'd7908, 16'd43907, 16'd37920, 16'd4643, 16'd22094, 16'd64022});
	test_expansion(128'hc4dfca0cd43edffe1e34467491a21d8f, {16'd14043, 16'd53820, 16'd20819, 16'd26479, 16'd27019, 16'd56109, 16'd39643, 16'd29460, 16'd40666, 16'd9205, 16'd59204, 16'd36594, 16'd43503, 16'd50388, 16'd56826, 16'd36465, 16'd32202, 16'd19899, 16'd57279, 16'd7450, 16'd27569, 16'd53480, 16'd3304, 16'd17387, 16'd37413, 16'd9108});
	test_expansion(128'h7c150f00e4307a2466f9bc5361a79a2a, {16'd16854, 16'd34360, 16'd24172, 16'd33242, 16'd34098, 16'd55306, 16'd29126, 16'd11891, 16'd28898, 16'd3156, 16'd64050, 16'd883, 16'd36672, 16'd37387, 16'd10065, 16'd30917, 16'd65508, 16'd58903, 16'd35348, 16'd39098, 16'd61518, 16'd42928, 16'd29037, 16'd39210, 16'd54754, 16'd4596});
	test_expansion(128'h6cc3ef055185acd7039d9b30aae34adb, {16'd54639, 16'd25121, 16'd62785, 16'd31054, 16'd26517, 16'd51143, 16'd6231, 16'd63249, 16'd50807, 16'd13079, 16'd34540, 16'd56826, 16'd33340, 16'd37360, 16'd18892, 16'd11240, 16'd48007, 16'd38854, 16'd22107, 16'd15028, 16'd31018, 16'd27548, 16'd23271, 16'd24550, 16'd48465, 16'd63173});
	test_expansion(128'ha34bf5b54c0d96adaa9693a38f5778e0, {16'd8527, 16'd41434, 16'd7767, 16'd29994, 16'd32481, 16'd28651, 16'd52615, 16'd30339, 16'd11855, 16'd35671, 16'd55033, 16'd2023, 16'd3243, 16'd40283, 16'd21639, 16'd53951, 16'd36740, 16'd14356, 16'd3308, 16'd27288, 16'd23358, 16'd34950, 16'd36006, 16'd59727, 16'd33860, 16'd39142});
	test_expansion(128'h35da1a61136bc31fe0fa35564f870199, {16'd12482, 16'd27787, 16'd4003, 16'd47338, 16'd60946, 16'd10309, 16'd17084, 16'd11406, 16'd61675, 16'd52696, 16'd31697, 16'd44500, 16'd60185, 16'd50516, 16'd43154, 16'd21588, 16'd50153, 16'd5481, 16'd26224, 16'd10216, 16'd56936, 16'd55760, 16'd13659, 16'd28327, 16'd14061, 16'd24712});
	test_expansion(128'h7997396ce246440b955a3c3b9b2bb4dd, {16'd35975, 16'd65126, 16'd36545, 16'd58640, 16'd24323, 16'd35121, 16'd45087, 16'd61665, 16'd42211, 16'd55093, 16'd37899, 16'd46763, 16'd47498, 16'd58565, 16'd59930, 16'd6505, 16'd49897, 16'd62854, 16'd58844, 16'd59347, 16'd20846, 16'd25983, 16'd39622, 16'd21858, 16'd3233, 16'd26257});
	test_expansion(128'hd45470b36277b7f5f839be907ebeb9ba, {16'd34248, 16'd45537, 16'd65431, 16'd21534, 16'd11648, 16'd3880, 16'd19237, 16'd42118, 16'd55795, 16'd4236, 16'd41880, 16'd61646, 16'd55008, 16'd6594, 16'd24195, 16'd35590, 16'd51008, 16'd16419, 16'd39794, 16'd55239, 16'd22464, 16'd16194, 16'd26195, 16'd57406, 16'd63371, 16'd30815});
	test_expansion(128'h239ca3f5b28395ddd8ae256c0e34ec39, {16'd36210, 16'd12047, 16'd38949, 16'd15984, 16'd3546, 16'd40636, 16'd50595, 16'd52655, 16'd62628, 16'd23375, 16'd8237, 16'd11930, 16'd41714, 16'd51250, 16'd38121, 16'd29470, 16'd15623, 16'd44749, 16'd13119, 16'd5057, 16'd1971, 16'd30022, 16'd7713, 16'd4706, 16'd27259, 16'd64062});
	test_expansion(128'hbc4eb08172635943135735df23ce2f89, {16'd27533, 16'd12308, 16'd6277, 16'd47025, 16'd60004, 16'd48216, 16'd46802, 16'd43898, 16'd58462, 16'd13229, 16'd37456, 16'd51352, 16'd59668, 16'd51961, 16'd1098, 16'd21380, 16'd16628, 16'd12045, 16'd8679, 16'd825, 16'd17974, 16'd6525, 16'd21316, 16'd46456, 16'd9669, 16'd48351});
	test_expansion(128'h603500d0fde9f2aca40bf1ede7a0fd2b, {16'd50815, 16'd59805, 16'd28590, 16'd19392, 16'd48736, 16'd40068, 16'd7342, 16'd16750, 16'd3851, 16'd38801, 16'd52086, 16'd4709, 16'd56371, 16'd34221, 16'd10528, 16'd12977, 16'd30282, 16'd50014, 16'd19028, 16'd25604, 16'd39918, 16'd41280, 16'd18648, 16'd31700, 16'd32393, 16'd58380});
	test_expansion(128'hb91948847918a83d421b0d3b97257b1d, {16'd22903, 16'd62147, 16'd4221, 16'd31627, 16'd10009, 16'd24234, 16'd42360, 16'd8601, 16'd27616, 16'd30784, 16'd58343, 16'd22026, 16'd13235, 16'd45745, 16'd58704, 16'd63203, 16'd46581, 16'd32935, 16'd35639, 16'd58602, 16'd64879, 16'd62587, 16'd50474, 16'd37589, 16'd59834, 16'd12460});
	test_expansion(128'h3e748559da37430e49e5f3357eb46d8d, {16'd38881, 16'd42616, 16'd4442, 16'd59681, 16'd21616, 16'd30126, 16'd64080, 16'd46315, 16'd9706, 16'd29873, 16'd13147, 16'd37628, 16'd61180, 16'd16050, 16'd24782, 16'd5109, 16'd19381, 16'd40237, 16'd17160, 16'd25, 16'd33939, 16'd37499, 16'd25641, 16'd37869, 16'd54021, 16'd13751});
	test_expansion(128'h3416dfdf4d735f946d1d7e832cc05bf7, {16'd48888, 16'd54374, 16'd6957, 16'd14118, 16'd53377, 16'd41958, 16'd60193, 16'd17659, 16'd541, 16'd55188, 16'd43916, 16'd49817, 16'd1703, 16'd31254, 16'd233, 16'd32456, 16'd26575, 16'd1295, 16'd50958, 16'd11937, 16'd8409, 16'd64916, 16'd61272, 16'd42460, 16'd21704, 16'd34769});
	test_expansion(128'h64fc075e47a9dbe1067195c1ee0f92bf, {16'd44798, 16'd39044, 16'd10579, 16'd43333, 16'd14720, 16'd30004, 16'd63198, 16'd51098, 16'd49634, 16'd58410, 16'd3775, 16'd44067, 16'd52470, 16'd59155, 16'd23882, 16'd13538, 16'd18525, 16'd61984, 16'd32227, 16'd25908, 16'd46011, 16'd51516, 16'd8785, 16'd51808, 16'd5893, 16'd61063});
	test_expansion(128'hfe016aae68c8bbfcee714747490b4055, {16'd61186, 16'd20496, 16'd22873, 16'd4299, 16'd24825, 16'd65298, 16'd44257, 16'd52110, 16'd13547, 16'd33339, 16'd7738, 16'd26887, 16'd62266, 16'd14488, 16'd5192, 16'd4222, 16'd3795, 16'd60331, 16'd7206, 16'd60922, 16'd42052, 16'd61231, 16'd18936, 16'd23576, 16'd56349, 16'd19263});
	test_expansion(128'h610bec892b1a7d9c445246fdefeaaa97, {16'd32432, 16'd17379, 16'd45993, 16'd11642, 16'd20959, 16'd62357, 16'd51111, 16'd53394, 16'd52118, 16'd206, 16'd7602, 16'd47009, 16'd16187, 16'd54693, 16'd1873, 16'd28226, 16'd46590, 16'd52964, 16'd23289, 16'd17402, 16'd24319, 16'd30709, 16'd17400, 16'd51580, 16'd21396, 16'd63068});
	test_expansion(128'h25654ed10b8d963215f01eddc7cf9f53, {16'd42307, 16'd1103, 16'd23291, 16'd15358, 16'd6849, 16'd21744, 16'd7022, 16'd29917, 16'd15912, 16'd61465, 16'd36676, 16'd17206, 16'd47761, 16'd65263, 16'd29981, 16'd56140, 16'd55917, 16'd19772, 16'd2239, 16'd12297, 16'd12695, 16'd1785, 16'd33816, 16'd19311, 16'd13386, 16'd60766});
	test_expansion(128'h726f0c04cd2a91f2c8a051964248f6e5, {16'd44441, 16'd53686, 16'd30706, 16'd34076, 16'd6179, 16'd24587, 16'd33170, 16'd21275, 16'd4594, 16'd58687, 16'd1175, 16'd25427, 16'd27982, 16'd28098, 16'd38684, 16'd48795, 16'd11600, 16'd20875, 16'd1733, 16'd55696, 16'd22746, 16'd57403, 16'd56767, 16'd2700, 16'd10462, 16'd55366});
	test_expansion(128'h72e4168ddc8032ccc11d9151356fc123, {16'd4674, 16'd13619, 16'd24027, 16'd39088, 16'd3100, 16'd57932, 16'd30454, 16'd43182, 16'd53658, 16'd60418, 16'd48905, 16'd52236, 16'd13735, 16'd53574, 16'd527, 16'd60609, 16'd45210, 16'd55442, 16'd19371, 16'd36468, 16'd37058, 16'd28795, 16'd20143, 16'd25902, 16'd22034, 16'd15117});
	test_expansion(128'h4dd7b2ea1dd2b2ceaff0bc2a5fdefe96, {16'd35862, 16'd53200, 16'd10886, 16'd47104, 16'd50260, 16'd20808, 16'd596, 16'd12358, 16'd61053, 16'd8306, 16'd64249, 16'd20911, 16'd30832, 16'd46766, 16'd27599, 16'd17900, 16'd42095, 16'd11526, 16'd62247, 16'd11724, 16'd58997, 16'd36617, 16'd21480, 16'd26248, 16'd4641, 16'd50630});
	test_expansion(128'h0f189bd83fcb1a29e95aff6bdbb81261, {16'd32176, 16'd65459, 16'd44829, 16'd22270, 16'd64382, 16'd53544, 16'd56233, 16'd3172, 16'd944, 16'd58761, 16'd23213, 16'd60611, 16'd16154, 16'd22893, 16'd42707, 16'd37629, 16'd19673, 16'd36702, 16'd2333, 16'd27546, 16'd54210, 16'd8731, 16'd42126, 16'd23777, 16'd36550, 16'd4014});
	test_expansion(128'hedf9dab3a0f18a805e6c756f9ecc2e7d, {16'd52975, 16'd36885, 16'd41355, 16'd36197, 16'd30737, 16'd24824, 16'd56077, 16'd53343, 16'd28780, 16'd46486, 16'd11717, 16'd26481, 16'd63885, 16'd8975, 16'd20523, 16'd10107, 16'd17400, 16'd23797, 16'd30899, 16'd26519, 16'd37966, 16'd52017, 16'd18987, 16'd15629, 16'd58860, 16'd12728});
	test_expansion(128'h44ec9cc9e8dd15b47b599965e56ab590, {16'd3032, 16'd14063, 16'd13776, 16'd6760, 16'd30495, 16'd52707, 16'd4726, 16'd46649, 16'd1257, 16'd31861, 16'd62962, 16'd33110, 16'd32055, 16'd46720, 16'd42152, 16'd35450, 16'd5555, 16'd11155, 16'd48470, 16'd37901, 16'd4476, 16'd34082, 16'd33062, 16'd11346, 16'd60394, 16'd25459});
	test_expansion(128'h6d00fcd40236de970be5cafde707ca04, {16'd48410, 16'd57246, 16'd25978, 16'd13138, 16'd16703, 16'd6225, 16'd27881, 16'd408, 16'd62705, 16'd33936, 16'd43487, 16'd4919, 16'd59704, 16'd12453, 16'd47702, 16'd10683, 16'd46879, 16'd36749, 16'd2754, 16'd65306, 16'd60650, 16'd16612, 16'd1696, 16'd64561, 16'd53990, 16'd34437});
	test_expansion(128'hddb00b81c5b1ee59eb77934b36666f23, {16'd27658, 16'd27504, 16'd42243, 16'd54487, 16'd30753, 16'd37036, 16'd21429, 16'd19101, 16'd16670, 16'd19406, 16'd22069, 16'd5526, 16'd39578, 16'd30635, 16'd38824, 16'd61402, 16'd7746, 16'd47822, 16'd7211, 16'd30386, 16'd9605, 16'd23096, 16'd56736, 16'd13964, 16'd30263, 16'd30953});
	test_expansion(128'h3ebefb8dac60cb80c9c03c3627768218, {16'd29418, 16'd47045, 16'd22560, 16'd63143, 16'd56935, 16'd46264, 16'd43751, 16'd41523, 16'd27903, 16'd63178, 16'd60080, 16'd61742, 16'd5845, 16'd29933, 16'd14505, 16'd58792, 16'd44150, 16'd2070, 16'd54773, 16'd28563, 16'd61528, 16'd57484, 16'd60957, 16'd53670, 16'd63074, 16'd35220});
	test_expansion(128'hb4f50f8108d62b218721d2eb8dd2fc46, {16'd54849, 16'd29318, 16'd7496, 16'd28513, 16'd3502, 16'd14731, 16'd26083, 16'd48029, 16'd46471, 16'd41192, 16'd24224, 16'd52847, 16'd6740, 16'd49500, 16'd42247, 16'd686, 16'd51917, 16'd47907, 16'd42026, 16'd44941, 16'd4147, 16'd31044, 16'd25411, 16'd31998, 16'd55668, 16'd2924});
	test_expansion(128'h68a3f029833cb8f4c80dca7f7a117a35, {16'd51492, 16'd26076, 16'd31618, 16'd314, 16'd65124, 16'd61553, 16'd22903, 16'd26396, 16'd24816, 16'd4694, 16'd49868, 16'd7377, 16'd35939, 16'd7114, 16'd60812, 16'd26377, 16'd22608, 16'd10110, 16'd62205, 16'd61715, 16'd23658, 16'd42244, 16'd18138, 16'd59139, 16'd7715, 16'd1118});
	test_expansion(128'he1b1ba586e92a176518035d0ab246f0e, {16'd61168, 16'd13022, 16'd28802, 16'd33413, 16'd43900, 16'd351, 16'd32131, 16'd48560, 16'd49008, 16'd39315, 16'd37683, 16'd62587, 16'd56325, 16'd36419, 16'd59867, 16'd30921, 16'd61054, 16'd27642, 16'd3007, 16'd15984, 16'd54438, 16'd7784, 16'd21904, 16'd52480, 16'd45001, 16'd4675});
	test_expansion(128'h788bbaae00faafb7b16fc92539c3edc5, {16'd2241, 16'd27860, 16'd51877, 16'd10126, 16'd3907, 16'd22521, 16'd39981, 16'd12066, 16'd9607, 16'd2279, 16'd2084, 16'd56995, 16'd29752, 16'd34078, 16'd7497, 16'd24579, 16'd27850, 16'd21680, 16'd26718, 16'd24196, 16'd9494, 16'd52366, 16'd20529, 16'd65494, 16'd45494, 16'd7070});
	test_expansion(128'he31a66eba0796e1215e9c9fea60d0b62, {16'd193, 16'd48253, 16'd48598, 16'd61908, 16'd9058, 16'd29166, 16'd12235, 16'd28110, 16'd19693, 16'd24839, 16'd54862, 16'd59694, 16'd33798, 16'd14270, 16'd13847, 16'd33932, 16'd44362, 16'd55079, 16'd5813, 16'd2999, 16'd55694, 16'd28417, 16'd57469, 16'd2006, 16'd36209, 16'd10601});
	test_expansion(128'h7e054e8601e32fb6f2f33a57814dd14e, {16'd34480, 16'd38873, 16'd39738, 16'd31314, 16'd5202, 16'd10092, 16'd14811, 16'd2795, 16'd8319, 16'd64131, 16'd43481, 16'd2236, 16'd40690, 16'd51141, 16'd22035, 16'd37250, 16'd11015, 16'd12564, 16'd47813, 16'd52680, 16'd36718, 16'd9409, 16'd65241, 16'd45245, 16'd40768, 16'd15264});
	test_expansion(128'h8716ad28ab4b73f9f6759d204d167496, {16'd48852, 16'd60570, 16'd8155, 16'd25492, 16'd5744, 16'd18168, 16'd4281, 16'd10503, 16'd9003, 16'd16266, 16'd45088, 16'd44820, 16'd6788, 16'd10640, 16'd26021, 16'd38156, 16'd22494, 16'd8300, 16'd32253, 16'd54596, 16'd4383, 16'd32348, 16'd50657, 16'd52402, 16'd23965, 16'd28145});
	test_expansion(128'h050ba61f13a6b0bef0274ca6331fa039, {16'd20073, 16'd14358, 16'd64545, 16'd13601, 16'd56758, 16'd60185, 16'd20203, 16'd49857, 16'd10603, 16'd1483, 16'd32674, 16'd46792, 16'd690, 16'd59287, 16'd50762, 16'd26718, 16'd57257, 16'd12788, 16'd28297, 16'd9755, 16'd37100, 16'd61187, 16'd35885, 16'd34755, 16'd63912, 16'd12306});
	test_expansion(128'h04886640077abd4567983e40c4696969, {16'd51963, 16'd56886, 16'd54777, 16'd55217, 16'd16111, 16'd23811, 16'd62087, 16'd26807, 16'd7160, 16'd37943, 16'd62886, 16'd8823, 16'd35844, 16'd40018, 16'd7160, 16'd55796, 16'd36922, 16'd63559, 16'd4597, 16'd25399, 16'd51405, 16'd57026, 16'd63213, 16'd43866, 16'd3081, 16'd9040});
	test_expansion(128'h6f884a74ee9e4e0877849a331392e8bf, {16'd31211, 16'd37475, 16'd36204, 16'd62841, 16'd11398, 16'd27103, 16'd1318, 16'd61469, 16'd40293, 16'd755, 16'd39733, 16'd58975, 16'd46938, 16'd37365, 16'd4191, 16'd17158, 16'd2957, 16'd42634, 16'd57921, 16'd40639, 16'd39152, 16'd60151, 16'd18863, 16'd2203, 16'd46525, 16'd37429});
	test_expansion(128'h21d3f09037127ea08da2bbb7d1bc04fd, {16'd25272, 16'd9282, 16'd38290, 16'd55888, 16'd8441, 16'd13771, 16'd12617, 16'd50978, 16'd54559, 16'd55747, 16'd38498, 16'd63356, 16'd50159, 16'd38346, 16'd18558, 16'd38953, 16'd39033, 16'd6829, 16'd2563, 16'd60024, 16'd55485, 16'd1239, 16'd35252, 16'd57170, 16'd38744, 16'd61327});
	test_expansion(128'he0e9918eb03ee1972c5a16d9c9123a31, {16'd3045, 16'd3223, 16'd63168, 16'd37979, 16'd51480, 16'd24968, 16'd34854, 16'd60530, 16'd61014, 16'd53054, 16'd29005, 16'd47543, 16'd3543, 16'd27569, 16'd7356, 16'd47167, 16'd45187, 16'd3679, 16'd9897, 16'd62594, 16'd40864, 16'd9025, 16'd38665, 16'd31981, 16'd22312, 16'd7546});
	test_expansion(128'hfd4d03fdf8179c67e5da7bece93cda13, {16'd18556, 16'd45807, 16'd20367, 16'd3185, 16'd17130, 16'd54153, 16'd65469, 16'd53790, 16'd38237, 16'd31709, 16'd50563, 16'd7666, 16'd46052, 16'd27826, 16'd13090, 16'd58035, 16'd9992, 16'd31614, 16'd39692, 16'd27645, 16'd51734, 16'd12940, 16'd32553, 16'd56467, 16'd33952, 16'd51277});
	test_expansion(128'h523a6d0c427c57d230d658e07314b2ad, {16'd20620, 16'd51897, 16'd35380, 16'd29071, 16'd435, 16'd7004, 16'd8886, 16'd26827, 16'd20136, 16'd17154, 16'd212, 16'd10122, 16'd35294, 16'd5976, 16'd63183, 16'd32035, 16'd20286, 16'd65314, 16'd61449, 16'd64815, 16'd45144, 16'd34675, 16'd41422, 16'd61471, 16'd57014, 16'd27698});
	test_expansion(128'h22a967af0d1d3e65b2c0b754dc49c94a, {16'd58518, 16'd24325, 16'd7504, 16'd56585, 16'd10596, 16'd45420, 16'd16776, 16'd42906, 16'd7323, 16'd28798, 16'd26660, 16'd9246, 16'd801, 16'd1082, 16'd16789, 16'd13502, 16'd40848, 16'd7158, 16'd43894, 16'd47998, 16'd21621, 16'd65277, 16'd32822, 16'd26299, 16'd50069, 16'd40191});
	test_expansion(128'h6f8fbd9af478e48d8737903e134f7faf, {16'd40224, 16'd22451, 16'd48515, 16'd62820, 16'd39264, 16'd29785, 16'd48461, 16'd943, 16'd1598, 16'd36794, 16'd55036, 16'd3177, 16'd44922, 16'd56962, 16'd44965, 16'd28493, 16'd10821, 16'd4620, 16'd3596, 16'd19605, 16'd40164, 16'd7689, 16'd210, 16'd64689, 16'd3150, 16'd18754});
	test_expansion(128'hb042dd2ffd6c24b5eec0bd35880d3380, {16'd41379, 16'd48910, 16'd44493, 16'd50100, 16'd65218, 16'd43265, 16'd22427, 16'd54927, 16'd37460, 16'd20177, 16'd48940, 16'd59022, 16'd49213, 16'd25160, 16'd5125, 16'd63094, 16'd51185, 16'd38483, 16'd22827, 16'd14283, 16'd24374, 16'd53829, 16'd11114, 16'd23745, 16'd64871, 16'd58537});
	test_expansion(128'h5b142cf36f686699bf9e13fea3b62396, {16'd27437, 16'd58038, 16'd38957, 16'd57277, 16'd22406, 16'd39565, 16'd17099, 16'd62754, 16'd40335, 16'd5830, 16'd31899, 16'd30667, 16'd18677, 16'd34294, 16'd32253, 16'd62923, 16'd64903, 16'd23439, 16'd9703, 16'd56869, 16'd42448, 16'd9623, 16'd20315, 16'd11331, 16'd63053, 16'd21006});
	test_expansion(128'h3f875f96b28935b2128b972a9ea06e34, {16'd15596, 16'd30879, 16'd30461, 16'd48817, 16'd47772, 16'd30837, 16'd63151, 16'd39182, 16'd37442, 16'd3354, 16'd1482, 16'd10078, 16'd43124, 16'd49170, 16'd45807, 16'd34734, 16'd28138, 16'd23625, 16'd26195, 16'd11922, 16'd63129, 16'd60333, 16'd18532, 16'd31844, 16'd16417, 16'd44323});
	test_expansion(128'h27cd60c82973e59feb41ea36f29b4d3c, {16'd53232, 16'd45879, 16'd53384, 16'd49059, 16'd25318, 16'd43737, 16'd12082, 16'd47199, 16'd14516, 16'd43772, 16'd56610, 16'd21135, 16'd18240, 16'd11685, 16'd59764, 16'd55089, 16'd8153, 16'd52801, 16'd3058, 16'd36818, 16'd57136, 16'd52320, 16'd57342, 16'd29161, 16'd19419, 16'd3655});
	test_expansion(128'h7357f6c166f74dec0415a95e7419cc47, {16'd6336, 16'd51628, 16'd35292, 16'd27824, 16'd33035, 16'd11237, 16'd36084, 16'd41905, 16'd14158, 16'd15923, 16'd17305, 16'd28416, 16'd30077, 16'd24247, 16'd65144, 16'd49733, 16'd48008, 16'd91, 16'd64202, 16'd1957, 16'd54483, 16'd48184, 16'd34375, 16'd4895, 16'd49400, 16'd429});
	test_expansion(128'h0dab930511b85097058017502bfff1d9, {16'd55157, 16'd22844, 16'd25188, 16'd16188, 16'd41055, 16'd45851, 16'd27296, 16'd52258, 16'd2012, 16'd14370, 16'd8346, 16'd34602, 16'd11771, 16'd54684, 16'd6668, 16'd201, 16'd44051, 16'd716, 16'd56100, 16'd36383, 16'd44026, 16'd38023, 16'd11224, 16'd26766, 16'd11773, 16'd26538});
	test_expansion(128'he10317f92bf92b73836f389fb28248ed, {16'd1566, 16'd53512, 16'd6148, 16'd61630, 16'd29072, 16'd35688, 16'd6307, 16'd21873, 16'd12045, 16'd35593, 16'd34317, 16'd21987, 16'd54125, 16'd4035, 16'd6530, 16'd50786, 16'd21376, 16'd51655, 16'd50855, 16'd41168, 16'd15915, 16'd44393, 16'd41949, 16'd45149, 16'd60842, 16'd8366});
	test_expansion(128'h1806c319041133d9f99177c6506225f2, {16'd3358, 16'd57368, 16'd11053, 16'd52786, 16'd40840, 16'd48084, 16'd34709, 16'd19383, 16'd22469, 16'd26558, 16'd7370, 16'd40630, 16'd14876, 16'd1594, 16'd12991, 16'd12369, 16'd42914, 16'd32902, 16'd14646, 16'd10470, 16'd39354, 16'd27214, 16'd14624, 16'd4999, 16'd20960, 16'd32563});
	test_expansion(128'h4072e6516c8dae296b15dbf75aade512, {16'd34569, 16'd32672, 16'd40427, 16'd23080, 16'd26719, 16'd36332, 16'd45473, 16'd56539, 16'd47922, 16'd44794, 16'd2238, 16'd49566, 16'd59356, 16'd13217, 16'd30542, 16'd46022, 16'd20270, 16'd279, 16'd54033, 16'd53078, 16'd37018, 16'd19670, 16'd22000, 16'd13352, 16'd35903, 16'd56998});
	test_expansion(128'h9c0c3b47c2ada59c89529be54d7591a2, {16'd10995, 16'd20523, 16'd29798, 16'd27732, 16'd7596, 16'd59729, 16'd64904, 16'd53408, 16'd23693, 16'd4442, 16'd39610, 16'd57395, 16'd25172, 16'd8733, 16'd3286, 16'd34330, 16'd2138, 16'd49237, 16'd28998, 16'd29845, 16'd12923, 16'd31111, 16'd64733, 16'd13775, 16'd15755, 16'd25166});
	test_expansion(128'h4e4405c2e772791c38375d54c0833a73, {16'd28828, 16'd7686, 16'd60330, 16'd20494, 16'd10414, 16'd32969, 16'd54990, 16'd25348, 16'd32836, 16'd9554, 16'd62930, 16'd50486, 16'd40823, 16'd6517, 16'd1653, 16'd32010, 16'd3452, 16'd56896, 16'd49006, 16'd2426, 16'd18650, 16'd12798, 16'd42876, 16'd32084, 16'd16558, 16'd4936});
	test_expansion(128'hc42f84eb082f8f61380aa2ba4f5c4fff, {16'd30908, 16'd32734, 16'd52104, 16'd26786, 16'd60012, 16'd30763, 16'd57893, 16'd56352, 16'd6245, 16'd1865, 16'd24768, 16'd51000, 16'd51425, 16'd1452, 16'd5911, 16'd10475, 16'd12966, 16'd9645, 16'd2855, 16'd22015, 16'd32695, 16'd29255, 16'd34387, 16'd942, 16'd6673, 16'd1867});
	test_expansion(128'h02daeb33c3ac3d0ed09cb72777a786b7, {16'd17346, 16'd7819, 16'd34918, 16'd40309, 16'd40311, 16'd10954, 16'd53078, 16'd56281, 16'd60136, 16'd42343, 16'd18350, 16'd30925, 16'd33381, 16'd32787, 16'd1948, 16'd14480, 16'd54105, 16'd6503, 16'd29033, 16'd28112, 16'd18212, 16'd23228, 16'd48305, 16'd46810, 16'd56512, 16'd35142});
	test_expansion(128'hfc643630a6d897e16cc5006e54d4586f, {16'd48914, 16'd54368, 16'd10447, 16'd42486, 16'd37339, 16'd18010, 16'd28056, 16'd27780, 16'd6390, 16'd10233, 16'd10157, 16'd57830, 16'd39995, 16'd27286, 16'd64658, 16'd62995, 16'd5750, 16'd61622, 16'd43441, 16'd39293, 16'd8503, 16'd53437, 16'd26259, 16'd3471, 16'd63396, 16'd24977});
	test_expansion(128'h49f04f6177ea4cfaba8115f2d3b95c63, {16'd728, 16'd40667, 16'd11127, 16'd14836, 16'd16737, 16'd16106, 16'd30574, 16'd4240, 16'd27131, 16'd41629, 16'd22681, 16'd11343, 16'd15515, 16'd5137, 16'd39612, 16'd11189, 16'd30338, 16'd63746, 16'd6951, 16'd64505, 16'd39425, 16'd21923, 16'd36526, 16'd61097, 16'd59878, 16'd5074});
	test_expansion(128'hebd737b099718e688bf54306ab24cce9, {16'd34845, 16'd23389, 16'd41925, 16'd21628, 16'd21025, 16'd65398, 16'd8179, 16'd19405, 16'd23712, 16'd33266, 16'd49251, 16'd37492, 16'd60790, 16'd33342, 16'd60101, 16'd20489, 16'd29690, 16'd56850, 16'd20722, 16'd11063, 16'd16096, 16'd32967, 16'd55271, 16'd48659, 16'd35996, 16'd64916});
	test_expansion(128'hadd036bc8bb5ef0979a02bd74c33c4b0, {16'd25205, 16'd44398, 16'd38453, 16'd44164, 16'd43336, 16'd28201, 16'd20523, 16'd26790, 16'd52938, 16'd58626, 16'd775, 16'd30886, 16'd28734, 16'd21765, 16'd44158, 16'd19672, 16'd6438, 16'd10287, 16'd51244, 16'd58271, 16'd50853, 16'd55404, 16'd57356, 16'd64555, 16'd22234, 16'd25935});
	test_expansion(128'h717b5be658c4225bf28b484b4809289b, {16'd29002, 16'd25317, 16'd36430, 16'd53801, 16'd16106, 16'd23127, 16'd17049, 16'd10260, 16'd13506, 16'd6465, 16'd18840, 16'd800, 16'd50184, 16'd23955, 16'd16814, 16'd26611, 16'd39570, 16'd23572, 16'd40500, 16'd20078, 16'd4481, 16'd33090, 16'd35031, 16'd61326, 16'd47105, 16'd30616});
	test_expansion(128'h3d5f4c00a588efcaa97eaee9aa29b2e1, {16'd13856, 16'd65510, 16'd51773, 16'd56669, 16'd46498, 16'd10849, 16'd50941, 16'd20824, 16'd30319, 16'd54573, 16'd24274, 16'd14954, 16'd50896, 16'd16161, 16'd60134, 16'd12233, 16'd34086, 16'd53086, 16'd51065, 16'd50375, 16'd53327, 16'd53521, 16'd40847, 16'd51181, 16'd64419, 16'd3903});
	test_expansion(128'h19c51c41bc7d67a61f124fba8a690176, {16'd55514, 16'd16684, 16'd32063, 16'd55058, 16'd12591, 16'd10857, 16'd13424, 16'd30589, 16'd63756, 16'd16519, 16'd9603, 16'd31582, 16'd13612, 16'd14436, 16'd20078, 16'd39180, 16'd12377, 16'd49110, 16'd2098, 16'd47709, 16'd50845, 16'd25142, 16'd57307, 16'd45525, 16'd33600, 16'd37528});
	test_expansion(128'h4fa87f982b3c4033784cae937c2f7fe8, {16'd11527, 16'd50938, 16'd6001, 16'd9489, 16'd22791, 16'd57591, 16'd29546, 16'd30483, 16'd22200, 16'd28653, 16'd38284, 16'd49601, 16'd64364, 16'd1825, 16'd7060, 16'd11883, 16'd52680, 16'd42247, 16'd13960, 16'd59558, 16'd64004, 16'd38590, 16'd37971, 16'd41231, 16'd11143, 16'd20092});
	test_expansion(128'h5aeaccc734d53c7f7b2851f2ef554af5, {16'd58078, 16'd63358, 16'd57133, 16'd54891, 16'd35001, 16'd45385, 16'd60863, 16'd51625, 16'd21571, 16'd5068, 16'd39774, 16'd58222, 16'd52343, 16'd19734, 16'd52867, 16'd19730, 16'd48240, 16'd26327, 16'd57799, 16'd64404, 16'd27007, 16'd53315, 16'd2164, 16'd61326, 16'd7777, 16'd51014});
	test_expansion(128'h876c273d3a25f9ecf06ab5a5231f80eb, {16'd64161, 16'd47535, 16'd55046, 16'd53770, 16'd41798, 16'd45654, 16'd29142, 16'd52788, 16'd38950, 16'd5361, 16'd47028, 16'd25363, 16'd62619, 16'd50096, 16'd61055, 16'd42989, 16'd60633, 16'd46959, 16'd45836, 16'd44879, 16'd3969, 16'd63479, 16'd63501, 16'd12143, 16'd44818, 16'd16593});
	test_expansion(128'hb034b2d39f51f5812f6cc216ce858301, {16'd51854, 16'd11452, 16'd30012, 16'd49842, 16'd56234, 16'd63626, 16'd3424, 16'd57759, 16'd31669, 16'd48240, 16'd43479, 16'd48554, 16'd32087, 16'd19598, 16'd14606, 16'd25179, 16'd29857, 16'd20758, 16'd64267, 16'd63608, 16'd30046, 16'd32195, 16'd63718, 16'd3487, 16'd15228, 16'd49753});
	test_expansion(128'h86c80f197fe2061e727aba28e378fed8, {16'd47478, 16'd19914, 16'd13043, 16'd19972, 16'd29962, 16'd63619, 16'd25320, 16'd50137, 16'd50754, 16'd41738, 16'd31071, 16'd49750, 16'd63888, 16'd1166, 16'd39156, 16'd22559, 16'd55558, 16'd61741, 16'd60392, 16'd59387, 16'd19777, 16'd39911, 16'd64796, 16'd41741, 16'd46115, 16'd61355});
	test_expansion(128'h4fe7ef900d61185173236e34c54ddb49, {16'd45299, 16'd8836, 16'd60998, 16'd30864, 16'd50240, 16'd62659, 16'd35314, 16'd8503, 16'd18350, 16'd41974, 16'd53277, 16'd39899, 16'd1455, 16'd53259, 16'd5164, 16'd21964, 16'd659, 16'd13907, 16'd19732, 16'd10253, 16'd44780, 16'd61598, 16'd59034, 16'd29331, 16'd8696, 16'd45140});
	test_expansion(128'hd01b09e012e3a0383cc58e8837c5b9cc, {16'd10988, 16'd65116, 16'd20887, 16'd1024, 16'd42390, 16'd58395, 16'd58118, 16'd49927, 16'd38702, 16'd27616, 16'd10309, 16'd7817, 16'd26854, 16'd25472, 16'd23602, 16'd3223, 16'd25529, 16'd3831, 16'd22941, 16'd12679, 16'd55632, 16'd13869, 16'd48224, 16'd62954, 16'd61108, 16'd47358});
	test_expansion(128'hdceda91086c343dca51aa637a81cf9fc, {16'd37439, 16'd62009, 16'd62987, 16'd23520, 16'd16764, 16'd9617, 16'd46731, 16'd28810, 16'd24823, 16'd61160, 16'd27126, 16'd65288, 16'd7063, 16'd14634, 16'd40980, 16'd16337, 16'd12774, 16'd28746, 16'd41015, 16'd50486, 16'd41120, 16'd51559, 16'd32927, 16'd52472, 16'd64545, 16'd49191});
	test_expansion(128'h8ff2510ef811d81d7ae9d3c208e9c766, {16'd46073, 16'd48615, 16'd29382, 16'd29739, 16'd59542, 16'd47392, 16'd17672, 16'd28291, 16'd24799, 16'd43972, 16'd55353, 16'd30922, 16'd25746, 16'd44513, 16'd58843, 16'd22691, 16'd39938, 16'd3619, 16'd46217, 16'd12403, 16'd34027, 16'd44725, 16'd52828, 16'd54222, 16'd42209, 16'd11607});
	test_expansion(128'h0d1d79d01c5e0aa922c4972b07bd6c1b, {16'd62333, 16'd15560, 16'd46435, 16'd42445, 16'd19587, 16'd45477, 16'd52732, 16'd13041, 16'd62767, 16'd21876, 16'd45334, 16'd18628, 16'd25559, 16'd44241, 16'd30919, 16'd41925, 16'd36215, 16'd8535, 16'd7485, 16'd42128, 16'd13869, 16'd920, 16'd4985, 16'd62065, 16'd43757, 16'd56143});
	test_expansion(128'hb090660e86df5883418c7fa2eec43a3f, {16'd18033, 16'd48701, 16'd12388, 16'd13303, 16'd55873, 16'd36656, 16'd32384, 16'd28253, 16'd47592, 16'd51071, 16'd37407, 16'd32848, 16'd21173, 16'd19805, 16'd14822, 16'd24100, 16'd22056, 16'd64327, 16'd35047, 16'd42875, 16'd6007, 16'd61352, 16'd28553, 16'd36011, 16'd32010, 16'd24485});
	test_expansion(128'hb9024a0a233d11da4d00703b8f4db68f, {16'd60099, 16'd47474, 16'd4936, 16'd22470, 16'd23667, 16'd63113, 16'd12730, 16'd16133, 16'd29598, 16'd50342, 16'd44963, 16'd54, 16'd13935, 16'd10211, 16'd9471, 16'd36735, 16'd57492, 16'd14446, 16'd24137, 16'd51905, 16'd20134, 16'd3358, 16'd47193, 16'd35765, 16'd60319, 16'd42973});
	test_expansion(128'h8b374dda90f24065240e3c1a7bbe9a32, {16'd48060, 16'd55577, 16'd17539, 16'd1766, 16'd20563, 16'd51647, 16'd21220, 16'd42627, 16'd53833, 16'd16220, 16'd16257, 16'd10365, 16'd15161, 16'd17459, 16'd7297, 16'd3937, 16'd6702, 16'd51902, 16'd11583, 16'd27860, 16'd51931, 16'd43668, 16'd45062, 16'd62635, 16'd61403, 16'd57633});
	test_expansion(128'hc23f55df7251f5cb1fde3e4a8306cd3a, {16'd61189, 16'd29835, 16'd2211, 16'd42183, 16'd12607, 16'd46690, 16'd26402, 16'd41413, 16'd81, 16'd26367, 16'd33684, 16'd14170, 16'd47800, 16'd17347, 16'd16557, 16'd37642, 16'd17697, 16'd56186, 16'd36304, 16'd11225, 16'd18087, 16'd64605, 16'd49070, 16'd37180, 16'd33989, 16'd50060});
	test_expansion(128'h3042433880850030c87130399c5456b2, {16'd806, 16'd37878, 16'd19226, 16'd51396, 16'd50255, 16'd63742, 16'd63754, 16'd55710, 16'd13264, 16'd44260, 16'd23687, 16'd43391, 16'd31221, 16'd54566, 16'd10818, 16'd34068, 16'd59780, 16'd49329, 16'd7989, 16'd31960, 16'd42850, 16'd15604, 16'd5731, 16'd23229, 16'd2128, 16'd18762});
	test_expansion(128'h3c1bc70e77659a11c732bb871c6862d8, {16'd59100, 16'd50567, 16'd65515, 16'd44850, 16'd35280, 16'd59126, 16'd29204, 16'd5094, 16'd1088, 16'd19610, 16'd22109, 16'd1402, 16'd1417, 16'd53867, 16'd58998, 16'd44058, 16'd24589, 16'd23634, 16'd1510, 16'd32684, 16'd9373, 16'd61627, 16'd35444, 16'd142, 16'd51556, 16'd31817});
	test_expansion(128'h38885bb263675da473af77f3cc039ec7, {16'd9396, 16'd22430, 16'd65229, 16'd5622, 16'd56018, 16'd52487, 16'd63663, 16'd38424, 16'd11930, 16'd3498, 16'd47836, 16'd1062, 16'd27105, 16'd11722, 16'd20479, 16'd60537, 16'd4804, 16'd49632, 16'd40635, 16'd43985, 16'd57616, 16'd30545, 16'd44583, 16'd22178, 16'd8760, 16'd29309});
	test_expansion(128'h4ed5f274ee1c8b4dd38328c76fb98783, {16'd43709, 16'd31975, 16'd32201, 16'd23583, 16'd17298, 16'd20382, 16'd62308, 16'd135, 16'd60968, 16'd32792, 16'd30855, 16'd42562, 16'd44700, 16'd1196, 16'd4859, 16'd31977, 16'd59969, 16'd5038, 16'd973, 16'd47772, 16'd16143, 16'd26518, 16'd20170, 16'd52518, 16'd21699, 16'd39246});
	test_expansion(128'h61575d5b834b242f606262eee8d7add3, {16'd24949, 16'd770, 16'd20570, 16'd62805, 16'd26099, 16'd11771, 16'd6524, 16'd3792, 16'd63106, 16'd52965, 16'd10622, 16'd28622, 16'd52054, 16'd5640, 16'd12500, 16'd10587, 16'd29151, 16'd59080, 16'd52442, 16'd52599, 16'd55972, 16'd36536, 16'd16908, 16'd9184, 16'd2083, 16'd12829});
	test_expansion(128'h2419eaa89704c71ab0375e86efe0e023, {16'd53440, 16'd35393, 16'd24898, 16'd30792, 16'd14213, 16'd25868, 16'd29631, 16'd33928, 16'd57328, 16'd43375, 16'd36563, 16'd9634, 16'd1899, 16'd6280, 16'd45321, 16'd29700, 16'd11974, 16'd44631, 16'd59659, 16'd5553, 16'd20316, 16'd10780, 16'd5006, 16'd35836, 16'd43005, 16'd18303});
	test_expansion(128'h2dc880f41808b34e9e89e13785f7105e, {16'd42168, 16'd18208, 16'd6943, 16'd21602, 16'd55776, 16'd33200, 16'd44124, 16'd23033, 16'd27924, 16'd19880, 16'd27010, 16'd16129, 16'd35453, 16'd35002, 16'd12087, 16'd56265, 16'd19295, 16'd32257, 16'd32010, 16'd32068, 16'd22921, 16'd18178, 16'd52594, 16'd50167, 16'd4108, 16'd54421});
	test_expansion(128'h70b3d91d28834121e66466b3dd1ac831, {16'd14213, 16'd43039, 16'd42952, 16'd16347, 16'd53451, 16'd2497, 16'd37865, 16'd33946, 16'd37779, 16'd62287, 16'd7544, 16'd39128, 16'd49430, 16'd51687, 16'd3312, 16'd56526, 16'd44988, 16'd61693, 16'd20210, 16'd4518, 16'd6620, 16'd36130, 16'd12965, 16'd25949, 16'd5720, 16'd22541});
	test_expansion(128'hd733b7028e4edfc27ff6b91c37a58fb1, {16'd41114, 16'd46957, 16'd43329, 16'd5178, 16'd51092, 16'd17058, 16'd38524, 16'd43943, 16'd46609, 16'd52155, 16'd27980, 16'd846, 16'd14474, 16'd27956, 16'd20627, 16'd17737, 16'd50127, 16'd18758, 16'd15355, 16'd61551, 16'd31216, 16'd15940, 16'd64983, 16'd54450, 16'd1553, 16'd39110});
	test_expansion(128'h17d9cbb939ec7aca4993bf1ca070c7cf, {16'd63537, 16'd53388, 16'd45569, 16'd64957, 16'd35546, 16'd21846, 16'd8901, 16'd798, 16'd17780, 16'd63294, 16'd34123, 16'd57064, 16'd47999, 16'd44929, 16'd62651, 16'd47341, 16'd6178, 16'd18595, 16'd31648, 16'd31476, 16'd24683, 16'd42821, 16'd39434, 16'd49896, 16'd6607, 16'd32170});
	test_expansion(128'hd01efbbea1e4f4d0958d0bea4dd6b6e7, {16'd42568, 16'd13102, 16'd17562, 16'd14070, 16'd367, 16'd19714, 16'd5688, 16'd39798, 16'd64491, 16'd55355, 16'd36980, 16'd45149, 16'd57053, 16'd2938, 16'd60332, 16'd27964, 16'd7895, 16'd3691, 16'd63682, 16'd12191, 16'd46557, 16'd2122, 16'd47272, 16'd22358, 16'd37979, 16'd22640});
	test_expansion(128'hdee9396f372adeabf5ea6621217b2bc0, {16'd28294, 16'd59474, 16'd8627, 16'd12572, 16'd8252, 16'd28706, 16'd53698, 16'd49619, 16'd54045, 16'd46517, 16'd34636, 16'd55362, 16'd59953, 16'd35859, 16'd21270, 16'd17011, 16'd37938, 16'd53511, 16'd61695, 16'd12217, 16'd17408, 16'd21320, 16'd9970, 16'd47214, 16'd55849, 16'd12003});
	test_expansion(128'h74abd4508605d8bc23db69aae283005c, {16'd49156, 16'd48988, 16'd47774, 16'd36635, 16'd6334, 16'd12009, 16'd51623, 16'd54726, 16'd16418, 16'd4297, 16'd6462, 16'd50038, 16'd18193, 16'd36413, 16'd12309, 16'd49167, 16'd49508, 16'd56771, 16'd17552, 16'd13483, 16'd42567, 16'd52919, 16'd6428, 16'd15770, 16'd11581, 16'd1262});
	test_expansion(128'h3fadcbeb6f72de3c7a550729c12cd1b3, {16'd29562, 16'd61770, 16'd60268, 16'd12984, 16'd6375, 16'd24170, 16'd57023, 16'd63488, 16'd48112, 16'd10154, 16'd56050, 16'd37549, 16'd21450, 16'd47235, 16'd42569, 16'd658, 16'd19496, 16'd15684, 16'd20163, 16'd49813, 16'd59817, 16'd39376, 16'd36354, 16'd20000, 16'd32350, 16'd31994});
	test_expansion(128'h6a1d57912ada7fc77c8501e1a14bb0a0, {16'd35378, 16'd2568, 16'd27428, 16'd26170, 16'd3797, 16'd47003, 16'd62894, 16'd32182, 16'd26443, 16'd18189, 16'd5551, 16'd30264, 16'd9886, 16'd26329, 16'd48667, 16'd23285, 16'd18032, 16'd41563, 16'd28757, 16'd36297, 16'd62663, 16'd17409, 16'd19825, 16'd4251, 16'd54438, 16'd17201});
	test_expansion(128'hd97739aef9a7df95abc925ffd7cf4a16, {16'd60998, 16'd51907, 16'd46845, 16'd32697, 16'd31055, 16'd15475, 16'd53420, 16'd43123, 16'd64037, 16'd18501, 16'd40729, 16'd54085, 16'd32416, 16'd1425, 16'd50853, 16'd20641, 16'd22505, 16'd59103, 16'd22070, 16'd34288, 16'd15077, 16'd43355, 16'd18250, 16'd46399, 16'd64314, 16'd22000});
	test_expansion(128'hc691d39f335be6890bc259ead597a6f7, {16'd45186, 16'd20867, 16'd3213, 16'd25950, 16'd56637, 16'd54831, 16'd52411, 16'd25641, 16'd60493, 16'd57879, 16'd10733, 16'd42315, 16'd43730, 16'd40147, 16'd23170, 16'd21193, 16'd39592, 16'd38983, 16'd38962, 16'd22584, 16'd47428, 16'd15236, 16'd41529, 16'd63118, 16'd33311, 16'd12156});
	test_expansion(128'h21834e9a56888f62281fd7039dff2204, {16'd5550, 16'd51443, 16'd22029, 16'd47507, 16'd2409, 16'd48962, 16'd9809, 16'd11960, 16'd57494, 16'd52803, 16'd873, 16'd6532, 16'd17391, 16'd48031, 16'd31950, 16'd18118, 16'd11034, 16'd57490, 16'd9004, 16'd8352, 16'd17410, 16'd27596, 16'd13664, 16'd12010, 16'd48551, 16'd51139});
	test_expansion(128'h9e53a98e53e63b1359830ff944722355, {16'd52398, 16'd62767, 16'd52992, 16'd32220, 16'd55361, 16'd62404, 16'd63336, 16'd22286, 16'd9872, 16'd42100, 16'd8322, 16'd40498, 16'd48717, 16'd46184, 16'd40570, 16'd35192, 16'd41778, 16'd54354, 16'd4329, 16'd13337, 16'd56740, 16'd7853, 16'd43875, 16'd23932, 16'd15088, 16'd50069});
	test_expansion(128'hefd76c562f3c5fe6c1a0d7872ae85970, {16'd28069, 16'd1109, 16'd28109, 16'd48093, 16'd32142, 16'd17003, 16'd30744, 16'd33233, 16'd52869, 16'd29856, 16'd39796, 16'd13493, 16'd49395, 16'd63727, 16'd31821, 16'd27976, 16'd19912, 16'd59695, 16'd26688, 16'd32225, 16'd18213, 16'd39764, 16'd59652, 16'd11968, 16'd30628, 16'd42938});
	test_expansion(128'hdc14c0b371598c44f0c3874370e43ba3, {16'd33220, 16'd4469, 16'd22992, 16'd36999, 16'd56801, 16'd22022, 16'd49806, 16'd11466, 16'd44612, 16'd21938, 16'd33234, 16'd49290, 16'd13122, 16'd64558, 16'd55343, 16'd64904, 16'd62921, 16'd55350, 16'd59212, 16'd55452, 16'd53644, 16'd59616, 16'd36496, 16'd5849, 16'd53075, 16'd57289});
	test_expansion(128'ha44da5dfcd19d8780e4e418baa018912, {16'd30253, 16'd40090, 16'd11720, 16'd37325, 16'd7350, 16'd61087, 16'd45794, 16'd22337, 16'd23690, 16'd30776, 16'd43540, 16'd52177, 16'd14946, 16'd59722, 16'd39879, 16'd38530, 16'd13017, 16'd5296, 16'd24162, 16'd16014, 16'd25813, 16'd50030, 16'd5734, 16'd36616, 16'd42177, 16'd34639});
	test_expansion(128'h5a44a469bafe1ae079654e0f63f6e2f6, {16'd54728, 16'd20302, 16'd41635, 16'd65216, 16'd46060, 16'd5964, 16'd43376, 16'd26414, 16'd26387, 16'd21490, 16'd55039, 16'd27053, 16'd266, 16'd29193, 16'd51196, 16'd45573, 16'd47865, 16'd59383, 16'd50725, 16'd44830, 16'd53135, 16'd38928, 16'd8673, 16'd32617, 16'd30084, 16'd46581});
	test_expansion(128'hf52a0deca2519b4fe9d567978a3f9634, {16'd43920, 16'd43958, 16'd46646, 16'd58271, 16'd32135, 16'd39165, 16'd30725, 16'd28068, 16'd38902, 16'd17511, 16'd15078, 16'd54178, 16'd39350, 16'd9777, 16'd41683, 16'd40993, 16'd41031, 16'd7780, 16'd62966, 16'd20134, 16'd35440, 16'd33109, 16'd24929, 16'd57494, 16'd30070, 16'd13506});
	test_expansion(128'hd9461749dc2dfd5f4ed8f391007dbd57, {16'd33961, 16'd20551, 16'd13857, 16'd54244, 16'd25246, 16'd3917, 16'd62465, 16'd13540, 16'd62168, 16'd61437, 16'd1145, 16'd30218, 16'd48176, 16'd22670, 16'd57668, 16'd14758, 16'd32918, 16'd5811, 16'd46036, 16'd35320, 16'd40095, 16'd30270, 16'd17780, 16'd62479, 16'd31762, 16'd52380});
	test_expansion(128'hf7a466ecd5476296cdd3cfae43956142, {16'd576, 16'd17353, 16'd36326, 16'd878, 16'd60994, 16'd25014, 16'd41920, 16'd4105, 16'd30511, 16'd1017, 16'd42803, 16'd42049, 16'd56565, 16'd21363, 16'd42281, 16'd54776, 16'd10969, 16'd29367, 16'd65423, 16'd52864, 16'd52348, 16'd14385, 16'd31831, 16'd57998, 16'd34389, 16'd45840});
	test_expansion(128'h8ea0f79c2386ecaf5315caa1bd750671, {16'd28310, 16'd16363, 16'd22400, 16'd21299, 16'd44241, 16'd59659, 16'd13816, 16'd916, 16'd50709, 16'd6736, 16'd61060, 16'd22857, 16'd34515, 16'd41118, 16'd30089, 16'd58763, 16'd23467, 16'd34676, 16'd61592, 16'd50341, 16'd55411, 16'd35279, 16'd54680, 16'd41999, 16'd60300, 16'd29939});
	test_expansion(128'h863a177f5ec8c63613be5c4e810f201d, {16'd47242, 16'd41788, 16'd50721, 16'd8408, 16'd3728, 16'd48264, 16'd49031, 16'd48785, 16'd47185, 16'd30361, 16'd36486, 16'd21490, 16'd53235, 16'd55855, 16'd42240, 16'd33634, 16'd57088, 16'd8978, 16'd26294, 16'd32011, 16'd64782, 16'd28255, 16'd62898, 16'd24944, 16'd30378, 16'd57160});
	test_expansion(128'h5c4afebd2c992f4b0f4cfdc226e8f4d2, {16'd40011, 16'd63981, 16'd32800, 16'd29730, 16'd3533, 16'd13163, 16'd18967, 16'd27466, 16'd16977, 16'd50856, 16'd27707, 16'd41101, 16'd64256, 16'd26382, 16'd14850, 16'd9931, 16'd56380, 16'd60617, 16'd19623, 16'd25126, 16'd60499, 16'd57072, 16'd25525, 16'd9948, 16'd41514, 16'd24732});
	test_expansion(128'h01102ba830634424e5888f51b7747e5b, {16'd59663, 16'd53875, 16'd16662, 16'd39662, 16'd11195, 16'd24569, 16'd1489, 16'd2940, 16'd59353, 16'd26400, 16'd45088, 16'd53468, 16'd51245, 16'd28686, 16'd64708, 16'd14772, 16'd59051, 16'd57770, 16'd55715, 16'd51408, 16'd61496, 16'd11130, 16'd44244, 16'd64010, 16'd26434, 16'd17803});
	test_expansion(128'h2620ac80f0da5b2f03c1c853cd858a1a, {16'd38347, 16'd8443, 16'd11892, 16'd50406, 16'd50096, 16'd35866, 16'd62954, 16'd2457, 16'd39606, 16'd22133, 16'd57123, 16'd2438, 16'd370, 16'd2665, 16'd28135, 16'd11650, 16'd15327, 16'd49805, 16'd37765, 16'd11167, 16'd62671, 16'd27873, 16'd14106, 16'd7, 16'd15597, 16'd60157});
	test_expansion(128'h5ab295d8da0c30730b5f9628c102da41, {16'd59991, 16'd40722, 16'd25147, 16'd62921, 16'd49178, 16'd1460, 16'd43557, 16'd53726, 16'd23574, 16'd651, 16'd28992, 16'd20139, 16'd60604, 16'd20694, 16'd42281, 16'd35388, 16'd47877, 16'd5346, 16'd49581, 16'd29899, 16'd34979, 16'd34589, 16'd35774, 16'd11945, 16'd41113, 16'd25140});
	test_expansion(128'hf29ac4709210496cc6f0a0af990ed3cb, {16'd53402, 16'd10650, 16'd26049, 16'd17296, 16'd13372, 16'd4323, 16'd30855, 16'd25032, 16'd4532, 16'd24535, 16'd33027, 16'd33140, 16'd10920, 16'd36352, 16'd22384, 16'd48816, 16'd38431, 16'd36277, 16'd16968, 16'd1264, 16'd35517, 16'd63552, 16'd11908, 16'd63182, 16'd38701, 16'd37087});
	test_expansion(128'hdb64fd990e1ee038c2c027b3b011292f, {16'd8223, 16'd41058, 16'd59128, 16'd31683, 16'd61994, 16'd7253, 16'd5949, 16'd5000, 16'd45988, 16'd27367, 16'd256, 16'd60116, 16'd50491, 16'd22898, 16'd25467, 16'd47116, 16'd11909, 16'd52422, 16'd46353, 16'd33292, 16'd4537, 16'd60906, 16'd16799, 16'd44073, 16'd4761, 16'd37484});
	test_expansion(128'h14884c7733a040970e8c2545063ac319, {16'd47509, 16'd21776, 16'd34289, 16'd667, 16'd4054, 16'd23425, 16'd61986, 16'd1056, 16'd37525, 16'd64143, 16'd64105, 16'd59129, 16'd18610, 16'd11599, 16'd63586, 16'd65357, 16'd21738, 16'd25983, 16'd32867, 16'd43541, 16'd47233, 16'd11390, 16'd43593, 16'd47142, 16'd57655, 16'd41699});
	test_expansion(128'h879ab4225fd56f5289ff9cc7871477b9, {16'd31357, 16'd32552, 16'd11625, 16'd24197, 16'd21966, 16'd54753, 16'd34985, 16'd42800, 16'd48822, 16'd6049, 16'd41642, 16'd16127, 16'd1700, 16'd54326, 16'd20075, 16'd16200, 16'd15943, 16'd719, 16'd13011, 16'd18789, 16'd62960, 16'd55890, 16'd477, 16'd60783, 16'd5136, 16'd61787});
	test_expansion(128'ha685abafab81e245f232066b0f5f6208, {16'd57131, 16'd57208, 16'd24844, 16'd4742, 16'd30291, 16'd60584, 16'd39096, 16'd12938, 16'd53044, 16'd30803, 16'd15162, 16'd31872, 16'd3134, 16'd18732, 16'd8812, 16'd42699, 16'd21742, 16'd2733, 16'd17161, 16'd14649, 16'd3132, 16'd34059, 16'd35479, 16'd52936, 16'd15783, 16'd61772});
	test_expansion(128'h91b2f155130cc3e39ce0bed13801c88a, {16'd56139, 16'd2684, 16'd61885, 16'd56949, 16'd60854, 16'd36236, 16'd39309, 16'd5957, 16'd14566, 16'd62754, 16'd4803, 16'd49070, 16'd58278, 16'd8692, 16'd20547, 16'd40519, 16'd19672, 16'd46192, 16'd60437, 16'd10643, 16'd33518, 16'd51972, 16'd5845, 16'd47715, 16'd29836, 16'd56078});
	test_expansion(128'h202384022fd4bb14bf480f90239e3ba7, {16'd4194, 16'd35533, 16'd39825, 16'd6021, 16'd15864, 16'd9538, 16'd8958, 16'd62812, 16'd47793, 16'd25234, 16'd37899, 16'd21808, 16'd63934, 16'd43148, 16'd46613, 16'd31754, 16'd19959, 16'd16100, 16'd38875, 16'd43005, 16'd15172, 16'd22291, 16'd396, 16'd56779, 16'd29744, 16'd47018});
	test_expansion(128'h4c16c379b648a32ae7dfc48893ee0696, {16'd48959, 16'd17829, 16'd28230, 16'd23759, 16'd3084, 16'd45348, 16'd9321, 16'd28289, 16'd44410, 16'd14609, 16'd57767, 16'd22746, 16'd15434, 16'd11605, 16'd32679, 16'd59645, 16'd15148, 16'd2031, 16'd44256, 16'd60878, 16'd60425, 16'd26917, 16'd58277, 16'd45729, 16'd57128, 16'd6426});
	test_expansion(128'hc6fb255ddbbb3124e82ec79bd470bae1, {16'd52578, 16'd14560, 16'd61618, 16'd7203, 16'd18818, 16'd56021, 16'd49953, 16'd38276, 16'd41141, 16'd19283, 16'd42040, 16'd53275, 16'd2924, 16'd46434, 16'd59636, 16'd1301, 16'd23515, 16'd15982, 16'd7098, 16'd18810, 16'd9758, 16'd5705, 16'd31959, 16'd45738, 16'd42213, 16'd70});
	test_expansion(128'h5284684b836070be6b18a08bea9f5b8a, {16'd40973, 16'd35825, 16'd49489, 16'd13791, 16'd60405, 16'd27166, 16'd15318, 16'd33888, 16'd21405, 16'd23231, 16'd25694, 16'd42529, 16'd22577, 16'd46197, 16'd13723, 16'd31405, 16'd3719, 16'd55970, 16'd52789, 16'd370, 16'd51784, 16'd29830, 16'd62765, 16'd32827, 16'd50969, 16'd53846});
	test_expansion(128'hf1720857c2787d4f0902c945b25f46d3, {16'd64774, 16'd32143, 16'd25919, 16'd22568, 16'd63732, 16'd18812, 16'd1981, 16'd11427, 16'd32866, 16'd7275, 16'd8768, 16'd16265, 16'd44233, 16'd22222, 16'd12601, 16'd9265, 16'd37441, 16'd5037, 16'd20152, 16'd21203, 16'd17042, 16'd44609, 16'd14661, 16'd46299, 16'd20047, 16'd2729});
	test_expansion(128'hb69cd985d194a9d7d07ca828d30fb989, {16'd14236, 16'd27574, 16'd30685, 16'd52859, 16'd23868, 16'd26007, 16'd5607, 16'd42654, 16'd37623, 16'd1244, 16'd31750, 16'd43822, 16'd46946, 16'd24961, 16'd14273, 16'd47313, 16'd37129, 16'd57644, 16'd18588, 16'd49541, 16'd26637, 16'd30654, 16'd35136, 16'd1956, 16'd64584, 16'd47564});
	test_expansion(128'h71f6e700412785b6eebc89529182987a, {16'd59068, 16'd21016, 16'd45983, 16'd32487, 16'd41069, 16'd1746, 16'd49011, 16'd44186, 16'd20145, 16'd9475, 16'd16875, 16'd642, 16'd19785, 16'd12057, 16'd21424, 16'd29299, 16'd23384, 16'd47383, 16'd7202, 16'd25589, 16'd19150, 16'd39564, 16'd47674, 16'd20038, 16'd33112, 16'd33230});
	test_expansion(128'h5bb7ddbb63264405ce3f47cf9b18152c, {16'd29911, 16'd55666, 16'd38574, 16'd18426, 16'd5199, 16'd8556, 16'd3280, 16'd50744, 16'd37365, 16'd20143, 16'd37461, 16'd59060, 16'd41223, 16'd23216, 16'd19044, 16'd54767, 16'd63071, 16'd5444, 16'd8691, 16'd30360, 16'd52338, 16'd14894, 16'd40755, 16'd51639, 16'd13476, 16'd55587});
	test_expansion(128'h129d20351c79bc36e38ba376ff666a80, {16'd57602, 16'd18007, 16'd19660, 16'd4421, 16'd54387, 16'd28942, 16'd10500, 16'd12300, 16'd21318, 16'd16503, 16'd39128, 16'd38927, 16'd27265, 16'd39611, 16'd46089, 16'd40814, 16'd38013, 16'd51981, 16'd12362, 16'd2290, 16'd42622, 16'd10149, 16'd5916, 16'd21811, 16'd5945, 16'd18846});
	test_expansion(128'h24581b45ef910a024a07b5a17e035846, {16'd6057, 16'd25047, 16'd28743, 16'd14555, 16'd4745, 16'd22377, 16'd46116, 16'd10841, 16'd46490, 16'd46518, 16'd3813, 16'd39603, 16'd64316, 16'd52701, 16'd5562, 16'd63590, 16'd5175, 16'd33661, 16'd2197, 16'd18613, 16'd39110, 16'd65097, 16'd58154, 16'd58000, 16'd52937, 16'd41362});
	test_expansion(128'hdaf1d8255bc43d1ad5a0a4e5d6c13f77, {16'd52564, 16'd35468, 16'd30010, 16'd19221, 16'd38020, 16'd57001, 16'd37304, 16'd42664, 16'd49205, 16'd7907, 16'd23585, 16'd14690, 16'd52194, 16'd19567, 16'd12624, 16'd20726, 16'd55100, 16'd39299, 16'd62268, 16'd37895, 16'd59340, 16'd10502, 16'd7164, 16'd3682, 16'd57926, 16'd42648});
	test_expansion(128'h425dba3ef17268ee7c788222781cd753, {16'd15010, 16'd26713, 16'd41344, 16'd2226, 16'd55678, 16'd6204, 16'd58275, 16'd10626, 16'd9137, 16'd42892, 16'd63951, 16'd5957, 16'd59482, 16'd60885, 16'd46561, 16'd40294, 16'd27035, 16'd32655, 16'd16391, 16'd31202, 16'd62476, 16'd27287, 16'd48438, 16'd35916, 16'd22846, 16'd225});
	test_expansion(128'h922a61127074cdafb3cd0d687468833c, {16'd56058, 16'd21279, 16'd33116, 16'd17235, 16'd30530, 16'd48633, 16'd31122, 16'd43111, 16'd43884, 16'd39238, 16'd32612, 16'd32555, 16'd59399, 16'd51243, 16'd25674, 16'd19003, 16'd16495, 16'd3185, 16'd55875, 16'd45254, 16'd8518, 16'd571, 16'd10834, 16'd4773, 16'd35446, 16'd6604});
	test_expansion(128'hf61a5c65f700edfbf6e1fd59d9a7d227, {16'd15471, 16'd6990, 16'd700, 16'd52041, 16'd28231, 16'd49304, 16'd60876, 16'd56015, 16'd36131, 16'd31757, 16'd56438, 16'd40443, 16'd1857, 16'd19470, 16'd33452, 16'd39856, 16'd44718, 16'd59854, 16'd44665, 16'd46755, 16'd37444, 16'd25761, 16'd24468, 16'd22108, 16'd131, 16'd17299});
	test_expansion(128'h2c05248c3c0316460e84ecd9dedd53dd, {16'd26579, 16'd23792, 16'd28562, 16'd26317, 16'd45314, 16'd61439, 16'd58443, 16'd25446, 16'd65008, 16'd6196, 16'd18351, 16'd49666, 16'd25774, 16'd23910, 16'd8130, 16'd13916, 16'd53800, 16'd43358, 16'd24469, 16'd52451, 16'd44022, 16'd43517, 16'd30690, 16'd55212, 16'd60902, 16'd1468});
	test_expansion(128'h4eddddea743a8d19243e4a3592547a8c, {16'd60791, 16'd34337, 16'd39283, 16'd31771, 16'd55737, 16'd32644, 16'd12095, 16'd8939, 16'd28380, 16'd12445, 16'd43813, 16'd4016, 16'd21818, 16'd64270, 16'd52097, 16'd33617, 16'd36787, 16'd42086, 16'd26981, 16'd65270, 16'd32145, 16'd12723, 16'd31952, 16'd35215, 16'd15748, 16'd8159});
	test_expansion(128'h8d5eb78677b94aa1928ed27eaf9a1561, {16'd57277, 16'd63084, 16'd38787, 16'd19961, 16'd63182, 16'd38219, 16'd49165, 16'd58524, 16'd1163, 16'd26344, 16'd33775, 16'd2294, 16'd24145, 16'd39373, 16'd22616, 16'd15918, 16'd47325, 16'd51950, 16'd6532, 16'd42784, 16'd14551, 16'd1931, 16'd10213, 16'd24626, 16'd63849, 16'd37699});
	test_expansion(128'h7b055c429c35c758eb2fa9ca644d809f, {16'd39770, 16'd15666, 16'd2781, 16'd51884, 16'd4343, 16'd62012, 16'd25929, 16'd38208, 16'd31045, 16'd28205, 16'd7471, 16'd62908, 16'd12697, 16'd35268, 16'd50184, 16'd22357, 16'd41402, 16'd23838, 16'd17340, 16'd9504, 16'd59563, 16'd22253, 16'd24579, 16'd4979, 16'd44474, 16'd51513});
	test_expansion(128'h9b91708ad6d982dd993bfcf4739ba2fc, {16'd48130, 16'd34333, 16'd22667, 16'd24537, 16'd17060, 16'd32653, 16'd45203, 16'd19517, 16'd43145, 16'd35464, 16'd11488, 16'd28529, 16'd40759, 16'd24292, 16'd31237, 16'd11983, 16'd45807, 16'd13671, 16'd59600, 16'd39830, 16'd364, 16'd9085, 16'd60157, 16'd62336, 16'd13432, 16'd59077});
	test_expansion(128'he468acaa0d34db34313fa8a02e0def18, {16'd51589, 16'd56931, 16'd41124, 16'd51702, 16'd58283, 16'd62991, 16'd17091, 16'd34749, 16'd26804, 16'd24578, 16'd65112, 16'd3057, 16'd18267, 16'd41622, 16'd62648, 16'd44191, 16'd5062, 16'd39118, 16'd39437, 16'd21677, 16'd16706, 16'd32146, 16'd61126, 16'd8188, 16'd39224, 16'd18935});
	test_expansion(128'h28681af97821d601de3cec198db65a2e, {16'd41093, 16'd51322, 16'd26001, 16'd19060, 16'd64243, 16'd36707, 16'd37201, 16'd45554, 16'd17682, 16'd58341, 16'd45353, 16'd57011, 16'd2813, 16'd297, 16'd24023, 16'd52206, 16'd51903, 16'd4113, 16'd56247, 16'd52365, 16'd27838, 16'd47670, 16'd5492, 16'd42470, 16'd17944, 16'd28389});
	test_expansion(128'h7807e3bbcda0f4d7a75d901af07d9e0e, {16'd18889, 16'd50522, 16'd46311, 16'd26667, 16'd16636, 16'd55257, 16'd24321, 16'd45906, 16'd36145, 16'd35523, 16'd59981, 16'd12280, 16'd10725, 16'd1943, 16'd37168, 16'd38843, 16'd34149, 16'd51232, 16'd42071, 16'd57562, 16'd26964, 16'd63154, 16'd50342, 16'd8910, 16'd33972, 16'd56904});
	test_expansion(128'hfe2cea3c2bcf7faf3efc691ecc999a85, {16'd21818, 16'd22383, 16'd4921, 16'd48500, 16'd32409, 16'd2893, 16'd54115, 16'd40787, 16'd3007, 16'd60841, 16'd51254, 16'd58879, 16'd36427, 16'd43473, 16'd10990, 16'd51256, 16'd59621, 16'd34706, 16'd35584, 16'd48294, 16'd37365, 16'd59033, 16'd37886, 16'd45647, 16'd8679, 16'd17472});
	test_expansion(128'h9156f92a319901675252e3de229d21b3, {16'd7698, 16'd20766, 16'd58005, 16'd43294, 16'd4480, 16'd29509, 16'd23679, 16'd37446, 16'd14674, 16'd50162, 16'd63596, 16'd9681, 16'd7678, 16'd51820, 16'd36035, 16'd33095, 16'd17845, 16'd797, 16'd53278, 16'd4012, 16'd37997, 16'd51954, 16'd32574, 16'd63492, 16'd22673, 16'd30339});
	test_expansion(128'h690e0f132f0e9853c40f82bfea784d5e, {16'd28904, 16'd1198, 16'd40458, 16'd1142, 16'd18810, 16'd3015, 16'd53352, 16'd47414, 16'd20993, 16'd12571, 16'd4935, 16'd26715, 16'd34787, 16'd28035, 16'd12437, 16'd36996, 16'd4459, 16'd56953, 16'd10564, 16'd41725, 16'd39252, 16'd19897, 16'd64965, 16'd36159, 16'd16428, 16'd9854});
	test_expansion(128'h36adf6d1a221ed325c9edd9feda1f6e7, {16'd56638, 16'd12861, 16'd31728, 16'd37555, 16'd13542, 16'd29935, 16'd16498, 16'd54549, 16'd15130, 16'd55598, 16'd12036, 16'd36927, 16'd39995, 16'd28793, 16'd14254, 16'd36662, 16'd39628, 16'd18893, 16'd48642, 16'd42640, 16'd56106, 16'd37968, 16'd20334, 16'd2575, 16'd12627, 16'd14456});
	test_expansion(128'h9ebe692355fff64ba50818b332b53063, {16'd46083, 16'd39053, 16'd21821, 16'd39514, 16'd46711, 16'd12513, 16'd51361, 16'd56060, 16'd39897, 16'd21468, 16'd2250, 16'd55803, 16'd64810, 16'd62817, 16'd55561, 16'd42203, 16'd22517, 16'd25855, 16'd22354, 16'd44868, 16'd54810, 16'd22291, 16'd43996, 16'd29599, 16'd7005, 16'd23964});
	test_expansion(128'h097fb55fee1050db17847dd7263c2c68, {16'd28615, 16'd27282, 16'd48206, 16'd25354, 16'd64186, 16'd4867, 16'd7981, 16'd25086, 16'd35347, 16'd8404, 16'd49556, 16'd23047, 16'd54911, 16'd817, 16'd47067, 16'd64123, 16'd55053, 16'd11453, 16'd30255, 16'd72, 16'd10666, 16'd65518, 16'd16671, 16'd53333, 16'd36045, 16'd25320});
	test_expansion(128'h29d4b33d558246c62d3d89b1df359d2a, {16'd46491, 16'd15301, 16'd42464, 16'd60825, 16'd56884, 16'd38266, 16'd24130, 16'd49403, 16'd40444, 16'd23266, 16'd58922, 16'd44185, 16'd39593, 16'd6261, 16'd31414, 16'd641, 16'd594, 16'd59477, 16'd59480, 16'd60742, 16'd36965, 16'd40613, 16'd15842, 16'd52798, 16'd56310, 16'd12499});
	test_expansion(128'hc2fed046a59263ad1e5f0112bbd97600, {16'd41470, 16'd22122, 16'd18468, 16'd46768, 16'd50761, 16'd22067, 16'd48585, 16'd55588, 16'd50592, 16'd10403, 16'd11983, 16'd19679, 16'd33596, 16'd34441, 16'd18511, 16'd10696, 16'd20496, 16'd39749, 16'd29802, 16'd51044, 16'd21458, 16'd21463, 16'd32848, 16'd51569, 16'd15616, 16'd54202});
	test_expansion(128'h47ccc4a3457f37052c8d07fbf97e825a, {16'd64584, 16'd36065, 16'd13619, 16'd13713, 16'd50962, 16'd11609, 16'd4007, 16'd60005, 16'd28379, 16'd18740, 16'd27662, 16'd22411, 16'd1721, 16'd3363, 16'd64639, 16'd3817, 16'd12256, 16'd62042, 16'd43062, 16'd1601, 16'd9650, 16'd15077, 16'd35126, 16'd24041, 16'd47039, 16'd12807});
	test_expansion(128'h702a4dfddf14774f824df0279119aa83, {16'd52577, 16'd57170, 16'd30750, 16'd39340, 16'd6364, 16'd32860, 16'd51784, 16'd34713, 16'd3276, 16'd54714, 16'd16056, 16'd56003, 16'd11867, 16'd27964, 16'd27543, 16'd18200, 16'd7052, 16'd19838, 16'd5913, 16'd9324, 16'd49529, 16'd7285, 16'd45878, 16'd23925, 16'd8072, 16'd49478});
	test_expansion(128'h3c224076d15a18fdd623dd6e5fc81456, {16'd22013, 16'd42838, 16'd20850, 16'd15468, 16'd60254, 16'd44809, 16'd12293, 16'd30624, 16'd12581, 16'd64412, 16'd55990, 16'd15435, 16'd10229, 16'd58259, 16'd51596, 16'd54408, 16'd35357, 16'd1957, 16'd41376, 16'd9100, 16'd42938, 16'd59192, 16'd299, 16'd51003, 16'd30905, 16'd9520});
	test_expansion(128'h2e33828d4dc200ca196f23ac0f99ed9a, {16'd42008, 16'd64822, 16'd48461, 16'd41694, 16'd47027, 16'd16509, 16'd21371, 16'd51359, 16'd38486, 16'd14288, 16'd9216, 16'd3162, 16'd47762, 16'd9462, 16'd47127, 16'd60369, 16'd30558, 16'd21207, 16'd31218, 16'd51244, 16'd46471, 16'd54001, 16'd3355, 16'd11760, 16'd38282, 16'd38143});
	test_expansion(128'hf6a2a9c1d0b008b4f1894b68f25db230, {16'd21648, 16'd30829, 16'd26074, 16'd57683, 16'd28509, 16'd11860, 16'd39449, 16'd47999, 16'd34238, 16'd41597, 16'd49317, 16'd55900, 16'd61354, 16'd41915, 16'd23159, 16'd59715, 16'd48992, 16'd36258, 16'd17421, 16'd46931, 16'd50142, 16'd20780, 16'd53980, 16'd27441, 16'd12341, 16'd13017});
	test_expansion(128'h8b8a524495e6160769f9cb57d04db25b, {16'd57568, 16'd61906, 16'd42961, 16'd41394, 16'd173, 16'd116, 16'd28342, 16'd58705, 16'd48249, 16'd19780, 16'd44169, 16'd30123, 16'd39989, 16'd7140, 16'd27531, 16'd21605, 16'd48270, 16'd25780, 16'd36215, 16'd44005, 16'd28472, 16'd24666, 16'd22821, 16'd59934, 16'd16617, 16'd39767});
	test_expansion(128'hc3313cab1551fd9143c54e9e2c0eda06, {16'd37183, 16'd40397, 16'd52511, 16'd58349, 16'd20100, 16'd51284, 16'd5325, 16'd57988, 16'd59503, 16'd45042, 16'd28733, 16'd4274, 16'd29671, 16'd27617, 16'd11718, 16'd39232, 16'd61692, 16'd2958, 16'd39843, 16'd22463, 16'd192, 16'd42298, 16'd44875, 16'd5476, 16'd2584, 16'd62979});
	test_expansion(128'h02ec8d25605cbf8a1e8256892fa2c978, {16'd39971, 16'd42463, 16'd24743, 16'd20996, 16'd12618, 16'd9473, 16'd4344, 16'd49133, 16'd44099, 16'd7770, 16'd24920, 16'd63497, 16'd20719, 16'd17295, 16'd27178, 16'd24224, 16'd33743, 16'd33847, 16'd5916, 16'd22462, 16'd55330, 16'd13923, 16'd24670, 16'd11438, 16'd43287, 16'd61264});
	test_expansion(128'h26bc1acdc323384ae65586d15be0490e, {16'd45694, 16'd61292, 16'd49961, 16'd47417, 16'd17597, 16'd60758, 16'd3104, 16'd55376, 16'd38133, 16'd41830, 16'd51521, 16'd7361, 16'd32902, 16'd2512, 16'd39203, 16'd5518, 16'd15182, 16'd11638, 16'd35302, 16'd57546, 16'd49133, 16'd24300, 16'd61569, 16'd5907, 16'd18904, 16'd43287});
	test_expansion(128'h9ffec046806fc49a0d3068ba6bf71a83, {16'd17315, 16'd2395, 16'd12409, 16'd26454, 16'd58822, 16'd29886, 16'd32370, 16'd32546, 16'd44345, 16'd58117, 16'd52888, 16'd8969, 16'd16621, 16'd37873, 16'd45757, 16'd27366, 16'd41344, 16'd49284, 16'd37240, 16'd56587, 16'd4617, 16'd7543, 16'd4819, 16'd51968, 16'd61093, 16'd64997});
	test_expansion(128'h427d0f84b8f6c8f176b833edf3e70c7a, {16'd54280, 16'd1154, 16'd43801, 16'd19163, 16'd48241, 16'd45246, 16'd61827, 16'd4938, 16'd61652, 16'd5571, 16'd57577, 16'd42711, 16'd64968, 16'd3847, 16'd29324, 16'd26189, 16'd23515, 16'd40808, 16'd6121, 16'd17651, 16'd35636, 16'd9442, 16'd13067, 16'd22076, 16'd46001, 16'd26546});
	test_expansion(128'hfb526a1aeb23e219dfb717dfd9c96049, {16'd15100, 16'd55751, 16'd36390, 16'd34863, 16'd58522, 16'd58784, 16'd45447, 16'd25866, 16'd58219, 16'd56883, 16'd43815, 16'd46813, 16'd4447, 16'd49865, 16'd2836, 16'd18841, 16'd20946, 16'd50484, 16'd40672, 16'd15183, 16'd25944, 16'd31257, 16'd35516, 16'd5155, 16'd1994, 16'd31898});
	test_expansion(128'hfa268af01af3efceb702a473cb170d74, {16'd27320, 16'd48748, 16'd41652, 16'd23923, 16'd59657, 16'd6027, 16'd63936, 16'd29079, 16'd20963, 16'd6059, 16'd30687, 16'd25280, 16'd8979, 16'd45778, 16'd54490, 16'd1673, 16'd29906, 16'd34312, 16'd2102, 16'd6211, 16'd30354, 16'd57482, 16'd58883, 16'd18915, 16'd51072, 16'd33596});
	test_expansion(128'h938eda2f0445a6d81c421b22ba34354a, {16'd46922, 16'd42623, 16'd40718, 16'd21986, 16'd9320, 16'd65184, 16'd16568, 16'd63394, 16'd14709, 16'd38563, 16'd44446, 16'd4675, 16'd44765, 16'd63224, 16'd1417, 16'd22207, 16'd35637, 16'd44654, 16'd8424, 16'd12323, 16'd27756, 16'd40797, 16'd14272, 16'd1628, 16'd10495, 16'd32075});
	test_expansion(128'hdc124cb0b3074b21c1a789dbed6fde69, {16'd11631, 16'd62339, 16'd40658, 16'd46950, 16'd24484, 16'd24688, 16'd1360, 16'd61085, 16'd51214, 16'd20431, 16'd24820, 16'd9514, 16'd23466, 16'd4320, 16'd47161, 16'd25973, 16'd46917, 16'd13980, 16'd38336, 16'd26344, 16'd13943, 16'd27307, 16'd39059, 16'd11649, 16'd24253, 16'd54723});
	test_expansion(128'h83539886460dd5cfa52fa6b6bec6ecb3, {16'd8182, 16'd49435, 16'd65450, 16'd11531, 16'd14120, 16'd63031, 16'd54162, 16'd29568, 16'd40239, 16'd58201, 16'd29901, 16'd39845, 16'd42335, 16'd52037, 16'd48264, 16'd21969, 16'd32512, 16'd5182, 16'd17527, 16'd33858, 16'd13671, 16'd18158, 16'd26849, 16'd39896, 16'd39237, 16'd5985});
	test_expansion(128'h7116f5d126ec688c4cabf5b5e839fc31, {16'd37437, 16'd12616, 16'd36591, 16'd27869, 16'd34592, 16'd57249, 16'd61686, 16'd21246, 16'd37324, 16'd48645, 16'd35566, 16'd56427, 16'd27341, 16'd10090, 16'd12611, 16'd23980, 16'd50055, 16'd51203, 16'd10357, 16'd49467, 16'd22195, 16'd7895, 16'd47128, 16'd53091, 16'd63032, 16'd31292});
	test_expansion(128'h58272ef6ffd68d06916abb7c4270114f, {16'd40929, 16'd64333, 16'd40859, 16'd3238, 16'd46869, 16'd7583, 16'd45994, 16'd59057, 16'd2570, 16'd20525, 16'd25836, 16'd631, 16'd17961, 16'd59117, 16'd44066, 16'd4089, 16'd26231, 16'd1651, 16'd27798, 16'd34876, 16'd20011, 16'd25005, 16'd38062, 16'd22665, 16'd39078, 16'd26204});
	test_expansion(128'h3359b472b04df05aa1ec24a4f344cb7a, {16'd6411, 16'd60466, 16'd58619, 16'd4125, 16'd24390, 16'd28401, 16'd58619, 16'd11530, 16'd18512, 16'd26355, 16'd52991, 16'd9586, 16'd4456, 16'd58252, 16'd54902, 16'd12022, 16'd30226, 16'd31894, 16'd34091, 16'd25925, 16'd6582, 16'd64799, 16'd9293, 16'd61912, 16'd31691, 16'd41053});
	test_expansion(128'ha5e8c72b167450e7abb106bb135bf3b5, {16'd42104, 16'd58993, 16'd61400, 16'd63134, 16'd65177, 16'd7442, 16'd55804, 16'd22076, 16'd39517, 16'd55965, 16'd41853, 16'd32704, 16'd14297, 16'd10297, 16'd3966, 16'd64851, 16'd32122, 16'd60133, 16'd56671, 16'd45058, 16'd34627, 16'd65162, 16'd19498, 16'd39445, 16'd23845, 16'd33201});
	test_expansion(128'h7b92932724521f6f34e51db021ef873d, {16'd41970, 16'd1137, 16'd15913, 16'd38469, 16'd37129, 16'd65151, 16'd10908, 16'd9009, 16'd37779, 16'd8359, 16'd12148, 16'd25669, 16'd8352, 16'd56926, 16'd13127, 16'd58212, 16'd1322, 16'd49076, 16'd894, 16'd40041, 16'd24126, 16'd7903, 16'd2795, 16'd30244, 16'd58227, 16'd29709});
	test_expansion(128'h9ffb475137cd5cf15639c54f537e9b61, {16'd1274, 16'd5000, 16'd22395, 16'd63664, 16'd23982, 16'd12521, 16'd32738, 16'd30431, 16'd58362, 16'd41362, 16'd44466, 16'd38015, 16'd28046, 16'd23547, 16'd10601, 16'd42401, 16'd14370, 16'd25503, 16'd26899, 16'd3520, 16'd46967, 16'd39591, 16'd60655, 16'd36048, 16'd34629, 16'd17385});
	test_expansion(128'h060ecfe235c92a76054d86a87b0053a0, {16'd43678, 16'd179, 16'd43189, 16'd27509, 16'd58183, 16'd33525, 16'd49826, 16'd47941, 16'd54717, 16'd55009, 16'd29639, 16'd60408, 16'd43688, 16'd25503, 16'd41174, 16'd11348, 16'd40169, 16'd17613, 16'd11525, 16'd10781, 16'd47653, 16'd20076, 16'd4528, 16'd47055, 16'd9848, 16'd24431});
	test_expansion(128'h809d1248b46258783af7f91a25fe8e0e, {16'd21554, 16'd8749, 16'd5015, 16'd29483, 16'd15477, 16'd18917, 16'd6015, 16'd59089, 16'd24276, 16'd48212, 16'd17417, 16'd55346, 16'd3865, 16'd30180, 16'd16009, 16'd19097, 16'd32622, 16'd43303, 16'd18559, 16'd8230, 16'd34931, 16'd16785, 16'd43391, 16'd17422, 16'd16849, 16'd18368});
	test_expansion(128'h059625d9f97df43288ac2c7f9c4e4760, {16'd51380, 16'd55672, 16'd13112, 16'd11432, 16'd35302, 16'd33813, 16'd23622, 16'd48811, 16'd33205, 16'd9432, 16'd17246, 16'd20852, 16'd989, 16'd22738, 16'd56735, 16'd41699, 16'd61223, 16'd50246, 16'd63206, 16'd11998, 16'd48908, 16'd10896, 16'd9699, 16'd10479, 16'd29800, 16'd62771});
	test_expansion(128'h0b729d344bd812840d56f6ac111f0ffb, {16'd63487, 16'd41826, 16'd55809, 16'd17317, 16'd29970, 16'd56619, 16'd34761, 16'd27415, 16'd39404, 16'd48604, 16'd28293, 16'd47261, 16'd43138, 16'd59228, 16'd21843, 16'd26536, 16'd61866, 16'd20243, 16'd26505, 16'd5935, 16'd28304, 16'd52999, 16'd47111, 16'd23490, 16'd9795, 16'd49613});
	test_expansion(128'h35442137ca7df00f9e0252a2504dc8ab, {16'd42746, 16'd4864, 16'd61392, 16'd43358, 16'd31524, 16'd57520, 16'd57132, 16'd55926, 16'd26609, 16'd10527, 16'd29554, 16'd31864, 16'd62351, 16'd62101, 16'd18747, 16'd48385, 16'd25464, 16'd18522, 16'd52809, 16'd58856, 16'd12245, 16'd53896, 16'd59950, 16'd34514, 16'd18245, 16'd14399});
	test_expansion(128'h1247a0a9837d71c4b5105ee602477453, {16'd11923, 16'd29199, 16'd35365, 16'd62904, 16'd19517, 16'd6014, 16'd55544, 16'd52952, 16'd62844, 16'd41385, 16'd61724, 16'd27271, 16'd29226, 16'd65454, 16'd50154, 16'd17601, 16'd11988, 16'd10922, 16'd54776, 16'd25735, 16'd14994, 16'd58979, 16'd29548, 16'd29047, 16'd28820, 16'd58186});
	test_expansion(128'hf2182c46226a2e052f761954b819c782, {16'd33126, 16'd20505, 16'd7820, 16'd24648, 16'd19654, 16'd31582, 16'd53863, 16'd27481, 16'd32733, 16'd57189, 16'd60578, 16'd31569, 16'd29584, 16'd14810, 16'd64771, 16'd61262, 16'd16757, 16'd247, 16'd5694, 16'd62680, 16'd58404, 16'd40180, 16'd41266, 16'd49398, 16'd40017, 16'd63171});
	test_expansion(128'h20c87a8826cc2e2bea34a9879b851996, {16'd52769, 16'd44400, 16'd46731, 16'd27267, 16'd29695, 16'd53235, 16'd16794, 16'd44380, 16'd43105, 16'd63753, 16'd53387, 16'd37827, 16'd23199, 16'd9022, 16'd3111, 16'd62655, 16'd19841, 16'd253, 16'd53127, 16'd8718, 16'd64233, 16'd33725, 16'd26445, 16'd34796, 16'd58007, 16'd61530});
	test_expansion(128'hcfac6028c707a70e65d4764fc6f12ee3, {16'd29029, 16'd58890, 16'd32670, 16'd37381, 16'd29849, 16'd59742, 16'd52416, 16'd38018, 16'd19351, 16'd40106, 16'd6964, 16'd54967, 16'd10743, 16'd29178, 16'd47090, 16'd23861, 16'd32715, 16'd59858, 16'd54951, 16'd51292, 16'd13764, 16'd18907, 16'd23888, 16'd39522, 16'd3539, 16'd2427});
	test_expansion(128'hf0cd2b2042a30f5ed7b099af6d1a405e, {16'd18446, 16'd58506, 16'd58434, 16'd23920, 16'd12282, 16'd31036, 16'd45931, 16'd3325, 16'd13734, 16'd63046, 16'd19309, 16'd53289, 16'd11641, 16'd16095, 16'd11931, 16'd22634, 16'd56095, 16'd16507, 16'd19805, 16'd49863, 16'd28846, 16'd52851, 16'd62537, 16'd47496, 16'd1859, 16'd55487});
	test_expansion(128'h8010fed1ac33a75bbd52aa633f0f88a7, {16'd56184, 16'd26459, 16'd6379, 16'd22542, 16'd28946, 16'd15148, 16'd29247, 16'd51352, 16'd55623, 16'd16901, 16'd64089, 16'd6894, 16'd32998, 16'd46532, 16'd38148, 16'd48597, 16'd48710, 16'd17373, 16'd44131, 16'd63037, 16'd12325, 16'd30821, 16'd39471, 16'd64691, 16'd55179, 16'd43770});
	test_expansion(128'h4aa2ae13646b91087c5046c8de2acf96, {16'd34038, 16'd16397, 16'd23359, 16'd24427, 16'd50431, 16'd35782, 16'd18913, 16'd15807, 16'd54591, 16'd5540, 16'd15019, 16'd49286, 16'd22670, 16'd7066, 16'd63425, 16'd22516, 16'd4985, 16'd1851, 16'd47169, 16'd45806, 16'd56789, 16'd40210, 16'd40583, 16'd34887, 16'd39231, 16'd28696});
	test_expansion(128'h4aa8657e809f28f81c35eb8b29b3097d, {16'd53690, 16'd20257, 16'd35980, 16'd15344, 16'd51285, 16'd30939, 16'd21245, 16'd30327, 16'd46273, 16'd55153, 16'd18540, 16'd65247, 16'd47395, 16'd874, 16'd47760, 16'd26356, 16'd57046, 16'd40578, 16'd53424, 16'd56275, 16'd2053, 16'd14702, 16'd21827, 16'd55626, 16'd21594, 16'd13307});
	test_expansion(128'h964f102eb067c0a638c166f5f2fad5e1, {16'd8029, 16'd43785, 16'd59608, 16'd51561, 16'd17288, 16'd16328, 16'd14934, 16'd61713, 16'd58923, 16'd40886, 16'd50641, 16'd21643, 16'd4569, 16'd39392, 16'd13152, 16'd7325, 16'd36964, 16'd16944, 16'd20306, 16'd61224, 16'd46634, 16'd64523, 16'd26062, 16'd34095, 16'd16373, 16'd1856});
	test_expansion(128'he2a28951d00fa2d230617cddc5ffefa2, {16'd37658, 16'd46391, 16'd12567, 16'd29162, 16'd58721, 16'd3544, 16'd12910, 16'd55937, 16'd53394, 16'd37510, 16'd57264, 16'd48841, 16'd25801, 16'd1435, 16'd11123, 16'd29778, 16'd14144, 16'd22297, 16'd45539, 16'd53677, 16'd4674, 16'd40477, 16'd12246, 16'd32891, 16'd27705, 16'd27955});
	test_expansion(128'h7c910f89e77dda478e40d8f9564970b0, {16'd49477, 16'd17024, 16'd9066, 16'd51715, 16'd4475, 16'd22311, 16'd11126, 16'd49392, 16'd10147, 16'd35975, 16'd36221, 16'd59898, 16'd10083, 16'd62317, 16'd30461, 16'd6592, 16'd18034, 16'd21930, 16'd23725, 16'd29420, 16'd51318, 16'd35346, 16'd33883, 16'd61541, 16'd30943, 16'd33001});
	test_expansion(128'h755223cc63f3017736d107752f1b7c42, {16'd34032, 16'd52321, 16'd38688, 16'd64557, 16'd49642, 16'd17275, 16'd2002, 16'd45582, 16'd26759, 16'd59866, 16'd33615, 16'd18257, 16'd5118, 16'd11673, 16'd26965, 16'd6268, 16'd29747, 16'd12519, 16'd10104, 16'd51519, 16'd34024, 16'd23413, 16'd57947, 16'd62757, 16'd30001, 16'd51436});
	test_expansion(128'h049dd09b8d13d23e03ee1cfe9a0b21b1, {16'd49578, 16'd37305, 16'd58251, 16'd4577, 16'd28449, 16'd18636, 16'd36371, 16'd13834, 16'd14763, 16'd17693, 16'd41677, 16'd26498, 16'd15295, 16'd17005, 16'd22941, 16'd27166, 16'd62145, 16'd26919, 16'd24882, 16'd25343, 16'd44642, 16'd30895, 16'd465, 16'd55750, 16'd44550, 16'd65430});
	test_expansion(128'haa4db199a0c747dfcaf9a6bf228c1376, {16'd3509, 16'd41192, 16'd13221, 16'd12126, 16'd17943, 16'd17304, 16'd26922, 16'd33146, 16'd24741, 16'd3676, 16'd6805, 16'd35308, 16'd26828, 16'd36789, 16'd61848, 16'd59246, 16'd13173, 16'd31177, 16'd17968, 16'd33659, 16'd60765, 16'd34320, 16'd59702, 16'd10533, 16'd58849, 16'd22169});
	test_expansion(128'hc5a3a66140b55751d54d1dd611ffbcdb, {16'd58365, 16'd46774, 16'd35664, 16'd23194, 16'd5773, 16'd43066, 16'd39074, 16'd65292, 16'd32642, 16'd55925, 16'd41431, 16'd39802, 16'd39199, 16'd55120, 16'd57987, 16'd60019, 16'd65460, 16'd59596, 16'd27964, 16'd37837, 16'd52890, 16'd4387, 16'd29085, 16'd18998, 16'd29683, 16'd31679});
	test_expansion(128'h75b307cff8270e4d4eca0ba34ccd0a2c, {16'd3934, 16'd33026, 16'd50754, 16'd58484, 16'd38595, 16'd34121, 16'd23415, 16'd3435, 16'd5782, 16'd13771, 16'd62348, 16'd425, 16'd6654, 16'd8622, 16'd13880, 16'd23695, 16'd19426, 16'd5775, 16'd46892, 16'd59004, 16'd11062, 16'd21400, 16'd28345, 16'd3556, 16'd17825, 16'd58475});
	test_expansion(128'h27abcc535e69b3d45037b6d19b4f5162, {16'd12652, 16'd27076, 16'd41608, 16'd65137, 16'd11788, 16'd21168, 16'd62217, 16'd13160, 16'd52239, 16'd5362, 16'd14640, 16'd17920, 16'd10400, 16'd18931, 16'd57258, 16'd7225, 16'd290, 16'd1038, 16'd49490, 16'd17500, 16'd56365, 16'd43249, 16'd11059, 16'd12218, 16'd41508, 16'd37942});
	test_expansion(128'h75141fc767e33202f101fd61c8cfb23f, {16'd65046, 16'd8369, 16'd60105, 16'd39384, 16'd46745, 16'd30023, 16'd36745, 16'd42662, 16'd36428, 16'd43753, 16'd6443, 16'd7768, 16'd64306, 16'd23866, 16'd48634, 16'd24706, 16'd31916, 16'd16737, 16'd11263, 16'd2236, 16'd16332, 16'd57500, 16'd32556, 16'd49846, 16'd18514, 16'd1584});
	test_expansion(128'h0d6dd0649fc3624d8372a2921f7f5228, {16'd49812, 16'd51962, 16'd16440, 16'd42647, 16'd22488, 16'd12377, 16'd33858, 16'd22995, 16'd57070, 16'd46236, 16'd26631, 16'd43892, 16'd4630, 16'd32477, 16'd11595, 16'd12223, 16'd62602, 16'd894, 16'd52485, 16'd12903, 16'd14621, 16'd44048, 16'd54295, 16'd15283, 16'd7323, 16'd60714});
	test_expansion(128'h6ba85e799f80998c1566fde645770a86, {16'd44507, 16'd44034, 16'd58840, 16'd5908, 16'd40421, 16'd32690, 16'd33518, 16'd22572, 16'd4155, 16'd26032, 16'd21174, 16'd27176, 16'd64205, 16'd22535, 16'd42888, 16'd24837, 16'd30835, 16'd53910, 16'd17650, 16'd42486, 16'd36394, 16'd56774, 16'd5884, 16'd56928, 16'd20982, 16'd20395});
	test_expansion(128'hfdb5ec844fc820b40ae53a2c399a5155, {16'd13138, 16'd21417, 16'd35653, 16'd33608, 16'd45989, 16'd811, 16'd59903, 16'd7848, 16'd48610, 16'd3811, 16'd36628, 16'd972, 16'd36032, 16'd24215, 16'd50717, 16'd1990, 16'd50020, 16'd24556, 16'd58616, 16'd12133, 16'd54923, 16'd38805, 16'd8532, 16'd5892, 16'd28831, 16'd2341});
	test_expansion(128'hdc7436a5016286928b8acdff48f9c8c5, {16'd2551, 16'd38634, 16'd61322, 16'd55320, 16'd48831, 16'd59287, 16'd9097, 16'd50785, 16'd8174, 16'd13599, 16'd37113, 16'd57514, 16'd5955, 16'd42021, 16'd4502, 16'd15865, 16'd39519, 16'd46554, 16'd58886, 16'd22608, 16'd31223, 16'd13632, 16'd16382, 16'd51077, 16'd54438, 16'd25926});
	test_expansion(128'hf7e70801458f2fb91c955f4881c75f90, {16'd35531, 16'd7599, 16'd13849, 16'd17792, 16'd34053, 16'd14880, 16'd58303, 16'd24929, 16'd43077, 16'd2827, 16'd61149, 16'd22156, 16'd3595, 16'd28654, 16'd27298, 16'd52642, 16'd45870, 16'd63779, 16'd43416, 16'd15033, 16'd39345, 16'd8875, 16'd54894, 16'd34609, 16'd35289, 16'd53268});
	test_expansion(128'haa860377619644dae71b04d1cd456659, {16'd36757, 16'd32054, 16'd26966, 16'd64113, 16'd23456, 16'd58399, 16'd47505, 16'd31669, 16'd50022, 16'd28774, 16'd35968, 16'd11488, 16'd10395, 16'd55781, 16'd23773, 16'd7893, 16'd26770, 16'd21730, 16'd46885, 16'd56965, 16'd31042, 16'd51745, 16'd46858, 16'd48628, 16'd52256, 16'd13190});
	test_expansion(128'h3b69c3b9c5cd13a6d9997aa895be47d7, {16'd34606, 16'd53927, 16'd50440, 16'd1102, 16'd11420, 16'd16262, 16'd24590, 16'd55095, 16'd50643, 16'd54812, 16'd56499, 16'd6652, 16'd45326, 16'd4279, 16'd34711, 16'd58521, 16'd22252, 16'd49926, 16'd25500, 16'd9040, 16'd26787, 16'd16516, 16'd17734, 16'd48135, 16'd31915, 16'd10515});
	test_expansion(128'h8967417b8037bfeb3271a401469428b2, {16'd62440, 16'd13106, 16'd10012, 16'd7957, 16'd57807, 16'd3611, 16'd9082, 16'd46104, 16'd14669, 16'd9771, 16'd36148, 16'd23763, 16'd18987, 16'd10627, 16'd23341, 16'd19033, 16'd6415, 16'd20174, 16'd32009, 16'd51800, 16'd15456, 16'd51087, 16'd39291, 16'd62637, 16'd49555, 16'd57491});
	test_expansion(128'h4fe160fb052a33952282431272f90311, {16'd29085, 16'd12590, 16'd29145, 16'd45039, 16'd53916, 16'd61112, 16'd52446, 16'd2879, 16'd9057, 16'd44447, 16'd18259, 16'd15050, 16'd32503, 16'd317, 16'd32378, 16'd44319, 16'd16881, 16'd63394, 16'd14055, 16'd32622, 16'd37789, 16'd2928, 16'd14504, 16'd4009, 16'd7216, 16'd1125});
	test_expansion(128'h9089d4fba51ea2415ab845ad5d7c55a3, {16'd35976, 16'd49164, 16'd29899, 16'd40227, 16'd4603, 16'd44576, 16'd28419, 16'd32562, 16'd16541, 16'd25146, 16'd60943, 16'd58901, 16'd25628, 16'd23442, 16'd14413, 16'd37999, 16'd65455, 16'd29792, 16'd60073, 16'd8473, 16'd54284, 16'd53358, 16'd47368, 16'd12984, 16'd21177, 16'd37492});
	test_expansion(128'h6a048a725678e071a49f28619a64346e, {16'd59617, 16'd54764, 16'd33955, 16'd60125, 16'd43722, 16'd38191, 16'd13818, 16'd57700, 16'd37911, 16'd25035, 16'd2710, 16'd13686, 16'd43420, 16'd7365, 16'd1322, 16'd49916, 16'd25756, 16'd49014, 16'd46368, 16'd45292, 16'd61864, 16'd38444, 16'd40022, 16'd26202, 16'd23969, 16'd17610});
	test_expansion(128'h6561ae4071eaf853143705acbdf22dc9, {16'd51200, 16'd55555, 16'd32460, 16'd14786, 16'd54349, 16'd61305, 16'd30732, 16'd42182, 16'd41781, 16'd51872, 16'd44021, 16'd32479, 16'd10216, 16'd3000, 16'd31436, 16'd9893, 16'd13751, 16'd26748, 16'd2716, 16'd18780, 16'd6772, 16'd11167, 16'd7696, 16'd35301, 16'd9042, 16'd4891});
	test_expansion(128'h13bd59d21fc0db5800c5d280c0165491, {16'd18421, 16'd939, 16'd26053, 16'd21722, 16'd17276, 16'd59438, 16'd26142, 16'd20108, 16'd12889, 16'd41906, 16'd56222, 16'd15993, 16'd47277, 16'd19891, 16'd5373, 16'd59329, 16'd53685, 16'd18109, 16'd41164, 16'd24523, 16'd61952, 16'd54910, 16'd4974, 16'd62404, 16'd45469, 16'd19477});
	test_expansion(128'hfa89ff3a79f8ebe46de542989c2a0e6b, {16'd39911, 16'd52910, 16'd24759, 16'd61547, 16'd46742, 16'd16556, 16'd30737, 16'd64448, 16'd27936, 16'd43362, 16'd45285, 16'd8085, 16'd16104, 16'd16460, 16'd59732, 16'd47147, 16'd25824, 16'd328, 16'd31411, 16'd25509, 16'd61910, 16'd14706, 16'd57038, 16'd56702, 16'd50556, 16'd29036});
	test_expansion(128'h979fae7d640e3e87e859f820b16cf2ad, {16'd14988, 16'd64575, 16'd9655, 16'd7548, 16'd34083, 16'd37539, 16'd34254, 16'd38277, 16'd60961, 16'd33668, 16'd49285, 16'd55244, 16'd30145, 16'd16546, 16'd5980, 16'd5394, 16'd13181, 16'd33456, 16'd5241, 16'd54558, 16'd56706, 16'd51547, 16'd53154, 16'd63266, 16'd48046, 16'd12144});
	test_expansion(128'h76f1fadbf8b3103a84d7d217b6893d94, {16'd12012, 16'd47611, 16'd35000, 16'd12885, 16'd4523, 16'd34631, 16'd34560, 16'd48294, 16'd13919, 16'd18001, 16'd23615, 16'd22449, 16'd49438, 16'd53479, 16'd17974, 16'd26453, 16'd25188, 16'd45686, 16'd22737, 16'd2775, 16'd29692, 16'd43860, 16'd8437, 16'd7131, 16'd27256, 16'd5417});
	test_expansion(128'h93da09caed06b67184a122dd7c71c80b, {16'd54961, 16'd61998, 16'd9749, 16'd43367, 16'd20260, 16'd22633, 16'd53950, 16'd23441, 16'd50330, 16'd46026, 16'd13333, 16'd12051, 16'd59109, 16'd4515, 16'd24518, 16'd31288, 16'd50527, 16'd35167, 16'd44638, 16'd10647, 16'd26533, 16'd22411, 16'd20585, 16'd44597, 16'd44527, 16'd2940});
	test_expansion(128'h63105c807442837c607bbdc01c8e731f, {16'd62067, 16'd33842, 16'd10619, 16'd49269, 16'd14832, 16'd37029, 16'd64247, 16'd33596, 16'd11490, 16'd30981, 16'd64675, 16'd44665, 16'd10204, 16'd12309, 16'd8112, 16'd64510, 16'd59180, 16'd32997, 16'd30652, 16'd44588, 16'd16942, 16'd19578, 16'd38781, 16'd11316, 16'd53684, 16'd40041});
	test_expansion(128'h3f62524bcc80ed509d7fcd11b15e782f, {16'd28671, 16'd63312, 16'd43064, 16'd36580, 16'd29540, 16'd48988, 16'd35727, 16'd12228, 16'd8196, 16'd51669, 16'd52292, 16'd19730, 16'd55347, 16'd54256, 16'd16386, 16'd50268, 16'd7622, 16'd3589, 16'd55320, 16'd378, 16'd5132, 16'd63312, 16'd60476, 16'd13995, 16'd15681, 16'd63852});
	test_expansion(128'h2e844990e6c225cbb86ff06427eef2a5, {16'd35132, 16'd13335, 16'd58260, 16'd6494, 16'd8010, 16'd31068, 16'd47461, 16'd37020, 16'd29980, 16'd17058, 16'd46077, 16'd40788, 16'd6801, 16'd53868, 16'd41588, 16'd2834, 16'd48215, 16'd10077, 16'd28579, 16'd13289, 16'd64824, 16'd32742, 16'd54007, 16'd49674, 16'd41540, 16'd46098});
	test_expansion(128'h4d37cf32e6a4bdad093b961cac172c67, {16'd19693, 16'd48975, 16'd38378, 16'd4008, 16'd32954, 16'd25255, 16'd9600, 16'd10243, 16'd65067, 16'd6350, 16'd42172, 16'd1321, 16'd21296, 16'd29415, 16'd29858, 16'd20231, 16'd58269, 16'd59361, 16'd128, 16'd21155, 16'd33803, 16'd36575, 16'd37525, 16'd16896, 16'd25825, 16'd46261});
	test_expansion(128'h3649e73474a3cc3d01a3ab907c513ebb, {16'd48359, 16'd54263, 16'd19795, 16'd42542, 16'd33287, 16'd32122, 16'd34326, 16'd57505, 16'd58467, 16'd27504, 16'd23648, 16'd59026, 16'd27875, 16'd15451, 16'd53163, 16'd22640, 16'd58527, 16'd61363, 16'd3031, 16'd39934, 16'd183, 16'd64573, 16'd25348, 16'd32179, 16'd33125, 16'd17893});
	test_expansion(128'h983976eb12b17e6278d0b00c2b44c11f, {16'd3307, 16'd57125, 16'd7811, 16'd38784, 16'd48366, 16'd28058, 16'd27622, 16'd28681, 16'd50438, 16'd62361, 16'd12484, 16'd45633, 16'd55776, 16'd63386, 16'd15739, 16'd18154, 16'd58151, 16'd6020, 16'd58401, 16'd11532, 16'd35013, 16'd1021, 16'd2997, 16'd56765, 16'd58023, 16'd48469});
	test_expansion(128'he4674b5f55ff8904d8d9ea98e8e5ec35, {16'd38678, 16'd42202, 16'd148, 16'd23081, 16'd36641, 16'd36667, 16'd25994, 16'd61660, 16'd14847, 16'd20835, 16'd22087, 16'd19649, 16'd27673, 16'd53144, 16'd11292, 16'd566, 16'd42133, 16'd19590, 16'd2339, 16'd43689, 16'd50009, 16'd45794, 16'd49475, 16'd54910, 16'd21169, 16'd59055});
	test_expansion(128'h43fbe307abbc645edf897a2a00348cd1, {16'd41820, 16'd42774, 16'd17984, 16'd49065, 16'd13982, 16'd54673, 16'd6937, 16'd36722, 16'd12886, 16'd19236, 16'd24436, 16'd31973, 16'd33031, 16'd21614, 16'd42773, 16'd11127, 16'd43276, 16'd2851, 16'd28332, 16'd59890, 16'd22667, 16'd789, 16'd31270, 16'd3770, 16'd11096, 16'd26416});
	test_expansion(128'h7de6fb63bb898d15bfb0da394aa611c4, {16'd44098, 16'd14694, 16'd36243, 16'd64833, 16'd58747, 16'd17305, 16'd30988, 16'd25974, 16'd47618, 16'd42829, 16'd25584, 16'd7128, 16'd50888, 16'd16649, 16'd36105, 16'd63320, 16'd28514, 16'd57148, 16'd32108, 16'd15289, 16'd2526, 16'd39914, 16'd21980, 16'd5330, 16'd53982, 16'd2515});
	test_expansion(128'h8f4191d6c41a0b3e0e2e944aeb8e0e71, {16'd10696, 16'd11696, 16'd10123, 16'd32533, 16'd40440, 16'd56924, 16'd51577, 16'd43859, 16'd47165, 16'd36610, 16'd59852, 16'd1247, 16'd23103, 16'd22646, 16'd45477, 16'd63389, 16'd37607, 16'd32144, 16'd46966, 16'd6151, 16'd3463, 16'd33859, 16'd3046, 16'd46067, 16'd8608, 16'd39570});
	test_expansion(128'h83263b223d1e05834b5c214c5d406db3, {16'd21775, 16'd59523, 16'd59960, 16'd63815, 16'd31613, 16'd20220, 16'd8793, 16'd49156, 16'd6642, 16'd19547, 16'd38815, 16'd29203, 16'd43484, 16'd53349, 16'd9773, 16'd51181, 16'd56611, 16'd59120, 16'd3806, 16'd32545, 16'd48575, 16'd11631, 16'd10262, 16'd50211, 16'd53413, 16'd43752});
	test_expansion(128'h8c64410b9fe2ff7f91b018d5e537bd55, {16'd9464, 16'd58371, 16'd4095, 16'd3901, 16'd46241, 16'd39177, 16'd48351, 16'd14274, 16'd16505, 16'd11874, 16'd35209, 16'd54267, 16'd46431, 16'd25917, 16'd35585, 16'd26776, 16'd7666, 16'd56998, 16'd17827, 16'd15788, 16'd21476, 16'd58709, 16'd25288, 16'd31107, 16'd19611, 16'd41871});
	test_expansion(128'ha5f5a58db14c044fbd4215d68e4ed854, {16'd76, 16'd65284, 16'd11544, 16'd51480, 16'd11313, 16'd31880, 16'd7129, 16'd61630, 16'd23106, 16'd36747, 16'd32655, 16'd42474, 16'd32294, 16'd60323, 16'd13001, 16'd11152, 16'd9110, 16'd36797, 16'd39428, 16'd19190, 16'd34218, 16'd57090, 16'd60155, 16'd34702, 16'd25833, 16'd30547});
	test_expansion(128'h742a855a5b01f7127091412ff18de943, {16'd19038, 16'd50780, 16'd22267, 16'd50774, 16'd8526, 16'd39234, 16'd51165, 16'd4380, 16'd55832, 16'd41546, 16'd18072, 16'd14695, 16'd40992, 16'd64644, 16'd669, 16'd29856, 16'd9209, 16'd45715, 16'd26557, 16'd49832, 16'd26880, 16'd23680, 16'd16430, 16'd26110, 16'd61268, 16'd47812});
	test_expansion(128'h0c9248571d6016164177d031912df6cc, {16'd43316, 16'd62301, 16'd10729, 16'd20609, 16'd1608, 16'd20763, 16'd12735, 16'd53865, 16'd39246, 16'd7233, 16'd20827, 16'd38185, 16'd17271, 16'd46031, 16'd3984, 16'd29786, 16'd33335, 16'd23668, 16'd48253, 16'd6999, 16'd47604, 16'd56318, 16'd34292, 16'd60230, 16'd40750, 16'd41662});
	test_expansion(128'hfa0294fdea9485a10f7c22772d9f65f1, {16'd13563, 16'd41992, 16'd44340, 16'd37062, 16'd26208, 16'd9414, 16'd38368, 16'd2295, 16'd9497, 16'd51359, 16'd48765, 16'd15269, 16'd30012, 16'd5454, 16'd25916, 16'd52296, 16'd54477, 16'd61112, 16'd11767, 16'd11184, 16'd43133, 16'd37791, 16'd49220, 16'd18473, 16'd45965, 16'd27070});
	test_expansion(128'h32b0e6b3b2001489d6e28a11b51e4b0e, {16'd63623, 16'd2755, 16'd23593, 16'd24138, 16'd53154, 16'd32740, 16'd19001, 16'd29238, 16'd53991, 16'd55800, 16'd40707, 16'd23704, 16'd10335, 16'd14696, 16'd9954, 16'd48202, 16'd24727, 16'd65339, 16'd35992, 16'd37459, 16'd22672, 16'd52379, 16'd23792, 16'd44692, 16'd779, 16'd3354});
	test_expansion(128'h008f145a8b415afd31e8c6da5135a2f2, {16'd6932, 16'd62400, 16'd46516, 16'd13571, 16'd36594, 16'd30435, 16'd22329, 16'd22909, 16'd48417, 16'd58564, 16'd53966, 16'd33061, 16'd7914, 16'd59883, 16'd36146, 16'd58620, 16'd139, 16'd52657, 16'd41284, 16'd47726, 16'd49508, 16'd57778, 16'd55578, 16'd36744, 16'd23684, 16'd994});
	test_expansion(128'h49c6b6cb039e72def3d3b327f7deef20, {16'd17762, 16'd13385, 16'd42603, 16'd30458, 16'd16775, 16'd38866, 16'd53916, 16'd26403, 16'd6474, 16'd45803, 16'd58626, 16'd39972, 16'd24186, 16'd43166, 16'd62672, 16'd59413, 16'd49462, 16'd63806, 16'd18330, 16'd6662, 16'd24556, 16'd50390, 16'd60158, 16'd2118, 16'd27196, 16'd50261});
	test_expansion(128'h9b734a156544576e14d27591f8d7244c, {16'd26410, 16'd49940, 16'd43579, 16'd8272, 16'd39089, 16'd36687, 16'd5096, 16'd35547, 16'd14532, 16'd14351, 16'd21529, 16'd7548, 16'd64270, 16'd35645, 16'd50458, 16'd23769, 16'd4599, 16'd14707, 16'd18217, 16'd59554, 16'd62458, 16'd20246, 16'd8301, 16'd2945, 16'd11377, 16'd652});
	test_expansion(128'hf1ab3f9a170609bc30bfd698c5157acd, {16'd56965, 16'd37516, 16'd40385, 16'd49204, 16'd50192, 16'd11931, 16'd36394, 16'd41760, 16'd56796, 16'd4942, 16'd21637, 16'd21356, 16'd58132, 16'd46645, 16'd5054, 16'd54335, 16'd9172, 16'd46581, 16'd46360, 16'd49251, 16'd48534, 16'd29547, 16'd32129, 16'd57331, 16'd61003, 16'd18000});
	test_expansion(128'he6077fd4d042df8ad83c8c17b2b940a4, {16'd15646, 16'd1875, 16'd8965, 16'd15188, 16'd9809, 16'd21284, 16'd44181, 16'd1028, 16'd43721, 16'd54074, 16'd36628, 16'd39369, 16'd23944, 16'd43591, 16'd41871, 16'd30941, 16'd51385, 16'd26568, 16'd45368, 16'd58920, 16'd54094, 16'd50678, 16'd53775, 16'd63039, 16'd40162, 16'd56022});
	test_expansion(128'hfe269b733383dc1b370619a35465d38c, {16'd14210, 16'd19940, 16'd47708, 16'd49961, 16'd20299, 16'd26950, 16'd23609, 16'd15117, 16'd55767, 16'd44640, 16'd43115, 16'd60190, 16'd20877, 16'd15368, 16'd27665, 16'd22747, 16'd64740, 16'd6823, 16'd62880, 16'd62020, 16'd10470, 16'd64801, 16'd32627, 16'd59121, 16'd16076, 16'd7487});
	test_expansion(128'h0d70975f6f34726fbf64fce67d656e36, {16'd45259, 16'd4719, 16'd26449, 16'd4713, 16'd39100, 16'd49531, 16'd58398, 16'd37884, 16'd38782, 16'd22102, 16'd48434, 16'd38709, 16'd62382, 16'd38249, 16'd29368, 16'd55367, 16'd12967, 16'd45650, 16'd61273, 16'd59934, 16'd46970, 16'd21953, 16'd33958, 16'd21726, 16'd32356, 16'd42563});
	test_expansion(128'hd7cb9de881d0d7ea134f20f249276977, {16'd446, 16'd17103, 16'd60097, 16'd41730, 16'd47460, 16'd56384, 16'd11493, 16'd18204, 16'd56786, 16'd41835, 16'd52014, 16'd43485, 16'd9221, 16'd56651, 16'd61762, 16'd21228, 16'd7103, 16'd9619, 16'd5475, 16'd19980, 16'd11804, 16'd49389, 16'd44703, 16'd64725, 16'd15548, 16'd3306});
	test_expansion(128'hab92db8cd60cc9eb19d9e93708d0b1c4, {16'd23235, 16'd55388, 16'd1118, 16'd34090, 16'd45438, 16'd46168, 16'd47336, 16'd10669, 16'd27484, 16'd54848, 16'd31507, 16'd27278, 16'd39967, 16'd65428, 16'd49627, 16'd50290, 16'd8330, 16'd11766, 16'd40716, 16'd7311, 16'd8916, 16'd56743, 16'd38260, 16'd45547, 16'd17276, 16'd42190});
	test_expansion(128'h1ce67856683664302a37ea8b75458dcc, {16'd674, 16'd23690, 16'd43770, 16'd61188, 16'd11955, 16'd1905, 16'd55446, 16'd45943, 16'd62862, 16'd2759, 16'd45058, 16'd64420, 16'd38339, 16'd40008, 16'd15502, 16'd26922, 16'd10709, 16'd20747, 16'd15724, 16'd18241, 16'd35640, 16'd55939, 16'd39942, 16'd60980, 16'd30802, 16'd31152});
	test_expansion(128'h5206a264ec7a1f8ebdc756d0744c4605, {16'd33592, 16'd63606, 16'd39554, 16'd44495, 16'd23771, 16'd36537, 16'd31884, 16'd12019, 16'd8075, 16'd24408, 16'd42871, 16'd6873, 16'd41448, 16'd6670, 16'd24216, 16'd33102, 16'd24466, 16'd27463, 16'd44297, 16'd27954, 16'd48411, 16'd34086, 16'd44887, 16'd46231, 16'd41104, 16'd26757});
	test_expansion(128'h3230b9f054925eaba32d694168090a76, {16'd60865, 16'd11888, 16'd25549, 16'd45651, 16'd58041, 16'd55394, 16'd56138, 16'd13097, 16'd46214, 16'd23876, 16'd39132, 16'd34286, 16'd7256, 16'd35065, 16'd884, 16'd22711, 16'd22744, 16'd56029, 16'd54123, 16'd10512, 16'd43876, 16'd1425, 16'd36980, 16'd25529, 16'd25209, 16'd26134});
	test_expansion(128'h618a24614ba65352d201d31dddf6db61, {16'd45121, 16'd49102, 16'd21645, 16'd41859, 16'd11832, 16'd28268, 16'd32573, 16'd26838, 16'd57700, 16'd22840, 16'd22734, 16'd16877, 16'd55580, 16'd19526, 16'd51135, 16'd23934, 16'd42318, 16'd41886, 16'd21578, 16'd44998, 16'd55343, 16'd46362, 16'd54596, 16'd45992, 16'd715, 16'd65331});
	test_expansion(128'hcd1c983977c72d199b51eed1d2522d67, {16'd35981, 16'd40908, 16'd24925, 16'd7189, 16'd14447, 16'd29085, 16'd10573, 16'd41472, 16'd2385, 16'd43987, 16'd53892, 16'd28982, 16'd63237, 16'd32883, 16'd26600, 16'd55486, 16'd33290, 16'd16707, 16'd14777, 16'd41484, 16'd25224, 16'd18947, 16'd25952, 16'd58597, 16'd33927, 16'd12052});
	test_expansion(128'h32a19cfbc77e605781ebc8c5fc7e42dd, {16'd19821, 16'd49955, 16'd54932, 16'd13742, 16'd40828, 16'd37801, 16'd56378, 16'd28627, 16'd58166, 16'd1542, 16'd55718, 16'd24139, 16'd35266, 16'd897, 16'd58039, 16'd9600, 16'd51726, 16'd40025, 16'd48524, 16'd58114, 16'd12488, 16'd34619, 16'd17072, 16'd41421, 16'd62910, 16'd32163});
	test_expansion(128'hb00f118f46744fa1b716755e8bee55f7, {16'd55112, 16'd52270, 16'd34584, 16'd51967, 16'd46750, 16'd42767, 16'd52829, 16'd2893, 16'd3845, 16'd19485, 16'd38759, 16'd53523, 16'd39449, 16'd62059, 16'd33143, 16'd65238, 16'd26949, 16'd43226, 16'd19725, 16'd7723, 16'd63077, 16'd11934, 16'd28783, 16'd21736, 16'd16172, 16'd13772});
	test_expansion(128'ha38cd1962a3436f832aa11f5f080b59e, {16'd23046, 16'd51537, 16'd53328, 16'd62041, 16'd15182, 16'd10996, 16'd36431, 16'd51590, 16'd40613, 16'd50505, 16'd51790, 16'd50318, 16'd53191, 16'd57495, 16'd8775, 16'd26350, 16'd13260, 16'd12424, 16'd60691, 16'd60539, 16'd20512, 16'd51423, 16'd11286, 16'd42447, 16'd52806, 16'd43396});
	test_expansion(128'h714befcbcf102fa6f29c1a3225b12c35, {16'd62161, 16'd43671, 16'd23392, 16'd22873, 16'd60385, 16'd1968, 16'd8300, 16'd60433, 16'd29638, 16'd38510, 16'd28881, 16'd29359, 16'd32624, 16'd39898, 16'd27889, 16'd42549, 16'd44752, 16'd22106, 16'd48435, 16'd36042, 16'd23412, 16'd11160, 16'd42557, 16'd23252, 16'd63323, 16'd26186});
	test_expansion(128'h0fc28a5ab01bb02d80763455866f7fff, {16'd46088, 16'd51567, 16'd53727, 16'd924, 16'd26588, 16'd55070, 16'd31750, 16'd34563, 16'd5446, 16'd3033, 16'd28245, 16'd21590, 16'd39287, 16'd39374, 16'd35840, 16'd6124, 16'd13671, 16'd49909, 16'd38651, 16'd46049, 16'd46743, 16'd28323, 16'd65346, 16'd36590, 16'd557, 16'd59});
	test_expansion(128'h0ed7aaa8b6576f275ab1cb53d2230c3e, {16'd27513, 16'd7590, 16'd26603, 16'd40072, 16'd39109, 16'd11089, 16'd22737, 16'd48106, 16'd324, 16'd44744, 16'd36572, 16'd12573, 16'd690, 16'd8655, 16'd12358, 16'd23747, 16'd60609, 16'd65504, 16'd40362, 16'd35607, 16'd61166, 16'd41189, 16'd60903, 16'd5568, 16'd39115, 16'd12386});
	test_expansion(128'h37a7306e033fe11ec76392c70f984bfb, {16'd14532, 16'd5147, 16'd46754, 16'd59233, 16'd29798, 16'd47262, 16'd47625, 16'd2902, 16'd25033, 16'd2038, 16'd54662, 16'd38908, 16'd4100, 16'd59586, 16'd40020, 16'd56212, 16'd50026, 16'd56124, 16'd33046, 16'd26772, 16'd40379, 16'd31205, 16'd15398, 16'd16885, 16'd16762, 16'd42189});
	test_expansion(128'h8653394a8d538d4dde916005d9a93ac0, {16'd50402, 16'd42679, 16'd64688, 16'd19961, 16'd1968, 16'd56640, 16'd27846, 16'd371, 16'd14548, 16'd5658, 16'd46151, 16'd47560, 16'd59391, 16'd12939, 16'd36773, 16'd21665, 16'd10220, 16'd135, 16'd61044, 16'd63122, 16'd16118, 16'd63285, 16'd44585, 16'd21738, 16'd49907, 16'd52146});
	test_expansion(128'h86f68ef7594a5835b1d22c90acf7126c, {16'd47240, 16'd29036, 16'd10178, 16'd9022, 16'd45534, 16'd61197, 16'd25225, 16'd49666, 16'd45653, 16'd5298, 16'd34718, 16'd52750, 16'd48666, 16'd26993, 16'd16915, 16'd15995, 16'd64298, 16'd34661, 16'd44446, 16'd62274, 16'd3351, 16'd37326, 16'd3145, 16'd56047, 16'd33712, 16'd32061});
	test_expansion(128'hfa5df4aca4a900131091dd61dfc6e5d3, {16'd3102, 16'd33018, 16'd45489, 16'd32298, 16'd59262, 16'd61916, 16'd50006, 16'd4250, 16'd22991, 16'd43473, 16'd2418, 16'd48289, 16'd62830, 16'd46331, 16'd64843, 16'd32706, 16'd64352, 16'd55882, 16'd42501, 16'd36847, 16'd13057, 16'd1668, 16'd15762, 16'd12947, 16'd22484, 16'd18900});
	test_expansion(128'h6e0754c234bd11005a11d81f99ca6966, {16'd38068, 16'd65440, 16'd48599, 16'd36090, 16'd19031, 16'd43803, 16'd6465, 16'd65445, 16'd11022, 16'd11161, 16'd30468, 16'd10840, 16'd17058, 16'd16629, 16'd21773, 16'd7632, 16'd63718, 16'd42845, 16'd54607, 16'd18722, 16'd58901, 16'd46033, 16'd11351, 16'd58359, 16'd10157, 16'd48187});
	test_expansion(128'h66af144eee7624892b054d0e76defd66, {16'd17843, 16'd52683, 16'd59945, 16'd62021, 16'd195, 16'd132, 16'd31127, 16'd4416, 16'd29690, 16'd34473, 16'd51340, 16'd25502, 16'd34589, 16'd59568, 16'd65005, 16'd42629, 16'd59067, 16'd4441, 16'd54807, 16'd8370, 16'd20589, 16'd24933, 16'd25756, 16'd5952, 16'd1328, 16'd29414});
	test_expansion(128'h275b1d4a85c9c31085eb1387af241f6b, {16'd34359, 16'd36007, 16'd18672, 16'd27235, 16'd19773, 16'd15546, 16'd43822, 16'd34448, 16'd49938, 16'd15154, 16'd44857, 16'd38830, 16'd31698, 16'd30151, 16'd38319, 16'd35459, 16'd6935, 16'd49563, 16'd6531, 16'd58459, 16'd24588, 16'd8704, 16'd7555, 16'd27538, 16'd63210, 16'd31314});
	test_expansion(128'h3810879172b7cc4e7952c94b0ae0a044, {16'd54337, 16'd49583, 16'd39912, 16'd34590, 16'd61295, 16'd43767, 16'd49797, 16'd33507, 16'd15863, 16'd20845, 16'd54798, 16'd51780, 16'd2423, 16'd26165, 16'd44599, 16'd52176, 16'd50101, 16'd36549, 16'd57121, 16'd63306, 16'd21389, 16'd49786, 16'd29886, 16'd9612, 16'd2480, 16'd7520});
	test_expansion(128'h428f53118a4d575d7682f70cbe4bbe4a, {16'd29605, 16'd6602, 16'd19530, 16'd5370, 16'd34332, 16'd31839, 16'd41653, 16'd24686, 16'd56447, 16'd47315, 16'd34619, 16'd25186, 16'd54385, 16'd13668, 16'd64988, 16'd22909, 16'd50393, 16'd1378, 16'd31119, 16'd38048, 16'd21744, 16'd22995, 16'd48253, 16'd33195, 16'd43199, 16'd49263});
	test_expansion(128'h27cc96baf6ae2c11b36be2c9ce4f16e1, {16'd36124, 16'd3940, 16'd29987, 16'd28690, 16'd18087, 16'd19911, 16'd3861, 16'd18611, 16'd22607, 16'd50082, 16'd63740, 16'd61705, 16'd46123, 16'd22735, 16'd61576, 16'd4575, 16'd59925, 16'd60654, 16'd15564, 16'd58743, 16'd33264, 16'd51333, 16'd25578, 16'd24641, 16'd30804, 16'd44633});
	test_expansion(128'haec1063eea9c5f37ab90965099f1fd31, {16'd28853, 16'd16067, 16'd31731, 16'd420, 16'd59557, 16'd34579, 16'd35140, 16'd61041, 16'd5744, 16'd30254, 16'd56014, 16'd3294, 16'd31276, 16'd29460, 16'd58923, 16'd16870, 16'd34024, 16'd60263, 16'd49519, 16'd2700, 16'd3426, 16'd8584, 16'd49643, 16'd45797, 16'd24632, 16'd9673});
	test_expansion(128'he269e743f6e621a299463190fc737219, {16'd37475, 16'd51728, 16'd21980, 16'd39179, 16'd29856, 16'd47004, 16'd15230, 16'd14598, 16'd45980, 16'd36252, 16'd61210, 16'd23944, 16'd36551, 16'd26837, 16'd24203, 16'd26106, 16'd44117, 16'd6691, 16'd18745, 16'd25096, 16'd44896, 16'd20033, 16'd31907, 16'd52611, 16'd58916, 16'd36285});
	test_expansion(128'h30b2864cf8af483d855123487a50492f, {16'd28080, 16'd40087, 16'd600, 16'd53615, 16'd19323, 16'd14617, 16'd37962, 16'd6335, 16'd28827, 16'd19152, 16'd35382, 16'd22511, 16'd6546, 16'd33667, 16'd19034, 16'd36049, 16'd34241, 16'd64016, 16'd26424, 16'd20246, 16'd59020, 16'd57464, 16'd17825, 16'd65117, 16'd58379, 16'd47744});
	test_expansion(128'h87c1b580c4d19c6e36e99bb4edb76f38, {16'd4361, 16'd41513, 16'd25211, 16'd63629, 16'd16283, 16'd20902, 16'd34772, 16'd12362, 16'd44532, 16'd26229, 16'd52738, 16'd9343, 16'd12501, 16'd61772, 16'd55520, 16'd62299, 16'd64262, 16'd47964, 16'd64289, 16'd25699, 16'd3314, 16'd35610, 16'd7530, 16'd39438, 16'd34414, 16'd30169});
	test_expansion(128'hf582af76d226c2b73b2a188a2cb62cc2, {16'd34620, 16'd49094, 16'd33095, 16'd23927, 16'd13008, 16'd49871, 16'd35013, 16'd30098, 16'd59701, 16'd62713, 16'd873, 16'd33546, 16'd38694, 16'd5674, 16'd26717, 16'd44350, 16'd64387, 16'd61333, 16'd23000, 16'd41162, 16'd43946, 16'd59162, 16'd45416, 16'd45037, 16'd7566, 16'd8882});
	test_expansion(128'hd9430026d9f8b473a76b177471549e81, {16'd62050, 16'd4743, 16'd48449, 16'd63079, 16'd40836, 16'd30559, 16'd48441, 16'd20104, 16'd16758, 16'd61210, 16'd10702, 16'd60748, 16'd57018, 16'd43886, 16'd20064, 16'd58516, 16'd50021, 16'd46005, 16'd63174, 16'd55916, 16'd37990, 16'd3238, 16'd3231, 16'd45816, 16'd40693, 16'd57120});
	test_expansion(128'hd2de1f86e3c8a34431d76de604f85b1d, {16'd9909, 16'd17300, 16'd55809, 16'd14594, 16'd42518, 16'd55374, 16'd1642, 16'd58914, 16'd18646, 16'd60344, 16'd45138, 16'd8831, 16'd35262, 16'd59048, 16'd22418, 16'd43747, 16'd12970, 16'd29377, 16'd64466, 16'd43255, 16'd22631, 16'd7842, 16'd38068, 16'd32483, 16'd60506, 16'd8807});
	test_expansion(128'hf2b3c5ecdcf1e61a836820598e1c20ac, {16'd9239, 16'd35796, 16'd46888, 16'd30399, 16'd25017, 16'd32388, 16'd15849, 16'd61159, 16'd65357, 16'd3368, 16'd27265, 16'd22254, 16'd58823, 16'd11019, 16'd8448, 16'd62241, 16'd42924, 16'd6284, 16'd21333, 16'd50787, 16'd60356, 16'd13454, 16'd63866, 16'd14516, 16'd26764, 16'd38034});
	test_expansion(128'hf5ba84b3dfb3c728f0580f403ec0a5f9, {16'd34777, 16'd9918, 16'd23600, 16'd12820, 16'd15805, 16'd24956, 16'd41088, 16'd10502, 16'd25642, 16'd63038, 16'd9513, 16'd45545, 16'd47248, 16'd56719, 16'd50076, 16'd34210, 16'd57530, 16'd8593, 16'd40033, 16'd32974, 16'd31159, 16'd26835, 16'd49985, 16'd49073, 16'd6911, 16'd13719});
	test_expansion(128'h55201461ef6d9fffa5056d6fb84fda50, {16'd28072, 16'd38555, 16'd36613, 16'd15674, 16'd28677, 16'd51555, 16'd9124, 16'd22353, 16'd20277, 16'd30665, 16'd39955, 16'd50296, 16'd29884, 16'd19984, 16'd8976, 16'd8269, 16'd24068, 16'd48523, 16'd2966, 16'd28262, 16'd19642, 16'd62168, 16'd46204, 16'd14214, 16'd59247, 16'd56237});
	test_expansion(128'h5eaf42223ecd30b48d17f2b8346b9f3d, {16'd60277, 16'd4479, 16'd27211, 16'd63521, 16'd30345, 16'd16319, 16'd12552, 16'd35196, 16'd32590, 16'd1620, 16'd1113, 16'd50273, 16'd49849, 16'd2501, 16'd11927, 16'd54823, 16'd10548, 16'd14255, 16'd62769, 16'd42290, 16'd12668, 16'd39296, 16'd27241, 16'd38486, 16'd45575, 16'd25761});
	test_expansion(128'ha2a7f96a27f0903e3e65fa8138103b34, {16'd37583, 16'd23712, 16'd61216, 16'd28858, 16'd56576, 16'd6847, 16'd52858, 16'd3554, 16'd7976, 16'd25945, 16'd13853, 16'd4697, 16'd22235, 16'd16651, 16'd41536, 16'd61016, 16'd32237, 16'd21630, 16'd49198, 16'd12160, 16'd26384, 16'd26547, 16'd16909, 16'd48760, 16'd51050, 16'd31240});
	test_expansion(128'h1cfe54c44c2eba03fb5ff552c2ace061, {16'd17489, 16'd38212, 16'd61391, 16'd54803, 16'd23768, 16'd10130, 16'd62225, 16'd57516, 16'd28955, 16'd28712, 16'd8804, 16'd1847, 16'd43807, 16'd56160, 16'd9436, 16'd1747, 16'd61393, 16'd3553, 16'd36508, 16'd2503, 16'd31085, 16'd63608, 16'd26988, 16'd19993, 16'd21116, 16'd65439});
	test_expansion(128'hfbbfe612918cfc41940cc937ff1f3a71, {16'd39091, 16'd44007, 16'd60916, 16'd18689, 16'd13787, 16'd53097, 16'd50399, 16'd26130, 16'd40004, 16'd3133, 16'd59074, 16'd14284, 16'd5337, 16'd58584, 16'd772, 16'd32894, 16'd41004, 16'd45467, 16'd11831, 16'd64344, 16'd37495, 16'd40151, 16'd64850, 16'd19385, 16'd28456, 16'd47797});
	test_expansion(128'he8e9bd02336a38edcfe3821560c5917f, {16'd4795, 16'd60476, 16'd35816, 16'd5831, 16'd59950, 16'd18396, 16'd21155, 16'd35008, 16'd50630, 16'd12019, 16'd51368, 16'd57673, 16'd8799, 16'd35809, 16'd12792, 16'd430, 16'd58512, 16'd22062, 16'd40431, 16'd42011, 16'd23796, 16'd3331, 16'd34654, 16'd21598, 16'd564, 16'd2552});
	test_expansion(128'hc7c4568fb877d94050431ebfd032481b, {16'd41455, 16'd48371, 16'd47043, 16'd52166, 16'd20180, 16'd44314, 16'd38929, 16'd3102, 16'd11946, 16'd54598, 16'd33519, 16'd38843, 16'd56230, 16'd8923, 16'd8428, 16'd19795, 16'd59590, 16'd46603, 16'd4492, 16'd24564, 16'd11612, 16'd48771, 16'd5063, 16'd55189, 16'd62658, 16'd40672});
	test_expansion(128'h47f160c4dc09f9955908d105562a99c8, {16'd57941, 16'd55783, 16'd49840, 16'd2608, 16'd39940, 16'd12558, 16'd3906, 16'd21069, 16'd17708, 16'd14078, 16'd45590, 16'd11635, 16'd45683, 16'd47390, 16'd9166, 16'd46796, 16'd21874, 16'd12659, 16'd58741, 16'd45668, 16'd3219, 16'd61373, 16'd3386, 16'd55517, 16'd53056, 16'd42864});
	test_expansion(128'h3e99496a06be912fc6e10cb414aa73c1, {16'd31187, 16'd64977, 16'd45870, 16'd65070, 16'd18241, 16'd47769, 16'd52337, 16'd42293, 16'd28238, 16'd41086, 16'd24681, 16'd13298, 16'd48380, 16'd30128, 16'd36468, 16'd24130, 16'd10260, 16'd13059, 16'd30173, 16'd4656, 16'd15836, 16'd21684, 16'd63298, 16'd48873, 16'd38488, 16'd36397});
	test_expansion(128'h4a6da2ded0840e2710656ba673795fec, {16'd30056, 16'd13111, 16'd12151, 16'd44456, 16'd59636, 16'd54256, 16'd46221, 16'd60333, 16'd10390, 16'd50267, 16'd38049, 16'd12779, 16'd15605, 16'd57094, 16'd13061, 16'd18888, 16'd60184, 16'd38130, 16'd17213, 16'd61413, 16'd43020, 16'd51473, 16'd7529, 16'd64625, 16'd51144, 16'd30553});
	test_expansion(128'h441e20d211e25b3b17c1986851499b24, {16'd41942, 16'd53807, 16'd40854, 16'd12044, 16'd15854, 16'd27185, 16'd34506, 16'd27810, 16'd19755, 16'd7400, 16'd22591, 16'd4742, 16'd3026, 16'd64242, 16'd26444, 16'd18927, 16'd28267, 16'd22653, 16'd3260, 16'd43286, 16'd4226, 16'd27068, 16'd48109, 16'd57740, 16'd63143, 16'd21079});
	test_expansion(128'h77ee54b3731bf6023b8a2e61bdac984c, {16'd22738, 16'd29642, 16'd3766, 16'd1617, 16'd39886, 16'd769, 16'd5684, 16'd50815, 16'd42256, 16'd33549, 16'd45247, 16'd23121, 16'd31480, 16'd7025, 16'd32661, 16'd31560, 16'd27270, 16'd51722, 16'd43902, 16'd41801, 16'd1270, 16'd2061, 16'd24895, 16'd17651, 16'd47518, 16'd56445});
	test_expansion(128'h080e61f665d86b1756bb735b12d1f9a2, {16'd28465, 16'd2220, 16'd51952, 16'd58757, 16'd16548, 16'd22733, 16'd52676, 16'd19239, 16'd3216, 16'd4601, 16'd13131, 16'd6956, 16'd18136, 16'd973, 16'd54483, 16'd10496, 16'd38178, 16'd51805, 16'd4349, 16'd33068, 16'd5798, 16'd59621, 16'd4015, 16'd15621, 16'd19047, 16'd23978});
	test_expansion(128'he4ad45bb3c6f5e74b874aebcf8d26bfb, {16'd37481, 16'd11313, 16'd11232, 16'd60251, 16'd36386, 16'd17493, 16'd34248, 16'd3745, 16'd23532, 16'd41749, 16'd817, 16'd64846, 16'd53644, 16'd15040, 16'd57539, 16'd18672, 16'd29198, 16'd4811, 16'd56740, 16'd32468, 16'd46443, 16'd54366, 16'd14244, 16'd60445, 16'd55437, 16'd40061});
	test_expansion(128'h918f6a3ba33b7a4119a33d33f6e2beb7, {16'd65463, 16'd29873, 16'd8147, 16'd17348, 16'd53210, 16'd16699, 16'd20282, 16'd34798, 16'd49960, 16'd564, 16'd23067, 16'd36143, 16'd32026, 16'd44217, 16'd52368, 16'd55781, 16'd11123, 16'd28620, 16'd62175, 16'd43594, 16'd58180, 16'd1219, 16'd30603, 16'd20084, 16'd10311, 16'd26010});
	test_expansion(128'hb8c3b3b4e715e3ae0ec2e35af0a3305e, {16'd21566, 16'd49754, 16'd2693, 16'd8811, 16'd35855, 16'd336, 16'd49566, 16'd54196, 16'd3104, 16'd27850, 16'd17068, 16'd3217, 16'd56766, 16'd46007, 16'd32667, 16'd40962, 16'd9648, 16'd24707, 16'd14480, 16'd24902, 16'd33394, 16'd46499, 16'd11128, 16'd5476, 16'd35200, 16'd28006});
	test_expansion(128'h79f764e45011f84b9df86fc771a2951b, {16'd22315, 16'd44690, 16'd21796, 16'd21849, 16'd28563, 16'd32650, 16'd19859, 16'd7755, 16'd45689, 16'd35872, 16'd12520, 16'd13525, 16'd60414, 16'd24744, 16'd39636, 16'd25970, 16'd16361, 16'd5372, 16'd52801, 16'd55204, 16'd21174, 16'd22228, 16'd7259, 16'd4137, 16'd19790, 16'd4819});
	test_expansion(128'h20c06af5894220c6f5ddf368791aec02, {16'd27678, 16'd57048, 16'd18288, 16'd49696, 16'd13258, 16'd55010, 16'd33301, 16'd8919, 16'd48825, 16'd40207, 16'd4283, 16'd46983, 16'd1139, 16'd7571, 16'd49171, 16'd47589, 16'd57454, 16'd55254, 16'd7120, 16'd56017, 16'd47309, 16'd37200, 16'd16135, 16'd58764, 16'd7881, 16'd25142});
	test_expansion(128'hcd20b564205fe8bb52340ef8b4260817, {16'd64738, 16'd14865, 16'd1983, 16'd46575, 16'd42621, 16'd5140, 16'd33971, 16'd29233, 16'd40825, 16'd19317, 16'd27318, 16'd6551, 16'd18036, 16'd39459, 16'd7199, 16'd60809, 16'd1620, 16'd49389, 16'd61591, 16'd19370, 16'd47350, 16'd20458, 16'd24751, 16'd34810, 16'd59529, 16'd50948});
	test_expansion(128'hfc87e279347f6559e702e0bfc5bacc2f, {16'd11928, 16'd32474, 16'd48490, 16'd57546, 16'd16932, 16'd34104, 16'd46151, 16'd18400, 16'd1844, 16'd45333, 16'd58666, 16'd55419, 16'd29235, 16'd53853, 16'd17132, 16'd31168, 16'd30605, 16'd60420, 16'd26199, 16'd43271, 16'd23401, 16'd41255, 16'd14389, 16'd49642, 16'd19972, 16'd6042});
	test_expansion(128'he33c999b8a4b71ab52ac037ed1e2585f, {16'd36930, 16'd46752, 16'd6920, 16'd6428, 16'd32252, 16'd29890, 16'd46400, 16'd16035, 16'd26149, 16'd60033, 16'd26729, 16'd37539, 16'd4195, 16'd50462, 16'd13123, 16'd29397, 16'd55960, 16'd53369, 16'd18460, 16'd37567, 16'd54423, 16'd17696, 16'd13057, 16'd46704, 16'd1302, 16'd52466});
	test_expansion(128'h68b2994bca4699e356f679ae48d023d3, {16'd54023, 16'd17652, 16'd21881, 16'd38095, 16'd36940, 16'd15110, 16'd7409, 16'd3501, 16'd48748, 16'd4469, 16'd57778, 16'd59584, 16'd7278, 16'd48168, 16'd6589, 16'd38674, 16'd3116, 16'd42387, 16'd60924, 16'd37616, 16'd60799, 16'd6736, 16'd49227, 16'd64819, 16'd64682, 16'd11385});
	test_expansion(128'h63ab51ec54915180135c740b28631ee7, {16'd53040, 16'd62060, 16'd64695, 16'd26278, 16'd63418, 16'd8820, 16'd51010, 16'd20138, 16'd35041, 16'd48407, 16'd57956, 16'd9258, 16'd53179, 16'd18585, 16'd13866, 16'd60036, 16'd47309, 16'd59794, 16'd916, 16'd51267, 16'd2541, 16'd34316, 16'd1365, 16'd30931, 16'd27629, 16'd49845});
	test_expansion(128'h5715c073275c1040295c8bc0e03e2af6, {16'd50768, 16'd24142, 16'd53616, 16'd50095, 16'd2729, 16'd49197, 16'd43055, 16'd49068, 16'd6050, 16'd37665, 16'd50287, 16'd25965, 16'd10682, 16'd56102, 16'd37133, 16'd33005, 16'd37042, 16'd59844, 16'd62200, 16'd53009, 16'd711, 16'd34810, 16'd37939, 16'd50104, 16'd16840, 16'd12906});
	test_expansion(128'hea65fc9a79b42128df567c96957fabec, {16'd38093, 16'd49598, 16'd13148, 16'd39330, 16'd26668, 16'd20407, 16'd23185, 16'd20326, 16'd40560, 16'd30469, 16'd29598, 16'd10992, 16'd38477, 16'd41596, 16'd39430, 16'd19851, 16'd36320, 16'd10101, 16'd24381, 16'd27824, 16'd22881, 16'd32820, 16'd37298, 16'd9509, 16'd30490, 16'd25425});
	test_expansion(128'h86c5c18718c69a916f32ad2911f2c1b4, {16'd29771, 16'd11895, 16'd53533, 16'd30438, 16'd27431, 16'd13621, 16'd1569, 16'd39542, 16'd8358, 16'd50887, 16'd10213, 16'd23795, 16'd3254, 16'd14166, 16'd28072, 16'd53990, 16'd4168, 16'd32811, 16'd64243, 16'd32740, 16'd45564, 16'd53535, 16'd60045, 16'd37852, 16'd47999, 16'd50905});
	test_expansion(128'he4b654860afbbebc88e13e2c18a67c46, {16'd45506, 16'd51541, 16'd46011, 16'd15634, 16'd52104, 16'd22408, 16'd2892, 16'd28697, 16'd12511, 16'd61870, 16'd33276, 16'd29357, 16'd50820, 16'd28517, 16'd22585, 16'd3409, 16'd20046, 16'd44596, 16'd48732, 16'd44511, 16'd21634, 16'd199, 16'd42766, 16'd3542, 16'd58011, 16'd38944});
	test_expansion(128'h369102ee19768b6b0a839386d25c4111, {16'd10884, 16'd15733, 16'd11540, 16'd22066, 16'd51882, 16'd59784, 16'd9696, 16'd27441, 16'd17953, 16'd1234, 16'd44944, 16'd45050, 16'd2532, 16'd10637, 16'd24609, 16'd60152, 16'd18276, 16'd4467, 16'd42794, 16'd27034, 16'd50218, 16'd24746, 16'd36126, 16'd24070, 16'd22576, 16'd60993});
	test_expansion(128'hd689836925397b0c07bb862fb4c6631a, {16'd43148, 16'd17666, 16'd24744, 16'd50960, 16'd32557, 16'd41627, 16'd1366, 16'd40551, 16'd21703, 16'd16971, 16'd62215, 16'd4828, 16'd17970, 16'd54944, 16'd21728, 16'd60651, 16'd6155, 16'd25708, 16'd33072, 16'd30925, 16'd20147, 16'd18193, 16'd3423, 16'd31155, 16'd40063, 16'd37128});
	test_expansion(128'haae915f90b6c0f177602441a2b88001a, {16'd48382, 16'd42116, 16'd26127, 16'd18322, 16'd36511, 16'd49439, 16'd26676, 16'd33891, 16'd47211, 16'd53669, 16'd4261, 16'd21748, 16'd44775, 16'd10144, 16'd52427, 16'd62394, 16'd22020, 16'd31020, 16'd50602, 16'd58525, 16'd13709, 16'd44329, 16'd54263, 16'd57550, 16'd44099, 16'd31094});
	test_expansion(128'hf11176db9e1e5eb7a3850916bf6f04ca, {16'd14928, 16'd14603, 16'd55808, 16'd52778, 16'd33718, 16'd60713, 16'd58878, 16'd24154, 16'd44314, 16'd48244, 16'd48640, 16'd19456, 16'd38157, 16'd19780, 16'd58767, 16'd29432, 16'd28955, 16'd14505, 16'd15076, 16'd48579, 16'd25662, 16'd56179, 16'd51353, 16'd32210, 16'd24623, 16'd16836});
	test_expansion(128'h51288dda0d55b061906956d88d973e90, {16'd41667, 16'd15082, 16'd40436, 16'd24842, 16'd46291, 16'd57331, 16'd6089, 16'd9867, 16'd25840, 16'd22167, 16'd59289, 16'd42414, 16'd50019, 16'd55566, 16'd57104, 16'd50750, 16'd18648, 16'd30877, 16'd41192, 16'd35047, 16'd22298, 16'd18708, 16'd27474, 16'd36081, 16'd31122, 16'd38950});
	test_expansion(128'h0e1ae7ee31bd456aa2d5addf62270694, {16'd21223, 16'd51847, 16'd8484, 16'd54379, 16'd50135, 16'd63044, 16'd52989, 16'd57228, 16'd23374, 16'd64524, 16'd24410, 16'd31931, 16'd47807, 16'd54728, 16'd57508, 16'd2782, 16'd14894, 16'd52287, 16'd61235, 16'd53482, 16'd37675, 16'd65060, 16'd10703, 16'd40983, 16'd8360, 16'd36335});
	test_expansion(128'h1ac1df1ebec0f502589b50b60e25dd99, {16'd48175, 16'd60045, 16'd50271, 16'd34090, 16'd31575, 16'd18851, 16'd12154, 16'd63976, 16'd61209, 16'd9585, 16'd19401, 16'd58780, 16'd43719, 16'd36331, 16'd4566, 16'd3905, 16'd6453, 16'd22622, 16'd44344, 16'd54321, 16'd27686, 16'd21404, 16'd28342, 16'd29734, 16'd63359, 16'd13980});
	test_expansion(128'h83240402ea71e90e47e0104dae932b45, {16'd25847, 16'd2174, 16'd64913, 16'd811, 16'd58359, 16'd4925, 16'd62233, 16'd4692, 16'd16593, 16'd29695, 16'd33592, 16'd31506, 16'd49603, 16'd37015, 16'd11344, 16'd4543, 16'd47211, 16'd14130, 16'd61089, 16'd10758, 16'd23484, 16'd25397, 16'd63155, 16'd47914, 16'd49487, 16'd33139});
	test_expansion(128'h9ce65c6996576018183c72f6698f0860, {16'd478, 16'd16471, 16'd49638, 16'd47301, 16'd5788, 16'd47872, 16'd61256, 16'd22643, 16'd44175, 16'd6896, 16'd3125, 16'd14864, 16'd45042, 16'd63750, 16'd56641, 16'd17723, 16'd28275, 16'd11563, 16'd57054, 16'd16446, 16'd690, 16'd47680, 16'd24680, 16'd27500, 16'd5643, 16'd30743});
	test_expansion(128'ha55e918422466b5f93d087c224c2249f, {16'd49513, 16'd3659, 16'd55085, 16'd56595, 16'd57349, 16'd60064, 16'd38405, 16'd62037, 16'd12579, 16'd16298, 16'd35754, 16'd37627, 16'd21415, 16'd7313, 16'd26536, 16'd60527, 16'd1823, 16'd1524, 16'd27593, 16'd9620, 16'd31624, 16'd62825, 16'd11639, 16'd28043, 16'd8329, 16'd13037});
	test_expansion(128'h15d4e86c19c8a4af89400e79fb98adc9, {16'd8778, 16'd48865, 16'd580, 16'd28596, 16'd52775, 16'd53260, 16'd25657, 16'd40714, 16'd59017, 16'd55692, 16'd16377, 16'd39598, 16'd24920, 16'd26592, 16'd19266, 16'd13395, 16'd58512, 16'd7951, 16'd12101, 16'd53226, 16'd28078, 16'd13840, 16'd42652, 16'd48945, 16'd57706, 16'd28590});
	test_expansion(128'h7833f38899c3832c3e1d46b64a6818ad, {16'd8676, 16'd36404, 16'd59581, 16'd59868, 16'd24734, 16'd54827, 16'd38377, 16'd25331, 16'd47354, 16'd16571, 16'd41852, 16'd20960, 16'd40120, 16'd1724, 16'd54692, 16'd60062, 16'd56284, 16'd17552, 16'd42847, 16'd61294, 16'd5940, 16'd34631, 16'd50519, 16'd48223, 16'd13944, 16'd21371});
	test_expansion(128'hc4a2d8c5380dd2d5e48848e2520cca6e, {16'd33461, 16'd26326, 16'd10688, 16'd34924, 16'd41845, 16'd48459, 16'd48736, 16'd38722, 16'd5323, 16'd63937, 16'd59801, 16'd50398, 16'd13752, 16'd35153, 16'd36289, 16'd27656, 16'd21116, 16'd34917, 16'd33623, 16'd15540, 16'd34755, 16'd16098, 16'd56513, 16'd31682, 16'd65227, 16'd28764});
	test_expansion(128'h56937b5b343d3af2130a5b2d3024e44d, {16'd39360, 16'd13012, 16'd60790, 16'd22101, 16'd47656, 16'd53546, 16'd40872, 16'd19969, 16'd13101, 16'd21870, 16'd13554, 16'd14045, 16'd9747, 16'd37466, 16'd2094, 16'd49789, 16'd27156, 16'd1194, 16'd24673, 16'd30828, 16'd14262, 16'd23004, 16'd19827, 16'd827, 16'd37726, 16'd30154});
	test_expansion(128'h0653b07b9ade75915875033fd47ce9a5, {16'd6885, 16'd1096, 16'd32526, 16'd40999, 16'd45066, 16'd32839, 16'd16273, 16'd28214, 16'd59634, 16'd51797, 16'd26876, 16'd48218, 16'd45990, 16'd8451, 16'd55718, 16'd42734, 16'd55209, 16'd50019, 16'd9928, 16'd912, 16'd7081, 16'd3248, 16'd23369, 16'd3804, 16'd38606, 16'd60541});
	test_expansion(128'h1aefaf34523a37867d93aa1f1fb82440, {16'd63129, 16'd41741, 16'd51199, 16'd49185, 16'd4261, 16'd4818, 16'd4076, 16'd22245, 16'd23693, 16'd61768, 16'd44170, 16'd30894, 16'd5446, 16'd22142, 16'd26900, 16'd63543, 16'd330, 16'd8135, 16'd10804, 16'd16959, 16'd4272, 16'd40538, 16'd38729, 16'd24039, 16'd5583, 16'd15015});
	test_expansion(128'ha1902b75a0ee626cba934011f0346e00, {16'd36316, 16'd17015, 16'd46277, 16'd26060, 16'd55224, 16'd28257, 16'd19120, 16'd16189, 16'd64736, 16'd30479, 16'd41479, 16'd58788, 16'd50168, 16'd21122, 16'd43854, 16'd33622, 16'd14239, 16'd34304, 16'd62051, 16'd24371, 16'd23985, 16'd23963, 16'd3321, 16'd59180, 16'd47034, 16'd13942});
	test_expansion(128'h44345fdb5889bc7861a31d9b92abdd9a, {16'd42021, 16'd55859, 16'd8853, 16'd9763, 16'd1104, 16'd35143, 16'd15771, 16'd59495, 16'd58783, 16'd7452, 16'd34915, 16'd37834, 16'd13280, 16'd26899, 16'd42691, 16'd23228, 16'd54151, 16'd26896, 16'd29707, 16'd58291, 16'd797, 16'd1737, 16'd56665, 16'd29243, 16'd4485, 16'd20422});
	test_expansion(128'h57840b9784be36b7ea56517740378a27, {16'd41642, 16'd13946, 16'd27315, 16'd19384, 16'd17852, 16'd31170, 16'd12730, 16'd3049, 16'd43695, 16'd44602, 16'd25968, 16'd42644, 16'd24591, 16'd32729, 16'd56325, 16'd27299, 16'd56950, 16'd43928, 16'd53553, 16'd25592, 16'd64382, 16'd18586, 16'd50904, 16'd36504, 16'd40777, 16'd8550});
	test_expansion(128'h85339b8841a7862614369d4d4b49331e, {16'd9682, 16'd21000, 16'd59359, 16'd27798, 16'd23236, 16'd37848, 16'd6387, 16'd25665, 16'd65130, 16'd32010, 16'd40453, 16'd24687, 16'd22880, 16'd54773, 16'd2120, 16'd36986, 16'd39696, 16'd38889, 16'd49184, 16'd43051, 16'd1719, 16'd61696, 16'd37146, 16'd5975, 16'd35652, 16'd23229});
	test_expansion(128'hc929e7ca6f4b6f99589959708702b41f, {16'd4983, 16'd56629, 16'd2492, 16'd8011, 16'd6103, 16'd51833, 16'd51619, 16'd64419, 16'd20190, 16'd41462, 16'd36800, 16'd23975, 16'd46564, 16'd10746, 16'd32201, 16'd47295, 16'd28913, 16'd13408, 16'd26427, 16'd5349, 16'd47458, 16'd24726, 16'd20783, 16'd20054, 16'd24058, 16'd31774});
	test_expansion(128'hc0bd503f33da1754f540dd6fdd932ca3, {16'd19167, 16'd63169, 16'd45784, 16'd13808, 16'd47768, 16'd42134, 16'd47266, 16'd40022, 16'd21259, 16'd30005, 16'd23153, 16'd45551, 16'd27449, 16'd14575, 16'd1114, 16'd64121, 16'd24088, 16'd2104, 16'd63347, 16'd56565, 16'd11221, 16'd64461, 16'd2182, 16'd22954, 16'd61812, 16'd29458});
	test_expansion(128'h10426940f54fb14d87ce5c1848a01e1e, {16'd62025, 16'd55188, 16'd33258, 16'd25659, 16'd6370, 16'd46503, 16'd26946, 16'd34975, 16'd25380, 16'd9871, 16'd30608, 16'd10549, 16'd18810, 16'd65361, 16'd60171, 16'd33844, 16'd38411, 16'd22393, 16'd62655, 16'd30835, 16'd25065, 16'd41981, 16'd60389, 16'd52243, 16'd1845, 16'd36921});
	test_expansion(128'h6db1665cb493bc504065502a033f8d5c, {16'd34247, 16'd25699, 16'd38604, 16'd54341, 16'd33528, 16'd33389, 16'd48563, 16'd63128, 16'd19661, 16'd18322, 16'd18455, 16'd878, 16'd17433, 16'd25302, 16'd34405, 16'd25748, 16'd30172, 16'd62448, 16'd21195, 16'd45150, 16'd32144, 16'd36478, 16'd51599, 16'd64093, 16'd41062, 16'd91});
	test_expansion(128'h8ab1f3e2a4a89305c0fea44cddb05016, {16'd18944, 16'd33744, 16'd35778, 16'd47204, 16'd2673, 16'd61985, 16'd31807, 16'd35907, 16'd59965, 16'd16654, 16'd27754, 16'd59762, 16'd48624, 16'd15270, 16'd55679, 16'd36101, 16'd53098, 16'd33701, 16'd63271, 16'd42157, 16'd48719, 16'd29665, 16'd59158, 16'd41655, 16'd999, 16'd20758});
	test_expansion(128'h609131739483adc073425f0af1cc49ad, {16'd56306, 16'd51046, 16'd33084, 16'd34063, 16'd4290, 16'd37267, 16'd21319, 16'd63748, 16'd29357, 16'd20534, 16'd48394, 16'd42810, 16'd44185, 16'd61010, 16'd25063, 16'd55026, 16'd12077, 16'd628, 16'd1625, 16'd12569, 16'd27890, 16'd47190, 16'd17713, 16'd43375, 16'd13576, 16'd44063});
	test_expansion(128'hd0c93c1892b565c5ef68d51b787a9062, {16'd53793, 16'd30147, 16'd57896, 16'd36033, 16'd14993, 16'd63194, 16'd29062, 16'd404, 16'd9554, 16'd45473, 16'd5546, 16'd19523, 16'd39034, 16'd56051, 16'd14368, 16'd36973, 16'd34778, 16'd42509, 16'd8107, 16'd28146, 16'd62053, 16'd28156, 16'd57405, 16'd36090, 16'd22667, 16'd61869});
	test_expansion(128'hf2956e627cf728de806ce7f769e1aaef, {16'd26440, 16'd24190, 16'd25179, 16'd64273, 16'd6080, 16'd3459, 16'd39304, 16'd46640, 16'd7415, 16'd9504, 16'd38485, 16'd41436, 16'd16015, 16'd3431, 16'd62801, 16'd38777, 16'd56052, 16'd34512, 16'd3325, 16'd26293, 16'd53004, 16'd40783, 16'd13589, 16'd16475, 16'd2073, 16'd27082});
	test_expansion(128'h37204c86531353f679430c24a0c3f27d, {16'd6979, 16'd459, 16'd54265, 16'd20560, 16'd7702, 16'd12345, 16'd42077, 16'd55431, 16'd27421, 16'd38376, 16'd52492, 16'd50395, 16'd61628, 16'd53720, 16'd980, 16'd11586, 16'd27207, 16'd49256, 16'd32733, 16'd12332, 16'd40926, 16'd26342, 16'd8119, 16'd23531, 16'd23727, 16'd30824});
	test_expansion(128'h8785862de29e4ae86be5c51527e5b1f3, {16'd35672, 16'd3620, 16'd25894, 16'd34312, 16'd54612, 16'd8097, 16'd42609, 16'd2519, 16'd6859, 16'd23907, 16'd22788, 16'd18825, 16'd6954, 16'd25813, 16'd17769, 16'd5610, 16'd19296, 16'd2361, 16'd18184, 16'd2928, 16'd16230, 16'd8938, 16'd23853, 16'd45069, 16'd42239, 16'd32306});
	test_expansion(128'hcb3778e907de18678657c6e55e8a4ff8, {16'd30055, 16'd227, 16'd9771, 16'd25754, 16'd5663, 16'd36816, 16'd40862, 16'd32841, 16'd4762, 16'd30023, 16'd26657, 16'd12768, 16'd54378, 16'd28082, 16'd5377, 16'd11031, 16'd23697, 16'd8008, 16'd10324, 16'd20247, 16'd20258, 16'd54748, 16'd3834, 16'd47978, 16'd60919, 16'd47878});
	test_expansion(128'hb1aa6e060b1ed2bbf67882660fe4fe3e, {16'd14429, 16'd63825, 16'd48425, 16'd19166, 16'd63879, 16'd53912, 16'd63762, 16'd5707, 16'd61693, 16'd59016, 16'd2893, 16'd42750, 16'd31993, 16'd719, 16'd33654, 16'd57787, 16'd40315, 16'd6550, 16'd28020, 16'd4701, 16'd64189, 16'd18036, 16'd49998, 16'd17635, 16'd14516, 16'd30004});
	test_expansion(128'he2d709dd29219b6e0a63733b8385fcf7, {16'd23583, 16'd38725, 16'd51640, 16'd50590, 16'd54397, 16'd64143, 16'd4977, 16'd31115, 16'd45415, 16'd46628, 16'd14249, 16'd64282, 16'd7734, 16'd55948, 16'd12652, 16'd7978, 16'd49811, 16'd15089, 16'd64041, 16'd3953, 16'd45116, 16'd5604, 16'd39326, 16'd49074, 16'd37251, 16'd54254});
	test_expansion(128'h07c8cb182de3b3d7eb26d0e0882de5ff, {16'd45475, 16'd15623, 16'd51376, 16'd25762, 16'd42188, 16'd2294, 16'd64868, 16'd15741, 16'd31897, 16'd38032, 16'd23263, 16'd48921, 16'd8669, 16'd59854, 16'd30805, 16'd38780, 16'd22769, 16'd64058, 16'd59470, 16'd25543, 16'd11002, 16'd55628, 16'd39839, 16'd36069, 16'd42538, 16'd18348});
	test_expansion(128'h80a3dfce000c7283561b836e2d7501fd, {16'd40076, 16'd17176, 16'd56769, 16'd35158, 16'd40847, 16'd63187, 16'd38269, 16'd50420, 16'd47733, 16'd52947, 16'd24670, 16'd21824, 16'd10986, 16'd31606, 16'd16905, 16'd29186, 16'd7441, 16'd20328, 16'd45537, 16'd52299, 16'd53867, 16'd8427, 16'd33798, 16'd42005, 16'd4561, 16'd34229});
	test_expansion(128'h4f61ad04236f1a1938dc93078a98be03, {16'd51508, 16'd44909, 16'd20072, 16'd30502, 16'd32645, 16'd52556, 16'd41338, 16'd34836, 16'd31126, 16'd64423, 16'd29608, 16'd31787, 16'd46801, 16'd8415, 16'd45350, 16'd34931, 16'd40023, 16'd58169, 16'd7481, 16'd25870, 16'd14434, 16'd42584, 16'd19794, 16'd51876, 16'd36772, 16'd29949});
	test_expansion(128'hb94692dd95c0bf9a16e21accacfe47f7, {16'd6426, 16'd14328, 16'd30768, 16'd18360, 16'd20781, 16'd43240, 16'd55738, 16'd49363, 16'd45192, 16'd10049, 16'd25873, 16'd35539, 16'd18614, 16'd14360, 16'd61262, 16'd26620, 16'd34994, 16'd26234, 16'd31411, 16'd44449, 16'd23602, 16'd5892, 16'd52615, 16'd7757, 16'd33433, 16'd8921});
	test_expansion(128'h051bc68b9991c61a7baf27fbc57553d7, {16'd9405, 16'd49990, 16'd26238, 16'd44669, 16'd61453, 16'd56609, 16'd535, 16'd5356, 16'd13445, 16'd10400, 16'd46816, 16'd50272, 16'd54102, 16'd43639, 16'd27008, 16'd26098, 16'd9726, 16'd39241, 16'd33187, 16'd32075, 16'd10179, 16'd8106, 16'd33285, 16'd38728, 16'd61572, 16'd26175});
	test_expansion(128'hae4ed35056203de58c5f3c8e36c95a3a, {16'd56599, 16'd98, 16'd6846, 16'd11346, 16'd47799, 16'd37015, 16'd51524, 16'd19067, 16'd58536, 16'd65428, 16'd6457, 16'd16009, 16'd10091, 16'd7887, 16'd45060, 16'd5573, 16'd58607, 16'd32638, 16'd56305, 16'd65147, 16'd21609, 16'd34775, 16'd50192, 16'd41210, 16'd59454, 16'd569});
	test_expansion(128'h296ef660ce22a5684c880926fc0a1e49, {16'd22751, 16'd8936, 16'd51214, 16'd31494, 16'd48171, 16'd52624, 16'd58482, 16'd36173, 16'd14337, 16'd933, 16'd20975, 16'd23162, 16'd54315, 16'd36152, 16'd10415, 16'd17584, 16'd52007, 16'd2426, 16'd46780, 16'd37263, 16'd52945, 16'd28721, 16'd25883, 16'd65215, 16'd3839, 16'd430});
	test_expansion(128'h27cf0c81be49accf815dde08647ea16c, {16'd39313, 16'd43460, 16'd50490, 16'd34790, 16'd12214, 16'd27699, 16'd29720, 16'd8261, 16'd38431, 16'd43517, 16'd34303, 16'd64540, 16'd2264, 16'd7882, 16'd24736, 16'd18946, 16'd17486, 16'd41815, 16'd6431, 16'd28201, 16'd34730, 16'd42717, 16'd42258, 16'd3580, 16'd7961, 16'd12572});
	test_expansion(128'h09a31f0c0c3dc42b968a328c803a9343, {16'd19386, 16'd56374, 16'd36244, 16'd42179, 16'd22562, 16'd35713, 16'd52282, 16'd21726, 16'd51057, 16'd15696, 16'd14349, 16'd2791, 16'd3557, 16'd51159, 16'd41234, 16'd50116, 16'd25107, 16'd3136, 16'd36988, 16'd45518, 16'd29666, 16'd40172, 16'd44645, 16'd57564, 16'd34842, 16'd38211});
	test_expansion(128'h0ad290cd6f7bd43e3b9ff32891a7046a, {16'd32438, 16'd26819, 16'd3733, 16'd62828, 16'd33974, 16'd11506, 16'd65194, 16'd40578, 16'd44281, 16'd1582, 16'd33718, 16'd57503, 16'd55104, 16'd19549, 16'd30423, 16'd48147, 16'd35184, 16'd5254, 16'd33000, 16'd28864, 16'd49356, 16'd37788, 16'd2808, 16'd58411, 16'd63586, 16'd48731});
	test_expansion(128'hc8404f33ef7e5005a030954cb520ac49, {16'd44490, 16'd63957, 16'd58438, 16'd25712, 16'd31017, 16'd38917, 16'd31087, 16'd21247, 16'd47376, 16'd56234, 16'd36804, 16'd19701, 16'd50032, 16'd4370, 16'd43120, 16'd9679, 16'd64023, 16'd62573, 16'd18898, 16'd44832, 16'd420, 16'd34571, 16'd36318, 16'd37019, 16'd61318, 16'd9711});
	test_expansion(128'hefd7167198445fc35ec5119ddfb03fa5, {16'd63731, 16'd18267, 16'd61986, 16'd64529, 16'd30018, 16'd30709, 16'd21932, 16'd45403, 16'd63962, 16'd19384, 16'd38928, 16'd5512, 16'd63483, 16'd61476, 16'd10736, 16'd47373, 16'd41966, 16'd14115, 16'd26165, 16'd49056, 16'd55574, 16'd44390, 16'd36848, 16'd17443, 16'd21571, 16'd9384});
	test_expansion(128'h63d3cd80f1bc1b78eba1bccfb87739d6, {16'd60514, 16'd44188, 16'd15147, 16'd32959, 16'd33545, 16'd37473, 16'd60370, 16'd53686, 16'd64341, 16'd65482, 16'd63435, 16'd20799, 16'd47684, 16'd32771, 16'd6336, 16'd49167, 16'd5723, 16'd38625, 16'd25625, 16'd16661, 16'd15390, 16'd16932, 16'd35043, 16'd51263, 16'd21757, 16'd32975});
	test_expansion(128'h5d4fd546d3b82f2b22dd671e997f2ccc, {16'd7570, 16'd17004, 16'd42008, 16'd64438, 16'd4194, 16'd33725, 16'd58719, 16'd42998, 16'd41967, 16'd57476, 16'd29942, 16'd50229, 16'd63101, 16'd55022, 16'd28733, 16'd57025, 16'd13182, 16'd59480, 16'd42692, 16'd22111, 16'd10456, 16'd58262, 16'd14859, 16'd40507, 16'd43588, 16'd14481});
	test_expansion(128'h6e2affb92a7b786c45d938877aa6aaf4, {16'd2773, 16'd2779, 16'd15768, 16'd40595, 16'd21774, 16'd17651, 16'd57853, 16'd37935, 16'd63937, 16'd36063, 16'd1268, 16'd17313, 16'd64523, 16'd32985, 16'd14475, 16'd22759, 16'd12206, 16'd1374, 16'd4673, 16'd60248, 16'd49461, 16'd5318, 16'd3651, 16'd11307, 16'd33847, 16'd27317});
	test_expansion(128'ha19f4ed0e15c714f2954df12f7418db0, {16'd6838, 16'd36814, 16'd38165, 16'd44957, 16'd48622, 16'd23879, 16'd28523, 16'd10967, 16'd50844, 16'd3258, 16'd494, 16'd48044, 16'd17999, 16'd17253, 16'd51443, 16'd47428, 16'd45532, 16'd27233, 16'd50835, 16'd59855, 16'd57106, 16'd14043, 16'd50385, 16'd32040, 16'd46038, 16'd42587});
	test_expansion(128'h2bb338a08c2c6e652847a130b80bdbc1, {16'd39484, 16'd14448, 16'd15430, 16'd4814, 16'd63806, 16'd35258, 16'd24678, 16'd8714, 16'd20155, 16'd9921, 16'd26412, 16'd13407, 16'd25987, 16'd31654, 16'd22441, 16'd19005, 16'd25347, 16'd183, 16'd13251, 16'd16558, 16'd54514, 16'd33044, 16'd5507, 16'd49070, 16'd59943, 16'd22266});
	test_expansion(128'h1c6fce82c7a008c31e6a934dd1cbbc08, {16'd19950, 16'd60984, 16'd14292, 16'd47983, 16'd25862, 16'd51872, 16'd30342, 16'd32116, 16'd50253, 16'd15013, 16'd40526, 16'd4713, 16'd20117, 16'd1442, 16'd44432, 16'd57182, 16'd21922, 16'd38910, 16'd12678, 16'd58597, 16'd19752, 16'd52695, 16'd39351, 16'd39474, 16'd43276, 16'd26624});
	test_expansion(128'h75e7cbbec11028ce4a96a163ad30f33c, {16'd572, 16'd17159, 16'd12717, 16'd29645, 16'd58529, 16'd29453, 16'd5974, 16'd17884, 16'd63371, 16'd12749, 16'd63232, 16'd28792, 16'd39342, 16'd29818, 16'd7665, 16'd39864, 16'd22544, 16'd53821, 16'd3476, 16'd59257, 16'd60399, 16'd35830, 16'd8926, 16'd50390, 16'd19057, 16'd8607});
	test_expansion(128'hb25d44492401d42d1af4ae477041c10b, {16'd48205, 16'd59604, 16'd30083, 16'd1764, 16'd28780, 16'd25902, 16'd23966, 16'd37743, 16'd3468, 16'd17157, 16'd51172, 16'd15800, 16'd4751, 16'd30194, 16'd39698, 16'd38573, 16'd16868, 16'd32436, 16'd11220, 16'd57225, 16'd41664, 16'd19761, 16'd51251, 16'd51120, 16'd61169, 16'd237});
	test_expansion(128'h2dfbdd3bb1e767553e5a0e7065255740, {16'd48695, 16'd53856, 16'd9603, 16'd30877, 16'd29236, 16'd36700, 16'd7613, 16'd3943, 16'd18928, 16'd60803, 16'd57205, 16'd41918, 16'd37437, 16'd4124, 16'd1484, 16'd62194, 16'd55537, 16'd42165, 16'd49114, 16'd52388, 16'd62350, 16'd62043, 16'd41053, 16'd27555, 16'd10104, 16'd10332});
	test_expansion(128'hfe4ee7645afd2d86773cc6d515a86c2d, {16'd11395, 16'd7515, 16'd9910, 16'd13641, 16'd660, 16'd3876, 16'd29388, 16'd17054, 16'd29634, 16'd649, 16'd36733, 16'd53200, 16'd2100, 16'd54690, 16'd6172, 16'd41416, 16'd3033, 16'd23145, 16'd58259, 16'd33265, 16'd48466, 16'd4080, 16'd10090, 16'd8855, 16'd48212, 16'd36382});
	test_expansion(128'hbdd37134aec2bd6aa62a980115532707, {16'd19693, 16'd44635, 16'd16770, 16'd12810, 16'd59012, 16'd18318, 16'd57994, 16'd2878, 16'd61790, 16'd9113, 16'd40034, 16'd17687, 16'd46219, 16'd49946, 16'd56554, 16'd9792, 16'd29253, 16'd34058, 16'd14845, 16'd1954, 16'd47976, 16'd10281, 16'd62009, 16'd46958, 16'd47468, 16'd26849});
	test_expansion(128'h09f92eb69120ec480c0cdf7cb7ebbea5, {16'd45668, 16'd62334, 16'd16060, 16'd43251, 16'd27248, 16'd18530, 16'd28492, 16'd48673, 16'd58976, 16'd13262, 16'd27531, 16'd43115, 16'd16325, 16'd40316, 16'd34061, 16'd6312, 16'd49878, 16'd52733, 16'd49887, 16'd37491, 16'd25130, 16'd55961, 16'd54703, 16'd49441, 16'd46167, 16'd29607});
	test_expansion(128'h63a66f21604648cd1c9a8629b066092b, {16'd16392, 16'd61679, 16'd44342, 16'd43898, 16'd42856, 16'd5391, 16'd53907, 16'd32145, 16'd47110, 16'd1650, 16'd44670, 16'd35183, 16'd37515, 16'd45534, 16'd62677, 16'd16503, 16'd13446, 16'd7304, 16'd38349, 16'd62205, 16'd53104, 16'd17208, 16'd33669, 16'd14112, 16'd48190, 16'd31482});
	test_expansion(128'h6fcb40e222050bf8cac8740c38666942, {16'd59526, 16'd34741, 16'd8981, 16'd15390, 16'd59479, 16'd28910, 16'd28125, 16'd63905, 16'd38295, 16'd63863, 16'd65336, 16'd35504, 16'd20881, 16'd37045, 16'd60266, 16'd21016, 16'd13754, 16'd51885, 16'd818, 16'd31793, 16'd17379, 16'd39317, 16'd18492, 16'd26199, 16'd27404, 16'd6621});
	test_expansion(128'h4f6eeb43086b483e98723012a94232f0, {16'd21783, 16'd64610, 16'd31872, 16'd3301, 16'd2903, 16'd55951, 16'd29070, 16'd5094, 16'd17114, 16'd21246, 16'd36375, 16'd22262, 16'd65491, 16'd5585, 16'd43239, 16'd53676, 16'd47338, 16'd51877, 16'd759, 16'd17244, 16'd28927, 16'd882, 16'd61096, 16'd4167, 16'd34920, 16'd7584});
	test_expansion(128'h6b248714dcb46393631493e6e89422fa, {16'd40160, 16'd12553, 16'd28184, 16'd41402, 16'd52679, 16'd3764, 16'd36280, 16'd29338, 16'd15454, 16'd22604, 16'd12115, 16'd52820, 16'd43350, 16'd8990, 16'd5499, 16'd58264, 16'd41050, 16'd40755, 16'd39642, 16'd24326, 16'd24076, 16'd59494, 16'd14398, 16'd13869, 16'd36027, 16'd59386});
	test_expansion(128'he32b9fc5ae7f6d1d1dd9f32c59bf86d4, {16'd58706, 16'd3976, 16'd58540, 16'd17837, 16'd1791, 16'd38064, 16'd37810, 16'd63130, 16'd8644, 16'd57930, 16'd931, 16'd33632, 16'd61045, 16'd60988, 16'd52243, 16'd28970, 16'd36864, 16'd26472, 16'd27527, 16'd47726, 16'd38053, 16'd64466, 16'd29669, 16'd24761, 16'd33349, 16'd11830});
	test_expansion(128'he6ef5177939d69852a6d8a7af1653df6, {16'd30542, 16'd10606, 16'd39768, 16'd20899, 16'd56249, 16'd15689, 16'd24025, 16'd7896, 16'd16539, 16'd26857, 16'd62696, 16'd32553, 16'd3044, 16'd61344, 16'd22902, 16'd39816, 16'd62559, 16'd20196, 16'd61567, 16'd47842, 16'd24398, 16'd15609, 16'd57502, 16'd52229, 16'd60609, 16'd5937});
	test_expansion(128'hf42183879d761935ccd6f13cf0fed73f, {16'd45233, 16'd36737, 16'd46727, 16'd53993, 16'd27316, 16'd24448, 16'd39901, 16'd6198, 16'd7993, 16'd56200, 16'd7458, 16'd56208, 16'd38417, 16'd11683, 16'd45346, 16'd13728, 16'd36423, 16'd36957, 16'd44909, 16'd14838, 16'd49734, 16'd37010, 16'd45031, 16'd10155, 16'd62746, 16'd31403});
	test_expansion(128'h79c584737e4545b47c10fdd69f5e55b8, {16'd50895, 16'd23886, 16'd40445, 16'd3971, 16'd48039, 16'd27652, 16'd37894, 16'd33744, 16'd31369, 16'd2777, 16'd61318, 16'd26357, 16'd44199, 16'd57215, 16'd42029, 16'd53278, 16'd3684, 16'd44448, 16'd46618, 16'd34150, 16'd55332, 16'd45099, 16'd39941, 16'd5390, 16'd14477, 16'd23849});
	test_expansion(128'h9276e2b47bb2562ae17be56805c09eea, {16'd36185, 16'd3988, 16'd56632, 16'd19935, 16'd59850, 16'd7908, 16'd7116, 16'd54088, 16'd34597, 16'd1257, 16'd45808, 16'd702, 16'd33598, 16'd7491, 16'd4332, 16'd2538, 16'd40083, 16'd25620, 16'd6403, 16'd49882, 16'd33915, 16'd33118, 16'd47263, 16'd33934, 16'd28480, 16'd54390});
	test_expansion(128'h2ebf2e8df65ff1464f43b5986e900221, {16'd5423, 16'd58207, 16'd10035, 16'd43672, 16'd62818, 16'd45995, 16'd50648, 16'd44187, 16'd52312, 16'd56829, 16'd29806, 16'd15964, 16'd28291, 16'd35430, 16'd59945, 16'd39146, 16'd34016, 16'd15325, 16'd38893, 16'd12024, 16'd44005, 16'd54089, 16'd37339, 16'd60453, 16'd44945, 16'd38952});
	test_expansion(128'h3c69f8c4a2047536ba97a20e0d687f9e, {16'd43170, 16'd5035, 16'd18672, 16'd49522, 16'd50717, 16'd62072, 16'd2618, 16'd15097, 16'd62777, 16'd36504, 16'd3324, 16'd64652, 16'd1258, 16'd9951, 16'd40317, 16'd31759, 16'd48846, 16'd60129, 16'd39056, 16'd20138, 16'd1467, 16'd25236, 16'd22373, 16'd15251, 16'd44945, 16'd27196});
	test_expansion(128'hed437d8b5130e07cd7b3577f241133dc, {16'd50078, 16'd28954, 16'd47160, 16'd21664, 16'd62440, 16'd32425, 16'd10014, 16'd5169, 16'd63730, 16'd16389, 16'd5044, 16'd15277, 16'd26310, 16'd24872, 16'd6906, 16'd10799, 16'd27518, 16'd32178, 16'd57192, 16'd25176, 16'd57865, 16'd43204, 16'd47811, 16'd61793, 16'd50517, 16'd20417});
	test_expansion(128'h56fb39e5b662bf55945833b8101eb044, {16'd17378, 16'd9153, 16'd18031, 16'd30099, 16'd26382, 16'd8114, 16'd31650, 16'd41097, 16'd51624, 16'd24334, 16'd23715, 16'd48089, 16'd34512, 16'd41623, 16'd38811, 16'd49978, 16'd4451, 16'd20059, 16'd41950, 16'd8317, 16'd20568, 16'd49046, 16'd61309, 16'd15215, 16'd20095, 16'd63739});
	test_expansion(128'h8132be79223d87ead18617aa601295d3, {16'd28967, 16'd44003, 16'd28810, 16'd4800, 16'd28206, 16'd17750, 16'd37304, 16'd11269, 16'd52234, 16'd20384, 16'd12369, 16'd12318, 16'd38553, 16'd11412, 16'd18281, 16'd57976, 16'd30177, 16'd41129, 16'd60666, 16'd8145, 16'd58917, 16'd54378, 16'd11071, 16'd21613, 16'd30869, 16'd20421});
	test_expansion(128'h5196b856f8bf0f3e4fe473a0ab9ecc38, {16'd42477, 16'd23123, 16'd10691, 16'd40907, 16'd25255, 16'd44889, 16'd39511, 16'd13268, 16'd26813, 16'd21954, 16'd10687, 16'd985, 16'd47085, 16'd57347, 16'd54819, 16'd24029, 16'd49199, 16'd41938, 16'd41182, 16'd16242, 16'd14033, 16'd65364, 16'd10217, 16'd4289, 16'd16396, 16'd42293});
	test_expansion(128'he08f1686a4ea51841369414b324ca29e, {16'd65380, 16'd15809, 16'd1593, 16'd41014, 16'd56727, 16'd23963, 16'd51550, 16'd64902, 16'd50190, 16'd27013, 16'd23998, 16'd14270, 16'd32632, 16'd56560, 16'd35481, 16'd19150, 16'd45611, 16'd60461, 16'd14695, 16'd49811, 16'd49314, 16'd5945, 16'd5333, 16'd47765, 16'd47885, 16'd37916});
	test_expansion(128'hb3afab8e9189625237670dee298eb85c, {16'd64872, 16'd59345, 16'd1450, 16'd10089, 16'd57435, 16'd18540, 16'd4436, 16'd35133, 16'd65008, 16'd64299, 16'd9427, 16'd49253, 16'd10543, 16'd23108, 16'd9498, 16'd41093, 16'd42097, 16'd53315, 16'd43233, 16'd55264, 16'd2017, 16'd53170, 16'd2923, 16'd8685, 16'd10844, 16'd41452});
	test_expansion(128'he8b2457733bf86805ac4d4c996281cc1, {16'd16836, 16'd23060, 16'd30175, 16'd42293, 16'd39249, 16'd438, 16'd57326, 16'd18016, 16'd644, 16'd20145, 16'd7623, 16'd32090, 16'd37312, 16'd13351, 16'd24664, 16'd7586, 16'd14044, 16'd49851, 16'd62548, 16'd44537, 16'd19771, 16'd61264, 16'd33495, 16'd3953, 16'd57752, 16'd24931});
	test_expansion(128'h52a8517c99d8844df325b0ff64521815, {16'd49650, 16'd40364, 16'd1709, 16'd50662, 16'd48893, 16'd45761, 16'd29226, 16'd17413, 16'd8200, 16'd39168, 16'd50935, 16'd12692, 16'd34132, 16'd2669, 16'd42300, 16'd1212, 16'd17464, 16'd45395, 16'd62393, 16'd46209, 16'd13063, 16'd53652, 16'd51061, 16'd39942, 16'd8956, 16'd1902});
	test_expansion(128'h9a896813b69bac697d605564ad41fbe4, {16'd52985, 16'd26978, 16'd12734, 16'd61491, 16'd64873, 16'd11840, 16'd55817, 16'd14794, 16'd18560, 16'd44358, 16'd60643, 16'd3797, 16'd26349, 16'd58954, 16'd23798, 16'd44601, 16'd59668, 16'd43377, 16'd51754, 16'd30508, 16'd61497, 16'd11615, 16'd52393, 16'd27111, 16'd38072, 16'd11463});
	test_expansion(128'he59b40c65d5014bcecc6e38d2151302a, {16'd6605, 16'd47322, 16'd7057, 16'd10518, 16'd2453, 16'd44723, 16'd35295, 16'd18210, 16'd6049, 16'd20594, 16'd16397, 16'd9251, 16'd34428, 16'd6992, 16'd14496, 16'd11814, 16'd30080, 16'd43312, 16'd3023, 16'd36408, 16'd52829, 16'd4316, 16'd47465, 16'd56653, 16'd55293, 16'd25289});
	test_expansion(128'hf243e0273a97e181c7447944bd7d7c7c, {16'd1502, 16'd58076, 16'd65302, 16'd12116, 16'd24220, 16'd16631, 16'd10814, 16'd41303, 16'd60062, 16'd7670, 16'd51523, 16'd9988, 16'd2828, 16'd33316, 16'd22251, 16'd25891, 16'd10339, 16'd62365, 16'd53894, 16'd16337, 16'd30984, 16'd17732, 16'd38255, 16'd64035, 16'd32935, 16'd56285});
	test_expansion(128'h115c0a8421ae34b6d01c5bec411d7b10, {16'd12501, 16'd23116, 16'd65067, 16'd40028, 16'd26931, 16'd9590, 16'd33475, 16'd2540, 16'd47935, 16'd9686, 16'd5489, 16'd25179, 16'd31318, 16'd46316, 16'd51536, 16'd27826, 16'd13780, 16'd24085, 16'd17857, 16'd50088, 16'd14276, 16'd25458, 16'd3122, 16'd1525, 16'd5493, 16'd41274});
	test_expansion(128'h527cb16a8746867d289d253bbd8866f1, {16'd39313, 16'd26823, 16'd33462, 16'd25077, 16'd33395, 16'd2619, 16'd33376, 16'd60869, 16'd7858, 16'd55836, 16'd25971, 16'd9207, 16'd58837, 16'd14683, 16'd56357, 16'd12330, 16'd30605, 16'd55565, 16'd22551, 16'd9620, 16'd57456, 16'd45704, 16'd58079, 16'd27554, 16'd55446, 16'd16356});
	test_expansion(128'h4a36852b3092238f74b418a92336d16c, {16'd31319, 16'd38031, 16'd20615, 16'd41799, 16'd4420, 16'd58624, 16'd44339, 16'd15488, 16'd31804, 16'd9257, 16'd29850, 16'd4406, 16'd14711, 16'd43923, 16'd58027, 16'd34351, 16'd41642, 16'd17226, 16'd18295, 16'd46741, 16'd54651, 16'd38061, 16'd52787, 16'd64683, 16'd55325, 16'd8504});
	test_expansion(128'h7ae7b2523590bdd04cba5322bdbe0b35, {16'd64467, 16'd28907, 16'd36165, 16'd55066, 16'd24804, 16'd15162, 16'd18126, 16'd23687, 16'd60248, 16'd47608, 16'd45381, 16'd6933, 16'd32197, 16'd16441, 16'd33830, 16'd38695, 16'd56785, 16'd30745, 16'd53113, 16'd51891, 16'd3249, 16'd8922, 16'd8019, 16'd5594, 16'd52324, 16'd26811});
	test_expansion(128'h3a4793eefbf092c127aaa60a536f44b8, {16'd22529, 16'd41599, 16'd3737, 16'd52276, 16'd52209, 16'd11217, 16'd44889, 16'd18251, 16'd36845, 16'd45532, 16'd13158, 16'd19956, 16'd18569, 16'd14983, 16'd7439, 16'd45279, 16'd1691, 16'd5719, 16'd48916, 16'd13323, 16'd10515, 16'd13797, 16'd21153, 16'd45482, 16'd52677, 16'd5207});
	test_expansion(128'h4962ad26d411b765dc7670bf8658d9b6, {16'd38679, 16'd42723, 16'd27185, 16'd40448, 16'd17958, 16'd54034, 16'd41076, 16'd18301, 16'd25585, 16'd21420, 16'd50543, 16'd55250, 16'd16061, 16'd50454, 16'd45233, 16'd43287, 16'd17358, 16'd45237, 16'd13882, 16'd49127, 16'd20946, 16'd34744, 16'd58014, 16'd57032, 16'd50006, 16'd12776});
	test_expansion(128'h80c75c492ddb2eb1dfd37a8f9ec9eef6, {16'd26684, 16'd14861, 16'd2612, 16'd4376, 16'd21124, 16'd24653, 16'd57252, 16'd18912, 16'd19903, 16'd18395, 16'd58057, 16'd20080, 16'd56972, 16'd47743, 16'd14197, 16'd6637, 16'd51564, 16'd15982, 16'd20611, 16'd26422, 16'd2505, 16'd55994, 16'd50361, 16'd12158, 16'd49179, 16'd18665});
	test_expansion(128'h2404765ac3863e7565e2f6c79c8a711b, {16'd50596, 16'd51470, 16'd45822, 16'd45295, 16'd10351, 16'd62743, 16'd17561, 16'd30922, 16'd40406, 16'd17961, 16'd15908, 16'd20916, 16'd18752, 16'd4736, 16'd1097, 16'd36340, 16'd7075, 16'd14453, 16'd50415, 16'd19828, 16'd30079, 16'd22475, 16'd54825, 16'd40938, 16'd37783, 16'd10374});
	test_expansion(128'hef7def1f782046d8376939a4db179335, {16'd60892, 16'd34469, 16'd3081, 16'd11781, 16'd48113, 16'd28467, 16'd39428, 16'd8070, 16'd56926, 16'd47407, 16'd16460, 16'd51008, 16'd50318, 16'd16463, 16'd10240, 16'd15753, 16'd47732, 16'd42833, 16'd52604, 16'd16958, 16'd38354, 16'd12432, 16'd17045, 16'd23127, 16'd39306, 16'd56671});
	test_expansion(128'h058a37bbc0c120218942e1eb24c89a6a, {16'd54913, 16'd16235, 16'd58338, 16'd8241, 16'd61266, 16'd48028, 16'd3213, 16'd57339, 16'd29491, 16'd54225, 16'd22336, 16'd28616, 16'd38991, 16'd10845, 16'd109, 16'd48527, 16'd33683, 16'd28422, 16'd29403, 16'd6901, 16'd63748, 16'd37667, 16'd53517, 16'd64240, 16'd14452, 16'd28476});
	test_expansion(128'h6e127bcacadd4082facb8ffb2d8de15b, {16'd17952, 16'd17906, 16'd30310, 16'd5525, 16'd9005, 16'd18473, 16'd55805, 16'd3130, 16'd49666, 16'd10159, 16'd6997, 16'd11936, 16'd41053, 16'd49739, 16'd491, 16'd7164, 16'd18668, 16'd21719, 16'd33288, 16'd2089, 16'd15824, 16'd48405, 16'd42254, 16'd3722, 16'd50851, 16'd56481});
	test_expansion(128'hfa947630040b85322e10ac3fee937085, {16'd8184, 16'd26504, 16'd54706, 16'd5620, 16'd47475, 16'd35603, 16'd44702, 16'd34248, 16'd30562, 16'd4504, 16'd31799, 16'd61471, 16'd60042, 16'd28343, 16'd18308, 16'd20859, 16'd35734, 16'd50267, 16'd12621, 16'd12083, 16'd41080, 16'd56901, 16'd20600, 16'd50494, 16'd49803, 16'd44906});
	test_expansion(128'h271164f3be626d3ea24d76ae92396cdf, {16'd47698, 16'd59431, 16'd36657, 16'd6950, 16'd38308, 16'd24795, 16'd65051, 16'd6378, 16'd5593, 16'd53062, 16'd13659, 16'd35965, 16'd51808, 16'd33166, 16'd38036, 16'd58301, 16'd58107, 16'd51455, 16'd30089, 16'd54535, 16'd35513, 16'd36120, 16'd28134, 16'd9031, 16'd7087, 16'd58580});
	test_expansion(128'hb3f56accdd14c8a0f5aa5670ef37e423, {16'd20146, 16'd14665, 16'd24427, 16'd4063, 16'd48896, 16'd48089, 16'd8125, 16'd40220, 16'd21902, 16'd55824, 16'd27899, 16'd47928, 16'd4467, 16'd8652, 16'd33803, 16'd8982, 16'd57761, 16'd42482, 16'd47536, 16'd5896, 16'd51483, 16'd29787, 16'd6210, 16'd16683, 16'd57266, 16'd39816});
	test_expansion(128'h8f2171f6dd1328ad6414a744086e8228, {16'd25901, 16'd38457, 16'd44637, 16'd47930, 16'd42866, 16'd30047, 16'd59309, 16'd20900, 16'd32957, 16'd46933, 16'd53662, 16'd18521, 16'd18618, 16'd51494, 16'd30846, 16'd57477, 16'd61355, 16'd52334, 16'd29806, 16'd63497, 16'd45465, 16'd52134, 16'd54671, 16'd19559, 16'd28910, 16'd14919});
	test_expansion(128'hb2b115fa9d7a206301a46b6ffabdc17a, {16'd59176, 16'd30185, 16'd36347, 16'd49722, 16'd46954, 16'd52577, 16'd45234, 16'd28071, 16'd28442, 16'd16130, 16'd51982, 16'd17005, 16'd41151, 16'd39283, 16'd20011, 16'd42042, 16'd224, 16'd1975, 16'd51612, 16'd25031, 16'd34952, 16'd53470, 16'd7859, 16'd35868, 16'd26886, 16'd55564});
	test_expansion(128'h5e52c4d9327f13cb522e308bb2f88a69, {16'd31517, 16'd7300, 16'd10038, 16'd688, 16'd17844, 16'd16467, 16'd37218, 16'd28939, 16'd27001, 16'd19614, 16'd61230, 16'd64525, 16'd59753, 16'd2027, 16'd37771, 16'd20955, 16'd60006, 16'd21692, 16'd11631, 16'd3326, 16'd35389, 16'd57145, 16'd63931, 16'd1149, 16'd1972, 16'd25630});
	test_expansion(128'haba87429226ed45bd80c68365ce54cf7, {16'd28930, 16'd2742, 16'd22402, 16'd7500, 16'd18203, 16'd36928, 16'd59317, 16'd2461, 16'd15185, 16'd64082, 16'd13253, 16'd23092, 16'd19818, 16'd35378, 16'd27056, 16'd64206, 16'd60291, 16'd48887, 16'd59311, 16'd46475, 16'd306, 16'd2633, 16'd37772, 16'd43133, 16'd64683, 16'd55171});
	test_expansion(128'ha47c4fb7f82eab40a3e26a3d3f6fffea, {16'd57642, 16'd5873, 16'd31796, 16'd21618, 16'd4521, 16'd37986, 16'd49655, 16'd64069, 16'd63860, 16'd1582, 16'd1042, 16'd65334, 16'd61807, 16'd26742, 16'd63192, 16'd53624, 16'd21252, 16'd30204, 16'd49575, 16'd63064, 16'd41778, 16'd64717, 16'd12121, 16'd57975, 16'd4818, 16'd86});
	test_expansion(128'h0a0316ebc2b7f5a8dfde3188a1806ffb, {16'd18020, 16'd26571, 16'd36242, 16'd32081, 16'd29861, 16'd24596, 16'd46592, 16'd28321, 16'd51141, 16'd15720, 16'd17597, 16'd13961, 16'd45171, 16'd17620, 16'd54988, 16'd8691, 16'd40239, 16'd1028, 16'd36869, 16'd49996, 16'd41878, 16'd57328, 16'd52144, 16'd47919, 16'd33590, 16'd60895});
	test_expansion(128'h1120f9a4e12441e688a8a3316d336d80, {16'd6125, 16'd15166, 16'd214, 16'd25587, 16'd50926, 16'd4864, 16'd47788, 16'd31564, 16'd55962, 16'd23364, 16'd15464, 16'd64981, 16'd45835, 16'd47886, 16'd43444, 16'd50787, 16'd49425, 16'd13929, 16'd19525, 16'd15205, 16'd60311, 16'd53720, 16'd63329, 16'd44524, 16'd16094, 16'd35762});
	test_expansion(128'h79bdcb01f866cea48e5288a335b4e3c0, {16'd31902, 16'd1268, 16'd34040, 16'd36919, 16'd59125, 16'd46728, 16'd46329, 16'd49630, 16'd512, 16'd3517, 16'd8781, 16'd37042, 16'd38552, 16'd22906, 16'd45857, 16'd16364, 16'd5342, 16'd54640, 16'd50155, 16'd57540, 16'd27086, 16'd3469, 16'd37295, 16'd16095, 16'd34997, 16'd46637});
	test_expansion(128'h51e04521b42695d359818b6afaea4e1d, {16'd49952, 16'd31262, 16'd52392, 16'd8660, 16'd41973, 16'd5812, 16'd39819, 16'd10834, 16'd63419, 16'd14023, 16'd7319, 16'd40674, 16'd38033, 16'd37898, 16'd37564, 16'd17871, 16'd61772, 16'd8247, 16'd16407, 16'd65300, 16'd18894, 16'd384, 16'd11170, 16'd61167, 16'd37511, 16'd40235});
	test_expansion(128'hcca7c55bf3ed623f46f83919f656d78c, {16'd16810, 16'd28939, 16'd6160, 16'd39749, 16'd28201, 16'd30104, 16'd28648, 16'd14458, 16'd12374, 16'd30006, 16'd54719, 16'd18189, 16'd64447, 16'd16933, 16'd21995, 16'd24253, 16'd11852, 16'd21913, 16'd54461, 16'd13252, 16'd37996, 16'd44201, 16'd25584, 16'd36886, 16'd43722, 16'd17246});
	test_expansion(128'h0322f2bdb722195343c6f61964339ef9, {16'd21619, 16'd47058, 16'd24409, 16'd12671, 16'd62724, 16'd38258, 16'd14663, 16'd2562, 16'd5540, 16'd58637, 16'd57314, 16'd51873, 16'd42123, 16'd57828, 16'd49204, 16'd18503, 16'd12378, 16'd54294, 16'd32164, 16'd58497, 16'd42283, 16'd3131, 16'd2357, 16'd24402, 16'd54035, 16'd32754});
	test_expansion(128'h418ad6cf822e08dd9eca886a4dc1e77e, {16'd58239, 16'd17308, 16'd63571, 16'd16041, 16'd64859, 16'd44788, 16'd34931, 16'd41891, 16'd28837, 16'd39692, 16'd17381, 16'd42274, 16'd51137, 16'd29356, 16'd48431, 16'd60807, 16'd13348, 16'd3849, 16'd52090, 16'd20084, 16'd52255, 16'd47910, 16'd57354, 16'd8406, 16'd18346, 16'd6265});
	test_expansion(128'h6825a806aa1a7622fbd25dad37a0d7f8, {16'd32892, 16'd58019, 16'd52126, 16'd49895, 16'd1907, 16'd56626, 16'd9499, 16'd2644, 16'd58469, 16'd36988, 16'd45828, 16'd31952, 16'd37715, 16'd41501, 16'd45254, 16'd32979, 16'd55118, 16'd64086, 16'd24528, 16'd47022, 16'd20187, 16'd24239, 16'd60270, 16'd60847, 16'd509, 16'd24562});
	test_expansion(128'h2f4024facd97978aa75d93f3da50018f, {16'd65339, 16'd6718, 16'd43902, 16'd63116, 16'd12758, 16'd18597, 16'd36027, 16'd48561, 16'd57642, 16'd57806, 16'd48801, 16'd2162, 16'd19299, 16'd4167, 16'd57016, 16'd11702, 16'd4692, 16'd40336, 16'd33688, 16'd16758, 16'd4245, 16'd6893, 16'd20972, 16'd17926, 16'd52882, 16'd46738});
	test_expansion(128'h8bfbbc16af771896006f1a77ea230e6c, {16'd32491, 16'd17245, 16'd28866, 16'd61918, 16'd52191, 16'd33563, 16'd20203, 16'd44060, 16'd3337, 16'd25199, 16'd43636, 16'd24867, 16'd64420, 16'd41873, 16'd1371, 16'd13327, 16'd59117, 16'd59442, 16'd23394, 16'd48409, 16'd11358, 16'd50658, 16'd53144, 16'd21509, 16'd1747, 16'd52359});
	test_expansion(128'h5ad14d432fa38e663a08bfe479500a6a, {16'd47445, 16'd38500, 16'd13051, 16'd36685, 16'd19981, 16'd21020, 16'd15897, 16'd54670, 16'd18074, 16'd7579, 16'd13678, 16'd60646, 16'd29061, 16'd42312, 16'd15020, 16'd13951, 16'd22041, 16'd22685, 16'd31379, 16'd56437, 16'd62802, 16'd24056, 16'd16203, 16'd60346, 16'd16197, 16'd18499});
	test_expansion(128'h73fa2af6774569a116b74f51293694fb, {16'd34336, 16'd32039, 16'd24005, 16'd61682, 16'd41536, 16'd1021, 16'd57047, 16'd53092, 16'd36891, 16'd65248, 16'd25710, 16'd33595, 16'd4719, 16'd47723, 16'd35926, 16'd33344, 16'd52246, 16'd7911, 16'd6235, 16'd34209, 16'd12172, 16'd14683, 16'd31615, 16'd17886, 16'd10879, 16'd32847});
	test_expansion(128'hab8764119ab024599adfc2c9b8bb45e9, {16'd21734, 16'd1957, 16'd5764, 16'd51868, 16'd43195, 16'd12367, 16'd55685, 16'd62079, 16'd3431, 16'd40574, 16'd57362, 16'd1926, 16'd31011, 16'd8967, 16'd56229, 16'd26153, 16'd53608, 16'd31358, 16'd30018, 16'd57715, 16'd26388, 16'd44031, 16'd51674, 16'd51307, 16'd30003, 16'd17385});
	test_expansion(128'ha939c4c2b75a4cef87b3f53a7c496fa2, {16'd8641, 16'd25658, 16'd36072, 16'd36720, 16'd33752, 16'd49265, 16'd38094, 16'd46531, 16'd9121, 16'd24869, 16'd35074, 16'd44773, 16'd10460, 16'd58746, 16'd23024, 16'd30764, 16'd26695, 16'd51654, 16'd33458, 16'd1670, 16'd59278, 16'd5272, 16'd48160, 16'd31247, 16'd32908, 16'd10117});
	test_expansion(128'h3ae9d879f5d93efc8d9d173769a43ebe, {16'd4963, 16'd3951, 16'd15108, 16'd8856, 16'd64731, 16'd18357, 16'd17380, 16'd44204, 16'd34436, 16'd28801, 16'd55954, 16'd63426, 16'd19891, 16'd56342, 16'd54313, 16'd16916, 16'd27212, 16'd24815, 16'd7036, 16'd33126, 16'd7526, 16'd54408, 16'd7429, 16'd55156, 16'd52777, 16'd46663});
	test_expansion(128'h27925758e054dcd621bb80a9638c7c99, {16'd36250, 16'd58613, 16'd59229, 16'd56145, 16'd53317, 16'd39112, 16'd6053, 16'd11806, 16'd22698, 16'd44450, 16'd17792, 16'd57950, 16'd52006, 16'd48972, 16'd8224, 16'd20282, 16'd33998, 16'd48747, 16'd20857, 16'd28349, 16'd59081, 16'd51367, 16'd30847, 16'd8803, 16'd42003, 16'd18473});
	test_expansion(128'h1b5a2b0b187b3b430b353b55b49e60ae, {16'd19355, 16'd17166, 16'd38955, 16'd43962, 16'd42390, 16'd51345, 16'd10102, 16'd12891, 16'd58975, 16'd12412, 16'd38471, 16'd11441, 16'd46521, 16'd43638, 16'd1621, 16'd14776, 16'd11980, 16'd42035, 16'd26016, 16'd23053, 16'd23762, 16'd42979, 16'd2323, 16'd34655, 16'd13636, 16'd50600});
	test_expansion(128'hc44122ece8fe8d965f5edb9f93155fac, {16'd20108, 16'd21256, 16'd13726, 16'd38519, 16'd32327, 16'd49967, 16'd57282, 16'd29541, 16'd46624, 16'd39885, 16'd50003, 16'd53916, 16'd38464, 16'd34043, 16'd32489, 16'd55432, 16'd51240, 16'd36537, 16'd41402, 16'd55814, 16'd54879, 16'd16088, 16'd22050, 16'd11715, 16'd52884, 16'd64325});
	test_expansion(128'hd41b0e4fc1e5dc76be814c5d59172d42, {16'd4643, 16'd11537, 16'd20239, 16'd61600, 16'd39226, 16'd36783, 16'd45679, 16'd51829, 16'd24407, 16'd11969, 16'd29355, 16'd38713, 16'd4280, 16'd33507, 16'd33143, 16'd21717, 16'd5827, 16'd15282, 16'd60236, 16'd35799, 16'd63248, 16'd42711, 16'd30822, 16'd33545, 16'd23217, 16'd29559});
	test_expansion(128'h344fc9d30762f21488640c1ecccea681, {16'd32414, 16'd42479, 16'd27899, 16'd62830, 16'd43982, 16'd33176, 16'd46934, 16'd64914, 16'd46511, 16'd19125, 16'd34274, 16'd2398, 16'd3788, 16'd48170, 16'd49692, 16'd49470, 16'd48898, 16'd813, 16'd54747, 16'd53865, 16'd29280, 16'd64310, 16'd62937, 16'd35354, 16'd2092, 16'd3793});
	test_expansion(128'hdc77cfaedc214d0ad89b1270c27425fa, {16'd425, 16'd8417, 16'd55922, 16'd10320, 16'd61563, 16'd35321, 16'd60116, 16'd43356, 16'd20415, 16'd8009, 16'd52958, 16'd30470, 16'd24707, 16'd43498, 16'd65465, 16'd7316, 16'd14600, 16'd62766, 16'd10133, 16'd53971, 16'd8820, 16'd18056, 16'd17667, 16'd8391, 16'd11215, 16'd48236});
	test_expansion(128'h66e458fd320a231fed0be0665452c3a1, {16'd35793, 16'd45813, 16'd2434, 16'd45764, 16'd46810, 16'd60387, 16'd2508, 16'd4241, 16'd23321, 16'd35370, 16'd35366, 16'd38146, 16'd16957, 16'd11918, 16'd60017, 16'd26618, 16'd52897, 16'd8735, 16'd55928, 16'd11265, 16'd46181, 16'd35300, 16'd20102, 16'd41336, 16'd65480, 16'd9080});
	test_expansion(128'h8b84294318ee6e4823606fefbd421a8a, {16'd53492, 16'd38773, 16'd36675, 16'd58413, 16'd45840, 16'd63520, 16'd37741, 16'd23742, 16'd45818, 16'd15755, 16'd14512, 16'd62850, 16'd6937, 16'd16111, 16'd44078, 16'd54497, 16'd25044, 16'd17358, 16'd42748, 16'd8525, 16'd9464, 16'd23895, 16'd17427, 16'd54059, 16'd13234, 16'd16339});
	test_expansion(128'h17cd4d87561693f40670f37328728aea, {16'd4385, 16'd34285, 16'd23188, 16'd48582, 16'd46961, 16'd19435, 16'd40888, 16'd37466, 16'd43248, 16'd62505, 16'd36677, 16'd6320, 16'd24642, 16'd44000, 16'd8672, 16'd4845, 16'd56642, 16'd45490, 16'd10947, 16'd63105, 16'd45824, 16'd61671, 16'd15158, 16'd16133, 16'd33936, 16'd40916});
	test_expansion(128'hfb9d3baa73a926caaa26cfe4502c9fef, {16'd23923, 16'd65080, 16'd55582, 16'd65094, 16'd34, 16'd25016, 16'd11077, 16'd26138, 16'd52465, 16'd28109, 16'd32520, 16'd64454, 16'd14093, 16'd21935, 16'd18534, 16'd8335, 16'd13489, 16'd22898, 16'd41700, 16'd38728, 16'd4947, 16'd45917, 16'd52221, 16'd30407, 16'd57974, 16'd23199});
	test_expansion(128'h6659f8d6704439fd25bb02cd8a5c2cc3, {16'd52425, 16'd62291, 16'd25854, 16'd116, 16'd40790, 16'd36749, 16'd29375, 16'd26327, 16'd8399, 16'd35144, 16'd44353, 16'd15706, 16'd19814, 16'd2011, 16'd41745, 16'd55783, 16'd22133, 16'd29402, 16'd49700, 16'd51360, 16'd46184, 16'd16689, 16'd48997, 16'd1984, 16'd22149, 16'd56789});
	test_expansion(128'hc6d2824b390489c9b7495af2aeae1b1e, {16'd50312, 16'd16591, 16'd48500, 16'd4173, 16'd13381, 16'd15202, 16'd56240, 16'd21055, 16'd41632, 16'd58984, 16'd54817, 16'd53877, 16'd41549, 16'd27596, 16'd30078, 16'd56914, 16'd13208, 16'd30230, 16'd9181, 16'd9092, 16'd29745, 16'd54564, 16'd45260, 16'd29114, 16'd46331, 16'd19135});
	test_expansion(128'h026f9bda389e24278f43dd873f1095ac, {16'd19190, 16'd43673, 16'd18078, 16'd2443, 16'd29925, 16'd37781, 16'd33073, 16'd64770, 16'd53329, 16'd38002, 16'd40272, 16'd19392, 16'd37901, 16'd58595, 16'd14230, 16'd9157, 16'd9639, 16'd49440, 16'd37175, 16'd38909, 16'd65180, 16'd52553, 16'd53054, 16'd19713, 16'd6834, 16'd32136});
	test_expansion(128'haaf2dc9bf72cd3d13dd5f61033c85bee, {16'd20317, 16'd18727, 16'd25878, 16'd5680, 16'd9441, 16'd59564, 16'd19235, 16'd46513, 16'd58688, 16'd14649, 16'd31587, 16'd60816, 16'd34936, 16'd49270, 16'd15032, 16'd28850, 16'd49697, 16'd45995, 16'd20781, 16'd19266, 16'd21569, 16'd46694, 16'd17417, 16'd43037, 16'd46169, 16'd17238});
	test_expansion(128'h1beff77d127d236c40f971a4603d522e, {16'd12699, 16'd36809, 16'd20133, 16'd56527, 16'd3825, 16'd24122, 16'd3120, 16'd3273, 16'd39214, 16'd48513, 16'd18427, 16'd39538, 16'd25876, 16'd29267, 16'd33526, 16'd39031, 16'd61985, 16'd24144, 16'd12512, 16'd51126, 16'd7925, 16'd60088, 16'd49433, 16'd23903, 16'd11657, 16'd41296});
	test_expansion(128'hb7c251eb1cb0ee4d27af52ace1768ee8, {16'd58824, 16'd4230, 16'd41077, 16'd36970, 16'd17612, 16'd2104, 16'd17487, 16'd828, 16'd3150, 16'd41850, 16'd16973, 16'd44612, 16'd33694, 16'd13463, 16'd31583, 16'd63693, 16'd64394, 16'd28321, 16'd39886, 16'd18068, 16'd38355, 16'd14639, 16'd3371, 16'd5368, 16'd50936, 16'd2378});
	test_expansion(128'h8ec7cc16f351a081672ac19f8416bffb, {16'd16792, 16'd12042, 16'd10085, 16'd8320, 16'd377, 16'd57465, 16'd37459, 16'd52298, 16'd49784, 16'd53434, 16'd35321, 16'd29107, 16'd796, 16'd39399, 16'd34263, 16'd17979, 16'd25476, 16'd27206, 16'd4040, 16'd61069, 16'd38495, 16'd28199, 16'd57157, 16'd25585, 16'd41920, 16'd55581});
	test_expansion(128'h5ef026c7e7ed5b1fe27c6aaf947fe991, {16'd33902, 16'd8375, 16'd28776, 16'd57557, 16'd25580, 16'd26822, 16'd22086, 16'd5905, 16'd21541, 16'd51047, 16'd11330, 16'd38064, 16'd12816, 16'd63375, 16'd52241, 16'd25323, 16'd35501, 16'd61888, 16'd25420, 16'd56686, 16'd41385, 16'd8055, 16'd20309, 16'd19202, 16'd9299, 16'd52351});
	test_expansion(128'hda69370cea0c1ee88ddc7447cd3b28e8, {16'd25999, 16'd35145, 16'd56650, 16'd26997, 16'd23361, 16'd1634, 16'd18352, 16'd4405, 16'd45298, 16'd27169, 16'd40192, 16'd54376, 16'd60782, 16'd32941, 16'd12131, 16'd22305, 16'd51422, 16'd56738, 16'd31025, 16'd6213, 16'd41774, 16'd22452, 16'd60465, 16'd60072, 16'd32721, 16'd33100});
	test_expansion(128'h80736bcfaa14e5db7a94b9b17e04cd30, {16'd60616, 16'd11144, 16'd11251, 16'd43108, 16'd38569, 16'd57810, 16'd19129, 16'd21675, 16'd48753, 16'd14229, 16'd54435, 16'd58953, 16'd2398, 16'd30852, 16'd13629, 16'd4148, 16'd33860, 16'd29934, 16'd10790, 16'd15779, 16'd48580, 16'd62855, 16'd14123, 16'd4540, 16'd24851, 16'd32506});
	test_expansion(128'h88e55e04c3c3e7c30b92ef1e7a60b4c2, {16'd1709, 16'd18617, 16'd46935, 16'd57257, 16'd29269, 16'd25934, 16'd18710, 16'd17949, 16'd10928, 16'd34372, 16'd8645, 16'd54625, 16'd17807, 16'd9730, 16'd42158, 16'd56353, 16'd42635, 16'd32274, 16'd21179, 16'd14115, 16'd14190, 16'd12775, 16'd21473, 16'd56366, 16'd57721, 16'd57209});
	test_expansion(128'h6904b397cbcf6fd470df07f3a0320ca3, {16'd40633, 16'd2393, 16'd44103, 16'd23502, 16'd13426, 16'd19459, 16'd9639, 16'd51599, 16'd6614, 16'd26512, 16'd37214, 16'd59534, 16'd22107, 16'd13916, 16'd19404, 16'd33330, 16'd3346, 16'd42983, 16'd43972, 16'd8340, 16'd49092, 16'd15305, 16'd8559, 16'd62297, 16'd24058, 16'd25559});
	test_expansion(128'h6f048613745af23aa79cc103f573a730, {16'd35461, 16'd8270, 16'd45666, 16'd49986, 16'd33441, 16'd18782, 16'd43173, 16'd37813, 16'd63182, 16'd46412, 16'd21276, 16'd36413, 16'd2409, 16'd5304, 16'd30033, 16'd9887, 16'd30291, 16'd22585, 16'd43672, 16'd28807, 16'd40478, 16'd56101, 16'd9148, 16'd45718, 16'd53670, 16'd41573});
	test_expansion(128'h6d491b672a7a282ec78de7e2f81e518c, {16'd52152, 16'd8516, 16'd400, 16'd47236, 16'd6975, 16'd54803, 16'd9838, 16'd31288, 16'd9672, 16'd42505, 16'd9470, 16'd6732, 16'd63020, 16'd45127, 16'd23431, 16'd48696, 16'd24005, 16'd41619, 16'd3220, 16'd22673, 16'd36608, 16'd51588, 16'd614, 16'd184, 16'd16440, 16'd19032});
	test_expansion(128'h45f361da081c59471e5588ef96f65d6d, {16'd55562, 16'd17578, 16'd58184, 16'd52219, 16'd34632, 16'd27396, 16'd39789, 16'd42151, 16'd23724, 16'd3192, 16'd2798, 16'd29593, 16'd16083, 16'd61810, 16'd27863, 16'd1378, 16'd33719, 16'd10222, 16'd8916, 16'd20416, 16'd47294, 16'd29590, 16'd48526, 16'd45184, 16'd36522, 16'd58893});
	test_expansion(128'h7e1c08f2311c1c1c7fbe71c78c973201, {16'd29588, 16'd58087, 16'd34801, 16'd16865, 16'd14662, 16'd53585, 16'd39247, 16'd9615, 16'd38690, 16'd19373, 16'd63921, 16'd21539, 16'd21912, 16'd27249, 16'd53809, 16'd11280, 16'd48855, 16'd60106, 16'd8853, 16'd44428, 16'd8059, 16'd38797, 16'd4157, 16'd61466, 16'd36517, 16'd57873});
	test_expansion(128'ha33502f3ba6895608d65a5b70d7f025a, {16'd35440, 16'd21867, 16'd31869, 16'd47692, 16'd36656, 16'd18752, 16'd21997, 16'd42448, 16'd58224, 16'd10594, 16'd33289, 16'd19594, 16'd44366, 16'd17434, 16'd65083, 16'd56944, 16'd5646, 16'd27733, 16'd19089, 16'd64424, 16'd12528, 16'd62401, 16'd9440, 16'd10150, 16'd18724, 16'd18036});
	test_expansion(128'h05e475439af3277e82ca36822f46e0fc, {16'd55065, 16'd4194, 16'd47562, 16'd35483, 16'd54198, 16'd25675, 16'd54212, 16'd64906, 16'd17274, 16'd55232, 16'd36673, 16'd5743, 16'd41654, 16'd34681, 16'd52061, 16'd26085, 16'd28353, 16'd42300, 16'd43065, 16'd25334, 16'd24424, 16'd18446, 16'd17961, 16'd26529, 16'd55333, 16'd60484});
	test_expansion(128'h69a6daf77e3b4763e77386e3a7a9ca0b, {16'd32743, 16'd54689, 16'd33078, 16'd22950, 16'd29208, 16'd17903, 16'd51891, 16'd43224, 16'd2919, 16'd54771, 16'd37938, 16'd5262, 16'd1267, 16'd9192, 16'd31119, 16'd60154, 16'd63170, 16'd12701, 16'd34988, 16'd7895, 16'd10876, 16'd51841, 16'd45915, 16'd3437, 16'd38062, 16'd8752});
	test_expansion(128'h71f4e3ddd456d46a5e32efff4e61f15d, {16'd62380, 16'd35469, 16'd64868, 16'd33590, 16'd37999, 16'd60136, 16'd49705, 16'd9463, 16'd36530, 16'd27229, 16'd34363, 16'd25748, 16'd18239, 16'd26729, 16'd18083, 16'd12682, 16'd21925, 16'd58030, 16'd27156, 16'd16480, 16'd53974, 16'd54345, 16'd7620, 16'd56472, 16'd51045, 16'd32453});
	test_expansion(128'h14b9db47bc0459d3b95a73a50be166b4, {16'd4865, 16'd46155, 16'd15936, 16'd29864, 16'd22128, 16'd18815, 16'd65303, 16'd20949, 16'd9375, 16'd6010, 16'd57226, 16'd30712, 16'd53036, 16'd21378, 16'd48633, 16'd4993, 16'd55512, 16'd49572, 16'd38221, 16'd42576, 16'd13376, 16'd43202, 16'd62420, 16'd19775, 16'd24754, 16'd45113});
	test_expansion(128'h8fcf70f1335054977c290e54a030bdae, {16'd64553, 16'd55113, 16'd5458, 16'd4367, 16'd1506, 16'd28385, 16'd1612, 16'd51417, 16'd9209, 16'd26328, 16'd29240, 16'd42874, 16'd16769, 16'd3134, 16'd62345, 16'd17086, 16'd17899, 16'd36785, 16'd49308, 16'd14228, 16'd58022, 16'd27096, 16'd34469, 16'd23194, 16'd35910, 16'd39733});
	test_expansion(128'hb6b6095813274fabad39c6f060f58ae8, {16'd14209, 16'd37166, 16'd35847, 16'd48375, 16'd30055, 16'd39503, 16'd63122, 16'd28172, 16'd26092, 16'd61694, 16'd22498, 16'd33370, 16'd6955, 16'd29412, 16'd58838, 16'd17333, 16'd34464, 16'd35542, 16'd25298, 16'd48081, 16'd45130, 16'd25844, 16'd3906, 16'd9789, 16'd51057, 16'd8339});
	test_expansion(128'h9efc39e4d921c34c6cf8c7517349f15c, {16'd62659, 16'd25171, 16'd31304, 16'd11588, 16'd20296, 16'd39213, 16'd23872, 16'd27758, 16'd6560, 16'd55810, 16'd49614, 16'd53063, 16'd54672, 16'd42650, 16'd25631, 16'd58994, 16'd2367, 16'd61103, 16'd33921, 16'd50517, 16'd42818, 16'd43423, 16'd16358, 16'd61682, 16'd29493, 16'd46333});
	test_expansion(128'h22b2722b470b2f2b0523262b192ef12a, {16'd35056, 16'd58092, 16'd15491, 16'd9584, 16'd57391, 16'd5637, 16'd58, 16'd11367, 16'd2084, 16'd4118, 16'd64434, 16'd58876, 16'd22053, 16'd61796, 16'd24563, 16'd42429, 16'd764, 16'd48938, 16'd25587, 16'd29661, 16'd41990, 16'd47516, 16'd11503, 16'd2470, 16'd10159, 16'd60721});
	test_expansion(128'hc0a1c565cd1f4a578f223932a881bc14, {16'd36087, 16'd14564, 16'd32978, 16'd52668, 16'd13041, 16'd3064, 16'd34849, 16'd6478, 16'd29184, 16'd13093, 16'd44820, 16'd40390, 16'd43982, 16'd4526, 16'd24202, 16'd25623, 16'd4048, 16'd19956, 16'd64603, 16'd123, 16'd47087, 16'd27235, 16'd63240, 16'd45795, 16'd59183, 16'd14371});
	test_expansion(128'h79562435c50986bd8f5864f49d716f0a, {16'd1113, 16'd57947, 16'd34952, 16'd37517, 16'd2941, 16'd30178, 16'd21279, 16'd59361, 16'd28183, 16'd31491, 16'd48778, 16'd63566, 16'd15197, 16'd35562, 16'd47637, 16'd24800, 16'd42047, 16'd9393, 16'd59466, 16'd2373, 16'd35335, 16'd20490, 16'd37381, 16'd26127, 16'd797, 16'd51943});
	test_expansion(128'hac9eee0d4fe4e94d96f7c6a3980fb0e6, {16'd2219, 16'd13424, 16'd58020, 16'd58171, 16'd343, 16'd10829, 16'd26839, 16'd5803, 16'd21298, 16'd48457, 16'd53343, 16'd9493, 16'd42361, 16'd45205, 16'd40710, 16'd60901, 16'd62601, 16'd58072, 16'd40440, 16'd2099, 16'd567, 16'd14077, 16'd37432, 16'd13866, 16'd5309, 16'd23127});
	test_expansion(128'hf2fc8746a310273d97db85b3f2fa0a4c, {16'd252, 16'd57861, 16'd47796, 16'd15741, 16'd55045, 16'd28705, 16'd31591, 16'd58521, 16'd45899, 16'd26775, 16'd523, 16'd19123, 16'd36842, 16'd53911, 16'd27132, 16'd35177, 16'd35978, 16'd9349, 16'd44856, 16'd51287, 16'd3738, 16'd45636, 16'd23585, 16'd11793, 16'd29193, 16'd28138});
	test_expansion(128'h97ed8743cdf907ea5a9eac7e80361d79, {16'd19056, 16'd38894, 16'd44824, 16'd62680, 16'd10628, 16'd2520, 16'd9732, 16'd48398, 16'd46386, 16'd44065, 16'd23003, 16'd20367, 16'd16391, 16'd6413, 16'd22224, 16'd13166, 16'd11244, 16'd31861, 16'd28055, 16'd14356, 16'd18781, 16'd41425, 16'd15921, 16'd53033, 16'd26809, 16'd59303});
	test_expansion(128'hbcb852dd03797a9794e39c7d6b02cde7, {16'd42587, 16'd44368, 16'd58636, 16'd36823, 16'd9579, 16'd51715, 16'd38771, 16'd721, 16'd40440, 16'd20328, 16'd20619, 16'd49540, 16'd32003, 16'd9396, 16'd6931, 16'd57275, 16'd22038, 16'd19257, 16'd44955, 16'd40906, 16'd5481, 16'd21961, 16'd63586, 16'd35834, 16'd57394, 16'd11110});
	test_expansion(128'h84e27d707405bcdd0659b36da6dd7d7d, {16'd50626, 16'd36091, 16'd36020, 16'd1631, 16'd3949, 16'd54818, 16'd36889, 16'd7526, 16'd21379, 16'd15883, 16'd32998, 16'd21912, 16'd29659, 16'd19674, 16'd3796, 16'd64080, 16'd25262, 16'd40063, 16'd46168, 16'd28569, 16'd19880, 16'd43856, 16'd32358, 16'd15913, 16'd5557, 16'd38713});
	test_expansion(128'hac425a5564abc554b72082b5d0594e36, {16'd58105, 16'd57046, 16'd10398, 16'd56614, 16'd15972, 16'd14099, 16'd53290, 16'd9424, 16'd695, 16'd40497, 16'd52628, 16'd16967, 16'd29000, 16'd60605, 16'd30933, 16'd59695, 16'd61259, 16'd43929, 16'd4640, 16'd22266, 16'd27550, 16'd58412, 16'd7837, 16'd54771, 16'd43954, 16'd7332});
	test_expansion(128'hdabeba95553022d68e535aff79cdf7da, {16'd28360, 16'd51216, 16'd20219, 16'd47335, 16'd8191, 16'd37069, 16'd47767, 16'd60280, 16'd61232, 16'd7632, 16'd19316, 16'd57505, 16'd61066, 16'd22255, 16'd38686, 16'd11378, 16'd17583, 16'd19430, 16'd31437, 16'd25860, 16'd43192, 16'd12119, 16'd56756, 16'd963, 16'd50716, 16'd8521});
	test_expansion(128'h3640cac219f7835759f497a333e99c10, {16'd29855, 16'd28788, 16'd2726, 16'd55967, 16'd49979, 16'd9764, 16'd57101, 16'd50947, 16'd64255, 16'd36007, 16'd38205, 16'd6233, 16'd60969, 16'd53347, 16'd57977, 16'd13332, 16'd8418, 16'd42348, 16'd6635, 16'd8389, 16'd64447, 16'd10973, 16'd1877, 16'd1209, 16'd37976, 16'd13183});
	test_expansion(128'hc70c5fdee21ef62abf29157550a63792, {16'd5468, 16'd2846, 16'd34718, 16'd50694, 16'd41349, 16'd51034, 16'd9720, 16'd41459, 16'd49542, 16'd64369, 16'd48308, 16'd56025, 16'd40455, 16'd60610, 16'd17098, 16'd5136, 16'd41113, 16'd46880, 16'd22164, 16'd19877, 16'd48642, 16'd34384, 16'd18155, 16'd37786, 16'd57819, 16'd27870});
	test_expansion(128'h64ba6735ec6dc523f3632d8197f6e5e8, {16'd1787, 16'd50929, 16'd58381, 16'd38563, 16'd16213, 16'd8787, 16'd45322, 16'd2534, 16'd10818, 16'd64106, 16'd23572, 16'd21251, 16'd19649, 16'd23368, 16'd6592, 16'd38000, 16'd53107, 16'd37203, 16'd64177, 16'd61305, 16'd33063, 16'd10462, 16'd14245, 16'd34186, 16'd30549, 16'd13786});
	test_expansion(128'h7bd15b5b94652fcb63b520ab722431fa, {16'd19908, 16'd29359, 16'd1372, 16'd5496, 16'd2195, 16'd588, 16'd44922, 16'd65220, 16'd57737, 16'd15498, 16'd2418, 16'd58176, 16'd29049, 16'd28953, 16'd18241, 16'd47343, 16'd43714, 16'd35589, 16'd28717, 16'd56454, 16'd13381, 16'd31171, 16'd50419, 16'd11724, 16'd53693, 16'd63072});
	test_expansion(128'h6df70bc60a2d22c30163edef0937fe6d, {16'd37801, 16'd42691, 16'd13686, 16'd47641, 16'd15159, 16'd32763, 16'd44585, 16'd21580, 16'd57355, 16'd38221, 16'd55350, 16'd50720, 16'd3464, 16'd56340, 16'd48520, 16'd64282, 16'd26309, 16'd56699, 16'd12178, 16'd34388, 16'd37133, 16'd33615, 16'd19562, 16'd61857, 16'd33465, 16'd53021});
	test_expansion(128'h192cb218b68e58910ccdf5f39f6e9272, {16'd42054, 16'd25236, 16'd53873, 16'd54173, 16'd47682, 16'd26557, 16'd28244, 16'd41676, 16'd37599, 16'd14857, 16'd44960, 16'd8913, 16'd10516, 16'd57016, 16'd32337, 16'd7676, 16'd63290, 16'd60076, 16'd19492, 16'd55623, 16'd8381, 16'd25061, 16'd43133, 16'd23716, 16'd26393, 16'd45998});
	test_expansion(128'h0dad5e0ec2d449d0dab1cedb5ee703d4, {16'd62286, 16'd57364, 16'd44571, 16'd24919, 16'd2188, 16'd6279, 16'd12032, 16'd39892, 16'd52026, 16'd6049, 16'd57531, 16'd14387, 16'd14651, 16'd65006, 16'd4381, 16'd51494, 16'd51704, 16'd43410, 16'd27739, 16'd60381, 16'd58246, 16'd58898, 16'd47721, 16'd41960, 16'd22134, 16'd46104});
	test_expansion(128'h5974902121809d70afff772a3949bc3d, {16'd43282, 16'd53824, 16'd39760, 16'd21031, 16'd13466, 16'd5093, 16'd14058, 16'd43526, 16'd59975, 16'd3220, 16'd22161, 16'd24377, 16'd63632, 16'd5378, 16'd20854, 16'd13801, 16'd49676, 16'd26513, 16'd324, 16'd3329, 16'd27019, 16'd392, 16'd26746, 16'd54612, 16'd40729, 16'd17935});
	test_expansion(128'ha44cd3e72f949afa636f300f446e97b9, {16'd2533, 16'd2816, 16'd37304, 16'd40888, 16'd36881, 16'd57749, 16'd24294, 16'd64520, 16'd20028, 16'd35467, 16'd18541, 16'd43006, 16'd26349, 16'd61853, 16'd45309, 16'd58795, 16'd58108, 16'd26270, 16'd9099, 16'd5818, 16'd9593, 16'd4086, 16'd44752, 16'd64853, 16'd56776, 16'd54738});
	test_expansion(128'he2b4ab65ac8b4f49dd6c8bea7b2bdab2, {16'd29618, 16'd32785, 16'd32720, 16'd10448, 16'd63131, 16'd14612, 16'd35931, 16'd35067, 16'd36076, 16'd1859, 16'd16489, 16'd35499, 16'd25370, 16'd49079, 16'd32399, 16'd29998, 16'd6259, 16'd11477, 16'd42525, 16'd47738, 16'd60858, 16'd38951, 16'd50746, 16'd35529, 16'd56217, 16'd9071});
	test_expansion(128'h0e124433ff092a54796dc55c91a055d3, {16'd56597, 16'd45507, 16'd19752, 16'd39541, 16'd5568, 16'd63140, 16'd36235, 16'd38387, 16'd55295, 16'd27745, 16'd8620, 16'd36774, 16'd42296, 16'd41077, 16'd64185, 16'd39119, 16'd15195, 16'd7717, 16'd47156, 16'd20974, 16'd17573, 16'd18694, 16'd31901, 16'd9113, 16'd4607, 16'd3238});
	test_expansion(128'h1167889a10fcfd34af39c6b2880d432c, {16'd10020, 16'd32970, 16'd18440, 16'd7039, 16'd12847, 16'd29642, 16'd6675, 16'd34275, 16'd4667, 16'd34423, 16'd43939, 16'd24519, 16'd18610, 16'd35214, 16'd4240, 16'd2045, 16'd16942, 16'd65283, 16'd40662, 16'd64373, 16'd23322, 16'd18070, 16'd14318, 16'd37586, 16'd23300, 16'd50376});
	test_expansion(128'h944bbabf2cd969a29ed611e086f62e40, {16'd3167, 16'd61800, 16'd46832, 16'd51754, 16'd24200, 16'd44237, 16'd11745, 16'd40374, 16'd34631, 16'd42411, 16'd2173, 16'd43950, 16'd26019, 16'd41940, 16'd21798, 16'd38507, 16'd46658, 16'd23537, 16'd1955, 16'd33514, 16'd54073, 16'd7088, 16'd49464, 16'd62392, 16'd48410, 16'd10537});
	test_expansion(128'hb40d688930dd4128a1f7c544dac02bef, {16'd15529, 16'd36582, 16'd54542, 16'd65207, 16'd11883, 16'd33425, 16'd32082, 16'd7816, 16'd18266, 16'd8791, 16'd24270, 16'd40545, 16'd4999, 16'd5221, 16'd63053, 16'd35064, 16'd4795, 16'd45363, 16'd61155, 16'd49184, 16'd60129, 16'd32354, 16'd45702, 16'd56441, 16'd41827, 16'd62121});
	test_expansion(128'h13199dc182503bdebb140c5256f5e4dd, {16'd11021, 16'd6215, 16'd25452, 16'd28158, 16'd38583, 16'd39448, 16'd51111, 16'd46699, 16'd44505, 16'd19004, 16'd43980, 16'd7895, 16'd41000, 16'd57310, 16'd59367, 16'd40148, 16'd65040, 16'd65286, 16'd64757, 16'd27838, 16'd42993, 16'd46367, 16'd23362, 16'd12034, 16'd65524, 16'd8309});
	test_expansion(128'hf09a0ae19ca3f2ddd4a9f288804f2014, {16'd44098, 16'd52166, 16'd11166, 16'd17584, 16'd24105, 16'd61490, 16'd16167, 16'd23284, 16'd32775, 16'd64960, 16'd36852, 16'd55385, 16'd33394, 16'd43866, 16'd53000, 16'd28568, 16'd29060, 16'd38030, 16'd63822, 16'd63361, 16'd19853, 16'd30683, 16'd17559, 16'd25066, 16'd37411, 16'd22399});
	test_expansion(128'h463efdc8b4a42c265f94b7b7ba4835ef, {16'd63421, 16'd30268, 16'd36115, 16'd21157, 16'd44611, 16'd16247, 16'd46480, 16'd24541, 16'd63154, 16'd49684, 16'd62050, 16'd42340, 16'd18931, 16'd21928, 16'd13190, 16'd62710, 16'd47318, 16'd46169, 16'd5955, 16'd16057, 16'd43663, 16'd500, 16'd25399, 16'd53082, 16'd58923, 16'd23000});
	test_expansion(128'hbdb76720bda642fb180b1b14547bcb09, {16'd17536, 16'd64463, 16'd17936, 16'd29088, 16'd43558, 16'd6866, 16'd24775, 16'd50442, 16'd17399, 16'd54502, 16'd8120, 16'd41239, 16'd16624, 16'd3002, 16'd12977, 16'd34200, 16'd57582, 16'd46687, 16'd4925, 16'd38433, 16'd708, 16'd64303, 16'd48640, 16'd39854, 16'd47724, 16'd26905});
	test_expansion(128'hc1662d92c6bd06e85511d91ed46d655d, {16'd48827, 16'd32880, 16'd43816, 16'd1479, 16'd27630, 16'd44205, 16'd44282, 16'd34398, 16'd27253, 16'd50579, 16'd60303, 16'd17507, 16'd17008, 16'd35221, 16'd59910, 16'd3988, 16'd65316, 16'd31607, 16'd15542, 16'd10320, 16'd20271, 16'd30213, 16'd61094, 16'd38543, 16'd7705, 16'd26505});
	test_expansion(128'h168d90cf7b36098b8bad65a0aa8c3c2b, {16'd10298, 16'd20057, 16'd57300, 16'd28586, 16'd63499, 16'd54103, 16'd61300, 16'd20460, 16'd46184, 16'd41754, 16'd28289, 16'd114, 16'd8671, 16'd27562, 16'd15504, 16'd19611, 16'd6558, 16'd61631, 16'd32822, 16'd47844, 16'd4067, 16'd31203, 16'd31699, 16'd30507, 16'd50412, 16'd41849});
	test_expansion(128'h0320194f39d9813fa9e7ded01e9c3337, {16'd35500, 16'd18519, 16'd62942, 16'd61441, 16'd50320, 16'd11105, 16'd31854, 16'd24479, 16'd40967, 16'd60318, 16'd13357, 16'd14400, 16'd17788, 16'd30038, 16'd27629, 16'd1585, 16'd30144, 16'd29972, 16'd55662, 16'd42293, 16'd59063, 16'd53579, 16'd24501, 16'd52759, 16'd1327, 16'd12872});
	test_expansion(128'h69ec734ef5072c40321873bc52dd37eb, {16'd5784, 16'd14691, 16'd57082, 16'd62150, 16'd49080, 16'd23587, 16'd37993, 16'd14424, 16'd56973, 16'd5065, 16'd64028, 16'd25246, 16'd46, 16'd61534, 16'd24869, 16'd62546, 16'd40912, 16'd11827, 16'd9255, 16'd59510, 16'd15785, 16'd4213, 16'd59695, 16'd15118, 16'd63178, 16'd60237});
	test_expansion(128'h8255ef5ec99c5227fa44cc69ea4e0f86, {16'd23790, 16'd60048, 16'd40055, 16'd62627, 16'd1545, 16'd23480, 16'd62751, 16'd4406, 16'd59530, 16'd20022, 16'd51268, 16'd31577, 16'd8870, 16'd19386, 16'd51174, 16'd12984, 16'd60028, 16'd1861, 16'd55761, 16'd20086, 16'd1165, 16'd2027, 16'd13173, 16'd44938, 16'd50150, 16'd45280});
	test_expansion(128'hb881cf5ede4a909177a843d429128347, {16'd8278, 16'd6571, 16'd35721, 16'd9116, 16'd789, 16'd52297, 16'd42006, 16'd23745, 16'd8058, 16'd58499, 16'd43149, 16'd18678, 16'd9961, 16'd43088, 16'd49286, 16'd61606, 16'd53601, 16'd45257, 16'd33024, 16'd1721, 16'd59596, 16'd6703, 16'd13905, 16'd47879, 16'd49160, 16'd5393});
	test_expansion(128'h20ed8efa08d157cb9e62eb438c175a85, {16'd42456, 16'd58551, 16'd7839, 16'd1269, 16'd14337, 16'd3611, 16'd4756, 16'd3109, 16'd24543, 16'd3223, 16'd8712, 16'd11971, 16'd28410, 16'd7337, 16'd23053, 16'd32398, 16'd36147, 16'd57365, 16'd22498, 16'd11629, 16'd15488, 16'd12201, 16'd34925, 16'd30922, 16'd719, 16'd22118});
	test_expansion(128'h08f4c867bc30ff8ef944f5edd33c4c17, {16'd44889, 16'd9677, 16'd4015, 16'd16474, 16'd51222, 16'd22951, 16'd33683, 16'd58927, 16'd48196, 16'd54822, 16'd41770, 16'd16501, 16'd7600, 16'd1392, 16'd57495, 16'd63078, 16'd29278, 16'd13656, 16'd51249, 16'd65339, 16'd23881, 16'd53978, 16'd10765, 16'd27632, 16'd47016, 16'd34800});
	test_expansion(128'hd1f71d9ee102ae75118bc05dde4169b0, {16'd37684, 16'd16163, 16'd9294, 16'd5468, 16'd61304, 16'd47986, 16'd55465, 16'd15160, 16'd5484, 16'd6494, 16'd44728, 16'd7196, 16'd42389, 16'd51472, 16'd14348, 16'd45582, 16'd23537, 16'd45584, 16'd23390, 16'd34405, 16'd55424, 16'd52203, 16'd28034, 16'd29444, 16'd28386, 16'd7825});
	test_expansion(128'h710b3d6ddbdc9dc13a6f0294770bfd49, {16'd54133, 16'd10606, 16'd48965, 16'd19177, 16'd3304, 16'd22577, 16'd218, 16'd48347, 16'd49046, 16'd39842, 16'd22690, 16'd26029, 16'd31560, 16'd42655, 16'd7644, 16'd19593, 16'd62850, 16'd43306, 16'd32977, 16'd9680, 16'd15694, 16'd44901, 16'd63155, 16'd45914, 16'd20404, 16'd13843});
	test_expansion(128'h2dfdaa427189fb6addd36817a42b5819, {16'd14352, 16'd53092, 16'd30012, 16'd55465, 16'd37620, 16'd45085, 16'd62836, 16'd51209, 16'd586, 16'd9781, 16'd46577, 16'd2394, 16'd62269, 16'd33402, 16'd41366, 16'd5401, 16'd4746, 16'd58927, 16'd21614, 16'd23474, 16'd31495, 16'd28681, 16'd55202, 16'd18187, 16'd20188, 16'd29212});
	test_expansion(128'hf067ed3406339f9c20e436337542a411, {16'd5822, 16'd21239, 16'd61166, 16'd34253, 16'd61795, 16'd62176, 16'd4598, 16'd36919, 16'd54460, 16'd64366, 16'd13256, 16'd31403, 16'd23094, 16'd47852, 16'd52781, 16'd32088, 16'd32275, 16'd40686, 16'd13458, 16'd24548, 16'd26895, 16'd29632, 16'd42700, 16'd17469, 16'd14710, 16'd47615});
	test_expansion(128'h895ea9d10c354603a372c2330b391073, {16'd56016, 16'd54834, 16'd28843, 16'd30788, 16'd3788, 16'd28210, 16'd29405, 16'd58568, 16'd54956, 16'd44272, 16'd19385, 16'd36161, 16'd29016, 16'd44659, 16'd22554, 16'd17131, 16'd28440, 16'd46110, 16'd24245, 16'd51902, 16'd27061, 16'd38214, 16'd39517, 16'd25876, 16'd5617, 16'd9811});
	test_expansion(128'h4ecc8590cc3d9187513fe94e8c09485b, {16'd2305, 16'd60141, 16'd54049, 16'd23459, 16'd1439, 16'd48548, 16'd35138, 16'd37974, 16'd17244, 16'd46108, 16'd54545, 16'd19884, 16'd7314, 16'd28679, 16'd8502, 16'd6628, 16'd2023, 16'd6878, 16'd24290, 16'd14215, 16'd58588, 16'd55074, 16'd7333, 16'd59991, 16'd34457, 16'd54876});
	test_expansion(128'ha4b1ba5c1fe0a8a9eccc7f3913c494be, {16'd37798, 16'd2095, 16'd13989, 16'd45995, 16'd8875, 16'd40360, 16'd46753, 16'd36522, 16'd64, 16'd28724, 16'd53475, 16'd51036, 16'd10427, 16'd57524, 16'd24798, 16'd46678, 16'd42011, 16'd59372, 16'd13012, 16'd55354, 16'd59020, 16'd5347, 16'd50543, 16'd47399, 16'd39759, 16'd61440});
	test_expansion(128'h532c07d86a532a5a08ea1bc69dec6cdb, {16'd6811, 16'd47356, 16'd238, 16'd44471, 16'd62185, 16'd51056, 16'd16385, 16'd4085, 16'd31292, 16'd21544, 16'd28056, 16'd22294, 16'd45147, 16'd17143, 16'd2637, 16'd31150, 16'd32036, 16'd11573, 16'd25050, 16'd57094, 16'd46244, 16'd38107, 16'd25593, 16'd23192, 16'd34238, 16'd27478});
	test_expansion(128'h9f9d73bca20d202d7125e547e6e21aff, {16'd8342, 16'd23449, 16'd23182, 16'd49298, 16'd25429, 16'd38320, 16'd51532, 16'd7172, 16'd51817, 16'd25866, 16'd1839, 16'd4088, 16'd28432, 16'd32476, 16'd25457, 16'd44801, 16'd414, 16'd42333, 16'd23891, 16'd33532, 16'd19525, 16'd28301, 16'd1334, 16'd52528, 16'd35670, 16'd54145});
	test_expansion(128'h0fe7241999515b508c7ebb76e166cd7d, {16'd54993, 16'd21769, 16'd14632, 16'd21140, 16'd23849, 16'd44883, 16'd32904, 16'd60925, 16'd52671, 16'd19711, 16'd52089, 16'd39548, 16'd21425, 16'd33287, 16'd32789, 16'd6740, 16'd53049, 16'd43758, 16'd24615, 16'd16213, 16'd55558, 16'd43734, 16'd46903, 16'd47921, 16'd40038, 16'd36384});
	test_expansion(128'hce2dd15666416c8677f6064b46e88265, {16'd52110, 16'd10833, 16'd64868, 16'd21629, 16'd63987, 16'd26792, 16'd43045, 16'd32970, 16'd43936, 16'd39187, 16'd52986, 16'd4291, 16'd21969, 16'd61953, 16'd31514, 16'd44002, 16'd10144, 16'd25044, 16'd45295, 16'd8825, 16'd56227, 16'd51275, 16'd26777, 16'd34386, 16'd34899, 16'd63448});
	test_expansion(128'h861191e02d275ddf60fe52bc00f69ba4, {16'd38463, 16'd20518, 16'd44240, 16'd29820, 16'd15070, 16'd61685, 16'd22234, 16'd13227, 16'd55530, 16'd35490, 16'd38429, 16'd29554, 16'd44643, 16'd48661, 16'd3137, 16'd36321, 16'd63969, 16'd62664, 16'd25697, 16'd24785, 16'd27091, 16'd4300, 16'd62696, 16'd15278, 16'd20100, 16'd16504});
	test_expansion(128'hc98c81268a32aa430bb3f3b93abe9ab9, {16'd19614, 16'd27875, 16'd5729, 16'd44183, 16'd30022, 16'd1171, 16'd34945, 16'd28632, 16'd4863, 16'd9326, 16'd45874, 16'd23508, 16'd20890, 16'd14020, 16'd27150, 16'd62694, 16'd4501, 16'd26881, 16'd12093, 16'd61743, 16'd52641, 16'd38886, 16'd2601, 16'd30848, 16'd11514, 16'd13834});
	test_expansion(128'hc543a01dcb271834bc88a84935f7f357, {16'd2653, 16'd5110, 16'd38160, 16'd25777, 16'd9512, 16'd50182, 16'd11604, 16'd11753, 16'd49627, 16'd27959, 16'd53366, 16'd2095, 16'd32839, 16'd46960, 16'd49059, 16'd61351, 16'd36834, 16'd59705, 16'd55067, 16'd53217, 16'd36847, 16'd48019, 16'd64644, 16'd20734, 16'd37717, 16'd31687});
	test_expansion(128'h1a49e923848f610cad9d017867c2c72d, {16'd56939, 16'd24421, 16'd14133, 16'd29995, 16'd49445, 16'd34549, 16'd58608, 16'd10338, 16'd14613, 16'd62744, 16'd2377, 16'd8227, 16'd19465, 16'd44044, 16'd51371, 16'd50161, 16'd38160, 16'd19850, 16'd16516, 16'd56744, 16'd43226, 16'd8399, 16'd12364, 16'd9157, 16'd59678, 16'd3800});
	test_expansion(128'ha2ba979f031bba80991ca9d49d000047, {16'd47325, 16'd15922, 16'd62496, 16'd11645, 16'd39467, 16'd2848, 16'd65064, 16'd27300, 16'd64364, 16'd46307, 16'd20509, 16'd27423, 16'd16464, 16'd7806, 16'd25789, 16'd48012, 16'd45238, 16'd38538, 16'd19949, 16'd22234, 16'd49593, 16'd4503, 16'd53996, 16'd55941, 16'd41755, 16'd4958});
	test_expansion(128'h7d72234ff46d0096031cfca78aa0103e, {16'd8904, 16'd10918, 16'd14485, 16'd43513, 16'd53313, 16'd1771, 16'd57678, 16'd45, 16'd22520, 16'd15043, 16'd38203, 16'd30110, 16'd29348, 16'd38947, 16'd54144, 16'd32237, 16'd4707, 16'd14357, 16'd53159, 16'd14612, 16'd37245, 16'd13392, 16'd49194, 16'd39491, 16'd32815, 16'd18268});
	test_expansion(128'h9bab51a3a6d51212661a1905742f1da8, {16'd42945, 16'd17360, 16'd21983, 16'd40894, 16'd20378, 16'd55120, 16'd62191, 16'd14173, 16'd42280, 16'd21300, 16'd20213, 16'd63099, 16'd45718, 16'd53104, 16'd46551, 16'd65282, 16'd44085, 16'd58570, 16'd32041, 16'd63948, 16'd19921, 16'd36321, 16'd47789, 16'd17079, 16'd10260, 16'd13668});
	test_expansion(128'hcdd282abb36987c36c49160b63ecba44, {16'd44017, 16'd15881, 16'd28913, 16'd40156, 16'd63876, 16'd3587, 16'd40920, 16'd29055, 16'd43403, 16'd55366, 16'd19294, 16'd5531, 16'd1641, 16'd4838, 16'd50661, 16'd39256, 16'd33146, 16'd58023, 16'd51654, 16'd51265, 16'd57086, 16'd63908, 16'd12839, 16'd21583, 16'd19671, 16'd30772});
	test_expansion(128'hc8ce68e4fdd9ae548e023822c22500c4, {16'd43131, 16'd55486, 16'd54694, 16'd36069, 16'd14968, 16'd8984, 16'd7485, 16'd38679, 16'd12072, 16'd23715, 16'd8430, 16'd50842, 16'd39091, 16'd22912, 16'd58651, 16'd49176, 16'd65275, 16'd37668, 16'd19109, 16'd9889, 16'd65280, 16'd28013, 16'd34423, 16'd63966, 16'd14890, 16'd41289});
	test_expansion(128'h957ae28c9613b18dcdbb26adba8858fb, {16'd56595, 16'd41526, 16'd35616, 16'd49675, 16'd50595, 16'd5042, 16'd29355, 16'd26621, 16'd37893, 16'd21634, 16'd31316, 16'd31870, 16'd62603, 16'd4894, 16'd486, 16'd56306, 16'd248, 16'd22346, 16'd39031, 16'd11839, 16'd57514, 16'd62282, 16'd63443, 16'd54942, 16'd47015, 16'd28109});
	test_expansion(128'hd9c38f7f38844284bdeb88bed5aeb8b4, {16'd60320, 16'd19567, 16'd43726, 16'd29015, 16'd26257, 16'd57706, 16'd65246, 16'd36040, 16'd42425, 16'd24377, 16'd64178, 16'd53976, 16'd32217, 16'd35295, 16'd53738, 16'd18003, 16'd31822, 16'd54768, 16'd24451, 16'd64725, 16'd62850, 16'd61358, 16'd23109, 16'd9562, 16'd54351, 16'd4581});
	test_expansion(128'hf317d2f113170162f3354fc7f68c641e, {16'd23121, 16'd63672, 16'd18801, 16'd29471, 16'd44445, 16'd2574, 16'd55162, 16'd27461, 16'd42542, 16'd48441, 16'd35812, 16'd27298, 16'd12853, 16'd59422, 16'd51975, 16'd32625, 16'd13499, 16'd31277, 16'd50837, 16'd45551, 16'd28363, 16'd50816, 16'd210, 16'd9643, 16'd26386, 16'd54848});
	test_expansion(128'h7648ccdb096d290f382c7b2d6fed1be5, {16'd38661, 16'd56987, 16'd3656, 16'd6140, 16'd26903, 16'd52447, 16'd38781, 16'd16949, 16'd23032, 16'd55717, 16'd35825, 16'd41479, 16'd23506, 16'd21672, 16'd39516, 16'd50536, 16'd959, 16'd13663, 16'd15520, 16'd19298, 16'd5795, 16'd12300, 16'd10545, 16'd49692, 16'd4651, 16'd3686});
	test_expansion(128'h0f334a1ef8b82f4917cf32e0bda42f51, {16'd13908, 16'd23468, 16'd53249, 16'd15128, 16'd12658, 16'd53799, 16'd30640, 16'd32136, 16'd65501, 16'd39342, 16'd3070, 16'd7672, 16'd1564, 16'd10344, 16'd45132, 16'd22514, 16'd3383, 16'd17521, 16'd26315, 16'd20531, 16'd39888, 16'd10365, 16'd4098, 16'd33923, 16'd65189, 16'd10081});
	test_expansion(128'hc5b1998f9b972f93a79e4dd1358b1104, {16'd58084, 16'd63105, 16'd8421, 16'd62557, 16'd24882, 16'd59415, 16'd30457, 16'd42061, 16'd14443, 16'd3484, 16'd25239, 16'd15946, 16'd30186, 16'd2435, 16'd38166, 16'd38305, 16'd11081, 16'd61016, 16'd44912, 16'd36785, 16'd62682, 16'd54082, 16'd6878, 16'd60761, 16'd25711, 16'd63374});
	test_expansion(128'ha9e55631a81f254743fedcb08486f78e, {16'd47819, 16'd54727, 16'd9851, 16'd12721, 16'd24223, 16'd26272, 16'd48846, 16'd43646, 16'd13007, 16'd58796, 16'd55420, 16'd32189, 16'd25407, 16'd52264, 16'd11377, 16'd59107, 16'd39549, 16'd42088, 16'd56067, 16'd61423, 16'd2389, 16'd50171, 16'd7947, 16'd10698, 16'd13203, 16'd52399});
	test_expansion(128'hb64e5444b1a86418eba33afa20fa9992, {16'd26420, 16'd53794, 16'd42848, 16'd3117, 16'd65187, 16'd9319, 16'd37048, 16'd5600, 16'd36441, 16'd10835, 16'd30472, 16'd42469, 16'd7715, 16'd49364, 16'd52071, 16'd35796, 16'd29177, 16'd13221, 16'd59807, 16'd18211, 16'd16704, 16'd44354, 16'd47908, 16'd31570, 16'd20556, 16'd36540});
	test_expansion(128'h22eea582d1e989ae772283e4b438182e, {16'd21117, 16'd36764, 16'd14952, 16'd15685, 16'd47746, 16'd61809, 16'd51336, 16'd25292, 16'd15044, 16'd3711, 16'd21190, 16'd45971, 16'd13043, 16'd60416, 16'd48020, 16'd60183, 16'd49208, 16'd38002, 16'd4064, 16'd41351, 16'd30024, 16'd15366, 16'd10632, 16'd13015, 16'd25264, 16'd62979});
	test_expansion(128'hef030c9b847ba2c22026408cdbc19d07, {16'd20653, 16'd52014, 16'd37471, 16'd61641, 16'd13308, 16'd44795, 16'd35549, 16'd17637, 16'd10238, 16'd64012, 16'd31095, 16'd52058, 16'd5502, 16'd22524, 16'd46536, 16'd16274, 16'd1438, 16'd61792, 16'd3296, 16'd41928, 16'd57311, 16'd50088, 16'd1097, 16'd47172, 16'd19261, 16'd58148});
	test_expansion(128'h71aeb25477b0dac4139a8b9b042fb564, {16'd46906, 16'd53250, 16'd48950, 16'd4004, 16'd6608, 16'd34465, 16'd64219, 16'd63079, 16'd33282, 16'd10272, 16'd41645, 16'd56654, 16'd28364, 16'd16439, 16'd5760, 16'd18710, 16'd45559, 16'd21359, 16'd4563, 16'd22695, 16'd16895, 16'd5161, 16'd55526, 16'd1598, 16'd19179, 16'd16548});
	test_expansion(128'h89e9e97d6abe52421618ff78219417db, {16'd20554, 16'd44481, 16'd7992, 16'd45231, 16'd40653, 16'd16141, 16'd28630, 16'd52504, 16'd63564, 16'd40673, 16'd30642, 16'd16345, 16'd23076, 16'd32009, 16'd14955, 16'd61188, 16'd50030, 16'd64279, 16'd34440, 16'd58529, 16'd5668, 16'd19812, 16'd48917, 16'd22282, 16'd21862, 16'd65350});
	test_expansion(128'hc03f6146d5724b0f5de9e75990871693, {16'd62887, 16'd59534, 16'd30364, 16'd60008, 16'd58342, 16'd40793, 16'd12607, 16'd8460, 16'd57864, 16'd28479, 16'd53427, 16'd60175, 16'd56332, 16'd11507, 16'd33424, 16'd51322, 16'd60704, 16'd9937, 16'd45670, 16'd2378, 16'd59690, 16'd11085, 16'd7799, 16'd1551, 16'd17458, 16'd635});
	test_expansion(128'h738387e1ae3afdf3460a9062d2dbe471, {16'd28911, 16'd62729, 16'd43408, 16'd37884, 16'd48460, 16'd20811, 16'd44301, 16'd18432, 16'd31501, 16'd27230, 16'd51665, 16'd26821, 16'd16437, 16'd16988, 16'd48397, 16'd33844, 16'd48858, 16'd11463, 16'd24938, 16'd63299, 16'd4176, 16'd48290, 16'd14334, 16'd43029, 16'd48816, 16'd34612});
	test_expansion(128'he566220fffafd3fd8af6d1328714a014, {16'd48729, 16'd46333, 16'd20477, 16'd65174, 16'd24277, 16'd9206, 16'd31389, 16'd63314, 16'd59811, 16'd52906, 16'd4017, 16'd53987, 16'd50626, 16'd5990, 16'd36560, 16'd1995, 16'd57661, 16'd34627, 16'd33037, 16'd34654, 16'd45480, 16'd41273, 16'd42437, 16'd28210, 16'd62945, 16'd56122});
	test_expansion(128'hc8c6ef6f680b30f9aa9d1ebdbee4ecd7, {16'd52290, 16'd19947, 16'd34954, 16'd64166, 16'd59380, 16'd41418, 16'd23411, 16'd40516, 16'd46684, 16'd44027, 16'd64121, 16'd51903, 16'd40344, 16'd15915, 16'd21803, 16'd18439, 16'd30878, 16'd4414, 16'd6675, 16'd44247, 16'd34058, 16'd34396, 16'd41015, 16'd46022, 16'd61324, 16'd64201});
	test_expansion(128'hfc99f484d9470fcbc770d521fda48926, {16'd13744, 16'd60927, 16'd17294, 16'd59617, 16'd40888, 16'd32908, 16'd39649, 16'd18584, 16'd24606, 16'd62297, 16'd59580, 16'd45367, 16'd22169, 16'd9774, 16'd62806, 16'd37442, 16'd64084, 16'd4832, 16'd64123, 16'd33670, 16'd8084, 16'd21942, 16'd54662, 16'd48872, 16'd2146, 16'd46786});
	test_expansion(128'h64a972d1c9264fa03546668304a0acd5, {16'd40773, 16'd40472, 16'd33487, 16'd8522, 16'd62611, 16'd47409, 16'd21715, 16'd20939, 16'd40891, 16'd52496, 16'd56956, 16'd13656, 16'd36057, 16'd35923, 16'd44439, 16'd46532, 16'd7948, 16'd53144, 16'd43250, 16'd20731, 16'd64625, 16'd1337, 16'd56336, 16'd29346, 16'd55727, 16'd4563});
	test_expansion(128'hf1fd125edd8658223c52ed045810f6db, {16'd45540, 16'd48695, 16'd2505, 16'd52117, 16'd6442, 16'd61366, 16'd9609, 16'd47736, 16'd37756, 16'd489, 16'd32998, 16'd9729, 16'd32171, 16'd9901, 16'd10272, 16'd41538, 16'd60087, 16'd49379, 16'd26163, 16'd58472, 16'd7970, 16'd45995, 16'd41306, 16'd61487, 16'd60909, 16'd13828});
	test_expansion(128'h6ed539046091088a63d3e673e8371770, {16'd12030, 16'd55360, 16'd60871, 16'd16961, 16'd33615, 16'd18395, 16'd56912, 16'd65488, 16'd8918, 16'd39053, 16'd37142, 16'd38622, 16'd1601, 16'd19485, 16'd29422, 16'd55054, 16'd30571, 16'd36648, 16'd16254, 16'd60836, 16'd12784, 16'd25085, 16'd55206, 16'd50742, 16'd45678, 16'd54005});
	test_expansion(128'h94a0bb9cdb558749020b8a00e6e39320, {16'd20308, 16'd32968, 16'd42182, 16'd18724, 16'd49984, 16'd16781, 16'd59365, 16'd62271, 16'd29793, 16'd34886, 16'd28165, 16'd10261, 16'd25787, 16'd50012, 16'd55380, 16'd13953, 16'd21340, 16'd42197, 16'd1160, 16'd10767, 16'd48988, 16'd61224, 16'd26869, 16'd9514, 16'd53763, 16'd2515});
	test_expansion(128'hf72294dea2f6974595b2d5bc1f4bbaa8, {16'd23696, 16'd21980, 16'd34348, 16'd12272, 16'd39796, 16'd56192, 16'd27479, 16'd12086, 16'd2625, 16'd42458, 16'd5618, 16'd55317, 16'd18839, 16'd590, 16'd53299, 16'd36827, 16'd11088, 16'd26300, 16'd64332, 16'd38909, 16'd33976, 16'd45268, 16'd3952, 16'd24458, 16'd41100, 16'd25437});
	test_expansion(128'h6ff438c0e391517016a79f726a2da316, {16'd38709, 16'd45893, 16'd34912, 16'd20987, 16'd9814, 16'd8624, 16'd58659, 16'd51738, 16'd48603, 16'd55495, 16'd62655, 16'd3503, 16'd29252, 16'd44373, 16'd27436, 16'd38228, 16'd11778, 16'd55604, 16'd59418, 16'd26153, 16'd38414, 16'd16099, 16'd54918, 16'd1215, 16'd59634, 16'd3357});
	test_expansion(128'h37be2191087519a4862857e24c1cd8eb, {16'd64793, 16'd7368, 16'd34867, 16'd12434, 16'd37373, 16'd19340, 16'd7324, 16'd53982, 16'd1731, 16'd56478, 16'd48002, 16'd37828, 16'd54175, 16'd35562, 16'd45307, 16'd44682, 16'd65317, 16'd59213, 16'd32586, 16'd21710, 16'd4925, 16'd34491, 16'd17553, 16'd29787, 16'd58748, 16'd29287});
	test_expansion(128'hb54ccab43a9b15010ee91caaed45ebd9, {16'd18200, 16'd30846, 16'd51372, 16'd23859, 16'd54065, 16'd613, 16'd30973, 16'd20129, 16'd3012, 16'd7313, 16'd40562, 16'd9176, 16'd38674, 16'd26595, 16'd38391, 16'd58711, 16'd25394, 16'd49331, 16'd47839, 16'd5837, 16'd52256, 16'd12494, 16'd58458, 16'd61957, 16'd46044, 16'd30340});
	test_expansion(128'hfeba3976322fa0e2876801d502e2f7b3, {16'd29414, 16'd36741, 16'd81, 16'd1436, 16'd1529, 16'd62804, 16'd7648, 16'd57850, 16'd38127, 16'd44864, 16'd51886, 16'd30850, 16'd61135, 16'd12581, 16'd29506, 16'd65093, 16'd36369, 16'd45723, 16'd33650, 16'd23176, 16'd9604, 16'd54573, 16'd38472, 16'd1052, 16'd54743, 16'd10583});
	test_expansion(128'h3e2b82bdb13bf5ad7342f65fb1829aa2, {16'd4317, 16'd15033, 16'd56549, 16'd5508, 16'd52330, 16'd15857, 16'd40374, 16'd52190, 16'd60704, 16'd526, 16'd60922, 16'd8142, 16'd911, 16'd16300, 16'd37819, 16'd4696, 16'd57162, 16'd14857, 16'd38524, 16'd1409, 16'd32255, 16'd10514, 16'd36750, 16'd51024, 16'd22025, 16'd39750});
	test_expansion(128'hb36d33a7a72677f658a3cf11a9baee8d, {16'd1195, 16'd8076, 16'd61407, 16'd55286, 16'd59779, 16'd8923, 16'd5785, 16'd43055, 16'd48529, 16'd17312, 16'd44931, 16'd43206, 16'd57071, 16'd65312, 16'd33422, 16'd11595, 16'd28032, 16'd706, 16'd37460, 16'd45257, 16'd19584, 16'd36304, 16'd20160, 16'd25716, 16'd45697, 16'd53556});
	test_expansion(128'h0769c4dd79a55b86306464b0c25c9100, {16'd59291, 16'd20608, 16'd33501, 16'd58255, 16'd8236, 16'd26570, 16'd56894, 16'd51189, 16'd27216, 16'd24299, 16'd47940, 16'd58695, 16'd24808, 16'd57789, 16'd59899, 16'd46426, 16'd51860, 16'd60588, 16'd29712, 16'd64448, 16'd18780, 16'd42142, 16'd24960, 16'd53057, 16'd13516, 16'd21526});
	test_expansion(128'h32a4fcf82953d2407d755067ff410905, {16'd14241, 16'd45693, 16'd40661, 16'd65097, 16'd23680, 16'd55535, 16'd21104, 16'd28281, 16'd39871, 16'd47329, 16'd56867, 16'd3557, 16'd47435, 16'd63879, 16'd19844, 16'd30498, 16'd26919, 16'd49988, 16'd4312, 16'd49111, 16'd30709, 16'd20765, 16'd56277, 16'd6486, 16'd23431, 16'd15084});
	test_expansion(128'hbe3b73282379460e6a6d8fafaf564f97, {16'd60861, 16'd8275, 16'd17880, 16'd46760, 16'd42074, 16'd20886, 16'd5306, 16'd3655, 16'd42517, 16'd62330, 16'd56073, 16'd46971, 16'd49532, 16'd63174, 16'd29885, 16'd62107, 16'd46055, 16'd57552, 16'd34934, 16'd32027, 16'd38639, 16'd32911, 16'd60405, 16'd50232, 16'd9171, 16'd12028});
	test_expansion(128'h94fdfd9bbf8f7b654779081f1ed83016, {16'd50630, 16'd61083, 16'd17452, 16'd21585, 16'd56614, 16'd61496, 16'd22254, 16'd60655, 16'd30117, 16'd43084, 16'd50345, 16'd56861, 16'd55684, 16'd526, 16'd59401, 16'd27900, 16'd2468, 16'd11397, 16'd55587, 16'd20302, 16'd36078, 16'd16012, 16'd52205, 16'd44595, 16'd51985, 16'd52800});
	test_expansion(128'hb70ddc7c98b09175af7f6fbe9371def8, {16'd11219, 16'd7737, 16'd50127, 16'd38427, 16'd52766, 16'd51125, 16'd9717, 16'd22599, 16'd59050, 16'd20417, 16'd1590, 16'd59364, 16'd28650, 16'd28641, 16'd532, 16'd36017, 16'd42850, 16'd34402, 16'd54427, 16'd39843, 16'd7591, 16'd53470, 16'd30128, 16'd39169, 16'd6783, 16'd26643});
	test_expansion(128'h4cafa60ab059f90b125dc705cc6d3437, {16'd41378, 16'd22922, 16'd7512, 16'd59830, 16'd23422, 16'd30476, 16'd18810, 16'd48880, 16'd36596, 16'd51391, 16'd31891, 16'd11181, 16'd2076, 16'd36548, 16'd19941, 16'd34932, 16'd10527, 16'd27696, 16'd52058, 16'd1446, 16'd6475, 16'd63809, 16'd42515, 16'd2931, 16'd58514, 16'd47189});
	test_expansion(128'h637d0083f4fe905ae6dcd6b469ae9f75, {16'd60118, 16'd11426, 16'd58823, 16'd19870, 16'd61063, 16'd62501, 16'd25258, 16'd18062, 16'd22375, 16'd58196, 16'd4628, 16'd14582, 16'd37826, 16'd23984, 16'd3371, 16'd64221, 16'd19900, 16'd65381, 16'd30974, 16'd30626, 16'd57744, 16'd18379, 16'd20061, 16'd10761, 16'd13451, 16'd5216});
	test_expansion(128'haaedd12a5292d980b4618248e08313b8, {16'd32369, 16'd31748, 16'd34553, 16'd56709, 16'd22211, 16'd19225, 16'd56177, 16'd31058, 16'd15086, 16'd22675, 16'd34126, 16'd3549, 16'd53651, 16'd877, 16'd26067, 16'd37451, 16'd32258, 16'd34601, 16'd13521, 16'd29118, 16'd50731, 16'd32186, 16'd31089, 16'd51982, 16'd22288, 16'd20431});
	test_expansion(128'hca5c6a735920a7afef98141b9bc79c8f, {16'd10847, 16'd241, 16'd5724, 16'd21356, 16'd21695, 16'd27873, 16'd40291, 16'd61735, 16'd31430, 16'd17027, 16'd63719, 16'd33133, 16'd43366, 16'd24239, 16'd7026, 16'd4697, 16'd27869, 16'd35279, 16'd51355, 16'd29914, 16'd60748, 16'd29589, 16'd33479, 16'd57016, 16'd58782, 16'd18841});
	test_expansion(128'h452865e707061172e26277e2349fc2e8, {16'd25269, 16'd16179, 16'd55631, 16'd45447, 16'd17488, 16'd63514, 16'd42601, 16'd49583, 16'd48795, 16'd46097, 16'd12956, 16'd56077, 16'd11928, 16'd25297, 16'd10701, 16'd51619, 16'd19206, 16'd42529, 16'd15831, 16'd10676, 16'd61802, 16'd25766, 16'd12866, 16'd7874, 16'd53437, 16'd45095});
	test_expansion(128'h90c5fc5973cfcb6dbbd685ed1f012602, {16'd35175, 16'd35819, 16'd49979, 16'd11347, 16'd25190, 16'd13664, 16'd4492, 16'd24349, 16'd26907, 16'd26348, 16'd16468, 16'd49566, 16'd2264, 16'd8657, 16'd64623, 16'd30424, 16'd3755, 16'd27664, 16'd45317, 16'd6134, 16'd12679, 16'd15772, 16'd4447, 16'd46583, 16'd51573, 16'd13921});
	test_expansion(128'he634312d167dd5726dfdd1aa28dd8cf3, {16'd62460, 16'd33058, 16'd57884, 16'd42992, 16'd52853, 16'd29964, 16'd36802, 16'd15295, 16'd60674, 16'd43086, 16'd26363, 16'd61022, 16'd6761, 16'd63777, 16'd481, 16'd55003, 16'd54146, 16'd37974, 16'd38354, 16'd33501, 16'd33248, 16'd37051, 16'd20716, 16'd43649, 16'd44124, 16'd23217});
	test_expansion(128'h40dbb71675841e2b489d9b8f9afa4151, {16'd62585, 16'd40546, 16'd22938, 16'd11751, 16'd56476, 16'd31675, 16'd33235, 16'd51078, 16'd16236, 16'd63531, 16'd8007, 16'd9768, 16'd54112, 16'd26487, 16'd52628, 16'd55522, 16'd41297, 16'd8983, 16'd44057, 16'd29513, 16'd19182, 16'd3198, 16'd8109, 16'd40434, 16'd40471, 16'd11503});
	test_expansion(128'h50a1de14ec9565d55870fc26bf7e1317, {16'd57282, 16'd250, 16'd24504, 16'd36332, 16'd21030, 16'd19673, 16'd11287, 16'd12031, 16'd56912, 16'd48812, 16'd24655, 16'd51333, 16'd23968, 16'd36148, 16'd51608, 16'd13412, 16'd15382, 16'd55775, 16'd43194, 16'd59865, 16'd2727, 16'd32567, 16'd8387, 16'd26313, 16'd49622, 16'd51299});
	test_expansion(128'h26ab3eaeba7af825eb19293f79a6d46d, {16'd21045, 16'd43409, 16'd8173, 16'd3258, 16'd63530, 16'd24164, 16'd26753, 16'd62148, 16'd2932, 16'd11541, 16'd29693, 16'd30369, 16'd5873, 16'd58610, 16'd38525, 16'd34318, 16'd2584, 16'd55696, 16'd58671, 16'd29576, 16'd37743, 16'd24735, 16'd16653, 16'd24028, 16'd307, 16'd56502});
	test_expansion(128'hd4398589f8db637f61266491a8e5272c, {16'd29251, 16'd53532, 16'd36656, 16'd19775, 16'd8474, 16'd34991, 16'd38398, 16'd27932, 16'd9611, 16'd17725, 16'd56040, 16'd7048, 16'd22774, 16'd30304, 16'd21329, 16'd21110, 16'd37678, 16'd560, 16'd52125, 16'd48230, 16'd18851, 16'd18424, 16'd5278, 16'd41748, 16'd12992, 16'd62366});
	test_expansion(128'hdb09c14f7545e8beff898203294930a0, {16'd46538, 16'd11997, 16'd59503, 16'd27751, 16'd17430, 16'd47848, 16'd6325, 16'd63713, 16'd11905, 16'd2198, 16'd40357, 16'd33475, 16'd2570, 16'd17362, 16'd1629, 16'd1480, 16'd65383, 16'd49013, 16'd27152, 16'd37596, 16'd20362, 16'd65412, 16'd56700, 16'd61988, 16'd29829, 16'd51511});
	test_expansion(128'h3f822f9fc4da3971bc479fefc763f9ce, {16'd64199, 16'd12131, 16'd58424, 16'd9353, 16'd4635, 16'd6076, 16'd34746, 16'd41298, 16'd19037, 16'd338, 16'd27786, 16'd5691, 16'd37574, 16'd24089, 16'd19699, 16'd11125, 16'd24036, 16'd8093, 16'd9957, 16'd20188, 16'd36538, 16'd38640, 16'd42588, 16'd21445, 16'd30419, 16'd15967});
	test_expansion(128'h85eec97b573448fb1ad9bd2a9f32bd3c, {16'd21803, 16'd46692, 16'd22555, 16'd51686, 16'd43656, 16'd15453, 16'd15671, 16'd52687, 16'd47320, 16'd65054, 16'd29811, 16'd38562, 16'd34261, 16'd42526, 16'd13137, 16'd10408, 16'd30060, 16'd36863, 16'd31371, 16'd45094, 16'd39634, 16'd43875, 16'd50630, 16'd14323, 16'd16392, 16'd63403});
	test_expansion(128'h285c2f668260117cdb33c523b0b66e8e, {16'd36363, 16'd7646, 16'd51476, 16'd11671, 16'd60837, 16'd37533, 16'd61272, 16'd30250, 16'd61929, 16'd14125, 16'd29932, 16'd53331, 16'd25304, 16'd1393, 16'd30819, 16'd22001, 16'd18994, 16'd17101, 16'd27818, 16'd64220, 16'd283, 16'd21758, 16'd26229, 16'd8101, 16'd32337, 16'd8929});
	test_expansion(128'h4754bdb4a52e1701aaaf6f40b6c5a582, {16'd31856, 16'd52852, 16'd4186, 16'd27771, 16'd13534, 16'd15371, 16'd18116, 16'd44152, 16'd24681, 16'd34797, 16'd5845, 16'd44393, 16'd36953, 16'd46525, 16'd26948, 16'd42327, 16'd50323, 16'd23424, 16'd58925, 16'd64327, 16'd13577, 16'd26710, 16'd14519, 16'd49291, 16'd48451, 16'd48529});
	test_expansion(128'hcb48dc10fbb3d22e04a7ab1190081d32, {16'd60290, 16'd25259, 16'd42620, 16'd37578, 16'd11680, 16'd41562, 16'd11880, 16'd4581, 16'd52024, 16'd9223, 16'd20060, 16'd41985, 16'd5217, 16'd15558, 16'd29812, 16'd48196, 16'd52006, 16'd22173, 16'd6512, 16'd50696, 16'd8324, 16'd51640, 16'd18086, 16'd9130, 16'd12372, 16'd23055});
	test_expansion(128'ha15e0b33920eb6421daf3445c4e595cc, {16'd62979, 16'd4311, 16'd25058, 16'd29355, 16'd45699, 16'd41145, 16'd3110, 16'd20539, 16'd44966, 16'd4016, 16'd53580, 16'd43619, 16'd56072, 16'd59957, 16'd52716, 16'd6544, 16'd60293, 16'd55160, 16'd41055, 16'd63270, 16'd57461, 16'd37680, 16'd59050, 16'd42233, 16'd62931, 16'd58105});
	test_expansion(128'he270845d3afda34a7c869058385df4d8, {16'd4001, 16'd21064, 16'd20726, 16'd49941, 16'd6458, 16'd23216, 16'd17708, 16'd44171, 16'd34084, 16'd44547, 16'd18143, 16'd20629, 16'd37929, 16'd42140, 16'd31876, 16'd10829, 16'd23180, 16'd21944, 16'd40253, 16'd56307, 16'd53661, 16'd22499, 16'd14455, 16'd3598, 16'd28224, 16'd45978});
	test_expansion(128'h8eaf919ed1c968f2ca0433366166b33e, {16'd7962, 16'd48750, 16'd12922, 16'd17023, 16'd28472, 16'd19226, 16'd52052, 16'd20607, 16'd50611, 16'd6690, 16'd15470, 16'd4006, 16'd35685, 16'd57009, 16'd57641, 16'd47792, 16'd11271, 16'd46787, 16'd49552, 16'd54793, 16'd10565, 16'd62993, 16'd8964, 16'd49909, 16'd62267, 16'd42307});
	test_expansion(128'hbaaeddba05bd2078d28a6ee48160dbd1, {16'd27452, 16'd12619, 16'd7187, 16'd63305, 16'd53230, 16'd14232, 16'd26960, 16'd29397, 16'd10449, 16'd51009, 16'd5213, 16'd13563, 16'd26413, 16'd33092, 16'd62396, 16'd60067, 16'd65435, 16'd725, 16'd31491, 16'd49303, 16'd11840, 16'd45470, 16'd50177, 16'd56476, 16'd55468, 16'd46996});
	test_expansion(128'h882b1acd63b15bf19ca7292ac06a9319, {16'd4885, 16'd57731, 16'd60927, 16'd42067, 16'd53646, 16'd3240, 16'd33709, 16'd853, 16'd3317, 16'd45991, 16'd48656, 16'd42163, 16'd19148, 16'd38243, 16'd30627, 16'd18892, 16'd58630, 16'd3386, 16'd51376, 16'd29946, 16'd46519, 16'd49768, 16'd1909, 16'd7489, 16'd60649, 16'd35643});
	test_expansion(128'h0f3214853be320af05d7ecbb8ff896e6, {16'd16201, 16'd20685, 16'd8671, 16'd38481, 16'd13353, 16'd58947, 16'd53468, 16'd9564, 16'd33635, 16'd55518, 16'd16206, 16'd25974, 16'd10923, 16'd40414, 16'd28471, 16'd29258, 16'd34180, 16'd34476, 16'd22296, 16'd65358, 16'd65353, 16'd17826, 16'd52382, 16'd48678, 16'd35703, 16'd57701});
	test_expansion(128'h9f74ed99958d7d278e676ec3bdb6b81a, {16'd27702, 16'd14465, 16'd44898, 16'd43626, 16'd15204, 16'd2106, 16'd2158, 16'd20850, 16'd64500, 16'd48674, 16'd31166, 16'd25084, 16'd65073, 16'd2776, 16'd30659, 16'd14725, 16'd59451, 16'd51451, 16'd37157, 16'd17260, 16'd60810, 16'd50975, 16'd63992, 16'd40532, 16'd64570, 16'd16908});
	test_expansion(128'h6e0a15d11a7aed3701b958102e474bcb, {16'd62067, 16'd37209, 16'd37791, 16'd23399, 16'd14504, 16'd58767, 16'd48661, 16'd20, 16'd57362, 16'd15275, 16'd31187, 16'd25519, 16'd18192, 16'd25336, 16'd22709, 16'd13339, 16'd25043, 16'd58087, 16'd20557, 16'd37601, 16'd20739, 16'd18305, 16'd59132, 16'd6295, 16'd44445, 16'd39096});
	test_expansion(128'h06512fb93afd91acc88a045751934513, {16'd4268, 16'd44852, 16'd40912, 16'd33698, 16'd21629, 16'd21830, 16'd19495, 16'd18061, 16'd26289, 16'd4104, 16'd40225, 16'd64377, 16'd62697, 16'd33622, 16'd33942, 16'd31735, 16'd24575, 16'd41667, 16'd55922, 16'd55308, 16'd7305, 16'd25429, 16'd23922, 16'd37335, 16'd65473, 16'd21689});
	test_expansion(128'h749372edb741470a840c65b920038b2f, {16'd40570, 16'd42150, 16'd38479, 16'd9532, 16'd642, 16'd40511, 16'd39029, 16'd60857, 16'd59349, 16'd43814, 16'd45799, 16'd28620, 16'd45705, 16'd60926, 16'd50196, 16'd22639, 16'd30188, 16'd21057, 16'd28483, 16'd634, 16'd60342, 16'd20692, 16'd16682, 16'd31188, 16'd39070, 16'd8325});
	test_expansion(128'ha9e0e4951dfc02ad621200a9421a1320, {16'd11293, 16'd54694, 16'd54165, 16'd26279, 16'd25420, 16'd36943, 16'd20541, 16'd27492, 16'd24823, 16'd5094, 16'd57496, 16'd57550, 16'd64876, 16'd46362, 16'd18457, 16'd43469, 16'd63628, 16'd2558, 16'd14262, 16'd58647, 16'd33939, 16'd24086, 16'd21378, 16'd43109, 16'd64326, 16'd16773});
	test_expansion(128'h4ac23b0d6ac5f14aff3bd8f3ebe904e3, {16'd25460, 16'd50085, 16'd51061, 16'd11034, 16'd24383, 16'd4198, 16'd54918, 16'd10489, 16'd41021, 16'd5250, 16'd62222, 16'd60960, 16'd49223, 16'd46952, 16'd17880, 16'd4201, 16'd13672, 16'd44059, 16'd52202, 16'd64483, 16'd21332, 16'd42476, 16'd4043, 16'd47701, 16'd5117, 16'd15429});
	test_expansion(128'heb36df81efba08b0fbd0809a247bc540, {16'd35446, 16'd62377, 16'd47636, 16'd28253, 16'd9034, 16'd53060, 16'd7314, 16'd36708, 16'd46848, 16'd60189, 16'd36823, 16'd41668, 16'd45348, 16'd52822, 16'd55882, 16'd34777, 16'd29640, 16'd18405, 16'd6178, 16'd31044, 16'd56240, 16'd43038, 16'd64598, 16'd45397, 16'd57994, 16'd16960});
	test_expansion(128'h8dc42cf89992e43ea37e9d1e2283c197, {16'd10986, 16'd17458, 16'd51075, 16'd56702, 16'd21003, 16'd52468, 16'd64716, 16'd38238, 16'd61504, 16'd10868, 16'd25599, 16'd11751, 16'd10926, 16'd42084, 16'd1700, 16'd57346, 16'd52203, 16'd51235, 16'd24893, 16'd25010, 16'd3711, 16'd29653, 16'd19270, 16'd5585, 16'd57986, 16'd39301});
	test_expansion(128'h898efabc95649bdc76533b06212fe9c4, {16'd55966, 16'd36494, 16'd53653, 16'd8108, 16'd26596, 16'd42329, 16'd63048, 16'd23248, 16'd10001, 16'd12422, 16'd61867, 16'd54054, 16'd10871, 16'd64044, 16'd22017, 16'd20219, 16'd38604, 16'd6354, 16'd64229, 16'd65334, 16'd48786, 16'd32458, 16'd1167, 16'd15085, 16'd23215, 16'd11188});
	test_expansion(128'hb92ea0306b552c8bf8e70d8d8e0f82dc, {16'd5932, 16'd51074, 16'd46896, 16'd4035, 16'd26603, 16'd44109, 16'd27301, 16'd55376, 16'd22253, 16'd9771, 16'd19322, 16'd35718, 16'd47083, 16'd51026, 16'd4765, 16'd30990, 16'd17727, 16'd41533, 16'd1812, 16'd16970, 16'd28105, 16'd14040, 16'd56650, 16'd12608, 16'd63529, 16'd49058});
	test_expansion(128'h76a3c7ae93f4bcf0a35b68335d3f1f56, {16'd8663, 16'd32693, 16'd20886, 16'd8232, 16'd22114, 16'd40550, 16'd32092, 16'd1880, 16'd32242, 16'd8908, 16'd58778, 16'd58473, 16'd13991, 16'd58113, 16'd14782, 16'd49711, 16'd50954, 16'd45329, 16'd30938, 16'd45416, 16'd53985, 16'd63351, 16'd16986, 16'd42380, 16'd29168, 16'd44816});
	test_expansion(128'h9768fb80aeeded29b9be7342b9b85781, {16'd56516, 16'd53857, 16'd51338, 16'd32643, 16'd848, 16'd41055, 16'd21512, 16'd46764, 16'd14510, 16'd8880, 16'd37774, 16'd65460, 16'd19318, 16'd42957, 16'd39954, 16'd41161, 16'd56871, 16'd5900, 16'd56587, 16'd41884, 16'd56996, 16'd24454, 16'd26220, 16'd40896, 16'd43794, 16'd59760});
	test_expansion(128'hc19b41495453f2a892010a57fd095035, {16'd4481, 16'd42023, 16'd54167, 16'd58847, 16'd17291, 16'd22228, 16'd37765, 16'd55488, 16'd57628, 16'd31593, 16'd1607, 16'd9337, 16'd22189, 16'd54592, 16'd15622, 16'd36341, 16'd41932, 16'd8707, 16'd24420, 16'd13631, 16'd28775, 16'd49095, 16'd14253, 16'd9737, 16'd15983, 16'd3495});
	test_expansion(128'h12174bcb96ecc60db4dd6c4f480123dc, {16'd31466, 16'd59193, 16'd23855, 16'd34429, 16'd30059, 16'd23359, 16'd16550, 16'd10929, 16'd39421, 16'd16546, 16'd35751, 16'd41292, 16'd52069, 16'd20979, 16'd9103, 16'd4240, 16'd25687, 16'd41669, 16'd41163, 16'd63706, 16'd14513, 16'd58845, 16'd58033, 16'd1106, 16'd52695, 16'd45807});
	test_expansion(128'hb2ff4f4f746aa02b34b7f26076e7a6b2, {16'd36266, 16'd30434, 16'd63080, 16'd53715, 16'd21216, 16'd24622, 16'd38316, 16'd38224, 16'd16742, 16'd10508, 16'd38517, 16'd21242, 16'd48202, 16'd3709, 16'd7699, 16'd24570, 16'd17508, 16'd15100, 16'd26634, 16'd20787, 16'd7539, 16'd46607, 16'd56410, 16'd7916, 16'd2765, 16'd56800});
	test_expansion(128'h3e658346f4c49709d2fe4f528d4b7b37, {16'd62501, 16'd23412, 16'd15571, 16'd38613, 16'd50367, 16'd38769, 16'd46545, 16'd61364, 16'd35043, 16'd28043, 16'd9210, 16'd13157, 16'd38658, 16'd59248, 16'd41435, 16'd28183, 16'd18611, 16'd9686, 16'd5152, 16'd34263, 16'd17693, 16'd13396, 16'd22587, 16'd29782, 16'd60233, 16'd19745});
	test_expansion(128'he3a124271f42cdd83c3a8d98e1b51875, {16'd46545, 16'd8718, 16'd17221, 16'd30451, 16'd50069, 16'd13734, 16'd31181, 16'd27648, 16'd48772, 16'd42488, 16'd19612, 16'd39550, 16'd54456, 16'd38614, 16'd58231, 16'd59040, 16'd34373, 16'd23662, 16'd35079, 16'd5650, 16'd23320, 16'd63726, 16'd24300, 16'd45259, 16'd32762, 16'd9819});
	test_expansion(128'hd78234399ae8fae50f1ddd9f4294347c, {16'd29408, 16'd27176, 16'd26083, 16'd44977, 16'd10360, 16'd37278, 16'd30562, 16'd55926, 16'd1586, 16'd34345, 16'd42718, 16'd45465, 16'd50913, 16'd5854, 16'd19789, 16'd53670, 16'd53802, 16'd31597, 16'd35157, 16'd59682, 16'd19893, 16'd5305, 16'd13421, 16'd50943, 16'd18934, 16'd23808});
	test_expansion(128'h666c0a61859f5aa37793230f0521f273, {16'd20060, 16'd34428, 16'd21355, 16'd26401, 16'd32941, 16'd65118, 16'd47130, 16'd748, 16'd15958, 16'd59042, 16'd64072, 16'd2776, 16'd13300, 16'd47491, 16'd44688, 16'd36832, 16'd46724, 16'd52444, 16'd63729, 16'd53455, 16'd42866, 16'd3126, 16'd50705, 16'd10093, 16'd6709, 16'd1369});
	test_expansion(128'hd582daedf340c38c4fba8e990daba0d6, {16'd44715, 16'd26756, 16'd1238, 16'd19845, 16'd10200, 16'd13213, 16'd6222, 16'd14311, 16'd4631, 16'd39667, 16'd4441, 16'd8484, 16'd44400, 16'd764, 16'd812, 16'd64735, 16'd41586, 16'd6652, 16'd55152, 16'd63582, 16'd30208, 16'd8887, 16'd15268, 16'd11821, 16'd7881, 16'd64109});
	test_expansion(128'hc3e95ea3d4b79a96ba43a9cd58247d1f, {16'd41537, 16'd13931, 16'd26258, 16'd17768, 16'd29820, 16'd60349, 16'd65181, 16'd49177, 16'd8515, 16'd2283, 16'd22868, 16'd29615, 16'd23036, 16'd31222, 16'd16968, 16'd45592, 16'd34304, 16'd3292, 16'd47033, 16'd38344, 16'd3546, 16'd9138, 16'd12082, 16'd19154, 16'd45834, 16'd52822});
	test_expansion(128'hac98ccaa3298b7654afc691f5b28948d, {16'd21481, 16'd36142, 16'd3747, 16'd10782, 16'd52273, 16'd51348, 16'd62958, 16'd12212, 16'd64835, 16'd3691, 16'd13343, 16'd55147, 16'd27472, 16'd10682, 16'd2005, 16'd40049, 16'd28383, 16'd58816, 16'd62777, 16'd60696, 16'd3672, 16'd43679, 16'd13215, 16'd34275, 16'd64700, 16'd60604});
	test_expansion(128'h6b9524b31df44e0ae6c2acde5740e69b, {16'd30211, 16'd30222, 16'd20309, 16'd62873, 16'd39231, 16'd3886, 16'd50385, 16'd62369, 16'd53689, 16'd52411, 16'd21048, 16'd34268, 16'd44965, 16'd48631, 16'd22813, 16'd50852, 16'd63992, 16'd42321, 16'd10022, 16'd3058, 16'd16016, 16'd37158, 16'd7839, 16'd62199, 16'd42577, 16'd36103});
	test_expansion(128'h164ec1a3c26135fe032cad987ce38f07, {16'd38122, 16'd24704, 16'd5549, 16'd6871, 16'd47511, 16'd54308, 16'd29394, 16'd2978, 16'd38531, 16'd64456, 16'd59862, 16'd56096, 16'd60903, 16'd3116, 16'd29239, 16'd60625, 16'd8219, 16'd58314, 16'd45817, 16'd44813, 16'd60908, 16'd40984, 16'd63256, 16'd35995, 16'd20643, 16'd11588});
	test_expansion(128'hd42496e3eff717a63947ee6333cd02b3, {16'd52428, 16'd58328, 16'd1008, 16'd9210, 16'd54389, 16'd51972, 16'd30723, 16'd23720, 16'd1495, 16'd9422, 16'd6821, 16'd19531, 16'd24123, 16'd33501, 16'd49135, 16'd37406, 16'd21747, 16'd28143, 16'd15012, 16'd19684, 16'd3563, 16'd58726, 16'd42917, 16'd53378, 16'd27825, 16'd23913});
	test_expansion(128'h10d416d52fd11af5a7ff24263a95b20d, {16'd6581, 16'd17560, 16'd29263, 16'd20630, 16'd52072, 16'd40493, 16'd60763, 16'd18971, 16'd4093, 16'd15159, 16'd62906, 16'd13462, 16'd29356, 16'd51180, 16'd32932, 16'd40646, 16'd40724, 16'd15917, 16'd44760, 16'd55419, 16'd2883, 16'd65290, 16'd11729, 16'd10912, 16'd2225, 16'd61814});
	test_expansion(128'h7d40aee5731b6e98943ab83aadf16a55, {16'd49488, 16'd1755, 16'd22690, 16'd36135, 16'd35687, 16'd5164, 16'd577, 16'd48042, 16'd41408, 16'd58131, 16'd28780, 16'd30321, 16'd61540, 16'd57242, 16'd11159, 16'd32420, 16'd45134, 16'd17044, 16'd14745, 16'd32471, 16'd58833, 16'd8377, 16'd36981, 16'd25180, 16'd57692, 16'd33208});
	test_expansion(128'h34bfac78a8768a709caf43a626e9ea50, {16'd15626, 16'd54128, 16'd58218, 16'd37259, 16'd24937, 16'd51452, 16'd37290, 16'd60722, 16'd21334, 16'd60109, 16'd60813, 16'd45921, 16'd10975, 16'd1900, 16'd5310, 16'd5311, 16'd46185, 16'd28674, 16'd44154, 16'd33450, 16'd34280, 16'd50214, 16'd24751, 16'd54175, 16'd33763, 16'd9110});
	test_expansion(128'h69aa2774403b0cf03f3a77225b60a1ad, {16'd2804, 16'd51912, 16'd18525, 16'd52463, 16'd10283, 16'd37306, 16'd65024, 16'd12899, 16'd20450, 16'd38981, 16'd32367, 16'd6510, 16'd38571, 16'd15341, 16'd36237, 16'd21650, 16'd17960, 16'd41384, 16'd54460, 16'd39742, 16'd36110, 16'd34719, 16'd50020, 16'd20856, 16'd2099, 16'd33946});
	test_expansion(128'h9bd09a3e9d634df8cf8c24a81c59c97c, {16'd27188, 16'd65003, 16'd8662, 16'd58037, 16'd53626, 16'd4340, 16'd5379, 16'd59496, 16'd63784, 16'd14647, 16'd20717, 16'd14374, 16'd4302, 16'd8390, 16'd9076, 16'd58070, 16'd4827, 16'd88, 16'd31471, 16'd2387, 16'd55655, 16'd37490, 16'd13543, 16'd47147, 16'd2403, 16'd40609});
	test_expansion(128'hcb938fc60b390ab0aaa3cf82660e26b5, {16'd8534, 16'd22195, 16'd12320, 16'd1189, 16'd16800, 16'd8880, 16'd55790, 16'd22053, 16'd29440, 16'd65406, 16'd8235, 16'd43516, 16'd6184, 16'd8410, 16'd14252, 16'd62431, 16'd59469, 16'd60962, 16'd32820, 16'd47251, 16'd2735, 16'd26538, 16'd10125, 16'd18967, 16'd50807, 16'd18671});
	test_expansion(128'h82a37a44a6f6b1ed72c74ad227b01d4c, {16'd7562, 16'd43638, 16'd21267, 16'd47209, 16'd63852, 16'd36125, 16'd24576, 16'd11836, 16'd1393, 16'd54555, 16'd36647, 16'd64917, 16'd24647, 16'd62759, 16'd54403, 16'd29446, 16'd872, 16'd42602, 16'd40062, 16'd11363, 16'd14908, 16'd24236, 16'd50180, 16'd61573, 16'd13976, 16'd61308});
	test_expansion(128'h1750c583e186660bcc0286c52997e3ac, {16'd41796, 16'd31813, 16'd6226, 16'd17550, 16'd21962, 16'd40009, 16'd10756, 16'd34015, 16'd40635, 16'd10089, 16'd33553, 16'd55820, 16'd9972, 16'd6579, 16'd64582, 16'd39015, 16'd61629, 16'd1149, 16'd63942, 16'd11824, 16'd58133, 16'd46825, 16'd40998, 16'd59534, 16'd35088, 16'd17747});
	test_expansion(128'h4dc9fe5455ada40946121c386e4e2fd3, {16'd18423, 16'd55119, 16'd28914, 16'd16312, 16'd30736, 16'd50188, 16'd47156, 16'd60039, 16'd29583, 16'd15792, 16'd59036, 16'd4967, 16'd38509, 16'd2017, 16'd15960, 16'd9740, 16'd24991, 16'd36835, 16'd24606, 16'd33874, 16'd63167, 16'd25785, 16'd53070, 16'd6048, 16'd35189, 16'd27557});
	test_expansion(128'hbcc3ae9168ef6e62855390c469e8fdf4, {16'd27129, 16'd59203, 16'd15752, 16'd58144, 16'd46558, 16'd45520, 16'd32060, 16'd1927, 16'd26859, 16'd59378, 16'd13204, 16'd43810, 16'd7312, 16'd41635, 16'd42195, 16'd62486, 16'd31889, 16'd35763, 16'd38421, 16'd22725, 16'd65269, 16'd53818, 16'd44615, 16'd37004, 16'd674, 16'd12093});
	test_expansion(128'h52a644d0f3ebf90fc17ec564d4b30997, {16'd19860, 16'd61425, 16'd54126, 16'd39292, 16'd14480, 16'd320, 16'd38642, 16'd12259, 16'd48503, 16'd35013, 16'd2019, 16'd10958, 16'd53143, 16'd3613, 16'd49585, 16'd7310, 16'd23863, 16'd26965, 16'd33502, 16'd34880, 16'd27238, 16'd48439, 16'd57898, 16'd13328, 16'd64598, 16'd52420});
	test_expansion(128'hea504d47b217e947b300174431e87730, {16'd32033, 16'd51578, 16'd53644, 16'd50526, 16'd27223, 16'd8804, 16'd64793, 16'd11960, 16'd9464, 16'd36983, 16'd40342, 16'd26860, 16'd22741, 16'd46189, 16'd2655, 16'd5513, 16'd60079, 16'd61664, 16'd42395, 16'd4062, 16'd49797, 16'd7897, 16'd31879, 16'd28956, 16'd43690, 16'd41524});
	test_expansion(128'h23e598ea746a8a869107511f886a103b, {16'd36952, 16'd58706, 16'd5613, 16'd51328, 16'd11000, 16'd29798, 16'd18197, 16'd4910, 16'd37352, 16'd63206, 16'd7952, 16'd41560, 16'd56839, 16'd43377, 16'd13729, 16'd26099, 16'd39564, 16'd38009, 16'd31990, 16'd3812, 16'd27780, 16'd57258, 16'd48565, 16'd57536, 16'd48962, 16'd44463});
	test_expansion(128'h830804028134ceb027a01306e8acbb39, {16'd18423, 16'd12439, 16'd1364, 16'd578, 16'd60118, 16'd29083, 16'd65339, 16'd64413, 16'd1540, 16'd10608, 16'd40478, 16'd41695, 16'd32864, 16'd35199, 16'd64533, 16'd5290, 16'd2977, 16'd47009, 16'd44092, 16'd37101, 16'd10070, 16'd5448, 16'd18292, 16'd43125, 16'd1670, 16'd39583});
	test_expansion(128'h7cf51ef6455eedf36b9bd3add45273b1, {16'd36350, 16'd56003, 16'd32063, 16'd698, 16'd52200, 16'd33417, 16'd31476, 16'd51878, 16'd56088, 16'd14777, 16'd14180, 16'd58094, 16'd60419, 16'd5606, 16'd12894, 16'd42248, 16'd19420, 16'd23264, 16'd21015, 16'd53063, 16'd19440, 16'd42319, 16'd35224, 16'd19180, 16'd12353, 16'd33344});
	test_expansion(128'he9b1fb220f51b58e7c6e0de1228f68fd, {16'd19274, 16'd43056, 16'd52979, 16'd1032, 16'd10262, 16'd6857, 16'd54635, 16'd30610, 16'd25950, 16'd46174, 16'd3130, 16'd53384, 16'd44178, 16'd52798, 16'd14412, 16'd49724, 16'd45631, 16'd20703, 16'd48038, 16'd11976, 16'd45121, 16'd30842, 16'd16401, 16'd45598, 16'd9747, 16'd60524});
	test_expansion(128'h1cafe7bb437dc96a4c8537493679f4fe, {16'd12167, 16'd10138, 16'd30157, 16'd2798, 16'd44063, 16'd59605, 16'd9124, 16'd64350, 16'd17979, 16'd8568, 16'd48020, 16'd6568, 16'd47750, 16'd22923, 16'd42538, 16'd31574, 16'd45909, 16'd19069, 16'd52613, 16'd59206, 16'd27473, 16'd30455, 16'd27279, 16'd55097, 16'd15679, 16'd10761});
	test_expansion(128'h4ed445b9fda9c90bf164a7c6762ab852, {16'd26029, 16'd41015, 16'd65349, 16'd16440, 16'd24223, 16'd51628, 16'd41695, 16'd23220, 16'd38393, 16'd58986, 16'd41251, 16'd14797, 16'd53034, 16'd19247, 16'd44354, 16'd2489, 16'd25507, 16'd26003, 16'd20905, 16'd12387, 16'd8580, 16'd35724, 16'd65340, 16'd33530, 16'd29914, 16'd59092});
	test_expansion(128'h048d0fdc3c7a19036fd0aae296636cb9, {16'd64547, 16'd50014, 16'd25140, 16'd49675, 16'd41465, 16'd52548, 16'd62055, 16'd63592, 16'd38545, 16'd54546, 16'd58359, 16'd29957, 16'd51491, 16'd59893, 16'd51926, 16'd40467, 16'd63587, 16'd6024, 16'd51530, 16'd61961, 16'd21736, 16'd2856, 16'd49022, 16'd47529, 16'd32320, 16'd6592});
	test_expansion(128'h3615833aaec8f38e6aac29504189e9e5, {16'd2976, 16'd25251, 16'd36901, 16'd1792, 16'd47552, 16'd65473, 16'd20967, 16'd11413, 16'd16359, 16'd30553, 16'd53224, 16'd37687, 16'd38877, 16'd60979, 16'd46710, 16'd45574, 16'd51062, 16'd2834, 16'd5390, 16'd51307, 16'd37166, 16'd33758, 16'd18330, 16'd17810, 16'd14146, 16'd55496});
	test_expansion(128'hc04e70e40e399c7395a61bcc3b598451, {16'd24067, 16'd41442, 16'd46316, 16'd49860, 16'd38411, 16'd10630, 16'd26470, 16'd16508, 16'd31942, 16'd9981, 16'd55020, 16'd52982, 16'd17446, 16'd31370, 16'd3214, 16'd56644, 16'd19037, 16'd39009, 16'd29592, 16'd27586, 16'd28086, 16'd40074, 16'd7510, 16'd7993, 16'd48262, 16'd50276});
	test_expansion(128'h70dd70fddc34fba2404b8f2ea90a7682, {16'd27622, 16'd55705, 16'd16686, 16'd42170, 16'd20282, 16'd11617, 16'd55949, 16'd17229, 16'd35058, 16'd52680, 16'd649, 16'd14258, 16'd22215, 16'd59924, 16'd31089, 16'd54839, 16'd38791, 16'd59156, 16'd7871, 16'd5981, 16'd11147, 16'd8319, 16'd47320, 16'd28928, 16'd26032, 16'd24370});
	test_expansion(128'h4b5945aa84dc761ed6eaaa14dd7fcadc, {16'd14466, 16'd23431, 16'd15732, 16'd44479, 16'd40858, 16'd51302, 16'd10932, 16'd60273, 16'd36286, 16'd39626, 16'd49668, 16'd38198, 16'd12461, 16'd5703, 16'd58180, 16'd19040, 16'd43093, 16'd55770, 16'd44311, 16'd49105, 16'd59226, 16'd44959, 16'd7961, 16'd39208, 16'd41891, 16'd929});
	test_expansion(128'hdb99bf55dd314769e3cdc143da809bcf, {16'd9425, 16'd59920, 16'd30956, 16'd20927, 16'd50928, 16'd18986, 16'd55301, 16'd8135, 16'd8050, 16'd10611, 16'd10668, 16'd54660, 16'd7201, 16'd45967, 16'd59944, 16'd21275, 16'd15199, 16'd31407, 16'd53221, 16'd60345, 16'd3635, 16'd19981, 16'd56061, 16'd3873, 16'd42575, 16'd52769});
	test_expansion(128'hd013015977ce2bffcc4cecbea9377d7b, {16'd2005, 16'd41603, 16'd9595, 16'd24323, 16'd57218, 16'd3505, 16'd49704, 16'd33154, 16'd21836, 16'd41370, 16'd26835, 16'd25396, 16'd43488, 16'd24980, 16'd60009, 16'd50940, 16'd16824, 16'd43873, 16'd31248, 16'd64948, 16'd3397, 16'd37879, 16'd43801, 16'd14355, 16'd1295, 16'd57756});
	test_expansion(128'h7c8ff0bb7a822b3b67721f1967018d28, {16'd57266, 16'd32179, 16'd12638, 16'd15155, 16'd19082, 16'd64810, 16'd31896, 16'd6608, 16'd41282, 16'd44502, 16'd27747, 16'd52532, 16'd36062, 16'd17233, 16'd37702, 16'd9033, 16'd41045, 16'd60970, 16'd1312, 16'd62913, 16'd8351, 16'd44488, 16'd61179, 16'd34806, 16'd8754, 16'd65329});
	test_expansion(128'hd737b102e5068a538f6e7a007ee4b4ad, {16'd42295, 16'd53870, 16'd25502, 16'd51009, 16'd43473, 16'd51411, 16'd9804, 16'd4623, 16'd24932, 16'd34307, 16'd43820, 16'd64499, 16'd54046, 16'd34121, 16'd28278, 16'd60330, 16'd47567, 16'd31507, 16'd540, 16'd64978, 16'd43899, 16'd757, 16'd10008, 16'd41299, 16'd45469, 16'd40048});
	test_expansion(128'h5138a8baa469fbacbdffecd74de3b662, {16'd11951, 16'd13061, 16'd2691, 16'd22309, 16'd50598, 16'd37432, 16'd59658, 16'd28920, 16'd28329, 16'd24836, 16'd8380, 16'd64078, 16'd51935, 16'd49076, 16'd33378, 16'd18944, 16'd45704, 16'd6476, 16'd46904, 16'd20496, 16'd11993, 16'd890, 16'd49584, 16'd51310, 16'd58810, 16'd56336});
	test_expansion(128'h8dcd642a568e73e5264bc2883ab3d0cc, {16'd27995, 16'd57655, 16'd35532, 16'd29058, 16'd18173, 16'd42096, 16'd13857, 16'd28505, 16'd51817, 16'd5486, 16'd18003, 16'd20280, 16'd59060, 16'd37702, 16'd54560, 16'd54699, 16'd34297, 16'd52836, 16'd39798, 16'd21953, 16'd34092, 16'd14509, 16'd60647, 16'd15918, 16'd33867, 16'd20192});
	test_expansion(128'h48fb4a952ca7ada627ed0682a2d59a2e, {16'd34559, 16'd17764, 16'd49773, 16'd29000, 16'd10195, 16'd44208, 16'd10348, 16'd15817, 16'd3223, 16'd64884, 16'd17257, 16'd4519, 16'd13666, 16'd25302, 16'd6119, 16'd32981, 16'd17704, 16'd54795, 16'd49476, 16'd34754, 16'd57225, 16'd14410, 16'd23790, 16'd134, 16'd12284, 16'd57640});
	test_expansion(128'h1ebda9ba5d49542a6feff69d08a09060, {16'd55983, 16'd23968, 16'd60021, 16'd4375, 16'd49879, 16'd11250, 16'd35351, 16'd18632, 16'd3933, 16'd52381, 16'd6677, 16'd39633, 16'd7108, 16'd2690, 16'd46698, 16'd3941, 16'd29342, 16'd10016, 16'd7323, 16'd50337, 16'd12643, 16'd3841, 16'd40116, 16'd59988, 16'd32409, 16'd46270});
	test_expansion(128'hee5aa23b22f7b9e53df44b58375bc621, {16'd30968, 16'd19918, 16'd6115, 16'd32355, 16'd58544, 16'd33689, 16'd53974, 16'd41217, 16'd26997, 16'd56514, 16'd39156, 16'd52230, 16'd5911, 16'd40679, 16'd27906, 16'd28489, 16'd22767, 16'd14490, 16'd63613, 16'd19414, 16'd34628, 16'd56026, 16'd39616, 16'd34654, 16'd23557, 16'd14658});
	test_expansion(128'hf98a03462310895403c79b865e56c376, {16'd19492, 16'd19052, 16'd38975, 16'd32640, 16'd54018, 16'd59256, 16'd23882, 16'd63371, 16'd35219, 16'd9443, 16'd59488, 16'd21699, 16'd11524, 16'd4421, 16'd10260, 16'd60991, 16'd22136, 16'd61457, 16'd51987, 16'd64256, 16'd15663, 16'd18480, 16'd60947, 16'd56073, 16'd36527, 16'd6408});
	test_expansion(128'h74cd9065d360eadab0cc306c73373c37, {16'd59330, 16'd24693, 16'd28489, 16'd23157, 16'd60149, 16'd46414, 16'd14480, 16'd12273, 16'd19184, 16'd8321, 16'd7016, 16'd18667, 16'd52764, 16'd38955, 16'd25211, 16'd55452, 16'd25279, 16'd59008, 16'd25353, 16'd47915, 16'd47053, 16'd48732, 16'd51351, 16'd26551, 16'd49543, 16'd25841});
	test_expansion(128'he96e988c9ef3fc7e50eb4748a17c1c1b, {16'd52261, 16'd49431, 16'd11551, 16'd46727, 16'd23352, 16'd51148, 16'd12830, 16'd35424, 16'd56206, 16'd50080, 16'd34793, 16'd12157, 16'd63469, 16'd49113, 16'd33561, 16'd37563, 16'd62011, 16'd49303, 16'd11213, 16'd28012, 16'd13242, 16'd7058, 16'd57338, 16'd14653, 16'd12936, 16'd11918});
	test_expansion(128'h0516da5b4d49ca3063ca710d39d4fb5a, {16'd32964, 16'd39164, 16'd6911, 16'd16941, 16'd6379, 16'd38060, 16'd21761, 16'd26551, 16'd41821, 16'd55273, 16'd58674, 16'd34387, 16'd54917, 16'd20431, 16'd27307, 16'd55823, 16'd11294, 16'd22845, 16'd36500, 16'd58770, 16'd3902, 16'd38309, 16'd92, 16'd5346, 16'd49655, 16'd60547});
	test_expansion(128'h9a66a50c60290cc0f177a045e2b69c33, {16'd16700, 16'd21460, 16'd53025, 16'd16923, 16'd30136, 16'd39535, 16'd43448, 16'd20028, 16'd2542, 16'd62857, 16'd51540, 16'd8106, 16'd43841, 16'd39603, 16'd23647, 16'd33688, 16'd32759, 16'd34947, 16'd18222, 16'd21740, 16'd59659, 16'd10366, 16'd60342, 16'd39119, 16'd59620, 16'd4135});
	test_expansion(128'h1230790e580532b88c62a5a155df694d, {16'd41375, 16'd50901, 16'd16245, 16'd8455, 16'd17109, 16'd62876, 16'd5930, 16'd47671, 16'd52720, 16'd40785, 16'd37397, 16'd36924, 16'd5587, 16'd38049, 16'd40206, 16'd62451, 16'd4046, 16'd3583, 16'd17068, 16'd32700, 16'd49240, 16'd13752, 16'd46180, 16'd53065, 16'd54210, 16'd14342});
	test_expansion(128'h2931be22822a959c130290869557a1f4, {16'd23966, 16'd36147, 16'd25299, 16'd45572, 16'd41500, 16'd34872, 16'd20482, 16'd44141, 16'd5581, 16'd35479, 16'd37798, 16'd36338, 16'd6478, 16'd27424, 16'd28078, 16'd19220, 16'd42174, 16'd1028, 16'd18278, 16'd21395, 16'd55057, 16'd35737, 16'd26037, 16'd37181, 16'd24514, 16'd27072});
	test_expansion(128'hbb47f1562ad5045eb4942121cc414fdb, {16'd28286, 16'd27851, 16'd5859, 16'd56298, 16'd50909, 16'd61616, 16'd24152, 16'd40689, 16'd2177, 16'd21678, 16'd20358, 16'd27197, 16'd54284, 16'd376, 16'd51377, 16'd63715, 16'd55370, 16'd9726, 16'd10284, 16'd65284, 16'd5992, 16'd28584, 16'd61351, 16'd42699, 16'd49978, 16'd35820});
	test_expansion(128'h260a310e52a8d379112058b0c45fec10, {16'd38115, 16'd65164, 16'd38841, 16'd4034, 16'd47830, 16'd38513, 16'd3546, 16'd62375, 16'd12951, 16'd52410, 16'd22978, 16'd45281, 16'd14546, 16'd21542, 16'd21594, 16'd59673, 16'd34363, 16'd29473, 16'd9103, 16'd62341, 16'd41391, 16'd41282, 16'd32780, 16'd50775, 16'd19100, 16'd38399});
	test_expansion(128'ha2d1167c7bd7ea113ab259da01aad85c, {16'd63703, 16'd20722, 16'd2707, 16'd21431, 16'd11880, 16'd64234, 16'd37497, 16'd2156, 16'd12954, 16'd29008, 16'd14114, 16'd41778, 16'd26301, 16'd1514, 16'd2935, 16'd22957, 16'd63016, 16'd6959, 16'd61010, 16'd11854, 16'd65327, 16'd49583, 16'd14416, 16'd21096, 16'd56204, 16'd23215});
	test_expansion(128'hf19a803a26b156030b9eb4e0e103d4ad, {16'd62013, 16'd34081, 16'd26295, 16'd20488, 16'd14155, 16'd32262, 16'd52386, 16'd34523, 16'd24291, 16'd58598, 16'd20493, 16'd28469, 16'd46200, 16'd9107, 16'd53906, 16'd38841, 16'd35767, 16'd52418, 16'd36179, 16'd19679, 16'd27425, 16'd3452, 16'd30799, 16'd41181, 16'd5345, 16'd56839});
	test_expansion(128'h73e39caf7989ec8e0b23e3cbb5739ce2, {16'd15365, 16'd43991, 16'd52541, 16'd1441, 16'd8797, 16'd41767, 16'd28857, 16'd11053, 16'd6706, 16'd20386, 16'd40478, 16'd36966, 16'd50941, 16'd44847, 16'd37617, 16'd11570, 16'd4683, 16'd32208, 16'd64432, 16'd57345, 16'd55919, 16'd38989, 16'd60369, 16'd45989, 16'd56407, 16'd42646});
	test_expansion(128'h6f84b95847e2f678ca2a7952b29f11d1, {16'd787, 16'd57117, 16'd27422, 16'd61307, 16'd23888, 16'd39662, 16'd20846, 16'd38251, 16'd46881, 16'd12918, 16'd53772, 16'd54366, 16'd63357, 16'd8, 16'd48328, 16'd38757, 16'd8023, 16'd3253, 16'd58376, 16'd53655, 16'd17320, 16'd25580, 16'd55672, 16'd51909, 16'd63058, 16'd58292});
	test_expansion(128'h53c4aff8fd5123e62eed78cb02d7e156, {16'd8985, 16'd26964, 16'd28343, 16'd21678, 16'd27571, 16'd18339, 16'd54411, 16'd1616, 16'd11936, 16'd43390, 16'd4848, 16'd25678, 16'd20635, 16'd37535, 16'd43479, 16'd59527, 16'd59173, 16'd26148, 16'd36927, 16'd41280, 16'd39757, 16'd63643, 16'd24858, 16'd25427, 16'd15197, 16'd29728});
	test_expansion(128'hbb42c1a1bdad4ae7657f65e30af755ea, {16'd61262, 16'd19663, 16'd59963, 16'd55557, 16'd37461, 16'd36676, 16'd57226, 16'd43943, 16'd6710, 16'd19306, 16'd49701, 16'd50693, 16'd40254, 16'd46608, 16'd45359, 16'd16378, 16'd64748, 16'd41778, 16'd22282, 16'd59373, 16'd2401, 16'd9838, 16'd28753, 16'd55364, 16'd15237, 16'd59523});
	test_expansion(128'h734f0eb6bc1cbb58eb9a82e3bf2ddc06, {16'd18990, 16'd38506, 16'd57299, 16'd24998, 16'd48608, 16'd4203, 16'd60297, 16'd35222, 16'd13697, 16'd26081, 16'd36640, 16'd12377, 16'd63995, 16'd50406, 16'd59592, 16'd28767, 16'd26600, 16'd54883, 16'd17076, 16'd14612, 16'd36392, 16'd12393, 16'd35514, 16'd33135, 16'd19438, 16'd48741});
	test_expansion(128'h4a994ee90039e29153e610f5a229c239, {16'd52139, 16'd9668, 16'd23931, 16'd5653, 16'd56369, 16'd24846, 16'd41558, 16'd63586, 16'd51724, 16'd8286, 16'd54467, 16'd27181, 16'd45199, 16'd22446, 16'd34156, 16'd17239, 16'd22595, 16'd50095, 16'd11528, 16'd12454, 16'd62067, 16'd3405, 16'd33398, 16'd55965, 16'd33773, 16'd43902});
	test_expansion(128'h827a8f92598f57ece6ee49da3e691bd3, {16'd38393, 16'd4868, 16'd49646, 16'd42262, 16'd19177, 16'd26750, 16'd12014, 16'd310, 16'd32084, 16'd58969, 16'd20789, 16'd63200, 16'd52117, 16'd32655, 16'd56673, 16'd59463, 16'd10161, 16'd21213, 16'd10525, 16'd36928, 16'd19556, 16'd63054, 16'd2227, 16'd59496, 16'd10683, 16'd18278});
	test_expansion(128'hcffc1c1f762ed54670d82b081282f1ab, {16'd62361, 16'd56096, 16'd5040, 16'd35351, 16'd18530, 16'd43674, 16'd8357, 16'd54757, 16'd1641, 16'd54081, 16'd10839, 16'd4903, 16'd14079, 16'd55858, 16'd59855, 16'd30067, 16'd35170, 16'd60064, 16'd38306, 16'd58755, 16'd25310, 16'd12005, 16'd44402, 16'd41067, 16'd46100, 16'd7967});
	test_expansion(128'h69745d1fdc74b83f3f2ad81e10a52580, {16'd56366, 16'd62210, 16'd28651, 16'd53366, 16'd44810, 16'd35305, 16'd27688, 16'd27332, 16'd51190, 16'd41087, 16'd9186, 16'd50465, 16'd62628, 16'd40407, 16'd25592, 16'd34233, 16'd45222, 16'd12097, 16'd1489, 16'd28107, 16'd14387, 16'd20460, 16'd24787, 16'd47224, 16'd5659, 16'd35977});
	test_expansion(128'h522babf36e6c12c1961d919821c532e7, {16'd54107, 16'd17003, 16'd35354, 16'd21724, 16'd47501, 16'd5559, 16'd8022, 16'd55644, 16'd29698, 16'd58331, 16'd22793, 16'd89, 16'd32595, 16'd33976, 16'd49591, 16'd57591, 16'd25796, 16'd29527, 16'd18111, 16'd29616, 16'd39592, 16'd17342, 16'd15624, 16'd56447, 16'd3906, 16'd30316});
	test_expansion(128'h98f2cd5b70db3f3f252e12171ee2dab3, {16'd62137, 16'd46111, 16'd41207, 16'd35182, 16'd12326, 16'd59101, 16'd45715, 16'd32099, 16'd5237, 16'd47416, 16'd40195, 16'd32507, 16'd58893, 16'd37762, 16'd41830, 16'd29939, 16'd31439, 16'd23100, 16'd27612, 16'd4520, 16'd51118, 16'd15619, 16'd55075, 16'd10969, 16'd2503, 16'd60573});
	test_expansion(128'h7d50b171578ebe068e31cf9f71127b19, {16'd53299, 16'd30748, 16'd57331, 16'd44537, 16'd3992, 16'd13897, 16'd20322, 16'd59404, 16'd56626, 16'd33634, 16'd3015, 16'd26397, 16'd22190, 16'd32180, 16'd30767, 16'd17961, 16'd5170, 16'd24344, 16'd42634, 16'd2795, 16'd10513, 16'd27303, 16'd53558, 16'd59621, 16'd51787, 16'd50729});
	test_expansion(128'h60a027d49415fa53037d3c307c1c369a, {16'd10146, 16'd43474, 16'd28766, 16'd22396, 16'd2178, 16'd63248, 16'd15738, 16'd52583, 16'd11206, 16'd3406, 16'd61774, 16'd27769, 16'd59075, 16'd3849, 16'd36302, 16'd452, 16'd53159, 16'd46232, 16'd1319, 16'd14572, 16'd18559, 16'd44399, 16'd51567, 16'd61606, 16'd26887, 16'd65310});
	test_expansion(128'h2dffd108f183f7717797862deef0c8f6, {16'd16485, 16'd37227, 16'd7892, 16'd64815, 16'd5830, 16'd25081, 16'd42999, 16'd63561, 16'd38385, 16'd31399, 16'd24356, 16'd53584, 16'd3753, 16'd52794, 16'd39865, 16'd65350, 16'd39391, 16'd37683, 16'd44849, 16'd64829, 16'd9801, 16'd6500, 16'd9914, 16'd56045, 16'd18467, 16'd46183});
	test_expansion(128'hcbb4e10b88db538f745a821b275262b1, {16'd61198, 16'd59674, 16'd5707, 16'd20486, 16'd41109, 16'd18314, 16'd3123, 16'd63385, 16'd38645, 16'd22995, 16'd48228, 16'd6758, 16'd45893, 16'd10796, 16'd55861, 16'd10260, 16'd13991, 16'd54915, 16'd56711, 16'd63863, 16'd38783, 16'd29503, 16'd51797, 16'd1694, 16'd20962, 16'd44569});
	test_expansion(128'hbc0c845852812796defeee2a54b047c2, {16'd27812, 16'd19947, 16'd4979, 16'd32865, 16'd43775, 16'd32395, 16'd2480, 16'd11452, 16'd43824, 16'd334, 16'd5827, 16'd15509, 16'd15258, 16'd1728, 16'd36946, 16'd8016, 16'd11589, 16'd7501, 16'd60338, 16'd9638, 16'd59847, 16'd58813, 16'd38280, 16'd21007, 16'd46792, 16'd24326});
	test_expansion(128'h5c2c18a3ced15140b49638febdd2f391, {16'd2484, 16'd33255, 16'd52766, 16'd16437, 16'd6035, 16'd52015, 16'd64313, 16'd29319, 16'd20642, 16'd10265, 16'd19891, 16'd56328, 16'd11465, 16'd57939, 16'd36333, 16'd54825, 16'd4545, 16'd40355, 16'd38853, 16'd13924, 16'd50333, 16'd63428, 16'd58632, 16'd10801, 16'd64647, 16'd37111});
	test_expansion(128'he7fe9b8b6c6befcb223442851430d7a7, {16'd58208, 16'd48956, 16'd6711, 16'd33142, 16'd25242, 16'd64311, 16'd46006, 16'd50359, 16'd51585, 16'd47386, 16'd30446, 16'd41209, 16'd57429, 16'd10269, 16'd917, 16'd17728, 16'd52396, 16'd38996, 16'd65523, 16'd61745, 16'd53693, 16'd56370, 16'd11826, 16'd63022, 16'd47208, 16'd30517});
	test_expansion(128'ha6201ac117bb3fb8684160756dece35e, {16'd32534, 16'd17333, 16'd38516, 16'd11488, 16'd43720, 16'd59990, 16'd41587, 16'd42014, 16'd60634, 16'd8184, 16'd60632, 16'd29111, 16'd12189, 16'd26040, 16'd61562, 16'd56017, 16'd33457, 16'd19669, 16'd21678, 16'd40309, 16'd15787, 16'd268, 16'd57145, 16'd47559, 16'd26791, 16'd763});
	test_expansion(128'h7229e64a848222bd1c004751c9be0301, {16'd16183, 16'd40439, 16'd5566, 16'd11697, 16'd64865, 16'd46654, 16'd47676, 16'd53127, 16'd28319, 16'd33268, 16'd43459, 16'd42409, 16'd27517, 16'd29462, 16'd37564, 16'd18776, 16'd25978, 16'd57131, 16'd9387, 16'd19186, 16'd35834, 16'd30007, 16'd20721, 16'd19503, 16'd25068, 16'd5394});
	test_expansion(128'h412efbc676131ba8ab35b8fc5461cf58, {16'd9395, 16'd24372, 16'd26347, 16'd53237, 16'd23524, 16'd52826, 16'd19691, 16'd35290, 16'd11133, 16'd52263, 16'd26665, 16'd5650, 16'd30096, 16'd19694, 16'd10405, 16'd41885, 16'd19872, 16'd8865, 16'd5302, 16'd7170, 16'd3343, 16'd16592, 16'd34518, 16'd44181, 16'd25015, 16'd29649});
	test_expansion(128'h13ebfa06b0e5e27fec4685f3d57f0800, {16'd29303, 16'd32078, 16'd8754, 16'd3298, 16'd54371, 16'd6890, 16'd13665, 16'd54341, 16'd10196, 16'd38958, 16'd46434, 16'd2871, 16'd29859, 16'd8019, 16'd38535, 16'd287, 16'd43899, 16'd51681, 16'd6269, 16'd51394, 16'd24620, 16'd22632, 16'd34603, 16'd53791, 16'd7663, 16'd48542});
	test_expansion(128'hb5abad5b7aeb7d114a37e179e77e24a2, {16'd56572, 16'd29353, 16'd36773, 16'd48095, 16'd59968, 16'd43309, 16'd1767, 16'd48513, 16'd62918, 16'd33489, 16'd46807, 16'd58400, 16'd44011, 16'd51860, 16'd20198, 16'd59833, 16'd15345, 16'd25901, 16'd42917, 16'd47146, 16'd43902, 16'd27110, 16'd22504, 16'd21055, 16'd18430, 16'd6988});
	test_expansion(128'h84acdd071e9b0629dd718d3754e973f0, {16'd14447, 16'd45205, 16'd4277, 16'd28598, 16'd42709, 16'd5201, 16'd22768, 16'd59667, 16'd12651, 16'd1305, 16'd45136, 16'd8405, 16'd35489, 16'd59145, 16'd62867, 16'd35029, 16'd52772, 16'd32459, 16'd2791, 16'd121, 16'd3123, 16'd14168, 16'd37199, 16'd55368, 16'd18830, 16'd45404});
	test_expansion(128'h6799c723fcdc27285f544397809e4a63, {16'd30476, 16'd27575, 16'd18370, 16'd51372, 16'd27257, 16'd4052, 16'd51208, 16'd36303, 16'd32107, 16'd63410, 16'd50592, 16'd47984, 16'd46519, 16'd34178, 16'd57209, 16'd58374, 16'd29187, 16'd47698, 16'd55624, 16'd21749, 16'd42464, 16'd45747, 16'd3112, 16'd21602, 16'd54162, 16'd17327});
	test_expansion(128'hfea6091c4cc44bf2426edcfdce1f06eb, {16'd52343, 16'd22648, 16'd8225, 16'd38958, 16'd56129, 16'd42510, 16'd14130, 16'd38335, 16'd41925, 16'd38927, 16'd13929, 16'd44949, 16'd31237, 16'd3452, 16'd24311, 16'd14305, 16'd43400, 16'd30657, 16'd22606, 16'd19383, 16'd35, 16'd13603, 16'd42810, 16'd54979, 16'd47944, 16'd40872});
	test_expansion(128'h16d46492063ae2c0f6a891c1b7940e54, {16'd41705, 16'd6334, 16'd12342, 16'd35838, 16'd38292, 16'd47155, 16'd40449, 16'd64205, 16'd5542, 16'd28846, 16'd8706, 16'd18981, 16'd26103, 16'd14755, 16'd4425, 16'd17107, 16'd56109, 16'd10351, 16'd59052, 16'd55782, 16'd7698, 16'd45343, 16'd16574, 16'd8016, 16'd7175, 16'd56749});
	test_expansion(128'h3797f067dd624888a3c16b48906c8620, {16'd50579, 16'd26796, 16'd49466, 16'd13499, 16'd56377, 16'd1124, 16'd163, 16'd7267, 16'd34931, 16'd28314, 16'd59790, 16'd698, 16'd629, 16'd34324, 16'd32311, 16'd49685, 16'd58250, 16'd27995, 16'd5219, 16'd28668, 16'd50650, 16'd20376, 16'd33578, 16'd2740, 16'd26134, 16'd26645});
	test_expansion(128'hfc776500bef55f88acb8795558d5c3a3, {16'd2318, 16'd20728, 16'd57883, 16'd40538, 16'd26867, 16'd36800, 16'd30360, 16'd46176, 16'd4604, 16'd54545, 16'd32124, 16'd58062, 16'd36293, 16'd44429, 16'd7194, 16'd42709, 16'd6975, 16'd40770, 16'd35889, 16'd2310, 16'd22464, 16'd23355, 16'd22831, 16'd1645, 16'd16852, 16'd5325});
	test_expansion(128'hf082ee778fdf56d0639f582b7d37dc0c, {16'd53943, 16'd32342, 16'd2324, 16'd11359, 16'd28099, 16'd32956, 16'd47723, 16'd54808, 16'd8478, 16'd50993, 16'd39133, 16'd8622, 16'd15233, 16'd5762, 16'd16357, 16'd7036, 16'd51934, 16'd13227, 16'd50390, 16'd46933, 16'd65114, 16'd62906, 16'd40197, 16'd51948, 16'd36831, 16'd39536});
	test_expansion(128'h778d316ad50376550c1a997d0f711025, {16'd56633, 16'd62560, 16'd23162, 16'd26714, 16'd60159, 16'd39936, 16'd1814, 16'd60398, 16'd24808, 16'd59092, 16'd53019, 16'd35664, 16'd18961, 16'd35779, 16'd20027, 16'd18019, 16'd56761, 16'd15866, 16'd42856, 16'd11095, 16'd59929, 16'd39679, 16'd10953, 16'd970, 16'd34702, 16'd33379});
	test_expansion(128'h89b7d7f17d3df3667d556c6152ce0615, {16'd53340, 16'd154, 16'd4570, 16'd53057, 16'd25781, 16'd65407, 16'd7491, 16'd48630, 16'd60149, 16'd39105, 16'd62405, 16'd64810, 16'd17577, 16'd47680, 16'd15996, 16'd46843, 16'd45515, 16'd11994, 16'd38701, 16'd41685, 16'd17022, 16'd57611, 16'd54166, 16'd6394, 16'd65143, 16'd37216});
	test_expansion(128'h643fcace9c1f75b2a3fa6ce370679d33, {16'd56587, 16'd61148, 16'd64324, 16'd1312, 16'd8090, 16'd13846, 16'd19241, 16'd48527, 16'd19255, 16'd12178, 16'd17697, 16'd58379, 16'd17845, 16'd18403, 16'd40261, 16'd46422, 16'd39448, 16'd65307, 16'd23822, 16'd47683, 16'd18132, 16'd36237, 16'd64587, 16'd3183, 16'd11379, 16'd15713});
	test_expansion(128'hde1193347a3d910ae2ecd0a4d6097a42, {16'd8978, 16'd44602, 16'd63271, 16'd38280, 16'd2232, 16'd10591, 16'd11951, 16'd20107, 16'd12734, 16'd37559, 16'd15178, 16'd8357, 16'd17871, 16'd24040, 16'd4672, 16'd6693, 16'd23363, 16'd47028, 16'd28643, 16'd41350, 16'd45674, 16'd40796, 16'd64764, 16'd11684, 16'd5663, 16'd52297});
	test_expansion(128'h51135e23589438f0454dc6687996eca4, {16'd46155, 16'd54811, 16'd53992, 16'd5106, 16'd1370, 16'd19197, 16'd33806, 16'd62348, 16'd14248, 16'd28914, 16'd32053, 16'd2953, 16'd48934, 16'd131, 16'd21890, 16'd47460, 16'd16896, 16'd24082, 16'd2355, 16'd23607, 16'd38696, 16'd22866, 16'd17975, 16'd11164, 16'd47278, 16'd13299});
	test_expansion(128'h5987021c3ea61defd8d4bded4cb78786, {16'd32250, 16'd28935, 16'd32546, 16'd36621, 16'd55775, 16'd63909, 16'd14143, 16'd53351, 16'd30549, 16'd6778, 16'd32550, 16'd48204, 16'd61925, 16'd55271, 16'd31083, 16'd42949, 16'd9039, 16'd49890, 16'd61487, 16'd9232, 16'd23464, 16'd48492, 16'd20229, 16'd47793, 16'd61402, 16'd15433});
	test_expansion(128'hefa1f1ea96245eaab12e93fea19e80e6, {16'd20799, 16'd10638, 16'd50557, 16'd59640, 16'd13036, 16'd50355, 16'd52335, 16'd4104, 16'd22997, 16'd21378, 16'd31432, 16'd19532, 16'd14808, 16'd4133, 16'd49228, 16'd28244, 16'd57737, 16'd26961, 16'd5983, 16'd9457, 16'd59134, 16'd36699, 16'd3108, 16'd50240, 16'd36776, 16'd12464});
	test_expansion(128'hf2890a2b2cf29b8c9bd4edcb21cdb9af, {16'd16989, 16'd16042, 16'd47542, 16'd64292, 16'd35982, 16'd24452, 16'd4934, 16'd28684, 16'd7895, 16'd21578, 16'd19261, 16'd36330, 16'd64341, 16'd12095, 16'd12791, 16'd27856, 16'd12800, 16'd32922, 16'd52809, 16'd61854, 16'd54263, 16'd57224, 16'd19427, 16'd8105, 16'd40708, 16'd9277});
	test_expansion(128'h922ea1dfef0b70369fff50b69de5066d, {16'd45781, 16'd15783, 16'd11740, 16'd55433, 16'd30171, 16'd48649, 16'd44789, 16'd30011, 16'd5930, 16'd64309, 16'd39285, 16'd46733, 16'd2979, 16'd8653, 16'd2098, 16'd44631, 16'd1928, 16'd12174, 16'd54579, 16'd16417, 16'd14392, 16'd3285, 16'd28336, 16'd19885, 16'd15934, 16'd42958});
	test_expansion(128'h21d9f9873df64166222d001d575714b7, {16'd22124, 16'd21751, 16'd59382, 16'd18971, 16'd7275, 16'd53751, 16'd23196, 16'd14483, 16'd41216, 16'd59828, 16'd49383, 16'd48829, 16'd59596, 16'd61309, 16'd47512, 16'd14040, 16'd30358, 16'd2216, 16'd55302, 16'd36216, 16'd30604, 16'd55653, 16'd64686, 16'd2352, 16'd52637, 16'd28664});
	test_expansion(128'h3e3f799228f31ce5119935aeb1dc9374, {16'd64241, 16'd64650, 16'd14387, 16'd40420, 16'd15507, 16'd52732, 16'd18238, 16'd49188, 16'd53312, 16'd34046, 16'd59730, 16'd41802, 16'd65301, 16'd37678, 16'd14884, 16'd28641, 16'd38856, 16'd45848, 16'd24717, 16'd37368, 16'd26737, 16'd43376, 16'd48900, 16'd35282, 16'd27611, 16'd63640});
	test_expansion(128'ha6daea0961a8e01195ec55bd0a504c7d, {16'd63271, 16'd49996, 16'd6067, 16'd26004, 16'd23915, 16'd42844, 16'd4933, 16'd60928, 16'd58943, 16'd52729, 16'd37015, 16'd21943, 16'd28387, 16'd15708, 16'd19682, 16'd64325, 16'd3788, 16'd16088, 16'd27936, 16'd13635, 16'd22634, 16'd52323, 16'd49989, 16'd63945, 16'd11069, 16'd49875});
	test_expansion(128'h055e3f425e9604854533048970abb2fb, {16'd9353, 16'd25883, 16'd25693, 16'd32777, 16'd30963, 16'd11848, 16'd11675, 16'd2658, 16'd10482, 16'd22947, 16'd21306, 16'd40777, 16'd22001, 16'd17859, 16'd8936, 16'd36789, 16'd8116, 16'd65012, 16'd15816, 16'd50968, 16'd54341, 16'd31461, 16'd3051, 16'd12499, 16'd64483, 16'd48736});
	test_expansion(128'hb41073a252dea57d062b349a3af728b6, {16'd30123, 16'd64444, 16'd2002, 16'd28481, 16'd55848, 16'd56714, 16'd28998, 16'd43285, 16'd47886, 16'd13358, 16'd48158, 16'd34847, 16'd62163, 16'd14034, 16'd58636, 16'd59926, 16'd6273, 16'd58924, 16'd23733, 16'd2701, 16'd45242, 16'd23789, 16'd29624, 16'd21259, 16'd65346, 16'd54223});
	test_expansion(128'had6e9b544f8695e18f87dc7ea766f345, {16'd57208, 16'd61519, 16'd6495, 16'd55568, 16'd33080, 16'd2622, 16'd60915, 16'd31871, 16'd16000, 16'd52934, 16'd58587, 16'd31273, 16'd30943, 16'd13078, 16'd22814, 16'd40337, 16'd6879, 16'd54791, 16'd59619, 16'd4697, 16'd64526, 16'd52732, 16'd24928, 16'd957, 16'd155, 16'd41186});
	test_expansion(128'h7c6463a0bfd97d4d9d40adf1cc69a34c, {16'd30555, 16'd7008, 16'd24182, 16'd41808, 16'd53802, 16'd8908, 16'd1397, 16'd16277, 16'd58239, 16'd13338, 16'd31425, 16'd36423, 16'd19698, 16'd29160, 16'd19914, 16'd25997, 16'd24082, 16'd10970, 16'd25356, 16'd56356, 16'd44403, 16'd34703, 16'd7226, 16'd2425, 16'd25598, 16'd28426});
	test_expansion(128'hd28cc4308143f8822d5f064cf767683f, {16'd4250, 16'd29916, 16'd24163, 16'd43582, 16'd20872, 16'd20797, 16'd3571, 16'd16707, 16'd568, 16'd41659, 16'd62148, 16'd8845, 16'd16535, 16'd16734, 16'd44041, 16'd13841, 16'd60530, 16'd64361, 16'd33203, 16'd28897, 16'd38532, 16'd24966, 16'd19299, 16'd3919, 16'd13088, 16'd10489});
	test_expansion(128'hedb1166ea78f21f68f8dfb2c10ec4901, {16'd52430, 16'd47631, 16'd29898, 16'd10856, 16'd12847, 16'd45942, 16'd28088, 16'd53672, 16'd60297, 16'd40213, 16'd36537, 16'd35715, 16'd35921, 16'd55433, 16'd18866, 16'd58434, 16'd1082, 16'd10137, 16'd41196, 16'd10993, 16'd18633, 16'd42869, 16'd23048, 16'd57486, 16'd44476, 16'd29031});
	test_expansion(128'h0f0e1ff882ce0aef87db80fc5eb5f000, {16'd39623, 16'd58404, 16'd56366, 16'd54590, 16'd25584, 16'd57594, 16'd37188, 16'd49928, 16'd20291, 16'd30128, 16'd18072, 16'd52479, 16'd31063, 16'd12326, 16'd13476, 16'd47393, 16'd6212, 16'd46478, 16'd2265, 16'd20001, 16'd60798, 16'd25800, 16'd59891, 16'd10209, 16'd22508, 16'd33001});
	test_expansion(128'hb13d68e5f8a832da60ea466e5721f270, {16'd2895, 16'd42409, 16'd605, 16'd58509, 16'd45374, 16'd28564, 16'd3821, 16'd2705, 16'd22560, 16'd4357, 16'd61381, 16'd61978, 16'd12130, 16'd37176, 16'd15202, 16'd3645, 16'd60185, 16'd64371, 16'd8917, 16'd37107, 16'd48486, 16'd49248, 16'd64130, 16'd47851, 16'd46044, 16'd57278});
	test_expansion(128'hd3e8441520ce96880181da8843174f7f, {16'd57374, 16'd57503, 16'd55109, 16'd48466, 16'd49246, 16'd61542, 16'd35050, 16'd7629, 16'd4905, 16'd8971, 16'd5057, 16'd25305, 16'd59975, 16'd3299, 16'd51548, 16'd10640, 16'd18157, 16'd52434, 16'd35859, 16'd41334, 16'd65258, 16'd747, 16'd54182, 16'd55841, 16'd1464, 16'd45975});
	test_expansion(128'hd777ed9e0c332075f573e67d42be4138, {16'd65286, 16'd37556, 16'd56270, 16'd26050, 16'd20418, 16'd21116, 16'd18910, 16'd46553, 16'd49767, 16'd756, 16'd30027, 16'd59186, 16'd9077, 16'd46476, 16'd37929, 16'd20263, 16'd42329, 16'd56310, 16'd7099, 16'd29730, 16'd22009, 16'd5070, 16'd18368, 16'd50765, 16'd56620, 16'd36859});
	test_expansion(128'h1c16b2f04c5e0315299c9d6f8a5cb034, {16'd8101, 16'd33289, 16'd46692, 16'd19660, 16'd26501, 16'd63060, 16'd61623, 16'd25808, 16'd64923, 16'd16776, 16'd41954, 16'd26470, 16'd40026, 16'd53533, 16'd6768, 16'd43120, 16'd14921, 16'd5482, 16'd21456, 16'd53922, 16'd43703, 16'd36363, 16'd32686, 16'd7465, 16'd57019, 16'd48919});
	test_expansion(128'hbd028b0c5a6814ce46a5008a9f24f9b4, {16'd27208, 16'd14917, 16'd41284, 16'd15679, 16'd51822, 16'd20198, 16'd18822, 16'd18120, 16'd48527, 16'd63905, 16'd20361, 16'd1550, 16'd54176, 16'd52852, 16'd21425, 16'd7790, 16'd7670, 16'd30701, 16'd34551, 16'd9837, 16'd7013, 16'd22605, 16'd29096, 16'd42720, 16'd61273, 16'd65133});
	test_expansion(128'h120ee7d06b6751327f2fdd775228d2e2, {16'd60021, 16'd8694, 16'd51493, 16'd29267, 16'd6988, 16'd37340, 16'd9006, 16'd6202, 16'd19511, 16'd53429, 16'd50877, 16'd18558, 16'd42548, 16'd49403, 16'd7924, 16'd37098, 16'd31896, 16'd12924, 16'd42887, 16'd7624, 16'd8763, 16'd54202, 16'd4481, 16'd36660, 16'd33389, 16'd59597});
	test_expansion(128'h9cb732d9ed00b181135c0cc0b74aa181, {16'd14433, 16'd3583, 16'd38202, 16'd61256, 16'd27505, 16'd15052, 16'd54484, 16'd43324, 16'd7869, 16'd27032, 16'd49718, 16'd55235, 16'd30138, 16'd814, 16'd63002, 16'd27293, 16'd58323, 16'd19375, 16'd40445, 16'd2471, 16'd51840, 16'd26294, 16'd55977, 16'd42110, 16'd9659, 16'd60727});
	test_expansion(128'h9fad3bf488d3cc1e195386416699ab1b, {16'd60440, 16'd17808, 16'd7920, 16'd15554, 16'd39131, 16'd42098, 16'd34950, 16'd33166, 16'd26761, 16'd49949, 16'd11206, 16'd47904, 16'd59331, 16'd28013, 16'd63473, 16'd56501, 16'd35462, 16'd25941, 16'd12453, 16'd34217, 16'd54599, 16'd36559, 16'd60871, 16'd50647, 16'd35172, 16'd51273});
	test_expansion(128'h2d68758dddf13168f64877f4976c3578, {16'd19416, 16'd251, 16'd55716, 16'd54750, 16'd27170, 16'd2063, 16'd22131, 16'd8362, 16'd16421, 16'd29868, 16'd3339, 16'd7905, 16'd20747, 16'd61284, 16'd20841, 16'd13008, 16'd665, 16'd35185, 16'd57718, 16'd41813, 16'd31102, 16'd10815, 16'd22877, 16'd6266, 16'd21127, 16'd27198});
	test_expansion(128'hef5383fd0fc35a5dcb1acb2e3e461412, {16'd48505, 16'd1888, 16'd43146, 16'd17431, 16'd29294, 16'd15907, 16'd30814, 16'd33105, 16'd39963, 16'd40989, 16'd51297, 16'd25280, 16'd34057, 16'd18875, 16'd35892, 16'd12293, 16'd48648, 16'd44325, 16'd18210, 16'd9287, 16'd27517, 16'd8207, 16'd8673, 16'd65412, 16'd63274, 16'd29});
	test_expansion(128'h801d11611daf766006c5925530d200e5, {16'd61865, 16'd47844, 16'd6751, 16'd24586, 16'd16355, 16'd3331, 16'd63233, 16'd10037, 16'd22731, 16'd29148, 16'd24801, 16'd23395, 16'd44681, 16'd29711, 16'd53194, 16'd54640, 16'd50250, 16'd31056, 16'd56705, 16'd57460, 16'd46221, 16'd18172, 16'd48745, 16'd4287, 16'd14568, 16'd56207});
	test_expansion(128'hab15bd0e6b090a19b90a1d7c6c2757cc, {16'd34571, 16'd35318, 16'd32105, 16'd14670, 16'd31551, 16'd27862, 16'd56619, 16'd15954, 16'd5128, 16'd27463, 16'd60867, 16'd504, 16'd63567, 16'd26358, 16'd21569, 16'd34461, 16'd64152, 16'd30078, 16'd55712, 16'd36371, 16'd5432, 16'd50258, 16'd22507, 16'd60599, 16'd47933, 16'd53300});
	test_expansion(128'h8f34be7df91ecd293a52f9e384630f62, {16'd34387, 16'd33675, 16'd26141, 16'd20829, 16'd62007, 16'd59518, 16'd11765, 16'd64508, 16'd50945, 16'd11477, 16'd19898, 16'd48659, 16'd41913, 16'd23388, 16'd3417, 16'd27975, 16'd44362, 16'd61975, 16'd5411, 16'd23749, 16'd23979, 16'd15496, 16'd32706, 16'd22530, 16'd29627, 16'd63158});
	test_expansion(128'h41dc955ba75628abb1fe964672895ede, {16'd44383, 16'd24572, 16'd14345, 16'd64423, 16'd14012, 16'd31432, 16'd55748, 16'd57078, 16'd17483, 16'd35900, 16'd60006, 16'd63020, 16'd40002, 16'd17461, 16'd20915, 16'd62551, 16'd10978, 16'd40058, 16'd50415, 16'd1895, 16'd65231, 16'd51194, 16'd46341, 16'd14456, 16'd45080, 16'd10377});
	test_expansion(128'h15c6276e1a23f2883bef739ba5b610cb, {16'd55545, 16'd61516, 16'd59498, 16'd30901, 16'd3031, 16'd48550, 16'd26674, 16'd13200, 16'd46738, 16'd37892, 16'd4644, 16'd11103, 16'd18940, 16'd15791, 16'd25291, 16'd35278, 16'd35044, 16'd60672, 16'd17896, 16'd42119, 16'd63745, 16'd33741, 16'd57891, 16'd40991, 16'd63319, 16'd52001});
	test_expansion(128'he2a1954e030dd23564dd16ed563bfc70, {16'd41672, 16'd3806, 16'd20234, 16'd6265, 16'd53118, 16'd2031, 16'd46610, 16'd34121, 16'd40306, 16'd36340, 16'd62470, 16'd472, 16'd41330, 16'd49384, 16'd45505, 16'd54873, 16'd8443, 16'd19953, 16'd30901, 16'd8443, 16'd61261, 16'd18111, 16'd52266, 16'd13053, 16'd47512, 16'd45667});
	test_expansion(128'h559b57f9043d009bfb82e74185fc2780, {16'd29718, 16'd48441, 16'd39947, 16'd64881, 16'd34817, 16'd51846, 16'd45611, 16'd53330, 16'd31878, 16'd58680, 16'd60728, 16'd63800, 16'd27148, 16'd1096, 16'd4273, 16'd46678, 16'd40047, 16'd5572, 16'd3026, 16'd19373, 16'd34813, 16'd25479, 16'd8180, 16'd53298, 16'd14815, 16'd40960});
	test_expansion(128'h3050dfa8ddb1d47b5207f81c4e3d24db, {16'd12650, 16'd10330, 16'd19773, 16'd3091, 16'd49521, 16'd58941, 16'd28128, 16'd8039, 16'd36865, 16'd63384, 16'd60290, 16'd26561, 16'd8294, 16'd7754, 16'd21098, 16'd16765, 16'd19305, 16'd3906, 16'd26308, 16'd34825, 16'd54631, 16'd53867, 16'd10722, 16'd43601, 16'd14601, 16'd43832});
	test_expansion(128'he9cadda45f227fdb83294e01a6d886c4, {16'd47092, 16'd35709, 16'd37462, 16'd61403, 16'd10626, 16'd37061, 16'd43340, 16'd64596, 16'd60666, 16'd59144, 16'd53390, 16'd17318, 16'd53685, 16'd60391, 16'd33944, 16'd41677, 16'd3414, 16'd38676, 16'd59980, 16'd8569, 16'd57512, 16'd16740, 16'd38333, 16'd15849, 16'd53515, 16'd38211});
	test_expansion(128'h582f9c138681f5dcc1ad25796137579b, {16'd58482, 16'd17055, 16'd21388, 16'd46670, 16'd59106, 16'd28839, 16'd13715, 16'd12, 16'd51823, 16'd38279, 16'd21374, 16'd58607, 16'd27394, 16'd60435, 16'd26579, 16'd45374, 16'd50720, 16'd1027, 16'd38703, 16'd58332, 16'd14108, 16'd17814, 16'd8675, 16'd42759, 16'd35307, 16'd51802});
	test_expansion(128'h7d31de9cbc2992962e928d77d799b080, {16'd51510, 16'd55367, 16'd41507, 16'd7257, 16'd2081, 16'd13628, 16'd49160, 16'd18451, 16'd31604, 16'd48215, 16'd43476, 16'd31790, 16'd19766, 16'd7590, 16'd29039, 16'd53087, 16'd4681, 16'd28292, 16'd3999, 16'd63697, 16'd1646, 16'd64768, 16'd50949, 16'd23915, 16'd50120, 16'd6995});
	test_expansion(128'h92a4392f66a94aa15dabef64f86fcf21, {16'd50998, 16'd2055, 16'd37008, 16'd50170, 16'd18602, 16'd30731, 16'd52494, 16'd62339, 16'd61267, 16'd8590, 16'd64400, 16'd47014, 16'd33442, 16'd11694, 16'd54036, 16'd49158, 16'd11915, 16'd4697, 16'd14128, 16'd10969, 16'd62801, 16'd51177, 16'd50610, 16'd3807, 16'd58403, 16'd60414});
	test_expansion(128'h3efbd12332ff85a6887c30ef580fc788, {16'd33483, 16'd32756, 16'd5628, 16'd4310, 16'd21611, 16'd14058, 16'd564, 16'd45906, 16'd54578, 16'd33484, 16'd28585, 16'd50422, 16'd1410, 16'd30595, 16'd13882, 16'd13856, 16'd28095, 16'd49145, 16'd21787, 16'd60424, 16'd7426, 16'd62289, 16'd52941, 16'd27179, 16'd64668, 16'd42262});
	test_expansion(128'hd965737ebe82281ffd11c7c8fb819b3d, {16'd5783, 16'd56977, 16'd26068, 16'd1185, 16'd56033, 16'd30074, 16'd32671, 16'd52426, 16'd34594, 16'd16958, 16'd29576, 16'd17117, 16'd5406, 16'd9372, 16'd49662, 16'd44747, 16'd30644, 16'd34715, 16'd12647, 16'd46629, 16'd7700, 16'd20272, 16'd33052, 16'd44380, 16'd13391, 16'd49451});
	test_expansion(128'hee7cdd93e7e80ac7b4b3d3724990d84c, {16'd34271, 16'd57002, 16'd46871, 16'd61008, 16'd34724, 16'd45938, 16'd39536, 16'd8166, 16'd62352, 16'd59589, 16'd13115, 16'd38623, 16'd64148, 16'd11278, 16'd26048, 16'd40870, 16'd46963, 16'd38055, 16'd21907, 16'd35038, 16'd10819, 16'd15455, 16'd10279, 16'd19236, 16'd59412, 16'd18784});
	test_expansion(128'h21a9d9a1e17fca53dcb96674c42a1e1a, {16'd27203, 16'd11545, 16'd4806, 16'd18183, 16'd45900, 16'd7408, 16'd19478, 16'd47802, 16'd24293, 16'd36264, 16'd52505, 16'd38371, 16'd38240, 16'd16107, 16'd6047, 16'd20789, 16'd13507, 16'd56875, 16'd43764, 16'd14269, 16'd51255, 16'd11468, 16'd53235, 16'd4984, 16'd5495, 16'd20381});
	test_expansion(128'hb1463f4ffa35d51fb8e94fec10272143, {16'd10356, 16'd10272, 16'd60162, 16'd30950, 16'd36230, 16'd51541, 16'd8001, 16'd15838, 16'd60466, 16'd43912, 16'd16133, 16'd39219, 16'd41847, 16'd52265, 16'd30736, 16'd44716, 16'd40509, 16'd46426, 16'd49428, 16'd1130, 16'd20854, 16'd50381, 16'd37376, 16'd61894, 16'd46605, 16'd54611});
	test_expansion(128'hd4e459bf40489003201601352d805a43, {16'd6758, 16'd56442, 16'd4184, 16'd17682, 16'd55859, 16'd15924, 16'd60859, 16'd45651, 16'd42719, 16'd55211, 16'd28999, 16'd29544, 16'd20999, 16'd7892, 16'd46138, 16'd58496, 16'd30698, 16'd38498, 16'd54012, 16'd31108, 16'd52402, 16'd11838, 16'd44879, 16'd61516, 16'd21992, 16'd4668});
	test_expansion(128'h21ed5f9738d37db92e01b3fce98f0cfc, {16'd29031, 16'd8939, 16'd11386, 16'd8430, 16'd40595, 16'd48683, 16'd54362, 16'd41852, 16'd5004, 16'd46168, 16'd30700, 16'd37580, 16'd40258, 16'd7889, 16'd660, 16'd29030, 16'd17051, 16'd24873, 16'd8516, 16'd31942, 16'd61447, 16'd4568, 16'd52333, 16'd37835, 16'd60667, 16'd32840});
	test_expansion(128'hc5e213a44b02023f0bd84a1d5490f7f2, {16'd38913, 16'd22669, 16'd6727, 16'd63304, 16'd57731, 16'd43404, 16'd8015, 16'd49833, 16'd52366, 16'd23291, 16'd60285, 16'd3483, 16'd33700, 16'd17445, 16'd37322, 16'd30534, 16'd35283, 16'd26928, 16'd45446, 16'd16321, 16'd20641, 16'd3980, 16'd61058, 16'd43877, 16'd52581, 16'd36224});
	test_expansion(128'h3ef7c328fe5679de61fdf73ac15f8b36, {16'd59055, 16'd46622, 16'd52577, 16'd22741, 16'd11241, 16'd6777, 16'd48107, 16'd45798, 16'd51091, 16'd6043, 16'd42837, 16'd57967, 16'd35955, 16'd39822, 16'd25518, 16'd56376, 16'd46057, 16'd22094, 16'd60087, 16'd26015, 16'd56422, 16'd26090, 16'd56625, 16'd33984, 16'd51539, 16'd13622});
	test_expansion(128'h8f7b1ed95b562725cd65b2da46894e0f, {16'd20158, 16'd14464, 16'd50571, 16'd46859, 16'd316, 16'd18293, 16'd34547, 16'd36958, 16'd53481, 16'd19093, 16'd1612, 16'd55121, 16'd10696, 16'd20133, 16'd18292, 16'd37980, 16'd27838, 16'd10608, 16'd33148, 16'd6102, 16'd43470, 16'd40330, 16'd19974, 16'd12589, 16'd30800, 16'd36128});
	test_expansion(128'hf53fc5e923d731322419313f3c2b1d57, {16'd42184, 16'd13543, 16'd20917, 16'd24708, 16'd15636, 16'd48259, 16'd13, 16'd10055, 16'd23828, 16'd9841, 16'd57660, 16'd25962, 16'd56568, 16'd38051, 16'd34996, 16'd49512, 16'd48998, 16'd19864, 16'd43738, 16'd22721, 16'd19359, 16'd39064, 16'd31541, 16'd36153, 16'd38016, 16'd25427});
	test_expansion(128'h1b6efffd630a504ed7cfe36120532171, {16'd8416, 16'd19091, 16'd7471, 16'd9329, 16'd39923, 16'd56420, 16'd64602, 16'd3817, 16'd30956, 16'd48267, 16'd7552, 16'd58128, 16'd30668, 16'd60374, 16'd63, 16'd24840, 16'd15576, 16'd44148, 16'd8478, 16'd20396, 16'd9905, 16'd51571, 16'd58461, 16'd5340, 16'd51310, 16'd46080});
	test_expansion(128'h07b574b55801a7e20ef4e7a8d4d840fd, {16'd57781, 16'd58483, 16'd15043, 16'd40699, 16'd14949, 16'd65245, 16'd64631, 16'd26050, 16'd55413, 16'd13931, 16'd53638, 16'd55611, 16'd16154, 16'd58268, 16'd15254, 16'd52916, 16'd35011, 16'd20211, 16'd41123, 16'd58115, 16'd60170, 16'd14707, 16'd6553, 16'd49323, 16'd34463, 16'd36235});
	test_expansion(128'h755c7909ef8488edbe1db12ebd467252, {16'd40922, 16'd13552, 16'd44208, 16'd37169, 16'd52242, 16'd15641, 16'd30939, 16'd16744, 16'd40013, 16'd58947, 16'd4762, 16'd60321, 16'd25230, 16'd64355, 16'd21190, 16'd50004, 16'd20406, 16'd57534, 16'd36541, 16'd55800, 16'd65310, 16'd42024, 16'd2975, 16'd30420, 16'd17489, 16'd39149});
	test_expansion(128'h155b870931ac833f424a6ef516a6bc25, {16'd45274, 16'd54057, 16'd58588, 16'd33492, 16'd39521, 16'd28653, 16'd88, 16'd3716, 16'd55137, 16'd26075, 16'd26684, 16'd25332, 16'd33094, 16'd22827, 16'd36248, 16'd54499, 16'd41260, 16'd15997, 16'd49107, 16'd6463, 16'd37521, 16'd43899, 16'd52305, 16'd19074, 16'd64453, 16'd41178});
	test_expansion(128'h071baf9810a31adc3694556675abc1c5, {16'd20020, 16'd828, 16'd24747, 16'd42621, 16'd25375, 16'd4222, 16'd6315, 16'd22286, 16'd20572, 16'd18960, 16'd24641, 16'd43848, 16'd55090, 16'd25743, 16'd35918, 16'd16211, 16'd37296, 16'd8958, 16'd20764, 16'd27061, 16'd6861, 16'd29485, 16'd63047, 16'd21052, 16'd63770, 16'd37881});
	test_expansion(128'h6e1d814022345466ea57bd5bf670e5f3, {16'd53963, 16'd10115, 16'd2835, 16'd37960, 16'd17892, 16'd33298, 16'd15858, 16'd10457, 16'd6754, 16'd60151, 16'd25693, 16'd6086, 16'd9108, 16'd28046, 16'd54694, 16'd50145, 16'd55094, 16'd29860, 16'd29876, 16'd60442, 16'd15769, 16'd8432, 16'd26922, 16'd30710, 16'd63819, 16'd27623});
	test_expansion(128'hd844a122e2b741123bdfc0b0f7579e7b, {16'd28428, 16'd22186, 16'd14914, 16'd13123, 16'd63289, 16'd37148, 16'd55676, 16'd65160, 16'd26777, 16'd11779, 16'd40001, 16'd1814, 16'd27105, 16'd54792, 16'd14433, 16'd6806, 16'd37516, 16'd27940, 16'd51344, 16'd6425, 16'd11482, 16'd51661, 16'd28983, 16'd6939, 16'd41994, 16'd20766});
	test_expansion(128'h01897309f19cb4bbd41e9e77d5791d9b, {16'd10563, 16'd30246, 16'd38580, 16'd51729, 16'd36963, 16'd40528, 16'd58577, 16'd34332, 16'd8956, 16'd4745, 16'd1758, 16'd48872, 16'd13886, 16'd15121, 16'd43194, 16'd60690, 16'd62230, 16'd63670, 16'd49321, 16'd13274, 16'd8178, 16'd28994, 16'd58724, 16'd27363, 16'd13263, 16'd54536});
	test_expansion(128'hf98e9ab1d0a93c61bb6e7e8ef851364a, {16'd20836, 16'd47186, 16'd11154, 16'd57332, 16'd62506, 16'd32622, 16'd18978, 16'd32336, 16'd31287, 16'd3674, 16'd25325, 16'd50528, 16'd13057, 16'd55526, 16'd64245, 16'd65212, 16'd62703, 16'd11451, 16'd50068, 16'd21109, 16'd22662, 16'd57807, 16'd34197, 16'd61942, 16'd52591, 16'd29477});
	test_expansion(128'h9e1694e32ad45bb9e64e0918f05f5881, {16'd63680, 16'd51694, 16'd54985, 16'd8381, 16'd51295, 16'd48965, 16'd21140, 16'd34412, 16'd8912, 16'd33816, 16'd33307, 16'd61220, 16'd54518, 16'd664, 16'd46689, 16'd6505, 16'd13762, 16'd31559, 16'd46405, 16'd35973, 16'd887, 16'd35850, 16'd624, 16'd8702, 16'd25564, 16'd32865});
	test_expansion(128'hc3f9b12e9946a08dd1afb122b944a276, {16'd25821, 16'd8472, 16'd60590, 16'd54352, 16'd37136, 16'd52681, 16'd9971, 16'd20306, 16'd33890, 16'd41114, 16'd30115, 16'd31341, 16'd23336, 16'd49050, 16'd6357, 16'd35578, 16'd35888, 16'd27077, 16'd57065, 16'd14859, 16'd32261, 16'd21949, 16'd62521, 16'd47170, 16'd47291, 16'd33277});
	test_expansion(128'h78ac867c2c4ff0d2095e1f0d65ce10ef, {16'd48065, 16'd33144, 16'd18154, 16'd24441, 16'd8211, 16'd20189, 16'd50651, 16'd60949, 16'd31911, 16'd18989, 16'd32010, 16'd22643, 16'd9722, 16'd36973, 16'd21794, 16'd11374, 16'd19107, 16'd52362, 16'd40796, 16'd31804, 16'd19246, 16'd47631, 16'd9712, 16'd57542, 16'd32748, 16'd7293});
	test_expansion(128'hc3b21b86157674878cf86cba09624b68, {16'd61406, 16'd31866, 16'd12546, 16'd53923, 16'd45524, 16'd55811, 16'd50508, 16'd58758, 16'd49334, 16'd46196, 16'd2009, 16'd1085, 16'd55416, 16'd32364, 16'd38795, 16'd40815, 16'd23021, 16'd17148, 16'd33821, 16'd63541, 16'd47048, 16'd17057, 16'd45813, 16'd3988, 16'd38637, 16'd33809});
	test_expansion(128'h6a6ad7588d89a5cc8c72dc499bcdd0c4, {16'd12160, 16'd52101, 16'd7767, 16'd25851, 16'd59752, 16'd56039, 16'd33834, 16'd62209, 16'd2490, 16'd30766, 16'd29193, 16'd20262, 16'd32881, 16'd62152, 16'd14435, 16'd42811, 16'd10071, 16'd42559, 16'd47764, 16'd39348, 16'd5634, 16'd39792, 16'd20523, 16'd47809, 16'd15104, 16'd26116});
	test_expansion(128'hb3224b67fee35d0af6670496917ee2ea, {16'd6789, 16'd43348, 16'd867, 16'd26859, 16'd7321, 16'd20483, 16'd1959, 16'd63535, 16'd56874, 16'd51436, 16'd50463, 16'd2195, 16'd54395, 16'd36676, 16'd44115, 16'd54547, 16'd51986, 16'd15714, 16'd61204, 16'd63405, 16'd65137, 16'd30154, 16'd53726, 16'd62478, 16'd46911, 16'd60610});
	test_expansion(128'h226ba30f538e78c824c7a3e857a3118d, {16'd2658, 16'd62782, 16'd16988, 16'd48718, 16'd5982, 16'd3526, 16'd3049, 16'd45943, 16'd58924, 16'd39462, 16'd29864, 16'd45010, 16'd35063, 16'd6721, 16'd52465, 16'd36113, 16'd32779, 16'd63568, 16'd29678, 16'd923, 16'd38411, 16'd22877, 16'd3856, 16'd30873, 16'd48129, 16'd5070});
	test_expansion(128'h5d86560140ec5138f40a2fc6ec3d6b80, {16'd59434, 16'd3705, 16'd20072, 16'd34834, 16'd21681, 16'd16395, 16'd55170, 16'd43333, 16'd35458, 16'd25259, 16'd59415, 16'd31126, 16'd26382, 16'd28855, 16'd2610, 16'd26337, 16'd41971, 16'd9929, 16'd36957, 16'd52304, 16'd28587, 16'd29335, 16'd5814, 16'd30778, 16'd62447, 16'd44990});
	test_expansion(128'h6b1d1e8bdd4de04a6b0e03ee20151ac2, {16'd57216, 16'd27483, 16'd53930, 16'd10926, 16'd975, 16'd60492, 16'd1100, 16'd57153, 16'd12672, 16'd31569, 16'd14936, 16'd26878, 16'd2942, 16'd54977, 16'd50259, 16'd29990, 16'd22454, 16'd31557, 16'd59720, 16'd31754, 16'd65371, 16'd65100, 16'd30124, 16'd56954, 16'd16062, 16'd57607});
	test_expansion(128'h13d90a9573d278a36edadca602f8d50b, {16'd57901, 16'd27639, 16'd60932, 16'd19142, 16'd15399, 16'd50382, 16'd59530, 16'd52194, 16'd41402, 16'd39673, 16'd39407, 16'd19401, 16'd38896, 16'd3581, 16'd30744, 16'd50190, 16'd42973, 16'd61303, 16'd49908, 16'd65251, 16'd27949, 16'd31227, 16'd5067, 16'd44649, 16'd36088, 16'd29990});
	test_expansion(128'h1b0c7041736348d455c9e03116edc073, {16'd1281, 16'd35062, 16'd33967, 16'd51815, 16'd48984, 16'd46690, 16'd43484, 16'd36107, 16'd63970, 16'd15644, 16'd44070, 16'd46027, 16'd21536, 16'd19941, 16'd6082, 16'd8329, 16'd36228, 16'd41147, 16'd48674, 16'd64935, 16'd34477, 16'd30107, 16'd45194, 16'd55718, 16'd36228, 16'd47824});
	test_expansion(128'h4dc1d4a8699c1b1bd7beb60c0f1747af, {16'd24752, 16'd13199, 16'd44627, 16'd59445, 16'd53335, 16'd14515, 16'd52328, 16'd43565, 16'd33122, 16'd36061, 16'd10292, 16'd52782, 16'd19790, 16'd3784, 16'd59508, 16'd53637, 16'd3089, 16'd45808, 16'd24370, 16'd28923, 16'd4968, 16'd64768, 16'd6296, 16'd65465, 16'd36362, 16'd8612});
	test_expansion(128'h4aa2ec5da0b8ff5bfe08f865d916ee1a, {16'd30657, 16'd59781, 16'd11486, 16'd2318, 16'd10016, 16'd8975, 16'd55687, 16'd6164, 16'd3667, 16'd16043, 16'd16670, 16'd13422, 16'd4728, 16'd54724, 16'd65464, 16'd44249, 16'd44427, 16'd53990, 16'd46842, 16'd64309, 16'd47121, 16'd28991, 16'd23302, 16'd16101, 16'd21219, 16'd63294});
	test_expansion(128'he6c5e38671291834cdc0c536f908b80c, {16'd9542, 16'd20368, 16'd43502, 16'd1038, 16'd29742, 16'd31800, 16'd33866, 16'd20725, 16'd46679, 16'd31680, 16'd44335, 16'd65180, 16'd57190, 16'd12161, 16'd63589, 16'd48937, 16'd44251, 16'd57543, 16'd58489, 16'd52076, 16'd45201, 16'd17396, 16'd7451, 16'd34219, 16'd26833, 16'd43398});
	test_expansion(128'h3e510af271085cd5fc205d7de8e58457, {16'd29137, 16'd45712, 16'd6650, 16'd3233, 16'd44593, 16'd61810, 16'd5119, 16'd51815, 16'd8308, 16'd42133, 16'd1781, 16'd57123, 16'd49363, 16'd59266, 16'd27246, 16'd20401, 16'd22689, 16'd61035, 16'd19021, 16'd15265, 16'd2205, 16'd36595, 16'd62332, 16'd23841, 16'd61724, 16'd50462});
	test_expansion(128'hb11196d11a8a939459119697ce5a441d, {16'd19155, 16'd28370, 16'd30462, 16'd46670, 16'd17503, 16'd25392, 16'd10158, 16'd41540, 16'd15400, 16'd60486, 16'd17712, 16'd44081, 16'd23616, 16'd44635, 16'd22600, 16'd62389, 16'd55502, 16'd57838, 16'd61189, 16'd43897, 16'd64829, 16'd25934, 16'd46574, 16'd33213, 16'd8292, 16'd1057});
	test_expansion(128'hc82f6fdae9bbecb5e028af7e3070def0, {16'd34277, 16'd11893, 16'd16444, 16'd61447, 16'd53662, 16'd52804, 16'd30995, 16'd15849, 16'd17138, 16'd45845, 16'd36789, 16'd35656, 16'd28986, 16'd30682, 16'd29266, 16'd48976, 16'd274, 16'd33107, 16'd17614, 16'd55781, 16'd43147, 16'd47815, 16'd5223, 16'd38484, 16'd10344, 16'd35201});
	test_expansion(128'hbca3f9acb39f188101e657bb362209d1, {16'd21950, 16'd22638, 16'd11911, 16'd12103, 16'd49759, 16'd12208, 16'd1475, 16'd44796, 16'd29093, 16'd41298, 16'd40221, 16'd42706, 16'd35275, 16'd56634, 16'd17130, 16'd32184, 16'd38824, 16'd12321, 16'd45382, 16'd29601, 16'd39896, 16'd18618, 16'd43853, 16'd40755, 16'd37018, 16'd7702});
	test_expansion(128'h51f3a5486e4f5a5370782052a26f1156, {16'd44224, 16'd21999, 16'd262, 16'd61066, 16'd7344, 16'd59108, 16'd52063, 16'd22180, 16'd38932, 16'd21271, 16'd48935, 16'd49555, 16'd58356, 16'd23760, 16'd38189, 16'd40863, 16'd49518, 16'd35989, 16'd36603, 16'd54387, 16'd24328, 16'd49173, 16'd52601, 16'd61450, 16'd48505, 16'd25790});
	test_expansion(128'h16ed6cb0e277b63d2ed5bb2ebe6a27d4, {16'd9906, 16'd28990, 16'd64929, 16'd45480, 16'd26926, 16'd47215, 16'd26231, 16'd46313, 16'd62241, 16'd38838, 16'd58362, 16'd49676, 16'd30827, 16'd25994, 16'd6335, 16'd8599, 16'd24951, 16'd64806, 16'd24962, 16'd23788, 16'd21638, 16'd44121, 16'd33131, 16'd29874, 16'd7568, 16'd54240});
	test_expansion(128'h71fe60563c2441485688cee18b44be15, {16'd34904, 16'd28282, 16'd61092, 16'd56451, 16'd27516, 16'd62704, 16'd34495, 16'd2597, 16'd26723, 16'd59156, 16'd58536, 16'd13233, 16'd44260, 16'd60248, 16'd44255, 16'd51211, 16'd1047, 16'd8742, 16'd7166, 16'd30967, 16'd20060, 16'd53539, 16'd22571, 16'd1108, 16'd29812, 16'd27316});
	test_expansion(128'h6304a4d01372373ba012bd57ae72fa33, {16'd41376, 16'd48163, 16'd35491, 16'd4635, 16'd42087, 16'd18278, 16'd63892, 16'd12569, 16'd27107, 16'd33928, 16'd54105, 16'd8569, 16'd55836, 16'd38643, 16'd15894, 16'd56802, 16'd46189, 16'd5747, 16'd63466, 16'd36538, 16'd31116, 16'd48887, 16'd21675, 16'd24656, 16'd25918, 16'd20481});
	test_expansion(128'h9aed8d257f0aeab381716605ea219bd3, {16'd43740, 16'd21916, 16'd49612, 16'd55467, 16'd63015, 16'd5979, 16'd57230, 16'd55588, 16'd12634, 16'd46689, 16'd33138, 16'd59810, 16'd64703, 16'd16881, 16'd30512, 16'd59682, 16'd13439, 16'd24749, 16'd1716, 16'd61495, 16'd25543, 16'd20078, 16'd60768, 16'd35822, 16'd55721, 16'd509});
	test_expansion(128'hb85627f46793b615d7502bc71104072d, {16'd16318, 16'd24071, 16'd45345, 16'd53075, 16'd53574, 16'd17181, 16'd60962, 16'd53165, 16'd45826, 16'd46649, 16'd705, 16'd58392, 16'd58897, 16'd22409, 16'd34041, 16'd12365, 16'd19287, 16'd14306, 16'd43281, 16'd60150, 16'd32807, 16'd22463, 16'd46233, 16'd13251, 16'd63710, 16'd63933});
	test_expansion(128'h153fe91c7f321f89ea155e2b63cd23b9, {16'd1746, 16'd55666, 16'd43512, 16'd11477, 16'd28023, 16'd65234, 16'd42747, 16'd8826, 16'd18823, 16'd50413, 16'd44365, 16'd34853, 16'd12289, 16'd29772, 16'd26498, 16'd14982, 16'd44350, 16'd6874, 16'd53688, 16'd40077, 16'd4935, 16'd58381, 16'd51300, 16'd636, 16'd24697, 16'd48785});
	test_expansion(128'h234951a286fff9d4c1f87f6630c528f4, {16'd24634, 16'd38311, 16'd33935, 16'd7663, 16'd642, 16'd13458, 16'd41048, 16'd5318, 16'd19077, 16'd13388, 16'd33429, 16'd36707, 16'd11917, 16'd55575, 16'd40963, 16'd45141, 16'd50330, 16'd7766, 16'd28775, 16'd62968, 16'd51686, 16'd63484, 16'd63307, 16'd15309, 16'd51877, 16'd2182});
	test_expansion(128'hc5be06d6c8c4dd516314c1305a0f1127, {16'd36819, 16'd18040, 16'd51284, 16'd7054, 16'd34664, 16'd41153, 16'd34965, 16'd27575, 16'd9338, 16'd9592, 16'd15087, 16'd17495, 16'd25241, 16'd12075, 16'd54394, 16'd36626, 16'd15434, 16'd13270, 16'd29979, 16'd15587, 16'd37652, 16'd5387, 16'd29442, 16'd28859, 16'd61337, 16'd64422});
	test_expansion(128'hed61454881d3b5db1f5e80cd41bdd03d, {16'd37293, 16'd39867, 16'd52524, 16'd7647, 16'd61038, 16'd4, 16'd1152, 16'd18236, 16'd49426, 16'd13811, 16'd51642, 16'd25010, 16'd30260, 16'd28193, 16'd31131, 16'd45512, 16'd16619, 16'd16334, 16'd52780, 16'd61063, 16'd7244, 16'd16525, 16'd54754, 16'd5621, 16'd36405, 16'd2165});
	test_expansion(128'hd2519f3a82a518e50cd7dcdfd99c8bf0, {16'd4285, 16'd37776, 16'd21917, 16'd60159, 16'd48689, 16'd16355, 16'd40955, 16'd37371, 16'd37420, 16'd60468, 16'd23629, 16'd30585, 16'd60170, 16'd16294, 16'd65307, 16'd36485, 16'd63936, 16'd41937, 16'd14147, 16'd6288, 16'd36973, 16'd50396, 16'd36769, 16'd48824, 16'd37620, 16'd37819});
	test_expansion(128'ha5fc5048a439b32aadaed65a9eae4545, {16'd48345, 16'd27374, 16'd63626, 16'd38052, 16'd21666, 16'd24991, 16'd59934, 16'd47262, 16'd18586, 16'd55902, 16'd52354, 16'd9510, 16'd32955, 16'd60459, 16'd30241, 16'd33746, 16'd27796, 16'd52200, 16'd21957, 16'd57762, 16'd21706, 16'd63663, 16'd60803, 16'd40980, 16'd29139, 16'd22097});
	test_expansion(128'hfd5a6c96b7f738bb6d73e18e89c4f70e, {16'd54603, 16'd44414, 16'd37979, 16'd33783, 16'd52072, 16'd44457, 16'd49458, 16'd59058, 16'd57281, 16'd60443, 16'd20310, 16'd320, 16'd58533, 16'd42469, 16'd56793, 16'd16972, 16'd23988, 16'd30374, 16'd58339, 16'd35356, 16'd34481, 16'd12913, 16'd47463, 16'd13347, 16'd1773, 16'd5064});
	test_expansion(128'h3f8336fcf8cfb25270611a0451b1f80f, {16'd20976, 16'd36533, 16'd41620, 16'd46719, 16'd36912, 16'd23528, 16'd28799, 16'd22706, 16'd51396, 16'd160, 16'd57765, 16'd44542, 16'd58993, 16'd47026, 16'd9653, 16'd16403, 16'd65423, 16'd16448, 16'd998, 16'd41337, 16'd39004, 16'd26860, 16'd8082, 16'd14798, 16'd14609, 16'd59179});
	test_expansion(128'h0cdcb8fc294972c1aec2caa033e760d2, {16'd53744, 16'd37031, 16'd20744, 16'd43441, 16'd8030, 16'd9590, 16'd21219, 16'd60721, 16'd48512, 16'd31866, 16'd561, 16'd14736, 16'd32535, 16'd35066, 16'd58791, 16'd47270, 16'd41148, 16'd40304, 16'd8926, 16'd16461, 16'd25974, 16'd65025, 16'd38844, 16'd10680, 16'd2675, 16'd56053});
	test_expansion(128'hc26f93b3f9a6fe430c428840728a5ec4, {16'd44524, 16'd38071, 16'd21989, 16'd1327, 16'd32332, 16'd21754, 16'd11506, 16'd34598, 16'd57064, 16'd19687, 16'd36798, 16'd5079, 16'd36274, 16'd22811, 16'd49513, 16'd4810, 16'd26122, 16'd54379, 16'd5364, 16'd20126, 16'd14179, 16'd38650, 16'd36234, 16'd40083, 16'd40571, 16'd7285});
	test_expansion(128'hd70f7dad2b5f4f5f69cba919890b3269, {16'd5754, 16'd50141, 16'd15179, 16'd37908, 16'd4034, 16'd28477, 16'd50801, 16'd27691, 16'd55899, 16'd9952, 16'd18062, 16'd44812, 16'd43012, 16'd3400, 16'd52244, 16'd49649, 16'd9931, 16'd12106, 16'd19330, 16'd21144, 16'd50120, 16'd58729, 16'd48275, 16'd20223, 16'd28261, 16'd18887});
	test_expansion(128'h46a85fb6b2b93ae9d5786ee4eca061f8, {16'd60217, 16'd5675, 16'd2837, 16'd3881, 16'd31643, 16'd39819, 16'd3797, 16'd12052, 16'd51284, 16'd19769, 16'd20304, 16'd36427, 16'd27259, 16'd17628, 16'd18894, 16'd61322, 16'd19805, 16'd39198, 16'd25021, 16'd10852, 16'd3386, 16'd62073, 16'd26394, 16'd14349, 16'd32720, 16'd63446});
	test_expansion(128'h10e894cd0059b19a36ecdb9be14a04ea, {16'd42436, 16'd15988, 16'd51560, 16'd63725, 16'd7325, 16'd21133, 16'd45861, 16'd60771, 16'd12100, 16'd62871, 16'd47916, 16'd53075, 16'd57628, 16'd45505, 16'd18695, 16'd52104, 16'd9079, 16'd8492, 16'd56831, 16'd22085, 16'd55478, 16'd26966, 16'd23694, 16'd58914, 16'd6756, 16'd45172});
	test_expansion(128'h94f9314982d29fc4d21757989bb01f59, {16'd3521, 16'd23288, 16'd20131, 16'd57631, 16'd19151, 16'd47459, 16'd43867, 16'd58373, 16'd46620, 16'd48277, 16'd7399, 16'd25552, 16'd62094, 16'd24186, 16'd51153, 16'd41039, 16'd21156, 16'd53922, 16'd19202, 16'd17470, 16'd7294, 16'd60255, 16'd37196, 16'd16700, 16'd33091, 16'd28573});
	test_expansion(128'h58ae88ed9772d0397378dc9edc680ebf, {16'd17785, 16'd11128, 16'd20945, 16'd58155, 16'd30991, 16'd35777, 16'd991, 16'd53647, 16'd1589, 16'd11154, 16'd12778, 16'd33679, 16'd62290, 16'd8624, 16'd59961, 16'd19652, 16'd20462, 16'd11862, 16'd37110, 16'd31612, 16'd5809, 16'd24975, 16'd6591, 16'd21609, 16'd9019, 16'd10300});
	test_expansion(128'he7d7e9254aa1118dfcdc4164de7e830a, {16'd55970, 16'd20, 16'd61100, 16'd5373, 16'd45431, 16'd39295, 16'd30384, 16'd32022, 16'd10352, 16'd51885, 16'd23551, 16'd35225, 16'd5094, 16'd13392, 16'd22328, 16'd39203, 16'd65438, 16'd6434, 16'd57735, 16'd23297, 16'd32346, 16'd14409, 16'd46337, 16'd42714, 16'd28289, 16'd13716});
	test_expansion(128'h9e8ba293865d3ea814c5ecf74e038e7e, {16'd43220, 16'd27819, 16'd24406, 16'd2132, 16'd7912, 16'd32999, 16'd30898, 16'd19872, 16'd26905, 16'd7783, 16'd29121, 16'd26077, 16'd40546, 16'd12944, 16'd45200, 16'd2605, 16'd1189, 16'd10350, 16'd52028, 16'd22401, 16'd5016, 16'd53477, 16'd46851, 16'd50006, 16'd30974, 16'd31128});
	test_expansion(128'h61e8cf497128a34410b4a26e0a8a98a9, {16'd20341, 16'd7710, 16'd40926, 16'd16606, 16'd45442, 16'd32778, 16'd38797, 16'd60827, 16'd64457, 16'd27823, 16'd2191, 16'd50053, 16'd51247, 16'd42057, 16'd30499, 16'd25854, 16'd41568, 16'd23700, 16'd51046, 16'd19198, 16'd54679, 16'd35213, 16'd44339, 16'd11137, 16'd43399, 16'd17355});
	test_expansion(128'h46fe4772d0d067e9b66750a31dd611cc, {16'd39223, 16'd15716, 16'd175, 16'd29074, 16'd13743, 16'd18642, 16'd58048, 16'd14490, 16'd47192, 16'd2144, 16'd10893, 16'd1504, 16'd14471, 16'd10622, 16'd50129, 16'd30501, 16'd10030, 16'd1097, 16'd25109, 16'd62157, 16'd61064, 16'd48242, 16'd56390, 16'd20634, 16'd60911, 16'd3785});
	test_expansion(128'h356837e888b5077387177277fc26761c, {16'd64414, 16'd44724, 16'd6342, 16'd25525, 16'd37444, 16'd20163, 16'd39463, 16'd39452, 16'd43174, 16'd9350, 16'd20729, 16'd160, 16'd44606, 16'd57018, 16'd34775, 16'd32190, 16'd1888, 16'd29829, 16'd13820, 16'd61437, 16'd38962, 16'd7913, 16'd30894, 16'd23021, 16'd58231, 16'd28704});
	test_expansion(128'hb9fb79202755c2ae7d517fc2a930f322, {16'd63141, 16'd29788, 16'd9018, 16'd8409, 16'd1756, 16'd1672, 16'd27185, 16'd9208, 16'd1606, 16'd6339, 16'd53422, 16'd33134, 16'd57512, 16'd53281, 16'd29632, 16'd16613, 16'd58563, 16'd10785, 16'd5616, 16'd52699, 16'd12193, 16'd52620, 16'd31769, 16'd21331, 16'd14316, 16'd38931});
	test_expansion(128'h9af1fbda57ec7ab7b403c4e0d06ca161, {16'd31757, 16'd14950, 16'd52752, 16'd34293, 16'd60031, 16'd16252, 16'd19301, 16'd28545, 16'd51557, 16'd34726, 16'd20115, 16'd61738, 16'd2344, 16'd25625, 16'd57576, 16'd35154, 16'd25827, 16'd8014, 16'd1352, 16'd25793, 16'd56893, 16'd51239, 16'd53046, 16'd40825, 16'd33931, 16'd55339});
	test_expansion(128'h77f8986bf52a0f0057a1e23eccdf827f, {16'd19083, 16'd45282, 16'd23573, 16'd56131, 16'd14107, 16'd58834, 16'd32438, 16'd27063, 16'd35505, 16'd58482, 16'd39275, 16'd4193, 16'd37857, 16'd20434, 16'd39820, 16'd2462, 16'd10739, 16'd45266, 16'd32796, 16'd36818, 16'd2310, 16'd62760, 16'd64212, 16'd26520, 16'd13907, 16'd3897});
	test_expansion(128'hd4bb1a316ef5f9c0d6faf1bc13553558, {16'd62378, 16'd43609, 16'd47759, 16'd7981, 16'd58904, 16'd47107, 16'd695, 16'd16636, 16'd19413, 16'd54368, 16'd8994, 16'd59408, 16'd50873, 16'd58664, 16'd59251, 16'd29787, 16'd63805, 16'd1781, 16'd26954, 16'd40475, 16'd16135, 16'd11618, 16'd1466, 16'd26057, 16'd6666, 16'd504});
	test_expansion(128'he2da798d39b22c0528b25fb38cd9b92c, {16'd56924, 16'd57429, 16'd2497, 16'd21437, 16'd39085, 16'd23725, 16'd28481, 16'd8086, 16'd40391, 16'd51366, 16'd56222, 16'd50520, 16'd23948, 16'd6703, 16'd48057, 16'd56828, 16'd19764, 16'd56102, 16'd36275, 16'd5983, 16'd61885, 16'd13383, 16'd23430, 16'd35882, 16'd760, 16'd25946});
	test_expansion(128'hcde0b827672f2352c4ef700bee668c5d, {16'd9674, 16'd56850, 16'd11112, 16'd36357, 16'd49035, 16'd12502, 16'd24366, 16'd14895, 16'd36058, 16'd40715, 16'd17472, 16'd50794, 16'd47803, 16'd36731, 16'd4972, 16'd609, 16'd54888, 16'd43405, 16'd7863, 16'd43805, 16'd28139, 16'd55385, 16'd1739, 16'd1157, 16'd34906, 16'd12981});
	test_expansion(128'hba64443600fda43863879586e8ceb1a6, {16'd48045, 16'd453, 16'd51235, 16'd34501, 16'd50575, 16'd50970, 16'd25324, 16'd9560, 16'd42431, 16'd25863, 16'd36247, 16'd3164, 16'd16149, 16'd6745, 16'd59862, 16'd57781, 16'd42951, 16'd12535, 16'd59427, 16'd10690, 16'd36983, 16'd10656, 16'd61026, 16'd9743, 16'd47308, 16'd25387});
	test_expansion(128'hf87841af983b41f9d1b6615ae0520261, {16'd25410, 16'd44319, 16'd5399, 16'd1865, 16'd31169, 16'd34445, 16'd62276, 16'd53161, 16'd30953, 16'd3398, 16'd53778, 16'd43259, 16'd37088, 16'd58458, 16'd27810, 16'd16847, 16'd3464, 16'd33586, 16'd16740, 16'd4872, 16'd12430, 16'd63267, 16'd31906, 16'd9183, 16'd26019, 16'd11813});
	test_expansion(128'h3264aebdaea37f5c8fd0c21d6458b66b, {16'd35, 16'd16025, 16'd15694, 16'd36186, 16'd11192, 16'd3514, 16'd52885, 16'd47013, 16'd60029, 16'd64863, 16'd61185, 16'd42927, 16'd37526, 16'd5050, 16'd27232, 16'd43052, 16'd21483, 16'd43205, 16'd46532, 16'd2733, 16'd48190, 16'd20966, 16'd27210, 16'd47099, 16'd20154, 16'd34273});
	test_expansion(128'h304b106e50a3fe7a6332d44e22aee9af, {16'd56389, 16'd19790, 16'd24608, 16'd10124, 16'd36444, 16'd41864, 16'd61167, 16'd56164, 16'd12765, 16'd49622, 16'd14188, 16'd19948, 16'd41722, 16'd37335, 16'd61878, 16'd54391, 16'd17501, 16'd48457, 16'd16299, 16'd60379, 16'd58482, 16'd40948, 16'd39987, 16'd17223, 16'd57561, 16'd26517});
	test_expansion(128'h36c74f76f474fe62e8a071710acb7586, {16'd57078, 16'd37555, 16'd3415, 16'd46414, 16'd15252, 16'd3210, 16'd24567, 16'd14813, 16'd48665, 16'd33420, 16'd1944, 16'd33792, 16'd27683, 16'd39848, 16'd39721, 16'd3964, 16'd31381, 16'd65396, 16'd57728, 16'd5856, 16'd64411, 16'd7688, 16'd21301, 16'd37431, 16'd13666, 16'd59672});
	test_expansion(128'hb123049686fc5c1a28e03dd06bb53d1a, {16'd4515, 16'd5686, 16'd20594, 16'd33106, 16'd62609, 16'd29582, 16'd41959, 16'd7228, 16'd28560, 16'd28251, 16'd61703, 16'd55911, 16'd3002, 16'd5135, 16'd30097, 16'd64910, 16'd13616, 16'd51601, 16'd58199, 16'd18195, 16'd57100, 16'd12078, 16'd13966, 16'd48471, 16'd15046, 16'd31997});
	test_expansion(128'hfd9bf920b447b1a507529f5144dc57bd, {16'd24319, 16'd33239, 16'd51722, 16'd10575, 16'd20578, 16'd65354, 16'd56873, 16'd64122, 16'd8662, 16'd12630, 16'd52193, 16'd60461, 16'd19503, 16'd45232, 16'd48383, 16'd32326, 16'd39018, 16'd3511, 16'd53443, 16'd9038, 16'd48347, 16'd63450, 16'd45621, 16'd34905, 16'd31372, 16'd44373});
	test_expansion(128'h84aa1034827ff9a39de34a1e10f173e0, {16'd8071, 16'd51097, 16'd62935, 16'd11686, 16'd63942, 16'd19721, 16'd62832, 16'd63755, 16'd27721, 16'd58989, 16'd28029, 16'd42491, 16'd64776, 16'd54416, 16'd21064, 16'd18344, 16'd38008, 16'd37930, 16'd29115, 16'd17237, 16'd7668, 16'd33191, 16'd43623, 16'd32418, 16'd24406, 16'd63916});
	test_expansion(128'h348c1f03b22e468737731df7657f3528, {16'd33616, 16'd7542, 16'd38601, 16'd24747, 16'd18553, 16'd65070, 16'd48531, 16'd56594, 16'd47108, 16'd38435, 16'd30580, 16'd30129, 16'd59138, 16'd12096, 16'd49248, 16'd9378, 16'd18880, 16'd58390, 16'd28971, 16'd38083, 16'd8576, 16'd50370, 16'd17497, 16'd46872, 16'd45756, 16'd7113});
	test_expansion(128'hd483207cb21f5dd0bce1f8fd00c50882, {16'd21694, 16'd20598, 16'd25331, 16'd8818, 16'd18869, 16'd51257, 16'd60777, 16'd50851, 16'd28245, 16'd33214, 16'd65476, 16'd46104, 16'd31438, 16'd12077, 16'd61495, 16'd27329, 16'd20591, 16'd45710, 16'd47400, 16'd22572, 16'd850, 16'd3292, 16'd63367, 16'd27737, 16'd55687, 16'd490});
	test_expansion(128'h261c06dddf9af7f83bc337212e43de72, {16'd13521, 16'd40091, 16'd33845, 16'd4397, 16'd10439, 16'd16348, 16'd16702, 16'd43473, 16'd23824, 16'd49205, 16'd6751, 16'd38492, 16'd37097, 16'd2957, 16'd47364, 16'd2671, 16'd57847, 16'd46917, 16'd63493, 16'd55079, 16'd27556, 16'd61421, 16'd28140, 16'd37326, 16'd7689, 16'd34238});
	test_expansion(128'h48b59c7d01f0c8a5d51df673a813f660, {16'd1959, 16'd35225, 16'd26951, 16'd17648, 16'd60451, 16'd45046, 16'd39045, 16'd24319, 16'd19995, 16'd45861, 16'd4481, 16'd13197, 16'd34676, 16'd33712, 16'd14583, 16'd9729, 16'd53829, 16'd43509, 16'd5369, 16'd41012, 16'd35651, 16'd53153, 16'd30305, 16'd786, 16'd47353, 16'd54042});
	test_expansion(128'h98424c5f5375e86ffa4c17eefca26575, {16'd46211, 16'd11502, 16'd12440, 16'd14544, 16'd20611, 16'd63888, 16'd14971, 16'd59300, 16'd35080, 16'd37371, 16'd57695, 16'd36342, 16'd9993, 16'd32501, 16'd8121, 16'd53008, 16'd4874, 16'd39560, 16'd56370, 16'd19778, 16'd31435, 16'd25404, 16'd13303, 16'd9661, 16'd57955, 16'd14310});
	test_expansion(128'h8a1f05c584317064dbf8f4f22e592b29, {16'd1568, 16'd63112, 16'd61360, 16'd22062, 16'd4953, 16'd57950, 16'd36096, 16'd6708, 16'd5886, 16'd43822, 16'd59740, 16'd59424, 16'd40548, 16'd4402, 16'd8594, 16'd38404, 16'd49526, 16'd60717, 16'd30883, 16'd12624, 16'd16103, 16'd54147, 16'd32545, 16'd20417, 16'd36707, 16'd36621});
	test_expansion(128'hd3201718ed3e1f049ae4819f97474076, {16'd58029, 16'd29551, 16'd9577, 16'd13138, 16'd53726, 16'd45992, 16'd10413, 16'd11807, 16'd8952, 16'd60890, 16'd50194, 16'd32594, 16'd59589, 16'd52190, 16'd44047, 16'd32636, 16'd52138, 16'd32892, 16'd62382, 16'd11567, 16'd52440, 16'd40898, 16'd38236, 16'd60779, 16'd50423, 16'd17173});
	test_expansion(128'h5a74ea8846ab2ed5912b540accab7c4a, {16'd349, 16'd15281, 16'd6861, 16'd45829, 16'd35432, 16'd60440, 16'd19594, 16'd49512, 16'd25323, 16'd26841, 16'd2208, 16'd24925, 16'd49921, 16'd31664, 16'd24837, 16'd25614, 16'd46497, 16'd39072, 16'd42828, 16'd37194, 16'd57025, 16'd41898, 16'd26184, 16'd41820, 16'd36937, 16'd7063});
	test_expansion(128'h540f96a7de27b30b6fb58b1167e5256b, {16'd11030, 16'd21788, 16'd10967, 16'd36786, 16'd1984, 16'd10368, 16'd64404, 16'd2310, 16'd43009, 16'd28898, 16'd17376, 16'd33814, 16'd63060, 16'd35353, 16'd55528, 16'd33525, 16'd15254, 16'd13302, 16'd56739, 16'd14909, 16'd48749, 16'd55650, 16'd16676, 16'd4414, 16'd25401, 16'd7457});
	test_expansion(128'hc064f670e90d8113843e83821bcb9120, {16'd31622, 16'd40090, 16'd32418, 16'd64038, 16'd28971, 16'd19657, 16'd32719, 16'd4556, 16'd33066, 16'd53296, 16'd5977, 16'd20793, 16'd20814, 16'd34923, 16'd23798, 16'd45598, 16'd36200, 16'd37582, 16'd61725, 16'd16638, 16'd34553, 16'd15497, 16'd45758, 16'd4141, 16'd60659, 16'd37860});
	test_expansion(128'h48b92728bf55df067a04d8aba702f2b6, {16'd37477, 16'd62298, 16'd56298, 16'd25587, 16'd38020, 16'd41704, 16'd46150, 16'd3986, 16'd15184, 16'd4744, 16'd1794, 16'd60116, 16'd53598, 16'd50143, 16'd44768, 16'd21947, 16'd12030, 16'd8733, 16'd39687, 16'd22815, 16'd12281, 16'd3405, 16'd6611, 16'd3527, 16'd55287, 16'd18225});
	test_expansion(128'hc6f861f67a3cc8714c47ede0dbf4c115, {16'd29741, 16'd37474, 16'd15370, 16'd14615, 16'd18093, 16'd57956, 16'd10096, 16'd59219, 16'd43555, 16'd12753, 16'd39295, 16'd31254, 16'd33898, 16'd25253, 16'd10205, 16'd63750, 16'd41737, 16'd8589, 16'd29954, 16'd4963, 16'd22641, 16'd45239, 16'd40345, 16'd48405, 16'd38053, 16'd40480});
	test_expansion(128'h6e1512e1f0569dcf380b5960f45f8236, {16'd37380, 16'd38838, 16'd43455, 16'd22335, 16'd7453, 16'd49710, 16'd25041, 16'd1594, 16'd11038, 16'd36254, 16'd63664, 16'd27915, 16'd56836, 16'd32202, 16'd3421, 16'd53808, 16'd55496, 16'd46770, 16'd18379, 16'd64660, 16'd59178, 16'd28472, 16'd45359, 16'd4261, 16'd63064, 16'd939});
	test_expansion(128'h4afab593c6661470bc105799e3cdb457, {16'd20836, 16'd51048, 16'd45408, 16'd6890, 16'd37908, 16'd40517, 16'd61310, 16'd49744, 16'd27802, 16'd7574, 16'd50461, 16'd24333, 16'd62989, 16'd54938, 16'd54431, 16'd1814, 16'd39870, 16'd54157, 16'd47759, 16'd36827, 16'd46129, 16'd29155, 16'd31595, 16'd16960, 16'd45606, 16'd28260});
	test_expansion(128'h39a5a2b379fdffa800b584df06dc125c, {16'd33596, 16'd44905, 16'd40021, 16'd55875, 16'd27446, 16'd27967, 16'd59633, 16'd6546, 16'd63455, 16'd24255, 16'd6802, 16'd21526, 16'd19947, 16'd35626, 16'd39283, 16'd64813, 16'd46389, 16'd62879, 16'd28399, 16'd12188, 16'd38066, 16'd60278, 16'd43491, 16'd47509, 16'd9733, 16'd14104});
	test_expansion(128'h135183521e60b8a9a401f8d08609e3a3, {16'd37148, 16'd52274, 16'd1433, 16'd63797, 16'd26713, 16'd10437, 16'd1869, 16'd39622, 16'd58173, 16'd58142, 16'd10293, 16'd39669, 16'd17088, 16'd44612, 16'd37424, 16'd24686, 16'd34814, 16'd48040, 16'd29239, 16'd7817, 16'd40816, 16'd43846, 16'd61610, 16'd56168, 16'd38356, 16'd61121});
	test_expansion(128'he0b5a5531a1c28818890b35b15077181, {16'd53469, 16'd45645, 16'd29360, 16'd47540, 16'd45615, 16'd15879, 16'd19504, 16'd8203, 16'd44939, 16'd57432, 16'd63477, 16'd47986, 16'd8130, 16'd28682, 16'd9769, 16'd58635, 16'd38707, 16'd59042, 16'd24355, 16'd55932, 16'd38724, 16'd15125, 16'd27350, 16'd57443, 16'd14939, 16'd24166});
	test_expansion(128'hf339a7da70f2bdfcfbb0de48b0378b52, {16'd40853, 16'd19710, 16'd43837, 16'd43579, 16'd51607, 16'd675, 16'd46203, 16'd58089, 16'd55358, 16'd4386, 16'd64657, 16'd38215, 16'd9897, 16'd28604, 16'd52294, 16'd21205, 16'd51438, 16'd569, 16'd13165, 16'd47510, 16'd39836, 16'd37129, 16'd5780, 16'd37932, 16'd48299, 16'd1480});
	test_expansion(128'he690543103ad5648cddb41fb50feeaee, {16'd29021, 16'd60052, 16'd47930, 16'd25413, 16'd48316, 16'd40800, 16'd55222, 16'd8311, 16'd64123, 16'd31877, 16'd4321, 16'd5615, 16'd14424, 16'd12053, 16'd30444, 16'd58523, 16'd61845, 16'd58769, 16'd31114, 16'd42744, 16'd37768, 16'd3968, 16'd42245, 16'd32975, 16'd27185, 16'd52337});
	test_expansion(128'h8d4b42027e7e0a222b9e026c119e3340, {16'd54909, 16'd5546, 16'd46017, 16'd26258, 16'd61586, 16'd9837, 16'd9074, 16'd26649, 16'd62103, 16'd21851, 16'd21380, 16'd39113, 16'd37662, 16'd28318, 16'd26614, 16'd32905, 16'd12739, 16'd17019, 16'd44762, 16'd17576, 16'd40271, 16'd28860, 16'd30538, 16'd64268, 16'd8480, 16'd50183});
	test_expansion(128'h02f1870dc7f3bfd0d7cc59f0d2a71170, {16'd4065, 16'd624, 16'd40322, 16'd11582, 16'd51665, 16'd30485, 16'd53806, 16'd39836, 16'd2724, 16'd38506, 16'd35637, 16'd10104, 16'd26912, 16'd6118, 16'd14432, 16'd37706, 16'd44663, 16'd34090, 16'd36580, 16'd907, 16'd29884, 16'd25801, 16'd9971, 16'd2084, 16'd17819, 16'd6958});
	test_expansion(128'h04874564a854caa33534431ab26831b7, {16'd25371, 16'd38677, 16'd9581, 16'd59251, 16'd56297, 16'd18266, 16'd21091, 16'd20854, 16'd20763, 16'd50877, 16'd65101, 16'd40619, 16'd20834, 16'd55903, 16'd41252, 16'd19344, 16'd7438, 16'd22283, 16'd61792, 16'd6101, 16'd64287, 16'd20933, 16'd31687, 16'd40095, 16'd8189, 16'd5650});
	test_expansion(128'hb615a3ee2109ca31b776a43432f088fc, {16'd43462, 16'd62534, 16'd18832, 16'd24502, 16'd39427, 16'd50819, 16'd1787, 16'd24424, 16'd54185, 16'd28111, 16'd40924, 16'd57074, 16'd14828, 16'd17678, 16'd16382, 16'd9613, 16'd6185, 16'd63105, 16'd63494, 16'd57209, 16'd52502, 16'd45263, 16'd13103, 16'd20508, 16'd2884, 16'd51544});
	test_expansion(128'hb1fb84bd10fa9bf2bad26033ed259945, {16'd27239, 16'd19323, 16'd41686, 16'd39827, 16'd23631, 16'd26523, 16'd51814, 16'd17996, 16'd7793, 16'd5253, 16'd60743, 16'd30519, 16'd2633, 16'd34999, 16'd33359, 16'd9348, 16'd38739, 16'd28834, 16'd37269, 16'd10765, 16'd56789, 16'd58076, 16'd64029, 16'd22940, 16'd7414, 16'd11835});
	test_expansion(128'h1d1b498fb9fa3b6fd00a887da26bd059, {16'd20614, 16'd18563, 16'd14740, 16'd36689, 16'd15653, 16'd64535, 16'd9379, 16'd57843, 16'd64971, 16'd54924, 16'd19960, 16'd18377, 16'd12511, 16'd34626, 16'd17007, 16'd25706, 16'd35222, 16'd59253, 16'd2032, 16'd24715, 16'd22906, 16'd33506, 16'd57287, 16'd21359, 16'd54821, 16'd43568});
	test_expansion(128'h28ddd2fb883856a15a2b45263d14568c, {16'd3626, 16'd65331, 16'd29613, 16'd25382, 16'd53186, 16'd45012, 16'd24512, 16'd63972, 16'd901, 16'd22976, 16'd31739, 16'd42362, 16'd35629, 16'd39684, 16'd16476, 16'd17008, 16'd53992, 16'd8894, 16'd44299, 16'd19668, 16'd22347, 16'd10235, 16'd56330, 16'd47399, 16'd24162, 16'd11222});
	test_expansion(128'h7ca249bd09c4a5c14cbe732f266e689a, {16'd52755, 16'd28483, 16'd22490, 16'd25774, 16'd17498, 16'd49696, 16'd48614, 16'd26645, 16'd49766, 16'd46698, 16'd15742, 16'd25429, 16'd3074, 16'd20816, 16'd50687, 16'd29058, 16'd43849, 16'd48453, 16'd25775, 16'd51665, 16'd35124, 16'd27922, 16'd3940, 16'd46837, 16'd40076, 16'd24087});
	test_expansion(128'h802eab0715f31a959e3e21d9c4323877, {16'd18823, 16'd48145, 16'd54795, 16'd61122, 16'd47790, 16'd55125, 16'd23460, 16'd18894, 16'd14044, 16'd27516, 16'd25235, 16'd41154, 16'd41696, 16'd1086, 16'd16279, 16'd2242, 16'd53798, 16'd53922, 16'd55, 16'd62632, 16'd50087, 16'd30554, 16'd54170, 16'd3840, 16'd11950, 16'd11802});
	test_expansion(128'h7d6852de0f2a0d16443b959d4de0efce, {16'd10415, 16'd49300, 16'd3843, 16'd24647, 16'd63758, 16'd61444, 16'd34423, 16'd23447, 16'd53219, 16'd29136, 16'd12749, 16'd32288, 16'd28275, 16'd31204, 16'd40410, 16'd29029, 16'd32459, 16'd60395, 16'd37696, 16'd36422, 16'd3250, 16'd12457, 16'd57035, 16'd13894, 16'd1414, 16'd22677});
	test_expansion(128'hf5fccc03f9d51a4cd7f8a9b382f92613, {16'd12008, 16'd62694, 16'd54434, 16'd42433, 16'd24184, 16'd48108, 16'd50744, 16'd29697, 16'd32703, 16'd49906, 16'd52787, 16'd18031, 16'd44446, 16'd6346, 16'd34863, 16'd8335, 16'd62712, 16'd30311, 16'd31359, 16'd14570, 16'd38927, 16'd64774, 16'd13978, 16'd27627, 16'd16583, 16'd29929});
	test_expansion(128'h0f84585d22a0f869f5422c9cc71a1a7d, {16'd12756, 16'd36015, 16'd39487, 16'd10054, 16'd19206, 16'd9501, 16'd56255, 16'd23473, 16'd55392, 16'd46734, 16'd15037, 16'd53233, 16'd17502, 16'd18307, 16'd16700, 16'd20426, 16'd37512, 16'd9869, 16'd9091, 16'd61099, 16'd1810, 16'd37767, 16'd26528, 16'd39581, 16'd16459, 16'd43686});
	test_expansion(128'h6968ec78633cee690898a3be928f45a8, {16'd1341, 16'd39874, 16'd16172, 16'd36731, 16'd58023, 16'd56814, 16'd50309, 16'd54163, 16'd38371, 16'd49869, 16'd49659, 16'd8935, 16'd41679, 16'd16829, 16'd49734, 16'd34762, 16'd33420, 16'd16165, 16'd59637, 16'd42723, 16'd8168, 16'd30065, 16'd34775, 16'd52439, 16'd39908, 16'd37405});
	test_expansion(128'h28df47fdb2728cbd5dc084e36f3da59a, {16'd47761, 16'd11994, 16'd59580, 16'd49035, 16'd5708, 16'd6004, 16'd23144, 16'd54237, 16'd61379, 16'd45938, 16'd61430, 16'd51984, 16'd45614, 16'd8175, 16'd6955, 16'd17019, 16'd7856, 16'd32653, 16'd42423, 16'd1162, 16'd14118, 16'd31608, 16'd2834, 16'd62284, 16'd33845, 16'd21143});
	test_expansion(128'hd41547b5762f6f31e71b7258f2201a77, {16'd31224, 16'd61516, 16'd19340, 16'd63597, 16'd17266, 16'd36094, 16'd16931, 16'd20311, 16'd46631, 16'd31667, 16'd48766, 16'd50837, 16'd42427, 16'd18786, 16'd62750, 16'd60165, 16'd11011, 16'd62224, 16'd43589, 16'd46127, 16'd45058, 16'd112, 16'd42310, 16'd26091, 16'd4318, 16'd25814});
	test_expansion(128'hbc94bfb81df866078910fee23608499e, {16'd42523, 16'd56763, 16'd48244, 16'd27943, 16'd14643, 16'd37411, 16'd49227, 16'd3350, 16'd36669, 16'd23392, 16'd17972, 16'd63889, 16'd2725, 16'd10968, 16'd59632, 16'd17569, 16'd63234, 16'd8786, 16'd53775, 16'd25477, 16'd21275, 16'd25906, 16'd21873, 16'd42784, 16'd53805, 16'd21621});
	test_expansion(128'h216acbed9833c44ae5bebdc9d082737e, {16'd29889, 16'd60719, 16'd55477, 16'd37280, 16'd29426, 16'd65175, 16'd54415, 16'd64506, 16'd62869, 16'd57466, 16'd51553, 16'd57703, 16'd8659, 16'd56064, 16'd34996, 16'd56590, 16'd20635, 16'd57982, 16'd55999, 16'd26993, 16'd35643, 16'd53117, 16'd19184, 16'd51513, 16'd44007, 16'd2819});
	test_expansion(128'h1f27ec1a2da44599fbe5684cf48a0154, {16'd2600, 16'd18199, 16'd39694, 16'd34733, 16'd23728, 16'd42391, 16'd16920, 16'd47293, 16'd50395, 16'd33197, 16'd29831, 16'd42030, 16'd60118, 16'd55418, 16'd7498, 16'd17385, 16'd61404, 16'd19647, 16'd674, 16'd33563, 16'd53127, 16'd941, 16'd9771, 16'd65355, 16'd43141, 16'd29392});
	test_expansion(128'h93551d5815a189229c31985373b08c67, {16'd21593, 16'd40580, 16'd9722, 16'd25356, 16'd41521, 16'd54138, 16'd15719, 16'd26010, 16'd48766, 16'd38006, 16'd31531, 16'd20872, 16'd33280, 16'd53354, 16'd15191, 16'd47753, 16'd32475, 16'd5605, 16'd64271, 16'd45313, 16'd40457, 16'd11366, 16'd21550, 16'd2843, 16'd8197, 16'd38336});
	test_expansion(128'h88b613feeb283535cbb63f3e5fc76411, {16'd48539, 16'd15232, 16'd27442, 16'd26034, 16'd1193, 16'd59991, 16'd35898, 16'd24632, 16'd36727, 16'd18168, 16'd24790, 16'd34493, 16'd32031, 16'd50383, 16'd36625, 16'd48162, 16'd57019, 16'd59744, 16'd31243, 16'd36279, 16'd6488, 16'd20775, 16'd57093, 16'd8500, 16'd25245, 16'd37544});
	test_expansion(128'he142b55394c44aec3701c4fd5939b6c3, {16'd56289, 16'd43206, 16'd19361, 16'd36212, 16'd20365, 16'd2957, 16'd21478, 16'd5678, 16'd60487, 16'd32099, 16'd39458, 16'd47024, 16'd35410, 16'd61072, 16'd22754, 16'd31504, 16'd55295, 16'd15639, 16'd61218, 16'd26626, 16'd46340, 16'd25180, 16'd19216, 16'd30320, 16'd45373, 16'd26555});
	test_expansion(128'h91702eb1d71ea78a6be714efe8e6173e, {16'd4476, 16'd9000, 16'd43942, 16'd43106, 16'd59695, 16'd903, 16'd43033, 16'd59689, 16'd46918, 16'd28920, 16'd2532, 16'd29376, 16'd55525, 16'd17267, 16'd11308, 16'd61872, 16'd62346, 16'd23240, 16'd5000, 16'd62333, 16'd5735, 16'd51876, 16'd62367, 16'd62173, 16'd21039, 16'd53297});
	test_expansion(128'ha9ddd98684bd5960e65665986d0b58a3, {16'd58049, 16'd2112, 16'd2721, 16'd27697, 16'd30743, 16'd27664, 16'd23959, 16'd59224, 16'd27891, 16'd54359, 16'd55359, 16'd37984, 16'd44382, 16'd8659, 16'd47294, 16'd14957, 16'd27274, 16'd15489, 16'd23985, 16'd32067, 16'd44312, 16'd34165, 16'd58663, 16'd3215, 16'd10795, 16'd28204});
	test_expansion(128'h477cee36a5c391e8127835826b8f8bfb, {16'd59316, 16'd46109, 16'd41167, 16'd45903, 16'd39319, 16'd7955, 16'd52519, 16'd21529, 16'd29757, 16'd31009, 16'd43181, 16'd58923, 16'd37858, 16'd57826, 16'd54357, 16'd23172, 16'd13835, 16'd57676, 16'd17075, 16'd11495, 16'd57884, 16'd18016, 16'd17752, 16'd39505, 16'd73, 16'd24810});
	test_expansion(128'h55424015a04d9de0bf3f1ad1fbbb8ade, {16'd10320, 16'd33908, 16'd61291, 16'd24681, 16'd63079, 16'd6263, 16'd43220, 16'd34183, 16'd34448, 16'd6515, 16'd11452, 16'd53984, 16'd40159, 16'd50087, 16'd56094, 16'd35049, 16'd59484, 16'd58144, 16'd18376, 16'd65475, 16'd2669, 16'd43198, 16'd899, 16'd17222, 16'd57879, 16'd26972});
	test_expansion(128'h646be0a12c9ed8d4e05218fa3802ad3d, {16'd16203, 16'd9873, 16'd31502, 16'd28948, 16'd38188, 16'd45439, 16'd34226, 16'd39998, 16'd65360, 16'd51372, 16'd33041, 16'd30477, 16'd62896, 16'd17861, 16'd3851, 16'd38001, 16'd64059, 16'd60774, 16'd23220, 16'd44288, 16'd48162, 16'd36052, 16'd51386, 16'd11372, 16'd62377, 16'd39664});
	test_expansion(128'h13892e281eadbe5a16d118a4c58d5a19, {16'd43374, 16'd13312, 16'd4342, 16'd16505, 16'd61065, 16'd39392, 16'd29030, 16'd42769, 16'd30522, 16'd14902, 16'd16952, 16'd46390, 16'd33819, 16'd28985, 16'd43866, 16'd40125, 16'd34986, 16'd63851, 16'd10908, 16'd52710, 16'd6038, 16'd33084, 16'd60106, 16'd52375, 16'd22548, 16'd6303});
	test_expansion(128'h3175af73f8872d7f351bb17a3d956ff6, {16'd32994, 16'd36436, 16'd28132, 16'd53634, 16'd62945, 16'd28395, 16'd54910, 16'd29966, 16'd31904, 16'd28947, 16'd49727, 16'd14757, 16'd15025, 16'd53287, 16'd10846, 16'd16058, 16'd12496, 16'd29594, 16'd17008, 16'd38210, 16'd41211, 16'd42142, 16'd57382, 16'd39061, 16'd43565, 16'd5852});
	test_expansion(128'h967f1e38cdc177408ec3299ffd06b227, {16'd9598, 16'd56618, 16'd63106, 16'd24305, 16'd24357, 16'd58067, 16'd7076, 16'd31253, 16'd14091, 16'd32636, 16'd23870, 16'd30085, 16'd62965, 16'd12272, 16'd1750, 16'd46431, 16'd46507, 16'd64364, 16'd23642, 16'd37513, 16'd34100, 16'd12902, 16'd64453, 16'd56088, 16'd53867, 16'd39330});
	test_expansion(128'h2d560bef123a392059b1c80a953a7281, {16'd57355, 16'd23370, 16'd57799, 16'd7010, 16'd31466, 16'd49267, 16'd64900, 16'd17632, 16'd33802, 16'd8686, 16'd56009, 16'd16248, 16'd11163, 16'd12234, 16'd23271, 16'd40948, 16'd21747, 16'd6923, 16'd52382, 16'd49258, 16'd8281, 16'd55479, 16'd60054, 16'd36831, 16'd3108, 16'd27453});
	test_expansion(128'h0ed8937cf1c0763445be39286bddfaf2, {16'd47337, 16'd65413, 16'd1779, 16'd59359, 16'd36734, 16'd45681, 16'd45763, 16'd21341, 16'd41293, 16'd21093, 16'd35935, 16'd14453, 16'd1878, 16'd9802, 16'd11092, 16'd45218, 16'd16925, 16'd45987, 16'd4719, 16'd52363, 16'd10018, 16'd61482, 16'd43285, 16'd40794, 16'd63119, 16'd16463});
	test_expansion(128'hbea63b5e651d53ae1bce9205d7b4ea89, {16'd55742, 16'd26343, 16'd20146, 16'd40075, 16'd45660, 16'd23439, 16'd18019, 16'd47019, 16'd40539, 16'd13911, 16'd57882, 16'd21631, 16'd64874, 16'd60951, 16'd51498, 16'd21, 16'd40733, 16'd41233, 16'd48883, 16'd25521, 16'd40373, 16'd24604, 16'd60426, 16'd25737, 16'd19931, 16'd16777});
	test_expansion(128'hbb9fdbe100d4901b383ff5db6c016d94, {16'd16357, 16'd28761, 16'd58474, 16'd6414, 16'd60361, 16'd21936, 16'd5725, 16'd56423, 16'd64176, 16'd33264, 16'd37238, 16'd36668, 16'd52158, 16'd12174, 16'd52446, 16'd12785, 16'd58026, 16'd44377, 16'd28017, 16'd3712, 16'd49178, 16'd20370, 16'd53290, 16'd47693, 16'd34526, 16'd9090});
	test_expansion(128'h055efd618feac4ef227e6dc53aeb28cd, {16'd3140, 16'd3132, 16'd31805, 16'd41053, 16'd51973, 16'd55340, 16'd53633, 16'd33808, 16'd48881, 16'd22271, 16'd22209, 16'd18419, 16'd61712, 16'd54351, 16'd51109, 16'd18468, 16'd37781, 16'd24972, 16'd28783, 16'd50792, 16'd16149, 16'd34789, 16'd36326, 16'd56827, 16'd38806, 16'd42312});
	test_expansion(128'h990a11bbc019322d3b26d608f633d285, {16'd39030, 16'd63298, 16'd16445, 16'd41511, 16'd53399, 16'd17214, 16'd45088, 16'd23619, 16'd2898, 16'd58790, 16'd64359, 16'd19622, 16'd47543, 16'd9609, 16'd14952, 16'd56687, 16'd59179, 16'd54573, 16'd47024, 16'd39415, 16'd13669, 16'd56322, 16'd55789, 16'd61591, 16'd2311, 16'd35941});
	test_expansion(128'h44717de60bb3338f9fecae97854998c3, {16'd27527, 16'd35196, 16'd4770, 16'd15552, 16'd37779, 16'd57488, 16'd43601, 16'd51667, 16'd1290, 16'd53665, 16'd16598, 16'd16865, 16'd31798, 16'd50937, 16'd20845, 16'd63418, 16'd33119, 16'd33418, 16'd22231, 16'd3524, 16'd22236, 16'd19367, 16'd1753, 16'd49206, 16'd10898, 16'd42564});
	test_expansion(128'ha28c0db8d60769352442e88dff9a1dfd, {16'd55222, 16'd34645, 16'd4559, 16'd23860, 16'd62291, 16'd23760, 16'd7083, 16'd36066, 16'd64426, 16'd60851, 16'd45366, 16'd38209, 16'd61867, 16'd54699, 16'd49933, 16'd4886, 16'd40698, 16'd21484, 16'd30887, 16'd1570, 16'd6151, 16'd36515, 16'd34680, 16'd33987, 16'd7781, 16'd14631});
	test_expansion(128'h3dd18b7b5b1ebc8d9c7bc6c78ada3a32, {16'd36908, 16'd48418, 16'd53277, 16'd59962, 16'd61728, 16'd19307, 16'd4185, 16'd57806, 16'd56187, 16'd4257, 16'd37160, 16'd62479, 16'd51689, 16'd53825, 16'd47320, 16'd53489, 16'd174, 16'd34699, 16'd56685, 16'd21213, 16'd54117, 16'd46917, 16'd17258, 16'd18872, 16'd48495, 16'd2766});
	test_expansion(128'hd2c8adb0557ec983002a3ab7bf357e02, {16'd6250, 16'd55775, 16'd44820, 16'd48803, 16'd1842, 16'd40563, 16'd27130, 16'd30963, 16'd17082, 16'd7142, 16'd14846, 16'd23026, 16'd3395, 16'd40857, 16'd8760, 16'd45579, 16'd7614, 16'd1297, 16'd60653, 16'd60400, 16'd47416, 16'd64146, 16'd54000, 16'd60646, 16'd60022, 16'd9344});
	test_expansion(128'hf943f2cef9cc4c6282a6e831124700a4, {16'd12605, 16'd35471, 16'd23673, 16'd14999, 16'd29129, 16'd17813, 16'd61690, 16'd41054, 16'd61731, 16'd47467, 16'd42777, 16'd3563, 16'd53392, 16'd30536, 16'd15147, 16'd22435, 16'd24005, 16'd12641, 16'd64799, 16'd24486, 16'd57235, 16'd4845, 16'd5155, 16'd39075, 16'd20455, 16'd23555});
	test_expansion(128'hb3b3fd39ce17d843ec811937180354f2, {16'd9147, 16'd55001, 16'd56361, 16'd54946, 16'd27327, 16'd38894, 16'd48988, 16'd56683, 16'd6757, 16'd61070, 16'd10101, 16'd53963, 16'd1290, 16'd47183, 16'd13534, 16'd21249, 16'd14316, 16'd49051, 16'd63209, 16'd65310, 16'd44571, 16'd43251, 16'd40090, 16'd63284, 16'd5697, 16'd24571});
	test_expansion(128'h2cdb2630e63db9120965a8959aa1bad5, {16'd22572, 16'd13304, 16'd63517, 16'd13270, 16'd63776, 16'd15882, 16'd12064, 16'd28539, 16'd12648, 16'd40597, 16'd42594, 16'd64249, 16'd24978, 16'd21820, 16'd4073, 16'd52757, 16'd14723, 16'd52367, 16'd9401, 16'd62245, 16'd17459, 16'd2975, 16'd20094, 16'd13940, 16'd33510, 16'd42040});
	test_expansion(128'h660227a2f621fa4cf7b594998176c219, {16'd6369, 16'd20735, 16'd1008, 16'd582, 16'd57652, 16'd2642, 16'd22286, 16'd41358, 16'd1326, 16'd15404, 16'd49435, 16'd22797, 16'd61254, 16'd56521, 16'd10827, 16'd22791, 16'd20558, 16'd28230, 16'd21719, 16'd46151, 16'd6011, 16'd47769, 16'd30033, 16'd49668, 16'd11953, 16'd49443});
	test_expansion(128'h2afe500c0b1816b24bf5e3138d035afc, {16'd14822, 16'd60622, 16'd59401, 16'd64654, 16'd55452, 16'd37010, 16'd32290, 16'd47554, 16'd40226, 16'd19073, 16'd27304, 16'd11816, 16'd64943, 16'd6829, 16'd63508, 16'd28701, 16'd3347, 16'd44819, 16'd24057, 16'd38846, 16'd29547, 16'd14788, 16'd65477, 16'd56345, 16'd1985, 16'd46506});
	test_expansion(128'h8438e46dcd300b2843c03bc80a8b3b3e, {16'd64431, 16'd60978, 16'd18524, 16'd13921, 16'd48016, 16'd61271, 16'd58750, 16'd9531, 16'd58669, 16'd54509, 16'd51347, 16'd33603, 16'd19410, 16'd15990, 16'd62191, 16'd47799, 16'd15469, 16'd31043, 16'd22230, 16'd61692, 16'd19785, 16'd18531, 16'd16745, 16'd3172, 16'd59723, 16'd55082});
	test_expansion(128'h9852be3517d1be2292adf407bef645a9, {16'd33752, 16'd333, 16'd38437, 16'd10773, 16'd35137, 16'd62841, 16'd43882, 16'd39493, 16'd20249, 16'd35902, 16'd18661, 16'd64515, 16'd47820, 16'd59148, 16'd44664, 16'd17285, 16'd43686, 16'd52237, 16'd7680, 16'd60731, 16'd11018, 16'd28892, 16'd54454, 16'd55920, 16'd16561, 16'd47476});
	test_expansion(128'h009b1b441c4269ff8eacfd5fc6329803, {16'd50335, 16'd20768, 16'd44290, 16'd36677, 16'd4732, 16'd21691, 16'd10028, 16'd46724, 16'd17735, 16'd18769, 16'd27893, 16'd18943, 16'd35568, 16'd5753, 16'd37272, 16'd56354, 16'd59641, 16'd57453, 16'd61781, 16'd45130, 16'd47320, 16'd4944, 16'd62456, 16'd16626, 16'd40375, 16'd45309});
	test_expansion(128'h689ba289a17d130ad847934cb5e326fe, {16'd35670, 16'd10437, 16'd39, 16'd51237, 16'd59096, 16'd4022, 16'd46072, 16'd521, 16'd54456, 16'd30863, 16'd51769, 16'd9391, 16'd40795, 16'd6139, 16'd51385, 16'd63675, 16'd46703, 16'd18269, 16'd9432, 16'd26932, 16'd52348, 16'd65172, 16'd57221, 16'd41859, 16'd15852, 16'd63037});
	test_expansion(128'hdee0ec32272985c1a3d0ebb07d232c02, {16'd52043, 16'd62082, 16'd7490, 16'd14369, 16'd53642, 16'd59354, 16'd10281, 16'd33196, 16'd45503, 16'd31546, 16'd39566, 16'd25047, 16'd59513, 16'd6060, 16'd26864, 16'd16, 16'd14514, 16'd53039, 16'd42566, 16'd45354, 16'd49513, 16'd12796, 16'd34697, 16'd14313, 16'd1756, 16'd27740});
	test_expansion(128'hafd08577d97a7c8f75bcebf4f790a1cb, {16'd43694, 16'd33786, 16'd46358, 16'd36215, 16'd7429, 16'd9675, 16'd29324, 16'd54219, 16'd33008, 16'd41229, 16'd31767, 16'd33127, 16'd43907, 16'd48670, 16'd33978, 16'd25108, 16'd8504, 16'd40782, 16'd52352, 16'd25954, 16'd60864, 16'd18667, 16'd30433, 16'd55927, 16'd16881, 16'd59839});
	test_expansion(128'h95a112fef4e6a6140e9d49f2d3ca07dd, {16'd60256, 16'd34564, 16'd3984, 16'd63044, 16'd20264, 16'd54061, 16'd6421, 16'd24830, 16'd18726, 16'd5425, 16'd8413, 16'd37073, 16'd44337, 16'd56971, 16'd38217, 16'd37415, 16'd41710, 16'd10777, 16'd51188, 16'd58183, 16'd31342, 16'd56394, 16'd6075, 16'd43363, 16'd1643, 16'd27759});
	test_expansion(128'h8eb6ccbb02da80c5a81c74171f9507f5, {16'd48895, 16'd41891, 16'd60275, 16'd46716, 16'd2449, 16'd24136, 16'd44083, 16'd31900, 16'd53775, 16'd59785, 16'd27780, 16'd23825, 16'd32195, 16'd37782, 16'd43888, 16'd44010, 16'd16212, 16'd28376, 16'd48774, 16'd41694, 16'd7817, 16'd54808, 16'd30401, 16'd50958, 16'd55512, 16'd43843});
	test_expansion(128'h3be5419a19495fb54ec25548e4ed9116, {16'd32122, 16'd26164, 16'd8929, 16'd7685, 16'd32336, 16'd42267, 16'd966, 16'd4144, 16'd515, 16'd39903, 16'd37955, 16'd7405, 16'd19765, 16'd3323, 16'd18721, 16'd61006, 16'd18835, 16'd34153, 16'd17295, 16'd6595, 16'd43203, 16'd29129, 16'd24749, 16'd10458, 16'd60745, 16'd47557});
	test_expansion(128'h02e1967f8ec3991ccb5c07ff970ccf85, {16'd16275, 16'd36033, 16'd56379, 16'd36740, 16'd49443, 16'd43274, 16'd37414, 16'd39352, 16'd29839, 16'd51573, 16'd49458, 16'd20211, 16'd895, 16'd17809, 16'd61528, 16'd55319, 16'd5181, 16'd43380, 16'd44133, 16'd46362, 16'd53005, 16'd53637, 16'd22643, 16'd31633, 16'd53986, 16'd27902});
	test_expansion(128'h9fb08d91b753bca320bca03b218c2f16, {16'd45496, 16'd6577, 16'd14478, 16'd14572, 16'd54440, 16'd27686, 16'd41601, 16'd38088, 16'd4554, 16'd65239, 16'd43859, 16'd13227, 16'd64908, 16'd65530, 16'd36429, 16'd60717, 16'd63454, 16'd54036, 16'd52547, 16'd5010, 16'd7832, 16'd4842, 16'd63866, 16'd47641, 16'd53349, 16'd39634});
	test_expansion(128'h2ff452425b07ab16671e64578504cd61, {16'd45140, 16'd64, 16'd46370, 16'd59208, 16'd55189, 16'd2262, 16'd51334, 16'd28146, 16'd51211, 16'd26000, 16'd49491, 16'd31355, 16'd58885, 16'd34270, 16'd29638, 16'd41450, 16'd45383, 16'd31989, 16'd14600, 16'd32455, 16'd49024, 16'd23080, 16'd47279, 16'd43211, 16'd16883, 16'd62395});
	test_expansion(128'h7293d7d43833485b0fb212c2ad31e9ea, {16'd28779, 16'd22725, 16'd3919, 16'd24151, 16'd39944, 16'd3441, 16'd61673, 16'd53705, 16'd23234, 16'd22960, 16'd64005, 16'd61123, 16'd7346, 16'd41747, 16'd15705, 16'd30706, 16'd48542, 16'd59510, 16'd43366, 16'd16775, 16'd29854, 16'd25883, 16'd62116, 16'd61026, 16'd22420, 16'd14960});
	test_expansion(128'h1bb3c9c6402b48829a477e03da6e71e9, {16'd21932, 16'd52082, 16'd14376, 16'd57864, 16'd11229, 16'd386, 16'd13538, 16'd10167, 16'd12428, 16'd157, 16'd35929, 16'd18349, 16'd24951, 16'd11723, 16'd27360, 16'd36037, 16'd47976, 16'd2880, 16'd25775, 16'd670, 16'd2657, 16'd41101, 16'd14885, 16'd39096, 16'd32339, 16'd57790});
	test_expansion(128'h588ad03f8d7276aefb5e91298682bf97, {16'd6075, 16'd49293, 16'd2743, 16'd58541, 16'd6830, 16'd14112, 16'd42122, 16'd26203, 16'd44308, 16'd52394, 16'd39021, 16'd27657, 16'd61229, 16'd38311, 16'd23323, 16'd38471, 16'd12027, 16'd51368, 16'd516, 16'd42201, 16'd1225, 16'd46310, 16'd64538, 16'd20243, 16'd34629, 16'd50544});
	test_expansion(128'hfe6905ed15af5b1567ffe576770dc67b, {16'd59654, 16'd26087, 16'd44483, 16'd38580, 16'd10024, 16'd65248, 16'd54223, 16'd25537, 16'd13579, 16'd18016, 16'd18248, 16'd1060, 16'd45952, 16'd24291, 16'd51975, 16'd55661, 16'd64704, 16'd9456, 16'd8969, 16'd40950, 16'd33411, 16'd15435, 16'd30834, 16'd17926, 16'd49352, 16'd28844});
	test_expansion(128'h9c2826d8969b8c2436989655b760d614, {16'd1195, 16'd24899, 16'd52847, 16'd23890, 16'd727, 16'd63990, 16'd8774, 16'd55897, 16'd48646, 16'd56793, 16'd43973, 16'd25032, 16'd33653, 16'd26899, 16'd23422, 16'd5681, 16'd40905, 16'd42310, 16'd61652, 16'd44912, 16'd59012, 16'd47158, 16'd32828, 16'd25090, 16'd7720, 16'd6896});
	test_expansion(128'hebf3ec09de1f20543e3469d7cbeb3b17, {16'd50926, 16'd16582, 16'd30018, 16'd10838, 16'd48874, 16'd54509, 16'd22499, 16'd52901, 16'd13657, 16'd48832, 16'd10731, 16'd61153, 16'd61914, 16'd24287, 16'd59989, 16'd41730, 16'd32491, 16'd16944, 16'd6723, 16'd63666, 16'd58130, 16'd52706, 16'd19666, 16'd50345, 16'd31485, 16'd13069});
	test_expansion(128'hb075bbf7f8c555b0d41f99b18336a5a8, {16'd46285, 16'd31061, 16'd53653, 16'd43595, 16'd39406, 16'd6231, 16'd33636, 16'd63985, 16'd46965, 16'd5633, 16'd43663, 16'd23118, 16'd36844, 16'd48229, 16'd7884, 16'd41426, 16'd52363, 16'd31294, 16'd52619, 16'd14174, 16'd64984, 16'd26340, 16'd2650, 16'd24547, 16'd9399, 16'd24907});
	test_expansion(128'h0fa16fa28df765fc957bebea483a2c2a, {16'd33031, 16'd40722, 16'd57413, 16'd31605, 16'd11989, 16'd22254, 16'd60862, 16'd3756, 16'd48701, 16'd62075, 16'd21976, 16'd30136, 16'd10465, 16'd43376, 16'd38429, 16'd7059, 16'd58800, 16'd62636, 16'd53538, 16'd47263, 16'd46059, 16'd20008, 16'd4318, 16'd14877, 16'd12650, 16'd35099});
	test_expansion(128'hdb841b45834971398c8147f6a2144dd4, {16'd34274, 16'd21788, 16'd13067, 16'd63709, 16'd51057, 16'd49015, 16'd14459, 16'd15021, 16'd25229, 16'd10272, 16'd44478, 16'd45359, 16'd56474, 16'd57699, 16'd4446, 16'd50561, 16'd54770, 16'd22427, 16'd65212, 16'd46062, 16'd18790, 16'd11117, 16'd59599, 16'd26450, 16'd46509, 16'd24639});
	test_expansion(128'h98521dabb6167741e128f904f4c5e750, {16'd25392, 16'd44615, 16'd33629, 16'd54074, 16'd18921, 16'd23000, 16'd39257, 16'd34195, 16'd45421, 16'd2423, 16'd45599, 16'd44108, 16'd29500, 16'd56374, 16'd28518, 16'd16752, 16'd21256, 16'd31697, 16'd1379, 16'd5890, 16'd24792, 16'd62447, 16'd33525, 16'd41624, 16'd2224, 16'd19470});
	test_expansion(128'ha1562235a82616f351576d19cdfa0bb1, {16'd11593, 16'd13450, 16'd53578, 16'd30241, 16'd52032, 16'd15932, 16'd55020, 16'd14757, 16'd33200, 16'd36899, 16'd27047, 16'd5536, 16'd35524, 16'd8083, 16'd17520, 16'd64668, 16'd64331, 16'd58648, 16'd28448, 16'd25037, 16'd1172, 16'd19764, 16'd14467, 16'd64507, 16'd39282, 16'd21312});
	test_expansion(128'hd757906df603dd4c870746e32abd9ef2, {16'd19723, 16'd10032, 16'd18449, 16'd6389, 16'd33253, 16'd21186, 16'd30995, 16'd50226, 16'd42524, 16'd46177, 16'd50584, 16'd62561, 16'd23318, 16'd29490, 16'd17305, 16'd3269, 16'd27115, 16'd39363, 16'd59726, 16'd25772, 16'd57198, 16'd59357, 16'd56282, 16'd236, 16'd5019, 16'd64879});
	test_expansion(128'hab471a5633693bd7e3b705e3905df164, {16'd4237, 16'd62927, 16'd32891, 16'd32595, 16'd24946, 16'd25336, 16'd49949, 16'd56936, 16'd1782, 16'd4530, 16'd32170, 16'd15315, 16'd59515, 16'd30957, 16'd57753, 16'd51935, 16'd51919, 16'd2130, 16'd28418, 16'd31519, 16'd16343, 16'd22529, 16'd1914, 16'd24025, 16'd52418, 16'd34322});
	test_expansion(128'hab982282ab82c41513d6e6d238fb7c54, {16'd19239, 16'd53482, 16'd56364, 16'd32592, 16'd61905, 16'd41019, 16'd61717, 16'd47090, 16'd1734, 16'd64900, 16'd65533, 16'd44977, 16'd29350, 16'd812, 16'd45633, 16'd33658, 16'd17631, 16'd55961, 16'd64243, 16'd48386, 16'd8793, 16'd18094, 16'd21453, 16'd29292, 16'd63390, 16'd57310});
	test_expansion(128'hc2968474d1bd1f9db607f5c5a0276a58, {16'd33129, 16'd57521, 16'd48318, 16'd20085, 16'd43901, 16'd14855, 16'd58690, 16'd19969, 16'd13015, 16'd31982, 16'd50131, 16'd41159, 16'd65411, 16'd58331, 16'd46597, 16'd30460, 16'd33386, 16'd57546, 16'd24740, 16'd2296, 16'd31269, 16'd23683, 16'd35947, 16'd19277, 16'd34775, 16'd48418});
	test_expansion(128'h0c51f78358be00e8f80f37b9585ffdc6, {16'd9749, 16'd11743, 16'd59278, 16'd32594, 16'd53671, 16'd2606, 16'd15858, 16'd53971, 16'd65336, 16'd54581, 16'd32801, 16'd52249, 16'd45053, 16'd60385, 16'd54382, 16'd3726, 16'd36652, 16'd47790, 16'd23772, 16'd15191, 16'd29784, 16'd46341, 16'd19839, 16'd24374, 16'd24657, 16'd10671});
	test_expansion(128'h421b87d1300d2bb54f230e618a0e137b, {16'd59187, 16'd32714, 16'd10425, 16'd56681, 16'd54854, 16'd5702, 16'd28344, 16'd56687, 16'd35649, 16'd36152, 16'd52054, 16'd10873, 16'd38256, 16'd22120, 16'd3129, 16'd10043, 16'd58099, 16'd9377, 16'd2684, 16'd8077, 16'd46606, 16'd40434, 16'd50543, 16'd25381, 16'd51815, 16'd150});
	test_expansion(128'hf697db70e64e2780df82cac21ee1f6ea, {16'd56066, 16'd8801, 16'd25157, 16'd2905, 16'd29069, 16'd54147, 16'd30063, 16'd29660, 16'd22000, 16'd50201, 16'd24564, 16'd2885, 16'd40188, 16'd49770, 16'd13059, 16'd48082, 16'd32570, 16'd62648, 16'd16807, 16'd13212, 16'd18500, 16'd39832, 16'd37355, 16'd62728, 16'd44817, 16'd29393});
	test_expansion(128'h9f110af37724df5144275a639e68afeb, {16'd61185, 16'd47477, 16'd21991, 16'd33492, 16'd44265, 16'd42590, 16'd43398, 16'd1322, 16'd25543, 16'd54358, 16'd54238, 16'd55966, 16'd49469, 16'd47784, 16'd35087, 16'd62643, 16'd20017, 16'd62448, 16'd25853, 16'd44287, 16'd22056, 16'd35668, 16'd18137, 16'd43824, 16'd3132, 16'd61371});
	test_expansion(128'hc3c4b4a354483928eba5056a6f5c7d2b, {16'd42947, 16'd47657, 16'd19975, 16'd34893, 16'd8063, 16'd51689, 16'd46058, 16'd55678, 16'd22173, 16'd63723, 16'd25279, 16'd49901, 16'd21882, 16'd33348, 16'd30407, 16'd58420, 16'd49380, 16'd55735, 16'd28005, 16'd6687, 16'd47349, 16'd2131, 16'd53714, 16'd5753, 16'd1546, 16'd58932});
	test_expansion(128'h7f37305e48c689e9527e7df71cddb81d, {16'd43230, 16'd15555, 16'd30232, 16'd27354, 16'd56825, 16'd48424, 16'd40637, 16'd7691, 16'd33934, 16'd9767, 16'd13288, 16'd19117, 16'd41838, 16'd21275, 16'd44522, 16'd55408, 16'd18356, 16'd30135, 16'd5544, 16'd28537, 16'd29462, 16'd10965, 16'd62404, 16'd40774, 16'd34138, 16'd37620});
	test_expansion(128'hc68780d75fc89d08951fb01cddf79e87, {16'd2661, 16'd22184, 16'd14850, 16'd58139, 16'd12291, 16'd6660, 16'd43766, 16'd51223, 16'd20715, 16'd16820, 16'd34233, 16'd15798, 16'd55735, 16'd15001, 16'd1914, 16'd40726, 16'd59678, 16'd9826, 16'd13696, 16'd8931, 16'd37677, 16'd17575, 16'd8201, 16'd35664, 16'd56701, 16'd56979});
	test_expansion(128'hf114dccc487e10487ad72e01831f2aac, {16'd14509, 16'd30946, 16'd29350, 16'd50093, 16'd7759, 16'd6541, 16'd18343, 16'd27335, 16'd13248, 16'd63215, 16'd60202, 16'd37002, 16'd10654, 16'd21009, 16'd24151, 16'd52179, 16'd43570, 16'd21066, 16'd42298, 16'd19268, 16'd63769, 16'd24706, 16'd16993, 16'd16984, 16'd57219, 16'd280});
	test_expansion(128'h4648cd29e87dd3618247feaac4bd0d82, {16'd21703, 16'd45068, 16'd38070, 16'd20183, 16'd4447, 16'd34134, 16'd12017, 16'd26692, 16'd26448, 16'd8345, 16'd63789, 16'd43936, 16'd29767, 16'd10373, 16'd35789, 16'd50100, 16'd4588, 16'd21627, 16'd37256, 16'd16482, 16'd22056, 16'd53908, 16'd10853, 16'd5534, 16'd61717, 16'd6246});
	test_expansion(128'hc1a636a0787f20d14e241b41779c9497, {16'd16954, 16'd34351, 16'd10449, 16'd51325, 16'd50351, 16'd61367, 16'd53771, 16'd2612, 16'd9969, 16'd43366, 16'd7843, 16'd11928, 16'd46686, 16'd44354, 16'd59125, 16'd26105, 16'd27381, 16'd57693, 16'd46189, 16'd46540, 16'd58307, 16'd9181, 16'd62153, 16'd58409, 16'd26868, 16'd26756});
	test_expansion(128'he7b4915a25ef04b8f630d539ad562fa1, {16'd55302, 16'd40383, 16'd4538, 16'd35505, 16'd27058, 16'd46498, 16'd9346, 16'd20021, 16'd17486, 16'd38616, 16'd60861, 16'd34071, 16'd53735, 16'd25284, 16'd35358, 16'd16017, 16'd48452, 16'd46813, 16'd19068, 16'd58645, 16'd48775, 16'd22483, 16'd35268, 16'd64783, 16'd62347, 16'd35940});
	test_expansion(128'h271ab6e4a4abf4a32cac094f2ba06c8e, {16'd52775, 16'd6733, 16'd8179, 16'd2605, 16'd37738, 16'd46609, 16'd59456, 16'd38975, 16'd3106, 16'd45222, 16'd55019, 16'd57339, 16'd18650, 16'd62302, 16'd38117, 16'd60545, 16'd22320, 16'd7285, 16'd60457, 16'd11152, 16'd46135, 16'd49967, 16'd61543, 16'd14138, 16'd27772, 16'd36766});
	test_expansion(128'ha92e2e585e46bf5d463038de60113749, {16'd10955, 16'd1369, 16'd25481, 16'd8613, 16'd28548, 16'd10913, 16'd29807, 16'd17300, 16'd7563, 16'd43041, 16'd23094, 16'd46532, 16'd9310, 16'd42404, 16'd2821, 16'd7853, 16'd56563, 16'd35366, 16'd46537, 16'd46690, 16'd21347, 16'd29666, 16'd2233, 16'd15417, 16'd64465, 16'd36349});
	test_expansion(128'h16fb711fc9a652ad36815058f926b99e, {16'd62251, 16'd39627, 16'd19336, 16'd64673, 16'd34148, 16'd59404, 16'd2082, 16'd21372, 16'd18114, 16'd58555, 16'd46329, 16'd43292, 16'd16043, 16'd22416, 16'd35531, 16'd15348, 16'd19726, 16'd57631, 16'd62297, 16'd6613, 16'd12005, 16'd35706, 16'd8059, 16'd27716, 16'd39145, 16'd52865});
	test_expansion(128'hf9cb24cf8d9b406b3a3388c5cb76ba70, {16'd46861, 16'd42388, 16'd55598, 16'd50242, 16'd63287, 16'd742, 16'd64600, 16'd55056, 16'd44480, 16'd40912, 16'd54245, 16'd60427, 16'd64115, 16'd12793, 16'd52517, 16'd60918, 16'd55602, 16'd7609, 16'd45962, 16'd35451, 16'd25593, 16'd35468, 16'd49325, 16'd12206, 16'd21499, 16'd38735});
	test_expansion(128'h2d6c0ee6be2f97c07c1e3bdad6f49923, {16'd35070, 16'd46042, 16'd23413, 16'd33168, 16'd46122, 16'd11731, 16'd52655, 16'd28699, 16'd50404, 16'd30223, 16'd27656, 16'd23970, 16'd28041, 16'd61607, 16'd4720, 16'd62562, 16'd23291, 16'd16037, 16'd28206, 16'd11820, 16'd58789, 16'd21244, 16'd58008, 16'd17082, 16'd55379, 16'd44272});
	test_expansion(128'h032a06990cb4b60d1431c1d78b1dce08, {16'd58164, 16'd59088, 16'd37869, 16'd10502, 16'd32254, 16'd34949, 16'd34914, 16'd62417, 16'd1818, 16'd48366, 16'd5362, 16'd63300, 16'd39548, 16'd29199, 16'd61089, 16'd41396, 16'd227, 16'd5099, 16'd39312, 16'd21773, 16'd4085, 16'd25532, 16'd33926, 16'd52962, 16'd5686, 16'd38155});
	test_expansion(128'he0c9d9437943a29b098cbe59bd21e861, {16'd4966, 16'd6080, 16'd18236, 16'd5694, 16'd11286, 16'd44893, 16'd7220, 16'd28839, 16'd22777, 16'd63064, 16'd1213, 16'd13111, 16'd33783, 16'd14119, 16'd44443, 16'd41747, 16'd7537, 16'd55550, 16'd59340, 16'd5498, 16'd30105, 16'd9120, 16'd64730, 16'd26929, 16'd25142, 16'd9376});
	test_expansion(128'h1ec4dabe865bfb0387a96bed7a786f13, {16'd22546, 16'd37932, 16'd15339, 16'd45907, 16'd58056, 16'd14571, 16'd39509, 16'd26986, 16'd39137, 16'd38578, 16'd14330, 16'd12646, 16'd58236, 16'd53335, 16'd6355, 16'd19746, 16'd4279, 16'd43975, 16'd16015, 16'd31594, 16'd22945, 16'd13646, 16'd40298, 16'd17392, 16'd30654, 16'd43902});
	test_expansion(128'h1c3832ceb7575a71189e162ac6a1e358, {16'd55927, 16'd58894, 16'd43281, 16'd52433, 16'd50714, 16'd15617, 16'd38195, 16'd36032, 16'd9734, 16'd47186, 16'd43489, 16'd13670, 16'd43414, 16'd7342, 16'd31277, 16'd44494, 16'd10415, 16'd50113, 16'd53191, 16'd35392, 16'd8448, 16'd19751, 16'd2525, 16'd45944, 16'd37918, 16'd38856});
	test_expansion(128'hb925360a6fb50ac1837bbf8a9646cb8c, {16'd43167, 16'd26288, 16'd6862, 16'd18441, 16'd50928, 16'd57503, 16'd20222, 16'd34743, 16'd20244, 16'd3932, 16'd42661, 16'd53404, 16'd54644, 16'd5708, 16'd42600, 16'd17270, 16'd53810, 16'd6513, 16'd36459, 16'd64865, 16'd3083, 16'd21700, 16'd18106, 16'd17313, 16'd64917, 16'd53974});
	test_expansion(128'hd26072ffd2094d58d5215714ea5585f5, {16'd50418, 16'd29669, 16'd13551, 16'd27157, 16'd42022, 16'd56498, 16'd28156, 16'd56180, 16'd25150, 16'd52005, 16'd56337, 16'd21527, 16'd56945, 16'd22733, 16'd32479, 16'd14016, 16'd45168, 16'd14697, 16'd57660, 16'd23929, 16'd64223, 16'd1991, 16'd50883, 16'd26031, 16'd49527, 16'd27294});
	test_expansion(128'h5157baf22b40e8993f6323cd197d01c1, {16'd62317, 16'd20889, 16'd62044, 16'd58373, 16'd6263, 16'd40058, 16'd34271, 16'd22254, 16'd37324, 16'd39023, 16'd49726, 16'd14179, 16'd7040, 16'd56524, 16'd27385, 16'd51875, 16'd42244, 16'd14912, 16'd64515, 16'd53860, 16'd57198, 16'd53847, 16'd59950, 16'd62477, 16'd56249, 16'd32713});
	test_expansion(128'h2af2a5e07ec0bc7e0dd7606957e63ad4, {16'd56291, 16'd25694, 16'd22947, 16'd55174, 16'd33223, 16'd23485, 16'd24682, 16'd64975, 16'd29068, 16'd55521, 16'd46164, 16'd59816, 16'd35540, 16'd29903, 16'd46570, 16'd33625, 16'd63104, 16'd8413, 16'd31890, 16'd4690, 16'd30897, 16'd35542, 16'd9109, 16'd1332, 16'd27427, 16'd44992});
	test_expansion(128'hbe624127449ea7b1e4f9a5797b9836cc, {16'd46182, 16'd64373, 16'd17864, 16'd45990, 16'd36333, 16'd51858, 16'd65519, 16'd41735, 16'd64004, 16'd44633, 16'd53583, 16'd62371, 16'd4942, 16'd19319, 16'd24972, 16'd60211, 16'd56807, 16'd23981, 16'd51988, 16'd53121, 16'd31226, 16'd29688, 16'd6902, 16'd43202, 16'd17441, 16'd6000});
	test_expansion(128'ha9af5888adef7f0821f9aacfdeeb493b, {16'd42928, 16'd45604, 16'd6511, 16'd7922, 16'd36586, 16'd3701, 16'd22646, 16'd15328, 16'd523, 16'd31797, 16'd48862, 16'd17227, 16'd1796, 16'd49228, 16'd38910, 16'd57755, 16'd46973, 16'd16056, 16'd31121, 16'd44574, 16'd10974, 16'd26492, 16'd65038, 16'd38512, 16'd32311, 16'd19956});
	test_expansion(128'h8b8eca746f4c63d56763a605a199292c, {16'd59737, 16'd36631, 16'd4176, 16'd44172, 16'd34918, 16'd45828, 16'd42850, 16'd19646, 16'd19262, 16'd49399, 16'd16636, 16'd49192, 16'd43467, 16'd3727, 16'd62716, 16'd698, 16'd22564, 16'd62695, 16'd37326, 16'd51898, 16'd58242, 16'd12589, 16'd37885, 16'd1200, 16'd54525, 16'd23857});
	test_expansion(128'h9f92ad758770ac803c8dd39471cc4cc0, {16'd29176, 16'd5257, 16'd42660, 16'd54804, 16'd7222, 16'd33181, 16'd63022, 16'd35645, 16'd4294, 16'd33472, 16'd26409, 16'd50427, 16'd60686, 16'd21368, 16'd59140, 16'd64389, 16'd62527, 16'd1767, 16'd15448, 16'd4974, 16'd42909, 16'd24350, 16'd55059, 16'd15817, 16'd54630, 16'd1934});
	test_expansion(128'h21586257db1621a6308a8851af886f29, {16'd14269, 16'd31953, 16'd59419, 16'd58188, 16'd13358, 16'd37438, 16'd26167, 16'd31790, 16'd24034, 16'd59100, 16'd30042, 16'd17107, 16'd14570, 16'd27732, 16'd23142, 16'd37159, 16'd9636, 16'd62736, 16'd15458, 16'd17132, 16'd1692, 16'd843, 16'd11139, 16'd16348, 16'd62976, 16'd62362});
	test_expansion(128'h6fd07de1232ea19b17f834d8d8b121c9, {16'd52961, 16'd15301, 16'd64413, 16'd15821, 16'd49123, 16'd53994, 16'd63042, 16'd37821, 16'd50469, 16'd27565, 16'd19328, 16'd22095, 16'd3851, 16'd10104, 16'd13599, 16'd24438, 16'd41993, 16'd33566, 16'd20346, 16'd45619, 16'd3628, 16'd24284, 16'd63024, 16'd65376, 16'd7764, 16'd35711});
	test_expansion(128'h60127a70112249cae1c71b21bfd1ce28, {16'd33871, 16'd49708, 16'd62466, 16'd18369, 16'd17243, 16'd42915, 16'd21180, 16'd48126, 16'd31142, 16'd17920, 16'd59235, 16'd43036, 16'd59996, 16'd22200, 16'd19917, 16'd25173, 16'd9761, 16'd1865, 16'd65272, 16'd11893, 16'd16985, 16'd1680, 16'd41115, 16'd42945, 16'd26317, 16'd30667});
	test_expansion(128'ha8601ae27d05b96f52b88798972a4790, {16'd4189, 16'd33028, 16'd51663, 16'd22219, 16'd51048, 16'd24334, 16'd42155, 16'd56296, 16'd43151, 16'd49684, 16'd10727, 16'd16740, 16'd54010, 16'd47431, 16'd11933, 16'd45343, 16'd1880, 16'd6002, 16'd32151, 16'd1458, 16'd31908, 16'd27787, 16'd25265, 16'd33962, 16'd4280, 16'd28263});
	test_expansion(128'h371de0a06dde05f1decca262a672f42d, {16'd15640, 16'd44409, 16'd50204, 16'd64246, 16'd8413, 16'd26097, 16'd53289, 16'd42747, 16'd57179, 16'd12990, 16'd39214, 16'd26843, 16'd158, 16'd2766, 16'd32119, 16'd65052, 16'd19973, 16'd15926, 16'd65317, 16'd58939, 16'd54066, 16'd39541, 16'd44077, 16'd4895, 16'd61010, 16'd64671});
	test_expansion(128'ha22a0c79d3ebd00b65cca6dc7be85508, {16'd21150, 16'd53473, 16'd56395, 16'd45755, 16'd2896, 16'd36292, 16'd7251, 16'd44439, 16'd56130, 16'd17108, 16'd63269, 16'd54640, 16'd60523, 16'd53191, 16'd46457, 16'd11923, 16'd55973, 16'd26768, 16'd53995, 16'd37569, 16'd50062, 16'd41437, 16'd36504, 16'd34117, 16'd10096, 16'd40763});
	test_expansion(128'h7bb684e2b3a76ea31315bc2014017899, {16'd297, 16'd8702, 16'd18038, 16'd8005, 16'd10985, 16'd38967, 16'd38217, 16'd21574, 16'd10277, 16'd7275, 16'd22345, 16'd24872, 16'd50637, 16'd59792, 16'd40339, 16'd10494, 16'd9255, 16'd32833, 16'd31851, 16'd37717, 16'd46370, 16'd23735, 16'd17904, 16'd1518, 16'd41001, 16'd18084});
	test_expansion(128'h9eecbfde82a51e1ad0b33ba9dd29810c, {16'd15502, 16'd43923, 16'd8170, 16'd8957, 16'd20706, 16'd33869, 16'd35047, 16'd54157, 16'd44737, 16'd49927, 16'd36764, 16'd19525, 16'd55106, 16'd20161, 16'd4018, 16'd38883, 16'd65348, 16'd52390, 16'd19888, 16'd10660, 16'd43486, 16'd19055, 16'd31749, 16'd22535, 16'd8740, 16'd56411});
	test_expansion(128'hbfe49bed050b0f1d06685a90d7377dbc, {16'd17259, 16'd61411, 16'd13136, 16'd29476, 16'd392, 16'd44617, 16'd47293, 16'd60593, 16'd27468, 16'd19162, 16'd13196, 16'd16619, 16'd50686, 16'd14663, 16'd62071, 16'd62697, 16'd20660, 16'd28005, 16'd43896, 16'd57489, 16'd20481, 16'd27684, 16'd41422, 16'd64742, 16'd39417, 16'd42459});
	test_expansion(128'h573d83274a62e70ac1fd8678223dcd73, {16'd63461, 16'd27012, 16'd45857, 16'd11913, 16'd47324, 16'd18002, 16'd727, 16'd37068, 16'd30809, 16'd55146, 16'd10418, 16'd44610, 16'd49145, 16'd13078, 16'd27712, 16'd2586, 16'd15475, 16'd15516, 16'd7772, 16'd33995, 16'd8244, 16'd64973, 16'd3935, 16'd60352, 16'd12788, 16'd20943});
	test_expansion(128'h4d5909ad51cd0cfde5d47189a0a9c3f7, {16'd57860, 16'd38514, 16'd53909, 16'd13004, 16'd64562, 16'd19715, 16'd9489, 16'd57627, 16'd60084, 16'd30887, 16'd39921, 16'd10527, 16'd38403, 16'd20414, 16'd31559, 16'd37009, 16'd38148, 16'd4370, 16'd25905, 16'd54270, 16'd26688, 16'd58229, 16'd14428, 16'd40282, 16'd19304, 16'd55962});
	test_expansion(128'hc6b14b619a4257e198bb8275d018ee96, {16'd21315, 16'd8539, 16'd63773, 16'd19541, 16'd8237, 16'd63046, 16'd21766, 16'd17823, 16'd28161, 16'd61990, 16'd65074, 16'd59247, 16'd49937, 16'd52438, 16'd48443, 16'd46328, 16'd5103, 16'd40152, 16'd15631, 16'd62957, 16'd39656, 16'd64860, 16'd32661, 16'd64535, 16'd4673, 16'd11917});
	test_expansion(128'h7301cc2f88ed0a68f1db3939c324c084, {16'd8272, 16'd61475, 16'd12315, 16'd62251, 16'd37566, 16'd58999, 16'd46259, 16'd49949, 16'd64788, 16'd31510, 16'd47469, 16'd48940, 16'd53628, 16'd55904, 16'd14866, 16'd9074, 16'd58349, 16'd29552, 16'd14585, 16'd25205, 16'd40677, 16'd17301, 16'd45126, 16'd36454, 16'd29555, 16'd28765});
	test_expansion(128'hc5e982e73919f607dbb4cd0c86846de6, {16'd1308, 16'd40822, 16'd4590, 16'd48577, 16'd12, 16'd5191, 16'd34625, 16'd36697, 16'd18986, 16'd48069, 16'd44870, 16'd5660, 16'd6684, 16'd8014, 16'd46051, 16'd22952, 16'd50675, 16'd29201, 16'd6476, 16'd59458, 16'd48883, 16'd8059, 16'd23685, 16'd64507, 16'd28240, 16'd5362});
	test_expansion(128'he452ce0127d2c870d381b8dd39a46dc0, {16'd53722, 16'd20348, 16'd50951, 16'd63535, 16'd19471, 16'd56838, 16'd40083, 16'd3129, 16'd25345, 16'd54333, 16'd43946, 16'd11785, 16'd51132, 16'd49098, 16'd56729, 16'd48105, 16'd52679, 16'd46963, 16'd1187, 16'd9092, 16'd49254, 16'd42618, 16'd49493, 16'd4199, 16'd59451, 16'd52383});
	test_expansion(128'h2fe5ef51f5b3fb58a3b12baa53671148, {16'd33697, 16'd5, 16'd4591, 16'd2883, 16'd45886, 16'd36290, 16'd56869, 16'd52666, 16'd53456, 16'd16911, 16'd36907, 16'd6092, 16'd33898, 16'd51335, 16'd11335, 16'd24181, 16'd33680, 16'd38351, 16'd22599, 16'd8985, 16'd17678, 16'd52020, 16'd33327, 16'd33793, 16'd60390, 16'd3498});
	test_expansion(128'h273d1c2ad8cc044d69aa9ef6cb46ed2e, {16'd390, 16'd17258, 16'd52679, 16'd45496, 16'd37558, 16'd49823, 16'd38259, 16'd41772, 16'd39029, 16'd50451, 16'd36990, 16'd28390, 16'd64615, 16'd29651, 16'd27592, 16'd63530, 16'd16642, 16'd34771, 16'd9684, 16'd22998, 16'd56885, 16'd10510, 16'd25736, 16'd44149, 16'd2456, 16'd11792});
	test_expansion(128'h3c01dd743f11ac42fd7f310fb210fd24, {16'd32829, 16'd62215, 16'd36230, 16'd34080, 16'd21413, 16'd41071, 16'd8756, 16'd49972, 16'd14155, 16'd54191, 16'd38010, 16'd40406, 16'd29623, 16'd13830, 16'd61137, 16'd30666, 16'd15239, 16'd14601, 16'd49832, 16'd47769, 16'd64923, 16'd17035, 16'd8592, 16'd34415, 16'd4480, 16'd40483});
	test_expansion(128'ha02de3b6608f22079f7566f24471c42d, {16'd60466, 16'd46288, 16'd6983, 16'd7618, 16'd43803, 16'd3016, 16'd920, 16'd7708, 16'd30399, 16'd34889, 16'd20984, 16'd14258, 16'd51693, 16'd47307, 16'd60724, 16'd15030, 16'd53764, 16'd61244, 16'd14613, 16'd14660, 16'd42703, 16'd26769, 16'd5562, 16'd30917, 16'd23572, 16'd31928});
	test_expansion(128'hfde0ecbf673e7d71747526a2456a824c, {16'd24031, 16'd26498, 16'd26576, 16'd30306, 16'd60530, 16'd54858, 16'd3058, 16'd34703, 16'd30710, 16'd49108, 16'd59659, 16'd28966, 16'd60777, 16'd55503, 16'd64347, 16'd23052, 16'd43987, 16'd25096, 16'd6585, 16'd41778, 16'd15226, 16'd61926, 16'd9617, 16'd14177, 16'd64321, 16'd39399});
	test_expansion(128'h35278c757c183d1217c996dc5b996812, {16'd533, 16'd55744, 16'd64802, 16'd9089, 16'd20154, 16'd11026, 16'd30780, 16'd51161, 16'd60951, 16'd45128, 16'd7733, 16'd58441, 16'd22306, 16'd27284, 16'd20317, 16'd33868, 16'd48566, 16'd13680, 16'd47361, 16'd56482, 16'd16695, 16'd35220, 16'd36362, 16'd9065, 16'd50287, 16'd46497});
	test_expansion(128'h6d84addfb9ae9a81dcb88aff0820cb4e, {16'd24152, 16'd43482, 16'd62075, 16'd42737, 16'd44493, 16'd12594, 16'd3504, 16'd12962, 16'd58710, 16'd10826, 16'd28295, 16'd39499, 16'd60622, 16'd59854, 16'd7800, 16'd22475, 16'd20406, 16'd29041, 16'd41364, 16'd37263, 16'd31028, 16'd20365, 16'd48290, 16'd39449, 16'd21556, 16'd50927});
	test_expansion(128'h5ecefce4c6fed354d205e9ecdf7965a4, {16'd56748, 16'd5712, 16'd49746, 16'd11090, 16'd28929, 16'd19586, 16'd64855, 16'd55977, 16'd46133, 16'd1437, 16'd27447, 16'd59997, 16'd35391, 16'd37995, 16'd44590, 16'd10704, 16'd53487, 16'd43466, 16'd33720, 16'd37005, 16'd12708, 16'd43567, 16'd24324, 16'd25127, 16'd4643, 16'd28268});
	test_expansion(128'hea1931a15ea0405a1aa1682aec475258, {16'd46979, 16'd3464, 16'd2442, 16'd64498, 16'd64225, 16'd42274, 16'd59337, 16'd10356, 16'd27949, 16'd22001, 16'd60023, 16'd17976, 16'd44726, 16'd53056, 16'd44810, 16'd53150, 16'd57590, 16'd63332, 16'd19797, 16'd23091, 16'd13208, 16'd40201, 16'd14512, 16'd4161, 16'd11930, 16'd17521});
	test_expansion(128'hf98128b9471d1eb3a722f6f3c6dfc387, {16'd429, 16'd62566, 16'd62005, 16'd44072, 16'd16833, 16'd26644, 16'd50342, 16'd42925, 16'd61973, 16'd9933, 16'd56390, 16'd10565, 16'd47168, 16'd37151, 16'd36282, 16'd6432, 16'd10503, 16'd26711, 16'd34397, 16'd29306, 16'd2424, 16'd38879, 16'd15106, 16'd58313, 16'd33417, 16'd62907});
	test_expansion(128'h4a037d963795674b0e933e866936ac95, {16'd13394, 16'd14986, 16'd38946, 16'd21351, 16'd36772, 16'd29461, 16'd24078, 16'd29750, 16'd20265, 16'd9186, 16'd39385, 16'd22840, 16'd39545, 16'd7258, 16'd10473, 16'd64963, 16'd39420, 16'd13615, 16'd45491, 16'd35735, 16'd37701, 16'd21550, 16'd56955, 16'd12756, 16'd38244, 16'd35872});
	test_expansion(128'hd55df483d23075f3f2e1a6dbc1428126, {16'd6920, 16'd3551, 16'd28314, 16'd64644, 16'd8636, 16'd49596, 16'd20135, 16'd49440, 16'd44238, 16'd64011, 16'd1118, 16'd14946, 16'd15084, 16'd37691, 16'd31471, 16'd15244, 16'd62788, 16'd10862, 16'd52977, 16'd13403, 16'd29219, 16'd49999, 16'd10593, 16'd47847, 16'd61443, 16'd47920});
	test_expansion(128'hbd59018d619e2184956a51b700d15535, {16'd43494, 16'd34821, 16'd28413, 16'd8539, 16'd35616, 16'd18441, 16'd20840, 16'd27631, 16'd25306, 16'd58157, 16'd54839, 16'd60567, 16'd21854, 16'd16836, 16'd57716, 16'd23103, 16'd59535, 16'd16025, 16'd6787, 16'd45709, 16'd59861, 16'd57592, 16'd626, 16'd33202, 16'd16381, 16'd64388});
	test_expansion(128'h38c222d7b704b0c1086b49c8b6ee429d, {16'd465, 16'd54594, 16'd6896, 16'd12736, 16'd25125, 16'd62136, 16'd12084, 16'd14755, 16'd37146, 16'd31465, 16'd33145, 16'd65282, 16'd10968, 16'd7648, 16'd41501, 16'd919, 16'd34678, 16'd8186, 16'd57555, 16'd25432, 16'd354, 16'd44707, 16'd65045, 16'd45068, 16'd36220, 16'd8413});
	test_expansion(128'h883115cc16cbd6d90590175226ae1261, {16'd57511, 16'd52402, 16'd17093, 16'd57699, 16'd54108, 16'd42494, 16'd51661, 16'd25617, 16'd63306, 16'd4918, 16'd30243, 16'd28201, 16'd20368, 16'd12019, 16'd25338, 16'd52874, 16'd44916, 16'd51765, 16'd6535, 16'd50855, 16'd13724, 16'd6034, 16'd45217, 16'd62047, 16'd2244, 16'd28914});
	test_expansion(128'ha5d769d44fb4e245be23127c62a4261e, {16'd44483, 16'd11638, 16'd61317, 16'd52821, 16'd47203, 16'd39924, 16'd44083, 16'd8902, 16'd58427, 16'd9057, 16'd60787, 16'd22975, 16'd6927, 16'd58718, 16'd55733, 16'd52723, 16'd14663, 16'd13854, 16'd9297, 16'd19806, 16'd44101, 16'd22498, 16'd12129, 16'd27023, 16'd37297, 16'd499});
	test_expansion(128'h2bdce1f660e8380866c813b055e19db5, {16'd59785, 16'd32092, 16'd23114, 16'd18894, 16'd28061, 16'd53695, 16'd20580, 16'd48003, 16'd64189, 16'd60001, 16'd52221, 16'd13820, 16'd27925, 16'd63524, 16'd10813, 16'd19508, 16'd39605, 16'd44769, 16'd8445, 16'd44048, 16'd57554, 16'd35100, 16'd57799, 16'd22599, 16'd47275, 16'd34762});
	test_expansion(128'h1db2d15f83c099e5ea872a3f8a9adf26, {16'd52697, 16'd48962, 16'd27143, 16'd21474, 16'd4372, 16'd2373, 16'd1286, 16'd31385, 16'd20425, 16'd17160, 16'd32773, 16'd51579, 16'd39224, 16'd45941, 16'd59056, 16'd62906, 16'd36998, 16'd20537, 16'd46634, 16'd43282, 16'd46663, 16'd38414, 16'd23954, 16'd5154, 16'd35621, 16'd55443});
	test_expansion(128'h6b96116bb20a26b00203d3a9f5fd010c, {16'd40687, 16'd1245, 16'd31861, 16'd56093, 16'd54519, 16'd26423, 16'd41491, 16'd54856, 16'd50284, 16'd5413, 16'd53896, 16'd56785, 16'd48483, 16'd50167, 16'd16870, 16'd23691, 16'd31326, 16'd59111, 16'd7067, 16'd18441, 16'd5314, 16'd37368, 16'd8776, 16'd7159, 16'd18031, 16'd6590});
	test_expansion(128'h7952ae02c3e2d6f58331c6f6f420801e, {16'd29183, 16'd59569, 16'd48114, 16'd42741, 16'd36066, 16'd16140, 16'd5339, 16'd43688, 16'd46894, 16'd58294, 16'd25507, 16'd32336, 16'd15870, 16'd39599, 16'd49965, 16'd45151, 16'd5440, 16'd62938, 16'd55739, 16'd39143, 16'd39317, 16'd50189, 16'd36722, 16'd7403, 16'd25373, 16'd55203});
	test_expansion(128'he8dfc7144f5ef43046c33247ca75f591, {16'd58778, 16'd39561, 16'd52233, 16'd36329, 16'd20013, 16'd2254, 16'd54219, 16'd42463, 16'd63481, 16'd17175, 16'd44660, 16'd59616, 16'd64577, 16'd58759, 16'd42227, 16'd3760, 16'd43812, 16'd30145, 16'd33618, 16'd51964, 16'd51395, 16'd43790, 16'd24259, 16'd15558, 16'd55851, 16'd36366});
	test_expansion(128'h4318fc76f0772bd167dc4edb159f2e11, {16'd37475, 16'd31845, 16'd31809, 16'd5757, 16'd45924, 16'd21248, 16'd3665, 16'd18335, 16'd22984, 16'd33591, 16'd38984, 16'd19913, 16'd30014, 16'd50785, 16'd63959, 16'd26120, 16'd64635, 16'd62341, 16'd60379, 16'd59224, 16'd269, 16'd36076, 16'd21737, 16'd14615, 16'd5006, 16'd62845});
	test_expansion(128'hbb4dbce8d95b03187c4ab23be9b369d3, {16'd56525, 16'd44432, 16'd6826, 16'd61482, 16'd26540, 16'd36198, 16'd38529, 16'd28861, 16'd53462, 16'd29837, 16'd15975, 16'd18657, 16'd23832, 16'd4873, 16'd43302, 16'd45098, 16'd16687, 16'd45541, 16'd24367, 16'd60799, 16'd45099, 16'd6904, 16'd37854, 16'd8176, 16'd57959, 16'd39680});
	test_expansion(128'h537390f36b16cb4cfad44c0f7c727a9d, {16'd47022, 16'd14681, 16'd27032, 16'd40890, 16'd9676, 16'd46887, 16'd33369, 16'd35272, 16'd19585, 16'd45231, 16'd2589, 16'd19709, 16'd53620, 16'd38655, 16'd49483, 16'd26081, 16'd34103, 16'd860, 16'd41489, 16'd47367, 16'd40972, 16'd59913, 16'd13459, 16'd21642, 16'd60630, 16'd33807});
	test_expansion(128'h537122ed8fc60e60792ac5f90c084019, {16'd22861, 16'd4273, 16'd40841, 16'd29712, 16'd46938, 16'd25045, 16'd54494, 16'd49190, 16'd44318, 16'd23183, 16'd16039, 16'd2593, 16'd43067, 16'd65105, 16'd64000, 16'd55988, 16'd37775, 16'd34207, 16'd5522, 16'd49829, 16'd4488, 16'd7308, 16'd46095, 16'd50163, 16'd29275, 16'd28561});
	test_expansion(128'h917915eb0ea7b939b3a99062df037e71, {16'd54507, 16'd3659, 16'd10741, 16'd28147, 16'd11181, 16'd2099, 16'd34830, 16'd21019, 16'd19543, 16'd59977, 16'd60431, 16'd61019, 16'd45470, 16'd16328, 16'd21652, 16'd45742, 16'd19914, 16'd26938, 16'd49356, 16'd57230, 16'd54214, 16'd39724, 16'd31941, 16'd48088, 16'd48470, 16'd37226});
	test_expansion(128'h2add3fc97018c960151ad01f989eb949, {16'd22384, 16'd49765, 16'd36041, 16'd16331, 16'd56609, 16'd39028, 16'd56881, 16'd15559, 16'd2782, 16'd17761, 16'd65492, 16'd10162, 16'd36692, 16'd7236, 16'd35719, 16'd64648, 16'd15635, 16'd57168, 16'd46135, 16'd61907, 16'd29943, 16'd10506, 16'd4132, 16'd19883, 16'd41209, 16'd64684});
	test_expansion(128'h0ef213606263461797622710a3852337, {16'd1619, 16'd33067, 16'd64670, 16'd41816, 16'd44560, 16'd575, 16'd8088, 16'd54035, 16'd20856, 16'd45957, 16'd28351, 16'd7624, 16'd712, 16'd61997, 16'd42756, 16'd49892, 16'd34209, 16'd57606, 16'd56810, 16'd17728, 16'd61641, 16'd51530, 16'd15525, 16'd20990, 16'd36833, 16'd41219});
	test_expansion(128'h370d49b1dbeededa9ef81debb185fb2d, {16'd24956, 16'd63291, 16'd19347, 16'd56636, 16'd12184, 16'd52854, 16'd56020, 16'd26650, 16'd3690, 16'd53143, 16'd24885, 16'd46401, 16'd37400, 16'd23349, 16'd52550, 16'd2228, 16'd11306, 16'd23658, 16'd8688, 16'd54982, 16'd56994, 16'd20977, 16'd38788, 16'd57893, 16'd65140, 16'd43232});
	test_expansion(128'h391dc706e3e6f3ec857f2f21fd870ba9, {16'd22446, 16'd36784, 16'd63239, 16'd55778, 16'd7107, 16'd30362, 16'd16118, 16'd10479, 16'd53174, 16'd31169, 16'd23654, 16'd50492, 16'd41233, 16'd63137, 16'd27974, 16'd49665, 16'd32662, 16'd58399, 16'd15534, 16'd16234, 16'd51664, 16'd43453, 16'd28922, 16'd40311, 16'd1041, 16'd2536});
	test_expansion(128'ha44ddb347aa0d095d068fcf7c71e88b2, {16'd27276, 16'd63590, 16'd6913, 16'd13627, 16'd17983, 16'd11441, 16'd36613, 16'd64155, 16'd21963, 16'd8698, 16'd46246, 16'd59110, 16'd19167, 16'd32901, 16'd5446, 16'd31107, 16'd33497, 16'd28086, 16'd2687, 16'd50514, 16'd60255, 16'd14920, 16'd23199, 16'd39751, 16'd7421, 16'd37428});
	test_expansion(128'h940fc633367b618986b88a8b8fac9e6e, {16'd22749, 16'd3922, 16'd26566, 16'd36355, 16'd19115, 16'd44940, 16'd36573, 16'd23046, 16'd63692, 16'd56843, 16'd18356, 16'd39716, 16'd29128, 16'd65249, 16'd33368, 16'd29183, 16'd65246, 16'd63817, 16'd20858, 16'd45669, 16'd12636, 16'd32835, 16'd60149, 16'd49972, 16'd53854, 16'd20982});
	test_expansion(128'hfdd4cf3f43e8ac30b2a72f33b87f7ed2, {16'd61552, 16'd33190, 16'd56255, 16'd62585, 16'd41994, 16'd44487, 16'd60604, 16'd51645, 16'd13380, 16'd16352, 16'd11692, 16'd6088, 16'd35090, 16'd34282, 16'd41039, 16'd30211, 16'd6109, 16'd30650, 16'd17262, 16'd4326, 16'd64002, 16'd46929, 16'd31655, 16'd35706, 16'd35963, 16'd22704});
	test_expansion(128'h20d1631821295f8e119b26ceeca30d47, {16'd5713, 16'd39357, 16'd1049, 16'd20722, 16'd44025, 16'd12150, 16'd34275, 16'd55261, 16'd13397, 16'd24304, 16'd44404, 16'd14763, 16'd3939, 16'd54656, 16'd31452, 16'd34902, 16'd16486, 16'd41707, 16'd15884, 16'd9281, 16'd48248, 16'd16016, 16'd31410, 16'd55762, 16'd25656, 16'd43374});
	test_expansion(128'hcd00ad29633fce4585ab1c41a40cdf6e, {16'd21951, 16'd21015, 16'd48427, 16'd11079, 16'd40648, 16'd18180, 16'd29113, 16'd33108, 16'd53364, 16'd21837, 16'd43431, 16'd33622, 16'd61919, 16'd38646, 16'd28738, 16'd13798, 16'd9059, 16'd64090, 16'd35213, 16'd22792, 16'd58848, 16'd11897, 16'd53872, 16'd64227, 16'd44211, 16'd46359});
	test_expansion(128'h63ab683ab47a80b49983bddd27d0c260, {16'd53060, 16'd664, 16'd41714, 16'd5868, 16'd59935, 16'd26130, 16'd11047, 16'd22561, 16'd23861, 16'd4471, 16'd53956, 16'd3437, 16'd47010, 16'd34340, 16'd22946, 16'd459, 16'd63464, 16'd24380, 16'd46305, 16'd27866, 16'd53798, 16'd58765, 16'd10082, 16'd57278, 16'd62774, 16'd33497});
	test_expansion(128'hcd4ae0766ecfd05700d15c36cff7c4d7, {16'd37859, 16'd7869, 16'd64501, 16'd12896, 16'd20380, 16'd61970, 16'd58546, 16'd26007, 16'd2828, 16'd32939, 16'd12336, 16'd22491, 16'd19779, 16'd16084, 16'd61440, 16'd21734, 16'd57859, 16'd19177, 16'd58822, 16'd21010, 16'd41777, 16'd52133, 16'd10109, 16'd12703, 16'd6305, 16'd17200});
	test_expansion(128'hf49e41c889f7bdfc81550589cf4a6110, {16'd53486, 16'd7607, 16'd47771, 16'd2176, 16'd16782, 16'd10197, 16'd58586, 16'd65503, 16'd25170, 16'd13954, 16'd56867, 16'd3805, 16'd30377, 16'd45919, 16'd55824, 16'd15326, 16'd48309, 16'd24806, 16'd33513, 16'd8543, 16'd28637, 16'd28438, 16'd59539, 16'd49760, 16'd63626, 16'd2977});
	test_expansion(128'h33399b0145790a54cba98e0da2ce807d, {16'd56660, 16'd14762, 16'd35941, 16'd58, 16'd5527, 16'd26482, 16'd24126, 16'd61621, 16'd41204, 16'd63946, 16'd48887, 16'd50336, 16'd27617, 16'd57666, 16'd58361, 16'd65500, 16'd27512, 16'd35184, 16'd30093, 16'd65295, 16'd57972, 16'd18504, 16'd33290, 16'd62768, 16'd41614, 16'd54350});
	test_expansion(128'h4f7f5af526b8eec396f8414d9d0f8eb6, {16'd22555, 16'd57350, 16'd42391, 16'd55930, 16'd38333, 16'd19681, 16'd7553, 16'd48388, 16'd62817, 16'd61412, 16'd44176, 16'd51255, 16'd4559, 16'd58739, 16'd3177, 16'd23690, 16'd59834, 16'd63016, 16'd11545, 16'd25832, 16'd40597, 16'd63786, 16'd62177, 16'd51907, 16'd6466, 16'd22332});
	test_expansion(128'hfa32b1e21c46b30df4e271a09622bade, {16'd38115, 16'd47044, 16'd19823, 16'd35304, 16'd4348, 16'd759, 16'd53748, 16'd30430, 16'd51879, 16'd27067, 16'd8544, 16'd62872, 16'd45220, 16'd31520, 16'd50609, 16'd42291, 16'd38160, 16'd56496, 16'd32501, 16'd45767, 16'd4521, 16'd34347, 16'd23303, 16'd47343, 16'd20901, 16'd14288});
	test_expansion(128'he2256319052b77f7b2c9ea46f07b8976, {16'd62490, 16'd62564, 16'd63225, 16'd21796, 16'd42258, 16'd23192, 16'd32417, 16'd47542, 16'd41316, 16'd52703, 16'd2801, 16'd16982, 16'd3117, 16'd21273, 16'd26374, 16'd25421, 16'd58091, 16'd2343, 16'd59318, 16'd40200, 16'd1455, 16'd29841, 16'd62682, 16'd52088, 16'd55792, 16'd18148});
	test_expansion(128'h8de1323550aaac62cb71ee3905307347, {16'd11148, 16'd64425, 16'd7844, 16'd53927, 16'd18045, 16'd589, 16'd40625, 16'd33741, 16'd26285, 16'd37688, 16'd10239, 16'd49139, 16'd35744, 16'd32513, 16'd15763, 16'd9222, 16'd34533, 16'd47930, 16'd57065, 16'd58954, 16'd5865, 16'd41226, 16'd58210, 16'd22791, 16'd51909, 16'd58527});
	test_expansion(128'he898612e2a08f6d7312c4ce1b9e33b22, {16'd49277, 16'd43247, 16'd40332, 16'd16980, 16'd60379, 16'd39510, 16'd21834, 16'd35730, 16'd9986, 16'd10288, 16'd51652, 16'd58330, 16'd6147, 16'd26525, 16'd10483, 16'd56911, 16'd9227, 16'd3529, 16'd34448, 16'd55997, 16'd22097, 16'd23429, 16'd36512, 16'd20591, 16'd12940, 16'd58355});
	test_expansion(128'h19c3487ac68fca086f4e6780250f69c0, {16'd42377, 16'd8113, 16'd23435, 16'd6493, 16'd31762, 16'd6313, 16'd24461, 16'd24898, 16'd39119, 16'd19887, 16'd8008, 16'd40983, 16'd15304, 16'd27345, 16'd27880, 16'd60795, 16'd15929, 16'd51097, 16'd28230, 16'd22253, 16'd50420, 16'd2824, 16'd47093, 16'd19826, 16'd64477, 16'd19910});
	test_expansion(128'h7b265ea71ba902effe30233f72017799, {16'd21996, 16'd7770, 16'd55395, 16'd40034, 16'd25064, 16'd966, 16'd63398, 16'd30414, 16'd39179, 16'd53461, 16'd36838, 16'd43345, 16'd6333, 16'd44849, 16'd53785, 16'd22145, 16'd44384, 16'd38189, 16'd28181, 16'd65391, 16'd21349, 16'd60182, 16'd16060, 16'd60990, 16'd15, 16'd60244});
	test_expansion(128'h6e4a432bed3ded1affa23ae40ac76b16, {16'd38847, 16'd45680, 16'd56505, 16'd31535, 16'd50229, 16'd40983, 16'd24634, 16'd43202, 16'd8647, 16'd47184, 16'd64139, 16'd52680, 16'd1751, 16'd39517, 16'd64565, 16'd51765, 16'd5882, 16'd13677, 16'd7731, 16'd59878, 16'd34584, 16'd21596, 16'd49399, 16'd9845, 16'd30891, 16'd45146});
	test_expansion(128'h10213d27d58a74db446a93b141a7e52a, {16'd55569, 16'd52851, 16'd4633, 16'd18965, 16'd63015, 16'd19924, 16'd31256, 16'd32533, 16'd48263, 16'd56422, 16'd4097, 16'd437, 16'd206, 16'd57969, 16'd17299, 16'd64730, 16'd5805, 16'd29531, 16'd36223, 16'd22368, 16'd33243, 16'd64743, 16'd49396, 16'd28207, 16'd46797, 16'd9611});
	test_expansion(128'h2b945a23e367849de615bfce03f33b5c, {16'd41186, 16'd15300, 16'd58783, 16'd36101, 16'd22334, 16'd10244, 16'd42701, 16'd64572, 16'd26614, 16'd37841, 16'd43721, 16'd59745, 16'd30895, 16'd41175, 16'd38348, 16'd62095, 16'd30176, 16'd60607, 16'd41101, 16'd5436, 16'd44524, 16'd38715, 16'd47687, 16'd37550, 16'd41455, 16'd43261});
	test_expansion(128'h9862f4b6ac4a0f905c6bff934784c77a, {16'd21031, 16'd39274, 16'd21147, 16'd47106, 16'd46115, 16'd50120, 16'd23976, 16'd60523, 16'd32821, 16'd4234, 16'd32312, 16'd44363, 16'd7604, 16'd30254, 16'd24653, 16'd48935, 16'd37710, 16'd40479, 16'd18157, 16'd13895, 16'd56198, 16'd18070, 16'd13391, 16'd10993, 16'd42212, 16'd44901});
	test_expansion(128'hd89bbb5be53ec81f73f3e386d4778c4f, {16'd37765, 16'd61569, 16'd64842, 16'd10689, 16'd21176, 16'd45730, 16'd47212, 16'd61316, 16'd27718, 16'd15533, 16'd46259, 16'd63003, 16'd33406, 16'd56163, 16'd57550, 16'd58598, 16'd5361, 16'd14529, 16'd10049, 16'd28526, 16'd7947, 16'd49556, 16'd1818, 16'd40504, 16'd38284, 16'd40617});
	test_expansion(128'hafff337a8bbe41c66fec1c9eec454540, {16'd21980, 16'd2331, 16'd40195, 16'd19068, 16'd21524, 16'd12604, 16'd39276, 16'd41696, 16'd28317, 16'd9858, 16'd41057, 16'd41922, 16'd27012, 16'd49354, 16'd17919, 16'd20879, 16'd7880, 16'd23259, 16'd49362, 16'd55152, 16'd40398, 16'd47965, 16'd14647, 16'd40330, 16'd3188, 16'd59021});
	test_expansion(128'h96850ceee169ef1be8499e5b141ba5d4, {16'd265, 16'd57016, 16'd47781, 16'd28293, 16'd11605, 16'd33898, 16'd14629, 16'd8718, 16'd4801, 16'd8803, 16'd57811, 16'd48336, 16'd11661, 16'd42476, 16'd40326, 16'd27086, 16'd31416, 16'd17950, 16'd56470, 16'd62586, 16'd24561, 16'd62994, 16'd52247, 16'd47258, 16'd5792, 16'd49632});
	test_expansion(128'h5ad9c8896f43c904e877d7150195baab, {16'd55810, 16'd49426, 16'd23111, 16'd51988, 16'd56525, 16'd53581, 16'd13288, 16'd30957, 16'd13358, 16'd49977, 16'd21157, 16'd31761, 16'd41496, 16'd27963, 16'd20440, 16'd27914, 16'd6378, 16'd39865, 16'd12543, 16'd19661, 16'd8903, 16'd45494, 16'd24665, 16'd53023, 16'd59411, 16'd9905});
	test_expansion(128'hc7dbf7e1aacbe5c1fa66aecc9914170a, {16'd32212, 16'd47450, 16'd50098, 16'd36178, 16'd57949, 16'd54615, 16'd18044, 16'd3978, 16'd5198, 16'd59088, 16'd61161, 16'd12678, 16'd30354, 16'd4197, 16'd52003, 16'd27913, 16'd48229, 16'd2713, 16'd50694, 16'd63689, 16'd3998, 16'd63888, 16'd1898, 16'd39447, 16'd20879, 16'd29712});
	test_expansion(128'h6db86f3205ce8c3e8bd97e39492cc8d5, {16'd47555, 16'd2383, 16'd2728, 16'd2453, 16'd31235, 16'd24157, 16'd14554, 16'd42662, 16'd36250, 16'd52439, 16'd1416, 16'd46902, 16'd39406, 16'd15599, 16'd45056, 16'd55960, 16'd17515, 16'd55431, 16'd33059, 16'd39679, 16'd29317, 16'd17180, 16'd60824, 16'd6792, 16'd46509, 16'd21073});
	test_expansion(128'hf7ceca740d6dd7d577cb3ee27b908409, {16'd25016, 16'd9611, 16'd48924, 16'd51107, 16'd64445, 16'd2280, 16'd56973, 16'd24378, 16'd30428, 16'd25511, 16'd35750, 16'd39232, 16'd22651, 16'd59461, 16'd63134, 16'd43629, 16'd21845, 16'd5041, 16'd19990, 16'd18281, 16'd14220, 16'd20815, 16'd17158, 16'd56485, 16'd30039, 16'd60436});
	test_expansion(128'hb858852feca5cc8087abdf662c34052e, {16'd32774, 16'd63460, 16'd802, 16'd35869, 16'd18357, 16'd30354, 16'd43982, 16'd48169, 16'd18697, 16'd40680, 16'd62986, 16'd16217, 16'd19911, 16'd36318, 16'd55522, 16'd2241, 16'd61963, 16'd19744, 16'd38924, 16'd16248, 16'd19736, 16'd35391, 16'd9379, 16'd50858, 16'd42088, 16'd21048});
	test_expansion(128'h89294ee050947819df2ed9caa6c2a847, {16'd53431, 16'd44606, 16'd3558, 16'd18729, 16'd44031, 16'd53515, 16'd52224, 16'd58786, 16'd34902, 16'd58007, 16'd61763, 16'd42369, 16'd42934, 16'd29752, 16'd34136, 16'd6071, 16'd63859, 16'd10585, 16'd24006, 16'd31856, 16'd26198, 16'd46193, 16'd38771, 16'd18143, 16'd8774, 16'd17292});
	test_expansion(128'hc286a1defffc9d5454f2d3ba7abaa10f, {16'd21172, 16'd6103, 16'd27763, 16'd4991, 16'd55457, 16'd58202, 16'd17459, 16'd11282, 16'd48489, 16'd50995, 16'd41280, 16'd27422, 16'd40710, 16'd53634, 16'd61333, 16'd9014, 16'd15359, 16'd36884, 16'd21958, 16'd4910, 16'd5078, 16'd16487, 16'd5406, 16'd39565, 16'd17975, 16'd32206});
	test_expansion(128'he3666e14a29990ae352a1e6b64216b64, {16'd58225, 16'd54750, 16'd38227, 16'd41989, 16'd15421, 16'd51427, 16'd48921, 16'd24272, 16'd43667, 16'd46017, 16'd1663, 16'd60120, 16'd64463, 16'd52025, 16'd38779, 16'd50256, 16'd27317, 16'd10714, 16'd43692, 16'd13056, 16'd39029, 16'd7689, 16'd28978, 16'd46885, 16'd4465, 16'd37403});
	test_expansion(128'h2b3dcfc8103fc6edf07e46313c94e746, {16'd23788, 16'd20203, 16'd44772, 16'd11754, 16'd6555, 16'd38736, 16'd47100, 16'd58988, 16'd49327, 16'd455, 16'd36964, 16'd10103, 16'd17692, 16'd31003, 16'd25538, 16'd30796, 16'd29874, 16'd62463, 16'd63720, 16'd61670, 16'd12980, 16'd53809, 16'd12994, 16'd49748, 16'd48386, 16'd28466});
	test_expansion(128'h11b7ae2c42817a674a05836114509120, {16'd63783, 16'd23712, 16'd24765, 16'd63724, 16'd26442, 16'd43031, 16'd2279, 16'd6857, 16'd53015, 16'd52759, 16'd12212, 16'd42853, 16'd56955, 16'd7958, 16'd4511, 16'd52047, 16'd9887, 16'd27261, 16'd49819, 16'd6847, 16'd53990, 16'd57455, 16'd32564, 16'd61577, 16'd24674, 16'd49514});
	test_expansion(128'h32e7ba064d2f2e9f41263ee040c286ee, {16'd52141, 16'd37262, 16'd19605, 16'd43804, 16'd20656, 16'd60310, 16'd56554, 16'd13692, 16'd46538, 16'd37887, 16'd63951, 16'd33129, 16'd21283, 16'd44878, 16'd21154, 16'd9918, 16'd36775, 16'd27877, 16'd36193, 16'd10870, 16'd49934, 16'd46586, 16'd19232, 16'd59839, 16'd14140, 16'd44001});
	test_expansion(128'h19bedcd4798afaa046e1087b766ef7ad, {16'd47316, 16'd63578, 16'd938, 16'd60670, 16'd56709, 16'd491, 16'd48505, 16'd2070, 16'd13312, 16'd62580, 16'd58724, 16'd40483, 16'd23933, 16'd13342, 16'd22980, 16'd5840, 16'd53051, 16'd24324, 16'd57996, 16'd35975, 16'd61461, 16'd16935, 16'd26788, 16'd32613, 16'd7597, 16'd20454});
	test_expansion(128'h6fb197155d5ab54bde54abc71cd2fbce, {16'd44010, 16'd3647, 16'd16261, 16'd16894, 16'd9847, 16'd57883, 16'd25191, 16'd15154, 16'd19585, 16'd48773, 16'd35578, 16'd51457, 16'd11723, 16'd46262, 16'd19262, 16'd5325, 16'd13337, 16'd18766, 16'd2008, 16'd56803, 16'd35707, 16'd34105, 16'd13360, 16'd57187, 16'd46227, 16'd56466});
	test_expansion(128'h8fed87327aeb272dfebe253c9d9c0752, {16'd919, 16'd46013, 16'd22999, 16'd133, 16'd51617, 16'd32808, 16'd19588, 16'd6781, 16'd8592, 16'd50547, 16'd63909, 16'd45654, 16'd54162, 16'd30679, 16'd26697, 16'd62335, 16'd5817, 16'd20145, 16'd53373, 16'd58917, 16'd15383, 16'd54178, 16'd62347, 16'd28897, 16'd58768, 16'd16957});
	test_expansion(128'h31ca1e34d88dda143efee4b1f242085a, {16'd48988, 16'd247, 16'd3570, 16'd59034, 16'd30153, 16'd3170, 16'd21303, 16'd5421, 16'd46927, 16'd42832, 16'd7294, 16'd53711, 16'd1843, 16'd5285, 16'd25006, 16'd31535, 16'd6759, 16'd5400, 16'd23114, 16'd31139, 16'd6932, 16'd62503, 16'd4347, 16'd1309, 16'd4979, 16'd29644});
	test_expansion(128'h0d150783e9e40604d63084387de8659c, {16'd31321, 16'd58500, 16'd3174, 16'd37308, 16'd32462, 16'd50688, 16'd17446, 16'd11427, 16'd48251, 16'd35024, 16'd6868, 16'd20348, 16'd13531, 16'd51274, 16'd17807, 16'd58402, 16'd8921, 16'd52575, 16'd44436, 16'd3106, 16'd15108, 16'd27793, 16'd2147, 16'd12661, 16'd41402, 16'd29400});
	test_expansion(128'hfc6f818a36236d66cc1efdd988c5b14f, {16'd56231, 16'd59828, 16'd14927, 16'd21038, 16'd30168, 16'd50568, 16'd20709, 16'd41055, 16'd13108, 16'd14599, 16'd52745, 16'd35059, 16'd35039, 16'd30653, 16'd56932, 16'd33112, 16'd47130, 16'd13383, 16'd54726, 16'd40872, 16'd14567, 16'd43739, 16'd12597, 16'd11256, 16'd15745, 16'd54132});
	test_expansion(128'h21de6d02ce0864b5d28c0872f87dbf17, {16'd62586, 16'd46571, 16'd8920, 16'd47984, 16'd13593, 16'd10784, 16'd26986, 16'd55632, 16'd13906, 16'd35067, 16'd57255, 16'd37354, 16'd19700, 16'd9400, 16'd58177, 16'd44978, 16'd44380, 16'd18519, 16'd57729, 16'd44514, 16'd727, 16'd35804, 16'd34411, 16'd57714, 16'd53497, 16'd2770});
	test_expansion(128'ha004b1913ee2ab50a78e0c4fc37e369d, {16'd60964, 16'd61835, 16'd34601, 16'd42272, 16'd46972, 16'd16457, 16'd7995, 16'd45643, 16'd53103, 16'd20683, 16'd27563, 16'd58718, 16'd38558, 16'd25051, 16'd61404, 16'd63059, 16'd65131, 16'd25342, 16'd6937, 16'd22852, 16'd15372, 16'd64614, 16'd15891, 16'd21383, 16'd48152, 16'd44090});
	test_expansion(128'h3d7d121857e9bf7fd170f3be6b2dc913, {16'd12308, 16'd59045, 16'd17889, 16'd56214, 16'd15769, 16'd9280, 16'd1145, 16'd36388, 16'd51894, 16'd63018, 16'd15608, 16'd23144, 16'd1123, 16'd27416, 16'd35992, 16'd37097, 16'd35047, 16'd60517, 16'd37364, 16'd31920, 16'd51318, 16'd30748, 16'd24941, 16'd34631, 16'd12177, 16'd45604});
	test_expansion(128'hc700dc91b487a9813dfd0a4555ddfe32, {16'd47181, 16'd61615, 16'd21351, 16'd40877, 16'd44007, 16'd49322, 16'd61191, 16'd37707, 16'd60079, 16'd3851, 16'd13, 16'd41364, 16'd7660, 16'd31735, 16'd40551, 16'd54777, 16'd48360, 16'd37693, 16'd55204, 16'd51119, 16'd21450, 16'd10927, 16'd25752, 16'd34929, 16'd43001, 16'd7398});
	test_expansion(128'hc64296d85bb37eb5d2d67f15c6194cb2, {16'd64535, 16'd48521, 16'd23699, 16'd47471, 16'd64311, 16'd36764, 16'd2654, 16'd7883, 16'd63412, 16'd46471, 16'd3130, 16'd42405, 16'd22367, 16'd39523, 16'd47549, 16'd35311, 16'd58575, 16'd58770, 16'd57122, 16'd21938, 16'd38745, 16'd10488, 16'd3692, 16'd43411, 16'd51054, 16'd39665});
	test_expansion(128'ha3db6e9a750e715cf71f9839ec4c8090, {16'd17314, 16'd18259, 16'd46122, 16'd50532, 16'd55908, 16'd46803, 16'd62086, 16'd34378, 16'd18737, 16'd12473, 16'd53938, 16'd19690, 16'd34612, 16'd31090, 16'd6485, 16'd55928, 16'd116, 16'd5863, 16'd52587, 16'd14488, 16'd46656, 16'd6418, 16'd53913, 16'd59393, 16'd10621, 16'd21881});
	test_expansion(128'hc7a4195d9ff6324a1cc3f6da4532d80a, {16'd40560, 16'd15687, 16'd21963, 16'd27275, 16'd4821, 16'd21339, 16'd39105, 16'd28249, 16'd64016, 16'd3779, 16'd1019, 16'd8933, 16'd44768, 16'd41896, 16'd15676, 16'd42019, 16'd41298, 16'd59257, 16'd23327, 16'd14956, 16'd47094, 16'd61336, 16'd40483, 16'd43189, 16'd30293, 16'd65054});
	test_expansion(128'h5260b5c2d5289c7d7b70b7365cf77a87, {16'd36006, 16'd13809, 16'd43686, 16'd63267, 16'd58267, 16'd56606, 16'd34872, 16'd18653, 16'd44089, 16'd20384, 16'd48193, 16'd54095, 16'd40922, 16'd30904, 16'd32481, 16'd25165, 16'd25610, 16'd52104, 16'd54247, 16'd10564, 16'd39744, 16'd36156, 16'd63284, 16'd45317, 16'd20215, 16'd29115});
	test_expansion(128'h0150b72543bd5b5dc0be550cc6908483, {16'd34248, 16'd43765, 16'd7413, 16'd31798, 16'd22721, 16'd61596, 16'd60442, 16'd45290, 16'd46, 16'd5775, 16'd41003, 16'd25346, 16'd42290, 16'd63767, 16'd52338, 16'd8446, 16'd9298, 16'd49229, 16'd1897, 16'd16889, 16'd41812, 16'd31791, 16'd19126, 16'd6614, 16'd31087, 16'd64246});
	test_expansion(128'hbef3be8bbd6362e4fb0a43267718aafe, {16'd58232, 16'd34605, 16'd53413, 16'd971, 16'd61236, 16'd41190, 16'd56884, 16'd38467, 16'd6657, 16'd48605, 16'd31731, 16'd56830, 16'd1242, 16'd34279, 16'd1013, 16'd44760, 16'd34991, 16'd53356, 16'd62382, 16'd48715, 16'd63657, 16'd41545, 16'd5836, 16'd64551, 16'd11533, 16'd43298});
	test_expansion(128'h96aa6bb3eea6a3d5905e3e026cc1e730, {16'd60582, 16'd41763, 16'd23728, 16'd55658, 16'd3213, 16'd12285, 16'd64771, 16'd47915, 16'd59073, 16'd28199, 16'd44783, 16'd28991, 16'd53268, 16'd25550, 16'd55874, 16'd7784, 16'd14306, 16'd52792, 16'd57307, 16'd44896, 16'd23713, 16'd25280, 16'd22789, 16'd47728, 16'd9632, 16'd14711});
	test_expansion(128'h0b59c1ba38b67d14fa935108d2891989, {16'd36908, 16'd45700, 16'd45520, 16'd25831, 16'd64605, 16'd38448, 16'd27936, 16'd8902, 16'd14575, 16'd30020, 16'd11393, 16'd40112, 16'd64038, 16'd54286, 16'd52739, 16'd32267, 16'd26911, 16'd51676, 16'd18591, 16'd35840, 16'd52451, 16'd21825, 16'd43675, 16'd55093, 16'd37385, 16'd7896});
	test_expansion(128'h709a32e55ecfaf266e19057a1db5c349, {16'd30280, 16'd154, 16'd37533, 16'd321, 16'd48258, 16'd36712, 16'd23079, 16'd5148, 16'd50811, 16'd11487, 16'd5124, 16'd3574, 16'd36314, 16'd3084, 16'd40841, 16'd13324, 16'd47863, 16'd33173, 16'd19938, 16'd23752, 16'd7025, 16'd13840, 16'd36589, 16'd49592, 16'd22413, 16'd23623});
	test_expansion(128'h6159c936834092b181c8f084ea040213, {16'd40836, 16'd30893, 16'd7927, 16'd41301, 16'd50059, 16'd2154, 16'd38055, 16'd32024, 16'd64551, 16'd9398, 16'd15306, 16'd19188, 16'd48567, 16'd35945, 16'd34220, 16'd9491, 16'd8645, 16'd54203, 16'd56118, 16'd31319, 16'd49421, 16'd28288, 16'd15560, 16'd21350, 16'd47077, 16'd46719});
	test_expansion(128'hab362e170a9ff9f2e0ed4b8c1dc569a5, {16'd63545, 16'd41190, 16'd64285, 16'd48311, 16'd19270, 16'd22931, 16'd52213, 16'd47926, 16'd36635, 16'd43963, 16'd15862, 16'd4640, 16'd40854, 16'd65023, 16'd24569, 16'd23272, 16'd3417, 16'd6574, 16'd6165, 16'd38837, 16'd20860, 16'd9925, 16'd49222, 16'd26124, 16'd42205, 16'd32481});
	test_expansion(128'h7b09ac1ae5795efd4b02d87a7b0233fd, {16'd29010, 16'd16966, 16'd28763, 16'd16435, 16'd30131, 16'd56418, 16'd1698, 16'd41079, 16'd7609, 16'd21810, 16'd24243, 16'd34753, 16'd16719, 16'd52178, 16'd62324, 16'd28981, 16'd1608, 16'd27865, 16'd34174, 16'd18572, 16'd4707, 16'd12025, 16'd55614, 16'd23481, 16'd32698, 16'd39728});
	test_expansion(128'h0aa96d436f8739230badf55d96396560, {16'd65448, 16'd60514, 16'd57597, 16'd33269, 16'd53182, 16'd24528, 16'd51067, 16'd7515, 16'd43412, 16'd63508, 16'd33870, 16'd10475, 16'd36536, 16'd60816, 16'd39930, 16'd33491, 16'd54998, 16'd6237, 16'd7564, 16'd15877, 16'd15567, 16'd5190, 16'd36292, 16'd4690, 16'd6303, 16'd33469});
	test_expansion(128'h4c77e9562e409767f019cff176d15c7e, {16'd10758, 16'd49978, 16'd52056, 16'd44335, 16'd45930, 16'd50991, 16'd39859, 16'd46859, 16'd12061, 16'd25422, 16'd4647, 16'd31161, 16'd32206, 16'd41737, 16'd34353, 16'd54307, 16'd37310, 16'd47820, 16'd15831, 16'd56774, 16'd8970, 16'd29971, 16'd52667, 16'd55845, 16'd32092, 16'd4409});
	test_expansion(128'h766f1b828a50a57604270b18435d9153, {16'd3608, 16'd9400, 16'd60036, 16'd64444, 16'd40947, 16'd51224, 16'd24439, 16'd63548, 16'd22659, 16'd14017, 16'd51037, 16'd52142, 16'd39019, 16'd38531, 16'd33348, 16'd39397, 16'd65530, 16'd54515, 16'd5361, 16'd39415, 16'd28530, 16'd32586, 16'd6461, 16'd44749, 16'd39768, 16'd27422});
	test_expansion(128'h96e1698832450afdecb9f600e985fae8, {16'd49516, 16'd44868, 16'd32570, 16'd2303, 16'd38881, 16'd43644, 16'd1030, 16'd44312, 16'd49458, 16'd9473, 16'd40525, 16'd36395, 16'd1638, 16'd50688, 16'd20701, 16'd18136, 16'd55998, 16'd7187, 16'd54037, 16'd55947, 16'd6757, 16'd47650, 16'd48304, 16'd9008, 16'd11183, 16'd44246});
	test_expansion(128'h1c33a74d071e680490cadebf6674918d, {16'd53633, 16'd15647, 16'd3285, 16'd32635, 16'd16924, 16'd20930, 16'd36663, 16'd7180, 16'd19810, 16'd15064, 16'd61400, 16'd60936, 16'd62496, 16'd55624, 16'd17702, 16'd27023, 16'd48023, 16'd54870, 16'd30253, 16'd27698, 16'd19654, 16'd19513, 16'd50972, 16'd55616, 16'd37056, 16'd27566});
	test_expansion(128'h02c2dfda152fb2c53a8f10c7bee68f8b, {16'd31351, 16'd31212, 16'd41538, 16'd43298, 16'd21080, 16'd46933, 16'd46174, 16'd55464, 16'd42828, 16'd49385, 16'd58269, 16'd62434, 16'd21870, 16'd62133, 16'd42872, 16'd35607, 16'd35826, 16'd58626, 16'd42185, 16'd17841, 16'd3750, 16'd31318, 16'd9492, 16'd48485, 16'd47074, 16'd45449});
	test_expansion(128'h38b2430c51f72b6aae9149f3e0f80b14, {16'd63478, 16'd3701, 16'd55473, 16'd54114, 16'd46260, 16'd27260, 16'd57281, 16'd22817, 16'd8941, 16'd543, 16'd19658, 16'd22115, 16'd35228, 16'd55022, 16'd6762, 16'd3391, 16'd205, 16'd35492, 16'd688, 16'd9972, 16'd31465, 16'd43467, 16'd11406, 16'd29101, 16'd5466, 16'd14056});
	test_expansion(128'h6f2dc3d2af3146bd3acc03c9a0974871, {16'd36562, 16'd2438, 16'd20205, 16'd10463, 16'd11250, 16'd13777, 16'd44740, 16'd61436, 16'd11700, 16'd57831, 16'd21878, 16'd41807, 16'd12448, 16'd56329, 16'd47056, 16'd16137, 16'd26711, 16'd9259, 16'd50237, 16'd24235, 16'd58212, 16'd33629, 16'd23445, 16'd31707, 16'd13833, 16'd54043});
	test_expansion(128'hba8ea7a72426d54aa77f26aa82453404, {16'd48469, 16'd4664, 16'd46356, 16'd42806, 16'd62232, 16'd62991, 16'd10860, 16'd5433, 16'd37429, 16'd25865, 16'd36982, 16'd29901, 16'd11189, 16'd45559, 16'd15342, 16'd3182, 16'd11341, 16'd47403, 16'd7879, 16'd32160, 16'd58280, 16'd29001, 16'd7988, 16'd4921, 16'd43742, 16'd43266});
	test_expansion(128'he95d5b20c3aa5e0b24b3e294300ef531, {16'd63057, 16'd1378, 16'd54084, 16'd53017, 16'd58940, 16'd51635, 16'd14566, 16'd13106, 16'd36179, 16'd40252, 16'd2044, 16'd56764, 16'd35592, 16'd39651, 16'd41309, 16'd39475, 16'd40203, 16'd65378, 16'd51667, 16'd39057, 16'd17413, 16'd23584, 16'd48732, 16'd10901, 16'd64280, 16'd33290});
	test_expansion(128'hbe56273b4d3be361f940ff4602fc7eec, {16'd289, 16'd51801, 16'd20827, 16'd15736, 16'd59675, 16'd25805, 16'd64149, 16'd63067, 16'd59876, 16'd60539, 16'd9989, 16'd17800, 16'd33098, 16'd26851, 16'd37198, 16'd63734, 16'd65258, 16'd25070, 16'd9986, 16'd33359, 16'd13581, 16'd1839, 16'd17213, 16'd11646, 16'd20724, 16'd32647});
	test_expansion(128'had1819649f3df208da0ce6a0b8ce310a, {16'd33894, 16'd25662, 16'd12560, 16'd45847, 16'd63119, 16'd47375, 16'd29425, 16'd37712, 16'd50504, 16'd28433, 16'd34224, 16'd951, 16'd18519, 16'd26755, 16'd33166, 16'd18235, 16'd49276, 16'd26629, 16'd40800, 16'd34477, 16'd23689, 16'd17621, 16'd6025, 16'd50945, 16'd50878, 16'd15645});
	test_expansion(128'h49ecbc78c1dc2b784080f12e8f7b0257, {16'd34778, 16'd38236, 16'd11168, 16'd35570, 16'd24437, 16'd38928, 16'd18414, 16'd51328, 16'd34442, 16'd28451, 16'd10375, 16'd8322, 16'd24741, 16'd46727, 16'd23310, 16'd28705, 16'd7587, 16'd53727, 16'd43896, 16'd32501, 16'd34455, 16'd11599, 16'd10566, 16'd44628, 16'd49042, 16'd25820});
	test_expansion(128'h5d7beb6d8d7f79b2a387a13ab70986d7, {16'd13233, 16'd55792, 16'd26217, 16'd8614, 16'd6945, 16'd18663, 16'd26332, 16'd33054, 16'd49670, 16'd14249, 16'd43446, 16'd33687, 16'd25158, 16'd50446, 16'd3520, 16'd3843, 16'd3941, 16'd23827, 16'd18484, 16'd45527, 16'd52, 16'd48122, 16'd15202, 16'd35599, 16'd19147, 16'd30283});
	test_expansion(128'h5fd8082c1856551b64e352d4994206b9, {16'd65133, 16'd38535, 16'd47147, 16'd16504, 16'd45948, 16'd4764, 16'd15749, 16'd48130, 16'd25189, 16'd9109, 16'd28586, 16'd34781, 16'd48610, 16'd7039, 16'd40893, 16'd14079, 16'd39464, 16'd24277, 16'd48950, 16'd61105, 16'd1718, 16'd2212, 16'd3352, 16'd7486, 16'd52920, 16'd18377});
	test_expansion(128'h5efa3be7356f4da2d10b1f61dfbcb6c5, {16'd2124, 16'd48368, 16'd41798, 16'd17559, 16'd28812, 16'd24654, 16'd65084, 16'd28757, 16'd8630, 16'd9478, 16'd44253, 16'd53519, 16'd49626, 16'd65453, 16'd31206, 16'd47279, 16'd39407, 16'd57644, 16'd23419, 16'd37097, 16'd43825, 16'd64732, 16'd44164, 16'd23510, 16'd22744, 16'd37305});
	test_expansion(128'h5d1e50e6b1da99463edbf9226cd65d4a, {16'd46873, 16'd55387, 16'd20009, 16'd779, 16'd7177, 16'd46096, 16'd1954, 16'd49757, 16'd46227, 16'd5726, 16'd35411, 16'd3670, 16'd37035, 16'd33806, 16'd56002, 16'd23915, 16'd63985, 16'd54854, 16'd43094, 16'd41741, 16'd49753, 16'd32053, 16'd2407, 16'd37375, 16'd28033, 16'd20667});
	test_expansion(128'ha0078f536534324a7a1934fc8431187d, {16'd22349, 16'd411, 16'd42821, 16'd23865, 16'd32546, 16'd36653, 16'd22695, 16'd26824, 16'd22321, 16'd4614, 16'd3726, 16'd210, 16'd11696, 16'd6462, 16'd18370, 16'd65462, 16'd27720, 16'd20138, 16'd54547, 16'd52404, 16'd47396, 16'd11190, 16'd18484, 16'd9082, 16'd59632, 16'd33433});
	test_expansion(128'h3ca630e24ab8709c9f8a61a16d686215, {16'd4895, 16'd54933, 16'd19880, 16'd50229, 16'd43985, 16'd13859, 16'd18496, 16'd187, 16'd41630, 16'd4021, 16'd62754, 16'd45779, 16'd35673, 16'd57446, 16'd19116, 16'd38927, 16'd24921, 16'd2646, 16'd1581, 16'd11104, 16'd100, 16'd14931, 16'd26894, 16'd59102, 16'd17829, 16'd34763});
	test_expansion(128'ha1429c03a40caf15b8f731f664fe24ce, {16'd14493, 16'd61366, 16'd57129, 16'd48071, 16'd61356, 16'd42028, 16'd29018, 16'd8634, 16'd34928, 16'd36826, 16'd2671, 16'd56874, 16'd53523, 16'd17470, 16'd23542, 16'd39504, 16'd12727, 16'd13245, 16'd14370, 16'd39080, 16'd4542, 16'd25102, 16'd19539, 16'd7128, 16'd6209, 16'd2613});
	test_expansion(128'hdf447333e739db9093e3e6dea44fd8b5, {16'd12221, 16'd10158, 16'd34366, 16'd44243, 16'd5067, 16'd6493, 16'd28510, 16'd33175, 16'd52453, 16'd44972, 16'd58684, 16'd17306, 16'd52649, 16'd59958, 16'd40339, 16'd318, 16'd23749, 16'd21055, 16'd9940, 16'd29566, 16'd19556, 16'd45477, 16'd33868, 16'd50811, 16'd51049, 16'd5901});
	test_expansion(128'h91f26868ba2dc9ce42513bb4e00910ce, {16'd20050, 16'd22724, 16'd18401, 16'd36199, 16'd4862, 16'd55615, 16'd33817, 16'd28541, 16'd55002, 16'd51343, 16'd57824, 16'd26584, 16'd23570, 16'd49083, 16'd40181, 16'd1141, 16'd53260, 16'd26914, 16'd50218, 16'd64754, 16'd39825, 16'd20358, 16'd61344, 16'd15706, 16'd36977, 16'd49710});
	test_expansion(128'hd89634ec985ae1f9e4d3642494aa8aed, {16'd10788, 16'd32837, 16'd19099, 16'd59966, 16'd26625, 16'd49708, 16'd14837, 16'd21169, 16'd12958, 16'd30382, 16'd29292, 16'd54149, 16'd15206, 16'd21619, 16'd34628, 16'd11021, 16'd45649, 16'd55772, 16'd19067, 16'd18160, 16'd25649, 16'd59318, 16'd34951, 16'd42086, 16'd31098, 16'd29446});
	test_expansion(128'hbd46309a89db376bacff77687e84b52a, {16'd34911, 16'd20054, 16'd35405, 16'd46484, 16'd61083, 16'd29787, 16'd26852, 16'd26698, 16'd51382, 16'd54217, 16'd46883, 16'd44594, 16'd17404, 16'd44746, 16'd17148, 16'd8980, 16'd20773, 16'd23252, 16'd51818, 16'd44749, 16'd65510, 16'd16302, 16'd57392, 16'd60051, 16'd49722, 16'd36241});
	test_expansion(128'hd1e1876d4de3d64fdb068f8a2432cdfc, {16'd9819, 16'd18098, 16'd62231, 16'd50204, 16'd10784, 16'd46431, 16'd36594, 16'd16590, 16'd26569, 16'd53668, 16'd58170, 16'd11708, 16'd34647, 16'd20728, 16'd23918, 16'd10018, 16'd2381, 16'd47741, 16'd45036, 16'd14280, 16'd55008, 16'd28317, 16'd25547, 16'd8551, 16'd14672, 16'd49146});
	test_expansion(128'h1d273d108cf1af340d14f542d192ba73, {16'd30308, 16'd56669, 16'd41457, 16'd32877, 16'd29205, 16'd58879, 16'd46101, 16'd59188, 16'd32565, 16'd56222, 16'd22787, 16'd55957, 16'd3781, 16'd11009, 16'd7059, 16'd20769, 16'd43542, 16'd14135, 16'd15068, 16'd52551, 16'd38747, 16'd45997, 16'd7260, 16'd17430, 16'd51467, 16'd52163});
	test_expansion(128'h531d487d70d265217ff0d665f825bc76, {16'd55314, 16'd39978, 16'd20798, 16'd22833, 16'd738, 16'd44769, 16'd57686, 16'd61875, 16'd14872, 16'd57928, 16'd9309, 16'd33546, 16'd49023, 16'd20920, 16'd3835, 16'd40654, 16'd37110, 16'd44654, 16'd28298, 16'd1986, 16'd26471, 16'd36354, 16'd35662, 16'd17828, 16'd52754, 16'd12250});
	test_expansion(128'h54ccdb7d76a66b538f7b42bdf0bd376b, {16'd57529, 16'd20650, 16'd34755, 16'd16017, 16'd10068, 16'd8454, 16'd51541, 16'd7098, 16'd17710, 16'd43905, 16'd25523, 16'd53457, 16'd22442, 16'd32967, 16'd1753, 16'd6534, 16'd27893, 16'd20358, 16'd48103, 16'd9259, 16'd12521, 16'd710, 16'd63462, 16'd4703, 16'd17384, 16'd31548});
	test_expansion(128'h58f021f3ac50d58d71578dce876cc328, {16'd51005, 16'd8010, 16'd28997, 16'd3625, 16'd50701, 16'd20669, 16'd23183, 16'd62676, 16'd47569, 16'd19184, 16'd11072, 16'd44795, 16'd28288, 16'd39720, 16'd7955, 16'd29664, 16'd53663, 16'd25398, 16'd43413, 16'd60953, 16'd38904, 16'd43855, 16'd27648, 16'd28270, 16'd6681, 16'd16920});
	test_expansion(128'hafac945693a21314f8b78c8d9cb42f66, {16'd15699, 16'd51946, 16'd28340, 16'd22878, 16'd32800, 16'd57162, 16'd9250, 16'd46969, 16'd20446, 16'd50980, 16'd9523, 16'd49573, 16'd19447, 16'd47806, 16'd38853, 16'd64715, 16'd22444, 16'd55955, 16'd23239, 16'd1546, 16'd12634, 16'd13782, 16'd55371, 16'd12076, 16'd65090, 16'd5204});
	test_expansion(128'h34a574ff68f0b2deb2d62d1a2eee92dc, {16'd47784, 16'd26186, 16'd26382, 16'd45065, 16'd27012, 16'd48102, 16'd10533, 16'd6743, 16'd23600, 16'd34230, 16'd39824, 16'd54815, 16'd19802, 16'd65313, 16'd3264, 16'd60422, 16'd37251, 16'd40829, 16'd25922, 16'd47732, 16'd39214, 16'd34430, 16'd59486, 16'd59217, 16'd42077, 16'd35996});
	test_expansion(128'h887024b796284e795bf2c87b8783e6ea, {16'd49317, 16'd31537, 16'd41671, 16'd54221, 16'd43524, 16'd39532, 16'd26259, 16'd39236, 16'd53016, 16'd32647, 16'd3742, 16'd56985, 16'd9813, 16'd4012, 16'd47082, 16'd21790, 16'd14645, 16'd27345, 16'd56348, 16'd63485, 16'd16135, 16'd1250, 16'd6366, 16'd14016, 16'd48990, 16'd53137});
	test_expansion(128'h2cbd5c1fae6d30b9e74250d8933927b2, {16'd848, 16'd36115, 16'd23350, 16'd58320, 16'd50997, 16'd38253, 16'd64492, 16'd20909, 16'd58867, 16'd50333, 16'd64339, 16'd53084, 16'd3854, 16'd32440, 16'd43521, 16'd57422, 16'd57352, 16'd65437, 16'd63021, 16'd6667, 16'd36325, 16'd34213, 16'd35305, 16'd24675, 16'd6216, 16'd63279});
	test_expansion(128'he664921798614be54801317f2d60095b, {16'd33369, 16'd33981, 16'd6871, 16'd1446, 16'd18912, 16'd64747, 16'd18590, 16'd15464, 16'd21196, 16'd8237, 16'd19431, 16'd30522, 16'd37691, 16'd14751, 16'd37168, 16'd162, 16'd31891, 16'd8042, 16'd10068, 16'd26410, 16'd4957, 16'd13241, 16'd51453, 16'd9696, 16'd47563, 16'd46558});
	test_expansion(128'h0fd3e915cc98dce6589fe000846c730a, {16'd24272, 16'd38016, 16'd37055, 16'd50066, 16'd5351, 16'd43490, 16'd59005, 16'd14330, 16'd27926, 16'd41761, 16'd8190, 16'd61101, 16'd35319, 16'd46103, 16'd53958, 16'd38575, 16'd14545, 16'd7103, 16'd45520, 16'd41622, 16'd17558, 16'd6749, 16'd3176, 16'd37855, 16'd53068, 16'd20844});
	test_expansion(128'h215ad8bb559b0bfed4a9e547af4724c6, {16'd37557, 16'd52636, 16'd13075, 16'd3822, 16'd6844, 16'd36568, 16'd23142, 16'd5601, 16'd1618, 16'd49437, 16'd62939, 16'd35592, 16'd59186, 16'd51432, 16'd62228, 16'd58561, 16'd31286, 16'd18255, 16'd42837, 16'd42383, 16'd17636, 16'd1806, 16'd45518, 16'd57881, 16'd37631, 16'd19438});
	test_expansion(128'h70f09dd608a4585f443e110b61a6978c, {16'd63604, 16'd65125, 16'd51148, 16'd26639, 16'd2853, 16'd53409, 16'd8134, 16'd22626, 16'd62082, 16'd52034, 16'd62923, 16'd2647, 16'd29198, 16'd36567, 16'd37681, 16'd35598, 16'd3820, 16'd60112, 16'd36730, 16'd36074, 16'd34203, 16'd43071, 16'd28721, 16'd52709, 16'd29988, 16'd22031});
	test_expansion(128'h3e43d38cef856d7d6a7cc4fd595f0c01, {16'd9230, 16'd50674, 16'd60222, 16'd40163, 16'd29475, 16'd49411, 16'd287, 16'd24611, 16'd36671, 16'd14568, 16'd51612, 16'd22026, 16'd30204, 16'd11093, 16'd57980, 16'd54314, 16'd52600, 16'd19775, 16'd47884, 16'd45377, 16'd35362, 16'd60548, 16'd41272, 16'd35814, 16'd44243, 16'd22927});
	test_expansion(128'h86f7ec02d983354b1dd388ebff627f8d, {16'd31148, 16'd3772, 16'd49288, 16'd51524, 16'd32346, 16'd30494, 16'd49951, 16'd34494, 16'd44765, 16'd1973, 16'd55349, 16'd52605, 16'd57216, 16'd56510, 16'd3970, 16'd57484, 16'd29244, 16'd40078, 16'd624, 16'd41966, 16'd25488, 16'd61194, 16'd63038, 16'd39956, 16'd27030, 16'd591});
	test_expansion(128'h4ba93701347616d89343344732b81a66, {16'd21626, 16'd29762, 16'd56621, 16'd39312, 16'd58808, 16'd44969, 16'd48934, 16'd62731, 16'd49096, 16'd10468, 16'd32998, 16'd15089, 16'd9586, 16'd16594, 16'd18305, 16'd2080, 16'd51533, 16'd32404, 16'd27127, 16'd33510, 16'd39737, 16'd27644, 16'd57729, 16'd5936, 16'd19216, 16'd30385});
	test_expansion(128'h488f104c0bfe41b4b2d238b5eb44e690, {16'd64643, 16'd17938, 16'd5603, 16'd39038, 16'd47559, 16'd50341, 16'd6529, 16'd52808, 16'd46865, 16'd56899, 16'd65327, 16'd17050, 16'd62664, 16'd27462, 16'd14878, 16'd42377, 16'd64558, 16'd64521, 16'd19486, 16'd64358, 16'd55409, 16'd31956, 16'd44883, 16'd51520, 16'd30809, 16'd32383});
	test_expansion(128'h3395d69ca21462edb25fd18843b3a3bb, {16'd4457, 16'd7368, 16'd59615, 16'd27687, 16'd39849, 16'd29581, 16'd22869, 16'd33981, 16'd40233, 16'd26721, 16'd19444, 16'd65279, 16'd4168, 16'd38448, 16'd39639, 16'd60775, 16'd22805, 16'd58145, 16'd58791, 16'd2703, 16'd47638, 16'd30028, 16'd7649, 16'd54694, 16'd12646, 16'd1153});
	test_expansion(128'hff31583c6f0a0c402cd9ffaba1db7100, {16'd47070, 16'd8671, 16'd4726, 16'd26456, 16'd14839, 16'd64169, 16'd59718, 16'd57135, 16'd23622, 16'd46142, 16'd64851, 16'd45271, 16'd27853, 16'd2749, 16'd32514, 16'd33875, 16'd22989, 16'd47890, 16'd65200, 16'd34806, 16'd42222, 16'd2820, 16'd43421, 16'd52607, 16'd64982, 16'd22653});
	test_expansion(128'h6ca315f20de9c76ad55c8c5641d8e3f5, {16'd24403, 16'd14655, 16'd18106, 16'd40422, 16'd13168, 16'd65019, 16'd37310, 16'd56119, 16'd47203, 16'd42058, 16'd40406, 16'd5118, 16'd5873, 16'd419, 16'd15046, 16'd11494, 16'd31967, 16'd22357, 16'd3559, 16'd9152, 16'd39993, 16'd17826, 16'd41799, 16'd39574, 16'd60248, 16'd63247});
	test_expansion(128'h133cb43de39c5b6e2afbb02e3ce8703d, {16'd61142, 16'd26952, 16'd19492, 16'd54852, 16'd18190, 16'd4943, 16'd30076, 16'd5840, 16'd21952, 16'd44267, 16'd29296, 16'd676, 16'd8714, 16'd36708, 16'd9345, 16'd6655, 16'd35181, 16'd54607, 16'd35429, 16'd37805, 16'd26174, 16'd19480, 16'd26113, 16'd19112, 16'd57564, 16'd41022});
	test_expansion(128'h2005936ab8105d64ec6d443bccca08ba, {16'd28220, 16'd15704, 16'd59332, 16'd41921, 16'd15474, 16'd40166, 16'd6258, 16'd41378, 16'd9338, 16'd8655, 16'd3531, 16'd57606, 16'd59866, 16'd51095, 16'd53363, 16'd3783, 16'd31237, 16'd1379, 16'd50622, 16'd27477, 16'd23681, 16'd50371, 16'd39359, 16'd38921, 16'd30014, 16'd51432});
	test_expansion(128'hdd254df9bcfbc448979c6f1f3583e8f1, {16'd11521, 16'd12728, 16'd17268, 16'd24339, 16'd53549, 16'd10468, 16'd56639, 16'd5758, 16'd39598, 16'd58265, 16'd30171, 16'd18812, 16'd34873, 16'd517, 16'd56184, 16'd64403, 16'd21415, 16'd29523, 16'd23084, 16'd10978, 16'd41332, 16'd65, 16'd26796, 16'd55376, 16'd16857, 16'd54313});
	test_expansion(128'hccac848c1df2b873c8ccae718367ec1d, {16'd28573, 16'd8419, 16'd5978, 16'd19474, 16'd54342, 16'd64340, 16'd58340, 16'd4801, 16'd42938, 16'd16245, 16'd44580, 16'd53354, 16'd16007, 16'd33790, 16'd6680, 16'd20551, 16'd51241, 16'd57517, 16'd31289, 16'd44599, 16'd5452, 16'd21315, 16'd60396, 16'd11274, 16'd2007, 16'd50623});
	test_expansion(128'habc4e4c9d5ccf5c8d9128d3199ec7d04, {16'd25519, 16'd41754, 16'd60171, 16'd42972, 16'd62214, 16'd11377, 16'd33067, 16'd65025, 16'd31653, 16'd42370, 16'd48620, 16'd34129, 16'd13797, 16'd22011, 16'd38869, 16'd8359, 16'd16186, 16'd9274, 16'd3368, 16'd35512, 16'd19178, 16'd50497, 16'd50289, 16'd51250, 16'd42708, 16'd8348});
	test_expansion(128'hd1542ee3c617f1f821ee096b203f608a, {16'd2833, 16'd55087, 16'd64524, 16'd32426, 16'd63614, 16'd41703, 16'd64193, 16'd41865, 16'd64398, 16'd45026, 16'd24846, 16'd23680, 16'd58236, 16'd13205, 16'd5688, 16'd56524, 16'd55922, 16'd3123, 16'd54387, 16'd55393, 16'd31426, 16'd60345, 16'd10199, 16'd1732, 16'd46541, 16'd29250});
	test_expansion(128'hcbca8d5aa80543a55d2b2ff223258105, {16'd39417, 16'd10259, 16'd10184, 16'd11898, 16'd30982, 16'd50432, 16'd22023, 16'd1010, 16'd41844, 16'd32091, 16'd404, 16'd25083, 16'd28281, 16'd1759, 16'd45090, 16'd53240, 16'd26467, 16'd1418, 16'd43657, 16'd55846, 16'd36695, 16'd11058, 16'd12855, 16'd7390, 16'd51624, 16'd24454});
	test_expansion(128'h770980a1069d76c23cb1478c5b7f5e69, {16'd51184, 16'd33988, 16'd53801, 16'd43254, 16'd15965, 16'd9460, 16'd53222, 16'd28121, 16'd24810, 16'd18215, 16'd22156, 16'd29719, 16'd54220, 16'd4797, 16'd40384, 16'd11406, 16'd34765, 16'd62004, 16'd50886, 16'd6728, 16'd17184, 16'd17066, 16'd36009, 16'd62887, 16'd63355, 16'd62462});
	test_expansion(128'h5a8bbcc23229c14d4ce656aae6a3a21e, {16'd51101, 16'd39207, 16'd49239, 16'd26594, 16'd8736, 16'd600, 16'd47159, 16'd54174, 16'd10619, 16'd58247, 16'd24460, 16'd7764, 16'd1794, 16'd15537, 16'd64448, 16'd41351, 16'd6945, 16'd43711, 16'd38640, 16'd39241, 16'd58278, 16'd39294, 16'd62701, 16'd4106, 16'd29188, 16'd40323});
	test_expansion(128'he27db1d3e4c9bb3ca54336975537af5c, {16'd42411, 16'd16599, 16'd37314, 16'd9746, 16'd44629, 16'd62056, 16'd13232, 16'd18071, 16'd35978, 16'd39230, 16'd9121, 16'd48778, 16'd10429, 16'd26659, 16'd10983, 16'd10400, 16'd12854, 16'd44627, 16'd1943, 16'd46147, 16'd32790, 16'd20583, 16'd48875, 16'd62182, 16'd46732, 16'd58170});
	test_expansion(128'h1f9179145e1eb2baa0fe3e1d1690d34c, {16'd28654, 16'd31676, 16'd64102, 16'd33871, 16'd56472, 16'd49570, 16'd12217, 16'd33916, 16'd16654, 16'd10012, 16'd550, 16'd20426, 16'd45895, 16'd17520, 16'd2472, 16'd36247, 16'd773, 16'd4544, 16'd31178, 16'd7826, 16'd31351, 16'd29784, 16'd39243, 16'd9974, 16'd33032, 16'd45983});
	test_expansion(128'hd72b111220f8789cc1d64960be38cb02, {16'd19902, 16'd9921, 16'd26226, 16'd40352, 16'd45928, 16'd917, 16'd56541, 16'd50001, 16'd34867, 16'd10490, 16'd24527, 16'd16464, 16'd24843, 16'd54194, 16'd30203, 16'd47932, 16'd2766, 16'd15378, 16'd5183, 16'd23530, 16'd26753, 16'd2254, 16'd35541, 16'd22967, 16'd7000, 16'd50495});
	test_expansion(128'h4ec79c887829124d2f06ce548d7f44af, {16'd42939, 16'd37765, 16'd27503, 16'd23723, 16'd14582, 16'd63731, 16'd16771, 16'd37335, 16'd29609, 16'd8100, 16'd47932, 16'd65061, 16'd37741, 16'd10297, 16'd27437, 16'd14131, 16'd46319, 16'd65129, 16'd54006, 16'd14823, 16'd43982, 16'd27948, 16'd16334, 16'd43053, 16'd5973, 16'd31333});
	test_expansion(128'h0493efbdc083aa396e063322d0d07b85, {16'd21857, 16'd39146, 16'd39795, 16'd42622, 16'd35313, 16'd6335, 16'd15106, 16'd52892, 16'd53975, 16'd19571, 16'd49144, 16'd39386, 16'd52513, 16'd37630, 16'd51004, 16'd54496, 16'd58231, 16'd27334, 16'd57962, 16'd46489, 16'd40569, 16'd35526, 16'd22499, 16'd39058, 16'd16079, 16'd13604});
	test_expansion(128'hc4316ea4b83b5958beead71468a1ee13, {16'd26133, 16'd22369, 16'd37260, 16'd56161, 16'd35032, 16'd56057, 16'd25540, 16'd59971, 16'd27277, 16'd21960, 16'd26165, 16'd8563, 16'd60987, 16'd30503, 16'd4925, 16'd7000, 16'd18705, 16'd27082, 16'd38258, 16'd18756, 16'd2373, 16'd42122, 16'd36448, 16'd29477, 16'd45058, 16'd4728});
	test_expansion(128'h7fb31e643c3c1597e0b2fe7de7fa585f, {16'd7980, 16'd38154, 16'd8030, 16'd40145, 16'd31072, 16'd9959, 16'd61688, 16'd6677, 16'd36652, 16'd39297, 16'd11914, 16'd17158, 16'd35623, 16'd10117, 16'd181, 16'd23110, 16'd34704, 16'd25965, 16'd2892, 16'd60183, 16'd55916, 16'd3240, 16'd5529, 16'd44132, 16'd21310, 16'd39199});
	test_expansion(128'h7adc7250081c50bdc7015454261be155, {16'd32396, 16'd12611, 16'd55386, 16'd18653, 16'd35385, 16'd47394, 16'd60889, 16'd26561, 16'd1600, 16'd51241, 16'd54161, 16'd26954, 16'd36236, 16'd56293, 16'd18483, 16'd27641, 16'd37847, 16'd13066, 16'd31388, 16'd61923, 16'd1753, 16'd36196, 16'd27943, 16'd11126, 16'd859, 16'd3808});
	test_expansion(128'h5ce4f8e78f9359ea3411a2bb721fa7fb, {16'd63429, 16'd13499, 16'd42417, 16'd41359, 16'd14933, 16'd63213, 16'd51521, 16'd56264, 16'd35652, 16'd60351, 16'd19959, 16'd37429, 16'd55294, 16'd21457, 16'd24666, 16'd10527, 16'd41778, 16'd63242, 16'd17148, 16'd34707, 16'd13726, 16'd16615, 16'd62168, 16'd8802, 16'd31744, 16'd22974});
	test_expansion(128'h34c466f9ea44b1e3e242f8c82fc0f156, {16'd21172, 16'd47798, 16'd8703, 16'd17858, 16'd36997, 16'd28420, 16'd56242, 16'd21575, 16'd47183, 16'd34900, 16'd35453, 16'd40945, 16'd42707, 16'd19744, 16'd15801, 16'd2240, 16'd54180, 16'd51370, 16'd24080, 16'd12991, 16'd3226, 16'd4133, 16'd15351, 16'd12859, 16'd27699, 16'd52532});
	test_expansion(128'hc28b2549893b7f8e71afcdf82d08a480, {16'd28146, 16'd50161, 16'd55355, 16'd59664, 16'd16605, 16'd41417, 16'd40188, 16'd16870, 16'd59640, 16'd53444, 16'd36405, 16'd29622, 16'd1670, 16'd37427, 16'd14388, 16'd20175, 16'd37344, 16'd50112, 16'd28779, 16'd21972, 16'd50683, 16'd44076, 16'd9394, 16'd8650, 16'd44442, 16'd16361});
	test_expansion(128'hb6eb7a58a7a096c95ff9f65e03171f6a, {16'd8092, 16'd19384, 16'd60123, 16'd27133, 16'd48658, 16'd39578, 16'd50338, 16'd26603, 16'd24630, 16'd2911, 16'd10927, 16'd26136, 16'd19256, 16'd55689, 16'd19875, 16'd740, 16'd49216, 16'd19084, 16'd56524, 16'd10549, 16'd22687, 16'd11917, 16'd25056, 16'd1266, 16'd36326, 16'd30765});
	test_expansion(128'h16f0939459acd9026808c558c7e671b3, {16'd61017, 16'd7813, 16'd20212, 16'd59621, 16'd32415, 16'd14727, 16'd1113, 16'd52067, 16'd32162, 16'd9457, 16'd59240, 16'd57393, 16'd10553, 16'd50996, 16'd51931, 16'd9501, 16'd523, 16'd33828, 16'd55868, 16'd21357, 16'd26524, 16'd55524, 16'd21441, 16'd42340, 16'd26195, 16'd1467});
	test_expansion(128'h0738cbf6e95b840524f96b34ae0307e1, {16'd4376, 16'd60861, 16'd52170, 16'd4604, 16'd23870, 16'd45213, 16'd14995, 16'd21960, 16'd45341, 16'd33722, 16'd7223, 16'd35127, 16'd325, 16'd41483, 16'd36365, 16'd52551, 16'd31958, 16'd18120, 16'd11444, 16'd42203, 16'd55150, 16'd31327, 16'd63575, 16'd25601, 16'd50944, 16'd33936});
	test_expansion(128'h06f1226924a5dd24c6a117d2b6f4f71a, {16'd37642, 16'd47686, 16'd1227, 16'd44641, 16'd2331, 16'd28827, 16'd42706, 16'd46693, 16'd30126, 16'd47129, 16'd38980, 16'd61655, 16'd61539, 16'd59055, 16'd27940, 16'd13495, 16'd35841, 16'd53774, 16'd27139, 16'd15444, 16'd46333, 16'd43675, 16'd56304, 16'd62958, 16'd12046, 16'd39016});
	test_expansion(128'h35be0cb846eb005e35b595408e88b050, {16'd13206, 16'd43211, 16'd35890, 16'd52406, 16'd36610, 16'd47774, 16'd22723, 16'd54551, 16'd16146, 16'd46875, 16'd56133, 16'd37758, 16'd44672, 16'd43508, 16'd33680, 16'd60709, 16'd13685, 16'd52607, 16'd49930, 16'd41116, 16'd44671, 16'd54954, 16'd10343, 16'd3174, 16'd10386, 16'd33540});
	test_expansion(128'h2fdfffcb74381188db49b1dcab518800, {16'd41884, 16'd34629, 16'd28800, 16'd30628, 16'd31221, 16'd51360, 16'd50551, 16'd30462, 16'd48196, 16'd24869, 16'd22222, 16'd56852, 16'd48860, 16'd28208, 16'd760, 16'd43748, 16'd30248, 16'd37215, 16'd5751, 16'd1689, 16'd51617, 16'd17010, 16'd47451, 16'd30537, 16'd41522, 16'd43103});
	test_expansion(128'h8feafb73b6d1247bddf15194f572186b, {16'd30422, 16'd51362, 16'd63066, 16'd96, 16'd42725, 16'd26314, 16'd9869, 16'd49128, 16'd34060, 16'd57599, 16'd53223, 16'd16629, 16'd57541, 16'd44074, 16'd53208, 16'd40449, 16'd42308, 16'd54037, 16'd39348, 16'd7918, 16'd21557, 16'd9727, 16'd43626, 16'd46335, 16'd60242, 16'd49911});
	test_expansion(128'hfa81f91f226ba3b0c5a38bfcec593d5c, {16'd24921, 16'd61769, 16'd9220, 16'd2093, 16'd15340, 16'd23277, 16'd20101, 16'd43949, 16'd40274, 16'd33754, 16'd385, 16'd24125, 16'd32799, 16'd64270, 16'd42875, 16'd47931, 16'd13223, 16'd62983, 16'd42937, 16'd21339, 16'd20811, 16'd48024, 16'd12441, 16'd1349, 16'd13610, 16'd11899});
	test_expansion(128'h07c9c0bf14854c868f289d0750a15ee2, {16'd9796, 16'd7752, 16'd59296, 16'd29009, 16'd28954, 16'd58625, 16'd40535, 16'd8481, 16'd4298, 16'd40240, 16'd8887, 16'd6087, 16'd25434, 16'd25738, 16'd40027, 16'd39923, 16'd29334, 16'd45497, 16'd2072, 16'd14392, 16'd13841, 16'd3595, 16'd63166, 16'd49918, 16'd45103, 16'd28455});
	test_expansion(128'h506bc5ffda61d05b022f112bfe2a5385, {16'd19175, 16'd41337, 16'd34302, 16'd59994, 16'd34134, 16'd34858, 16'd63837, 16'd33047, 16'd34621, 16'd50840, 16'd58885, 16'd44519, 16'd62121, 16'd11377, 16'd30433, 16'd13490, 16'd698, 16'd35776, 16'd57352, 16'd48651, 16'd14748, 16'd10581, 16'd24819, 16'd34416, 16'd20043, 16'd31852});
	test_expansion(128'h3b5861a092c88dc4243ebcd2d52bf09f, {16'd23379, 16'd1201, 16'd47540, 16'd13775, 16'd53829, 16'd25975, 16'd6080, 16'd6688, 16'd16070, 16'd65217, 16'd10163, 16'd39478, 16'd57458, 16'd40880, 16'd35237, 16'd27159, 16'd14359, 16'd14997, 16'd55222, 16'd49223, 16'd42838, 16'd8580, 16'd62533, 16'd34648, 16'd61543, 16'd4060});
	test_expansion(128'hb3158336371c4864f86cefd378c4e011, {16'd17029, 16'd48328, 16'd28864, 16'd62333, 16'd30715, 16'd15245, 16'd11594, 16'd38022, 16'd11069, 16'd28460, 16'd50225, 16'd25494, 16'd63054, 16'd50375, 16'd32561, 16'd1566, 16'd46710, 16'd37808, 16'd41864, 16'd19425, 16'd64426, 16'd17342, 16'd19245, 16'd46067, 16'd29703, 16'd34645});
	test_expansion(128'hf0e468b7dcb2144daad7c1c920db5d32, {16'd44715, 16'd10064, 16'd60560, 16'd61764, 16'd41572, 16'd3242, 16'd46408, 16'd17934, 16'd10185, 16'd12837, 16'd41520, 16'd6024, 16'd31392, 16'd22063, 16'd35562, 16'd18465, 16'd30575, 16'd31153, 16'd26004, 16'd59264, 16'd32262, 16'd32325, 16'd37037, 16'd37570, 16'd2086, 16'd47532});
	test_expansion(128'hbf6731e1867d70c425bc2b82a1da319b, {16'd63982, 16'd36140, 16'd56047, 16'd6970, 16'd7023, 16'd47447, 16'd750, 16'd19554, 16'd25234, 16'd22808, 16'd24618, 16'd39559, 16'd62886, 16'd41143, 16'd1403, 16'd32174, 16'd14817, 16'd29573, 16'd25030, 16'd25281, 16'd57601, 16'd12621, 16'd51939, 16'd58190, 16'd48696, 16'd10316});
	test_expansion(128'h915dd34e812b2720495cbed402129a0b, {16'd60937, 16'd10171, 16'd25635, 16'd54251, 16'd4613, 16'd60628, 16'd17512, 16'd36307, 16'd36690, 16'd48658, 16'd14024, 16'd29584, 16'd21980, 16'd33124, 16'd10057, 16'd56003, 16'd40781, 16'd14441, 16'd30171, 16'd46016, 16'd12091, 16'd14589, 16'd20756, 16'd1974, 16'd9466, 16'd58481});
	test_expansion(128'hcf7828e1d3bb5fbc32124468044ba580, {16'd1744, 16'd9371, 16'd10902, 16'd1483, 16'd50866, 16'd28287, 16'd1645, 16'd21766, 16'd58604, 16'd63210, 16'd44128, 16'd8416, 16'd47647, 16'd53789, 16'd50490, 16'd45760, 16'd11645, 16'd45365, 16'd11635, 16'd39020, 16'd60897, 16'd25291, 16'd58038, 16'd52658, 16'd43156, 16'd37229});
	test_expansion(128'hb25211927e1ff3b3c367c93c963e28f9, {16'd64445, 16'd2899, 16'd9249, 16'd58018, 16'd35859, 16'd54728, 16'd22542, 16'd48394, 16'd18838, 16'd49221, 16'd65412, 16'd43497, 16'd32452, 16'd43707, 16'd15543, 16'd39685, 16'd29350, 16'd25484, 16'd41245, 16'd40255, 16'd19396, 16'd5959, 16'd5642, 16'd610, 16'd48656, 16'd20901});
	test_expansion(128'h96e4ed6423313122345258edf7b2d4a6, {16'd8138, 16'd54679, 16'd8906, 16'd63905, 16'd9074, 16'd54, 16'd4071, 16'd19282, 16'd57634, 16'd47287, 16'd64154, 16'd39595, 16'd35108, 16'd58229, 16'd59345, 16'd46713, 16'd44417, 16'd9037, 16'd31922, 16'd54917, 16'd60571, 16'd28173, 16'd41309, 16'd14618, 16'd22849, 16'd55775});
	test_expansion(128'h0497f26052848f8a2812909d73350588, {16'd39654, 16'd56551, 16'd37829, 16'd60432, 16'd48632, 16'd22804, 16'd54934, 16'd57682, 16'd39285, 16'd48422, 16'd55591, 16'd18804, 16'd43590, 16'd43030, 16'd4186, 16'd22882, 16'd44324, 16'd15551, 16'd61586, 16'd46051, 16'd18736, 16'd23177, 16'd39615, 16'd50040, 16'd12548, 16'd59213});
	test_expansion(128'h75a653bf7c7917a709e9ed9f3dbe34ab, {16'd12690, 16'd59546, 16'd25983, 16'd5278, 16'd9551, 16'd63234, 16'd55077, 16'd18604, 16'd9541, 16'd46815, 16'd4874, 16'd52151, 16'd31498, 16'd65301, 16'd50622, 16'd64993, 16'd46886, 16'd2025, 16'd26047, 16'd23686, 16'd48588, 16'd30494, 16'd51978, 16'd51401, 16'd9397, 16'd34740});
	test_expansion(128'h3c59e35697a772e949b8b3e2ff801adb, {16'd11206, 16'd23253, 16'd49618, 16'd11396, 16'd64201, 16'd20012, 16'd14755, 16'd38032, 16'd7833, 16'd54271, 16'd63983, 16'd62889, 16'd46488, 16'd13451, 16'd14938, 16'd28720, 16'd3708, 16'd13912, 16'd50420, 16'd61828, 16'd60896, 16'd5913, 16'd61101, 16'd32716, 16'd39570, 16'd44691});
	test_expansion(128'h2081134a32ba8f3e1d9da646a9a91dac, {16'd10397, 16'd60746, 16'd44296, 16'd2119, 16'd34365, 16'd20369, 16'd38977, 16'd59948, 16'd21040, 16'd6540, 16'd25256, 16'd55224, 16'd60215, 16'd10228, 16'd2041, 16'd61305, 16'd58997, 16'd60198, 16'd12359, 16'd51871, 16'd608, 16'd11442, 16'd22714, 16'd18886, 16'd42554, 16'd61713});
	test_expansion(128'h4a25cab8042fa839f55ac82a1523462f, {16'd59242, 16'd61208, 16'd11095, 16'd11312, 16'd64835, 16'd48908, 16'd43, 16'd64438, 16'd6241, 16'd62590, 16'd885, 16'd35742, 16'd30138, 16'd49566, 16'd42649, 16'd32935, 16'd21580, 16'd49871, 16'd21491, 16'd63635, 16'd11000, 16'd62851, 16'd9647, 16'd8656, 16'd40536, 16'd23481});
	test_expansion(128'h72fb6f1230f9eda56b4552068d8d341c, {16'd63920, 16'd48773, 16'd20467, 16'd40620, 16'd12384, 16'd30667, 16'd11110, 16'd46676, 16'd19805, 16'd36390, 16'd50048, 16'd44899, 16'd53885, 16'd8219, 16'd43093, 16'd52106, 16'd47434, 16'd11049, 16'd1233, 16'd46680, 16'd48891, 16'd28684, 16'd58989, 16'd40558, 16'd9745, 16'd59299});
	test_expansion(128'h74725daeeafc1095f7143f7da1b81e0c, {16'd16321, 16'd47284, 16'd29043, 16'd2814, 16'd56826, 16'd41720, 16'd6758, 16'd54382, 16'd37436, 16'd7187, 16'd9631, 16'd51229, 16'd10311, 16'd21915, 16'd11439, 16'd51658, 16'd63993, 16'd20563, 16'd29929, 16'd36258, 16'd37115, 16'd60454, 16'd43534, 16'd65142, 16'd62760, 16'd50451});
	test_expansion(128'hf57b4407ce406bf7b37b04e6ae17dec1, {16'd44686, 16'd55236, 16'd32748, 16'd50834, 16'd32922, 16'd31001, 16'd51114, 16'd53386, 16'd29346, 16'd21002, 16'd29384, 16'd24309, 16'd847, 16'd43651, 16'd30487, 16'd55286, 16'd31783, 16'd12832, 16'd54764, 16'd46470, 16'd60813, 16'd40866, 16'd3542, 16'd18777, 16'd16429, 16'd7841});
	test_expansion(128'h7be136138aad5aea1304dc72e7083531, {16'd54956, 16'd13471, 16'd25312, 16'd57771, 16'd18151, 16'd47112, 16'd34609, 16'd55375, 16'd57267, 16'd32106, 16'd61631, 16'd60546, 16'd13542, 16'd31534, 16'd32332, 16'd15340, 16'd44818, 16'd19573, 16'd60298, 16'd3732, 16'd44214, 16'd14451, 16'd25925, 16'd18196, 16'd50326, 16'd30368});
	test_expansion(128'hc40a457040ca3325c36cb6e8057e619c, {16'd41380, 16'd62995, 16'd18935, 16'd3792, 16'd52982, 16'd60665, 16'd54847, 16'd21126, 16'd58908, 16'd17732, 16'd27438, 16'd24534, 16'd58143, 16'd27011, 16'd13489, 16'd39611, 16'd59452, 16'd50125, 16'd58335, 16'd18372, 16'd20593, 16'd50761, 16'd25444, 16'd14111, 16'd55479, 16'd28391});
	test_expansion(128'h2199c35acbd8300be8eaa91011882311, {16'd34112, 16'd14896, 16'd40380, 16'd54423, 16'd38884, 16'd50029, 16'd52175, 16'd45435, 16'd20615, 16'd7407, 16'd50612, 16'd4193, 16'd32732, 16'd48625, 16'd607, 16'd20528, 16'd56601, 16'd1332, 16'd24880, 16'd394, 16'd17965, 16'd8439, 16'd46937, 16'd41562, 16'd35803, 16'd7907});
	test_expansion(128'h0c1388abda66f5b333a10cc4d40fac72, {16'd22377, 16'd22920, 16'd30560, 16'd48312, 16'd31237, 16'd27628, 16'd63565, 16'd47542, 16'd65283, 16'd23815, 16'd55446, 16'd2853, 16'd35004, 16'd45881, 16'd58576, 16'd15386, 16'd43127, 16'd30343, 16'd63084, 16'd13652, 16'd41407, 16'd53132, 16'd27594, 16'd39142, 16'd2980, 16'd3932});
	test_expansion(128'h0a5c015699191365cc847e0e42e49591, {16'd52337, 16'd4043, 16'd6677, 16'd21821, 16'd29889, 16'd42270, 16'd43855, 16'd48167, 16'd2252, 16'd60414, 16'd53251, 16'd28450, 16'd58535, 16'd17450, 16'd58729, 16'd60073, 16'd39576, 16'd34262, 16'd59966, 16'd49379, 16'd21720, 16'd53317, 16'd55004, 16'd34591, 16'd60193, 16'd49139});
	test_expansion(128'hdfbfe6020d09d8d9b79fc10573eff636, {16'd34896, 16'd61344, 16'd28492, 16'd14713, 16'd51214, 16'd20375, 16'd34279, 16'd4750, 16'd9629, 16'd8399, 16'd33035, 16'd13659, 16'd7452, 16'd50832, 16'd26913, 16'd60494, 16'd29624, 16'd35905, 16'd41032, 16'd49185, 16'd6370, 16'd48929, 16'd32230, 16'd3158, 16'd58496, 16'd58600});
	test_expansion(128'hc4216d6877e8b315ed85421ef5dcf2ce, {16'd2507, 16'd41761, 16'd58384, 16'd29732, 16'd43060, 16'd4576, 16'd8673, 16'd3202, 16'd61695, 16'd6231, 16'd22523, 16'd580, 16'd42416, 16'd38562, 16'd42554, 16'd42379, 16'd51439, 16'd21372, 16'd65446, 16'd2773, 16'd30886, 16'd64918, 16'd5877, 16'd2080, 16'd59267, 16'd31224});
	test_expansion(128'hba86c515a968b31ddf94fb718b9161b4, {16'd61969, 16'd28312, 16'd16142, 16'd45901, 16'd59121, 16'd61910, 16'd7700, 16'd46252, 16'd6044, 16'd7206, 16'd41027, 16'd17399, 16'd29627, 16'd54297, 16'd48467, 16'd24207, 16'd14030, 16'd29435, 16'd12877, 16'd25546, 16'd26692, 16'd57847, 16'd12082, 16'd8053, 16'd52060, 16'd31043});
	test_expansion(128'h797a5bb340b37d6da13c62b27737efc9, {16'd36122, 16'd43651, 16'd43721, 16'd49267, 16'd61288, 16'd29501, 16'd36642, 16'd3020, 16'd14210, 16'd58261, 16'd38679, 16'd50244, 16'd6274, 16'd62055, 16'd41682, 16'd26731, 16'd26682, 16'd59832, 16'd14717, 16'd2479, 16'd4624, 16'd51071, 16'd34637, 16'd24043, 16'd54662, 16'd52004});
	test_expansion(128'h6449cd27462253f70e75f9229be02efe, {16'd49082, 16'd17448, 16'd10860, 16'd28291, 16'd50284, 16'd13565, 16'd3265, 16'd42302, 16'd42146, 16'd59276, 16'd15235, 16'd47735, 16'd30870, 16'd58897, 16'd65454, 16'd6526, 16'd32149, 16'd1694, 16'd51077, 16'd30600, 16'd59462, 16'd65228, 16'd55712, 16'd32572, 16'd46639, 16'd45317});
	test_expansion(128'h28a4d8437ba04212b26ce895d277942b, {16'd62095, 16'd31461, 16'd15613, 16'd44851, 16'd11898, 16'd17475, 16'd48532, 16'd2293, 16'd16096, 16'd37879, 16'd38614, 16'd61449, 16'd34008, 16'd59293, 16'd44280, 16'd39782, 16'd24557, 16'd45370, 16'd55794, 16'd51698, 16'd37843, 16'd51360, 16'd16588, 16'd58694, 16'd9463, 16'd7610});
	test_expansion(128'h3d887c68aaa7d2702c3452813bb55b36, {16'd32428, 16'd36234, 16'd52171, 16'd40182, 16'd8960, 16'd37344, 16'd32684, 16'd38224, 16'd33356, 16'd63380, 16'd8015, 16'd4883, 16'd5991, 16'd54011, 16'd7536, 16'd5741, 16'd1775, 16'd21970, 16'd42845, 16'd902, 16'd2079, 16'd64468, 16'd8140, 16'd41434, 16'd39537, 16'd53826});
	test_expansion(128'hf2e48256cd12cd63e35d2df71494fb27, {16'd45887, 16'd57140, 16'd50969, 16'd62194, 16'd1534, 16'd23773, 16'd20857, 16'd32422, 16'd49733, 16'd10243, 16'd30985, 16'd13382, 16'd28240, 16'd61070, 16'd34371, 16'd30462, 16'd21575, 16'd6095, 16'd7248, 16'd9479, 16'd62761, 16'd30643, 16'd54285, 16'd22189, 16'd57487, 16'd15112});
	test_expansion(128'hf75ccfe726fa506da0d5f0a29430969d, {16'd1463, 16'd18642, 16'd63425, 16'd33323, 16'd54273, 16'd29195, 16'd12775, 16'd37230, 16'd39633, 16'd15341, 16'd12006, 16'd46815, 16'd32553, 16'd22722, 16'd64243, 16'd12138, 16'd5358, 16'd13421, 16'd20257, 16'd31712, 16'd31515, 16'd62625, 16'd40950, 16'd13408, 16'd30049, 16'd31576});
	test_expansion(128'h944b611842764b1f9aab24f56506d841, {16'd46564, 16'd57113, 16'd4438, 16'd15605, 16'd63904, 16'd31878, 16'd28184, 16'd25831, 16'd29980, 16'd8898, 16'd19697, 16'd19896, 16'd13374, 16'd37595, 16'd21057, 16'd7406, 16'd56805, 16'd65260, 16'd60047, 16'd17589, 16'd6587, 16'd64738, 16'd16590, 16'd17880, 16'd62845, 16'd40614});
	test_expansion(128'h80b73b60dc62f218917dc19d60d10830, {16'd51911, 16'd28148, 16'd25427, 16'd51909, 16'd42416, 16'd31669, 16'd12643, 16'd4611, 16'd52237, 16'd21055, 16'd43744, 16'd15082, 16'd63470, 16'd12104, 16'd61843, 16'd5982, 16'd13720, 16'd57768, 16'd62114, 16'd441, 16'd7597, 16'd15316, 16'd18846, 16'd38771, 16'd63911, 16'd36823});
	test_expansion(128'h07221b09ac1c8e577f96bd4522b4d05d, {16'd1960, 16'd56548, 16'd4830, 16'd39884, 16'd41740, 16'd5493, 16'd51494, 16'd908, 16'd9303, 16'd43547, 16'd57863, 16'd35599, 16'd17863, 16'd15238, 16'd21470, 16'd53278, 16'd17597, 16'd61873, 16'd16786, 16'd7000, 16'd50251, 16'd15189, 16'd46677, 16'd1983, 16'd61818, 16'd30697});
	test_expansion(128'h7ca3960cb5edc4323cca2cbb0c0f2eb8, {16'd37115, 16'd41093, 16'd12538, 16'd22465, 16'd27692, 16'd9105, 16'd49868, 16'd28916, 16'd58563, 16'd24176, 16'd30613, 16'd27840, 16'd54843, 16'd33, 16'd10754, 16'd26722, 16'd56512, 16'd29538, 16'd33903, 16'd3202, 16'd14576, 16'd30571, 16'd51451, 16'd52275, 16'd36484, 16'd5160});
	test_expansion(128'h745dc33a9fd0f3fae2f9f611f2b2592c, {16'd31567, 16'd4728, 16'd39021, 16'd13412, 16'd29626, 16'd21927, 16'd55069, 16'd31346, 16'd50340, 16'd22100, 16'd27816, 16'd59178, 16'd47881, 16'd1919, 16'd11382, 16'd55575, 16'd56286, 16'd8603, 16'd9524, 16'd21336, 16'd7992, 16'd7859, 16'd17414, 16'd62904, 16'd11970, 16'd18323});
	test_expansion(128'h34cc87d6a1035ec198b8d27dde432086, {16'd47716, 16'd61476, 16'd12526, 16'd3006, 16'd65370, 16'd41720, 16'd44356, 16'd26313, 16'd36481, 16'd12066, 16'd22908, 16'd29236, 16'd46605, 16'd40282, 16'd13006, 16'd3602, 16'd1787, 16'd55190, 16'd58928, 16'd46646, 16'd12245, 16'd196, 16'd52149, 16'd25449, 16'd39634, 16'd27652});
	test_expansion(128'h9a56ce7abe7908d4ead1abf33aed3dcd, {16'd15973, 16'd59140, 16'd49323, 16'd1741, 16'd22248, 16'd29463, 16'd52814, 16'd16885, 16'd47054, 16'd20810, 16'd11396, 16'd34292, 16'd53678, 16'd35435, 16'd61021, 16'd33744, 16'd10426, 16'd4449, 16'd20793, 16'd21065, 16'd5474, 16'd6064, 16'd52305, 16'd17427, 16'd52875, 16'd52859});
	test_expansion(128'ha789b3b7f7ff58f49e187fe375e0029b, {16'd26544, 16'd52157, 16'd38107, 16'd39984, 16'd55013, 16'd47318, 16'd53748, 16'd62949, 16'd3415, 16'd51085, 16'd35052, 16'd58841, 16'd33625, 16'd4112, 16'd39045, 16'd23359, 16'd61261, 16'd3589, 16'd32472, 16'd4388, 16'd32642, 16'd2602, 16'd53125, 16'd19214, 16'd438, 16'd30639});
	test_expansion(128'hb6168d2b5c1543c4f8c971326f800793, {16'd3632, 16'd38346, 16'd18787, 16'd25914, 16'd43711, 16'd15638, 16'd10250, 16'd49836, 16'd16935, 16'd22360, 16'd6299, 16'd36461, 16'd18620, 16'd5233, 16'd9464, 16'd2729, 16'd6208, 16'd26528, 16'd20545, 16'd36231, 16'd31773, 16'd12753, 16'd29716, 16'd50762, 16'd20185, 16'd59036});
	test_expansion(128'hc454a0bb04ddf2700b4f2d73b318d92e, {16'd43676, 16'd63407, 16'd50065, 16'd43013, 16'd16915, 16'd53359, 16'd15697, 16'd362, 16'd44397, 16'd46569, 16'd38973, 16'd19663, 16'd23747, 16'd37318, 16'd8009, 16'd12208, 16'd20136, 16'd12000, 16'd60896, 16'd26175, 16'd64126, 16'd6688, 16'd4003, 16'd12465, 16'd43670, 16'd51110});
	test_expansion(128'h9169d7cd38ff2aeb3affb5eb73d66cec, {16'd2162, 16'd57011, 16'd28052, 16'd989, 16'd63295, 16'd58464, 16'd39018, 16'd44099, 16'd31835, 16'd55624, 16'd12118, 16'd62277, 16'd6736, 16'd57814, 16'd22003, 16'd58435, 16'd47773, 16'd52229, 16'd44879, 16'd61274, 16'd21312, 16'd51176, 16'd30731, 16'd17603, 16'd648, 16'd5519});
	test_expansion(128'h7dab6accba8869433639cf42b740a840, {16'd31165, 16'd57445, 16'd24787, 16'd11546, 16'd27203, 16'd11548, 16'd41781, 16'd26753, 16'd62373, 16'd38008, 16'd16411, 16'd59755, 16'd35703, 16'd48578, 16'd12664, 16'd50432, 16'd35171, 16'd44513, 16'd36931, 16'd16263, 16'd34432, 16'd25440, 16'd10558, 16'd43158, 16'd56283, 16'd648});
	test_expansion(128'hd4fad18211589033b5d467058a56c8a1, {16'd41949, 16'd55669, 16'd63849, 16'd14241, 16'd2954, 16'd56641, 16'd61381, 16'd22605, 16'd38112, 16'd25420, 16'd58757, 16'd54801, 16'd49556, 16'd37089, 16'd12808, 16'd45436, 16'd60174, 16'd61323, 16'd19986, 16'd29458, 16'd38909, 16'd43243, 16'd57658, 16'd35113, 16'd58009, 16'd16487});
	test_expansion(128'h82a059f692c06dfba7e478e834c221b5, {16'd15270, 16'd50905, 16'd38742, 16'd23158, 16'd40207, 16'd19834, 16'd71, 16'd7590, 16'd17525, 16'd46692, 16'd31812, 16'd19675, 16'd26362, 16'd14555, 16'd32694, 16'd43778, 16'd44280, 16'd28730, 16'd45658, 16'd45961, 16'd883, 16'd48444, 16'd34484, 16'd45780, 16'd25679, 16'd25721});
	test_expansion(128'h0f79fe4fb1a3c9b40ecd2d86236c9bf7, {16'd52283, 16'd15377, 16'd32019, 16'd26178, 16'd38274, 16'd58230, 16'd22748, 16'd53244, 16'd45015, 16'd48156, 16'd19984, 16'd61675, 16'd53522, 16'd16930, 16'd27808, 16'd31064, 16'd2431, 16'd34840, 16'd35132, 16'd20053, 16'd3425, 16'd36440, 16'd49892, 16'd28945, 16'd33457, 16'd45075});
	test_expansion(128'hfcc3fc89a826d6530f43ab15d4ab55a0, {16'd43792, 16'd15686, 16'd30792, 16'd33748, 16'd55612, 16'd5075, 16'd60111, 16'd3942, 16'd15756, 16'd28975, 16'd590, 16'd49406, 16'd10128, 16'd28367, 16'd6735, 16'd10636, 16'd52310, 16'd10006, 16'd3149, 16'd3403, 16'd63432, 16'd5482, 16'd44604, 16'd11586, 16'd13962, 16'd599});
	test_expansion(128'h84fb78fec15b8dac21a15dd6a8f4e27c, {16'd34478, 16'd58265, 16'd62176, 16'd1992, 16'd50770, 16'd56872, 16'd39750, 16'd37485, 16'd27026, 16'd36019, 16'd27124, 16'd31637, 16'd31643, 16'd50577, 16'd4381, 16'd7413, 16'd24721, 16'd37280, 16'd40917, 16'd12879, 16'd49670, 16'd18492, 16'd45898, 16'd64119, 16'd28326, 16'd53293});
	test_expansion(128'hf9f600feb08330d9fccef8694149c68f, {16'd19762, 16'd55387, 16'd26815, 16'd50124, 16'd1619, 16'd12027, 16'd28005, 16'd21875, 16'd13760, 16'd50662, 16'd28675, 16'd37189, 16'd35864, 16'd7419, 16'd36578, 16'd49876, 16'd54081, 16'd34388, 16'd11964, 16'd40397, 16'd33978, 16'd39700, 16'd24854, 16'd56801, 16'd45300, 16'd39231});
	test_expansion(128'h1e33f79c56af7a84e403836651362780, {16'd3004, 16'd62969, 16'd50431, 16'd36644, 16'd34897, 16'd57241, 16'd13476, 16'd45587, 16'd27701, 16'd29031, 16'd22281, 16'd36908, 16'd20670, 16'd4746, 16'd23876, 16'd18989, 16'd62758, 16'd27753, 16'd46877, 16'd31552, 16'd39306, 16'd55218, 16'd26500, 16'd56652, 16'd45539, 16'd29096});
	test_expansion(128'h579550631fb76cb7c8f39b21e32c2145, {16'd27009, 16'd60420, 16'd50236, 16'd42648, 16'd4200, 16'd55713, 16'd37489, 16'd16904, 16'd8922, 16'd27696, 16'd58014, 16'd43617, 16'd20727, 16'd47625, 16'd44814, 16'd713, 16'd20200, 16'd61379, 16'd43288, 16'd4178, 16'd34792, 16'd55831, 16'd24093, 16'd61734, 16'd3520, 16'd25227});
	test_expansion(128'h87ed8fcdca9f8d0a77026b5d0928823f, {16'd28325, 16'd60779, 16'd30658, 16'd18545, 16'd1378, 16'd35963, 16'd7711, 16'd13483, 16'd61168, 16'd27213, 16'd55692, 16'd33277, 16'd255, 16'd16903, 16'd52166, 16'd37371, 16'd1796, 16'd38417, 16'd36191, 16'd34570, 16'd63664, 16'd28759, 16'd59764, 16'd17197, 16'd62846, 16'd49214});
	test_expansion(128'h24a32ba94959b0bcb15eb0be6dfbb805, {16'd46352, 16'd667, 16'd10163, 16'd8986, 16'd954, 16'd18, 16'd42202, 16'd20460, 16'd35217, 16'd26053, 16'd59763, 16'd26931, 16'd20857, 16'd25230, 16'd6975, 16'd35641, 16'd41940, 16'd50184, 16'd29241, 16'd1999, 16'd10993, 16'd39601, 16'd25531, 16'd28374, 16'd43231, 16'd24021});
	test_expansion(128'h571a84cd4d1c17def2a285a381a13d16, {16'd31467, 16'd57768, 16'd47599, 16'd22519, 16'd35908, 16'd41765, 16'd40045, 16'd10547, 16'd13228, 16'd24328, 16'd47596, 16'd36358, 16'd25779, 16'd60224, 16'd61226, 16'd40245, 16'd35318, 16'd96, 16'd17890, 16'd47623, 16'd9722, 16'd31616, 16'd54323, 16'd248, 16'd24215, 16'd65186});
	test_expansion(128'hb0c22d0fe8f0ddb8ec191ae5858dc518, {16'd44565, 16'd37702, 16'd8427, 16'd32970, 16'd27472, 16'd1060, 16'd18196, 16'd48109, 16'd44327, 16'd34046, 16'd39232, 16'd57210, 16'd57587, 16'd59868, 16'd3831, 16'd26253, 16'd58524, 16'd12504, 16'd34107, 16'd17188, 16'd16218, 16'd5617, 16'd23412, 16'd28645, 16'd39721, 16'd28237});
	test_expansion(128'h6d03ff360f14599cef1af89341157536, {16'd43590, 16'd60542, 16'd28817, 16'd39178, 16'd28515, 16'd33560, 16'd59595, 16'd63881, 16'd9131, 16'd2172, 16'd5326, 16'd45574, 16'd40542, 16'd27098, 16'd35170, 16'd55064, 16'd55425, 16'd8315, 16'd45833, 16'd63455, 16'd7028, 16'd20492, 16'd64243, 16'd62780, 16'd24249, 16'd21407});
	test_expansion(128'hdca1afdf1dce5ff48317ff6f7c19d7ca, {16'd60766, 16'd8980, 16'd7435, 16'd43246, 16'd48012, 16'd25048, 16'd36932, 16'd10677, 16'd14377, 16'd17009, 16'd8581, 16'd41037, 16'd48398, 16'd44727, 16'd9154, 16'd12252, 16'd21011, 16'd44532, 16'd34663, 16'd13426, 16'd803, 16'd32233, 16'd22871, 16'd14376, 16'd7889, 16'd50621});
	test_expansion(128'h4c3bce9f2eb755c71c3417cd62d8d4fa, {16'd2814, 16'd40846, 16'd29961, 16'd48230, 16'd19322, 16'd38348, 16'd45463, 16'd54866, 16'd53144, 16'd51618, 16'd18875, 16'd34274, 16'd10023, 16'd64477, 16'd41143, 16'd28777, 16'd17687, 16'd59964, 16'd4814, 16'd22678, 16'd7856, 16'd60462, 16'd24784, 16'd22363, 16'd18092, 16'd2132});
	test_expansion(128'hdf92a17fc9e754678b5f5319bc9e5f80, {16'd15486, 16'd27871, 16'd32368, 16'd42875, 16'd26076, 16'd36098, 16'd57499, 16'd19449, 16'd21431, 16'd41107, 16'd58862, 16'd26029, 16'd44068, 16'd41173, 16'd38093, 16'd51297, 16'd11769, 16'd49315, 16'd42099, 16'd56540, 16'd50413, 16'd3405, 16'd2670, 16'd44310, 16'd62280, 16'd43610});
	test_expansion(128'h8a52ad073468d1b7fb8f61058908b2e4, {16'd34167, 16'd44634, 16'd9547, 16'd39415, 16'd3162, 16'd45936, 16'd30595, 16'd24509, 16'd20164, 16'd58610, 16'd55645, 16'd48449, 16'd63432, 16'd61786, 16'd29179, 16'd17114, 16'd35708, 16'd44208, 16'd24538, 16'd42246, 16'd29091, 16'd14939, 16'd20580, 16'd2326, 16'd53530, 16'd4227});
	test_expansion(128'h1f31a8f2afdac584860c986c5d45a662, {16'd48715, 16'd25305, 16'd43904, 16'd4331, 16'd18577, 16'd17778, 16'd32428, 16'd58027, 16'd41186, 16'd40945, 16'd17860, 16'd60607, 16'd41314, 16'd3337, 16'd51678, 16'd37075, 16'd7287, 16'd36266, 16'd32172, 16'd3873, 16'd32364, 16'd64795, 16'd35189, 16'd47707, 16'd19413, 16'd44237});
	test_expansion(128'hfcc25a9411653800d9537a95ed266a34, {16'd30748, 16'd47842, 16'd8324, 16'd39399, 16'd57199, 16'd41277, 16'd9128, 16'd19913, 16'd21640, 16'd59628, 16'd16949, 16'd9513, 16'd49350, 16'd36711, 16'd18793, 16'd36447, 16'd50265, 16'd53597, 16'd65226, 16'd56008, 16'd15891, 16'd39318, 16'd61308, 16'd26032, 16'd53109, 16'd56703});
	test_expansion(128'h9023180fb7d646388135622c79d709c1, {16'd18066, 16'd24276, 16'd18232, 16'd38563, 16'd57604, 16'd21746, 16'd38442, 16'd25930, 16'd8785, 16'd12308, 16'd23606, 16'd12124, 16'd16727, 16'd32289, 16'd62962, 16'd32043, 16'd16199, 16'd49064, 16'd22454, 16'd56435, 16'd15130, 16'd2231, 16'd6335, 16'd4778, 16'd51580, 16'd18981});
	test_expansion(128'h67e81622b469e5cc8fcafb2f41196938, {16'd26506, 16'd26829, 16'd33260, 16'd31043, 16'd50703, 16'd33033, 16'd42065, 16'd55446, 16'd63560, 16'd31261, 16'd9176, 16'd27592, 16'd22956, 16'd30011, 16'd27960, 16'd16778, 16'd11071, 16'd10181, 16'd44029, 16'd25198, 16'd2890, 16'd37442, 16'd43561, 16'd19169, 16'd45401, 16'd17786});
	test_expansion(128'h75a68ccccba12d3ac9664837631d2616, {16'd13983, 16'd41283, 16'd59306, 16'd63345, 16'd25836, 16'd719, 16'd61209, 16'd19812, 16'd27076, 16'd61641, 16'd60333, 16'd21035, 16'd54770, 16'd47293, 16'd7912, 16'd53187, 16'd25398, 16'd57869, 16'd25518, 16'd24946, 16'd48823, 16'd64812, 16'd20358, 16'd575, 16'd51525, 16'd56539});
	test_expansion(128'hc2888ff40f0b7f048e3ee07006c21dc3, {16'd15751, 16'd384, 16'd58755, 16'd26552, 16'd21944, 16'd20929, 16'd3027, 16'd61262, 16'd5558, 16'd46777, 16'd25548, 16'd58420, 16'd2023, 16'd58973, 16'd22026, 16'd58898, 16'd56462, 16'd15096, 16'd31451, 16'd13205, 16'd38947, 16'd61157, 16'd64789, 16'd56747, 16'd52480, 16'd22075});
	test_expansion(128'h8da02ae82ebd53bc233fef0cf5dc62b9, {16'd14704, 16'd4784, 16'd25583, 16'd28489, 16'd9635, 16'd3001, 16'd48018, 16'd39835, 16'd63014, 16'd9894, 16'd58828, 16'd25952, 16'd59366, 16'd35055, 16'd22796, 16'd47177, 16'd27432, 16'd12306, 16'd43622, 16'd39005, 16'd33828, 16'd33877, 16'd32221, 16'd65494, 16'd16426, 16'd45817});
	test_expansion(128'hc1634e1d8ad5e37cfffc2c7bb0ba527b, {16'd23021, 16'd40363, 16'd28256, 16'd24262, 16'd13071, 16'd26498, 16'd42874, 16'd29176, 16'd47895, 16'd21356, 16'd15405, 16'd13789, 16'd58322, 16'd37505, 16'd10443, 16'd51110, 16'd886, 16'd55124, 16'd25854, 16'd63658, 16'd30963, 16'd27512, 16'd30642, 16'd37947, 16'd25098, 16'd12324});
	test_expansion(128'hb2253a7a6b3237f8a00cd83fb903f5c2, {16'd2249, 16'd24613, 16'd64110, 16'd61762, 16'd1354, 16'd47962, 16'd9048, 16'd2354, 16'd30026, 16'd8652, 16'd18015, 16'd18745, 16'd21577, 16'd13183, 16'd29586, 16'd29760, 16'd24447, 16'd7232, 16'd36506, 16'd54651, 16'd25972, 16'd30416, 16'd29173, 16'd26965, 16'd45831, 16'd47387});
	test_expansion(128'h2b932c0f8c1a1945eb89060ad71c3c3f, {16'd27915, 16'd4155, 16'd10517, 16'd52350, 16'd23901, 16'd60164, 16'd29248, 16'd46388, 16'd64494, 16'd57371, 16'd32287, 16'd47395, 16'd49115, 16'd43087, 16'd25357, 16'd29501, 16'd10621, 16'd42253, 16'd17961, 16'd55713, 16'd32323, 16'd2059, 16'd15403, 16'd4471, 16'd38454, 16'd49626});
	test_expansion(128'hbb10d27bcc9b0a29f11ee3570d1bf51f, {16'd21769, 16'd57863, 16'd48603, 16'd27999, 16'd55180, 16'd29603, 16'd5608, 16'd10295, 16'd55487, 16'd64153, 16'd60688, 16'd25888, 16'd39412, 16'd56997, 16'd48169, 16'd61086, 16'd32495, 16'd63772, 16'd9534, 16'd26818, 16'd50196, 16'd13954, 16'd717, 16'd34516, 16'd41214, 16'd42274});
	test_expansion(128'h2267de54c88fb6e956364b9347454622, {16'd6769, 16'd58628, 16'd63936, 16'd26753, 16'd56193, 16'd36752, 16'd13205, 16'd52634, 16'd36983, 16'd13220, 16'd35308, 16'd45981, 16'd24476, 16'd27894, 16'd29605, 16'd54401, 16'd441, 16'd44916, 16'd12381, 16'd60081, 16'd33005, 16'd44767, 16'd19910, 16'd21836, 16'd31302, 16'd34174});
	test_expansion(128'h715d236d98514e5f99a09a7aabe9cc51, {16'd34478, 16'd6228, 16'd51836, 16'd55411, 16'd56750, 16'd9585, 16'd30635, 16'd49650, 16'd32584, 16'd10274, 16'd26986, 16'd36164, 16'd728, 16'd27958, 16'd39469, 16'd33343, 16'd25443, 16'd16644, 16'd62141, 16'd54781, 16'd9376, 16'd39019, 16'd65198, 16'd4581, 16'd41124, 16'd15786});
	test_expansion(128'h6b73d2f220e7c52aca88d2ea004e5018, {16'd35735, 16'd18588, 16'd15838, 16'd46139, 16'd36890, 16'd29872, 16'd51627, 16'd17277, 16'd7816, 16'd51731, 16'd19658, 16'd36631, 16'd12157, 16'd17311, 16'd31310, 16'd50776, 16'd16295, 16'd39267, 16'd26478, 16'd16960, 16'd9137, 16'd59193, 16'd50445, 16'd61499, 16'd62344, 16'd27316});
	test_expansion(128'h2fb196a7d756ad6c66baa771c0ed250a, {16'd3461, 16'd26942, 16'd53596, 16'd39, 16'd41379, 16'd64391, 16'd10684, 16'd2089, 16'd51557, 16'd31049, 16'd15271, 16'd14269, 16'd58287, 16'd40273, 16'd31654, 16'd51704, 16'd65211, 16'd46520, 16'd33686, 16'd49644, 16'd54997, 16'd34645, 16'd17760, 16'd19821, 16'd49265, 16'd2686});
	test_expansion(128'hde79c9eb80ab787c4b3a3a6aa0d117d1, {16'd47213, 16'd56604, 16'd58572, 16'd31178, 16'd35381, 16'd58265, 16'd30223, 16'd6296, 16'd18984, 16'd47544, 16'd18871, 16'd29251, 16'd40347, 16'd48243, 16'd21480, 16'd13075, 16'd47849, 16'd36741, 16'd52946, 16'd61943, 16'd42667, 16'd36876, 16'd7858, 16'd14110, 16'd50294, 16'd65092});
	test_expansion(128'hecbe95f15ecea4bf271a24e9b4d66693, {16'd396, 16'd24632, 16'd16493, 16'd2603, 16'd38697, 16'd50034, 16'd17974, 16'd5439, 16'd4705, 16'd17259, 16'd5613, 16'd38895, 16'd27408, 16'd41468, 16'd27956, 16'd28169, 16'd63788, 16'd61554, 16'd19412, 16'd36572, 16'd15445, 16'd13643, 16'd30187, 16'd44764, 16'd34782, 16'd11880});
	test_expansion(128'hd030f50a8d56b6284448aab22ac33c72, {16'd34074, 16'd52239, 16'd5852, 16'd1190, 16'd16050, 16'd15512, 16'd15206, 16'd48725, 16'd53756, 16'd64240, 16'd7399, 16'd22106, 16'd43463, 16'd62135, 16'd54334, 16'd45746, 16'd55096, 16'd14061, 16'd34263, 16'd30419, 16'd26040, 16'd34540, 16'd5418, 16'd29050, 16'd36770, 16'd14518});
	test_expansion(128'h8dd6863d18ef1dbe2c6cd661564a2cdf, {16'd581, 16'd64998, 16'd34711, 16'd43535, 16'd34761, 16'd22898, 16'd64731, 16'd20394, 16'd4018, 16'd62735, 16'd4309, 16'd8254, 16'd27095, 16'd9385, 16'd60934, 16'd27399, 16'd1781, 16'd30534, 16'd397, 16'd48607, 16'd54327, 16'd48914, 16'd30278, 16'd61357, 16'd11649, 16'd30946});
	test_expansion(128'h53be0e92652b4f13eff954efa2faa310, {16'd46757, 16'd2677, 16'd46127, 16'd20229, 16'd40900, 16'd11440, 16'd23116, 16'd21500, 16'd14307, 16'd25223, 16'd23129, 16'd201, 16'd8664, 16'd46038, 16'd37341, 16'd8306, 16'd6748, 16'd4325, 16'd5027, 16'd36320, 16'd51389, 16'd13770, 16'd37901, 16'd27477, 16'd9546, 16'd48741});
	test_expansion(128'hcf544944bc4fc2a12961bf2bcc445521, {16'd23273, 16'd24372, 16'd55698, 16'd23668, 16'd26372, 16'd18982, 16'd14044, 16'd61553, 16'd41625, 16'd18965, 16'd33763, 16'd3520, 16'd63718, 16'd17377, 16'd14420, 16'd63589, 16'd10184, 16'd60014, 16'd22106, 16'd9485, 16'd12730, 16'd62944, 16'd38052, 16'd36452, 16'd16738, 16'd9136});
	test_expansion(128'h7b92199b6c09dd64a865d0d6710cb75a, {16'd60424, 16'd8190, 16'd2361, 16'd60655, 16'd40735, 16'd46886, 16'd5076, 16'd57676, 16'd31659, 16'd7176, 16'd11034, 16'd54546, 16'd31519, 16'd33985, 16'd27894, 16'd8662, 16'd16265, 16'd1003, 16'd32040, 16'd20791, 16'd65449, 16'd38779, 16'd59463, 16'd45680, 16'd3143, 16'd57485});
	test_expansion(128'ha1f33c0afb2da1ec3e1333f5f9310aae, {16'd38570, 16'd58381, 16'd29433, 16'd6112, 16'd36509, 16'd26787, 16'd28012, 16'd349, 16'd62892, 16'd5055, 16'd23168, 16'd22156, 16'd18932, 16'd13986, 16'd43879, 16'd9185, 16'd47588, 16'd16918, 16'd2495, 16'd40758, 16'd35152, 16'd21152, 16'd42358, 16'd54885, 16'd54848, 16'd58619});
	test_expansion(128'hf12f92fc5ac155b215af2073231fefad, {16'd22562, 16'd65080, 16'd64396, 16'd32642, 16'd61336, 16'd29588, 16'd38128, 16'd12588, 16'd37699, 16'd1687, 16'd43824, 16'd7697, 16'd38486, 16'd47978, 16'd485, 16'd65005, 16'd48945, 16'd20732, 16'd60658, 16'd29586, 16'd20383, 16'd48463, 16'd60635, 16'd50066, 16'd53338, 16'd55314});
	test_expansion(128'h31d3b9b362e676252ba72e4eb29ef81a, {16'd33598, 16'd16077, 16'd31855, 16'd64787, 16'd54812, 16'd35555, 16'd18698, 16'd29627, 16'd9089, 16'd54314, 16'd6385, 16'd17963, 16'd9256, 16'd19168, 16'd11829, 16'd27776, 16'd54693, 16'd37625, 16'd14001, 16'd58805, 16'd3121, 16'd5087, 16'd45768, 16'd25913, 16'd39947, 16'd52764});
	test_expansion(128'ha648bcc46dce0d81e45556beec016fcb, {16'd37811, 16'd12644, 16'd56615, 16'd23979, 16'd23701, 16'd44614, 16'd30289, 16'd20124, 16'd63806, 16'd53837, 16'd14974, 16'd36873, 16'd27692, 16'd55326, 16'd15235, 16'd21395, 16'd36924, 16'd55186, 16'd6697, 16'd44428, 16'd429, 16'd11463, 16'd304, 16'd40160, 16'd49991, 16'd46824});
	test_expansion(128'h230ca86b074c7d99d54080aee73d7263, {16'd58712, 16'd30244, 16'd39102, 16'd49753, 16'd4142, 16'd30646, 16'd52365, 16'd4247, 16'd26272, 16'd48376, 16'd59005, 16'd29235, 16'd50381, 16'd63656, 16'd9367, 16'd18961, 16'd12565, 16'd63958, 16'd15530, 16'd58184, 16'd42288, 16'd9069, 16'd39094, 16'd1095, 16'd25263, 16'd12872});
	test_expansion(128'h681e941cb5c344b1d2424bf744d31d8a, {16'd14651, 16'd42812, 16'd42753, 16'd48059, 16'd39479, 16'd62239, 16'd8224, 16'd32006, 16'd29343, 16'd1229, 16'd62454, 16'd60061, 16'd5485, 16'd59219, 16'd18876, 16'd50293, 16'd23956, 16'd63554, 16'd11216, 16'd50037, 16'd35433, 16'd57092, 16'd41401, 16'd9816, 16'd55054, 16'd10528});
	test_expansion(128'h42c19e32d27322a03860cf94d499bf7c, {16'd11551, 16'd52172, 16'd65045, 16'd57934, 16'd62635, 16'd49892, 16'd2040, 16'd53340, 16'd37964, 16'd27617, 16'd46603, 16'd56244, 16'd39447, 16'd51955, 16'd42445, 16'd62191, 16'd43210, 16'd23487, 16'd20482, 16'd58035, 16'd31561, 16'd28295, 16'd63899, 16'd39462, 16'd7149, 16'd18081});
	test_expansion(128'h12edfa21d6ea9528665dfc84d3409cac, {16'd47432, 16'd62319, 16'd56832, 16'd25374, 16'd23537, 16'd12871, 16'd56290, 16'd31137, 16'd42693, 16'd10650, 16'd21313, 16'd18485, 16'd55377, 16'd32715, 16'd25180, 16'd42931, 16'd35268, 16'd15749, 16'd38915, 16'd48189, 16'd19604, 16'd31668, 16'd64112, 16'd13264, 16'd26346, 16'd57749});
	test_expansion(128'h584596d8bca09cb96b14e2ea12948631, {16'd5402, 16'd5318, 16'd55008, 16'd22153, 16'd51928, 16'd45698, 16'd63258, 16'd47581, 16'd2972, 16'd60099, 16'd43720, 16'd29638, 16'd32954, 16'd41580, 16'd39922, 16'd62169, 16'd15168, 16'd61508, 16'd8943, 16'd35040, 16'd53516, 16'd23354, 16'd37358, 16'd26764, 16'd43244, 16'd56295});
	test_expansion(128'h6635bab9a4ffa0fba4df9e29798126e9, {16'd37655, 16'd41490, 16'd64918, 16'd49565, 16'd15178, 16'd5181, 16'd14177, 16'd54925, 16'd35450, 16'd47263, 16'd61949, 16'd27533, 16'd12180, 16'd61958, 16'd61923, 16'd34539, 16'd49402, 16'd49167, 16'd1893, 16'd36102, 16'd49583, 16'd27829, 16'd38614, 16'd54151, 16'd30399, 16'd64636});
	test_expansion(128'hc12e2f046757a4040c9db59739649795, {16'd29385, 16'd29539, 16'd12998, 16'd28961, 16'd57993, 16'd18991, 16'd7656, 16'd48475, 16'd36971, 16'd13730, 16'd17502, 16'd35806, 16'd44446, 16'd28657, 16'd15944, 16'd62286, 16'd51955, 16'd26930, 16'd64501, 16'd7075, 16'd25763, 16'd59330, 16'd61513, 16'd15357, 16'd47824, 16'd52323});
	test_expansion(128'h3446efcc507aa3a5ed9bbe66cbe1bbdf, {16'd5214, 16'd56969, 16'd4460, 16'd30790, 16'd54147, 16'd19954, 16'd46771, 16'd53631, 16'd52407, 16'd45837, 16'd33727, 16'd5069, 16'd5209, 16'd29926, 16'd50731, 16'd1836, 16'd64989, 16'd40311, 16'd17219, 16'd12229, 16'd50311, 16'd41881, 16'd13705, 16'd9178, 16'd371, 16'd3161});
	test_expansion(128'h48f7b569bc9575c7e6d322ad7c09023a, {16'd26065, 16'd61325, 16'd18157, 16'd49653, 16'd2645, 16'd57013, 16'd45280, 16'd60581, 16'd35104, 16'd6958, 16'd40405, 16'd31647, 16'd23014, 16'd36210, 16'd26521, 16'd11647, 16'd25751, 16'd39510, 16'd46922, 16'd65015, 16'd38028, 16'd63952, 16'd38338, 16'd52890, 16'd3702, 16'd15569});
	test_expansion(128'hb76248d00f545cd139354b57a228329a, {16'd20392, 16'd34027, 16'd47961, 16'd20246, 16'd7383, 16'd11260, 16'd62886, 16'd18575, 16'd49145, 16'd23088, 16'd18276, 16'd45610, 16'd14258, 16'd54637, 16'd29153, 16'd55904, 16'd35445, 16'd21405, 16'd63181, 16'd44845, 16'd17009, 16'd63863, 16'd665, 16'd54337, 16'd44552, 16'd34710});
	test_expansion(128'hc15b6b25d78045a6f7f1bc1f1e2262bb, {16'd61203, 16'd59984, 16'd21973, 16'd51917, 16'd51359, 16'd12486, 16'd15430, 16'd34876, 16'd30910, 16'd24085, 16'd58828, 16'd49371, 16'd5340, 16'd50561, 16'd10310, 16'd31721, 16'd18167, 16'd52613, 16'd25569, 16'd58978, 16'd50934, 16'd21743, 16'd4483, 16'd823, 16'd58889, 16'd11911});
	test_expansion(128'h4335b5bb070b48cce95cdf815ba58721, {16'd35755, 16'd14545, 16'd38810, 16'd46444, 16'd45145, 16'd39999, 16'd46086, 16'd60658, 16'd31599, 16'd28842, 16'd23947, 16'd18266, 16'd272, 16'd9125, 16'd30013, 16'd39429, 16'd10102, 16'd57371, 16'd10014, 16'd36186, 16'd23807, 16'd27133, 16'd3675, 16'd52186, 16'd58833, 16'd39568});
	test_expansion(128'hda4dbc7f3a9456320d428c549666d032, {16'd1865, 16'd40186, 16'd55844, 16'd14782, 16'd28147, 16'd38351, 16'd44269, 16'd24402, 16'd33180, 16'd61407, 16'd51071, 16'd28934, 16'd37343, 16'd17712, 16'd19023, 16'd35942, 16'd60190, 16'd51789, 16'd46373, 16'd48248, 16'd6204, 16'd7112, 16'd49157, 16'd30560, 16'd4819, 16'd34428});
	test_expansion(128'h54016a0407494ac23237da16b4ae7b52, {16'd64931, 16'd34631, 16'd15578, 16'd43656, 16'd19870, 16'd53514, 16'd22397, 16'd18415, 16'd19486, 16'd5465, 16'd31983, 16'd54106, 16'd1168, 16'd65226, 16'd24597, 16'd3491, 16'd18340, 16'd18089, 16'd18673, 16'd61921, 16'd48817, 16'd2311, 16'd46383, 16'd57042, 16'd30647, 16'd23449});
	test_expansion(128'he22e3faaeb44b711fe549e702703d54d, {16'd8859, 16'd38873, 16'd15851, 16'd21165, 16'd20617, 16'd12642, 16'd46515, 16'd22830, 16'd28117, 16'd22368, 16'd5297, 16'd24187, 16'd17762, 16'd65300, 16'd19974, 16'd24351, 16'd24597, 16'd64557, 16'd60891, 16'd62208, 16'd7001, 16'd13690, 16'd19467, 16'd44954, 16'd12167, 16'd39513});
	test_expansion(128'h89f14004a0fee6879113f02d3cc66158, {16'd28251, 16'd44806, 16'd26008, 16'd52720, 16'd26638, 16'd16450, 16'd22223, 16'd32428, 16'd62621, 16'd5921, 16'd19866, 16'd40237, 16'd26438, 16'd21009, 16'd30795, 16'd46392, 16'd63538, 16'd51021, 16'd11705, 16'd4213, 16'd36639, 16'd34156, 16'd33142, 16'd14055, 16'd32619, 16'd43328});
	test_expansion(128'h5f992c03a585dcf25b2ebd83b9217e8c, {16'd39499, 16'd7389, 16'd11925, 16'd25077, 16'd44671, 16'd26691, 16'd62945, 16'd20320, 16'd31294, 16'd29403, 16'd34458, 16'd65381, 16'd31816, 16'd409, 16'd6772, 16'd57580, 16'd11030, 16'd28361, 16'd6403, 16'd19717, 16'd57688, 16'd51407, 16'd47746, 16'd2145, 16'd24114, 16'd43609});
	test_expansion(128'h76a2fc56ca641dd69c973342002ebe23, {16'd9022, 16'd58017, 16'd37232, 16'd21315, 16'd52523, 16'd61503, 16'd3339, 16'd13144, 16'd19970, 16'd28505, 16'd20792, 16'd18491, 16'd64242, 16'd2066, 16'd18107, 16'd501, 16'd45846, 16'd5102, 16'd59873, 16'd30388, 16'd63100, 16'd41077, 16'd30462, 16'd11952, 16'd7, 16'd49975});
	test_expansion(128'h7b28a2bcac28b1d427bb65bc869607c8, {16'd51799, 16'd24735, 16'd61897, 16'd6454, 16'd34903, 16'd14822, 16'd62350, 16'd40872, 16'd5919, 16'd11925, 16'd10312, 16'd41889, 16'd42458, 16'd51412, 16'd7224, 16'd60426, 16'd21678, 16'd30058, 16'd47757, 16'd25566, 16'd57775, 16'd60833, 16'd36478, 16'd49022, 16'd60604, 16'd63037});
	test_expansion(128'h3fed7744c6433f5df044d375b0d1879a, {16'd36649, 16'd22823, 16'd1209, 16'd43369, 16'd21906, 16'd26912, 16'd53689, 16'd36552, 16'd13068, 16'd23471, 16'd8622, 16'd26806, 16'd38560, 16'd25725, 16'd42751, 16'd64122, 16'd35929, 16'd25375, 16'd22040, 16'd64512, 16'd32174, 16'd18761, 16'd4240, 16'd64053, 16'd4458, 16'd9810});
	test_expansion(128'hbbbc2098b7a0d26769c6f23d4375bfa9, {16'd4020, 16'd5719, 16'd50194, 16'd16765, 16'd58366, 16'd52459, 16'd35016, 16'd42182, 16'd65385, 16'd12976, 16'd25638, 16'd63771, 16'd17482, 16'd49679, 16'd16126, 16'd63572, 16'd6634, 16'd29629, 16'd57113, 16'd50785, 16'd19399, 16'd23188, 16'd6913, 16'd17580, 16'd41373, 16'd26486});
	test_expansion(128'h91568400006801f5a190eca168321d0f, {16'd12821, 16'd22827, 16'd13342, 16'd42083, 16'd10989, 16'd5476, 16'd17303, 16'd8193, 16'd61360, 16'd48728, 16'd61841, 16'd27344, 16'd44003, 16'd19624, 16'd5231, 16'd13381, 16'd20261, 16'd1096, 16'd51565, 16'd48474, 16'd36086, 16'd50213, 16'd26198, 16'd21671, 16'd40075, 16'd20648});
	test_expansion(128'h920168a2caf120dc3cfd7d3093cc7ba7, {16'd63700, 16'd64997, 16'd42039, 16'd51542, 16'd28699, 16'd64225, 16'd32573, 16'd58413, 16'd60384, 16'd55587, 16'd60496, 16'd60417, 16'd21916, 16'd38449, 16'd24922, 16'd2797, 16'd55746, 16'd42555, 16'd57528, 16'd62070, 16'd8611, 16'd56154, 16'd28739, 16'd23402, 16'd27325, 16'd54028});
	test_expansion(128'hcba140d4ce937f6401d5946eb91ecd4a, {16'd45517, 16'd55552, 16'd61354, 16'd40988, 16'd34848, 16'd55598, 16'd21140, 16'd59932, 16'd64264, 16'd14230, 16'd42016, 16'd50005, 16'd4111, 16'd14393, 16'd12483, 16'd10438, 16'd24697, 16'd46104, 16'd20948, 16'd47824, 16'd4535, 16'd9378, 16'd31569, 16'd32954, 16'd9058, 16'd34172});
	test_expansion(128'hbface74ac065c8a47ebc977aa1215ed6, {16'd64610, 16'd2870, 16'd47952, 16'd62320, 16'd7462, 16'd50036, 16'd55886, 16'd22753, 16'd38567, 16'd9049, 16'd28838, 16'd6442, 16'd5967, 16'd44655, 16'd23901, 16'd53920, 16'd63802, 16'd4417, 16'd13474, 16'd45267, 16'd59533, 16'd60796, 16'd17883, 16'd24950, 16'd42620, 16'd46726});
	test_expansion(128'he5e3d11cef6a54c5609c5965c92bb20f, {16'd37493, 16'd4319, 16'd53084, 16'd21084, 16'd62997, 16'd31387, 16'd63700, 16'd13274, 16'd57570, 16'd1082, 16'd37887, 16'd48084, 16'd20584, 16'd5203, 16'd21385, 16'd48693, 16'd4456, 16'd26937, 16'd62790, 16'd5831, 16'd27326, 16'd51049, 16'd63069, 16'd40225, 16'd15841, 16'd14584});
	test_expansion(128'h37fbbbe4fadd3ba16ba412f71bc6f46f, {16'd36319, 16'd14950, 16'd24743, 16'd54675, 16'd27965, 16'd60648, 16'd5893, 16'd14076, 16'd9822, 16'd24388, 16'd18977, 16'd32320, 16'd46483, 16'd2134, 16'd35303, 16'd44935, 16'd62041, 16'd19878, 16'd57517, 16'd23396, 16'd14565, 16'd53664, 16'd24731, 16'd44950, 16'd23140, 16'd30019});
	test_expansion(128'hf3425ccd0db28c2b79e763c4c406b02a, {16'd43121, 16'd32133, 16'd37297, 16'd10438, 16'd1360, 16'd11355, 16'd49755, 16'd40642, 16'd39574, 16'd9879, 16'd60773, 16'd35496, 16'd7181, 16'd10249, 16'd49534, 16'd21173, 16'd56092, 16'd55496, 16'd50171, 16'd62446, 16'd20317, 16'd31793, 16'd37012, 16'd53407, 16'd18084, 16'd45092});
	test_expansion(128'h97548cf3f50587df3259959ac53a11d3, {16'd17954, 16'd19301, 16'd8278, 16'd15717, 16'd17562, 16'd8356, 16'd62159, 16'd32486, 16'd3047, 16'd27379, 16'd58386, 16'd54285, 16'd47388, 16'd34199, 16'd19188, 16'd3222, 16'd7375, 16'd54574, 16'd32970, 16'd23356, 16'd15942, 16'd9679, 16'd40101, 16'd52362, 16'd39371, 16'd65290});
	test_expansion(128'h230f8f8349cbf7cfd7af9a720b8c8d2f, {16'd56839, 16'd20894, 16'd55997, 16'd55385, 16'd16928, 16'd9995, 16'd30898, 16'd10910, 16'd19276, 16'd21590, 16'd1978, 16'd40856, 16'd16208, 16'd64319, 16'd60213, 16'd64940, 16'd33737, 16'd48811, 16'd15179, 16'd34330, 16'd31631, 16'd63870, 16'd47771, 16'd50319, 16'd24915, 16'd14055});
	test_expansion(128'h771581b516a8e0536a98d20a63ab7aa4, {16'd61004, 16'd44128, 16'd25286, 16'd14871, 16'd14998, 16'd4768, 16'd19077, 16'd30858, 16'd9376, 16'd32432, 16'd11579, 16'd47904, 16'd40673, 16'd22380, 16'd8675, 16'd47094, 16'd41553, 16'd31572, 16'd54090, 16'd51243, 16'd62828, 16'd382, 16'd18169, 16'd61319, 16'd41669, 16'd60307});
	test_expansion(128'hc649f3a52e67da9cbfe3a61872b77991, {16'd31917, 16'd43869, 16'd27874, 16'd21162, 16'd26489, 16'd34272, 16'd13165, 16'd45467, 16'd7160, 16'd45817, 16'd16590, 16'd10208, 16'd56511, 16'd18198, 16'd5420, 16'd17882, 16'd56576, 16'd51272, 16'd8554, 16'd42121, 16'd22702, 16'd22766, 16'd58949, 16'd8736, 16'd32048, 16'd15592});
	test_expansion(128'hedc62b6624988b6cd439693853e37463, {16'd3435, 16'd49796, 16'd245, 16'd494, 16'd37158, 16'd8281, 16'd9103, 16'd19544, 16'd32905, 16'd24729, 16'd9545, 16'd3384, 16'd49556, 16'd62303, 16'd59703, 16'd4695, 16'd59588, 16'd31269, 16'd42315, 16'd17870, 16'd24529, 16'd24259, 16'd57872, 16'd47682, 16'd19721, 16'd9726});
	test_expansion(128'h69a12997e74ba5bc780397a784663513, {16'd28025, 16'd10442, 16'd56579, 16'd25913, 16'd22542, 16'd22002, 16'd34903, 16'd32936, 16'd63856, 16'd44352, 16'd6511, 16'd35438, 16'd11778, 16'd21299, 16'd6826, 16'd25860, 16'd43442, 16'd16941, 16'd42129, 16'd41213, 16'd6366, 16'd18210, 16'd39856, 16'd27940, 16'd47900, 16'd4099});
	test_expansion(128'h63172c76f4aceb5bd256d10c8592511e, {16'd42652, 16'd10903, 16'd10704, 16'd57909, 16'd2934, 16'd8324, 16'd4191, 16'd44067, 16'd3133, 16'd31945, 16'd38353, 16'd21576, 16'd61582, 16'd40861, 16'd13535, 16'd4938, 16'd13192, 16'd29395, 16'd5160, 16'd65404, 16'd50677, 16'd64345, 16'd53093, 16'd15195, 16'd65138, 16'd48612});
	test_expansion(128'h751f8af800f8af7ade0e0672019c3841, {16'd63674, 16'd2998, 16'd59986, 16'd63856, 16'd34842, 16'd29093, 16'd50652, 16'd52503, 16'd12436, 16'd39399, 16'd24313, 16'd62275, 16'd56494, 16'd15076, 16'd16630, 16'd44899, 16'd16406, 16'd2730, 16'd24725, 16'd6488, 16'd22131, 16'd60769, 16'd39877, 16'd46130, 16'd12745, 16'd16934});
	test_expansion(128'h1eabc38dee9439ed4707902524856df1, {16'd18317, 16'd34541, 16'd36373, 16'd55059, 16'd64347, 16'd25961, 16'd33653, 16'd19019, 16'd23326, 16'd13024, 16'd40021, 16'd8711, 16'd19581, 16'd40896, 16'd23000, 16'd40476, 16'd49670, 16'd53089, 16'd5840, 16'd34393, 16'd44098, 16'd62998, 16'd38169, 16'd45404, 16'd63749, 16'd21377});
	test_expansion(128'hd7cb59223cfa28dc50580e8c15febd94, {16'd11090, 16'd6983, 16'd17568, 16'd61774, 16'd51295, 16'd23675, 16'd14107, 16'd21063, 16'd50982, 16'd11649, 16'd34447, 16'd45009, 16'd23526, 16'd37754, 16'd57779, 16'd1977, 16'd15037, 16'd9547, 16'd36033, 16'd1930, 16'd52951, 16'd9847, 16'd37191, 16'd52392, 16'd40765, 16'd274});
	test_expansion(128'h767b1fd261184452664bd64063042655, {16'd30968, 16'd10253, 16'd15873, 16'd25757, 16'd60444, 16'd3024, 16'd10819, 16'd10689, 16'd57923, 16'd14953, 16'd35016, 16'd22258, 16'd17497, 16'd51908, 16'd670, 16'd31225, 16'd8545, 16'd32101, 16'd49149, 16'd23288, 16'd15221, 16'd21729, 16'd59121, 16'd55269, 16'd14523, 16'd8018});
	test_expansion(128'h08289c89ddba01d61e11b980cb944e6c, {16'd49178, 16'd65532, 16'd28080, 16'd65376, 16'd50908, 16'd17681, 16'd35016, 16'd30628, 16'd23739, 16'd20475, 16'd6300, 16'd58144, 16'd56816, 16'd64307, 16'd6532, 16'd27021, 16'd42235, 16'd54325, 16'd54357, 16'd20107, 16'd35769, 16'd23241, 16'd28871, 16'd38817, 16'd35864, 16'd8620});
	test_expansion(128'hc4948e0b22a78eb2e7dbe356cc4fcf17, {16'd60487, 16'd26563, 16'd41995, 16'd4388, 16'd43387, 16'd5186, 16'd34416, 16'd65055, 16'd13499, 16'd53290, 16'd54501, 16'd42529, 16'd29056, 16'd9467, 16'd36387, 16'd18092, 16'd63195, 16'd31843, 16'd11185, 16'd41586, 16'd38773, 16'd64732, 16'd57656, 16'd35140, 16'd14752, 16'd46538});
	test_expansion(128'hd83263a8446cd2351b63e2dcb4d3368a, {16'd54499, 16'd55538, 16'd17801, 16'd39809, 16'd64344, 16'd62835, 16'd14230, 16'd37554, 16'd12546, 16'd15882, 16'd14877, 16'd3277, 16'd51272, 16'd46017, 16'd60368, 16'd58663, 16'd40992, 16'd35352, 16'd18218, 16'd36512, 16'd58801, 16'd47916, 16'd30734, 16'd12642, 16'd53700, 16'd52929});
	test_expansion(128'hdb16f30925d33e931e6838e014d5a986, {16'd11541, 16'd34588, 16'd41502, 16'd3347, 16'd37363, 16'd368, 16'd47233, 16'd24797, 16'd57671, 16'd50031, 16'd46337, 16'd18698, 16'd32585, 16'd44820, 16'd35619, 16'd39205, 16'd6700, 16'd65152, 16'd41058, 16'd490, 16'd47912, 16'd29550, 16'd42191, 16'd44288, 16'd30834, 16'd58207});
	test_expansion(128'h3b7c844b44b921e6ba5f17383bce2e1c, {16'd15951, 16'd59990, 16'd42816, 16'd35510, 16'd43295, 16'd30336, 16'd51537, 16'd59235, 16'd31975, 16'd14552, 16'd10017, 16'd11562, 16'd65034, 16'd27171, 16'd19375, 16'd33561, 16'd59938, 16'd40781, 16'd25337, 16'd33604, 16'd25084, 16'd49389, 16'd21669, 16'd54054, 16'd62257, 16'd44781});
	test_expansion(128'h46bf4545bfb6ff7db6d54592f4f82a0d, {16'd37678, 16'd27523, 16'd26284, 16'd52228, 16'd8521, 16'd56382, 16'd24342, 16'd62083, 16'd12525, 16'd49065, 16'd6248, 16'd7524, 16'd24433, 16'd47915, 16'd30044, 16'd9835, 16'd29720, 16'd12802, 16'd15803, 16'd40922, 16'd8426, 16'd33818, 16'd5423, 16'd52292, 16'd44625, 16'd58905});
	test_expansion(128'h1438054274f8ce0a090ebcf962f4db7d, {16'd49796, 16'd61492, 16'd51138, 16'd15422, 16'd23441, 16'd28397, 16'd6364, 16'd65335, 16'd15963, 16'd63588, 16'd51922, 16'd65058, 16'd7686, 16'd54795, 16'd46956, 16'd8298, 16'd6145, 16'd38464, 16'd65230, 16'd28006, 16'd55332, 16'd33710, 16'd27767, 16'd44871, 16'd36430, 16'd39843});
	test_expansion(128'h8c25d518e1eb61186397bef60a0139ad, {16'd15216, 16'd56286, 16'd59082, 16'd60859, 16'd37032, 16'd37701, 16'd53137, 16'd48308, 16'd960, 16'd8970, 16'd6975, 16'd32135, 16'd55840, 16'd53706, 16'd44659, 16'd48574, 16'd52400, 16'd42740, 16'd56959, 16'd48063, 16'd42898, 16'd34458, 16'd40748, 16'd55416, 16'd4915, 16'd23262});
	test_expansion(128'h76a9ee27ed5fd07750ce6f7dd4076bf5, {16'd12514, 16'd18737, 16'd28969, 16'd25998, 16'd24443, 16'd50782, 16'd25224, 16'd19812, 16'd49406, 16'd36084, 16'd59432, 16'd1042, 16'd46550, 16'd11013, 16'd62578, 16'd42189, 16'd25825, 16'd16817, 16'd61346, 16'd35685, 16'd28241, 16'd39100, 16'd54819, 16'd39086, 16'd22585, 16'd54354});
	test_expansion(128'hbcafe25e8db06484ee5bca4e04c37984, {16'd15428, 16'd63131, 16'd58549, 16'd16287, 16'd8917, 16'd61146, 16'd22261, 16'd26006, 16'd11672, 16'd29350, 16'd53590, 16'd27365, 16'd16545, 16'd1065, 16'd18500, 16'd25909, 16'd17586, 16'd16343, 16'd18226, 16'd52749, 16'd4026, 16'd47681, 16'd34927, 16'd20526, 16'd20332, 16'd46568});
	test_expansion(128'ha40455145d7c1b273820b449012dfa01, {16'd26921, 16'd41287, 16'd14167, 16'd53353, 16'd23566, 16'd24570, 16'd56425, 16'd60837, 16'd20026, 16'd42622, 16'd22228, 16'd53423, 16'd27663, 16'd29851, 16'd14895, 16'd41008, 16'd33765, 16'd3908, 16'd3143, 16'd36456, 16'd20538, 16'd5305, 16'd60947, 16'd4771, 16'd42423, 16'd50265});
	test_expansion(128'h91ff0d6bd6f5b280c39d3a0c1d58b1c6, {16'd35487, 16'd10966, 16'd11308, 16'd34810, 16'd27606, 16'd30848, 16'd14317, 16'd62930, 16'd60240, 16'd15713, 16'd57564, 16'd50238, 16'd13004, 16'd65183, 16'd56468, 16'd21123, 16'd24379, 16'd11346, 16'd19328, 16'd12870, 16'd11474, 16'd19265, 16'd17505, 16'd20036, 16'd42765, 16'd9863});
	test_expansion(128'h4dc0dbd7d10be65db7c26305a0ea4571, {16'd28147, 16'd34970, 16'd55076, 16'd40047, 16'd62025, 16'd44805, 16'd25850, 16'd4089, 16'd26021, 16'd47078, 16'd5361, 16'd2131, 16'd8710, 16'd23965, 16'd28617, 16'd64146, 16'd53288, 16'd27228, 16'd3722, 16'd3532, 16'd46498, 16'd34566, 16'd32511, 16'd34043, 16'd64367, 16'd16286});
	test_expansion(128'h70a3e4d7dace0475327ce2441f7b9cab, {16'd36342, 16'd33513, 16'd37421, 16'd9499, 16'd56918, 16'd62503, 16'd23339, 16'd23160, 16'd22819, 16'd45641, 16'd58619, 16'd23451, 16'd53141, 16'd9244, 16'd4750, 16'd14503, 16'd35699, 16'd51680, 16'd24825, 16'd8464, 16'd33054, 16'd10384, 16'd39136, 16'd26551, 16'd29517, 16'd8553});
	test_expansion(128'h471b07886fc57267ead86da6c07dfc08, {16'd19210, 16'd61833, 16'd3028, 16'd54689, 16'd35583, 16'd60495, 16'd44895, 16'd43247, 16'd29190, 16'd16416, 16'd9407, 16'd35260, 16'd58356, 16'd41585, 16'd35217, 16'd31689, 16'd61798, 16'd60798, 16'd50780, 16'd29633, 16'd63932, 16'd42321, 16'd13647, 16'd48751, 16'd40147, 16'd6720});
	test_expansion(128'h502d4d120c341406cfb6744e90c0db4d, {16'd49700, 16'd45868, 16'd4811, 16'd13554, 16'd3677, 16'd11769, 16'd55105, 16'd15217, 16'd38510, 16'd18081, 16'd44283, 16'd22603, 16'd53896, 16'd59797, 16'd25620, 16'd56987, 16'd12163, 16'd44258, 16'd31172, 16'd19705, 16'd44353, 16'd62627, 16'd24623, 16'd57940, 16'd20758, 16'd54062});
	test_expansion(128'h806f92c8529d0c966374f18f30802014, {16'd23625, 16'd34129, 16'd51042, 16'd27113, 16'd41783, 16'd54776, 16'd594, 16'd21097, 16'd8660, 16'd65285, 16'd47813, 16'd53200, 16'd48021, 16'd14213, 16'd19723, 16'd19956, 16'd53925, 16'd59594, 16'd50409, 16'd23669, 16'd39568, 16'd658, 16'd34041, 16'd30343, 16'd51453, 16'd21518});
	test_expansion(128'hd928a4cb90172b8929f63439d9aca5a5, {16'd55412, 16'd42737, 16'd58141, 16'd35987, 16'd62133, 16'd38621, 16'd26421, 16'd37598, 16'd20808, 16'd52881, 16'd46865, 16'd47502, 16'd27283, 16'd4673, 16'd2173, 16'd31762, 16'd20540, 16'd25867, 16'd56204, 16'd53458, 16'd2296, 16'd16556, 16'd41315, 16'd12857, 16'd16705, 16'd64295});
	test_expansion(128'h44834ebf0e9256e9a77ad734b3b279bb, {16'd35508, 16'd5723, 16'd40317, 16'd42844, 16'd5447, 16'd60776, 16'd48044, 16'd34589, 16'd17306, 16'd29199, 16'd37460, 16'd4845, 16'd24876, 16'd18837, 16'd26464, 16'd37355, 16'd14103, 16'd32763, 16'd36703, 16'd27439, 16'd55681, 16'd58420, 16'd21153, 16'd42414, 16'd33817, 16'd62246});
	test_expansion(128'h861f658ba58d69fba588c84123977b95, {16'd29067, 16'd3349, 16'd7833, 16'd32802, 16'd24137, 16'd10180, 16'd53347, 16'd24121, 16'd64729, 16'd52195, 16'd48743, 16'd21011, 16'd42798, 16'd61093, 16'd16857, 16'd16577, 16'd64048, 16'd49952, 16'd10820, 16'd41398, 16'd15565, 16'd1167, 16'd17257, 16'd26334, 16'd43967, 16'd40655});
	test_expansion(128'h42804ed6f175d0741b08666256995f44, {16'd65376, 16'd45311, 16'd3595, 16'd49407, 16'd17739, 16'd61052, 16'd12466, 16'd29679, 16'd63479, 16'd63616, 16'd631, 16'd8500, 16'd39178, 16'd14380, 16'd29717, 16'd11419, 16'd15884, 16'd29605, 16'd14066, 16'd38090, 16'd21374, 16'd52265, 16'd38638, 16'd14162, 16'd64000, 16'd10349});
	test_expansion(128'h5fce336ab5c31c7879d24d574c9d7a45, {16'd42759, 16'd5827, 16'd52293, 16'd52475, 16'd9453, 16'd12863, 16'd35058, 16'd64731, 16'd39071, 16'd32294, 16'd40784, 16'd20652, 16'd21032, 16'd49066, 16'd46834, 16'd48611, 16'd31733, 16'd20861, 16'd54380, 16'd46395, 16'd22377, 16'd10585, 16'd28966, 16'd5543, 16'd64338, 16'd23284});
	test_expansion(128'he23a6c02805b5c0b12961b8ae1d73abe, {16'd26458, 16'd35306, 16'd38864, 16'd5983, 16'd12063, 16'd14414, 16'd42625, 16'd35519, 16'd47968, 16'd8100, 16'd60539, 16'd51777, 16'd1300, 16'd3695, 16'd51211, 16'd13520, 16'd31242, 16'd28064, 16'd57887, 16'd57943, 16'd43743, 16'd41158, 16'd7807, 16'd64125, 16'd64145, 16'd46154});
	test_expansion(128'hac998762bce6a63204d1af27591d64c7, {16'd29121, 16'd450, 16'd8697, 16'd33608, 16'd6000, 16'd56387, 16'd55910, 16'd47110, 16'd32482, 16'd29266, 16'd6287, 16'd21344, 16'd63534, 16'd28542, 16'd58583, 16'd28905, 16'd54845, 16'd42487, 16'd8969, 16'd15138, 16'd21043, 16'd26515, 16'd18805, 16'd8965, 16'd4496, 16'd63041});
	test_expansion(128'ha8adbdd725c7f16fb6b693a3cbe951b4, {16'd33452, 16'd23908, 16'd38070, 16'd13867, 16'd61981, 16'd10130, 16'd18637, 16'd26318, 16'd13108, 16'd3093, 16'd28885, 16'd5888, 16'd43764, 16'd63928, 16'd18711, 16'd56830, 16'd10809, 16'd10181, 16'd53322, 16'd29376, 16'd31820, 16'd57811, 16'd47035, 16'd62981, 16'd9655, 16'd28691});
	test_expansion(128'h899c0ec55a89324150fa09d49c23be78, {16'd1987, 16'd24144, 16'd38837, 16'd22072, 16'd62900, 16'd38769, 16'd37741, 16'd35596, 16'd58761, 16'd27082, 16'd39599, 16'd13629, 16'd48571, 16'd27153, 16'd30345, 16'd44806, 16'd30204, 16'd48593, 16'd43838, 16'd6255, 16'd46970, 16'd58755, 16'd53938, 16'd31990, 16'd10178, 16'd58727});
	test_expansion(128'hf6bc15b753d22e9819a0a13c8f892b7d, {16'd44811, 16'd14506, 16'd49942, 16'd12585, 16'd35111, 16'd61129, 16'd59443, 16'd39340, 16'd53542, 16'd48750, 16'd53337, 16'd21292, 16'd10919, 16'd16027, 16'd33931, 16'd22247, 16'd14110, 16'd25160, 16'd29698, 16'd15058, 16'd7019, 16'd55573, 16'd31364, 16'd2065, 16'd29891, 16'd18931});
	test_expansion(128'h6d05b4cfcd18d8a45d2888a187733484, {16'd45240, 16'd42116, 16'd13879, 16'd53321, 16'd27130, 16'd52005, 16'd31049, 16'd63847, 16'd20582, 16'd30754, 16'd10312, 16'd57888, 16'd7623, 16'd4760, 16'd3099, 16'd3700, 16'd40943, 16'd7477, 16'd55686, 16'd43092, 16'd18025, 16'd36513, 16'd11959, 16'd42452, 16'd16452, 16'd10202});
	test_expansion(128'ha713512f76c73136656495465ab10a5c, {16'd55252, 16'd41152, 16'd63372, 16'd31338, 16'd19805, 16'd26483, 16'd28010, 16'd32333, 16'd52960, 16'd65073, 16'd56773, 16'd41682, 16'd16239, 16'd29977, 16'd40033, 16'd36726, 16'd18782, 16'd64861, 16'd42984, 16'd42282, 16'd12823, 16'd18989, 16'd10368, 16'd3006, 16'd2428, 16'd29694});
	test_expansion(128'h126b4a54012d2f58ab5cf37dd144fedc, {16'd52530, 16'd48381, 16'd51517, 16'd8948, 16'd16492, 16'd56288, 16'd54706, 16'd17584, 16'd14452, 16'd27568, 16'd31896, 16'd22482, 16'd11841, 16'd25207, 16'd16162, 16'd52243, 16'd65422, 16'd47093, 16'd31359, 16'd43822, 16'd28318, 16'd51300, 16'd2184, 16'd31080, 16'd7703, 16'd41015});
	test_expansion(128'h72c459498b94ca800d257da828a9d4f4, {16'd14318, 16'd28570, 16'd30223, 16'd34015, 16'd24, 16'd23385, 16'd30913, 16'd2527, 16'd6742, 16'd25629, 16'd6979, 16'd38606, 16'd15949, 16'd3889, 16'd5307, 16'd10701, 16'd32302, 16'd16743, 16'd33056, 16'd29845, 16'd40175, 16'd14346, 16'd6969, 16'd1918, 16'd47597, 16'd52326});
	test_expansion(128'hab8a0b07231e87c58704124002895817, {16'd44763, 16'd15217, 16'd47489, 16'd24937, 16'd7177, 16'd48398, 16'd32365, 16'd11035, 16'd50237, 16'd13317, 16'd60925, 16'd30921, 16'd5469, 16'd38212, 16'd63228, 16'd64700, 16'd26747, 16'd49628, 16'd25329, 16'd63531, 16'd12505, 16'd56976, 16'd41570, 16'd57760, 16'd49544, 16'd16887});
	test_expansion(128'hea8ba07825ce4872607f83aa09458dea, {16'd57229, 16'd46793, 16'd60680, 16'd44219, 16'd1473, 16'd60108, 16'd56989, 16'd24090, 16'd22577, 16'd50395, 16'd44607, 16'd18724, 16'd53996, 16'd48912, 16'd20584, 16'd1870, 16'd6615, 16'd52710, 16'd61375, 16'd43021, 16'd6981, 16'd6842, 16'd64419, 16'd40415, 16'd3879, 16'd33806});
	test_expansion(128'h8bcbd0323810ffec605789f75918376f, {16'd61348, 16'd38533, 16'd48589, 16'd34, 16'd37389, 16'd58806, 16'd51796, 16'd35273, 16'd54889, 16'd20779, 16'd31646, 16'd61228, 16'd8133, 16'd39738, 16'd49816, 16'd60405, 16'd22351, 16'd53696, 16'd14207, 16'd40154, 16'd13802, 16'd14567, 16'd49816, 16'd18792, 16'd12129, 16'd37878});
	test_expansion(128'h169068eb149eb971afe9fb31c74406b9, {16'd36113, 16'd18962, 16'd15176, 16'd64259, 16'd35372, 16'd40367, 16'd54063, 16'd31898, 16'd11717, 16'd38711, 16'd17012, 16'd21375, 16'd14891, 16'd58203, 16'd18402, 16'd35505, 16'd50065, 16'd7441, 16'd48718, 16'd26974, 16'd38053, 16'd63088, 16'd60943, 16'd36172, 16'd10417, 16'd10633});
	test_expansion(128'h672ddde65312192bca09e2ac789b838e, {16'd6939, 16'd15490, 16'd62460, 16'd25918, 16'd21631, 16'd7948, 16'd12034, 16'd45144, 16'd8952, 16'd19337, 16'd62946, 16'd9349, 16'd20897, 16'd2444, 16'd25858, 16'd17395, 16'd64402, 16'd19979, 16'd47790, 16'd37821, 16'd42937, 16'd30, 16'd30322, 16'd1866, 16'd22683, 16'd60445});
	test_expansion(128'hb4efde2c2a406bd0dd8c07488731a63a, {16'd58987, 16'd9003, 16'd39326, 16'd41163, 16'd51069, 16'd25173, 16'd30305, 16'd31322, 16'd44375, 16'd5356, 16'd14486, 16'd40699, 16'd33628, 16'd894, 16'd21437, 16'd62601, 16'd43611, 16'd36415, 16'd32820, 16'd62577, 16'd13800, 16'd18150, 16'd36640, 16'd56643, 16'd3286, 16'd27038});
	test_expansion(128'h5b037f2f044a71e38c66075ce474ff8a, {16'd32112, 16'd20478, 16'd59560, 16'd35257, 16'd62875, 16'd38892, 16'd37579, 16'd27081, 16'd49517, 16'd33857, 16'd16644, 16'd25528, 16'd31831, 16'd37119, 16'd43554, 16'd40480, 16'd11307, 16'd64392, 16'd15960, 16'd29045, 16'd40711, 16'd24938, 16'd62773, 16'd41134, 16'd30147, 16'd34692});
	test_expansion(128'hb9a5e90b59873595859f0e63186f271d, {16'd28210, 16'd46918, 16'd59159, 16'd21221, 16'd41393, 16'd15527, 16'd6746, 16'd18699, 16'd34181, 16'd23480, 16'd34134, 16'd29706, 16'd20209, 16'd58652, 16'd20239, 16'd11649, 16'd8022, 16'd23778, 16'd35229, 16'd10204, 16'd16157, 16'd36952, 16'd53197, 16'd28687, 16'd63945, 16'd47162});
	test_expansion(128'h5c5e2e42b9be2921337d6da97b630500, {16'd38350, 16'd39435, 16'd50301, 16'd34761, 16'd51069, 16'd25422, 16'd47221, 16'd20745, 16'd23915, 16'd63605, 16'd24020, 16'd40545, 16'd26987, 16'd15610, 16'd58402, 16'd9778, 16'd62749, 16'd26138, 16'd7238, 16'd17378, 16'd12828, 16'd63483, 16'd51848, 16'd15167, 16'd26267, 16'd26543});
	test_expansion(128'ha1c66ce64f5525eb7d563907aa6cba15, {16'd21028, 16'd44790, 16'd27447, 16'd47370, 16'd47767, 16'd5185, 16'd33208, 16'd19273, 16'd15869, 16'd3090, 16'd30375, 16'd49123, 16'd8004, 16'd10687, 16'd58118, 16'd8745, 16'd44311, 16'd29966, 16'd62148, 16'd36484, 16'd32717, 16'd38361, 16'd41667, 16'd25632, 16'd56637, 16'd16890});
	test_expansion(128'h03e810bb85efb27c4f702d8865c6603d, {16'd16579, 16'd3876, 16'd33906, 16'd33884, 16'd39157, 16'd9380, 16'd9155, 16'd34439, 16'd64985, 16'd1837, 16'd23425, 16'd29235, 16'd17732, 16'd30309, 16'd40193, 16'd46740, 16'd63257, 16'd58883, 16'd16450, 16'd53535, 16'd350, 16'd61060, 16'd60588, 16'd43193, 16'd12567, 16'd11084});
	test_expansion(128'hd77cbb5ce50b33718fa14340753b3829, {16'd20178, 16'd15037, 16'd5393, 16'd13965, 16'd65008, 16'd32425, 16'd47180, 16'd39309, 16'd36660, 16'd14043, 16'd14476, 16'd49247, 16'd46032, 16'd44338, 16'd37897, 16'd36678, 16'd61208, 16'd16953, 16'd50728, 16'd18914, 16'd5220, 16'd16006, 16'd18407, 16'd51931, 16'd32018, 16'd9447});
	test_expansion(128'h046ff3b40cde3c8b6233689a6e1563f0, {16'd15257, 16'd39187, 16'd43313, 16'd39903, 16'd48942, 16'd47442, 16'd18617, 16'd9903, 16'd59694, 16'd48209, 16'd53367, 16'd26032, 16'd8608, 16'd28304, 16'd3749, 16'd13969, 16'd52847, 16'd36084, 16'd14619, 16'd17657, 16'd46543, 16'd51106, 16'd10119, 16'd61474, 16'd11146, 16'd2390});
	test_expansion(128'h6d7de71c735b19937c2f763e42b8c84c, {16'd64596, 16'd20310, 16'd56971, 16'd8773, 16'd28863, 16'd56046, 16'd8507, 16'd21617, 16'd20253, 16'd13819, 16'd44046, 16'd24684, 16'd7793, 16'd15877, 16'd30097, 16'd28618, 16'd34708, 16'd38907, 16'd49042, 16'd56781, 16'd46746, 16'd55467, 16'd17063, 16'd55014, 16'd41817, 16'd27068});
	test_expansion(128'h5fb62888b3e2abe10341e1771ba987f8, {16'd45365, 16'd36968, 16'd65376, 16'd62060, 16'd35997, 16'd33831, 16'd52368, 16'd48305, 16'd25843, 16'd43373, 16'd7806, 16'd62720, 16'd19933, 16'd701, 16'd55426, 16'd28874, 16'd29784, 16'd18002, 16'd43354, 16'd20678, 16'd54289, 16'd59110, 16'd23563, 16'd22458, 16'd26379, 16'd62761});
	test_expansion(128'hc6ec902880fb5ed81acc06b250ac43da, {16'd37581, 16'd42069, 16'd5246, 16'd27516, 16'd44171, 16'd13827, 16'd21440, 16'd40294, 16'd41831, 16'd60001, 16'd26852, 16'd17635, 16'd63479, 16'd57040, 16'd25106, 16'd35792, 16'd35048, 16'd64670, 16'd19083, 16'd17792, 16'd18578, 16'd13399, 16'd54942, 16'd28204, 16'd56363, 16'd17142});
	test_expansion(128'h2833ee94236b0ebbf7299f2868053009, {16'd2842, 16'd4379, 16'd11817, 16'd5129, 16'd58807, 16'd25318, 16'd63714, 16'd34425, 16'd1978, 16'd15362, 16'd33534, 16'd15173, 16'd62669, 16'd3768, 16'd24241, 16'd3413, 16'd47617, 16'd60879, 16'd34057, 16'd14523, 16'd2513, 16'd484, 16'd29716, 16'd27047, 16'd61086, 16'd24841});
	test_expansion(128'ha5d2ecac7e6908edd937028628d75996, {16'd25815, 16'd23981, 16'd19257, 16'd1083, 16'd22326, 16'd40163, 16'd57867, 16'd53857, 16'd61774, 16'd11766, 16'd63461, 16'd29895, 16'd59376, 16'd21210, 16'd55893, 16'd15933, 16'd6357, 16'd44069, 16'd44703, 16'd31885, 16'd45303, 16'd20913, 16'd55287, 16'd15977, 16'd9835, 16'd17514});
	test_expansion(128'h895eccd4fb2f1bd854a31e56fd4bb6b0, {16'd9540, 16'd47232, 16'd348, 16'd55366, 16'd59145, 16'd39870, 16'd41790, 16'd19583, 16'd55228, 16'd45948, 16'd64842, 16'd32635, 16'd47033, 16'd26534, 16'd34475, 16'd48134, 16'd37488, 16'd41968, 16'd18704, 16'd38624, 16'd46256, 16'd40581, 16'd48198, 16'd21430, 16'd52160, 16'd44951});
	test_expansion(128'h40268f6787c1f708068cbbd66bb4f12d, {16'd2375, 16'd33711, 16'd49889, 16'd6625, 16'd31280, 16'd20089, 16'd8860, 16'd39047, 16'd35905, 16'd58578, 16'd64103, 16'd33514, 16'd4146, 16'd49944, 16'd40812, 16'd57840, 16'd57372, 16'd7420, 16'd30999, 16'd48356, 16'd61413, 16'd36745, 16'd43308, 16'd16462, 16'd34271, 16'd8215});
	test_expansion(128'ha1e5103a0bb5c717d3661c45cb95eb45, {16'd1064, 16'd34458, 16'd64901, 16'd20965, 16'd4774, 16'd53840, 16'd58002, 16'd14305, 16'd24422, 16'd32911, 16'd4431, 16'd36143, 16'd56487, 16'd12852, 16'd63738, 16'd6951, 16'd1508, 16'd43300, 16'd22096, 16'd1681, 16'd60390, 16'd16426, 16'd47746, 16'd38712, 16'd25521, 16'd15843});
	test_expansion(128'h92718b4eea3d392cea7154b11e0dce7e, {16'd22918, 16'd47531, 16'd35360, 16'd42803, 16'd16100, 16'd31540, 16'd20539, 16'd7237, 16'd16885, 16'd56595, 16'd48090, 16'd9886, 16'd17338, 16'd27736, 16'd10389, 16'd56456, 16'd15717, 16'd2192, 16'd28510, 16'd39618, 16'd8230, 16'd14161, 16'd48333, 16'd13774, 16'd18210, 16'd3092});
	test_expansion(128'hf3032af7bc376e1c0996559519fd6a80, {16'd23006, 16'd57059, 16'd27514, 16'd33058, 16'd51100, 16'd27730, 16'd16087, 16'd20313, 16'd19490, 16'd21705, 16'd48079, 16'd938, 16'd41812, 16'd29654, 16'd47449, 16'd46195, 16'd41684, 16'd44520, 16'd5157, 16'd8123, 16'd9984, 16'd38506, 16'd8101, 16'd39500, 16'd51890, 16'd30421});
	test_expansion(128'h8872439e10029d395d06204aa6daa331, {16'd11177, 16'd49410, 16'd20781, 16'd4139, 16'd7001, 16'd42971, 16'd59981, 16'd33183, 16'd20798, 16'd25413, 16'd33042, 16'd60926, 16'd38193, 16'd36217, 16'd36710, 16'd24957, 16'd28990, 16'd15365, 16'd37828, 16'd31885, 16'd62044, 16'd36575, 16'd44060, 16'd33038, 16'd6290, 16'd17201});
	test_expansion(128'hcf51d9b3d3ca6edbe0dad7fea98f521d, {16'd18995, 16'd20323, 16'd61706, 16'd8979, 16'd37546, 16'd61684, 16'd18584, 16'd18857, 16'd50810, 16'd9479, 16'd49719, 16'd26057, 16'd34676, 16'd47183, 16'd59507, 16'd21202, 16'd8177, 16'd56508, 16'd62913, 16'd33525, 16'd43465, 16'd41481, 16'd5783, 16'd8140, 16'd34910, 16'd9338});
	test_expansion(128'h4e88329dfd419a2366b6ab85233d6d6f, {16'd36893, 16'd47757, 16'd42221, 16'd60945, 16'd50562, 16'd30190, 16'd37199, 16'd2113, 16'd25260, 16'd56485, 16'd25288, 16'd55438, 16'd60863, 16'd27907, 16'd43060, 16'd45692, 16'd8334, 16'd51040, 16'd59110, 16'd60449, 16'd53770, 16'd9604, 16'd62541, 16'd37826, 16'd63612, 16'd55034});
	test_expansion(128'h2b79feacf861e76f85c91d5def5ae451, {16'd40583, 16'd12139, 16'd26799, 16'd58196, 16'd13472, 16'd11976, 16'd38914, 16'd13345, 16'd9234, 16'd12343, 16'd6034, 16'd2675, 16'd33691, 16'd15211, 16'd20185, 16'd48570, 16'd50950, 16'd41180, 16'd64785, 16'd25697, 16'd59439, 16'd27937, 16'd56980, 16'd344, 16'd11814, 16'd59671});
	test_expansion(128'h94b4a8d390a4b9f70a82003d905842bf, {16'd49742, 16'd37287, 16'd9769, 16'd5962, 16'd2557, 16'd51053, 16'd55219, 16'd891, 16'd15633, 16'd17232, 16'd63349, 16'd58608, 16'd33293, 16'd4827, 16'd14475, 16'd58802, 16'd15196, 16'd19883, 16'd46011, 16'd48726, 16'd3675, 16'd18958, 16'd28140, 16'd24104, 16'd23183, 16'd37613});
	test_expansion(128'hd123fb0d1a94d82f990085c9e45762ef, {16'd46857, 16'd20454, 16'd26268, 16'd31821, 16'd9111, 16'd11515, 16'd5450, 16'd45644, 16'd27314, 16'd14108, 16'd22934, 16'd6119, 16'd28437, 16'd49072, 16'd54529, 16'd41346, 16'd42225, 16'd33258, 16'd52904, 16'd61506, 16'd25227, 16'd18105, 16'd46515, 16'd31236, 16'd20734, 16'd13850});
	test_expansion(128'ha68d197af86e5dc90c448dad326450ff, {16'd50272, 16'd37218, 16'd8566, 16'd47842, 16'd34955, 16'd46229, 16'd20564, 16'd2733, 16'd5172, 16'd54155, 16'd35631, 16'd44078, 16'd60749, 16'd57392, 16'd53104, 16'd10579, 16'd16581, 16'd61326, 16'd168, 16'd19562, 16'd49375, 16'd17551, 16'd27884, 16'd17121, 16'd6077, 16'd41231});
	test_expansion(128'he94165ce63d7f69a723b3988756154cf, {16'd60965, 16'd65053, 16'd39680, 16'd36566, 16'd26360, 16'd51293, 16'd10228, 16'd44197, 16'd15774, 16'd26336, 16'd11146, 16'd11918, 16'd50293, 16'd30501, 16'd16209, 16'd47972, 16'd26318, 16'd33823, 16'd52740, 16'd6073, 16'd38498, 16'd48083, 16'd19875, 16'd36979, 16'd37932, 16'd43897});
	test_expansion(128'h0c71797bdab5abab8683c053e8ea032c, {16'd19053, 16'd32468, 16'd52211, 16'd59677, 16'd59015, 16'd57742, 16'd30380, 16'd7081, 16'd56427, 16'd19955, 16'd3656, 16'd30591, 16'd54441, 16'd49708, 16'd46897, 16'd5414, 16'd63217, 16'd3388, 16'd58816, 16'd50454, 16'd1345, 16'd7854, 16'd29101, 16'd61513, 16'd62257, 16'd49333});
	test_expansion(128'he5146bdade326bdc336d9a892196b478, {16'd18343, 16'd61447, 16'd63678, 16'd39430, 16'd44570, 16'd33777, 16'd16860, 16'd11397, 16'd41657, 16'd32415, 16'd33793, 16'd8196, 16'd60494, 16'd10867, 16'd55412, 16'd35626, 16'd57911, 16'd10934, 16'd32534, 16'd12956, 16'd20236, 16'd31841, 16'd61975, 16'd1492, 16'd34089, 16'd22406});
	test_expansion(128'hce98ce7c3a6d35949bf0bb6e1c3f515c, {16'd64242, 16'd54824, 16'd62306, 16'd41467, 16'd54169, 16'd26124, 16'd55626, 16'd19050, 16'd53409, 16'd51568, 16'd45473, 16'd43554, 16'd50923, 16'd215, 16'd1494, 16'd56046, 16'd46210, 16'd50788, 16'd63102, 16'd44264, 16'd40367, 16'd29957, 16'd37799, 16'd53808, 16'd18359, 16'd47692});
	test_expansion(128'hfc8ae45994abe6a63b05c79080c2dfe1, {16'd65339, 16'd17493, 16'd46117, 16'd64759, 16'd36591, 16'd6155, 16'd26320, 16'd41827, 16'd33705, 16'd53679, 16'd46716, 16'd24386, 16'd39448, 16'd20150, 16'd11428, 16'd34454, 16'd16825, 16'd30352, 16'd44391, 16'd57681, 16'd31521, 16'd21789, 16'd3602, 16'd59031, 16'd27654, 16'd63007});
	test_expansion(128'hf443761adaa3c36ee3dfc943f2c6b0d1, {16'd41505, 16'd55642, 16'd8204, 16'd57281, 16'd10308, 16'd57364, 16'd34848, 16'd14977, 16'd28902, 16'd23164, 16'd33152, 16'd34579, 16'd36432, 16'd31240, 16'd56326, 16'd31922, 16'd42057, 16'd6216, 16'd6778, 16'd57931, 16'd64818, 16'd17674, 16'd58568, 16'd31747, 16'd61706, 16'd3442});
	test_expansion(128'hdb799b52c8414a690e0f0295b12bb3b7, {16'd57962, 16'd34259, 16'd45385, 16'd26635, 16'd32948, 16'd55645, 16'd2767, 16'd27426, 16'd7469, 16'd20632, 16'd40455, 16'd41609, 16'd57201, 16'd30319, 16'd36221, 16'd56815, 16'd23785, 16'd63017, 16'd46413, 16'd44857, 16'd31345, 16'd45754, 16'd52807, 16'd13266, 16'd8913, 16'd24244});
	test_expansion(128'h8a3f2062accfd43d4f332fdeac432273, {16'd46484, 16'd41120, 16'd30396, 16'd28461, 16'd62121, 16'd25476, 16'd24574, 16'd63609, 16'd24813, 16'd30566, 16'd38313, 16'd52635, 16'd15433, 16'd48670, 16'd21920, 16'd23672, 16'd61726, 16'd39608, 16'd28656, 16'd52700, 16'd32210, 16'd1350, 16'd25543, 16'd646, 16'd56996, 16'd57760});
	test_expansion(128'had58791edf8ab9c40067a4b8a9f3412f, {16'd51758, 16'd36025, 16'd1149, 16'd20319, 16'd1463, 16'd40387, 16'd15053, 16'd41567, 16'd60851, 16'd2082, 16'd49410, 16'd23880, 16'd30858, 16'd3776, 16'd13004, 16'd12191, 16'd49041, 16'd65103, 16'd9239, 16'd7059, 16'd37765, 16'd435, 16'd45073, 16'd62985, 16'd17867, 16'd10972});
	test_expansion(128'ha6fe368fc65e3580ae4e3b140521fcbe, {16'd36661, 16'd52575, 16'd58430, 16'd65421, 16'd46626, 16'd1263, 16'd12872, 16'd4995, 16'd25794, 16'd10980, 16'd6226, 16'd18990, 16'd35346, 16'd59093, 16'd28768, 16'd51362, 16'd13169, 16'd15940, 16'd32807, 16'd39500, 16'd2984, 16'd43836, 16'd55632, 16'd11507, 16'd28753, 16'd46442});
	test_expansion(128'h377a02c9967bac6854c475690b295c60, {16'd19965, 16'd1459, 16'd20496, 16'd52997, 16'd37092, 16'd45285, 16'd50809, 16'd48878, 16'd8883, 16'd60271, 16'd25458, 16'd22561, 16'd16192, 16'd6265, 16'd13270, 16'd62936, 16'd6855, 16'd21888, 16'd55326, 16'd49587, 16'd38729, 16'd19696, 16'd61617, 16'd11878, 16'd55167, 16'd49394});
	test_expansion(128'hbd00ff0cace085902d3f9f8aac3e9a33, {16'd64357, 16'd16608, 16'd19180, 16'd4627, 16'd3215, 16'd45041, 16'd26202, 16'd25648, 16'd28907, 16'd3641, 16'd51619, 16'd8661, 16'd15791, 16'd29062, 16'd11752, 16'd1492, 16'd7628, 16'd8222, 16'd57004, 16'd1940, 16'd43850, 16'd52197, 16'd21271, 16'd51955, 16'd23154, 16'd61837});
	test_expansion(128'h48ea9e6b1c78aa5d376846a8830b2327, {16'd32442, 16'd11365, 16'd33630, 16'd13213, 16'd14526, 16'd36676, 16'd65487, 16'd33479, 16'd26359, 16'd49546, 16'd36833, 16'd35046, 16'd53029, 16'd59188, 16'd22451, 16'd2755, 16'd60263, 16'd30962, 16'd39198, 16'd12481, 16'd63906, 16'd32036, 16'd10999, 16'd45178, 16'd65081, 16'd4776});
	test_expansion(128'h67351898414e0c2d8d65b2157858ca14, {16'd22727, 16'd61291, 16'd35354, 16'd11900, 16'd49943, 16'd36339, 16'd11962, 16'd48561, 16'd14492, 16'd38189, 16'd47093, 16'd30617, 16'd63887, 16'd30183, 16'd42715, 16'd19281, 16'd29487, 16'd26134, 16'd45275, 16'd56334, 16'd36355, 16'd23432, 16'd17446, 16'd42966, 16'd29834, 16'd14515});
	test_expansion(128'h83b00125492bbe8cf6249745c317f904, {16'd65348, 16'd48299, 16'd14835, 16'd6907, 16'd36933, 16'd22495, 16'd33059, 16'd22594, 16'd59669, 16'd9890, 16'd58836, 16'd25688, 16'd5335, 16'd35088, 16'd50742, 16'd64074, 16'd20704, 16'd30292, 16'd11042, 16'd51862, 16'd42261, 16'd13130, 16'd55852, 16'd28433, 16'd62790, 16'd9788});
	test_expansion(128'h312b2a6a64703baa8e8e61d58416ce04, {16'd41801, 16'd39157, 16'd37635, 16'd33262, 16'd26937, 16'd31320, 16'd60247, 16'd2930, 16'd27144, 16'd53612, 16'd4317, 16'd42437, 16'd60662, 16'd19435, 16'd32439, 16'd8, 16'd11230, 16'd39362, 16'd26401, 16'd7066, 16'd16188, 16'd53143, 16'd14252, 16'd59974, 16'd26519, 16'd50977});
	test_expansion(128'h4dd0c50124ceb4df61ff581786af2f5b, {16'd62614, 16'd26755, 16'd3710, 16'd45659, 16'd18469, 16'd5386, 16'd11138, 16'd41382, 16'd3991, 16'd53295, 16'd16730, 16'd18202, 16'd10856, 16'd14469, 16'd36395, 16'd30399, 16'd37222, 16'd4341, 16'd26943, 16'd9796, 16'd63414, 16'd3658, 16'd33710, 16'd62808, 16'd32259, 16'd46073});
	test_expansion(128'h8db3461abf5a53162442b7c7dbdbff18, {16'd20527, 16'd44904, 16'd51691, 16'd63295, 16'd40442, 16'd26328, 16'd10608, 16'd42377, 16'd550, 16'd10095, 16'd58649, 16'd7520, 16'd54777, 16'd50335, 16'd45702, 16'd44793, 16'd26696, 16'd28467, 16'd16356, 16'd1641, 16'd47836, 16'd19117, 16'd59321, 16'd34662, 16'd3673, 16'd40977});
	test_expansion(128'h8d73669e729149471622d58c02d727dd, {16'd3391, 16'd51301, 16'd223, 16'd31425, 16'd29823, 16'd43249, 16'd21060, 16'd25173, 16'd47093, 16'd50852, 16'd24344, 16'd26244, 16'd55635, 16'd60099, 16'd42616, 16'd34475, 16'd38477, 16'd7240, 16'd26844, 16'd38070, 16'd15661, 16'd32547, 16'd35805, 16'd50620, 16'd36009, 16'd59839});
	test_expansion(128'h81a9c80e180961a27c59e7bc48e6f92e, {16'd60870, 16'd17357, 16'd45202, 16'd49610, 16'd3947, 16'd31447, 16'd37750, 16'd39803, 16'd62501, 16'd57005, 16'd59606, 16'd41955, 16'd21037, 16'd53528, 16'd42550, 16'd7082, 16'd24541, 16'd8566, 16'd44432, 16'd5295, 16'd7194, 16'd60597, 16'd14145, 16'd41451, 16'd26465, 16'd2741});
	test_expansion(128'hd0095caefa05222972ec2c1b5e5d67c2, {16'd62595, 16'd62451, 16'd2984, 16'd34446, 16'd64415, 16'd17394, 16'd1006, 16'd37126, 16'd51921, 16'd21294, 16'd53874, 16'd49407, 16'd14681, 16'd53587, 16'd16530, 16'd64014, 16'd61438, 16'd35015, 16'd5518, 16'd46747, 16'd1730, 16'd23989, 16'd36047, 16'd7182, 16'd17160, 16'd28160});
	test_expansion(128'h22e511453d6ba0e494ff6c9081e1baff, {16'd37558, 16'd43943, 16'd20784, 16'd50422, 16'd1828, 16'd48573, 16'd49467, 16'd27349, 16'd12491, 16'd27443, 16'd13903, 16'd57621, 16'd58245, 16'd47524, 16'd22955, 16'd54812, 16'd19590, 16'd4041, 16'd28056, 16'd6429, 16'd6118, 16'd50229, 16'd20433, 16'd9098, 16'd55220, 16'd59580});
	test_expansion(128'h99385f6b3d195c9de91d006d6c846792, {16'd29685, 16'd45427, 16'd18540, 16'd4130, 16'd33816, 16'd13804, 16'd35273, 16'd16659, 16'd58213, 16'd5710, 16'd16518, 16'd57342, 16'd53584, 16'd29228, 16'd38531, 16'd35616, 16'd47008, 16'd37061, 16'd52408, 16'd55473, 16'd2841, 16'd9946, 16'd26905, 16'd20459, 16'd54892, 16'd23857});
	test_expansion(128'h1925882afffed13495f1f2f030b75273, {16'd275, 16'd58702, 16'd25634, 16'd34091, 16'd24211, 16'd39752, 16'd2862, 16'd11060, 16'd6600, 16'd43965, 16'd53823, 16'd65530, 16'd25887, 16'd11340, 16'd7307, 16'd57729, 16'd46249, 16'd8440, 16'd19921, 16'd5326, 16'd49281, 16'd44468, 16'd24648, 16'd15225, 16'd164, 16'd30859});
	test_expansion(128'h6028c2a08a22cc4168302997c8d1f508, {16'd65444, 16'd8708, 16'd1109, 16'd31990, 16'd12337, 16'd9650, 16'd16101, 16'd40307, 16'd14132, 16'd34105, 16'd6862, 16'd35077, 16'd25941, 16'd57500, 16'd51191, 16'd50854, 16'd60086, 16'd29201, 16'd1080, 16'd4443, 16'd11891, 16'd55718, 16'd31776, 16'd27320, 16'd48312, 16'd22677});
	test_expansion(128'hcbdf43cd708512cb84ffd63b1050d2d4, {16'd54891, 16'd10542, 16'd39029, 16'd19591, 16'd12849, 16'd43848, 16'd23367, 16'd57170, 16'd4957, 16'd26545, 16'd37014, 16'd60442, 16'd35740, 16'd33807, 16'd43735, 16'd58750, 16'd11651, 16'd42650, 16'd59792, 16'd2601, 16'd32863, 16'd43629, 16'd46662, 16'd24249, 16'd20864, 16'd46431});
	test_expansion(128'h016c264653a02f31a4f8582a8969ea40, {16'd61733, 16'd24898, 16'd63764, 16'd65197, 16'd3809, 16'd37379, 16'd26345, 16'd37825, 16'd33103, 16'd45091, 16'd54622, 16'd35586, 16'd65405, 16'd43580, 16'd21592, 16'd54785, 16'd37706, 16'd34391, 16'd6904, 16'd17208, 16'd9468, 16'd938, 16'd32024, 16'd33662, 16'd6472, 16'd57882});
	test_expansion(128'h14f45100b27f494856bd85a958287149, {16'd56036, 16'd59067, 16'd54400, 16'd14864, 16'd16553, 16'd50868, 16'd7849, 16'd22142, 16'd19065, 16'd16576, 16'd34992, 16'd34664, 16'd65185, 16'd62521, 16'd56850, 16'd11267, 16'd50502, 16'd39617, 16'd60286, 16'd23913, 16'd38023, 16'd35590, 16'd19686, 16'd5465, 16'd54084, 16'd29910});
	test_expansion(128'hb38cb746a8bc0b6805855f3dfa2404fe, {16'd16252, 16'd38281, 16'd21724, 16'd13584, 16'd5354, 16'd5057, 16'd3639, 16'd53288, 16'd11902, 16'd55999, 16'd51691, 16'd12586, 16'd32818, 16'd58002, 16'd14871, 16'd62022, 16'd44965, 16'd51086, 16'd38335, 16'd7520, 16'd42076, 16'd44843, 16'd6838, 16'd41716, 16'd6498, 16'd30550});
	test_expansion(128'h888550bd51832fbfa25623409368aa0c, {16'd56226, 16'd34726, 16'd14138, 16'd1895, 16'd53638, 16'd14323, 16'd22652, 16'd55549, 16'd44573, 16'd29469, 16'd4478, 16'd63828, 16'd20255, 16'd64341, 16'd51274, 16'd26547, 16'd8409, 16'd37959, 16'd43237, 16'd49727, 16'd11898, 16'd16697, 16'd18441, 16'd33415, 16'd54694, 16'd130});
	test_expansion(128'hff749077128b2eb5b6d3658b9596ad98, {16'd16733, 16'd32682, 16'd63641, 16'd27150, 16'd2600, 16'd40939, 16'd63994, 16'd45484, 16'd26629, 16'd34745, 16'd22686, 16'd1183, 16'd49412, 16'd62023, 16'd3074, 16'd39434, 16'd35098, 16'd236, 16'd60340, 16'd40101, 16'd22636, 16'd26699, 16'd61588, 16'd5944, 16'd47286, 16'd54765});
	test_expansion(128'ha763b6f7f8afbc6562bdb1cde1d286c3, {16'd23669, 16'd2720, 16'd40222, 16'd61359, 16'd45695, 16'd578, 16'd7517, 16'd47652, 16'd59410, 16'd950, 16'd7897, 16'd3236, 16'd38122, 16'd33855, 16'd65404, 16'd11635, 16'd18321, 16'd16175, 16'd59215, 16'd13793, 16'd52310, 16'd59491, 16'd47926, 16'd36816, 16'd20325, 16'd59295});
	test_expansion(128'h084b4ec3ef8c39e24dc96a5be5702a3f, {16'd44144, 16'd9491, 16'd8949, 16'd64491, 16'd32922, 16'd51557, 16'd61486, 16'd27163, 16'd7903, 16'd36417, 16'd59118, 16'd45392, 16'd26195, 16'd25519, 16'd36478, 16'd25429, 16'd41609, 16'd29973, 16'd47152, 16'd59746, 16'd37195, 16'd34280, 16'd51911, 16'd63581, 16'd4060, 16'd3334});
	test_expansion(128'ha162c161d843698dedfd884e121d114e, {16'd15506, 16'd44716, 16'd32081, 16'd40738, 16'd65034, 16'd56840, 16'd63815, 16'd61726, 16'd27043, 16'd4438, 16'd21070, 16'd30980, 16'd53769, 16'd34979, 16'd29921, 16'd26102, 16'd12060, 16'd27188, 16'd32290, 16'd23533, 16'd52428, 16'd52072, 16'd59883, 16'd14388, 16'd19560, 16'd52480});
	test_expansion(128'h73a9586f2a1dd2c550a4543ee2e9d951, {16'd47217, 16'd15228, 16'd40447, 16'd27634, 16'd37056, 16'd54024, 16'd28803, 16'd17110, 16'd23967, 16'd10303, 16'd7933, 16'd34202, 16'd7331, 16'd6786, 16'd63171, 16'd40333, 16'd58450, 16'd53199, 16'd51957, 16'd57377, 16'd5478, 16'd5945, 16'd65008, 16'd34638, 16'd41664, 16'd55520});
	test_expansion(128'h0c599e68930b8d72e1a5b40632e935de, {16'd15727, 16'd38525, 16'd58533, 16'd38288, 16'd7592, 16'd36880, 16'd64902, 16'd3254, 16'd20598, 16'd42620, 16'd32792, 16'd3476, 16'd17004, 16'd21926, 16'd47234, 16'd36802, 16'd59863, 16'd49371, 16'd25387, 16'd5897, 16'd41791, 16'd60097, 16'd11285, 16'd51192, 16'd59022, 16'd34993});
	test_expansion(128'hce1988b5db6781224a7b06470c689b01, {16'd53055, 16'd13987, 16'd21244, 16'd43267, 16'd32520, 16'd24997, 16'd57016, 16'd45863, 16'd42896, 16'd381, 16'd31673, 16'd2643, 16'd42358, 16'd39618, 16'd43537, 16'd31093, 16'd15202, 16'd22248, 16'd44733, 16'd14748, 16'd22137, 16'd43638, 16'd5858, 16'd48766, 16'd22321, 16'd1734});
	test_expansion(128'h5258d6ed33c589b5abaf50621026e724, {16'd52180, 16'd6133, 16'd29814, 16'd12001, 16'd3566, 16'd48827, 16'd58978, 16'd45424, 16'd65238, 16'd34827, 16'd39765, 16'd59913, 16'd58947, 16'd40479, 16'd53425, 16'd3746, 16'd7113, 16'd10760, 16'd33732, 16'd23726, 16'd38447, 16'd23805, 16'd691, 16'd58722, 16'd62213, 16'd45660});
	test_expansion(128'hafd3b01a243180ef0c116a2ed022dd0c, {16'd27008, 16'd42328, 16'd40739, 16'd37138, 16'd40160, 16'd30126, 16'd17787, 16'd18546, 16'd43386, 16'd36070, 16'd53251, 16'd6404, 16'd13526, 16'd64583, 16'd31828, 16'd15255, 16'd13893, 16'd54819, 16'd18274, 16'd10655, 16'd4203, 16'd3367, 16'd40266, 16'd674, 16'd47327, 16'd10245});
	test_expansion(128'h9dfcbe470535a4aa60450675468743a8, {16'd62555, 16'd65134, 16'd15133, 16'd63904, 16'd42972, 16'd7317, 16'd2104, 16'd6415, 16'd4809, 16'd1842, 16'd43137, 16'd21251, 16'd5387, 16'd55464, 16'd18568, 16'd13131, 16'd30122, 16'd42135, 16'd17067, 16'd27088, 16'd34332, 16'd31797, 16'd41617, 16'd28894, 16'd38563, 16'd40895});
	test_expansion(128'he960f9566b85892bc5346b4dfa52eca4, {16'd37873, 16'd24911, 16'd28855, 16'd40869, 16'd49973, 16'd38524, 16'd16976, 16'd28332, 16'd43002, 16'd63676, 16'd9501, 16'd49115, 16'd22087, 16'd11357, 16'd57070, 16'd50972, 16'd21386, 16'd62999, 16'd65340, 16'd9046, 16'd33504, 16'd28899, 16'd65375, 16'd17434, 16'd10014, 16'd46170});
	test_expansion(128'h0f33fde6f6c185c544c8dffffd4a6efb, {16'd61777, 16'd37592, 16'd28586, 16'd54512, 16'd64216, 16'd33109, 16'd65377, 16'd47481, 16'd9916, 16'd27952, 16'd59707, 16'd44138, 16'd29265, 16'd12856, 16'd7607, 16'd60461, 16'd26927, 16'd23910, 16'd42584, 16'd63236, 16'd9907, 16'd14978, 16'd45996, 16'd43498, 16'd7565, 16'd53379});
	test_expansion(128'hb269d107c5d499b703f89ed0100d67eb, {16'd51104, 16'd57469, 16'd31126, 16'd41582, 16'd10357, 16'd59054, 16'd29201, 16'd15978, 16'd15937, 16'd25408, 16'd54071, 16'd17167, 16'd64209, 16'd47316, 16'd17675, 16'd28755, 16'd48847, 16'd61595, 16'd61384, 16'd7366, 16'd20303, 16'd49803, 16'd16972, 16'd20815, 16'd36118, 16'd16});
	test_expansion(128'h759b09ff55900db35169c6eb179aa180, {16'd961, 16'd42232, 16'd23023, 16'd1455, 16'd27307, 16'd40345, 16'd17396, 16'd15863, 16'd17593, 16'd50020, 16'd8247, 16'd26696, 16'd40370, 16'd55070, 16'd12075, 16'd35055, 16'd36545, 16'd59105, 16'd63016, 16'd9947, 16'd40648, 16'd62220, 16'd27762, 16'd60642, 16'd56498, 16'd42147});
	test_expansion(128'h2e539f5e1f3121dbf1e6b7a17b49c2af, {16'd18216, 16'd56649, 16'd56675, 16'd4286, 16'd3416, 16'd36216, 16'd10477, 16'd42604, 16'd63970, 16'd45189, 16'd57334, 16'd55382, 16'd49989, 16'd4294, 16'd36075, 16'd55389, 16'd57425, 16'd37715, 16'd28445, 16'd4561, 16'd13550, 16'd4154, 16'd4379, 16'd49213, 16'd41932, 16'd20823});
	test_expansion(128'h092ee9ea43b322b2a39cc9d2891cc130, {16'd18189, 16'd25503, 16'd33324, 16'd44321, 16'd58630, 16'd32946, 16'd35564, 16'd1813, 16'd3560, 16'd57803, 16'd22064, 16'd62191, 16'd60993, 16'd31342, 16'd48609, 16'd46201, 16'd63612, 16'd42037, 16'd61432, 16'd32611, 16'd35787, 16'd19893, 16'd5179, 16'd35720, 16'd15328, 16'd2315});
	test_expansion(128'h94c157d879e91b2bb2f009c4d52ab6e4, {16'd4513, 16'd3129, 16'd13713, 16'd10217, 16'd46592, 16'd61976, 16'd15575, 16'd10406, 16'd30594, 16'd18566, 16'd31506, 16'd10200, 16'd20918, 16'd20092, 16'd26883, 16'd52495, 16'd770, 16'd11949, 16'd12165, 16'd28296, 16'd65226, 16'd58015, 16'd31544, 16'd5417, 16'd51487, 16'd36603});
	test_expansion(128'heff8fb02fd0fd9259e543f302822401f, {16'd57529, 16'd12776, 16'd9198, 16'd37944, 16'd60852, 16'd29630, 16'd31807, 16'd45328, 16'd34778, 16'd23921, 16'd24931, 16'd35422, 16'd23360, 16'd30065, 16'd30277, 16'd45916, 16'd8899, 16'd28399, 16'd9201, 16'd39175, 16'd2862, 16'd55309, 16'd60338, 16'd43446, 16'd55496, 16'd13439});
	test_expansion(128'h28195c5c06f133362d5cd9840908cc1d, {16'd35076, 16'd39976, 16'd34155, 16'd1626, 16'd64222, 16'd7553, 16'd31924, 16'd24410, 16'd40107, 16'd47804, 16'd53335, 16'd47768, 16'd44041, 16'd9634, 16'd57803, 16'd45708, 16'd60695, 16'd54489, 16'd37153, 16'd36213, 16'd24001, 16'd19642, 16'd56635, 16'd65188, 16'd18628, 16'd26504});
	test_expansion(128'h92b640ba0eb9259f5b11f1a79e9fa997, {16'd16941, 16'd64225, 16'd46120, 16'd64376, 16'd60045, 16'd57438, 16'd14078, 16'd3517, 16'd53111, 16'd19914, 16'd10437, 16'd26142, 16'd50115, 16'd48621, 16'd51235, 16'd42966, 16'd63538, 16'd59001, 16'd33144, 16'd58126, 16'd56445, 16'd7770, 16'd45809, 16'd28982, 16'd769, 16'd40841});
	test_expansion(128'h05e87c3f60bcde6091b95a15b5f310f8, {16'd24545, 16'd9280, 16'd58526, 16'd18900, 16'd34836, 16'd56415, 16'd44343, 16'd50208, 16'd47443, 16'd7090, 16'd53535, 16'd62715, 16'd50701, 16'd40435, 16'd39738, 16'd6339, 16'd50964, 16'd27069, 16'd33713, 16'd22741, 16'd48297, 16'd17302, 16'd51666, 16'd10774, 16'd26195, 16'd4587});
	test_expansion(128'hff9b958923d67266dba12358c694366e, {16'd35631, 16'd18563, 16'd48417, 16'd30514, 16'd46199, 16'd58665, 16'd63520, 16'd22565, 16'd38650, 16'd26607, 16'd47515, 16'd21707, 16'd20509, 16'd44970, 16'd10775, 16'd2303, 16'd43559, 16'd31942, 16'd49654, 16'd24229, 16'd50916, 16'd19294, 16'd50010, 16'd54137, 16'd7167, 16'd32582});
	test_expansion(128'h5826fd8aa309313cb0ced509f17c6d72, {16'd40917, 16'd41685, 16'd58549, 16'd14551, 16'd19373, 16'd18310, 16'd36645, 16'd49628, 16'd45624, 16'd8753, 16'd3376, 16'd3788, 16'd6233, 16'd25682, 16'd47697, 16'd62004, 16'd5835, 16'd25187, 16'd33137, 16'd4557, 16'd53019, 16'd13070, 16'd27766, 16'd27179, 16'd16271, 16'd29042});
	test_expansion(128'h560308bf9fc788780066fa4592e9ec70, {16'd20477, 16'd8388, 16'd46921, 16'd46275, 16'd8227, 16'd5347, 16'd40328, 16'd40019, 16'd21879, 16'd59323, 16'd64155, 16'd19105, 16'd23044, 16'd20420, 16'd4893, 16'd24806, 16'd31524, 16'd24455, 16'd59176, 16'd22346, 16'd63576, 16'd21460, 16'd4260, 16'd50345, 16'd27145, 16'd43110});
	test_expansion(128'h42702526c75fefd9babb7fe49db965c3, {16'd23356, 16'd11880, 16'd60886, 16'd13562, 16'd14543, 16'd56882, 16'd37941, 16'd28145, 16'd57483, 16'd57737, 16'd7388, 16'd38967, 16'd53707, 16'd20319, 16'd10696, 16'd7564, 16'd12312, 16'd36859, 16'd31990, 16'd1504, 16'd8701, 16'd55485, 16'd13371, 16'd7023, 16'd12173, 16'd47334});
	test_expansion(128'h5f61d340d8f7ca6b0953ca95a7353976, {16'd4530, 16'd16510, 16'd55077, 16'd50569, 16'd39690, 16'd10853, 16'd57370, 16'd64806, 16'd18712, 16'd11305, 16'd9688, 16'd26886, 16'd65388, 16'd58806, 16'd44069, 16'd2697, 16'd33426, 16'd5567, 16'd45301, 16'd46679, 16'd60627, 16'd11753, 16'd48911, 16'd15145, 16'd39044, 16'd50222});
	test_expansion(128'h07e634315effa5238a68a2e10fb1f61e, {16'd33212, 16'd2874, 16'd45522, 16'd65031, 16'd38772, 16'd52897, 16'd56268, 16'd49265, 16'd39308, 16'd58395, 16'd1899, 16'd43012, 16'd8584, 16'd27827, 16'd30129, 16'd19314, 16'd33562, 16'd3519, 16'd61907, 16'd22895, 16'd3532, 16'd37460, 16'd48705, 16'd44184, 16'd61902, 16'd22108});
	test_expansion(128'haa02de448522f01942e97bb7093bb4dd, {16'd20159, 16'd19708, 16'd65280, 16'd801, 16'd29743, 16'd25296, 16'd9741, 16'd50839, 16'd59701, 16'd24561, 16'd60700, 16'd38449, 16'd34011, 16'd61284, 16'd50414, 16'd19904, 16'd60875, 16'd3996, 16'd42420, 16'd63970, 16'd25030, 16'd43761, 16'd63022, 16'd44744, 16'd47637, 16'd45861});
	test_expansion(128'h9ee7d1edea4e050ce43aa1d50fa8ab1d, {16'd6772, 16'd58878, 16'd62466, 16'd15515, 16'd6535, 16'd2712, 16'd52941, 16'd3143, 16'd6097, 16'd12525, 16'd15043, 16'd64999, 16'd61952, 16'd14334, 16'd58155, 16'd26638, 16'd23304, 16'd15652, 16'd30984, 16'd61989, 16'd39267, 16'd48680, 16'd54585, 16'd35179, 16'd65291, 16'd24968});
	test_expansion(128'h6757449704388196b67001f5125f0df8, {16'd45235, 16'd6503, 16'd10047, 16'd60999, 16'd22876, 16'd56149, 16'd11255, 16'd46566, 16'd8747, 16'd5820, 16'd60444, 16'd37358, 16'd2169, 16'd8081, 16'd64276, 16'd64992, 16'd3275, 16'd9795, 16'd5164, 16'd36934, 16'd25185, 16'd28099, 16'd47846, 16'd46213, 16'd56604, 16'd12763});
	test_expansion(128'hf88535a4af1176cf2e51edad9d518be2, {16'd15648, 16'd4042, 16'd23278, 16'd59936, 16'd17854, 16'd44905, 16'd32119, 16'd58657, 16'd13886, 16'd4464, 16'd27842, 16'd31560, 16'd25586, 16'd22153, 16'd36424, 16'd16664, 16'd26226, 16'd31545, 16'd3262, 16'd5281, 16'd5086, 16'd14034, 16'd44490, 16'd63064, 16'd40637, 16'd23947});
	test_expansion(128'h0f82195f38494cf6aec2286007efc010, {16'd32844, 16'd17818, 16'd42144, 16'd53963, 16'd40102, 16'd56203, 16'd9347, 16'd602, 16'd37547, 16'd38295, 16'd41184, 16'd63774, 16'd20380, 16'd55348, 16'd3005, 16'd22502, 16'd30720, 16'd27471, 16'd8194, 16'd38790, 16'd13834, 16'd56149, 16'd31181, 16'd5766, 16'd51878, 16'd17998});
	test_expansion(128'h5498e88683af1abf71ee19c13f32f129, {16'd39094, 16'd49143, 16'd61650, 16'd13132, 16'd64884, 16'd33769, 16'd4195, 16'd64903, 16'd1581, 16'd13721, 16'd64417, 16'd8449, 16'd41921, 16'd2392, 16'd33734, 16'd55193, 16'd42338, 16'd23644, 16'd43966, 16'd38444, 16'd30464, 16'd31849, 16'd27557, 16'd4835, 16'd27777, 16'd64837});
	test_expansion(128'hb221f4c7c9fadd06db9d02ce8352d996, {16'd23067, 16'd3818, 16'd18931, 16'd34697, 16'd51848, 16'd13374, 16'd39450, 16'd21892, 16'd9049, 16'd63200, 16'd19930, 16'd38244, 16'd28183, 16'd45418, 16'd48361, 16'd52245, 16'd23462, 16'd11043, 16'd59020, 16'd12892, 16'd24888, 16'd49495, 16'd65137, 16'd44494, 16'd41913, 16'd57444});
	test_expansion(128'hf4abf47765f181f180d6bca70d8f304a, {16'd38847, 16'd34638, 16'd23433, 16'd2683, 16'd41001, 16'd18439, 16'd60234, 16'd29246, 16'd36235, 16'd17804, 16'd14977, 16'd34599, 16'd41529, 16'd46694, 16'd28180, 16'd27350, 16'd16689, 16'd59388, 16'd7442, 16'd20867, 16'd17729, 16'd2928, 16'd2103, 16'd20066, 16'd39190, 16'd12263});
	test_expansion(128'h4f47dd500518054d027475986ea9afe3, {16'd1739, 16'd21201, 16'd14583, 16'd60006, 16'd274, 16'd4828, 16'd54168, 16'd29379, 16'd18188, 16'd63770, 16'd51621, 16'd11133, 16'd27759, 16'd35973, 16'd45081, 16'd18536, 16'd35832, 16'd59998, 16'd21323, 16'd21117, 16'd51483, 16'd33540, 16'd22706, 16'd17424, 16'd62427, 16'd41871});
	test_expansion(128'hfe0e48d6985b95e27896d058f665d788, {16'd43491, 16'd63295, 16'd21858, 16'd38513, 16'd47057, 16'd47871, 16'd751, 16'd20677, 16'd3348, 16'd45107, 16'd37407, 16'd60523, 16'd23010, 16'd21055, 16'd3067, 16'd37299, 16'd332, 16'd41306, 16'd21745, 16'd3313, 16'd23499, 16'd782, 16'd50428, 16'd7352, 16'd57493, 16'd54270});
	test_expansion(128'hb00bf3fb18b2a16315c2a0c6adb789c4, {16'd29062, 16'd37649, 16'd133, 16'd63129, 16'd13533, 16'd2276, 16'd51263, 16'd55677, 16'd3226, 16'd46258, 16'd3028, 16'd53432, 16'd23687, 16'd19337, 16'd10419, 16'd45861, 16'd64096, 16'd33668, 16'd56156, 16'd60101, 16'd33163, 16'd43315, 16'd22226, 16'd34490, 16'd5731, 16'd3264});
	test_expansion(128'hc5d6ac20ab1468b075ce5290e8f7443c, {16'd47833, 16'd45670, 16'd63583, 16'd177, 16'd37696, 16'd62616, 16'd21110, 16'd52152, 16'd26217, 16'd15779, 16'd39096, 16'd57084, 16'd39348, 16'd4740, 16'd61103, 16'd51556, 16'd48960, 16'd12377, 16'd47724, 16'd38332, 16'd41275, 16'd42434, 16'd29366, 16'd7791, 16'd5487, 16'd29445});
	test_expansion(128'h6574e31bb64bf4431278117abe5a73df, {16'd3361, 16'd50157, 16'd54277, 16'd53927, 16'd23653, 16'd4782, 16'd61075, 16'd28397, 16'd64952, 16'd7431, 16'd14600, 16'd30978, 16'd62866, 16'd13264, 16'd34126, 16'd62273, 16'd54795, 16'd38960, 16'd18991, 16'd36452, 16'd53247, 16'd32094, 16'd22951, 16'd26657, 16'd9630, 16'd54940});
	test_expansion(128'h6569b43a68252c0a3c62bb7900250c41, {16'd57837, 16'd18582, 16'd11846, 16'd22718, 16'd2218, 16'd50383, 16'd46095, 16'd24419, 16'd46836, 16'd50294, 16'd5112, 16'd51884, 16'd61303, 16'd39068, 16'd2659, 16'd25508, 16'd3652, 16'd53499, 16'd4297, 16'd35527, 16'd17950, 16'd47341, 16'd43701, 16'd4998, 16'd21779, 16'd24769});
	test_expansion(128'hbe0e42b01f49f864c13dbe5c96f92c80, {16'd11540, 16'd27960, 16'd42794, 16'd30007, 16'd17745, 16'd65152, 16'd50479, 16'd26604, 16'd17251, 16'd29874, 16'd22156, 16'd60289, 16'd29131, 16'd46188, 16'd51214, 16'd14721, 16'd20849, 16'd54774, 16'd13555, 16'd5504, 16'd36523, 16'd62983, 16'd54614, 16'd27383, 16'd11095, 16'd19989});
	test_expansion(128'h1a21137a8803c7b53735c90fa93f8ac3, {16'd37130, 16'd10588, 16'd30519, 16'd29016, 16'd40166, 16'd37461, 16'd32888, 16'd23004, 16'd60259, 16'd2600, 16'd31183, 16'd49839, 16'd45130, 16'd5432, 16'd10048, 16'd22528, 16'd39786, 16'd12112, 16'd56804, 16'd44137, 16'd36512, 16'd11145, 16'd62758, 16'd62834, 16'd17488, 16'd33483});
	test_expansion(128'h2db3a15ebcd7c1941db8aa26e3db2683, {16'd48432, 16'd37556, 16'd16021, 16'd61889, 16'd7442, 16'd63416, 16'd60398, 16'd53526, 16'd56695, 16'd39768, 16'd53373, 16'd26720, 16'd31016, 16'd48864, 16'd6747, 16'd22454, 16'd40871, 16'd54532, 16'd21730, 16'd28027, 16'd15732, 16'd39165, 16'd27292, 16'd46050, 16'd23459, 16'd45804});
	test_expansion(128'hb3fd2639ed40a7a860635823cfd456ae, {16'd60455, 16'd36293, 16'd55678, 16'd7260, 16'd6004, 16'd8503, 16'd38401, 16'd29682, 16'd40734, 16'd7545, 16'd43679, 16'd44270, 16'd24394, 16'd27353, 16'd720, 16'd62916, 16'd13788, 16'd2428, 16'd45043, 16'd51530, 16'd14640, 16'd65024, 16'd63492, 16'd62705, 16'd42658, 16'd42912});
	test_expansion(128'h0b139252162f44691e1f975e75b65a74, {16'd14145, 16'd2934, 16'd39183, 16'd59174, 16'd31090, 16'd42929, 16'd41019, 16'd16844, 16'd46331, 16'd61556, 16'd55723, 16'd58845, 16'd38093, 16'd11621, 16'd11543, 16'd33988, 16'd44749, 16'd52042, 16'd48317, 16'd9705, 16'd561, 16'd20700, 16'd15094, 16'd42442, 16'd29796, 16'd28301});
	test_expansion(128'hbc4c63119651cd9cc8cd961f13ddb778, {16'd44700, 16'd52610, 16'd44926, 16'd49659, 16'd7296, 16'd33107, 16'd43735, 16'd47938, 16'd22700, 16'd22100, 16'd37824, 16'd22628, 16'd63174, 16'd41369, 16'd55057, 16'd36659, 16'd31598, 16'd40760, 16'd42262, 16'd49219, 16'd5430, 16'd60275, 16'd21323, 16'd19529, 16'd51240, 16'd64637});
	test_expansion(128'h08d8272bdc3a41e347e018e916a4afa9, {16'd63415, 16'd35711, 16'd28270, 16'd60514, 16'd649, 16'd43661, 16'd13900, 16'd63295, 16'd54978, 16'd61733, 16'd7874, 16'd3879, 16'd59174, 16'd39972, 16'd11988, 16'd54467, 16'd33922, 16'd16893, 16'd10026, 16'd21329, 16'd11870, 16'd61794, 16'd38967, 16'd11255, 16'd16630, 16'd26451});
	test_expansion(128'he21b5367e40a0cce9dfad00fcfab2192, {16'd49502, 16'd3265, 16'd37448, 16'd24891, 16'd3755, 16'd7952, 16'd56213, 16'd45152, 16'd42904, 16'd32315, 16'd46288, 16'd23613, 16'd283, 16'd45335, 16'd20761, 16'd24277, 16'd13658, 16'd15805, 16'd30576, 16'd7493, 16'd49558, 16'd15114, 16'd15076, 16'd59617, 16'd64839, 16'd16692});
	test_expansion(128'h0f7a5d7578dbdd3c39e73e2e9f321682, {16'd48007, 16'd4336, 16'd155, 16'd59639, 16'd38512, 16'd45024, 16'd42229, 16'd29978, 16'd63380, 16'd33440, 16'd57825, 16'd33546, 16'd45845, 16'd21660, 16'd2245, 16'd22141, 16'd63760, 16'd55672, 16'd2127, 16'd8483, 16'd56803, 16'd55544, 16'd16386, 16'd13866, 16'd65121, 16'd53169});
	test_expansion(128'h922187d75682aa0108173ae4389fe3f6, {16'd39854, 16'd53878, 16'd45260, 16'd9396, 16'd22319, 16'd17630, 16'd52212, 16'd38625, 16'd10821, 16'd46908, 16'd5410, 16'd27710, 16'd14525, 16'd6333, 16'd61067, 16'd10198, 16'd53563, 16'd47874, 16'd10649, 16'd6006, 16'd1638, 16'd40452, 16'd27342, 16'd57862, 16'd54960, 16'd54642});
	test_expansion(128'h45a3cc6a5b60d710114cefaf15dbd323, {16'd7968, 16'd8744, 16'd37049, 16'd49365, 16'd35433, 16'd16883, 16'd41736, 16'd2072, 16'd8455, 16'd42859, 16'd42861, 16'd56128, 16'd55323, 16'd14003, 16'd13353, 16'd56118, 16'd50186, 16'd711, 16'd1515, 16'd22729, 16'd25806, 16'd63661, 16'd13279, 16'd27937, 16'd49034, 16'd10692});
	test_expansion(128'h14517ab8451a0112794383003bca7cad, {16'd25648, 16'd8566, 16'd54154, 16'd11091, 16'd14390, 16'd26004, 16'd275, 16'd40699, 16'd20466, 16'd35206, 16'd51120, 16'd9379, 16'd40508, 16'd20782, 16'd8400, 16'd33637, 16'd64142, 16'd31633, 16'd49213, 16'd62989, 16'd48, 16'd8970, 16'd24365, 16'd61996, 16'd29800, 16'd20993});
	test_expansion(128'hdf42fa07248bd70c9627019806d1e272, {16'd36352, 16'd46002, 16'd41587, 16'd49828, 16'd31555, 16'd46154, 16'd17, 16'd37850, 16'd58172, 16'd5888, 16'd65065, 16'd34369, 16'd16648, 16'd21382, 16'd33621, 16'd30737, 16'd14630, 16'd54468, 16'd56033, 16'd22796, 16'd6846, 16'd20203, 16'd61907, 16'd56759, 16'd53305, 16'd62157});
	test_expansion(128'h36cfaafc1c46e5caf2037da1700607d2, {16'd30265, 16'd47728, 16'd52124, 16'd43458, 16'd38853, 16'd65098, 16'd2430, 16'd14120, 16'd36085, 16'd63972, 16'd11035, 16'd18352, 16'd21684, 16'd24072, 16'd12741, 16'd694, 16'd62328, 16'd56843, 16'd58706, 16'd37149, 16'd15684, 16'd28606, 16'd43165, 16'd29482, 16'd42239, 16'd33737});
	test_expansion(128'h05880d799d929121efdeff8b0f305ed4, {16'd31276, 16'd10309, 16'd3298, 16'd1338, 16'd5188, 16'd40793, 16'd22013, 16'd1929, 16'd10555, 16'd38605, 16'd8606, 16'd16801, 16'd52308, 16'd55827, 16'd61483, 16'd15120, 16'd44901, 16'd13076, 16'd13551, 16'd23227, 16'd51221, 16'd39076, 16'd2476, 16'd12468, 16'd30118, 16'd63390});
	test_expansion(128'h7fe222345e8fa7f3098e56a82e84f052, {16'd17787, 16'd42013, 16'd12349, 16'd5227, 16'd64891, 16'd2243, 16'd63967, 16'd49026, 16'd29988, 16'd1837, 16'd60165, 16'd26620, 16'd15892, 16'd48397, 16'd28744, 16'd9642, 16'd24653, 16'd13716, 16'd25872, 16'd6344, 16'd12135, 16'd24721, 16'd42969, 16'd1261, 16'd206, 16'd47897});
	test_expansion(128'h98bf320f3153239e8543336f6bc81d46, {16'd56228, 16'd14564, 16'd63943, 16'd48733, 16'd41495, 16'd45022, 16'd355, 16'd3486, 16'd42835, 16'd38656, 16'd62997, 16'd45229, 16'd47776, 16'd32654, 16'd59829, 16'd61519, 16'd48634, 16'd6867, 16'd40611, 16'd171, 16'd52771, 16'd5079, 16'd34336, 16'd18435, 16'd11895, 16'd26786});
	test_expansion(128'h5556a02b86c60f7851eca5605abbf6a6, {16'd11054, 16'd61050, 16'd64728, 16'd21701, 16'd37500, 16'd24350, 16'd27224, 16'd10795, 16'd28165, 16'd25652, 16'd42774, 16'd44103, 16'd59236, 16'd34711, 16'd63746, 16'd46534, 16'd65346, 16'd59528, 16'd2797, 16'd38268, 16'd60588, 16'd49447, 16'd41276, 16'd19649, 16'd63394, 16'd32580});
	test_expansion(128'h6282b8b91ecda4cb3fcad477d7839f79, {16'd5276, 16'd6697, 16'd3666, 16'd28578, 16'd59004, 16'd26510, 16'd16588, 16'd28094, 16'd52845, 16'd50556, 16'd46974, 16'd6194, 16'd57771, 16'd3855, 16'd16667, 16'd423, 16'd16228, 16'd64540, 16'd53386, 16'd9482, 16'd48026, 16'd52343, 16'd61129, 16'd1525, 16'd3856, 16'd62882});
	test_expansion(128'h203834e71bc1965dc92e728533f69c99, {16'd32013, 16'd40849, 16'd43353, 16'd3156, 16'd26471, 16'd2161, 16'd19699, 16'd60524, 16'd43143, 16'd3891, 16'd50979, 16'd37360, 16'd61559, 16'd41729, 16'd50785, 16'd27918, 16'd56137, 16'd16909, 16'd19413, 16'd23351, 16'd56263, 16'd17527, 16'd23976, 16'd9708, 16'd28396, 16'd20599});
	test_expansion(128'hcdc28a2a466e5c71e313fb1c6377e0a7, {16'd55436, 16'd5080, 16'd50068, 16'd59950, 16'd6644, 16'd62944, 16'd18017, 16'd46533, 16'd34952, 16'd6817, 16'd38310, 16'd36163, 16'd18489, 16'd29208, 16'd29658, 16'd41087, 16'd45489, 16'd39715, 16'd19489, 16'd31775, 16'd34295, 16'd29249, 16'd12907, 16'd35468, 16'd7685, 16'd56100});
	test_expansion(128'h55650e5f6eb63d69c28212aabdbf6fbc, {16'd26126, 16'd41720, 16'd36411, 16'd4899, 16'd15088, 16'd12940, 16'd58742, 16'd14612, 16'd59252, 16'd4224, 16'd30996, 16'd27268, 16'd32248, 16'd4778, 16'd12142, 16'd11650, 16'd37235, 16'd8036, 16'd64648, 16'd28007, 16'd12780, 16'd8066, 16'd20772, 16'd35474, 16'd26476, 16'd3972});
	test_expansion(128'hc969773ac63779730d3fa4277c926607, {16'd1529, 16'd43705, 16'd64748, 16'd47576, 16'd22022, 16'd47606, 16'd44340, 16'd537, 16'd6426, 16'd33648, 16'd40166, 16'd2456, 16'd37408, 16'd64074, 16'd10496, 16'd22415, 16'd26733, 16'd24473, 16'd35858, 16'd44720, 16'd8669, 16'd55394, 16'd61250, 16'd3945, 16'd27675, 16'd32467});
	test_expansion(128'hf1455b5787692c10b0827de0d34cb19f, {16'd34625, 16'd31386, 16'd8124, 16'd3897, 16'd23705, 16'd38056, 16'd37435, 16'd35819, 16'd10402, 16'd1921, 16'd30102, 16'd64798, 16'd25432, 16'd34964, 16'd19760, 16'd50501, 16'd52657, 16'd64671, 16'd29476, 16'd3914, 16'd48184, 16'd5832, 16'd36152, 16'd29777, 16'd39471, 16'd8063});
	test_expansion(128'h1d411d2ba24fecfde501d332c646175b, {16'd33567, 16'd4258, 16'd48403, 16'd9204, 16'd41589, 16'd50909, 16'd56762, 16'd40320, 16'd11088, 16'd51499, 16'd28146, 16'd3094, 16'd7021, 16'd29159, 16'd48748, 16'd27748, 16'd7453, 16'd15448, 16'd25462, 16'd444, 16'd11424, 16'd31348, 16'd39671, 16'd22838, 16'd23349, 16'd11623});
	test_expansion(128'h27ea74637dd3048e804ba3056ef1967b, {16'd35167, 16'd56401, 16'd50582, 16'd2843, 16'd41504, 16'd40253, 16'd43232, 16'd61459, 16'd27809, 16'd49058, 16'd45025, 16'd65036, 16'd64794, 16'd28525, 16'd25996, 16'd27849, 16'd34917, 16'd41193, 16'd56646, 16'd11914, 16'd11731, 16'd37913, 16'd274, 16'd55966, 16'd50278, 16'd3239});
	test_expansion(128'h384f22bfb2757a72831c49005ede0f79, {16'd20671, 16'd29330, 16'd4386, 16'd5866, 16'd9156, 16'd64921, 16'd4478, 16'd63175, 16'd40303, 16'd59215, 16'd5480, 16'd38774, 16'd3073, 16'd10011, 16'd23725, 16'd11284, 16'd19479, 16'd30214, 16'd30213, 16'd48799, 16'd18976, 16'd63173, 16'd63014, 16'd42481, 16'd35921, 16'd62397});
	test_expansion(128'hf623fb88f55ff8924806df81ce3fc630, {16'd55132, 16'd2070, 16'd6976, 16'd57887, 16'd47814, 16'd59523, 16'd50259, 16'd62244, 16'd37660, 16'd4016, 16'd30413, 16'd26987, 16'd36971, 16'd41461, 16'd54447, 16'd25308, 16'd37738, 16'd28063, 16'd6832, 16'd59970, 16'd3586, 16'd61858, 16'd47229, 16'd38814, 16'd17685, 16'd3100});
	test_expansion(128'hbaf3a431188be99181ebcd4f6854df6d, {16'd7488, 16'd2227, 16'd40249, 16'd44613, 16'd60713, 16'd44424, 16'd34842, 16'd31328, 16'd61079, 16'd8958, 16'd24996, 16'd55658, 16'd58072, 16'd42061, 16'd16232, 16'd63854, 16'd35630, 16'd46763, 16'd41974, 16'd5994, 16'd41638, 16'd27405, 16'd5658, 16'd5124, 16'd6940, 16'd49195});
	test_expansion(128'h35bb3695f8bfa9fc70d0b3b99efd7502, {16'd6587, 16'd58415, 16'd21493, 16'd43698, 16'd29938, 16'd40232, 16'd48126, 16'd32760, 16'd34118, 16'd59430, 16'd6122, 16'd38643, 16'd44978, 16'd11451, 16'd45708, 16'd18914, 16'd50, 16'd30415, 16'd28396, 16'd4620, 16'd48339, 16'd60057, 16'd42378, 16'd291, 16'd29412, 16'd13781});
	test_expansion(128'he8b69fcca44450d1faaa02fc9e48a738, {16'd19674, 16'd829, 16'd40218, 16'd53645, 16'd8502, 16'd59609, 16'd20269, 16'd36868, 16'd5698, 16'd51542, 16'd56066, 16'd24803, 16'd5975, 16'd54328, 16'd29691, 16'd31841, 16'd30105, 16'd46785, 16'd32580, 16'd17537, 16'd62182, 16'd37567, 16'd18240, 16'd53830, 16'd47535, 16'd43500});
	test_expansion(128'hf9d5bda466f8dc4e38cd07020c3d48e1, {16'd15601, 16'd36283, 16'd47983, 16'd56138, 16'd59900, 16'd49705, 16'd62525, 16'd2502, 16'd20730, 16'd35277, 16'd44239, 16'd10158, 16'd1610, 16'd34678, 16'd56259, 16'd35544, 16'd3396, 16'd29330, 16'd34813, 16'd18928, 16'd13939, 16'd48782, 16'd23745, 16'd7366, 16'd44177, 16'd36884});
	test_expansion(128'h7ea05c833b4c7827abf325991ca99c00, {16'd18381, 16'd52078, 16'd25536, 16'd65213, 16'd28050, 16'd43374, 16'd24169, 16'd3018, 16'd7468, 16'd52172, 16'd61244, 16'd28751, 16'd60007, 16'd16550, 16'd50030, 16'd8282, 16'd28179, 16'd36916, 16'd44101, 16'd44769, 16'd64294, 16'd17990, 16'd6482, 16'd14846, 16'd31875, 16'd39907});
	test_expansion(128'ha59c43b5197865e76e15ff254c9dbe44, {16'd45773, 16'd57448, 16'd35922, 16'd48680, 16'd48061, 16'd2720, 16'd49354, 16'd62258, 16'd56954, 16'd52276, 16'd56061, 16'd62512, 16'd39996, 16'd52652, 16'd19622, 16'd55420, 16'd60676, 16'd1745, 16'd25454, 16'd25431, 16'd21748, 16'd10651, 16'd7281, 16'd43152, 16'd5054, 16'd11893});
	test_expansion(128'h5cb5d6b308872614f49e1ffa22ef00b3, {16'd33721, 16'd25283, 16'd48714, 16'd39310, 16'd13821, 16'd1674, 16'd47826, 16'd35732, 16'd7177, 16'd7133, 16'd4523, 16'd21024, 16'd5143, 16'd22315, 16'd65448, 16'd40049, 16'd26539, 16'd3727, 16'd11323, 16'd21610, 16'd40134, 16'd41421, 16'd11750, 16'd54058, 16'd4603, 16'd46305});
	test_expansion(128'h06067d9efd2053dd1eab22b0a919db55, {16'd6542, 16'd46350, 16'd49358, 16'd41395, 16'd31985, 16'd8416, 16'd64652, 16'd58595, 16'd16252, 16'd45304, 16'd20361, 16'd62693, 16'd41440, 16'd30252, 16'd52188, 16'd39288, 16'd35812, 16'd64390, 16'd59861, 16'd12370, 16'd57411, 16'd57407, 16'd9196, 16'd33480, 16'd20392, 16'd7748});
	test_expansion(128'hd2aaa2750e008af96bd4cee240b05323, {16'd15656, 16'd15523, 16'd41191, 16'd35145, 16'd27063, 16'd60325, 16'd7823, 16'd54722, 16'd60910, 16'd12646, 16'd56834, 16'd29513, 16'd39326, 16'd33241, 16'd58866, 16'd16814, 16'd63516, 16'd23771, 16'd1387, 16'd5117, 16'd51846, 16'd25542, 16'd46530, 16'd35620, 16'd17911, 16'd23088});
	test_expansion(128'he4b42457b5b0f63738d927152c2847c0, {16'd25586, 16'd42032, 16'd15259, 16'd2286, 16'd13513, 16'd1151, 16'd32259, 16'd100, 16'd44347, 16'd58516, 16'd33293, 16'd37996, 16'd31762, 16'd57546, 16'd23108, 16'd34069, 16'd16417, 16'd14095, 16'd52147, 16'd49164, 16'd56101, 16'd46299, 16'd15482, 16'd45761, 16'd13242, 16'd61379});
	test_expansion(128'heb88ab831494265c4d0e9c2cf3de81a6, {16'd39679, 16'd41673, 16'd54205, 16'd19634, 16'd34516, 16'd59736, 16'd46116, 16'd21392, 16'd23027, 16'd57477, 16'd16955, 16'd40409, 16'd3259, 16'd54405, 16'd31585, 16'd19138, 16'd25707, 16'd38385, 16'd32847, 16'd59329, 16'd33421, 16'd8544, 16'd13138, 16'd28103, 16'd34746, 16'd13377});
	test_expansion(128'hcc230c72be90ada49c29dce1d4c64ccf, {16'd23002, 16'd54456, 16'd52527, 16'd24332, 16'd3122, 16'd46417, 16'd5527, 16'd53247, 16'd38304, 16'd37384, 16'd15767, 16'd43924, 16'd13402, 16'd58759, 16'd39300, 16'd1546, 16'd20806, 16'd21576, 16'd9639, 16'd18250, 16'd29965, 16'd62255, 16'd42341, 16'd33162, 16'd4051, 16'd56880});
	test_expansion(128'h7f4f5307f86b5a77cefed583520bc52c, {16'd38182, 16'd23417, 16'd5050, 16'd46466, 16'd43965, 16'd53664, 16'd12424, 16'd60109, 16'd24594, 16'd11519, 16'd32715, 16'd65519, 16'd59096, 16'd33620, 16'd16692, 16'd32503, 16'd27141, 16'd46809, 16'd64739, 16'd7736, 16'd33457, 16'd22306, 16'd3940, 16'd9696, 16'd52747, 16'd33729});
	test_expansion(128'h00657b9e98671bc51ce40ed52fe260b4, {16'd51620, 16'd37663, 16'd50069, 16'd54812, 16'd30045, 16'd4157, 16'd63108, 16'd45299, 16'd33367, 16'd28273, 16'd59574, 16'd48639, 16'd9483, 16'd3971, 16'd59738, 16'd53144, 16'd3189, 16'd33321, 16'd39669, 16'd33716, 16'd35738, 16'd18985, 16'd8826, 16'd41919, 16'd42443, 16'd37786});
	test_expansion(128'hd5791f2b86bbbf276668e9f6463262bb, {16'd12641, 16'd42978, 16'd24239, 16'd61768, 16'd33253, 16'd46708, 16'd54823, 16'd39650, 16'd37893, 16'd46915, 16'd10140, 16'd32774, 16'd37937, 16'd11253, 16'd50143, 16'd28517, 16'd49217, 16'd47670, 16'd35404, 16'd58200, 16'd16638, 16'd1542, 16'd2611, 16'd8712, 16'd58440, 16'd10831});
	test_expansion(128'h61d7e24420f4c7c4acc23b8f1696ed48, {16'd19822, 16'd57636, 16'd10362, 16'd31551, 16'd36035, 16'd34173, 16'd24982, 16'd55668, 16'd56490, 16'd40404, 16'd6107, 16'd57927, 16'd19108, 16'd29629, 16'd38928, 16'd26708, 16'd41491, 16'd55521, 16'd32551, 16'd15115, 16'd29714, 16'd62817, 16'd44177, 16'd42149, 16'd50400, 16'd34820});
	test_expansion(128'h65365392b11277ed98497a593113da07, {16'd4153, 16'd64358, 16'd19021, 16'd7273, 16'd32229, 16'd46491, 16'd12848, 16'd2699, 16'd21178, 16'd10734, 16'd41007, 16'd16868, 16'd3194, 16'd21064, 16'd51740, 16'd10198, 16'd44570, 16'd13992, 16'd58901, 16'd60956, 16'd9275, 16'd19183, 16'd20491, 16'd11360, 16'd64861, 16'd39643});
	test_expansion(128'h115beedaf073c36d094d47943ffd0cc7, {16'd5505, 16'd27290, 16'd60810, 16'd28275, 16'd21058, 16'd14311, 16'd16502, 16'd1887, 16'd16380, 16'd49770, 16'd64768, 16'd28796, 16'd13099, 16'd37043, 16'd4334, 16'd46665, 16'd25724, 16'd11511, 16'd48930, 16'd10033, 16'd62972, 16'd45277, 16'd9065, 16'd49480, 16'd64808, 16'd22762});
	test_expansion(128'hec0ed6756c4c1fa89ef9981b2b5db817, {16'd31717, 16'd46410, 16'd10667, 16'd6524, 16'd50607, 16'd4336, 16'd58891, 16'd18882, 16'd35009, 16'd2158, 16'd61863, 16'd14407, 16'd47479, 16'd16478, 16'd40224, 16'd46518, 16'd18943, 16'd30705, 16'd22209, 16'd27193, 16'd47218, 16'd11468, 16'd56242, 16'd31603, 16'd21109, 16'd39491});
	test_expansion(128'hc2e341760d88ea580fbddc5f0b161e95, {16'd39522, 16'd6024, 16'd47271, 16'd37195, 16'd44348, 16'd56178, 16'd17165, 16'd51000, 16'd43906, 16'd46567, 16'd26597, 16'd51577, 16'd40102, 16'd20389, 16'd3997, 16'd3129, 16'd50909, 16'd20345, 16'd18027, 16'd19989, 16'd50227, 16'd23192, 16'd58740, 16'd18561, 16'd20649, 16'd23898});
	test_expansion(128'hf484cd98490b98534e3aeafa78fec44d, {16'd41388, 16'd15429, 16'd61792, 16'd13880, 16'd32683, 16'd51124, 16'd57579, 16'd39603, 16'd820, 16'd13573, 16'd41865, 16'd55353, 16'd63205, 16'd57507, 16'd8343, 16'd45275, 16'd23893, 16'd48957, 16'd21961, 16'd52611, 16'd60107, 16'd36753, 16'd26475, 16'd51231, 16'd28594, 16'd36357});
	test_expansion(128'he6961dcc95bba1da7343f57f3a05272e, {16'd9787, 16'd53605, 16'd39954, 16'd62268, 16'd40948, 16'd8391, 16'd7791, 16'd48022, 16'd5316, 16'd17866, 16'd34135, 16'd64598, 16'd33564, 16'd42825, 16'd63876, 16'd54602, 16'd4837, 16'd13136, 16'd53458, 16'd13971, 16'd12186, 16'd55058, 16'd22448, 16'd42295, 16'd58925, 16'd60925});
	test_expansion(128'h4991316ae7ea5bbefc32706c1a660436, {16'd36960, 16'd13825, 16'd17742, 16'd20953, 16'd15365, 16'd13079, 16'd61577, 16'd10892, 16'd53205, 16'd34595, 16'd17903, 16'd19135, 16'd56610, 16'd9158, 16'd34786, 16'd8196, 16'd44194, 16'd12214, 16'd23355, 16'd39454, 16'd22331, 16'd26334, 16'd37637, 16'd37224, 16'd51555, 16'd57932});
	test_expansion(128'h28765aff47e289d3f7000f58786c5a8b, {16'd2561, 16'd61000, 16'd30375, 16'd50730, 16'd18862, 16'd10758, 16'd53313, 16'd22281, 16'd33999, 16'd44756, 16'd38672, 16'd26280, 16'd15676, 16'd35153, 16'd3741, 16'd2568, 16'd3658, 16'd9145, 16'd38051, 16'd11780, 16'd62611, 16'd12251, 16'd16608, 16'd26131, 16'd3029, 16'd680});
	test_expansion(128'hb41bedfc260080bbe7d646125b6f717b, {16'd6255, 16'd19269, 16'd39315, 16'd33214, 16'd6970, 16'd58194, 16'd14639, 16'd48773, 16'd5489, 16'd16557, 16'd35077, 16'd31070, 16'd57716, 16'd39517, 16'd28597, 16'd58518, 16'd64493, 16'd45474, 16'd61310, 16'd34047, 16'd16292, 16'd37014, 16'd54366, 16'd39096, 16'd54798, 16'd13812});
	test_expansion(128'hbee8cf2034a65fb84f08a2feba83dd70, {16'd37879, 16'd37477, 16'd61281, 16'd22851, 16'd15607, 16'd3244, 16'd41461, 16'd27533, 16'd46957, 16'd11596, 16'd16566, 16'd36534, 16'd11652, 16'd55472, 16'd40288, 16'd8255, 16'd24284, 16'd50199, 16'd48353, 16'd2059, 16'd18867, 16'd56924, 16'd4037, 16'd10357, 16'd52617, 16'd52766});
	test_expansion(128'h38a1247af73c66f94f6aa7efa709c529, {16'd59230, 16'd45031, 16'd55022, 16'd41539, 16'd30192, 16'd43358, 16'd61086, 16'd10474, 16'd31464, 16'd56230, 16'd26245, 16'd33089, 16'd59054, 16'd48713, 16'd11577, 16'd44810, 16'd34339, 16'd15496, 16'd1143, 16'd9555, 16'd5747, 16'd2474, 16'd10745, 16'd16757, 16'd62646, 16'd33661});
	test_expansion(128'h19a8e303044e1ca3c348b2867d63c377, {16'd51605, 16'd10308, 16'd4976, 16'd24724, 16'd191, 16'd5316, 16'd21840, 16'd26794, 16'd15341, 16'd29152, 16'd44321, 16'd3429, 16'd47978, 16'd19095, 16'd43132, 16'd26532, 16'd37883, 16'd27772, 16'd42246, 16'd48568, 16'd26267, 16'd30129, 16'd64430, 16'd43522, 16'd28573, 16'd47139});
	test_expansion(128'he0ded111badf1958812137b9b3878106, {16'd19933, 16'd32517, 16'd43947, 16'd39684, 16'd47711, 16'd24823, 16'd54748, 16'd56545, 16'd62125, 16'd43335, 16'd50578, 16'd12326, 16'd46059, 16'd37418, 16'd60648, 16'd20971, 16'd36810, 16'd40331, 16'd57604, 16'd57435, 16'd39560, 16'd47855, 16'd39513, 16'd41551, 16'd9583, 16'd32994});
	test_expansion(128'h354910dbc324afa756f038872257a928, {16'd47534, 16'd31370, 16'd14803, 16'd51513, 16'd41428, 16'd53742, 16'd21562, 16'd18750, 16'd54350, 16'd32552, 16'd1195, 16'd15513, 16'd22323, 16'd25100, 16'd30144, 16'd3172, 16'd19389, 16'd30378, 16'd30466, 16'd1663, 16'd54266, 16'd12751, 16'd42693, 16'd27019, 16'd57059, 16'd59941});
	test_expansion(128'hf1684a00c2075a99f34af542832b6331, {16'd10869, 16'd57557, 16'd45400, 16'd8444, 16'd35163, 16'd24160, 16'd41005, 16'd14075, 16'd51308, 16'd20427, 16'd23716, 16'd7589, 16'd49612, 16'd43075, 16'd22902, 16'd52090, 16'd44782, 16'd947, 16'd14521, 16'd45700, 16'd12846, 16'd45846, 16'd64698, 16'd16674, 16'd28507, 16'd1140});
	test_expansion(128'h6fba792a9ed1f900fff4401a1dd8e632, {16'd54775, 16'd30127, 16'd23883, 16'd55719, 16'd2836, 16'd30109, 16'd17907, 16'd31236, 16'd54635, 16'd60627, 16'd29495, 16'd48346, 16'd17757, 16'd64022, 16'd59574, 16'd29183, 16'd7044, 16'd54686, 16'd9017, 16'd43416, 16'd61026, 16'd22746, 16'd10103, 16'd56560, 16'd8674, 16'd50562});
	test_expansion(128'hce65e1a43b92535c452ffb95e76a912e, {16'd42436, 16'd23431, 16'd42577, 16'd24155, 16'd44443, 16'd37687, 16'd59640, 16'd31125, 16'd54447, 16'd18537, 16'd35069, 16'd37937, 16'd873, 16'd3109, 16'd42551, 16'd45670, 16'd7939, 16'd22690, 16'd24151, 16'd14724, 16'd7689, 16'd54166, 16'd10081, 16'd4755, 16'd38123, 16'd8754});
	test_expansion(128'he21c730f156ccc8ce187ad50cf7a3543, {16'd55916, 16'd21705, 16'd34788, 16'd2991, 16'd21705, 16'd61222, 16'd58799, 16'd8993, 16'd21701, 16'd38856, 16'd17867, 16'd40616, 16'd50404, 16'd48553, 16'd19448, 16'd39687, 16'd27662, 16'd26413, 16'd19615, 16'd32819, 16'd9958, 16'd63934, 16'd26839, 16'd24020, 16'd32355, 16'd2148});
	test_expansion(128'he2ad4e0bfe6e501427325b2e30153c0f, {16'd6633, 16'd18655, 16'd45857, 16'd61995, 16'd51476, 16'd51178, 16'd26641, 16'd7724, 16'd30871, 16'd20047, 16'd32432, 16'd21647, 16'd8695, 16'd11894, 16'd64125, 16'd7472, 16'd35929, 16'd57565, 16'd20581, 16'd48111, 16'd29377, 16'd61354, 16'd31883, 16'd63733, 16'd25769, 16'd23066});
	test_expansion(128'hb2415199ff4f5a29ad9ff7d552774b55, {16'd45743, 16'd58520, 16'd29861, 16'd23844, 16'd44975, 16'd37904, 16'd709, 16'd61723, 16'd41509, 16'd10008, 16'd14742, 16'd18247, 16'd33503, 16'd17703, 16'd6873, 16'd4909, 16'd4538, 16'd40729, 16'd18934, 16'd58080, 16'd11011, 16'd57366, 16'd14031, 16'd14065, 16'd27475, 16'd34632});
	test_expansion(128'hf97c0755542c6c3aa3d2f9874675f411, {16'd7474, 16'd22865, 16'd19042, 16'd23948, 16'd40231, 16'd55346, 16'd31174, 16'd59034, 16'd64371, 16'd19210, 16'd45272, 16'd47609, 16'd23737, 16'd22610, 16'd37897, 16'd32289, 16'd56624, 16'd18317, 16'd26258, 16'd33931, 16'd53644, 16'd17363, 16'd26422, 16'd51423, 16'd30831, 16'd4032});
	test_expansion(128'h0f8af04f61fa6c0083e1a63a7ac5fae0, {16'd25910, 16'd43612, 16'd1156, 16'd5408, 16'd12680, 16'd49629, 16'd55387, 16'd35356, 16'd64468, 16'd24411, 16'd41958, 16'd19017, 16'd58432, 16'd5698, 16'd25557, 16'd63915, 16'd36689, 16'd18804, 16'd44930, 16'd23528, 16'd45302, 16'd63073, 16'd8885, 16'd37446, 16'd27530, 16'd33732});
	test_expansion(128'h7c757f6e5bd6590ad42f3852ba6e84ad, {16'd53602, 16'd2490, 16'd12567, 16'd40418, 16'd3124, 16'd51224, 16'd27947, 16'd15188, 16'd38007, 16'd57504, 16'd25242, 16'd56534, 16'd23655, 16'd4596, 16'd21126, 16'd48356, 16'd58048, 16'd51844, 16'd545, 16'd33286, 16'd51117, 16'd2888, 16'd16704, 16'd40330, 16'd13230, 16'd20294});
	test_expansion(128'hdd26141280f5694a6f1a163457b7860a, {16'd50555, 16'd41708, 16'd63489, 16'd4411, 16'd10788, 16'd9630, 16'd18151, 16'd63549, 16'd6798, 16'd59527, 16'd19532, 16'd2232, 16'd53135, 16'd13201, 16'd21241, 16'd22306, 16'd58537, 16'd14826, 16'd41958, 16'd5955, 16'd18681, 16'd43357, 16'd36729, 16'd54615, 16'd47762, 16'd36114});
	test_expansion(128'ha3372bc589bf3599e368201270de67ae, {16'd53083, 16'd19257, 16'd50120, 16'd57251, 16'd12980, 16'd52842, 16'd28785, 16'd7865, 16'd45443, 16'd23489, 16'd65333, 16'd51760, 16'd56114, 16'd54999, 16'd22514, 16'd47274, 16'd18191, 16'd15378, 16'd38291, 16'd63343, 16'd21433, 16'd34863, 16'd27530, 16'd19019, 16'd27833, 16'd24407});
	test_expansion(128'h19a3d293608ce270294aed298ea278f4, {16'd43725, 16'd18986, 16'd27352, 16'd45755, 16'd41740, 16'd25379, 16'd62667, 16'd20443, 16'd437, 16'd25037, 16'd39768, 16'd52339, 16'd38032, 16'd34835, 16'd28467, 16'd46926, 16'd31113, 16'd11468, 16'd33461, 16'd17867, 16'd62995, 16'd51411, 16'd15793, 16'd22482, 16'd61373, 16'd49419});
	test_expansion(128'h05c8465a50f97e7e058730393bae561a, {16'd37201, 16'd36414, 16'd32495, 16'd14298, 16'd28183, 16'd6207, 16'd41144, 16'd25883, 16'd32040, 16'd15844, 16'd20630, 16'd51489, 16'd20807, 16'd7531, 16'd63279, 16'd26429, 16'd39667, 16'd1566, 16'd48404, 16'd48839, 16'd14400, 16'd28732, 16'd4204, 16'd53514, 16'd64570, 16'd12727});
	test_expansion(128'hd3b50dc1eb71073c00f899773ed7849b, {16'd50263, 16'd38521, 16'd34830, 16'd61354, 16'd28497, 16'd19393, 16'd11911, 16'd37080, 16'd34416, 16'd7406, 16'd52273, 16'd22760, 16'd50622, 16'd44153, 16'd56176, 16'd4530, 16'd61163, 16'd33098, 16'd55508, 16'd24412, 16'd24450, 16'd54093, 16'd2507, 16'd25896, 16'd17945, 16'd19381});
	test_expansion(128'hbae318ab394b65aef859cec265c0da45, {16'd55307, 16'd43758, 16'd28397, 16'd62839, 16'd14271, 16'd7268, 16'd36182, 16'd38296, 16'd21508, 16'd40204, 16'd45546, 16'd4401, 16'd41877, 16'd62896, 16'd5692, 16'd29975, 16'd29348, 16'd12949, 16'd173, 16'd13640, 16'd49586, 16'd3013, 16'd56330, 16'd8008, 16'd6684, 16'd10887});
	test_expansion(128'hebcf1bb6ff285f8c3aa77fbeb6fa482b, {16'd44761, 16'd60958, 16'd61718, 16'd31467, 16'd25491, 16'd60202, 16'd44635, 16'd39586, 16'd59338, 16'd31957, 16'd44190, 16'd18369, 16'd41105, 16'd2664, 16'd20958, 16'd3404, 16'd51690, 16'd36844, 16'd18570, 16'd2682, 16'd26643, 16'd55503, 16'd29929, 16'd56626, 16'd3985, 16'd27557});
	test_expansion(128'h63be8182ee2d77f878f390176c682947, {16'd6697, 16'd32129, 16'd32761, 16'd48259, 16'd61729, 16'd36387, 16'd22178, 16'd8722, 16'd6778, 16'd37330, 16'd44498, 16'd57899, 16'd59619, 16'd42366, 16'd4827, 16'd9198, 16'd29979, 16'd30017, 16'd5904, 16'd13422, 16'd27513, 16'd2693, 16'd7525, 16'd17017, 16'd29874, 16'd61253});
	test_expansion(128'h4781b6f19dc3a727db1e0dfa22c033c4, {16'd3284, 16'd59837, 16'd16569, 16'd14019, 16'd14210, 16'd49798, 16'd51768, 16'd9536, 16'd56476, 16'd20483, 16'd55943, 16'd49678, 16'd1943, 16'd39948, 16'd21290, 16'd50225, 16'd34775, 16'd5461, 16'd44405, 16'd60314, 16'd65068, 16'd36405, 16'd39270, 16'd53547, 16'd50528, 16'd59952});
	test_expansion(128'h665c8818fbec46c4bcb5297e701b7fb0, {16'd10772, 16'd13699, 16'd24877, 16'd21762, 16'd23127, 16'd614, 16'd20470, 16'd9645, 16'd55696, 16'd32688, 16'd34928, 16'd14012, 16'd35205, 16'd21378, 16'd16439, 16'd29766, 16'd23389, 16'd21596, 16'd23509, 16'd8156, 16'd22730, 16'd51326, 16'd31355, 16'd58333, 16'd25665, 16'd4428});
	test_expansion(128'h9b98136ece72947cc832f7a2eb584900, {16'd14446, 16'd5078, 16'd19304, 16'd25436, 16'd43559, 16'd41055, 16'd30176, 16'd5966, 16'd53237, 16'd59888, 16'd3963, 16'd48495, 16'd2684, 16'd40652, 16'd23117, 16'd50947, 16'd18168, 16'd29628, 16'd60417, 16'd35782, 16'd59738, 16'd17324, 16'd19898, 16'd8160, 16'd50914, 16'd30123});
	test_expansion(128'h2fde358ef1b5cef81f619f6fd0c31297, {16'd4932, 16'd53061, 16'd42372, 16'd12028, 16'd22215, 16'd61495, 16'd60117, 16'd47941, 16'd36499, 16'd60303, 16'd39239, 16'd47244, 16'd57773, 16'd49717, 16'd18784, 16'd7464, 16'd35954, 16'd16496, 16'd9267, 16'd27675, 16'd51680, 16'd42650, 16'd12232, 16'd22318, 16'd2650, 16'd11201});
	test_expansion(128'h623b3bc96b9a3560c26ec2db48b18926, {16'd13502, 16'd53790, 16'd52887, 16'd8822, 16'd1029, 16'd42887, 16'd50159, 16'd46113, 16'd57936, 16'd50692, 16'd6858, 16'd34245, 16'd21316, 16'd55017, 16'd62487, 16'd61278, 16'd28562, 16'd62103, 16'd27692, 16'd48960, 16'd52439, 16'd12727, 16'd22475, 16'd39191, 16'd6079, 16'd55568});
	test_expansion(128'h33656fd1ac037201e2690641f8d0ba6b, {16'd3899, 16'd57292, 16'd24034, 16'd15451, 16'd32918, 16'd12844, 16'd63386, 16'd19045, 16'd58749, 16'd60192, 16'd58974, 16'd2552, 16'd16099, 16'd16091, 16'd36021, 16'd56697, 16'd25260, 16'd14590, 16'd2277, 16'd50778, 16'd10202, 16'd65331, 16'd11848, 16'd58163, 16'd23506, 16'd62777});
	test_expansion(128'he9aaee9076b4325efae45e312fa22203, {16'd57593, 16'd45130, 16'd24215, 16'd42092, 16'd30201, 16'd59654, 16'd1222, 16'd29957, 16'd63294, 16'd45612, 16'd53220, 16'd17321, 16'd63573, 16'd28418, 16'd24733, 16'd42652, 16'd20837, 16'd42561, 16'd52332, 16'd12428, 16'd14443, 16'd46238, 16'd13212, 16'd62028, 16'd24102, 16'd33858});
	test_expansion(128'hdad491f3d44b619dc9653be2d9537709, {16'd25772, 16'd8090, 16'd36629, 16'd49147, 16'd8955, 16'd65532, 16'd23746, 16'd13171, 16'd52669, 16'd41413, 16'd61570, 16'd51453, 16'd27336, 16'd9036, 16'd42786, 16'd41750, 16'd43845, 16'd18576, 16'd49874, 16'd18538, 16'd14815, 16'd58615, 16'd12549, 16'd7047, 16'd18413, 16'd23604});
	test_expansion(128'hac750cba70c853585297df04a6c8f342, {16'd22533, 16'd14170, 16'd38920, 16'd45256, 16'd34033, 16'd34356, 16'd54922, 16'd60685, 16'd59619, 16'd12589, 16'd7924, 16'd29472, 16'd13127, 16'd29222, 16'd13484, 16'd52703, 16'd13901, 16'd44676, 16'd38432, 16'd13046, 16'd34630, 16'd16962, 16'd544, 16'd9301, 16'd49787, 16'd4935});
	test_expansion(128'hddc806faae18105a185bad7f882a8d2d, {16'd4203, 16'd28845, 16'd56632, 16'd33760, 16'd2949, 16'd15574, 16'd54524, 16'd42850, 16'd10769, 16'd44302, 16'd23698, 16'd14887, 16'd2211, 16'd26862, 16'd30169, 16'd208, 16'd21305, 16'd62043, 16'd2365, 16'd23334, 16'd30182, 16'd45750, 16'd4884, 16'd62194, 16'd13729, 16'd1015});
	test_expansion(128'h472319398972e44898642fdc673e5668, {16'd44320, 16'd24753, 16'd64823, 16'd51549, 16'd14374, 16'd47487, 16'd726, 16'd31867, 16'd61133, 16'd14173, 16'd47200, 16'd4887, 16'd30327, 16'd29122, 16'd55562, 16'd4863, 16'd35305, 16'd9693, 16'd7086, 16'd64724, 16'd40597, 16'd61597, 16'd5787, 16'd7932, 16'd65389, 16'd31683});
	test_expansion(128'h920088086190e8286a26d6f6e552ce6c, {16'd52417, 16'd9745, 16'd46920, 16'd61169, 16'd38999, 16'd49603, 16'd3750, 16'd21743, 16'd61212, 16'd21992, 16'd17977, 16'd43305, 16'd3380, 16'd4019, 16'd58679, 16'd20392, 16'd25011, 16'd25338, 16'd1660, 16'd59427, 16'd49237, 16'd55429, 16'd5744, 16'd36960, 16'd37153, 16'd1884});
	test_expansion(128'h977fab6a5b48339e6a860283163ff5d5, {16'd40966, 16'd9253, 16'd4601, 16'd29791, 16'd54739, 16'd51126, 16'd28297, 16'd16174, 16'd50501, 16'd56502, 16'd44308, 16'd58763, 16'd4571, 16'd25876, 16'd48519, 16'd59582, 16'd23578, 16'd9638, 16'd53121, 16'd63202, 16'd27704, 16'd43152, 16'd63290, 16'd7710, 16'd54040, 16'd6306});
	test_expansion(128'hf9ae0be58564b2103d69a93f8ad5e46e, {16'd5363, 16'd37431, 16'd57462, 16'd35800, 16'd54501, 16'd2332, 16'd58907, 16'd29801, 16'd28344, 16'd8420, 16'd61645, 16'd48429, 16'd49109, 16'd7525, 16'd60481, 16'd53517, 16'd15671, 16'd30091, 16'd9944, 16'd50703, 16'd17950, 16'd65021, 16'd17307, 16'd53533, 16'd60462, 16'd24897});
	test_expansion(128'h54a10091d80a8a058ed63f19bd09eaf1, {16'd20862, 16'd56322, 16'd15446, 16'd47983, 16'd61814, 16'd57925, 16'd40138, 16'd20295, 16'd31627, 16'd50838, 16'd11041, 16'd7329, 16'd33578, 16'd55468, 16'd1431, 16'd63554, 16'd28144, 16'd20430, 16'd39112, 16'd25082, 16'd5376, 16'd65081, 16'd20259, 16'd61966, 16'd49686, 16'd3069});
	test_expansion(128'hd53fbb815af31e7429ff51652a4ff58c, {16'd32119, 16'd56025, 16'd23560, 16'd51183, 16'd49455, 16'd56317, 16'd63268, 16'd10568, 16'd20655, 16'd28780, 16'd60438, 16'd2716, 16'd14002, 16'd29499, 16'd9836, 16'd33728, 16'd4126, 16'd45408, 16'd22125, 16'd61173, 16'd40966, 16'd52110, 16'd58179, 16'd3503, 16'd33642, 16'd7362});
	test_expansion(128'ha47480bb993f4caeac0dcfb5b95f766c, {16'd17580, 16'd16836, 16'd30407, 16'd52697, 16'd14699, 16'd5634, 16'd16365, 16'd31287, 16'd21461, 16'd37034, 16'd25886, 16'd43002, 16'd8557, 16'd55760, 16'd5353, 16'd20150, 16'd30279, 16'd12240, 16'd23940, 16'd30777, 16'd26436, 16'd17047, 16'd15597, 16'd55992, 16'd33940, 16'd52606});
	test_expansion(128'h1f075b3c774e39654a6468b9ab65a0e7, {16'd65499, 16'd54433, 16'd57444, 16'd54807, 16'd59970, 16'd25257, 16'd1813, 16'd55875, 16'd41255, 16'd41944, 16'd8893, 16'd38120, 16'd33340, 16'd18937, 16'd63752, 16'd26225, 16'd8856, 16'd44931, 16'd39403, 16'd37627, 16'd6369, 16'd61035, 16'd37265, 16'd44392, 16'd35443, 16'd24282});
	test_expansion(128'h2e57a27b19a5ed877420c6c308f1ce33, {16'd29664, 16'd63506, 16'd41553, 16'd19668, 16'd6134, 16'd25974, 16'd30717, 16'd37580, 16'd51030, 16'd18213, 16'd27181, 16'd6656, 16'd17259, 16'd44314, 16'd1520, 16'd54985, 16'd6164, 16'd61554, 16'd48131, 16'd15999, 16'd12983, 16'd12564, 16'd63749, 16'd44185, 16'd24334, 16'd581});
	test_expansion(128'h960ea5d0939c8789732b595f1c3fb199, {16'd37480, 16'd63636, 16'd15734, 16'd27549, 16'd3872, 16'd16139, 16'd59978, 16'd11198, 16'd16256, 16'd51975, 16'd19468, 16'd31380, 16'd55821, 16'd26462, 16'd50672, 16'd29916, 16'd50349, 16'd24202, 16'd39149, 16'd22242, 16'd40336, 16'd43817, 16'd48575, 16'd57400, 16'd9801, 16'd23762});
	test_expansion(128'haf3ba0f0283313edab3382c779975d68, {16'd61381, 16'd32650, 16'd58890, 16'd41257, 16'd34143, 16'd53999, 16'd22749, 16'd57404, 16'd13487, 16'd19557, 16'd51761, 16'd55728, 16'd44205, 16'd47237, 16'd41414, 16'd50087, 16'd20424, 16'd49555, 16'd30410, 16'd64462, 16'd42264, 16'd47362, 16'd44839, 16'd58940, 16'd1936, 16'd30157});
	test_expansion(128'ha8ab48f80595fa70e71c993c19f6ec1e, {16'd3896, 16'd17965, 16'd7262, 16'd33308, 16'd27534, 16'd58221, 16'd39947, 16'd17314, 16'd47990, 16'd52349, 16'd30744, 16'd16879, 16'd52373, 16'd50090, 16'd51379, 16'd14979, 16'd7601, 16'd32005, 16'd1453, 16'd7986, 16'd26830, 16'd36059, 16'd12795, 16'd45816, 16'd4078, 16'd53181});
	test_expansion(128'hc9a8c5314a8a9a58525ec1d9c012e612, {16'd463, 16'd4694, 16'd57381, 16'd3001, 16'd31389, 16'd3071, 16'd39643, 16'd20206, 16'd61617, 16'd41111, 16'd4034, 16'd26508, 16'd15165, 16'd26390, 16'd65325, 16'd40566, 16'd15363, 16'd52986, 16'd63814, 16'd15021, 16'd23021, 16'd185, 16'd34699, 16'd65164, 16'd38601, 16'd33224});
	test_expansion(128'hfa697133ebd4cea215d6bcc1796528d3, {16'd39813, 16'd42091, 16'd12813, 16'd34439, 16'd18706, 16'd36526, 16'd40202, 16'd19766, 16'd2509, 16'd52045, 16'd26519, 16'd27913, 16'd31749, 16'd35190, 16'd60245, 16'd40792, 16'd51452, 16'd41543, 16'd4038, 16'd41364, 16'd58511, 16'd37733, 16'd40316, 16'd50862, 16'd49413, 16'd21518});
	test_expansion(128'h2f236dc4adf329a81b396e89746aa82f, {16'd35066, 16'd25175, 16'd58317, 16'd5808, 16'd15252, 16'd55007, 16'd9102, 16'd23280, 16'd39267, 16'd61905, 16'd12329, 16'd61104, 16'd47270, 16'd48186, 16'd26535, 16'd63112, 16'd29531, 16'd5021, 16'd37271, 16'd20786, 16'd45040, 16'd59464, 16'd34171, 16'd60458, 16'd60862, 16'd570});
	test_expansion(128'h0444e87c15d7374890abf648beaf5bcf, {16'd63951, 16'd13572, 16'd56196, 16'd32324, 16'd61967, 16'd24730, 16'd19780, 16'd24944, 16'd21493, 16'd9513, 16'd29940, 16'd63343, 16'd23169, 16'd42763, 16'd39567, 16'd30034, 16'd59681, 16'd22256, 16'd29598, 16'd2972, 16'd32640, 16'd10228, 16'd63711, 16'd39498, 16'd47782, 16'd31926});
	test_expansion(128'h0c853962fedb799199e1d753e2622f8a, {16'd63346, 16'd55469, 16'd29706, 16'd18713, 16'd10195, 16'd58692, 16'd44344, 16'd26595, 16'd4718, 16'd56659, 16'd45465, 16'd52560, 16'd32316, 16'd10802, 16'd58231, 16'd11123, 16'd7102, 16'd19965, 16'd33784, 16'd18461, 16'd8192, 16'd16098, 16'd45007, 16'd56883, 16'd23376, 16'd10658});
	test_expansion(128'h7120eda6904a0153b352f2981583a348, {16'd46464, 16'd52202, 16'd29188, 16'd26773, 16'd17640, 16'd1649, 16'd37719, 16'd24544, 16'd55244, 16'd9667, 16'd47418, 16'd42043, 16'd49080, 16'd5705, 16'd41872, 16'd27982, 16'd709, 16'd26915, 16'd52551, 16'd54497, 16'd47377, 16'd50651, 16'd36977, 16'd44084, 16'd5579, 16'd65191});
	test_expansion(128'h3645c81a12ba82af44d5ff7093642538, {16'd14751, 16'd41366, 16'd21395, 16'd7007, 16'd34700, 16'd29318, 16'd60163, 16'd6324, 16'd3807, 16'd61726, 16'd53296, 16'd5371, 16'd16598, 16'd26266, 16'd44575, 16'd14291, 16'd59773, 16'd32842, 16'd39379, 16'd3450, 16'd58829, 16'd34052, 16'd22246, 16'd38963, 16'd26457, 16'd56994});
	test_expansion(128'h500f7f6e3e95558859ca7e3195554a38, {16'd52186, 16'd7409, 16'd30617, 16'd22498, 16'd8396, 16'd41666, 16'd51053, 16'd3261, 16'd57234, 16'd9619, 16'd44113, 16'd50625, 16'd50675, 16'd15875, 16'd42387, 16'd54586, 16'd54597, 16'd61129, 16'd46926, 16'd60306, 16'd9588, 16'd61185, 16'd13567, 16'd22090, 16'd37052, 16'd41534});
	test_expansion(128'ha5b0115a2ae5623acbcd414897c5b1f2, {16'd28965, 16'd58975, 16'd33557, 16'd8290, 16'd15885, 16'd42749, 16'd14561, 16'd14099, 16'd39163, 16'd61508, 16'd44868, 16'd27341, 16'd10965, 16'd48133, 16'd13103, 16'd4220, 16'd56543, 16'd40983, 16'd8871, 16'd7394, 16'd19314, 16'd25544, 16'd53154, 16'd40921, 16'd4224, 16'd9476});
	test_expansion(128'h67ece5baf1004ca2d9c862805821940d, {16'd53856, 16'd31604, 16'd7796, 16'd10675, 16'd6719, 16'd17208, 16'd51701, 16'd3988, 16'd10590, 16'd58827, 16'd51213, 16'd52544, 16'd22739, 16'd7289, 16'd40581, 16'd56547, 16'd35856, 16'd33412, 16'd30697, 16'd32883, 16'd22144, 16'd20501, 16'd62801, 16'd17299, 16'd7420, 16'd449});
	test_expansion(128'ha5fa5eb119bd193c14404bb9ae729ca3, {16'd27826, 16'd23244, 16'd6247, 16'd34517, 16'd172, 16'd57155, 16'd43482, 16'd464, 16'd61531, 16'd56859, 16'd9436, 16'd26239, 16'd33701, 16'd36133, 16'd37913, 16'd33953, 16'd5397, 16'd36978, 16'd10479, 16'd41526, 16'd11445, 16'd11951, 16'd35735, 16'd44758, 16'd35537, 16'd50597});
	test_expansion(128'h213d97a59d49a4cb55d1162ce6c28cc2, {16'd27668, 16'd22475, 16'd33468, 16'd65040, 16'd22891, 16'd20880, 16'd1692, 16'd32336, 16'd11526, 16'd18481, 16'd53045, 16'd60100, 16'd36226, 16'd60250, 16'd61654, 16'd57268, 16'd54081, 16'd63072, 16'd51419, 16'd39491, 16'd51361, 16'd57098, 16'd22350, 16'd62683, 16'd27680, 16'd40712});
	test_expansion(128'h702cceb6ae0c50e903177cab4c6f66a5, {16'd3499, 16'd53904, 16'd49554, 16'd50143, 16'd55732, 16'd31083, 16'd22153, 16'd50364, 16'd57055, 16'd13900, 16'd4640, 16'd5751, 16'd61236, 16'd17757, 16'd46772, 16'd6195, 16'd7603, 16'd5299, 16'd9340, 16'd46453, 16'd37562, 16'd60894, 16'd13684, 16'd63222, 16'd42075, 16'd49811});
	test_expansion(128'h7bf57078cdd8474f7ef0ea29eb6b9798, {16'd64176, 16'd7295, 16'd30453, 16'd22267, 16'd13994, 16'd18503, 16'd4884, 16'd4585, 16'd23053, 16'd17294, 16'd25097, 16'd2436, 16'd29157, 16'd21847, 16'd57225, 16'd59342, 16'd43919, 16'd551, 16'd54198, 16'd19442, 16'd1816, 16'd2047, 16'd48429, 16'd10757, 16'd53835, 16'd19403});
	test_expansion(128'h7423858858a27db879c299029b44b438, {16'd49606, 16'd47559, 16'd39931, 16'd24969, 16'd6002, 16'd7229, 16'd48823, 16'd9078, 16'd39947, 16'd14254, 16'd6273, 16'd36392, 16'd47812, 16'd38955, 16'd30631, 16'd42562, 16'd59231, 16'd52516, 16'd48970, 16'd31381, 16'd54577, 16'd35101, 16'd10014, 16'd10905, 16'd61181, 16'd29534});
	test_expansion(128'h0a1ebf963264d8da1df3d6887ebe6a8b, {16'd57028, 16'd39573, 16'd23462, 16'd50454, 16'd32929, 16'd45566, 16'd2983, 16'd14956, 16'd20972, 16'd51706, 16'd3169, 16'd42015, 16'd61637, 16'd34539, 16'd61474, 16'd15024, 16'd16566, 16'd7169, 16'd29446, 16'd33356, 16'd3404, 16'd61495, 16'd21390, 16'd23280, 16'd49631, 16'd6874});
	test_expansion(128'h6a9423390abe7138e506ab61647cd94e, {16'd54822, 16'd52802, 16'd47578, 16'd17195, 16'd37943, 16'd59942, 16'd31709, 16'd6876, 16'd4387, 16'd26391, 16'd43924, 16'd33515, 16'd23181, 16'd11068, 16'd26455, 16'd22895, 16'd58154, 16'd25378, 16'd58176, 16'd25965, 16'd29452, 16'd8224, 16'd55149, 16'd41434, 16'd38107, 16'd36018});
	test_expansion(128'h29d1d54db499aa097a6d2a4c81265cdd, {16'd10191, 16'd60969, 16'd6625, 16'd52404, 16'd49687, 16'd44854, 16'd47487, 16'd63834, 16'd19901, 16'd31626, 16'd27431, 16'd33257, 16'd6806, 16'd8725, 16'd56385, 16'd14696, 16'd42379, 16'd65194, 16'd56176, 16'd24889, 16'd45146, 16'd58715, 16'd52552, 16'd24284, 16'd63309, 16'd65213});
	test_expansion(128'h952523fa108b83972024f5f4902914ae, {16'd51471, 16'd60510, 16'd34179, 16'd50064, 16'd13423, 16'd60181, 16'd3223, 16'd64246, 16'd3014, 16'd24154, 16'd15944, 16'd18264, 16'd3187, 16'd12942, 16'd24004, 16'd41226, 16'd41920, 16'd58669, 16'd22223, 16'd9364, 16'd34827, 16'd49494, 16'd34183, 16'd9917, 16'd18967, 16'd62571});
	test_expansion(128'hab7cea95c071daa37eaf5c9b251a492c, {16'd36473, 16'd56986, 16'd36447, 16'd18753, 16'd544, 16'd63979, 16'd65263, 16'd19046, 16'd4939, 16'd48051, 16'd16782, 16'd17584, 16'd38543, 16'd20139, 16'd6400, 16'd27919, 16'd53154, 16'd60462, 16'd55311, 16'd38018, 16'd28630, 16'd4177, 16'd38219, 16'd20155, 16'd20294, 16'd15419});
	test_expansion(128'h6e231c193e02752e154ac069819ccd61, {16'd48081, 16'd25187, 16'd22643, 16'd36271, 16'd14965, 16'd41204, 16'd17265, 16'd31790, 16'd8067, 16'd33381, 16'd5277, 16'd4618, 16'd10980, 16'd22496, 16'd44043, 16'd30675, 16'd21191, 16'd17293, 16'd45481, 16'd12104, 16'd31803, 16'd19220, 16'd63938, 16'd60399, 16'd722, 16'd29692});
	test_expansion(128'h4299240ae58f2f662a2116c3a8cb5ecc, {16'd59592, 16'd38197, 16'd59673, 16'd53615, 16'd38695, 16'd16082, 16'd5542, 16'd50357, 16'd42067, 16'd10398, 16'd35527, 16'd47631, 16'd4402, 16'd38491, 16'd41772, 16'd45239, 16'd24364, 16'd62776, 16'd40305, 16'd2380, 16'd36729, 16'd54138, 16'd10636, 16'd64619, 16'd49933, 16'd47694});
	test_expansion(128'hbe71efaa3245a6ccc64f04f136ecf6d0, {16'd17828, 16'd43224, 16'd20378, 16'd38567, 16'd660, 16'd12949, 16'd21155, 16'd21, 16'd1382, 16'd61624, 16'd48006, 16'd1688, 16'd41993, 16'd16606, 16'd39949, 16'd65104, 16'd24474, 16'd22267, 16'd186, 16'd14662, 16'd62132, 16'd34960, 16'd51599, 16'd18301, 16'd46579, 16'd35832});
	test_expansion(128'h2a314f232ca32292ae9b496fd22a60bd, {16'd41325, 16'd55995, 16'd31103, 16'd3203, 16'd29815, 16'd14301, 16'd28695, 16'd60258, 16'd37025, 16'd20909, 16'd13589, 16'd49523, 16'd18198, 16'd38880, 16'd18329, 16'd62662, 16'd16036, 16'd6317, 16'd37668, 16'd57230, 16'd34464, 16'd8646, 16'd39425, 16'd43935, 16'd4147, 16'd59964});
	test_expansion(128'h242ae70422fb018ffab3abd44e07dab1, {16'd301, 16'd22985, 16'd34084, 16'd2114, 16'd47878, 16'd15200, 16'd54768, 16'd13413, 16'd56412, 16'd24269, 16'd35740, 16'd50264, 16'd26787, 16'd34695, 16'd12320, 16'd62645, 16'd56866, 16'd24106, 16'd14682, 16'd47925, 16'd27672, 16'd9267, 16'd15589, 16'd43617, 16'd46148, 16'd43955});
	test_expansion(128'h89be7a06b532f223712f22504db5840a, {16'd2552, 16'd54038, 16'd3768, 16'd36391, 16'd37735, 16'd45393, 16'd55906, 16'd12535, 16'd65382, 16'd58020, 16'd29139, 16'd52748, 16'd1585, 16'd42527, 16'd20681, 16'd20159, 16'd19180, 16'd20847, 16'd38320, 16'd32261, 16'd57662, 16'd7499, 16'd43994, 16'd20540, 16'd4372, 16'd15169});
	test_expansion(128'h1d57df6f94ec525e43ea0de634f4eae8, {16'd7075, 16'd46820, 16'd32621, 16'd39007, 16'd33304, 16'd34769, 16'd63471, 16'd31555, 16'd1439, 16'd33966, 16'd21571, 16'd61672, 16'd8472, 16'd17246, 16'd16613, 16'd56213, 16'd29145, 16'd12750, 16'd52992, 16'd45119, 16'd12696, 16'd39069, 16'd63153, 16'd956, 16'd57015, 16'd49434});
	test_expansion(128'hcb78bf93f9a8dc618f82269237576f46, {16'd6067, 16'd59935, 16'd62631, 16'd59717, 16'd17883, 16'd22910, 16'd19854, 16'd44639, 16'd11899, 16'd52147, 16'd63415, 16'd10557, 16'd54510, 16'd18569, 16'd34477, 16'd35550, 16'd31843, 16'd46846, 16'd60307, 16'd846, 16'd48875, 16'd25937, 16'd10189, 16'd28923, 16'd40424, 16'd65401});
	test_expansion(128'h187b078fd6d15ff7dfb93c6d4f428b52, {16'd16106, 16'd6413, 16'd48277, 16'd52402, 16'd44926, 16'd19014, 16'd18093, 16'd21841, 16'd18601, 16'd21594, 16'd30711, 16'd61324, 16'd62349, 16'd25953, 16'd50479, 16'd27679, 16'd22607, 16'd2613, 16'd9986, 16'd55437, 16'd61457, 16'd45601, 16'd30791, 16'd51647, 16'd50790, 16'd34075});
	test_expansion(128'h23ebfc2f3eb37b8771fff01dc4f85aed, {16'd9948, 16'd13067, 16'd62259, 16'd50480, 16'd19993, 16'd22480, 16'd48026, 16'd39545, 16'd51676, 16'd57449, 16'd65070, 16'd33935, 16'd54436, 16'd35578, 16'd55994, 16'd32198, 16'd52858, 16'd48828, 16'd62057, 16'd40761, 16'd48650, 16'd5925, 16'd40181, 16'd50033, 16'd37566, 16'd58724});
	test_expansion(128'hb191cdb2889717ec51b6da8e1de09643, {16'd1781, 16'd4086, 16'd16456, 16'd29013, 16'd64428, 16'd4262, 16'd45910, 16'd497, 16'd41563, 16'd40782, 16'd44607, 16'd28302, 16'd62515, 16'd9941, 16'd32551, 16'd9990, 16'd44012, 16'd1209, 16'd47145, 16'd41147, 16'd2173, 16'd19691, 16'd47353, 16'd27189, 16'd35797, 16'd1265});
	test_expansion(128'h18358edd244781c0c8cf35494cd24012, {16'd62575, 16'd59638, 16'd11964, 16'd30121, 16'd15124, 16'd53598, 16'd27377, 16'd7919, 16'd64925, 16'd29609, 16'd2585, 16'd15830, 16'd63229, 16'd30456, 16'd7999, 16'd51653, 16'd5939, 16'd12784, 16'd30255, 16'd45119, 16'd10482, 16'd63258, 16'd61114, 16'd19485, 16'd16270, 16'd42586});
	test_expansion(128'hce0789f79501216bf7365d62efe79fb7, {16'd364, 16'd35096, 16'd64539, 16'd53360, 16'd22143, 16'd49296, 16'd53059, 16'd55227, 16'd37099, 16'd32090, 16'd24556, 16'd44911, 16'd17552, 16'd27814, 16'd11012, 16'd31319, 16'd6513, 16'd24799, 16'd38883, 16'd44369, 16'd58914, 16'd62658, 16'd54750, 16'd27455, 16'd38971, 16'd35011});
	test_expansion(128'haaf08a6d6dc1677ae61fe45b4693652c, {16'd51841, 16'd29789, 16'd58943, 16'd56067, 16'd33059, 16'd64946, 16'd26091, 16'd43076, 16'd41214, 16'd35834, 16'd23747, 16'd47683, 16'd41037, 16'd48578, 16'd13651, 16'd23190, 16'd56484, 16'd15367, 16'd2120, 16'd7002, 16'd830, 16'd49809, 16'd11592, 16'd39455, 16'd14520, 16'd24728});
	test_expansion(128'h42215542df75f317610fee49b8817229, {16'd10705, 16'd105, 16'd6080, 16'd5629, 16'd46408, 16'd58548, 16'd53679, 16'd56412, 16'd64688, 16'd20352, 16'd1252, 16'd31642, 16'd58120, 16'd53672, 16'd9857, 16'd39077, 16'd59768, 16'd15275, 16'd35711, 16'd64269, 16'd20550, 16'd48892, 16'd46357, 16'd44695, 16'd31126, 16'd63325});
	test_expansion(128'hb4d1058faa080a8f76926b44562dea99, {16'd21576, 16'd18360, 16'd62771, 16'd45565, 16'd30833, 16'd41535, 16'd42556, 16'd29139, 16'd30297, 16'd49925, 16'd25651, 16'd10084, 16'd33916, 16'd56364, 16'd57387, 16'd53880, 16'd1969, 16'd45175, 16'd29256, 16'd33649, 16'd17509, 16'd31440, 16'd30943, 16'd46436, 16'd28503, 16'd13282});
	test_expansion(128'hbc4d9a376d130961be96e403e33d79d9, {16'd12343, 16'd6175, 16'd4784, 16'd41644, 16'd18002, 16'd45087, 16'd59677, 16'd9205, 16'd42206, 16'd7212, 16'd14228, 16'd20059, 16'd15060, 16'd14697, 16'd32584, 16'd49089, 16'd27533, 16'd36942, 16'd19827, 16'd42730, 16'd6366, 16'd8938, 16'd3655, 16'd18009, 16'd41551, 16'd4956});
	test_expansion(128'h35c2b9e76010a6d7a6f6d2a3f2a82d58, {16'd63505, 16'd10184, 16'd749, 16'd11105, 16'd11658, 16'd63820, 16'd53186, 16'd307, 16'd1121, 16'd11575, 16'd60882, 16'd62914, 16'd35601, 16'd19458, 16'd63826, 16'd39317, 16'd17844, 16'd2899, 16'd55011, 16'd63287, 16'd45661, 16'd40550, 16'd39438, 16'd34145, 16'd14249, 16'd60558});
	test_expansion(128'h7babd9fa8c60d51385616be2937fc403, {16'd57257, 16'd50860, 16'd2148, 16'd10827, 16'd13054, 16'd21907, 16'd62927, 16'd51378, 16'd46693, 16'd693, 16'd39473, 16'd47075, 16'd16386, 16'd45584, 16'd50255, 16'd25135, 16'd30536, 16'd59797, 16'd62787, 16'd41118, 16'd53254, 16'd6459, 16'd29021, 16'd38057, 16'd28714, 16'd58974});
	test_expansion(128'hde0b905cbf8d405b37044045f3136ee8, {16'd32341, 16'd17041, 16'd50455, 16'd54338, 16'd50915, 16'd20906, 16'd12820, 16'd16512, 16'd25199, 16'd29988, 16'd36816, 16'd55064, 16'd17036, 16'd3779, 16'd9866, 16'd56097, 16'd38121, 16'd36316, 16'd1362, 16'd33397, 16'd58974, 16'd47332, 16'd33408, 16'd21008, 16'd35866, 16'd39979});
	test_expansion(128'hb3f3461c0817ce81b4ca5a1f05e5fa7f, {16'd33815, 16'd62011, 16'd54496, 16'd45112, 16'd54057, 16'd60320, 16'd656, 16'd496, 16'd14869, 16'd14288, 16'd53141, 16'd11053, 16'd36904, 16'd56654, 16'd36144, 16'd55130, 16'd39805, 16'd36211, 16'd52776, 16'd14553, 16'd59939, 16'd61875, 16'd55484, 16'd26580, 16'd53816, 16'd19448});
	test_expansion(128'h946dea89ae5d06bfa7f93f1e172a76fa, {16'd58889, 16'd58853, 16'd4101, 16'd61646, 16'd38067, 16'd34571, 16'd39552, 16'd43893, 16'd62664, 16'd65233, 16'd10289, 16'd61536, 16'd40372, 16'd9531, 16'd49124, 16'd49221, 16'd40172, 16'd47136, 16'd5775, 16'd50767, 16'd10780, 16'd51604, 16'd32375, 16'd56749, 16'd8723, 16'd25469});
	test_expansion(128'h1c1e3631526e9c2e5dc7d325cac06c25, {16'd5672, 16'd29771, 16'd49864, 16'd11, 16'd3399, 16'd18975, 16'd43764, 16'd40182, 16'd42265, 16'd16717, 16'd29018, 16'd23843, 16'd2903, 16'd12218, 16'd21498, 16'd40432, 16'd52769, 16'd17160, 16'd17894, 16'd30051, 16'd38476, 16'd9016, 16'd50147, 16'd56655, 16'd30317, 16'd12239});
	test_expansion(128'h679daa16b3ea57c98e66a86d49be8c04, {16'd24814, 16'd57140, 16'd24001, 16'd57647, 16'd38107, 16'd29784, 16'd28361, 16'd20062, 16'd64590, 16'd28507, 16'd24749, 16'd5398, 16'd42115, 16'd63203, 16'd37807, 16'd8538, 16'd41318, 16'd49779, 16'd64926, 16'd64576, 16'd21727, 16'd50624, 16'd57882, 16'd32478, 16'd14708, 16'd6822});
	test_expansion(128'h675e1ff87ff4c7ac153a23b601d3bf53, {16'd58143, 16'd30346, 16'd19900, 16'd14789, 16'd62570, 16'd47568, 16'd43280, 16'd349, 16'd34747, 16'd40297, 16'd21383, 16'd2858, 16'd18198, 16'd40090, 16'd44791, 16'd17123, 16'd44411, 16'd35575, 16'd31803, 16'd20427, 16'd58646, 16'd446, 16'd21913, 16'd63598, 16'd50375, 16'd55974});
	test_expansion(128'h4f676610bf85f55288118477ced196a1, {16'd28769, 16'd49013, 16'd37368, 16'd22647, 16'd32388, 16'd6319, 16'd18085, 16'd5425, 16'd60332, 16'd10476, 16'd22431, 16'd38319, 16'd15638, 16'd34012, 16'd40607, 16'd7683, 16'd15882, 16'd29291, 16'd37385, 16'd60575, 16'd60400, 16'd1822, 16'd62737, 16'd57023, 16'd55448, 16'd25840});
	test_expansion(128'h207fa9cd83af1c583803e708cde70422, {16'd11326, 16'd19256, 16'd11247, 16'd43242, 16'd52817, 16'd40171, 16'd8874, 16'd25533, 16'd13823, 16'd26086, 16'd22331, 16'd2949, 16'd60305, 16'd51508, 16'd50284, 16'd45687, 16'd19300, 16'd56888, 16'd1974, 16'd25512, 16'd39031, 16'd38036, 16'd27282, 16'd25823, 16'd24848, 16'd62453});
	test_expansion(128'h324f97c83499dcc64c63fa9c6376a508, {16'd27733, 16'd38170, 16'd32836, 16'd15133, 16'd29275, 16'd24536, 16'd42253, 16'd4503, 16'd17500, 16'd16906, 16'd62848, 16'd56831, 16'd10876, 16'd60003, 16'd56446, 16'd34119, 16'd53053, 16'd50002, 16'd30766, 16'd36832, 16'd9041, 16'd42191, 16'd7484, 16'd43417, 16'd61360, 16'd12832});
	test_expansion(128'hded609c235ee9afbe466a94193a2331e, {16'd13423, 16'd35243, 16'd35280, 16'd32844, 16'd44889, 16'd28598, 16'd14606, 16'd6531, 16'd11157, 16'd21270, 16'd25051, 16'd33823, 16'd35466, 16'd18448, 16'd2752, 16'd64345, 16'd34076, 16'd25975, 16'd1303, 16'd55192, 16'd48877, 16'd897, 16'd56812, 16'd55625, 16'd42363, 16'd43990});
	test_expansion(128'h84fac14d2b293fb762ade3dfe5a689e2, {16'd48723, 16'd42302, 16'd19300, 16'd15792, 16'd57026, 16'd58533, 16'd7412, 16'd79, 16'd34253, 16'd38281, 16'd8353, 16'd15393, 16'd34066, 16'd58863, 16'd55723, 16'd2762, 16'd60914, 16'd44293, 16'd30389, 16'd48935, 16'd22023, 16'd32416, 16'd44832, 16'd1512, 16'd43275, 16'd10236});
	test_expansion(128'h05bcc857d79ee942431b4c482b47cd29, {16'd42320, 16'd34849, 16'd5265, 16'd38821, 16'd12508, 16'd6599, 16'd29356, 16'd42335, 16'd34837, 16'd38124, 16'd26614, 16'd59720, 16'd49183, 16'd36690, 16'd62738, 16'd19088, 16'd21369, 16'd44556, 16'd48502, 16'd30257, 16'd26425, 16'd3181, 16'd59918, 16'd13068, 16'd8431, 16'd49551});
	test_expansion(128'he8af8a522b7edbb09a02ef2ec4480d02, {16'd36863, 16'd22638, 16'd6227, 16'd17738, 16'd42651, 16'd28902, 16'd41836, 16'd61264, 16'd2660, 16'd21780, 16'd17774, 16'd43825, 16'd36623, 16'd41490, 16'd45155, 16'd23905, 16'd52226, 16'd53700, 16'd12707, 16'd35303, 16'd16351, 16'd22357, 16'd59439, 16'd4835, 16'd54487, 16'd23210});
	test_expansion(128'ha4e4d802b6a7516cc8be899b0767ba8a, {16'd14251, 16'd23128, 16'd5104, 16'd35543, 16'd36072, 16'd53831, 16'd11995, 16'd36034, 16'd57578, 16'd63033, 16'd19566, 16'd4645, 16'd2384, 16'd24603, 16'd29805, 16'd27232, 16'd32699, 16'd13952, 16'd64088, 16'd23806, 16'd32700, 16'd45044, 16'd41416, 16'd32144, 16'd35009, 16'd27504});
	test_expansion(128'hc0a144783191d025ef6cce3b8805da40, {16'd17117, 16'd20676, 16'd50528, 16'd41437, 16'd29987, 16'd23065, 16'd21126, 16'd27475, 16'd47014, 16'd17700, 16'd29479, 16'd16408, 16'd61348, 16'd36487, 16'd44963, 16'd13803, 16'd51379, 16'd12824, 16'd39504, 16'd43933, 16'd27789, 16'd51856, 16'd25812, 16'd12529, 16'd19374, 16'd31248});
	test_expansion(128'h74856b1e2ca0c4d5210dfe95ce9c0aa2, {16'd19638, 16'd45125, 16'd53446, 16'd8519, 16'd48795, 16'd47230, 16'd35555, 16'd21721, 16'd64950, 16'd26264, 16'd39065, 16'd60780, 16'd40474, 16'd42295, 16'd63194, 16'd51292, 16'd6692, 16'd15743, 16'd63116, 16'd62768, 16'd31106, 16'd25239, 16'd16472, 16'd27616, 16'd46959, 16'd16713});
	test_expansion(128'h3cebe3ceaedee0c5d71df0656e93c4d2, {16'd49288, 16'd57446, 16'd8654, 16'd19513, 16'd10289, 16'd50164, 16'd39840, 16'd32121, 16'd31989, 16'd37276, 16'd19359, 16'd30754, 16'd11981, 16'd56858, 16'd51220, 16'd6945, 16'd3059, 16'd38511, 16'd27600, 16'd14376, 16'd28652, 16'd5012, 16'd1942, 16'd38279, 16'd39115, 16'd17885});
	test_expansion(128'h5b74ac4a5eedac6f7a37675387863a40, {16'd14799, 16'd9009, 16'd49236, 16'd30186, 16'd12513, 16'd9711, 16'd26244, 16'd20661, 16'd8241, 16'd44056, 16'd36298, 16'd5569, 16'd41459, 16'd32786, 16'd43521, 16'd10452, 16'd63890, 16'd24436, 16'd21349, 16'd39823, 16'd5945, 16'd23600, 16'd8184, 16'd3598, 16'd18230, 16'd35767});
	test_expansion(128'hcc08eed82ecd29ae2d2862b5f6658377, {16'd61793, 16'd16914, 16'd16830, 16'd59448, 16'd42087, 16'd28288, 16'd7964, 16'd48410, 16'd19018, 16'd10341, 16'd62871, 16'd56597, 16'd51325, 16'd51365, 16'd36955, 16'd43699, 16'd16505, 16'd3040, 16'd45432, 16'd32062, 16'd63977, 16'd4807, 16'd57589, 16'd62527, 16'd59977, 16'd3394});
	test_expansion(128'hc3c247a70b21f21384e02f7a56e047f9, {16'd34071, 16'd23095, 16'd12747, 16'd22971, 16'd20195, 16'd4271, 16'd46483, 16'd61473, 16'd49213, 16'd14059, 16'd2394, 16'd19906, 16'd52306, 16'd3624, 16'd62490, 16'd47603, 16'd16970, 16'd10341, 16'd26549, 16'd17067, 16'd9032, 16'd34078, 16'd6436, 16'd28834, 16'd40545, 16'd38056});
	test_expansion(128'hf41317a3885a865d7366d3e740d9f42a, {16'd7544, 16'd24327, 16'd18498, 16'd38223, 16'd9801, 16'd47151, 16'd12930, 16'd24897, 16'd48846, 16'd41693, 16'd5856, 16'd515, 16'd33563, 16'd20996, 16'd47325, 16'd50663, 16'd8674, 16'd51462, 16'd58098, 16'd60098, 16'd38432, 16'd29292, 16'd27213, 16'd64502, 16'd36665, 16'd50874});
	test_expansion(128'h361e7396da2a96b93915cb30b8cdc056, {16'd5130, 16'd49521, 16'd9456, 16'd47260, 16'd60027, 16'd30236, 16'd46995, 16'd35851, 16'd65336, 16'd26991, 16'd11145, 16'd56662, 16'd10184, 16'd19610, 16'd62358, 16'd53685, 16'd8930, 16'd24157, 16'd1226, 16'd21215, 16'd58215, 16'd38174, 16'd43984, 16'd11335, 16'd54945, 16'd57596});
	test_expansion(128'h387ed24a9048656be67937e8ea16eaae, {16'd36916, 16'd52215, 16'd11331, 16'd13329, 16'd60089, 16'd43238, 16'd2057, 16'd56396, 16'd25154, 16'd15330, 16'd63633, 16'd13807, 16'd19557, 16'd10524, 16'd57707, 16'd11719, 16'd41506, 16'd10108, 16'd17045, 16'd19666, 16'd46627, 16'd29047, 16'd35023, 16'd38625, 16'd59121, 16'd33684});
	test_expansion(128'h980b3289fb9751f4d17ab0df16b9c94d, {16'd32572, 16'd13646, 16'd3919, 16'd5982, 16'd60661, 16'd45643, 16'd5607, 16'd18369, 16'd36438, 16'd15260, 16'd30752, 16'd5581, 16'd29900, 16'd62546, 16'd61241, 16'd59501, 16'd14132, 16'd45741, 16'd16916, 16'd45154, 16'd61547, 16'd17400, 16'd44931, 16'd62985, 16'd36209, 16'd37409});
	test_expansion(128'he79ac3d31bde0e4c8f345fd010137b8a, {16'd43604, 16'd45693, 16'd48675, 16'd41253, 16'd623, 16'd26275, 16'd12805, 16'd39688, 16'd55098, 16'd1344, 16'd11662, 16'd25624, 16'd3818, 16'd853, 16'd44433, 16'd27840, 16'd60591, 16'd1765, 16'd33621, 16'd23212, 16'd50518, 16'd4890, 16'd40946, 16'd14243, 16'd62108, 16'd54861});
	test_expansion(128'h3be11a50ce9d4f6276b495cef2b24ab5, {16'd27167, 16'd20705, 16'd26982, 16'd4593, 16'd3046, 16'd22397, 16'd31671, 16'd18692, 16'd62367, 16'd13064, 16'd28389, 16'd2520, 16'd29690, 16'd38159, 16'd26752, 16'd19246, 16'd27474, 16'd39413, 16'd55141, 16'd1078, 16'd15260, 16'd44047, 16'd2830, 16'd12651, 16'd25459, 16'd38793});
	test_expansion(128'h2318646202476dda031426613f643f99, {16'd9841, 16'd27000, 16'd45695, 16'd18288, 16'd11618, 16'd12840, 16'd8180, 16'd811, 16'd15114, 16'd54495, 16'd52128, 16'd34857, 16'd40987, 16'd23801, 16'd53513, 16'd29919, 16'd42292, 16'd53013, 16'd36961, 16'd16828, 16'd12755, 16'd45508, 16'd5350, 16'd61988, 16'd35564, 16'd4809});
	test_expansion(128'hfc10e8232d44ca59a798185aa1f1b131, {16'd26556, 16'd50351, 16'd47814, 16'd23676, 16'd4890, 16'd19254, 16'd8985, 16'd50453, 16'd4954, 16'd47933, 16'd32835, 16'd57841, 16'd61699, 16'd40881, 16'd6239, 16'd5810, 16'd21913, 16'd12059, 16'd9428, 16'd30793, 16'd57059, 16'd39383, 16'd46352, 16'd23150, 16'd38025, 16'd39964});
	test_expansion(128'hc5264f8ed1887a16ecb5f9c232292d54, {16'd60573, 16'd37021, 16'd56284, 16'd28833, 16'd24358, 16'd32314, 16'd46979, 16'd17648, 16'd9637, 16'd28600, 16'd32334, 16'd23382, 16'd19155, 16'd9574, 16'd15504, 16'd36768, 16'd21347, 16'd62801, 16'd27533, 16'd19723, 16'd5038, 16'd47085, 16'd57505, 16'd54529, 16'd46544, 16'd28039});
	test_expansion(128'h8ecac3b0d76b18727b5d1dbe9e56b1df, {16'd8031, 16'd39438, 16'd6132, 16'd60214, 16'd54589, 16'd63406, 16'd35839, 16'd8391, 16'd57554, 16'd34989, 16'd14579, 16'd47933, 16'd41507, 16'd7806, 16'd34298, 16'd43992, 16'd41030, 16'd16196, 16'd6999, 16'd18780, 16'd58933, 16'd49882, 16'd61572, 16'd52471, 16'd47163, 16'd8816});
	test_expansion(128'h59fe26c423377de52b14c0438a8395eb, {16'd22492, 16'd20352, 16'd61380, 16'd48170, 16'd46697, 16'd42797, 16'd50440, 16'd62999, 16'd32350, 16'd34203, 16'd38314, 16'd2148, 16'd31135, 16'd32318, 16'd33673, 16'd37403, 16'd24996, 16'd47853, 16'd60409, 16'd57859, 16'd48517, 16'd63510, 16'd47173, 16'd30137, 16'd65210, 16'd42481});
	test_expansion(128'h55759a73e1c7dd4a7ac1e21546b5c78d, {16'd34649, 16'd910, 16'd33199, 16'd12751, 16'd54533, 16'd1709, 16'd44401, 16'd45054, 16'd61609, 16'd27417, 16'd30601, 16'd49963, 16'd32287, 16'd49006, 16'd12865, 16'd27670, 16'd42729, 16'd5408, 16'd50257, 16'd5274, 16'd310, 16'd54543, 16'd60136, 16'd46418, 16'd58650, 16'd51567});
	test_expansion(128'he910da2cf1fb369f21e2f8e313a0c452, {16'd55933, 16'd15976, 16'd2365, 16'd29779, 16'd12281, 16'd27436, 16'd31532, 16'd33564, 16'd41837, 16'd57376, 16'd33117, 16'd28317, 16'd26909, 16'd3023, 16'd58509, 16'd12010, 16'd20914, 16'd55260, 16'd27922, 16'd63320, 16'd28090, 16'd55110, 16'd33443, 16'd41901, 16'd7478, 16'd18090});
	test_expansion(128'hfc3b2c52391da058e0de49e2f687db11, {16'd30758, 16'd26556, 16'd18, 16'd38629, 16'd42097, 16'd26378, 16'd29456, 16'd24257, 16'd39440, 16'd26097, 16'd26002, 16'd59779, 16'd44704, 16'd22770, 16'd40292, 16'd47821, 16'd59960, 16'd14630, 16'd14071, 16'd55583, 16'd55680, 16'd44053, 16'd23532, 16'd61461, 16'd30655, 16'd16202});
	test_expansion(128'hb3c0ac0a0dec866b16bc65bd3d70ad60, {16'd44800, 16'd42085, 16'd52894, 16'd58926, 16'd32217, 16'd46443, 16'd51485, 16'd9886, 16'd32807, 16'd47299, 16'd22952, 16'd54953, 16'd60695, 16'd30259, 16'd36398, 16'd16995, 16'd2850, 16'd22355, 16'd52236, 16'd42478, 16'd36646, 16'd2208, 16'd17867, 16'd39882, 16'd9253, 16'd14035});
	test_expansion(128'h0c84ff03c646f63c5904e6aad9e4e56e, {16'd50692, 16'd17252, 16'd45296, 16'd56211, 16'd39047, 16'd25498, 16'd63510, 16'd9305, 16'd57738, 16'd58426, 16'd59824, 16'd56514, 16'd20217, 16'd27087, 16'd59207, 16'd37779, 16'd20815, 16'd22691, 16'd24121, 16'd64478, 16'd20946, 16'd29021, 16'd57811, 16'd40947, 16'd43147, 16'd62326});
	test_expansion(128'ha5c4f70ecc2c8b2baa8c7815968b450a, {16'd46966, 16'd21284, 16'd53601, 16'd46654, 16'd15437, 16'd61871, 16'd63420, 16'd37634, 16'd13998, 16'd47249, 16'd9090, 16'd22537, 16'd4917, 16'd31305, 16'd29949, 16'd6596, 16'd11289, 16'd228, 16'd64976, 16'd14982, 16'd35953, 16'd28116, 16'd36498, 16'd22403, 16'd29777, 16'd1894});
	test_expansion(128'h6ca5d49194e4edfd6c32b6420b031793, {16'd3278, 16'd6592, 16'd42775, 16'd900, 16'd43391, 16'd39948, 16'd14824, 16'd403, 16'd53244, 16'd38412, 16'd6937, 16'd16738, 16'd56657, 16'd851, 16'd31715, 16'd23298, 16'd44005, 16'd60166, 16'd3729, 16'd20465, 16'd28887, 16'd24452, 16'd31886, 16'd23151, 16'd46401, 16'd18396});
	test_expansion(128'h56cd6d6f01b19e6640bb89c52e5026c6, {16'd15914, 16'd57463, 16'd5843, 16'd55066, 16'd40321, 16'd5593, 16'd28273, 16'd10976, 16'd14141, 16'd54804, 16'd28353, 16'd12432, 16'd33127, 16'd62576, 16'd42200, 16'd1424, 16'd59648, 16'd3270, 16'd41918, 16'd11976, 16'd15071, 16'd22787, 16'd3614, 16'd13352, 16'd58199, 16'd56373});
	test_expansion(128'h93e8720b59cb0e0b2aec7d33f41187e1, {16'd38102, 16'd20243, 16'd58164, 16'd38414, 16'd10674, 16'd7593, 16'd44307, 16'd37604, 16'd54693, 16'd28565, 16'd45666, 16'd62036, 16'd8842, 16'd569, 16'd6460, 16'd60341, 16'd24864, 16'd41949, 16'd13744, 16'd11595, 16'd49125, 16'd17559, 16'd21411, 16'd20949, 16'd59200, 16'd62305});
	test_expansion(128'h14735b1e71cc805f005415d690500fb9, {16'd23294, 16'd19023, 16'd23026, 16'd17139, 16'd5942, 16'd15475, 16'd5093, 16'd13193, 16'd55964, 16'd15397, 16'd4619, 16'd18270, 16'd54976, 16'd7813, 16'd13917, 16'd28265, 16'd41384, 16'd15269, 16'd49250, 16'd33041, 16'd62613, 16'd50345, 16'd38491, 16'd1301, 16'd62374, 16'd40800});
	test_expansion(128'hce23953524f21e0ffd86adb36b4b07c8, {16'd4517, 16'd15395, 16'd8977, 16'd6796, 16'd22225, 16'd54181, 16'd61534, 16'd3711, 16'd63654, 16'd17698, 16'd26561, 16'd61085, 16'd46735, 16'd36788, 16'd38340, 16'd25452, 16'd6330, 16'd35524, 16'd37638, 16'd30278, 16'd30584, 16'd63365, 16'd37305, 16'd63125, 16'd27679, 16'd48517});
	test_expansion(128'h4439085d6e3c04c1d29a2a6349f10b19, {16'd30366, 16'd44870, 16'd47634, 16'd44465, 16'd23739, 16'd31757, 16'd23132, 16'd55380, 16'd32123, 16'd11846, 16'd61085, 16'd63041, 16'd41595, 16'd62633, 16'd62204, 16'd45978, 16'd36872, 16'd42087, 16'd32523, 16'd44912, 16'd48690, 16'd61549, 16'd48328, 16'd22883, 16'd9919, 16'd1571});
	test_expansion(128'hc482091896b1bfb5781f2ad58af5fd6f, {16'd7121, 16'd40809, 16'd62741, 16'd21526, 16'd24090, 16'd55095, 16'd52244, 16'd11345, 16'd54820, 16'd63436, 16'd59687, 16'd46872, 16'd63727, 16'd62503, 16'd32776, 16'd56877, 16'd21103, 16'd21893, 16'd48116, 16'd17478, 16'd38886, 16'd14151, 16'd6550, 16'd24731, 16'd30363, 16'd29510});
	test_expansion(128'hdc582f929193f895315473300c3d9529, {16'd41758, 16'd12131, 16'd39853, 16'd50315, 16'd33852, 16'd42952, 16'd23664, 16'd23034, 16'd42538, 16'd57452, 16'd61993, 16'd64299, 16'd15176, 16'd42969, 16'd21303, 16'd26905, 16'd28328, 16'd57665, 16'd8199, 16'd53127, 16'd58237, 16'd17080, 16'd26337, 16'd64550, 16'd43295, 16'd43342});
	test_expansion(128'h3710e899da2d8f46ff391971ae42af3c, {16'd41393, 16'd59179, 16'd40835, 16'd11974, 16'd64065, 16'd60696, 16'd24183, 16'd60479, 16'd26299, 16'd33181, 16'd51652, 16'd29633, 16'd9660, 16'd27866, 16'd52530, 16'd30087, 16'd62207, 16'd34684, 16'd19616, 16'd46520, 16'd49290, 16'd35956, 16'd6265, 16'd52369, 16'd3069, 16'd17551});
	test_expansion(128'h1985c1622d2dfe0c2bebc48a75d89701, {16'd52325, 16'd5886, 16'd54294, 16'd30512, 16'd20779, 16'd38577, 16'd22715, 16'd31654, 16'd44662, 16'd48929, 16'd14533, 16'd42244, 16'd34958, 16'd6215, 16'd56380, 16'd2484, 16'd3604, 16'd15288, 16'd8366, 16'd29558, 16'd9613, 16'd4384, 16'd40906, 16'd38031, 16'd45184, 16'd43159});
	test_expansion(128'h3ab6f1cf35f9004652065397f4b9f8ba, {16'd36085, 16'd60787, 16'd10170, 16'd24243, 16'd56743, 16'd10798, 16'd38135, 16'd38129, 16'd29506, 16'd4067, 16'd35801, 16'd29416, 16'd30028, 16'd7092, 16'd58597, 16'd10941, 16'd14412, 16'd22008, 16'd41433, 16'd39590, 16'd43287, 16'd39657, 16'd59519, 16'd22401, 16'd61334, 16'd17982});
	test_expansion(128'hd0351d2764e3e89b05d30c3dd3f666bc, {16'd7506, 16'd9681, 16'd55857, 16'd31135, 16'd41429, 16'd20138, 16'd46743, 16'd42572, 16'd41518, 16'd31546, 16'd9730, 16'd19966, 16'd12967, 16'd4182, 16'd60492, 16'd27984, 16'd21387, 16'd34709, 16'd37746, 16'd9537, 16'd57395, 16'd5644, 16'd58988, 16'd28375, 16'd64279, 16'd6994});
	test_expansion(128'habbb566322e4d20102f93ccdb1ad1aa8, {16'd38723, 16'd48842, 16'd60616, 16'd43572, 16'd37549, 16'd47304, 16'd1450, 16'd13115, 16'd27144, 16'd21006, 16'd2746, 16'd31565, 16'd64011, 16'd33817, 16'd5503, 16'd28496, 16'd15225, 16'd9884, 16'd63343, 16'd21297, 16'd52671, 16'd6011, 16'd54087, 16'd21737, 16'd63646, 16'd38838});
	test_expansion(128'h934dbf9ccddee54388c2417d43bfbd50, {16'd2120, 16'd3670, 16'd13325, 16'd33890, 16'd60457, 16'd12444, 16'd26043, 16'd12594, 16'd8502, 16'd51730, 16'd18194, 16'd28016, 16'd43642, 16'd61158, 16'd31903, 16'd30115, 16'd6311, 16'd7603, 16'd25479, 16'd57247, 16'd3108, 16'd2112, 16'd38032, 16'd9021, 16'd14246, 16'd27966});
	test_expansion(128'h2b7041907232cb190f122c7564985561, {16'd28887, 16'd6838, 16'd10395, 16'd59294, 16'd11080, 16'd61090, 16'd51723, 16'd34740, 16'd3113, 16'd13608, 16'd12523, 16'd41805, 16'd21985, 16'd12023, 16'd10240, 16'd5857, 16'd55777, 16'd14276, 16'd71, 16'd44633, 16'd23497, 16'd22396, 16'd58216, 16'd32905, 16'd18805, 16'd6899});
	test_expansion(128'ha0d893075cda68d8850b7d351bc30fe6, {16'd14687, 16'd34453, 16'd30862, 16'd42052, 16'd64461, 16'd62682, 16'd3708, 16'd18916, 16'd57534, 16'd64220, 16'd46322, 16'd25475, 16'd15827, 16'd21351, 16'd16338, 16'd29182, 16'd31292, 16'd45911, 16'd10129, 16'd28583, 16'd53152, 16'd57607, 16'd62672, 16'd6902, 16'd45321, 16'd35774});
	test_expansion(128'he490b607fc8fa72c6933fe5b2c1cbc78, {16'd43220, 16'd48601, 16'd32114, 16'd36869, 16'd10369, 16'd6461, 16'd53581, 16'd51390, 16'd61693, 16'd44204, 16'd18166, 16'd9963, 16'd57831, 16'd4060, 16'd9671, 16'd48445, 16'd33454, 16'd1190, 16'd1424, 16'd21002, 16'd220, 16'd65068, 16'd54470, 16'd36495, 16'd36494, 16'd59771});
	test_expansion(128'haa56a1c4248467b811b50d1acf00c7d4, {16'd18209, 16'd27415, 16'd45814, 16'd43826, 16'd62874, 16'd2809, 16'd40700, 16'd14002, 16'd29883, 16'd26319, 16'd6287, 16'd54658, 16'd37249, 16'd21439, 16'd36834, 16'd2915, 16'd60037, 16'd13772, 16'd58478, 16'd49089, 16'd50863, 16'd20760, 16'd61436, 16'd58594, 16'd49331, 16'd26711});
	test_expansion(128'hdaffd11129afc1ef073365b68192106e, {16'd1382, 16'd11666, 16'd24400, 16'd23800, 16'd28404, 16'd29726, 16'd18441, 16'd24850, 16'd5904, 16'd13340, 16'd27047, 16'd56462, 16'd5233, 16'd57337, 16'd54721, 16'd42603, 16'd34907, 16'd36344, 16'd55949, 16'd60758, 16'd46735, 16'd41936, 16'd52227, 16'd52219, 16'd35456, 16'd31035});
	test_expansion(128'hed1e12da15df5bd3c9b4ff13dacaa936, {16'd57743, 16'd52262, 16'd13987, 16'd31515, 16'd42219, 16'd59090, 16'd54437, 16'd36139, 16'd29582, 16'd55972, 16'd13007, 16'd52894, 16'd47390, 16'd56081, 16'd45172, 16'd22380, 16'd60606, 16'd64137, 16'd18167, 16'd26513, 16'd52573, 16'd28592, 16'd20645, 16'd19092, 16'd26063, 16'd64469});
	test_expansion(128'hdc003d570b34c6f602a25106894c917c, {16'd26631, 16'd53024, 16'd27929, 16'd44552, 16'd53913, 16'd37000, 16'd5288, 16'd14449, 16'd26258, 16'd43622, 16'd1399, 16'd63174, 16'd17222, 16'd31383, 16'd10465, 16'd35777, 16'd14387, 16'd33045, 16'd43488, 16'd9218, 16'd32045, 16'd55351, 16'd41948, 16'd35543, 16'd54114, 16'd25056});
	test_expansion(128'h56413c7e513175a12d7360c5e5c51aae, {16'd6704, 16'd56345, 16'd15075, 16'd49852, 16'd11604, 16'd14402, 16'd41561, 16'd16992, 16'd40104, 16'd46656, 16'd2379, 16'd54225, 16'd14728, 16'd58968, 16'd28948, 16'd40311, 16'd20973, 16'd6998, 16'd42420, 16'd48711, 16'd6960, 16'd31689, 16'd37121, 16'd5838, 16'd35291, 16'd37961});
	test_expansion(128'h3dc8f5e47f5417afb79facfb1135def9, {16'd60544, 16'd4899, 16'd48832, 16'd19788, 16'd17003, 16'd29673, 16'd15689, 16'd58305, 16'd8369, 16'd56402, 16'd21546, 16'd11733, 16'd5369, 16'd6950, 16'd29836, 16'd60118, 16'd48230, 16'd51266, 16'd54470, 16'd39632, 16'd1570, 16'd57219, 16'd39342, 16'd42400, 16'd33610, 16'd20652});
	test_expansion(128'heea2c7feb01571a9d6e9ae3c465828c1, {16'd62814, 16'd64714, 16'd2206, 16'd60323, 16'd44160, 16'd59674, 16'd46960, 16'd584, 16'd13258, 16'd434, 16'd22385, 16'd65020, 16'd56020, 16'd60365, 16'd52683, 16'd10453, 16'd11734, 16'd10359, 16'd63100, 16'd64755, 16'd55315, 16'd15162, 16'd5165, 16'd579, 16'd49770, 16'd47336});
	test_expansion(128'h697aeacd5075136097b6d0ffe94283a3, {16'd7581, 16'd11766, 16'd46498, 16'd20345, 16'd18364, 16'd12370, 16'd15867, 16'd20042, 16'd35654, 16'd41708, 16'd6578, 16'd58786, 16'd50750, 16'd27199, 16'd47272, 16'd38555, 16'd31872, 16'd60181, 16'd22844, 16'd21889, 16'd4972, 16'd11202, 16'd49467, 16'd7511, 16'd55630, 16'd32859});
	test_expansion(128'hf1ca1c0e4be20c2eaeaea32bd953feee, {16'd26340, 16'd52270, 16'd63550, 16'd27088, 16'd18590, 16'd13191, 16'd14605, 16'd59697, 16'd14108, 16'd23850, 16'd26276, 16'd36548, 16'd51780, 16'd59188, 16'd30872, 16'd41784, 16'd47687, 16'd49311, 16'd17053, 16'd10556, 16'd39403, 16'd56336, 16'd56570, 16'd40570, 16'd24749, 16'd51801});
	test_expansion(128'h07d98ec6c9e610e5b8c2e891efba3770, {16'd13186, 16'd48490, 16'd48744, 16'd29232, 16'd20072, 16'd29209, 16'd35572, 16'd25363, 16'd6115, 16'd277, 16'd39192, 16'd51970, 16'd43497, 16'd15547, 16'd17267, 16'd51966, 16'd28782, 16'd23837, 16'd35862, 16'd34546, 16'd39502, 16'd53917, 16'd50145, 16'd43913, 16'd123, 16'd27314});
	test_expansion(128'h88058320ec02dbe0ef98b75f071bf8ce, {16'd42665, 16'd13837, 16'd49701, 16'd22944, 16'd35409, 16'd38550, 16'd52607, 16'd39067, 16'd29374, 16'd16472, 16'd23937, 16'd51191, 16'd51060, 16'd54868, 16'd36370, 16'd18960, 16'd18811, 16'd8940, 16'd61279, 16'd25236, 16'd40937, 16'd64775, 16'd57937, 16'd46056, 16'd64314, 16'd48071});
	test_expansion(128'hb0c9093280383dc697568b63c281dd93, {16'd51081, 16'd48163, 16'd35239, 16'd4192, 16'd25918, 16'd45412, 16'd29896, 16'd40064, 16'd58066, 16'd1255, 16'd59450, 16'd70, 16'd7950, 16'd57227, 16'd19120, 16'd19792, 16'd57576, 16'd32554, 16'd18938, 16'd16404, 16'd10779, 16'd15946, 16'd49892, 16'd11034, 16'd7310, 16'd64029});
	test_expansion(128'h3c05699d303adf503b24adbd8928c8d4, {16'd34847, 16'd54934, 16'd26774, 16'd22370, 16'd62166, 16'd40271, 16'd17676, 16'd15209, 16'd23869, 16'd9172, 16'd57543, 16'd18682, 16'd55231, 16'd55913, 16'd56990, 16'd42435, 16'd41212, 16'd58193, 16'd39155, 16'd36821, 16'd58751, 16'd22564, 16'd45854, 16'd49783, 16'd18746, 16'd14923});
	test_expansion(128'h7c16442875475123385f5b9385913554, {16'd56729, 16'd29576, 16'd27396, 16'd13602, 16'd56536, 16'd54092, 16'd51319, 16'd52496, 16'd19409, 16'd13822, 16'd15, 16'd20708, 16'd64688, 16'd39987, 16'd34643, 16'd29471, 16'd50077, 16'd40836, 16'd25798, 16'd39929, 16'd22723, 16'd16522, 16'd32899, 16'd34321, 16'd6278, 16'd48});
	test_expansion(128'h17c5be19436b38f2f60dfb94d6b558ee, {16'd18125, 16'd17950, 16'd48628, 16'd11937, 16'd14204, 16'd24708, 16'd27818, 16'd21504, 16'd13000, 16'd48875, 16'd45826, 16'd30499, 16'd4432, 16'd2430, 16'd12476, 16'd64090, 16'd18838, 16'd60501, 16'd13192, 16'd58858, 16'd21977, 16'd9946, 16'd53997, 16'd41312, 16'd62736, 16'd40264});
	test_expansion(128'h2688661536c5d656c82b11b279e32877, {16'd9813, 16'd25683, 16'd710, 16'd7003, 16'd23946, 16'd5668, 16'd8883, 16'd3397, 16'd64643, 16'd41335, 16'd34863, 16'd36634, 16'd33647, 16'd13780, 16'd16313, 16'd51368, 16'd46822, 16'd7749, 16'd9639, 16'd1338, 16'd10446, 16'd63043, 16'd56440, 16'd29378, 16'd62535, 16'd25654});
	test_expansion(128'h76c286c41eb63f2a8cb705465ed0d9d7, {16'd52570, 16'd26585, 16'd564, 16'd21390, 16'd20738, 16'd27102, 16'd40880, 16'd46373, 16'd43045, 16'd60856, 16'd58572, 16'd12342, 16'd59584, 16'd46448, 16'd22037, 16'd51917, 16'd4455, 16'd49884, 16'd15468, 16'd30681, 16'd50005, 16'd48528, 16'd59480, 16'd35463, 16'd6096, 16'd259});
	test_expansion(128'h94e2b53fa5723e238146a12e790379c3, {16'd27720, 16'd58396, 16'd13452, 16'd7767, 16'd13954, 16'd23619, 16'd28954, 16'd14365, 16'd2922, 16'd14638, 16'd37752, 16'd29155, 16'd53559, 16'd10729, 16'd52453, 16'd58897, 16'd18862, 16'd47829, 16'd27203, 16'd44278, 16'd62864, 16'd36347, 16'd10286, 16'd33435, 16'd35928, 16'd24908});
	test_expansion(128'hfd6d101d7aa35f2cdcd5efa12d511b72, {16'd36438, 16'd47049, 16'd25734, 16'd13787, 16'd50394, 16'd57630, 16'd21941, 16'd38523, 16'd22388, 16'd47798, 16'd6023, 16'd31195, 16'd35314, 16'd60567, 16'd59845, 16'd50114, 16'd46431, 16'd35496, 16'd16951, 16'd41724, 16'd40338, 16'd56576, 16'd10712, 16'd38571, 16'd57152, 16'd24494});
	test_expansion(128'h4b4d0edb645356e2889a0790833637e7, {16'd51618, 16'd34342, 16'd58609, 16'd35778, 16'd47015, 16'd8421, 16'd27523, 16'd14462, 16'd63073, 16'd15722, 16'd996, 16'd21980, 16'd14682, 16'd47669, 16'd43780, 16'd58405, 16'd16829, 16'd38657, 16'd39517, 16'd32215, 16'd62644, 16'd30288, 16'd65478, 16'd10847, 16'd35252, 16'd3242});
	test_expansion(128'hffdb6a45181e408cece0828301095fc6, {16'd32094, 16'd6205, 16'd38013, 16'd31526, 16'd43136, 16'd7869, 16'd49476, 16'd17200, 16'd6909, 16'd45224, 16'd5761, 16'd53098, 16'd51327, 16'd47583, 16'd47613, 16'd63424, 16'd42970, 16'd26089, 16'd28453, 16'd44338, 16'd53726, 16'd65049, 16'd46329, 16'd19323, 16'd12607, 16'd15158});
	test_expansion(128'h3b93f70c9c6e44b3fd38864f21970089, {16'd23, 16'd34491, 16'd37763, 16'd9687, 16'd42040, 16'd14636, 16'd35939, 16'd38204, 16'd38236, 16'd15529, 16'd46648, 16'd60097, 16'd56846, 16'd8340, 16'd12049, 16'd27163, 16'd59580, 16'd2217, 16'd37894, 16'd19859, 16'd26424, 16'd50170, 16'd14016, 16'd13591, 16'd44504, 16'd61177});
	test_expansion(128'h230ed7c3da80e5936c5d698712c67957, {16'd20925, 16'd25106, 16'd23064, 16'd23933, 16'd53429, 16'd21445, 16'd26593, 16'd30048, 16'd35745, 16'd56247, 16'd10601, 16'd24785, 16'd856, 16'd46006, 16'd49435, 16'd26579, 16'd10754, 16'd23494, 16'd25064, 16'd59025, 16'd23122, 16'd11197, 16'd35761, 16'd25212, 16'd190, 16'd10707});
	test_expansion(128'h0757d12882311e11ff49ce4d9c976668, {16'd59780, 16'd37296, 16'd26722, 16'd61103, 16'd26878, 16'd33778, 16'd38231, 16'd33329, 16'd652, 16'd8921, 16'd45583, 16'd13502, 16'd45118, 16'd44326, 16'd57671, 16'd44382, 16'd22203, 16'd19230, 16'd40933, 16'd57459, 16'd13877, 16'd49324, 16'd56020, 16'd35380, 16'd44209, 16'd5778});
	test_expansion(128'hcbd995f199f011f12d7a371cd6d4aba4, {16'd22268, 16'd34776, 16'd49530, 16'd32203, 16'd56157, 16'd10998, 16'd48686, 16'd19988, 16'd20174, 16'd7365, 16'd8103, 16'd8479, 16'd25875, 16'd7929, 16'd52766, 16'd18834, 16'd11471, 16'd6531, 16'd52850, 16'd48388, 16'd39965, 16'd35131, 16'd26015, 16'd54202, 16'd1860, 16'd36611});
	test_expansion(128'h03b4a72bc25b973eef1dcb03012d4505, {16'd30583, 16'd3483, 16'd30260, 16'd40536, 16'd23289, 16'd19968, 16'd28015, 16'd9832, 16'd53787, 16'd25031, 16'd44437, 16'd56194, 16'd3353, 16'd14063, 16'd22439, 16'd2571, 16'd62728, 16'd44399, 16'd56759, 16'd8805, 16'd48498, 16'd9773, 16'd49064, 16'd6999, 16'd53828, 16'd33234});
	test_expansion(128'h98be04dcfe447700562dc0e86487520e, {16'd26230, 16'd6225, 16'd24534, 16'd21402, 16'd21698, 16'd14731, 16'd7247, 16'd1968, 16'd43878, 16'd17691, 16'd22714, 16'd15299, 16'd24370, 16'd14708, 16'd23181, 16'd28353, 16'd45784, 16'd15185, 16'd64520, 16'd10878, 16'd8524, 16'd23432, 16'd39375, 16'd7330, 16'd49661, 16'd49413});
	test_expansion(128'h2878259ce062545ccd1437722f48d8d4, {16'd23973, 16'd64832, 16'd4588, 16'd15169, 16'd47040, 16'd59078, 16'd47833, 16'd14277, 16'd22001, 16'd37908, 16'd65275, 16'd6584, 16'd54451, 16'd17791, 16'd50506, 16'd59452, 16'd32646, 16'd5101, 16'd48978, 16'd9547, 16'd63665, 16'd17334, 16'd16489, 16'd22142, 16'd23607, 16'd61060});
	test_expansion(128'hca18e6081705e69ea4897e6a67326291, {16'd55258, 16'd237, 16'd11595, 16'd29127, 16'd56391, 16'd28530, 16'd47469, 16'd6223, 16'd48784, 16'd53146, 16'd42701, 16'd41411, 16'd57462, 16'd58815, 16'd5709, 16'd12734, 16'd53089, 16'd34923, 16'd22021, 16'd13958, 16'd30719, 16'd41127, 16'd62614, 16'd11720, 16'd28210, 16'd42674});
	test_expansion(128'h7ce1117ba857951602099a7672dc6599, {16'd11716, 16'd60693, 16'd13236, 16'd54418, 16'd3864, 16'd46889, 16'd6583, 16'd59476, 16'd41100, 16'd20873, 16'd4157, 16'd1744, 16'd45700, 16'd43490, 16'd56780, 16'd51344, 16'd6768, 16'd36045, 16'd54314, 16'd38022, 16'd48258, 16'd31048, 16'd11912, 16'd26237, 16'd15352, 16'd50608});
	test_expansion(128'h1187ec445702d94a8dd7679187ea47d9, {16'd41521, 16'd60708, 16'd17719, 16'd32303, 16'd23806, 16'd41277, 16'd46713, 16'd22890, 16'd13323, 16'd10449, 16'd36117, 16'd31154, 16'd23452, 16'd57928, 16'd18504, 16'd50762, 16'd63898, 16'd38011, 16'd12441, 16'd48472, 16'd23174, 16'd20639, 16'd8049, 16'd4894, 16'd33633, 16'd47716});
	test_expansion(128'hf356d801a4615cc4b5b40f221e98fd49, {16'd63438, 16'd42300, 16'd46087, 16'd29366, 16'd40827, 16'd21202, 16'd22564, 16'd58171, 16'd48524, 16'd9216, 16'd36818, 16'd5977, 16'd49948, 16'd42010, 16'd57933, 16'd25196, 16'd59665, 16'd36371, 16'd63097, 16'd43109, 16'd7341, 16'd43794, 16'd14667, 16'd21486, 16'd20309, 16'd29601});
	test_expansion(128'h62f53444da9a0659e56fe4afac127000, {16'd24657, 16'd62461, 16'd6972, 16'd45352, 16'd8819, 16'd4384, 16'd23653, 16'd22479, 16'd36274, 16'd44575, 16'd28377, 16'd4378, 16'd38248, 16'd32587, 16'd65247, 16'd32708, 16'd32951, 16'd16778, 16'd35169, 16'd38940, 16'd63312, 16'd22333, 16'd53387, 16'd24844, 16'd46362, 16'd4472});
	test_expansion(128'hc497c28dfd02e9cfb798d4216aea1353, {16'd13447, 16'd14261, 16'd35008, 16'd23696, 16'd12782, 16'd13505, 16'd17037, 16'd18802, 16'd4214, 16'd59382, 16'd46776, 16'd4918, 16'd56512, 16'd25686, 16'd18374, 16'd21575, 16'd38864, 16'd3193, 16'd6653, 16'd17034, 16'd11421, 16'd41915, 16'd48349, 16'd58130, 16'd55990, 16'd16708});
	test_expansion(128'h4ed84fae86c3fcb35efe96b6731da69c, {16'd811, 16'd43549, 16'd45556, 16'd13992, 16'd22955, 16'd58517, 16'd38222, 16'd57377, 16'd65114, 16'd62799, 16'd371, 16'd38725, 16'd10607, 16'd16932, 16'd64264, 16'd61498, 16'd40238, 16'd62726, 16'd5552, 16'd26923, 16'd47205, 16'd6200, 16'd37813, 16'd14038, 16'd50757, 16'd32909});
	test_expansion(128'h3e5c68d0771149ba2b77be2a36fe89ca, {16'd43732, 16'd52813, 16'd4094, 16'd62322, 16'd18909, 16'd42177, 16'd57774, 16'd3403, 16'd49193, 16'd15910, 16'd63695, 16'd7347, 16'd65057, 16'd49869, 16'd36623, 16'd34376, 16'd52116, 16'd3663, 16'd56733, 16'd33314, 16'd23992, 16'd44631, 16'd22327, 16'd46057, 16'd49466, 16'd60550});
	test_expansion(128'h84d2bb2964191f96f9abbac09ee74c51, {16'd24626, 16'd16954, 16'd41242, 16'd29, 16'd51477, 16'd57319, 16'd13530, 16'd22174, 16'd17924, 16'd41519, 16'd62770, 16'd32355, 16'd48220, 16'd34367, 16'd21670, 16'd6822, 16'd52996, 16'd16844, 16'd35072, 16'd31485, 16'd12035, 16'd6994, 16'd11274, 16'd11705, 16'd29601, 16'd22862});
	test_expansion(128'h8112bc2b47f1bfc38ab27446e75e0717, {16'd61337, 16'd26372, 16'd20981, 16'd33232, 16'd35001, 16'd60158, 16'd49370, 16'd34832, 16'd9200, 16'd64503, 16'd48734, 16'd11693, 16'd49842, 16'd56036, 16'd19235, 16'd48936, 16'd51640, 16'd58357, 16'd7190, 16'd38724, 16'd21425, 16'd59545, 16'd48284, 16'd19880, 16'd37203, 16'd38874});
	test_expansion(128'h3fc9588d45e758a52f241b296f27d1ec, {16'd41915, 16'd51024, 16'd14834, 16'd8543, 16'd50629, 16'd22958, 16'd56111, 16'd25426, 16'd5912, 16'd33127, 16'd26199, 16'd11331, 16'd17604, 16'd48598, 16'd43461, 16'd226, 16'd34071, 16'd50061, 16'd11454, 16'd29480, 16'd62003, 16'd15819, 16'd32720, 16'd39276, 16'd40759, 16'd41047});
	test_expansion(128'h5be266131eda15c6815a736b101082ba, {16'd47126, 16'd18799, 16'd35717, 16'd64918, 16'd62474, 16'd21608, 16'd33372, 16'd45428, 16'd64398, 16'd13118, 16'd17643, 16'd63944, 16'd50514, 16'd38479, 16'd60441, 16'd35838, 16'd63093, 16'd57355, 16'd34329, 16'd32717, 16'd54329, 16'd53973, 16'd45988, 16'd4181, 16'd28396, 16'd30940});
	test_expansion(128'h43d04059b9a14fc58392899530458859, {16'd17309, 16'd6118, 16'd61447, 16'd43012, 16'd8624, 16'd1445, 16'd44503, 16'd42615, 16'd37151, 16'd62808, 16'd34330, 16'd53072, 16'd3006, 16'd38469, 16'd13771, 16'd37675, 16'd28277, 16'd8668, 16'd31696, 16'd38700, 16'd4965, 16'd58909, 16'd54343, 16'd49222, 16'd46184, 16'd23641});
	test_expansion(128'hcde622b1a264b44203e2664f4aa231a4, {16'd8830, 16'd62942, 16'd12957, 16'd5573, 16'd16815, 16'd51334, 16'd23721, 16'd15263, 16'd51977, 16'd45541, 16'd53959, 16'd7487, 16'd39513, 16'd3818, 16'd48068, 16'd52798, 16'd12222, 16'd54822, 16'd32864, 16'd37729, 16'd31236, 16'd23595, 16'd44552, 16'd28486, 16'd35130, 16'd7485});
	test_expansion(128'hd4770c41b24afd45d22d031fa53bc821, {16'd5036, 16'd40072, 16'd64738, 16'd45005, 16'd28846, 16'd33680, 16'd27662, 16'd4889, 16'd40902, 16'd55854, 16'd10635, 16'd33320, 16'd7128, 16'd55160, 16'd30759, 16'd56837, 16'd14881, 16'd54027, 16'd29310, 16'd38575, 16'd36140, 16'd35315, 16'd45639, 16'd53124, 16'd6286, 16'd4209});
	test_expansion(128'h4bffe95f88618b435f7cf8a940da27a7, {16'd29846, 16'd61145, 16'd61412, 16'd60178, 16'd6693, 16'd37274, 16'd20018, 16'd63204, 16'd33373, 16'd29008, 16'd38027, 16'd39295, 16'd48263, 16'd45009, 16'd26974, 16'd8896, 16'd29576, 16'd59870, 16'd31374, 16'd28435, 16'd4961, 16'd34590, 16'd957, 16'd34144, 16'd60447, 16'd63489});
	test_expansion(128'h308fb53b005496f0981dad746b225c71, {16'd53281, 16'd50162, 16'd18087, 16'd62271, 16'd47194, 16'd49731, 16'd58827, 16'd41576, 16'd53974, 16'd47053, 16'd32002, 16'd65142, 16'd62479, 16'd7275, 16'd61416, 16'd13978, 16'd44362, 16'd45732, 16'd14204, 16'd59127, 16'd27745, 16'd10774, 16'd54200, 16'd46751, 16'd11436, 16'd26934});
	test_expansion(128'h6ef744140b05bb80fa28eae03c6426ff, {16'd9571, 16'd62600, 16'd29079, 16'd19898, 16'd26563, 16'd17847, 16'd55384, 16'd42286, 16'd54708, 16'd29774, 16'd54790, 16'd38572, 16'd23467, 16'd10675, 16'd2617, 16'd2889, 16'd38888, 16'd40753, 16'd63855, 16'd28290, 16'd50013, 16'd35737, 16'd11075, 16'd54129, 16'd40745, 16'd3263});
	test_expansion(128'h950e451da27be8c5f9a0a36def6e047e, {16'd62801, 16'd61263, 16'd10329, 16'd30302, 16'd42010, 16'd56700, 16'd53533, 16'd63912, 16'd65490, 16'd7707, 16'd1746, 16'd7101, 16'd17416, 16'd39421, 16'd32209, 16'd24675, 16'd41877, 16'd2455, 16'd14727, 16'd59394, 16'd32404, 16'd2672, 16'd13288, 16'd65477, 16'd45861, 16'd57616});
	test_expansion(128'hde2be0c36e8da516c6157ac9a3a2c630, {16'd46858, 16'd2382, 16'd13878, 16'd11692, 16'd56892, 16'd54930, 16'd3428, 16'd62517, 16'd235, 16'd54233, 16'd27022, 16'd36605, 16'd56924, 16'd37691, 16'd31587, 16'd17243, 16'd58718, 16'd1380, 16'd34831, 16'd48156, 16'd50809, 16'd27785, 16'd63366, 16'd21314, 16'd46672, 16'd56370});
	test_expansion(128'h3eb424d13ec9d9217669f32076b40b7a, {16'd8813, 16'd48057, 16'd29173, 16'd7691, 16'd49611, 16'd48875, 16'd41666, 16'd29433, 16'd22429, 16'd29997, 16'd34314, 16'd32539, 16'd53960, 16'd35381, 16'd22313, 16'd53478, 16'd10273, 16'd44463, 16'd28748, 16'd17299, 16'd52458, 16'd20099, 16'd52202, 16'd49247, 16'd41366, 16'd50026});
	test_expansion(128'h049ca5bc07d2c41d274af7dd864485e1, {16'd43724, 16'd8116, 16'd5209, 16'd27222, 16'd35264, 16'd10306, 16'd59468, 16'd25592, 16'd35474, 16'd45906, 16'd16969, 16'd16698, 16'd57673, 16'd46264, 16'd42444, 16'd32710, 16'd3965, 16'd10487, 16'd39996, 16'd21889, 16'd31834, 16'd60881, 16'd46400, 16'd12535, 16'd60214, 16'd15845});
	test_expansion(128'h20621ad9cf11f3d4e8454006c7157ef7, {16'd4503, 16'd35751, 16'd27616, 16'd41680, 16'd39011, 16'd54456, 16'd3099, 16'd41634, 16'd59791, 16'd47957, 16'd5837, 16'd17890, 16'd47281, 16'd52528, 16'd54597, 16'd20589, 16'd20805, 16'd59731, 16'd1313, 16'd64042, 16'd10972, 16'd18159, 16'd46601, 16'd49175, 16'd42005, 16'd20704});
	test_expansion(128'h9dae6aac120e9e471642900fd4f5df5d, {16'd52111, 16'd48446, 16'd42846, 16'd58013, 16'd6861, 16'd8906, 16'd8928, 16'd54770, 16'd51213, 16'd39204, 16'd40948, 16'd42455, 16'd63868, 16'd45211, 16'd5041, 16'd37913, 16'd3240, 16'd51292, 16'd26403, 16'd2166, 16'd13718, 16'd3748, 16'd43818, 16'd15875, 16'd62706, 16'd57791});
	test_expansion(128'hbb74f53a515b7bc7f7c3f0c828f152fb, {16'd47023, 16'd23381, 16'd64406, 16'd57919, 16'd56525, 16'd11339, 16'd26030, 16'd9507, 16'd12573, 16'd29444, 16'd31908, 16'd45701, 16'd50416, 16'd22693, 16'd40492, 16'd28633, 16'd58436, 16'd27008, 16'd4772, 16'd51330, 16'd53071, 16'd12222, 16'd8942, 16'd28212, 16'd12526, 16'd39375});
	test_expansion(128'h1d83411d707d3404e509b46da3345f94, {16'd16468, 16'd57205, 16'd60815, 16'd26233, 16'd43368, 16'd51594, 16'd50994, 16'd22728, 16'd16883, 16'd21189, 16'd49758, 16'd46679, 16'd10930, 16'd41801, 16'd37537, 16'd35049, 16'd55847, 16'd54397, 16'd39213, 16'd55815, 16'd49464, 16'd3479, 16'd30588, 16'd65262, 16'd42255, 16'd28811});
	test_expansion(128'h91f3dafbba5d7c89f975c6b71e15eacc, {16'd11282, 16'd15202, 16'd23653, 16'd8343, 16'd45168, 16'd24147, 16'd64955, 16'd51364, 16'd27307, 16'd15780, 16'd60544, 16'd48508, 16'd31877, 16'd4893, 16'd32151, 16'd58842, 16'd16428, 16'd3994, 16'd2568, 16'd42756, 16'd40617, 16'd3854, 16'd31885, 16'd23027, 16'd64916, 16'd61089});
	test_expansion(128'h643d58790ed70a2d01d6a250aee7ab3e, {16'd35678, 16'd15028, 16'd26215, 16'd63664, 16'd4214, 16'd64802, 16'd57251, 16'd47116, 16'd10867, 16'd28668, 16'd37539, 16'd32837, 16'd22426, 16'd38658, 16'd48803, 16'd31982, 16'd49372, 16'd49845, 16'd58535, 16'd53040, 16'd63320, 16'd25014, 16'd32753, 16'd1388, 16'd17243, 16'd2663});
	test_expansion(128'h7f9b064c62c531878074a7b080b94458, {16'd40557, 16'd16531, 16'd30360, 16'd35998, 16'd21116, 16'd34946, 16'd51948, 16'd46171, 16'd4073, 16'd56602, 16'd48226, 16'd7195, 16'd4902, 16'd33561, 16'd57892, 16'd32025, 16'd35092, 16'd11983, 16'd44276, 16'd42070, 16'd48900, 16'd41477, 16'd2467, 16'd27195, 16'd26278, 16'd27467});
	test_expansion(128'h7c6e00b89c625054c020c1f088916da6, {16'd44936, 16'd37209, 16'd47664, 16'd34898, 16'd43205, 16'd23776, 16'd29730, 16'd947, 16'd5705, 16'd38472, 16'd42564, 16'd43562, 16'd20228, 16'd56430, 16'd10230, 16'd35920, 16'd21681, 16'd4633, 16'd24186, 16'd24686, 16'd3850, 16'd35972, 16'd40883, 16'd28412, 16'd51094, 16'd45659});
	test_expansion(128'had5be7d584f50a9a7e2a6b4cc213a0e2, {16'd20384, 16'd22241, 16'd43990, 16'd27439, 16'd58562, 16'd22359, 16'd36622, 16'd60994, 16'd36224, 16'd51434, 16'd44341, 16'd9974, 16'd1487, 16'd27753, 16'd62006, 16'd63985, 16'd45204, 16'd9147, 16'd43484, 16'd6989, 16'd7751, 16'd23079, 16'd35191, 16'd38391, 16'd2604, 16'd52634});
	test_expansion(128'ha0f610d09b287643830aefbdd2cd4fd8, {16'd23064, 16'd22507, 16'd51634, 16'd20892, 16'd35702, 16'd944, 16'd34170, 16'd38974, 16'd23806, 16'd313, 16'd37605, 16'd373, 16'd63435, 16'd24536, 16'd38269, 16'd7213, 16'd49098, 16'd34252, 16'd39457, 16'd60853, 16'd2434, 16'd53853, 16'd23747, 16'd63880, 16'd11227, 16'd43091});
	test_expansion(128'hf86b19a6b9501990a111bfc560c92921, {16'd45202, 16'd56867, 16'd57092, 16'd36528, 16'd19915, 16'd44789, 16'd8446, 16'd7345, 16'd33181, 16'd15450, 16'd14221, 16'd32260, 16'd4956, 16'd14637, 16'd477, 16'd48498, 16'd3955, 16'd41995, 16'd1370, 16'd25520, 16'd57062, 16'd37195, 16'd43905, 16'd27757, 16'd42473, 16'd5363});
	test_expansion(128'h3644e22f456085f42c8c04b30f55c3f6, {16'd41968, 16'd31683, 16'd21972, 16'd1506, 16'd22597, 16'd60071, 16'd4168, 16'd13858, 16'd14705, 16'd36091, 16'd43620, 16'd12625, 16'd14928, 16'd10385, 16'd47034, 16'd50521, 16'd24645, 16'd4095, 16'd38296, 16'd47382, 16'd3106, 16'd25521, 16'd51187, 16'd19354, 16'd18000, 16'd45375});
	test_expansion(128'hfaa7f59f590caf6856c22046552df815, {16'd14332, 16'd32409, 16'd20344, 16'd29158, 16'd55987, 16'd15794, 16'd24990, 16'd15283, 16'd48644, 16'd54774, 16'd38440, 16'd50822, 16'd51487, 16'd35336, 16'd32711, 16'd33508, 16'd5641, 16'd10263, 16'd23883, 16'd13594, 16'd54793, 16'd42390, 16'd29223, 16'd32688, 16'd37131, 16'd8330});
	test_expansion(128'h908289a67db72c1dcf29473a4eea4c87, {16'd1132, 16'd31419, 16'd15819, 16'd28441, 16'd27370, 16'd2911, 16'd9331, 16'd22638, 16'd49197, 16'd38934, 16'd50253, 16'd12142, 16'd45472, 16'd46098, 16'd46693, 16'd56630, 16'd24818, 16'd22215, 16'd2042, 16'd20221, 16'd35611, 16'd12331, 16'd8390, 16'd13541, 16'd60302, 16'd43324});
	test_expansion(128'h7301683d00d1c9744a5dc7a8f97747e6, {16'd29077, 16'd44516, 16'd10281, 16'd61169, 16'd23479, 16'd40595, 16'd43664, 16'd13704, 16'd50809, 16'd43057, 16'd38259, 16'd54523, 16'd6032, 16'd50375, 16'd42306, 16'd63704, 16'd3229, 16'd5600, 16'd53953, 16'd31878, 16'd6195, 16'd3856, 16'd65336, 16'd40822, 16'd25718, 16'd56308});
	test_expansion(128'h5555c25986cd22bfc85eb46ddba5c3bf, {16'd21411, 16'd43645, 16'd56592, 16'd42276, 16'd45291, 16'd38484, 16'd46524, 16'd5529, 16'd43637, 16'd15399, 16'd48300, 16'd39037, 16'd19176, 16'd22653, 16'd46661, 16'd30583, 16'd63166, 16'd65516, 16'd16011, 16'd48965, 16'd18075, 16'd26585, 16'd44803, 16'd51782, 16'd31263, 16'd60702});
	test_expansion(128'he17b11657e8aad9b13e9c66facf5cea5, {16'd43145, 16'd30878, 16'd63099, 16'd1996, 16'd57074, 16'd14366, 16'd63281, 16'd21266, 16'd51075, 16'd1999, 16'd56063, 16'd63568, 16'd49493, 16'd5571, 16'd10129, 16'd39019, 16'd45769, 16'd37651, 16'd4068, 16'd44837, 16'd11990, 16'd3275, 16'd54999, 16'd19838, 16'd6201, 16'd16389});
	test_expansion(128'h2535035d76337b1cf3bb171200fc4045, {16'd15052, 16'd11342, 16'd39299, 16'd45232, 16'd2372, 16'd38557, 16'd53401, 16'd55339, 16'd37108, 16'd16536, 16'd36480, 16'd16832, 16'd17342, 16'd10869, 16'd6399, 16'd15306, 16'd5271, 16'd54478, 16'd28738, 16'd51030, 16'd4539, 16'd39986, 16'd15168, 16'd20403, 16'd55279, 16'd34809});
	test_expansion(128'hb9853e9e1f9e5129aaaab2a4fb21e0e7, {16'd19746, 16'd47103, 16'd24494, 16'd19745, 16'd28562, 16'd12651, 16'd41228, 16'd4196, 16'd31979, 16'd9798, 16'd56807, 16'd52086, 16'd56110, 16'd12711, 16'd3952, 16'd58140, 16'd3128, 16'd37782, 16'd37060, 16'd36892, 16'd56683, 16'd2385, 16'd18477, 16'd52028, 16'd63303, 16'd49014});
	test_expansion(128'h3c753c4acde95059313be0060769cdcc, {16'd52125, 16'd22792, 16'd8452, 16'd17117, 16'd46088, 16'd17678, 16'd35308, 16'd39746, 16'd37073, 16'd39164, 16'd48403, 16'd17573, 16'd1318, 16'd34775, 16'd45328, 16'd52967, 16'd28321, 16'd24190, 16'd9900, 16'd19833, 16'd60316, 16'd47044, 16'd21562, 16'd48080, 16'd49958, 16'd24228});
	test_expansion(128'h33e0488bdfba0caa9c8409f08dae04ce, {16'd26479, 16'd64037, 16'd62372, 16'd18689, 16'd11862, 16'd26715, 16'd44032, 16'd39355, 16'd10233, 16'd7882, 16'd34231, 16'd16987, 16'd49337, 16'd6113, 16'd43476, 16'd58752, 16'd12741, 16'd16971, 16'd39141, 16'd52527, 16'd7557, 16'd29004, 16'd59302, 16'd36329, 16'd8557, 16'd33721});
	test_expansion(128'haf0d419c6a8f0066987433f5dcd025e9, {16'd20806, 16'd2421, 16'd54722, 16'd25627, 16'd15775, 16'd38271, 16'd51558, 16'd18617, 16'd65265, 16'd47949, 16'd1100, 16'd36161, 16'd57887, 16'd46597, 16'd42682, 16'd35840, 16'd34220, 16'd17166, 16'd52582, 16'd19975, 16'd63272, 16'd43818, 16'd6485, 16'd44498, 16'd35687, 16'd3312});
	test_expansion(128'h3b81cd38d5a329fb2748229e0a5cd6fa, {16'd21240, 16'd13991, 16'd48716, 16'd27129, 16'd32530, 16'd27328, 16'd57490, 16'd59054, 16'd22336, 16'd36735, 16'd39631, 16'd22548, 16'd57536, 16'd52981, 16'd29493, 16'd47512, 16'd35589, 16'd36666, 16'd32910, 16'd11872, 16'd38661, 16'd44086, 16'd3566, 16'd4032, 16'd54682, 16'd49965});
	test_expansion(128'he0d0439980013faa0d3e0524e0992229, {16'd884, 16'd59915, 16'd25643, 16'd29164, 16'd59210, 16'd2918, 16'd44095, 16'd14142, 16'd13434, 16'd58622, 16'd22090, 16'd2135, 16'd46830, 16'd613, 16'd60410, 16'd36360, 16'd35158, 16'd61851, 16'd33527, 16'd17600, 16'd56271, 16'd39412, 16'd64700, 16'd10719, 16'd30991, 16'd22386});
	test_expansion(128'hcef3519197da84685a87b8500200d8c1, {16'd37388, 16'd664, 16'd65228, 16'd34660, 16'd40147, 16'd8038, 16'd28872, 16'd55603, 16'd36989, 16'd45010, 16'd64566, 16'd62585, 16'd55528, 16'd6082, 16'd63871, 16'd42243, 16'd41139, 16'd18522, 16'd60810, 16'd64947, 16'd56093, 16'd4962, 16'd9055, 16'd42977, 16'd54772, 16'd21212});
	test_expansion(128'ha595ffb1e2a71c94a5207a8e51844d5d, {16'd20693, 16'd6400, 16'd39979, 16'd30560, 16'd30676, 16'd27643, 16'd53758, 16'd51394, 16'd22692, 16'd34812, 16'd41546, 16'd40661, 16'd8493, 16'd24082, 16'd9266, 16'd43420, 16'd18377, 16'd38376, 16'd43031, 16'd44105, 16'd4298, 16'd25934, 16'd36321, 16'd65158, 16'd48196, 16'd24472});
	test_expansion(128'h4a1eeefc489d85c1041611c73d1c901d, {16'd43845, 16'd27783, 16'd1653, 16'd35158, 16'd47117, 16'd31129, 16'd30302, 16'd44476, 16'd28614, 16'd27288, 16'd51355, 16'd18339, 16'd64706, 16'd36570, 16'd39268, 16'd35477, 16'd675, 16'd43183, 16'd64462, 16'd65298, 16'd35515, 16'd4738, 16'd63619, 16'd43099, 16'd9505, 16'd37942});
	test_expansion(128'h9efb444b59186ca79d09b9189d198b01, {16'd13687, 16'd43032, 16'd6768, 16'd52930, 16'd16890, 16'd36516, 16'd59652, 16'd6499, 16'd8090, 16'd63280, 16'd59523, 16'd22900, 16'd10357, 16'd51704, 16'd23879, 16'd32656, 16'd63814, 16'd47749, 16'd23698, 16'd58873, 16'd27920, 16'd53857, 16'd8007, 16'd8739, 16'd58053, 16'd10466});
	test_expansion(128'h820be099e67a7a839b75a5a8847ab9ed, {16'd22915, 16'd18978, 16'd39828, 16'd19993, 16'd26264, 16'd28437, 16'd20274, 16'd11038, 16'd1608, 16'd31200, 16'd46164, 16'd4665, 16'd19639, 16'd53649, 16'd12033, 16'd25428, 16'd8067, 16'd39177, 16'd10268, 16'd14607, 16'd3770, 16'd48211, 16'd39791, 16'd17498, 16'd48481, 16'd25455});
	test_expansion(128'h1058d2368edb6695adcb879dc16eaac9, {16'd46790, 16'd54339, 16'd34654, 16'd52048, 16'd59401, 16'd11614, 16'd54485, 16'd50410, 16'd42017, 16'd22555, 16'd45280, 16'd40839, 16'd60209, 16'd35546, 16'd9400, 16'd1533, 16'd63526, 16'd31506, 16'd30146, 16'd32440, 16'd48025, 16'd28083, 16'd59853, 16'd33372, 16'd64111, 16'd45356});
	test_expansion(128'hd5943f62c47e785a54de3b34bda13d11, {16'd8019, 16'd5993, 16'd22954, 16'd61353, 16'd44397, 16'd7727, 16'd26732, 16'd27852, 16'd56397, 16'd44671, 16'd50548, 16'd42659, 16'd38908, 16'd520, 16'd14799, 16'd11095, 16'd32743, 16'd22213, 16'd33720, 16'd13137, 16'd40242, 16'd26134, 16'd47249, 16'd22821, 16'd31757, 16'd36613});
	test_expansion(128'h18959cc06f62f483ef7267de5a36f5ff, {16'd62339, 16'd16604, 16'd58786, 16'd63380, 16'd55816, 16'd55040, 16'd5251, 16'd20526, 16'd59786, 16'd57864, 16'd1102, 16'd17076, 16'd64333, 16'd36847, 16'd45665, 16'd43355, 16'd20824, 16'd25287, 16'd30230, 16'd51624, 16'd13507, 16'd37061, 16'd27698, 16'd54041, 16'd17150, 16'd65282});
	test_expansion(128'h5807b546c3353fd2ce2e4af0926eb767, {16'd4818, 16'd56504, 16'd8522, 16'd46532, 16'd59504, 16'd64801, 16'd40626, 16'd8345, 16'd49638, 16'd6661, 16'd898, 16'd62282, 16'd1914, 16'd38850, 16'd4340, 16'd48577, 16'd15980, 16'd10274, 16'd43470, 16'd37758, 16'd43601, 16'd55578, 16'd50067, 16'd2457, 16'd49585, 16'd29463});
	test_expansion(128'h6f9e6910b7f2cc84a6c034715dc5e4c9, {16'd52551, 16'd8204, 16'd8355, 16'd57382, 16'd34693, 16'd11004, 16'd506, 16'd15641, 16'd3966, 16'd50721, 16'd15566, 16'd3339, 16'd43313, 16'd58469, 16'd41464, 16'd17451, 16'd19291, 16'd20829, 16'd34610, 16'd5063, 16'd20370, 16'd36932, 16'd10749, 16'd56442, 16'd52523, 16'd1406});
	test_expansion(128'hd380eaa91daffe8880934e67f2d937ce, {16'd5165, 16'd26110, 16'd21609, 16'd34459, 16'd2691, 16'd59390, 16'd61218, 16'd51428, 16'd17577, 16'd54491, 16'd42941, 16'd45321, 16'd42992, 16'd31976, 16'd3071, 16'd9637, 16'd5102, 16'd63618, 16'd25632, 16'd25644, 16'd36972, 16'd894, 16'd59307, 16'd45108, 16'd48846, 16'd18707});
	test_expansion(128'h0221c332b99721e2623b21a9821d0cf7, {16'd9840, 16'd44225, 16'd51117, 16'd39749, 16'd34371, 16'd15958, 16'd1675, 16'd46207, 16'd31783, 16'd3696, 16'd37370, 16'd20181, 16'd46644, 16'd31046, 16'd35786, 16'd43980, 16'd55059, 16'd64327, 16'd21275, 16'd55595, 16'd38420, 16'd42352, 16'd42160, 16'd47451, 16'd33101, 16'd47071});
	test_expansion(128'hb59144dbb590eec09c0bf757c17c2f7e, {16'd49943, 16'd40940, 16'd26091, 16'd9689, 16'd51592, 16'd46596, 16'd7515, 16'd21527, 16'd45547, 16'd10168, 16'd56326, 16'd64342, 16'd62268, 16'd63951, 16'd58709, 16'd43521, 16'd40300, 16'd16472, 16'd36591, 16'd55946, 16'd40049, 16'd41142, 16'd55543, 16'd14245, 16'd37699, 16'd57937});
	test_expansion(128'h9ad46e666b9f07b1baabf6c1654da9c5, {16'd2019, 16'd5470, 16'd6445, 16'd19774, 16'd26508, 16'd59581, 16'd45160, 16'd2836, 16'd59025, 16'd56966, 16'd20055, 16'd2920, 16'd51724, 16'd44627, 16'd28872, 16'd34714, 16'd50895, 16'd734, 16'd45089, 16'd42298, 16'd19145, 16'd62233, 16'd43073, 16'd53334, 16'd59089, 16'd58741});
	test_expansion(128'h51bd3487a924b4c9df7551f0dc616a72, {16'd37117, 16'd7541, 16'd6266, 16'd61605, 16'd14979, 16'd61276, 16'd46375, 16'd27198, 16'd57792, 16'd36067, 16'd36751, 16'd41727, 16'd59501, 16'd19962, 16'd29577, 16'd9046, 16'd51026, 16'd15246, 16'd9973, 16'd53613, 16'd29107, 16'd3029, 16'd10672, 16'd41849, 16'd63922, 16'd17999});
	test_expansion(128'h1dcaa4342f4dae659da81a9cc0f39717, {16'd49804, 16'd23105, 16'd58688, 16'd2188, 16'd16577, 16'd698, 16'd18122, 16'd61707, 16'd3222, 16'd46039, 16'd12475, 16'd33377, 16'd44336, 16'd59558, 16'd41907, 16'd31535, 16'd6493, 16'd19503, 16'd40735, 16'd14417, 16'd53345, 16'd16892, 16'd26189, 16'd36721, 16'd41033, 16'd62373});
	test_expansion(128'h7dd19fae942448106f4a164523ace046, {16'd47032, 16'd52697, 16'd17702, 16'd210, 16'd41753, 16'd8946, 16'd53365, 16'd25703, 16'd1202, 16'd49199, 16'd30953, 16'd46336, 16'd26464, 16'd44188, 16'd53209, 16'd62309, 16'd6098, 16'd45458, 16'd5625, 16'd52755, 16'd10728, 16'd2631, 16'd19069, 16'd14621, 16'd41180, 16'd37797});
	test_expansion(128'hd36d2e18dd1a1c91fe239ddf7522b6c3, {16'd17924, 16'd13712, 16'd38770, 16'd5095, 16'd50175, 16'd32123, 16'd1005, 16'd26123, 16'd18022, 16'd8483, 16'd62863, 16'd48191, 16'd24153, 16'd10655, 16'd27850, 16'd54651, 16'd27997, 16'd37554, 16'd62134, 16'd43717, 16'd5277, 16'd8010, 16'd41158, 16'd40310, 16'd43942, 16'd54617});
	test_expansion(128'hdde37c00f8d5f511d594905a8d077ea1, {16'd9796, 16'd40764, 16'd2460, 16'd41045, 16'd48853, 16'd31768, 16'd14984, 16'd37636, 16'd28173, 16'd14155, 16'd524, 16'd58586, 16'd60093, 16'd47911, 16'd27975, 16'd38710, 16'd27562, 16'd51773, 16'd28866, 16'd3935, 16'd21088, 16'd46950, 16'd51895, 16'd56596, 16'd36412, 16'd2926});
	test_expansion(128'hf0578ea2f024cf8b13886012b2f2efc4, {16'd9671, 16'd29837, 16'd17456, 16'd64083, 16'd40081, 16'd34387, 16'd45183, 16'd29961, 16'd2297, 16'd33717, 16'd17341, 16'd31619, 16'd11961, 16'd17539, 16'd22225, 16'd35326, 16'd56212, 16'd38211, 16'd16297, 16'd19040, 16'd29816, 16'd36762, 16'd13532, 16'd39752, 16'd54653, 16'd5237});
	test_expansion(128'h89c0a52bcfda88cd2dc7c9ca23d47cb6, {16'd55715, 16'd24860, 16'd64900, 16'd25023, 16'd32035, 16'd38484, 16'd56740, 16'd28920, 16'd12567, 16'd54096, 16'd5045, 16'd57249, 16'd55863, 16'd13816, 16'd52998, 16'd56191, 16'd35480, 16'd15713, 16'd6666, 16'd49606, 16'd26407, 16'd57166, 16'd63367, 16'd37925, 16'd48648, 16'd40952});
	test_expansion(128'h4cc9a3304d62350d01786ffbb267bf04, {16'd51714, 16'd44682, 16'd22692, 16'd3129, 16'd339, 16'd12602, 16'd35904, 16'd53441, 16'd56365, 16'd65462, 16'd55434, 16'd63022, 16'd55006, 16'd43542, 16'd42034, 16'd35966, 16'd20784, 16'd10807, 16'd5716, 16'd35615, 16'd50349, 16'd17590, 16'd24754, 16'd34375, 16'd38661, 16'd2010});
	test_expansion(128'h4ba1e80aec87e4c0f7c9d7b50f618c0d, {16'd12665, 16'd24731, 16'd12588, 16'd45738, 16'd38686, 16'd5657, 16'd15036, 16'd62299, 16'd1215, 16'd20296, 16'd6967, 16'd46396, 16'd41731, 16'd16532, 16'd24175, 16'd34940, 16'd40403, 16'd20336, 16'd4418, 16'd45829, 16'd41697, 16'd45696, 16'd53482, 16'd48828, 16'd15181, 16'd8484});
	test_expansion(128'ha8f3ba3a9d713ea31e728e570d85891c, {16'd62650, 16'd59994, 16'd2089, 16'd740, 16'd948, 16'd31112, 16'd52773, 16'd61294, 16'd16356, 16'd52215, 16'd31209, 16'd8875, 16'd9941, 16'd63614, 16'd8022, 16'd1905, 16'd8306, 16'd46151, 16'd29689, 16'd24625, 16'd25957, 16'd44027, 16'd13852, 16'd63029, 16'd30910, 16'd56752});
	test_expansion(128'h8f13e619605e02379a284e770bfdb9fc, {16'd62831, 16'd23893, 16'd10725, 16'd14596, 16'd23592, 16'd391, 16'd33872, 16'd2019, 16'd19806, 16'd31881, 16'd47357, 16'd45703, 16'd11038, 16'd20049, 16'd2286, 16'd7519, 16'd5047, 16'd58991, 16'd34510, 16'd64855, 16'd6768, 16'd56953, 16'd29131, 16'd32256, 16'd35851, 16'd20139});
	test_expansion(128'ha98f2b7fdc9c4a39145463d8bf03a70b, {16'd54996, 16'd48133, 16'd54070, 16'd33674, 16'd60392, 16'd57178, 16'd2985, 16'd1663, 16'd29063, 16'd34451, 16'd26203, 16'd36804, 16'd26463, 16'd22059, 16'd1573, 16'd18729, 16'd49811, 16'd27711, 16'd45417, 16'd26949, 16'd31242, 16'd13794, 16'd62549, 16'd34154, 16'd15285, 16'd43195});
	test_expansion(128'hca9ec8fa3947927ca39220d4d8e20f61, {16'd38679, 16'd55645, 16'd49809, 16'd44331, 16'd33834, 16'd26885, 16'd39254, 16'd19503, 16'd55817, 16'd37508, 16'd61702, 16'd42469, 16'd64689, 16'd301, 16'd27112, 16'd13615, 16'd15308, 16'd44524, 16'd11370, 16'd43323, 16'd44738, 16'd59444, 16'd26063, 16'd5252, 16'd11035, 16'd64097});
	test_expansion(128'h5b9c0aec7fd41293a58159ae501aee49, {16'd26063, 16'd15121, 16'd33866, 16'd26000, 16'd44976, 16'd56547, 16'd20949, 16'd45480, 16'd26120, 16'd52159, 16'd9150, 16'd65377, 16'd16118, 16'd9436, 16'd1426, 16'd6864, 16'd55631, 16'd13177, 16'd18462, 16'd58261, 16'd1921, 16'd45408, 16'd24781, 16'd46437, 16'd31519, 16'd8770});
	test_expansion(128'h50b4410c2a85b36632a0c15465915d99, {16'd18949, 16'd44728, 16'd10658, 16'd42714, 16'd47972, 16'd15839, 16'd62568, 16'd24816, 16'd35755, 16'd63963, 16'd23021, 16'd49658, 16'd18468, 16'd48428, 16'd6474, 16'd34230, 16'd56976, 16'd41778, 16'd14631, 16'd42007, 16'd19650, 16'd21799, 16'd33624, 16'd38429, 16'd15256, 16'd34330});
	test_expansion(128'hd4be4a750928dfa40d2b45bf1d7e907a, {16'd26118, 16'd44848, 16'd9690, 16'd27248, 16'd16455, 16'd33772, 16'd64772, 16'd8406, 16'd29103, 16'd60556, 16'd16386, 16'd48492, 16'd50330, 16'd49343, 16'd65296, 16'd30517, 16'd41890, 16'd19134, 16'd16488, 16'd19782, 16'd18777, 16'd8054, 16'd65004, 16'd26422, 16'd50869, 16'd8914});
	test_expansion(128'h252fcb0e122597302b113fea94b83c0c, {16'd29724, 16'd17152, 16'd22482, 16'd4231, 16'd117, 16'd32946, 16'd26112, 16'd8506, 16'd16574, 16'd20390, 16'd5, 16'd9486, 16'd9420, 16'd23688, 16'd57334, 16'd63638, 16'd25164, 16'd23004, 16'd63105, 16'd2255, 16'd6220, 16'd43184, 16'd56830, 16'd51751, 16'd62300, 16'd30343});
	test_expansion(128'h59c4eb97f42caf67bc0c425aa78eaeb2, {16'd9350, 16'd50368, 16'd34591, 16'd19557, 16'd58856, 16'd64662, 16'd49064, 16'd47826, 16'd64486, 16'd42618, 16'd56699, 16'd24307, 16'd43439, 16'd50237, 16'd13845, 16'd64444, 16'd39181, 16'd46621, 16'd4559, 16'd46633, 16'd56909, 16'd40537, 16'd50001, 16'd59759, 16'd51546, 16'd45105});
	test_expansion(128'h088dc1e6a316d5f03b3a88b35780b60c, {16'd62348, 16'd41457, 16'd11478, 16'd1149, 16'd33822, 16'd57514, 16'd23416, 16'd31961, 16'd47963, 16'd44519, 16'd31526, 16'd42384, 16'd38122, 16'd11620, 16'd59669, 16'd15661, 16'd3857, 16'd57552, 16'd56652, 16'd35905, 16'd10528, 16'd54112, 16'd32788, 16'd20402, 16'd815, 16'd44331});
	test_expansion(128'hbc04c2fbac96a1136f864327c26a597b, {16'd22424, 16'd11317, 16'd20069, 16'd25043, 16'd10038, 16'd54464, 16'd32542, 16'd9324, 16'd23480, 16'd36136, 16'd954, 16'd61727, 16'd17415, 16'd36647, 16'd51921, 16'd47654, 16'd518, 16'd36789, 16'd46154, 16'd10348, 16'd27883, 16'd41835, 16'd38347, 16'd27970, 16'd6649, 16'd55896});
	test_expansion(128'hfdf7fdb12ee2273d5c75c752e602635a, {16'd5501, 16'd16118, 16'd27102, 16'd37812, 16'd7123, 16'd13771, 16'd42164, 16'd46829, 16'd41630, 16'd42141, 16'd30449, 16'd48467, 16'd27324, 16'd25595, 16'd42023, 16'd62632, 16'd6906, 16'd23459, 16'd25255, 16'd34132, 16'd4736, 16'd13139, 16'd52704, 16'd8855, 16'd33886, 16'd21413});
	test_expansion(128'h0309d5cfb6cd11f03904fd2e5866c951, {16'd50498, 16'd24460, 16'd10491, 16'd33582, 16'd23229, 16'd29218, 16'd30186, 16'd9163, 16'd57941, 16'd13254, 16'd593, 16'd23710, 16'd31767, 16'd36316, 16'd51903, 16'd52872, 16'd55390, 16'd27303, 16'd35753, 16'd50589, 16'd28915, 16'd60797, 16'd61315, 16'd693, 16'd32206, 16'd16287});
	test_expansion(128'hef0f29ca997645bb9edc3df9f74ade93, {16'd29159, 16'd13796, 16'd1113, 16'd15245, 16'd12914, 16'd13078, 16'd40380, 16'd61834, 16'd5598, 16'd54210, 16'd32106, 16'd21653, 16'd41545, 16'd10306, 16'd48193, 16'd5217, 16'd1897, 16'd13172, 16'd29187, 16'd56149, 16'd8088, 16'd7084, 16'd54062, 16'd57984, 16'd56503, 16'd61540});
	test_expansion(128'h02382bc39b2a2e7445c028fd501dce56, {16'd62438, 16'd14828, 16'd32821, 16'd11151, 16'd48657, 16'd23115, 16'd21664, 16'd20358, 16'd316, 16'd38260, 16'd19901, 16'd2802, 16'd46200, 16'd21856, 16'd6900, 16'd54240, 16'd16909, 16'd25871, 16'd29946, 16'd3780, 16'd3158, 16'd21397, 16'd8670, 16'd54773, 16'd49823, 16'd8486});
	test_expansion(128'h5bdef338fb0231330b002af8d5767340, {16'd6055, 16'd52551, 16'd59507, 16'd29600, 16'd60154, 16'd22455, 16'd54236, 16'd39801, 16'd60642, 16'd46133, 16'd21738, 16'd56909, 16'd57264, 16'd47189, 16'd40348, 16'd58543, 16'd52222, 16'd61769, 16'd30741, 16'd31877, 16'd47801, 16'd29999, 16'd31698, 16'd52831, 16'd61465, 16'd10668});
	test_expansion(128'h64c4fbb4e4c3e5c326f92603608712e8, {16'd25446, 16'd55282, 16'd44476, 16'd56270, 16'd28139, 16'd61584, 16'd8648, 16'd33591, 16'd45311, 16'd57586, 16'd35823, 16'd13414, 16'd12505, 16'd64969, 16'd61032, 16'd11877, 16'd33568, 16'd11471, 16'd57814, 16'd31052, 16'd38401, 16'd15974, 16'd25979, 16'd2300, 16'd794, 16'd57882});
	test_expansion(128'h24e625f3a5cc58e8a783371560267ffb, {16'd30774, 16'd21435, 16'd61023, 16'd59818, 16'd32266, 16'd2410, 16'd54511, 16'd60049, 16'd39066, 16'd30411, 16'd46284, 16'd32659, 16'd57188, 16'd10272, 16'd14917, 16'd13616, 16'd38683, 16'd36422, 16'd34284, 16'd44815, 16'd12918, 16'd1256, 16'd49323, 16'd3695, 16'd46565, 16'd22763});
	test_expansion(128'h6425b56733cd395e45eab69be44b4c27, {16'd40529, 16'd29835, 16'd4160, 16'd4837, 16'd20746, 16'd24749, 16'd24502, 16'd51551, 16'd4469, 16'd38828, 16'd57515, 16'd15989, 16'd14743, 16'd20113, 16'd40788, 16'd24655, 16'd4700, 16'd649, 16'd5513, 16'd7499, 16'd64066, 16'd57907, 16'd3916, 16'd33638, 16'd34855, 16'd41656});
	test_expansion(128'h7cd6b417601edb060c70fc0847b4cd84, {16'd39649, 16'd39071, 16'd31786, 16'd14453, 16'd46804, 16'd41668, 16'd58485, 16'd39074, 16'd55085, 16'd32221, 16'd48071, 16'd13590, 16'd12016, 16'd34041, 16'd6003, 16'd51957, 16'd24637, 16'd30350, 16'd47738, 16'd1751, 16'd43484, 16'd19312, 16'd23479, 16'd37058, 16'd12857, 16'd46903});
	test_expansion(128'hf64dbfd92dec8b2cebe31bb50221870d, {16'd21872, 16'd41150, 16'd24421, 16'd23624, 16'd43828, 16'd51959, 16'd48749, 16'd17534, 16'd19849, 16'd42474, 16'd4691, 16'd13590, 16'd63594, 16'd34758, 16'd57385, 16'd60654, 16'd12602, 16'd37328, 16'd16765, 16'd54278, 16'd46565, 16'd35136, 16'd55439, 16'd35, 16'd61300, 16'd23015});
	test_expansion(128'h108bb42eee6075f0e476d4425ade8430, {16'd31191, 16'd58328, 16'd57197, 16'd34008, 16'd57533, 16'd17415, 16'd5221, 16'd43216, 16'd8494, 16'd25587, 16'd56621, 16'd13905, 16'd27719, 16'd22405, 16'd61100, 16'd28290, 16'd58498, 16'd46459, 16'd61855, 16'd62988, 16'd33223, 16'd64105, 16'd25793, 16'd4274, 16'd5228, 16'd32964});
	test_expansion(128'h91cc1b2977f924e274104769cf61a46d, {16'd14545, 16'd16690, 16'd33625, 16'd12794, 16'd6974, 16'd53039, 16'd61850, 16'd15985, 16'd27007, 16'd52387, 16'd25941, 16'd25629, 16'd54042, 16'd10929, 16'd47910, 16'd9391, 16'd27689, 16'd56088, 16'd47184, 16'd9071, 16'd19823, 16'd57517, 16'd5327, 16'd54444, 16'd17178, 16'd6160});
	test_expansion(128'h94c23599a6a68ef814163b16b93bd630, {16'd39684, 16'd7689, 16'd24982, 16'd50444, 16'd31023, 16'd8661, 16'd1402, 16'd24464, 16'd28216, 16'd41085, 16'd64182, 16'd64307, 16'd56674, 16'd29812, 16'd48137, 16'd39925, 16'd49535, 16'd33401, 16'd852, 16'd20170, 16'd15557, 16'd64050, 16'd2684, 16'd4931, 16'd25400, 16'd59752});
	test_expansion(128'hb2dcb01cefde07d9928af2523169b394, {16'd6814, 16'd4114, 16'd3254, 16'd63667, 16'd36787, 16'd2320, 16'd42116, 16'd9986, 16'd16224, 16'd62386, 16'd44712, 16'd5548, 16'd49981, 16'd17927, 16'd51087, 16'd4297, 16'd14182, 16'd10301, 16'd13800, 16'd64938, 16'd23815, 16'd58312, 16'd28439, 16'd14820, 16'd8772, 16'd30570});
	test_expansion(128'h8af7f40716338362755afe3ad2bb33f0, {16'd29588, 16'd2575, 16'd27615, 16'd8632, 16'd23939, 16'd1741, 16'd45213, 16'd33941, 16'd50689, 16'd16858, 16'd62496, 16'd44855, 16'd60915, 16'd24809, 16'd4794, 16'd52310, 16'd43581, 16'd11192, 16'd19044, 16'd17802, 16'd43744, 16'd14233, 16'd9502, 16'd17704, 16'd28467, 16'd49416});
	test_expansion(128'h4cd709e9573d6cc424a83b6c215558cb, {16'd42038, 16'd630, 16'd1223, 16'd13212, 16'd49910, 16'd48600, 16'd5340, 16'd40307, 16'd8604, 16'd16831, 16'd48604, 16'd30815, 16'd24566, 16'd7723, 16'd22677, 16'd37859, 16'd8004, 16'd57449, 16'd28863, 16'd62194, 16'd64113, 16'd52119, 16'd35197, 16'd10389, 16'd55344, 16'd17376});
	test_expansion(128'hadadf8c1ff3cc20933550c012cd0d294, {16'd39046, 16'd12657, 16'd51510, 16'd23134, 16'd44468, 16'd27045, 16'd13906, 16'd51104, 16'd63140, 16'd19294, 16'd27762, 16'd9476, 16'd41850, 16'd33822, 16'd26677, 16'd60698, 16'd42244, 16'd22656, 16'd21236, 16'd18085, 16'd58989, 16'd45773, 16'd48624, 16'd59374, 16'd28927, 16'd35939});
	test_expansion(128'hf060cdfa394f2a0fa921fe2e1a7e6096, {16'd50694, 16'd64451, 16'd680, 16'd27430, 16'd47020, 16'd3570, 16'd35588, 16'd15920, 16'd38835, 16'd16454, 16'd16499, 16'd45079, 16'd35384, 16'd42940, 16'd52805, 16'd3012, 16'd27138, 16'd60818, 16'd7904, 16'd58173, 16'd57353, 16'd45477, 16'd51232, 16'd15978, 16'd63282, 16'd38314});
	test_expansion(128'h53c998ad9169dc38b171514c18b6cfba, {16'd13828, 16'd57821, 16'd55747, 16'd22717, 16'd23172, 16'd61508, 16'd26928, 16'd10126, 16'd48839, 16'd51769, 16'd33716, 16'd44583, 16'd8883, 16'd7613, 16'd534, 16'd29089, 16'd21104, 16'd33534, 16'd53225, 16'd34276, 16'd58307, 16'd36974, 16'd32239, 16'd25944, 16'd53788, 16'd28492});
	test_expansion(128'h6cfdb910e38b19c13a5d2092ceb4bffe, {16'd29444, 16'd27496, 16'd40284, 16'd14506, 16'd49963, 16'd27288, 16'd53731, 16'd40187, 16'd47081, 16'd46902, 16'd61185, 16'd54889, 16'd6541, 16'd29832, 16'd1788, 16'd34104, 16'd37155, 16'd46944, 16'd29150, 16'd1054, 16'd55452, 16'd59547, 16'd21428, 16'd32044, 16'd24067, 16'd39322});
	test_expansion(128'h5ce4ede741d933663175b6991e4081a2, {16'd53444, 16'd34735, 16'd22017, 16'd32025, 16'd57974, 16'd63404, 16'd42711, 16'd19936, 16'd15832, 16'd34910, 16'd39426, 16'd37195, 16'd46893, 16'd59000, 16'd23718, 16'd57015, 16'd4660, 16'd2379, 16'd7790, 16'd21973, 16'd5882, 16'd11737, 16'd14916, 16'd54574, 16'd63025, 16'd27678});
	test_expansion(128'hccfbfafef71ee9f6f67b7679eeb0e75b, {16'd16124, 16'd8671, 16'd28867, 16'd33744, 16'd37550, 16'd577, 16'd55313, 16'd45172, 16'd58924, 16'd34497, 16'd44524, 16'd23682, 16'd38113, 16'd45698, 16'd46375, 16'd38233, 16'd45318, 16'd49457, 16'd64463, 16'd6870, 16'd44511, 16'd58279, 16'd15144, 16'd41077, 16'd12342, 16'd31140});
	test_expansion(128'h42bcd874b307e3bfec4d6299faaaba43, {16'd11158, 16'd60029, 16'd20537, 16'd20353, 16'd34955, 16'd34475, 16'd3632, 16'd27196, 16'd29990, 16'd41968, 16'd2931, 16'd56802, 16'd40798, 16'd921, 16'd51048, 16'd63540, 16'd21118, 16'd31782, 16'd21051, 16'd38709, 16'd51131, 16'd54315, 16'd39437, 16'd64485, 16'd5310, 16'd55052});
	test_expansion(128'he0437c1f47400715c8fcb92a5d817952, {16'd14870, 16'd10902, 16'd45061, 16'd49257, 16'd21730, 16'd6455, 16'd61449, 16'd61364, 16'd6527, 16'd39628, 16'd62105, 16'd56402, 16'd6495, 16'd34530, 16'd20896, 16'd22022, 16'd24080, 16'd15553, 16'd32397, 16'd12480, 16'd61707, 16'd26508, 16'd58186, 16'd30684, 16'd21792, 16'd13007});
	test_expansion(128'h984a95b8decf8b514bc9c835330b93eb, {16'd23063, 16'd61844, 16'd640, 16'd30911, 16'd2972, 16'd28774, 16'd35925, 16'd61175, 16'd19015, 16'd40279, 16'd54409, 16'd28376, 16'd7093, 16'd38557, 16'd48736, 16'd29819, 16'd18341, 16'd24157, 16'd32073, 16'd37507, 16'd55612, 16'd23992, 16'd51631, 16'd56802, 16'd63698, 16'd52668});
	test_expansion(128'hd5645802a5119917353bb044465d6521, {16'd22940, 16'd64079, 16'd31417, 16'd23739, 16'd56760, 16'd41181, 16'd29331, 16'd10421, 16'd8841, 16'd10813, 16'd52337, 16'd40544, 16'd28606, 16'd64053, 16'd27021, 16'd22094, 16'd55226, 16'd21339, 16'd40293, 16'd21572, 16'd10460, 16'd22639, 16'd45177, 16'd11295, 16'd12587, 16'd55918});
	test_expansion(128'h5bc307dce6d569495da8d1b844341d32, {16'd25051, 16'd45929, 16'd47852, 16'd6081, 16'd48504, 16'd49641, 16'd14144, 16'd12280, 16'd14616, 16'd21491, 16'd58194, 16'd33579, 16'd39350, 16'd7017, 16'd42491, 16'd29661, 16'd41886, 16'd60482, 16'd55970, 16'd53114, 16'd60525, 16'd5590, 16'd52254, 16'd52578, 16'd20490, 16'd39360});
	test_expansion(128'h3b318880605c40bec324d0b9412a9ed4, {16'd61347, 16'd35172, 16'd1194, 16'd60543, 16'd8407, 16'd52135, 16'd2224, 16'd44712, 16'd58741, 16'd37680, 16'd15863, 16'd36981, 16'd23273, 16'd46638, 16'd40190, 16'd3756, 16'd27032, 16'd17951, 16'd40282, 16'd23146, 16'd59237, 16'd39262, 16'd7420, 16'd59868, 16'd35559, 16'd45958});
	test_expansion(128'h88f99ddc1276a78d539a8ba10329437f, {16'd41442, 16'd34600, 16'd40071, 16'd31513, 16'd35998, 16'd23150, 16'd58010, 16'd42536, 16'd26107, 16'd12449, 16'd48161, 16'd61596, 16'd21017, 16'd45064, 16'd44521, 16'd59981, 16'd34509, 16'd16395, 16'd5137, 16'd56804, 16'd3900, 16'd1812, 16'd782, 16'd17642, 16'd10167, 16'd8432});
	test_expansion(128'hf20bbff61a030113e90917285c93d446, {16'd21330, 16'd33780, 16'd2476, 16'd22853, 16'd10502, 16'd63809, 16'd9472, 16'd11691, 16'd27538, 16'd6932, 16'd31643, 16'd8055, 16'd22402, 16'd31931, 16'd3919, 16'd31899, 16'd25446, 16'd41720, 16'd37130, 16'd59421, 16'd64555, 16'd13122, 16'd28798, 16'd61718, 16'd40213, 16'd51619});
	test_expansion(128'ha2fc0f14c3bc0c7c678805f532a0df7e, {16'd7960, 16'd53659, 16'd35282, 16'd27047, 16'd7451, 16'd32916, 16'd17370, 16'd29072, 16'd33172, 16'd1517, 16'd13133, 16'd12631, 16'd15374, 16'd53694, 16'd16715, 16'd52167, 16'd13694, 16'd58630, 16'd12587, 16'd7661, 16'd21343, 16'd40909, 16'd33244, 16'd15275, 16'd51394, 16'd7045});
	test_expansion(128'h67c33d7d5289398cedba95a9b129b888, {16'd23115, 16'd24349, 16'd59073, 16'd45426, 16'd6696, 16'd65503, 16'd16906, 16'd1800, 16'd8458, 16'd23990, 16'd10449, 16'd44724, 16'd16168, 16'd732, 16'd21037, 16'd20851, 16'd10966, 16'd36288, 16'd55369, 16'd56327, 16'd34009, 16'd38302, 16'd59911, 16'd56208, 16'd36322, 16'd30470});
	test_expansion(128'he04cb2508bc80383abde68708b78c48e, {16'd16253, 16'd4537, 16'd50828, 16'd13744, 16'd19748, 16'd15978, 16'd14569, 16'd57694, 16'd4172, 16'd63842, 16'd37843, 16'd35316, 16'd20865, 16'd54073, 16'd14160, 16'd54584, 16'd44247, 16'd22224, 16'd30304, 16'd54638, 16'd35980, 16'd18467, 16'd42416, 16'd17878, 16'd62031, 16'd30494});
	test_expansion(128'ha803dfd061586e35fa58d386f5fe8c13, {16'd63723, 16'd22220, 16'd10702, 16'd26910, 16'd56730, 16'd3393, 16'd25010, 16'd2760, 16'd21395, 16'd48301, 16'd22597, 16'd44951, 16'd5647, 16'd17623, 16'd43360, 16'd15998, 16'd59734, 16'd39117, 16'd46546, 16'd19742, 16'd48755, 16'd60329, 16'd46424, 16'd41568, 16'd30276, 16'd20856});
	test_expansion(128'hd6a2903ec84ba02d6a46003b0c7b4ca9, {16'd9122, 16'd63367, 16'd35146, 16'd63215, 16'd19866, 16'd54007, 16'd63402, 16'd53, 16'd22787, 16'd59373, 16'd20355, 16'd47455, 16'd11121, 16'd44314, 16'd31625, 16'd42608, 16'd42122, 16'd16769, 16'd37338, 16'd1737, 16'd7485, 16'd34304, 16'd25422, 16'd20158, 16'd26371, 16'd52887});
	test_expansion(128'h0776031ce89a48c1478f3986721b3341, {16'd11300, 16'd15317, 16'd63520, 16'd6708, 16'd56646, 16'd40031, 16'd52209, 16'd24544, 16'd9370, 16'd52173, 16'd4928, 16'd59430, 16'd51937, 16'd46529, 16'd4842, 16'd28333, 16'd6259, 16'd19140, 16'd32645, 16'd62676, 16'd47633, 16'd24083, 16'd58821, 16'd34022, 16'd54149, 16'd7146});
	test_expansion(128'hbcbe56e4498ed9c0d7f28232accf1b51, {16'd45200, 16'd65400, 16'd24581, 16'd11793, 16'd45411, 16'd38876, 16'd32984, 16'd30934, 16'd6014, 16'd24534, 16'd20133, 16'd29222, 16'd21037, 16'd28996, 16'd5598, 16'd8760, 16'd9950, 16'd55912, 16'd31229, 16'd28690, 16'd19053, 16'd27358, 16'd64683, 16'd40395, 16'd31364, 16'd41996});
	test_expansion(128'hf95bb3cd86279f8697ae4081a74fc5f3, {16'd7661, 16'd51753, 16'd61545, 16'd60955, 16'd18992, 16'd65299, 16'd63646, 16'd23312, 16'd37967, 16'd41960, 16'd39593, 16'd55856, 16'd62974, 16'd40750, 16'd13989, 16'd62265, 16'd18986, 16'd29144, 16'd10610, 16'd40350, 16'd60714, 16'd22111, 16'd6762, 16'd33181, 16'd46881, 16'd60299});
	test_expansion(128'h07bc216f2f3427616ac6335f51b61611, {16'd17686, 16'd57768, 16'd45370, 16'd30740, 16'd15637, 16'd9279, 16'd15844, 16'd32288, 16'd35251, 16'd18660, 16'd9706, 16'd35568, 16'd12962, 16'd24502, 16'd20794, 16'd6233, 16'd11196, 16'd60037, 16'd1469, 16'd14777, 16'd2355, 16'd53770, 16'd23047, 16'd47195, 16'd15536, 16'd24952});
	test_expansion(128'h65462c8431af72955ce8a72870e42f46, {16'd20078, 16'd39773, 16'd50308, 16'd37080, 16'd56876, 16'd34061, 16'd64951, 16'd50872, 16'd28882, 16'd36315, 16'd31573, 16'd30804, 16'd60203, 16'd61467, 16'd2193, 16'd11331, 16'd29142, 16'd40964, 16'd15259, 16'd7852, 16'd32158, 16'd16177, 16'd53276, 16'd54777, 16'd64464, 16'd11412});
	test_expansion(128'h161eb982988e2ad6ec92957d170a4ecf, {16'd13309, 16'd63868, 16'd33230, 16'd3641, 16'd56919, 16'd10166, 16'd16762, 16'd48240, 16'd61103, 16'd33598, 16'd6088, 16'd26074, 16'd47628, 16'd11761, 16'd17328, 16'd1277, 16'd19855, 16'd27522, 16'd43313, 16'd40305, 16'd31881, 16'd25176, 16'd54158, 16'd37221, 16'd65406, 16'd12409});
	test_expansion(128'hda693297dd6662dd5b00ee0820cb2875, {16'd21934, 16'd53313, 16'd29919, 16'd21322, 16'd30399, 16'd44229, 16'd53632, 16'd15327, 16'd16865, 16'd59094, 16'd57193, 16'd28170, 16'd57722, 16'd60587, 16'd28480, 16'd40329, 16'd12115, 16'd63517, 16'd55208, 16'd25680, 16'd26592, 16'd7649, 16'd10901, 16'd61985, 16'd60092, 16'd9786});
	test_expansion(128'ha3e7bfbcacd90f0658f042adb6e75cbf, {16'd31700, 16'd39963, 16'd35564, 16'd58152, 16'd59826, 16'd21230, 16'd52518, 16'd1417, 16'd45160, 16'd31073, 16'd44967, 16'd3284, 16'd53153, 16'd20246, 16'd22962, 16'd30995, 16'd7177, 16'd36687, 16'd2303, 16'd49386, 16'd21387, 16'd42731, 16'd44382, 16'd6729, 16'd59151, 16'd10047});
	test_expansion(128'h5425aa12acfb6ede584a972e2f90cbb7, {16'd38799, 16'd16596, 16'd61441, 16'd45944, 16'd21244, 16'd51261, 16'd35857, 16'd3648, 16'd30449, 16'd65478, 16'd33258, 16'd41522, 16'd46184, 16'd35160, 16'd52176, 16'd20947, 16'd3384, 16'd19213, 16'd55340, 16'd7795, 16'd39707, 16'd57036, 16'd19541, 16'd26603, 16'd59128, 16'd42772});
	test_expansion(128'hb0e4834b6b9ed3d80b44342295cf9dd6, {16'd14972, 16'd58838, 16'd580, 16'd21986, 16'd44375, 16'd36705, 16'd58137, 16'd60661, 16'd58594, 16'd52241, 16'd868, 16'd14744, 16'd9757, 16'd56634, 16'd11544, 16'd18760, 16'd53742, 16'd30479, 16'd39086, 16'd31813, 16'd23948, 16'd42056, 16'd18270, 16'd30465, 16'd60283, 16'd11471});
	test_expansion(128'hfe7f3607dfed62182fe12461e2747355, {16'd13494, 16'd27506, 16'd26500, 16'd22603, 16'd52594, 16'd33761, 16'd52987, 16'd7344, 16'd32205, 16'd21979, 16'd25962, 16'd64642, 16'd2223, 16'd23161, 16'd34703, 16'd18772, 16'd4703, 16'd56403, 16'd35368, 16'd40947, 16'd44631, 16'd5216, 16'd38695, 16'd34663, 16'd8174, 16'd20002});
	test_expansion(128'h2d28333259b891d87c8658005b05e1da, {16'd59259, 16'd59247, 16'd59755, 16'd38092, 16'd21733, 16'd2690, 16'd33770, 16'd49594, 16'd56187, 16'd24792, 16'd52134, 16'd21844, 16'd20595, 16'd6467, 16'd52567, 16'd27310, 16'd9859, 16'd52718, 16'd57233, 16'd41055, 16'd48360, 16'd11113, 16'd54130, 16'd46093, 16'd2990, 16'd57549});
	test_expansion(128'hd8a8e09e28e509a38e175d278a01b3bb, {16'd26417, 16'd17929, 16'd41426, 16'd22716, 16'd7085, 16'd56707, 16'd21531, 16'd28099, 16'd41579, 16'd37879, 16'd52766, 16'd50624, 16'd46373, 16'd39629, 16'd58219, 16'd42515, 16'd20247, 16'd45497, 16'd57231, 16'd25642, 16'd12822, 16'd59893, 16'd15275, 16'd7821, 16'd52381, 16'd51586});
	test_expansion(128'hbd0bed0b430027ddcc9f1ca2f35ea122, {16'd5635, 16'd57305, 16'd5725, 16'd28609, 16'd34225, 16'd35460, 16'd19792, 16'd41817, 16'd13570, 16'd46550, 16'd21958, 16'd28390, 16'd50361, 16'd4129, 16'd16755, 16'd62684, 16'd18965, 16'd47715, 16'd1083, 16'd28692, 16'd55614, 16'd56041, 16'd31915, 16'd48222, 16'd30957, 16'd1763});
	test_expansion(128'h2d72e7c42fd1eec7813a3642fd62c45c, {16'd41537, 16'd13846, 16'd58933, 16'd65535, 16'd57423, 16'd64794, 16'd18338, 16'd47613, 16'd40531, 16'd52564, 16'd36738, 16'd47767, 16'd34825, 16'd52726, 16'd5288, 16'd43829, 16'd20194, 16'd23482, 16'd16952, 16'd56981, 16'd47575, 16'd40288, 16'd51851, 16'd16404, 16'd23676, 16'd40876});
	test_expansion(128'h7f80b95d075c47da2d6f2acb281eb3b1, {16'd48139, 16'd53944, 16'd55611, 16'd26703, 16'd60187, 16'd35318, 16'd18237, 16'd31401, 16'd22655, 16'd10661, 16'd1273, 16'd47665, 16'd33724, 16'd24809, 16'd10291, 16'd801, 16'd22888, 16'd24154, 16'd45196, 16'd58638, 16'd9831, 16'd49683, 16'd13087, 16'd30275, 16'd30578, 16'd24170});
	test_expansion(128'h210d707f9996557d73357781204a5c38, {16'd21097, 16'd8105, 16'd17436, 16'd28762, 16'd46370, 16'd35303, 16'd25212, 16'd61898, 16'd41540, 16'd4285, 16'd58654, 16'd5465, 16'd10219, 16'd23199, 16'd50995, 16'd6544, 16'd1072, 16'd60729, 16'd27564, 16'd59647, 16'd19658, 16'd1921, 16'd58424, 16'd6515, 16'd34574, 16'd59263});
	test_expansion(128'hea74b89b67a57297ea0296194bc41b99, {16'd4746, 16'd6836, 16'd28592, 16'd29294, 16'd3223, 16'd32010, 16'd31430, 16'd16696, 16'd59628, 16'd31391, 16'd41633, 16'd24546, 16'd23233, 16'd59558, 16'd27176, 16'd10913, 16'd907, 16'd55706, 16'd21105, 16'd62736, 16'd43496, 16'd45639, 16'd44591, 16'd16231, 16'd63360, 16'd43409});
	test_expansion(128'hc1096d2e34288425ce34c1990e709f06, {16'd20031, 16'd64485, 16'd34274, 16'd38975, 16'd56697, 16'd45475, 16'd10039, 16'd9039, 16'd22708, 16'd61386, 16'd26660, 16'd45973, 16'd54001, 16'd60247, 16'd63518, 16'd48909, 16'd22157, 16'd25499, 16'd41580, 16'd20295, 16'd43119, 16'd9406, 16'd57330, 16'd48602, 16'd62722, 16'd24590});
	test_expansion(128'he4d12e32e51c4447cffc8ac1877e87d4, {16'd38034, 16'd23680, 16'd5183, 16'd56717, 16'd11700, 16'd38833, 16'd37846, 16'd1820, 16'd9387, 16'd36021, 16'd50974, 16'd62477, 16'd721, 16'd61353, 16'd60411, 16'd40792, 16'd10732, 16'd9580, 16'd23393, 16'd55678, 16'd40737, 16'd22064, 16'd56885, 16'd60736, 16'd8619, 16'd2639});
	test_expansion(128'hd446d88ab8bde8edcb952a9264bab979, {16'd53190, 16'd59263, 16'd24306, 16'd5940, 16'd13125, 16'd12736, 16'd52744, 16'd31557, 16'd45176, 16'd17250, 16'd51727, 16'd48115, 16'd24579, 16'd15516, 16'd60322, 16'd30163, 16'd16498, 16'd14298, 16'd42219, 16'd8972, 16'd30224, 16'd24074, 16'd39756, 16'd32264, 16'd52379, 16'd26177});
	test_expansion(128'h7c9997e86a949dcae249b85d88baf00e, {16'd21141, 16'd25899, 16'd59442, 16'd47051, 16'd19824, 16'd13196, 16'd17622, 16'd50853, 16'd30905, 16'd54119, 16'd3780, 16'd39479, 16'd17062, 16'd45210, 16'd11496, 16'd9545, 16'd19412, 16'd7682, 16'd63972, 16'd36133, 16'd38181, 16'd10534, 16'd35362, 16'd51535, 16'd4411, 16'd28503});
	test_expansion(128'h02970be0d6194e2a91910c54c3c78ce3, {16'd8804, 16'd9095, 16'd39135, 16'd45998, 16'd44508, 16'd51998, 16'd29787, 16'd2309, 16'd55646, 16'd30329, 16'd1544, 16'd54243, 16'd4121, 16'd16059, 16'd2112, 16'd43988, 16'd5295, 16'd5850, 16'd43614, 16'd54665, 16'd61616, 16'd16132, 16'd33432, 16'd32324, 16'd44576, 16'd38232});
	test_expansion(128'hf7846aa4b0bf114d1c1379219a6b6a62, {16'd64682, 16'd27689, 16'd105, 16'd316, 16'd9016, 16'd64839, 16'd55154, 16'd45653, 16'd48161, 16'd55483, 16'd23090, 16'd3363, 16'd24941, 16'd64017, 16'd41940, 16'd18911, 16'd10529, 16'd61486, 16'd61269, 16'd42283, 16'd24879, 16'd31746, 16'd53869, 16'd65174, 16'd63057, 16'd47461});
	test_expansion(128'h2b4fec0dff4cfedbec27fb449b5aafa9, {16'd23139, 16'd38022, 16'd43742, 16'd13148, 16'd46245, 16'd4503, 16'd2705, 16'd30536, 16'd41548, 16'd39480, 16'd37109, 16'd38420, 16'd56760, 16'd56320, 16'd42135, 16'd50537, 16'd53923, 16'd30601, 16'd20505, 16'd56055, 16'd20576, 16'd51662, 16'd5296, 16'd11239, 16'd28669, 16'd29594});
	test_expansion(128'h571b464d9f924e255528ef70cbbed5ff, {16'd28611, 16'd29790, 16'd43126, 16'd18788, 16'd11548, 16'd21370, 16'd2577, 16'd18536, 16'd40648, 16'd42999, 16'd52808, 16'd45040, 16'd36720, 16'd4524, 16'd32581, 16'd60214, 16'd58875, 16'd22705, 16'd48957, 16'd38912, 16'd355, 16'd45465, 16'd20314, 16'd28569, 16'd4509, 16'd5250});
	test_expansion(128'h2ba4065d182dbf0b5dc8b0ea415d86e4, {16'd49681, 16'd62449, 16'd47555, 16'd15417, 16'd65093, 16'd37161, 16'd61626, 16'd47214, 16'd52298, 16'd7559, 16'd63008, 16'd62927, 16'd38765, 16'd56680, 16'd43792, 16'd35505, 16'd3166, 16'd51911, 16'd52711, 16'd6348, 16'd4218, 16'd24060, 16'd19773, 16'd5344, 16'd45240, 16'd40468});
	test_expansion(128'h596800ffc8d928dbcbf1b865f84286c3, {16'd4653, 16'd39200, 16'd62070, 16'd30640, 16'd5468, 16'd57534, 16'd55807, 16'd28338, 16'd19090, 16'd30652, 16'd42790, 16'd266, 16'd60402, 16'd58143, 16'd12589, 16'd7773, 16'd31926, 16'd6850, 16'd56877, 16'd57538, 16'd24334, 16'd61023, 16'd61052, 16'd60922, 16'd9206, 16'd14282});
	test_expansion(128'hf36ab3e7cc3c84443aecd6455af41570, {16'd18516, 16'd9777, 16'd35598, 16'd51323, 16'd29940, 16'd3282, 16'd18213, 16'd43364, 16'd37366, 16'd4033, 16'd57572, 16'd1728, 16'd31473, 16'd63782, 16'd32297, 16'd44363, 16'd36838, 16'd63764, 16'd6353, 16'd40449, 16'd39319, 16'd13562, 16'd60979, 16'd10952, 16'd60141, 16'd60355});
	test_expansion(128'h403214ffe7dea4781e29655684279dcf, {16'd26307, 16'd62542, 16'd5989, 16'd31685, 16'd22587, 16'd36430, 16'd29392, 16'd18197, 16'd53401, 16'd50717, 16'd89, 16'd56637, 16'd13012, 16'd63853, 16'd3327, 16'd25431, 16'd21441, 16'd46336, 16'd56026, 16'd33676, 16'd1334, 16'd9874, 16'd50034, 16'd901, 16'd1821, 16'd40693});
	test_expansion(128'hcaf665d5a55700ba5eb28e9a696a6741, {16'd33090, 16'd33157, 16'd50263, 16'd52745, 16'd40745, 16'd7430, 16'd42543, 16'd59351, 16'd65321, 16'd9310, 16'd16042, 16'd55951, 16'd37290, 16'd8453, 16'd1304, 16'd7920, 16'd38083, 16'd4643, 16'd11752, 16'd23397, 16'd46935, 16'd27674, 16'd50566, 16'd25311, 16'd6365, 16'd35274});
	test_expansion(128'hcd5aed8b180febde54fba0fa7e1385cd, {16'd53049, 16'd2855, 16'd32053, 16'd48485, 16'd22442, 16'd39688, 16'd43259, 16'd30093, 16'd58719, 16'd62581, 16'd43177, 16'd44323, 16'd32544, 16'd34619, 16'd16366, 16'd17541, 16'd58626, 16'd36068, 16'd41968, 16'd45168, 16'd13219, 16'd22739, 16'd29769, 16'd21082, 16'd887, 16'd21717});
	test_expansion(128'hf560bfffdafc7db13e8332780e4a5460, {16'd39442, 16'd44029, 16'd60459, 16'd26171, 16'd39595, 16'd65421, 16'd61586, 16'd35054, 16'd27024, 16'd14167, 16'd35280, 16'd30185, 16'd34647, 16'd13184, 16'd59716, 16'd3102, 16'd35731, 16'd29357, 16'd17112, 16'd30474, 16'd30786, 16'd40576, 16'd19405, 16'd3819, 16'd40943, 16'd31841});
	test_expansion(128'h130dd1798cfa3ee70b2a1cc886eb6359, {16'd37790, 16'd52247, 16'd3112, 16'd18, 16'd20109, 16'd43546, 16'd60143, 16'd9806, 16'd15513, 16'd36755, 16'd2419, 16'd24574, 16'd17013, 16'd51564, 16'd32918, 16'd11357, 16'd2574, 16'd13314, 16'd37355, 16'd32155, 16'd65398, 16'd45664, 16'd5035, 16'd28786, 16'd15768, 16'd60929});
	test_expansion(128'h26b850daa1fa9490318963a238878247, {16'd55747, 16'd38937, 16'd56134, 16'd59032, 16'd48572, 16'd37630, 16'd31665, 16'd50920, 16'd53932, 16'd19661, 16'd35800, 16'd21537, 16'd54089, 16'd28790, 16'd49362, 16'd15683, 16'd11621, 16'd65020, 16'd63039, 16'd52534, 16'd53316, 16'd7293, 16'd3265, 16'd20316, 16'd35468, 16'd47299});
	test_expansion(128'h46e9e312b7ada7f0e5cd4b05cd760197, {16'd53710, 16'd59952, 16'd33658, 16'd13618, 16'd42785, 16'd54224, 16'd25248, 16'd14568, 16'd51680, 16'd17382, 16'd46848, 16'd61388, 16'd30415, 16'd26574, 16'd54442, 16'd7172, 16'd44479, 16'd35848, 16'd52081, 16'd24981, 16'd38487, 16'd20131, 16'd64799, 16'd125, 16'd11580, 16'd32553});
	test_expansion(128'h522dad589354723f5e4faebd590e464e, {16'd28176, 16'd19088, 16'd39812, 16'd4808, 16'd24603, 16'd13207, 16'd43532, 16'd21266, 16'd55407, 16'd48344, 16'd64428, 16'd16595, 16'd29831, 16'd38485, 16'd31140, 16'd63813, 16'd65060, 16'd9752, 16'd61699, 16'd20900, 16'd3328, 16'd62227, 16'd44080, 16'd24659, 16'd34297, 16'd634});
	test_expansion(128'h51e31a2a9c678c47bb79f38a5374b0ca, {16'd64186, 16'd62373, 16'd15942, 16'd18568, 16'd27107, 16'd12626, 16'd60447, 16'd43050, 16'd10048, 16'd23526, 16'd49568, 16'd20509, 16'd38438, 16'd11607, 16'd8617, 16'd3444, 16'd52638, 16'd19940, 16'd20566, 16'd30396, 16'd34034, 16'd6035, 16'd50850, 16'd54149, 16'd31457, 16'd41614});
	test_expansion(128'hc338e904c4f1c0512c0354ba21cb1e93, {16'd25341, 16'd8509, 16'd52013, 16'd58009, 16'd3249, 16'd24584, 16'd2819, 16'd11824, 16'd47904, 16'd2897, 16'd4719, 16'd188, 16'd38487, 16'd3150, 16'd25061, 16'd10635, 16'd58907, 16'd5172, 16'd41775, 16'd28353, 16'd40129, 16'd21064, 16'd36002, 16'd965, 16'd34354, 16'd63829});
	test_expansion(128'ha8371cdf6fd54a4500aadd05a56f6736, {16'd34550, 16'd47421, 16'd40660, 16'd45456, 16'd31199, 16'd23562, 16'd18571, 16'd64524, 16'd32768, 16'd10148, 16'd31399, 16'd29124, 16'd8576, 16'd54101, 16'd58534, 16'd19142, 16'd13477, 16'd2338, 16'd31048, 16'd14774, 16'd62386, 16'd25257, 16'd29055, 16'd17434, 16'd8137, 16'd52124});
	test_expansion(128'h9550d852ca01720072150302c29d22a8, {16'd24239, 16'd27748, 16'd16395, 16'd28942, 16'd1046, 16'd15713, 16'd1533, 16'd39266, 16'd60046, 16'd54075, 16'd54707, 16'd31290, 16'd45328, 16'd46284, 16'd47555, 16'd64553, 16'd4288, 16'd22251, 16'd1119, 16'd44092, 16'd794, 16'd1064, 16'd7250, 16'd55989, 16'd36381, 16'd44223});
	test_expansion(128'hdaff3bf24318f92823359594f60e98d9, {16'd40562, 16'd23097, 16'd1421, 16'd48246, 16'd16262, 16'd46562, 16'd39515, 16'd13169, 16'd64972, 16'd58634, 16'd26884, 16'd54022, 16'd23651, 16'd63677, 16'd40570, 16'd15173, 16'd11884, 16'd55796, 16'd53161, 16'd983, 16'd33255, 16'd47191, 16'd15388, 16'd8952, 16'd33444, 16'd8249});
	test_expansion(128'h7f506cdcb830394d2d8f966389f6b1cb, {16'd15830, 16'd34924, 16'd22343, 16'd24116, 16'd45643, 16'd17954, 16'd7548, 16'd21682, 16'd24863, 16'd54373, 16'd45609, 16'd9419, 16'd3935, 16'd39641, 16'd7453, 16'd59, 16'd61770, 16'd31801, 16'd13684, 16'd32648, 16'd47099, 16'd62894, 16'd5167, 16'd54468, 16'd29060, 16'd43054});
	test_expansion(128'hc2707bdf2c7f0189fde8104e29929d80, {16'd44159, 16'd22823, 16'd40907, 16'd15458, 16'd1269, 16'd26684, 16'd23980, 16'd27844, 16'd8170, 16'd61575, 16'd48650, 16'd18483, 16'd32986, 16'd43040, 16'd23127, 16'd39721, 16'd49553, 16'd33788, 16'd2131, 16'd4844, 16'd37089, 16'd31293, 16'd2127, 16'd34370, 16'd62366, 16'd25495});
	test_expansion(128'hafd9327c6a3d46defad1b3cc31f25a13, {16'd44085, 16'd48143, 16'd55642, 16'd59016, 16'd61831, 16'd22327, 16'd17261, 16'd5951, 16'd63998, 16'd61438, 16'd22559, 16'd58786, 16'd58161, 16'd61105, 16'd11695, 16'd50367, 16'd41856, 16'd27652, 16'd58701, 16'd59564, 16'd50566, 16'd6574, 16'd58136, 16'd14853, 16'd47548, 16'd48631});
	test_expansion(128'h57ab7e386dd589741d47b3bc917c19e6, {16'd32787, 16'd50402, 16'd12628, 16'd33666, 16'd58730, 16'd52541, 16'd9281, 16'd56793, 16'd32886, 16'd28228, 16'd24596, 16'd8702, 16'd7446, 16'd33911, 16'd37073, 16'd42636, 16'd62846, 16'd54634, 16'd22265, 16'd64402, 16'd12569, 16'd53683, 16'd20044, 16'd27862, 16'd54940, 16'd50236});
	test_expansion(128'hde7a0f218b2b7f4b4d38721d6f5db275, {16'd45795, 16'd57616, 16'd22744, 16'd34102, 16'd16159, 16'd13085, 16'd16747, 16'd47840, 16'd29206, 16'd29504, 16'd41858, 16'd7148, 16'd9494, 16'd25644, 16'd34647, 16'd4700, 16'd25057, 16'd52005, 16'd50009, 16'd47368, 16'd49197, 16'd10350, 16'd47645, 16'd17156, 16'd30665, 16'd8706});
	test_expansion(128'hab83215d7413d2e45c41c8a549dbf139, {16'd64980, 16'd36124, 16'd49687, 16'd59316, 16'd49028, 16'd61194, 16'd57217, 16'd28647, 16'd29758, 16'd6324, 16'd35044, 16'd42217, 16'd37633, 16'd19761, 16'd16046, 16'd47677, 16'd2494, 16'd667, 16'd54815, 16'd51157, 16'd26322, 16'd30070, 16'd41735, 16'd23130, 16'd433, 16'd34589});
	test_expansion(128'hd590d5058aad791a21a94977a8fae4f5, {16'd62860, 16'd28648, 16'd51406, 16'd3805, 16'd26721, 16'd29286, 16'd27182, 16'd39567, 16'd44657, 16'd6002, 16'd62424, 16'd17880, 16'd28163, 16'd8506, 16'd23003, 16'd31002, 16'd64927, 16'd16696, 16'd18182, 16'd53397, 16'd23671, 16'd61639, 16'd41234, 16'd52481, 16'd19095, 16'd33623});
	test_expansion(128'h1a846b3d326baa60a2de2a4784c020f0, {16'd23228, 16'd60130, 16'd27619, 16'd53746, 16'd32114, 16'd23424, 16'd26929, 16'd9619, 16'd9330, 16'd43160, 16'd52437, 16'd63842, 16'd60918, 16'd30686, 16'd39167, 16'd44602, 16'd50965, 16'd60643, 16'd45229, 16'd43266, 16'd13203, 16'd24305, 16'd17493, 16'd33879, 16'd2189, 16'd28118});
	test_expansion(128'h4371393c1c8a428fc5923e7a9cc6cb3c, {16'd41191, 16'd35255, 16'd33937, 16'd49563, 16'd56341, 16'd6505, 16'd37252, 16'd61758, 16'd49538, 16'd42761, 16'd55956, 16'd49088, 16'd38826, 16'd25134, 16'd54852, 16'd50416, 16'd25678, 16'd24919, 16'd41639, 16'd26892, 16'd27767, 16'd19872, 16'd27343, 16'd16007, 16'd60109, 16'd1968});
	test_expansion(128'h3d30d9ef0d096226e020291100b7814e, {16'd13849, 16'd45735, 16'd59901, 16'd56082, 16'd24592, 16'd37676, 16'd65244, 16'd45513, 16'd64791, 16'd58105, 16'd41874, 16'd50366, 16'd548, 16'd35064, 16'd56278, 16'd57662, 16'd420, 16'd53824, 16'd59770, 16'd8936, 16'd16370, 16'd4876, 16'd48114, 16'd26788, 16'd64856, 16'd18271});
	test_expansion(128'h1ce52b9a47190ffcf4455287329db1bf, {16'd6254, 16'd54068, 16'd30705, 16'd4491, 16'd17362, 16'd40744, 16'd12217, 16'd65305, 16'd40730, 16'd62964, 16'd57214, 16'd54992, 16'd51373, 16'd6077, 16'd30581, 16'd34286, 16'd20663, 16'd18980, 16'd30732, 16'd58226, 16'd45670, 16'd65445, 16'd34197, 16'd24843, 16'd2885, 16'd48677});
	test_expansion(128'he1264ef46ca9e54f637acf5f3bf32e1a, {16'd25203, 16'd36176, 16'd39405, 16'd55478, 16'd1457, 16'd38191, 16'd17999, 16'd55098, 16'd38001, 16'd52844, 16'd29605, 16'd37019, 16'd63416, 16'd25957, 16'd63425, 16'd21837, 16'd65228, 16'd39280, 16'd60686, 16'd9734, 16'd62400, 16'd10340, 16'd39479, 16'd48555, 16'd16586, 16'd36984});
	test_expansion(128'h241c5f4db5dbafff56523b3ae9daca14, {16'd62457, 16'd26476, 16'd12807, 16'd41052, 16'd35819, 16'd27727, 16'd3644, 16'd12841, 16'd39845, 16'd56536, 16'd65073, 16'd30446, 16'd107, 16'd5829, 16'd8485, 16'd35654, 16'd17966, 16'd12476, 16'd8570, 16'd7977, 16'd57986, 16'd48878, 16'd22710, 16'd23629, 16'd35217, 16'd33219});
	test_expansion(128'ha1cadf8410945132ea51ae4d08efc6c7, {16'd57882, 16'd46944, 16'd1722, 16'd37182, 16'd40101, 16'd18933, 16'd15741, 16'd64743, 16'd57451, 16'd17567, 16'd23413, 16'd17987, 16'd63755, 16'd5727, 16'd55405, 16'd47184, 16'd12976, 16'd57144, 16'd18273, 16'd53406, 16'd60144, 16'd53960, 16'd47767, 16'd18616, 16'd7333, 16'd8165});
	test_expansion(128'h39e8cd124245e11465d559862a6a321d, {16'd29210, 16'd45379, 16'd7725, 16'd10770, 16'd27154, 16'd11312, 16'd416, 16'd33411, 16'd38646, 16'd11547, 16'd52474, 16'd56181, 16'd39993, 16'd5390, 16'd51755, 16'd28322, 16'd14846, 16'd46676, 16'd13438, 16'd57549, 16'd63605, 16'd7872, 16'd13837, 16'd5296, 16'd45692, 16'd42850});
	test_expansion(128'h9db088f36c3172ec18e2c5e1a4948cea, {16'd30984, 16'd36690, 16'd37504, 16'd48684, 16'd65535, 16'd26456, 16'd3747, 16'd11524, 16'd35702, 16'd59966, 16'd2652, 16'd2635, 16'd42887, 16'd36313, 16'd63022, 16'd11152, 16'd30220, 16'd15972, 16'd52006, 16'd26414, 16'd53001, 16'd45583, 16'd15798, 16'd26787, 16'd50080, 16'd12675});
	test_expansion(128'h667ee76c23fe226e3d2abd6e71865b21, {16'd27797, 16'd57623, 16'd18945, 16'd55497, 16'd46665, 16'd51144, 16'd54432, 16'd28671, 16'd33917, 16'd58912, 16'd3577, 16'd18440, 16'd11691, 16'd16677, 16'd30124, 16'd14844, 16'd39781, 16'd1891, 16'd11485, 16'd35456, 16'd54484, 16'd45569, 16'd17205, 16'd1349, 16'd53908, 16'd36754});
	test_expansion(128'hf722808922a2423d30bdcf9cb1c16279, {16'd7778, 16'd33084, 16'd2503, 16'd54255, 16'd51912, 16'd38709, 16'd20939, 16'd59654, 16'd54446, 16'd16878, 16'd4829, 16'd43960, 16'd26386, 16'd38020, 16'd16318, 16'd49505, 16'd29177, 16'd12568, 16'd59608, 16'd53045, 16'd32758, 16'd2437, 16'd26735, 16'd35362, 16'd15930, 16'd3215});
	test_expansion(128'h2646e0ed614c8a086ea450059cd2e33e, {16'd13679, 16'd17725, 16'd45813, 16'd13933, 16'd5444, 16'd31606, 16'd8205, 16'd34751, 16'd39005, 16'd47011, 16'd21281, 16'd64594, 16'd14812, 16'd55244, 16'd6003, 16'd57046, 16'd64997, 16'd21016, 16'd49243, 16'd18879, 16'd31789, 16'd17420, 16'd3555, 16'd14261, 16'd33537, 16'd59078});
	test_expansion(128'haffb402e2d1befc7ccf00d643b0adccd, {16'd22996, 16'd54969, 16'd59479, 16'd23216, 16'd17848, 16'd59333, 16'd20439, 16'd11725, 16'd24405, 16'd29615, 16'd30136, 16'd62977, 16'd48530, 16'd50985, 16'd48351, 16'd32777, 16'd56392, 16'd20380, 16'd24128, 16'd57727, 16'd47367, 16'd18757, 16'd30876, 16'd48651, 16'd39170, 16'd41518});
	test_expansion(128'h4fc3332e09097d2297e2834c06b7076e, {16'd18334, 16'd54927, 16'd33010, 16'd38725, 16'd64896, 16'd30312, 16'd7768, 16'd23114, 16'd60412, 16'd55038, 16'd40951, 16'd43026, 16'd32, 16'd43370, 16'd9132, 16'd24948, 16'd61518, 16'd56736, 16'd24251, 16'd59964, 16'd28028, 16'd22772, 16'd61844, 16'd56618, 16'd58749, 16'd47715});
	test_expansion(128'hdb095f8d658b791d39020c32a1fbfe8b, {16'd61619, 16'd31224, 16'd30794, 16'd24450, 16'd63518, 16'd28319, 16'd19541, 16'd52341, 16'd40919, 16'd9386, 16'd18602, 16'd61380, 16'd39748, 16'd35331, 16'd7353, 16'd63679, 16'd61062, 16'd26733, 16'd25836, 16'd39010, 16'd7899, 16'd45986, 16'd54885, 16'd22287, 16'd35894, 16'd9915});
	test_expansion(128'hc4bea1869033c2d3ceae40f4b4c6b5df, {16'd63163, 16'd49177, 16'd37225, 16'd23705, 16'd55683, 16'd2132, 16'd30237, 16'd44832, 16'd4291, 16'd46320, 16'd29027, 16'd57600, 16'd26851, 16'd20399, 16'd46112, 16'd7869, 16'd41621, 16'd38796, 16'd39275, 16'd20765, 16'd45792, 16'd23097, 16'd48665, 16'd22383, 16'd26999, 16'd62044});
	test_expansion(128'h7a0dd0fff466521d65448b4eb381f622, {16'd4106, 16'd48310, 16'd42946, 16'd8383, 16'd58778, 16'd60819, 16'd41463, 16'd29959, 16'd14159, 16'd8431, 16'd27063, 16'd16083, 16'd49028, 16'd36781, 16'd5985, 16'd23176, 16'd56604, 16'd10117, 16'd18626, 16'd33151, 16'd50706, 16'd10450, 16'd24998, 16'd622, 16'd2318, 16'd45847});
	test_expansion(128'h19c631ed7d3c38f7c9eeb1cff7a9a4fb, {16'd33415, 16'd53267, 16'd53497, 16'd10957, 16'd35574, 16'd17321, 16'd28749, 16'd37768, 16'd9530, 16'd64722, 16'd26167, 16'd39226, 16'd7949, 16'd52282, 16'd5438, 16'd41054, 16'd64891, 16'd37768, 16'd38003, 16'd52305, 16'd55397, 16'd20565, 16'd57336, 16'd58710, 16'd51045, 16'd17847});
	test_expansion(128'hccebee4b2e2847948cb7ed690f9fa349, {16'd5565, 16'd8202, 16'd46117, 16'd40397, 16'd17882, 16'd13476, 16'd5519, 16'd50784, 16'd12235, 16'd20894, 16'd31387, 16'd32255, 16'd52923, 16'd12929, 16'd57604, 16'd44563, 16'd37915, 16'd3333, 16'd27145, 16'd27721, 16'd3007, 16'd25358, 16'd56325, 16'd7240, 16'd17946, 16'd7912});
	test_expansion(128'he40d96b8f9a83cd226b2ed7a5d419752, {16'd58465, 16'd5537, 16'd21726, 16'd21920, 16'd65079, 16'd36512, 16'd28986, 16'd8372, 16'd65474, 16'd57259, 16'd45916, 16'd5949, 16'd37045, 16'd39157, 16'd21427, 16'd25716, 16'd51722, 16'd45994, 16'd37321, 16'd3701, 16'd33692, 16'd2934, 16'd16760, 16'd25050, 16'd21486, 16'd38305});
	test_expansion(128'h326b0d73c37f3135a137eebd568273b5, {16'd47537, 16'd32116, 16'd17400, 16'd62995, 16'd42515, 16'd40475, 16'd26310, 16'd64057, 16'd3838, 16'd31389, 16'd26138, 16'd35087, 16'd15960, 16'd14872, 16'd38837, 16'd44748, 16'd28385, 16'd47499, 16'd7062, 16'd34125, 16'd24851, 16'd11142, 16'd60113, 16'd52677, 16'd24187, 16'd61505});
	test_expansion(128'h2edc5dfdb2eb4acff20527019c93d338, {16'd19994, 16'd60434, 16'd45307, 16'd38456, 16'd20152, 16'd55941, 16'd43490, 16'd24066, 16'd38925, 16'd22977, 16'd29000, 16'd52349, 16'd14340, 16'd25582, 16'd169, 16'd19125, 16'd10612, 16'd25514, 16'd60299, 16'd22842, 16'd12741, 16'd38505, 16'd49688, 16'd6149, 16'd29891, 16'd32505});
	test_expansion(128'hc5927307dbc2fd00d08e657dde4c65ba, {16'd27346, 16'd30921, 16'd20957, 16'd35276, 16'd3887, 16'd25830, 16'd50504, 16'd8123, 16'd25946, 16'd40653, 16'd64587, 16'd20700, 16'd24228, 16'd55989, 16'd18083, 16'd24309, 16'd57269, 16'd26617, 16'd64074, 16'd18961, 16'd7896, 16'd47633, 16'd15492, 16'd56878, 16'd44991, 16'd38978});
	test_expansion(128'hc1a232566ea562c353238a4937fbaa63, {16'd56323, 16'd2563, 16'd29968, 16'd43076, 16'd62948, 16'd63003, 16'd63090, 16'd61550, 16'd37429, 16'd17829, 16'd57256, 16'd13509, 16'd2514, 16'd12798, 16'd55468, 16'd54236, 16'd30577, 16'd27575, 16'd9092, 16'd28209, 16'd16381, 16'd7300, 16'd4893, 16'd62817, 16'd32394, 16'd30887});
	test_expansion(128'hd0d7dc3804a506d68d313ba88dc380c7, {16'd17686, 16'd43752, 16'd38821, 16'd11992, 16'd3048, 16'd54169, 16'd31418, 16'd2517, 16'd51013, 16'd35297, 16'd46374, 16'd30382, 16'd42012, 16'd29583, 16'd28561, 16'd48473, 16'd11402, 16'd64263, 16'd11987, 16'd4347, 16'd26668, 16'd10315, 16'd34408, 16'd41472, 16'd7950, 16'd28041});
	test_expansion(128'h95e6d85f4b3e06e840c2340f9caf054e, {16'd4398, 16'd30373, 16'd16740, 16'd15588, 16'd58461, 16'd30137, 16'd56208, 16'd13045, 16'd23755, 16'd63158, 16'd49163, 16'd26674, 16'd23546, 16'd59207, 16'd8035, 16'd60840, 16'd24315, 16'd29447, 16'd21226, 16'd9439, 16'd12528, 16'd23999, 16'd7437, 16'd48145, 16'd21524, 16'd33428});
	test_expansion(128'h90ea95921caf354a10438c8708359e53, {16'd50000, 16'd43310, 16'd48551, 16'd20578, 16'd29716, 16'd61787, 16'd61262, 16'd41259, 16'd40741, 16'd5603, 16'd17041, 16'd17758, 16'd29424, 16'd48141, 16'd38757, 16'd12697, 16'd7758, 16'd10946, 16'd37657, 16'd17955, 16'd34053, 16'd46160, 16'd28055, 16'd21267, 16'd23308, 16'd1082});
	test_expansion(128'h2acfbd83ba91de1fb8fdfa18c3bf2c38, {16'd19770, 16'd10698, 16'd43524, 16'd10075, 16'd6419, 16'd33648, 16'd39245, 16'd37361, 16'd5562, 16'd12072, 16'd22598, 16'd49711, 16'd18051, 16'd40999, 16'd62009, 16'd22250, 16'd8331, 16'd18519, 16'd35357, 16'd7909, 16'd63376, 16'd8835, 16'd6352, 16'd1042, 16'd48361, 16'd37361});
	test_expansion(128'h63024e0480a564c71f1d4dc4514beb5e, {16'd61181, 16'd27779, 16'd39155, 16'd55455, 16'd2382, 16'd14164, 16'd38397, 16'd33225, 16'd18026, 16'd39428, 16'd37256, 16'd53427, 16'd45105, 16'd58552, 16'd141, 16'd62627, 16'd3661, 16'd6214, 16'd29949, 16'd42618, 16'd9473, 16'd17307, 16'd52683, 16'd49097, 16'd16997, 16'd45255});
	test_expansion(128'h9aa5ce4f151ea2409f324fe2e7cfad50, {16'd52535, 16'd27593, 16'd18868, 16'd63767, 16'd42163, 16'd48710, 16'd63595, 16'd12210, 16'd55542, 16'd64894, 16'd41979, 16'd15063, 16'd46328, 16'd37144, 16'd39737, 16'd23927, 16'd761, 16'd25138, 16'd5440, 16'd41218, 16'd13082, 16'd744, 16'd5239, 16'd13505, 16'd37450, 16'd20414});
	test_expansion(128'h34fe85d7960bbd0c1d2bccb2d60dc7f7, {16'd32645, 16'd43805, 16'd13022, 16'd62175, 16'd34054, 16'd5889, 16'd52476, 16'd25780, 16'd44454, 16'd37241, 16'd62179, 16'd23054, 16'd7044, 16'd14932, 16'd31389, 16'd43052, 16'd34727, 16'd29517, 16'd33063, 16'd14100, 16'd15614, 16'd13066, 16'd6835, 16'd12588, 16'd28218, 16'd27009});
	test_expansion(128'h7fba3de39c8a8ca65d2108929ac4b742, {16'd19978, 16'd64160, 16'd17645, 16'd57426, 16'd21060, 16'd34927, 16'd15450, 16'd56568, 16'd63849, 16'd21136, 16'd45245, 16'd44466, 16'd59410, 16'd20539, 16'd52553, 16'd40406, 16'd42468, 16'd36459, 16'd18194, 16'd28923, 16'd51882, 16'd14844, 16'd37597, 16'd47077, 16'd44648, 16'd54040});
	test_expansion(128'h93895120bdc73c16eb2936ab4cf3720e, {16'd26343, 16'd35283, 16'd16802, 16'd49435, 16'd33006, 16'd56643, 16'd5370, 16'd10601, 16'd48859, 16'd37023, 16'd6275, 16'd36206, 16'd5987, 16'd18726, 16'd4597, 16'd50545, 16'd442, 16'd29642, 16'd61276, 16'd32433, 16'd14193, 16'd34785, 16'd51808, 16'd50236, 16'd62743, 16'd64362});
	test_expansion(128'h4e5e6b11da44e243852df9bac04f8297, {16'd56616, 16'd18182, 16'd10997, 16'd19841, 16'd45149, 16'd23352, 16'd31599, 16'd44023, 16'd53408, 16'd52685, 16'd48503, 16'd51670, 16'd4749, 16'd33044, 16'd56584, 16'd13503, 16'd14597, 16'd20119, 16'd20664, 16'd51875, 16'd51959, 16'd35205, 16'd61209, 16'd55965, 16'd45354, 16'd45187});
	test_expansion(128'h32361e75f4b718396cd6ddd437437fd1, {16'd57251, 16'd32292, 16'd30180, 16'd45152, 16'd39377, 16'd3369, 16'd42020, 16'd57469, 16'd8607, 16'd50332, 16'd64480, 16'd13049, 16'd29407, 16'd53604, 16'd62246, 16'd22624, 16'd34468, 16'd2791, 16'd29630, 16'd49079, 16'd37529, 16'd30027, 16'd23311, 16'd65237, 16'd60283, 16'd22188});
	test_expansion(128'h1972e0785c19744a2a75173bdf928522, {16'd10042, 16'd38736, 16'd60495, 16'd39284, 16'd59788, 16'd54442, 16'd31608, 16'd55781, 16'd55563, 16'd53205, 16'd52266, 16'd52861, 16'd47774, 16'd35944, 16'd54118, 16'd20963, 16'd40779, 16'd19279, 16'd28579, 16'd9103, 16'd56970, 16'd11612, 16'd11885, 16'd6184, 16'd61611, 16'd48857});
	test_expansion(128'h2a4d9e74c63d882646ffde11681a439f, {16'd27875, 16'd43874, 16'd27146, 16'd33227, 16'd7305, 16'd30181, 16'd62932, 16'd33696, 16'd27696, 16'd33988, 16'd13719, 16'd54088, 16'd17895, 16'd17294, 16'd8911, 16'd22808, 16'd40948, 16'd64523, 16'd49345, 16'd31466, 16'd26009, 16'd7307, 16'd62986, 16'd53646, 16'd2727, 16'd7629});
	test_expansion(128'h1147f0aff4aef9832591459fd3cb68e0, {16'd42195, 16'd6089, 16'd14298, 16'd28038, 16'd48312, 16'd30554, 16'd57073, 16'd28226, 16'd61138, 16'd54751, 16'd42569, 16'd29607, 16'd18095, 16'd57146, 16'd51994, 16'd62223, 16'd62316, 16'd36972, 16'd54037, 16'd13255, 16'd10113, 16'd13877, 16'd19818, 16'd43033, 16'd48368, 16'd27828});
	test_expansion(128'h686874bd4e77d05dd4749e317fcf9574, {16'd7592, 16'd26674, 16'd41691, 16'd19274, 16'd24911, 16'd1469, 16'd4093, 16'd3246, 16'd41924, 16'd3175, 16'd51271, 16'd31793, 16'd35256, 16'd27376, 16'd13894, 16'd28079, 16'd855, 16'd4315, 16'd25266, 16'd38411, 16'd17908, 16'd45886, 16'd9201, 16'd29430, 16'd55291, 16'd65459});
	test_expansion(128'he7cde723333c083add271f3c1fdafc68, {16'd12596, 16'd42923, 16'd19969, 16'd50483, 16'd56056, 16'd30653, 16'd37224, 16'd5102, 16'd47273, 16'd47721, 16'd57762, 16'd55859, 16'd48391, 16'd8639, 16'd40284, 16'd54541, 16'd3275, 16'd9634, 16'd19749, 16'd28370, 16'd7509, 16'd60868, 16'd3066, 16'd48798, 16'd63653, 16'd47140});
	test_expansion(128'h029d2699965622743646e2899c70d969, {16'd174, 16'd31780, 16'd39542, 16'd33947, 16'd36488, 16'd62290, 16'd54033, 16'd40461, 16'd48533, 16'd39102, 16'd18079, 16'd18508, 16'd51660, 16'd564, 16'd53225, 16'd52039, 16'd7320, 16'd51536, 16'd51014, 16'd55760, 16'd35437, 16'd45295, 16'd14097, 16'd54753, 16'd51981, 16'd30402});
	test_expansion(128'haa850931d4fe36340c854030a516f4f3, {16'd17781, 16'd50311, 16'd10067, 16'd56739, 16'd23946, 16'd52272, 16'd4133, 16'd30214, 16'd43487, 16'd3372, 16'd20467, 16'd55915, 16'd12754, 16'd30583, 16'd16219, 16'd13206, 16'd11713, 16'd8773, 16'd65329, 16'd60257, 16'd34803, 16'd53608, 16'd14736, 16'd54646, 16'd19666, 16'd27275});
	test_expansion(128'h3074177cc8c8c2a40811a84b0baaf8ef, {16'd38819, 16'd58713, 16'd50492, 16'd3858, 16'd15082, 16'd59701, 16'd60010, 16'd62073, 16'd43685, 16'd24431, 16'd16894, 16'd64406, 16'd12720, 16'd39964, 16'd5795, 16'd55613, 16'd59135, 16'd37628, 16'd434, 16'd51126, 16'd18530, 16'd57179, 16'd36459, 16'd27067, 16'd39190, 16'd2461});
	test_expansion(128'h0a9ce43040af27caf62ff2402399a462, {16'd33991, 16'd7600, 16'd1785, 16'd8728, 16'd53981, 16'd14527, 16'd26391, 16'd53945, 16'd37603, 16'd39466, 16'd53556, 16'd63847, 16'd16325, 16'd54026, 16'd28460, 16'd45080, 16'd13993, 16'd48053, 16'd493, 16'd61104, 16'd43722, 16'd24265, 16'd63025, 16'd29940, 16'd49815, 16'd39780});
	test_expansion(128'hf6fab02ef283e85685c9ed6495308131, {16'd2580, 16'd38357, 16'd57554, 16'd37372, 16'd38048, 16'd36540, 16'd42090, 16'd46652, 16'd28587, 16'd52069, 16'd57125, 16'd49828, 16'd29755, 16'd12974, 16'd40983, 16'd53997, 16'd55291, 16'd39057, 16'd19795, 16'd23569, 16'd39263, 16'd41342, 16'd5820, 16'd47948, 16'd33820, 16'd35939});
	test_expansion(128'h33e0630f29d4a2bb00865d48a29029a4, {16'd25049, 16'd15763, 16'd9823, 16'd36252, 16'd27661, 16'd17032, 16'd17362, 16'd21130, 16'd62961, 16'd4817, 16'd58360, 16'd41159, 16'd15251, 16'd53990, 16'd48748, 16'd36572, 16'd314, 16'd25941, 16'd51975, 16'd2775, 16'd64316, 16'd52103, 16'd20749, 16'd9592, 16'd17372, 16'd60684});
	test_expansion(128'h3e6ea649a74dda4b18698483b15e7274, {16'd17731, 16'd3676, 16'd58905, 16'd44047, 16'd52181, 16'd1272, 16'd29703, 16'd47937, 16'd29204, 16'd27058, 16'd28413, 16'd59937, 16'd49374, 16'd52127, 16'd5985, 16'd55629, 16'd54431, 16'd23515, 16'd56761, 16'd7159, 16'd22667, 16'd7558, 16'd46185, 16'd16900, 16'd38510, 16'd16176});
	test_expansion(128'h334e8dbd997a5853664dc4005e549803, {16'd3913, 16'd61737, 16'd35636, 16'd52187, 16'd23761, 16'd65121, 16'd36558, 16'd62500, 16'd52047, 16'd61146, 16'd9838, 16'd23674, 16'd18649, 16'd28735, 16'd57320, 16'd2209, 16'd49219, 16'd8938, 16'd64609, 16'd42524, 16'd35112, 16'd14076, 16'd62212, 16'd22281, 16'd45279, 16'd8070});
	test_expansion(128'h156283c88f8fe13620ff975ca7c6b278, {16'd24780, 16'd8195, 16'd50636, 16'd20383, 16'd17272, 16'd62062, 16'd31634, 16'd4416, 16'd30439, 16'd5782, 16'd22336, 16'd23662, 16'd63837, 16'd43673, 16'd20193, 16'd397, 16'd20953, 16'd16293, 16'd28010, 16'd43153, 16'd4321, 16'd22491, 16'd26435, 16'd31982, 16'd59596, 16'd47614});
	test_expansion(128'hab5e18220daced47b3dcc0a40eed5cb2, {16'd34571, 16'd54909, 16'd52348, 16'd27588, 16'd44917, 16'd29733, 16'd23578, 16'd19863, 16'd16381, 16'd62545, 16'd35792, 16'd58142, 16'd1342, 16'd52307, 16'd51997, 16'd48989, 16'd35080, 16'd51180, 16'd3335, 16'd52693, 16'd26491, 16'd47579, 16'd16173, 16'd4092, 16'd27124, 16'd19030});
	test_expansion(128'he27dbe23f6258e7dae0f715570fe24a2, {16'd19395, 16'd65374, 16'd47021, 16'd10358, 16'd3701, 16'd17064, 16'd45302, 16'd48429, 16'd61517, 16'd44510, 16'd19880, 16'd11219, 16'd34437, 16'd40651, 16'd56061, 16'd54991, 16'd43337, 16'd3458, 16'd6171, 16'd14641, 16'd45870, 16'd29390, 16'd21269, 16'd25460, 16'd10798, 16'd40911});
	test_expansion(128'h6c125dcf566b3f3433b1eae6dc69a3f5, {16'd8077, 16'd17419, 16'd50511, 16'd62813, 16'd3523, 16'd8255, 16'd36795, 16'd25790, 16'd6654, 16'd15818, 16'd41120, 16'd59558, 16'd54832, 16'd18218, 16'd22271, 16'd717, 16'd59304, 16'd20753, 16'd17064, 16'd38289, 16'd39104, 16'd60046, 16'd31502, 16'd4608, 16'd27251, 16'd36196});
	test_expansion(128'h827cdf78cc08f7157e4d96cdb4aae18e, {16'd25635, 16'd54385, 16'd50624, 16'd49409, 16'd3935, 16'd27649, 16'd40248, 16'd10408, 16'd14773, 16'd11007, 16'd59075, 16'd26883, 16'd32368, 16'd22027, 16'd10232, 16'd37223, 16'd1086, 16'd26558, 16'd60627, 16'd63431, 16'd17481, 16'd57905, 16'd46243, 16'd2104, 16'd12427, 16'd17914});
	test_expansion(128'hcd64c29e61029e4148eb10d7de881fee, {16'd49602, 16'd16469, 16'd56906, 16'd37399, 16'd29350, 16'd45482, 16'd17220, 16'd47064, 16'd45353, 16'd6435, 16'd31261, 16'd8435, 16'd33741, 16'd51994, 16'd61008, 16'd19636, 16'd36034, 16'd18056, 16'd51987, 16'd23003, 16'd57645, 16'd60996, 16'd35430, 16'd25731, 16'd46400, 16'd32153});
	test_expansion(128'hcea0fd734a247ba8e9bed203b1197bae, {16'd45410, 16'd44353, 16'd17337, 16'd22601, 16'd41129, 16'd15311, 16'd15087, 16'd65451, 16'd64376, 16'd47789, 16'd58800, 16'd43721, 16'd4206, 16'd11428, 16'd4663, 16'd62184, 16'd48718, 16'd11734, 16'd3124, 16'd53278, 16'd58207, 16'd48213, 16'd9914, 16'd34953, 16'd65297, 16'd19596});
	test_expansion(128'h6d7175582cfe25c9b8188c4551fedf4c, {16'd9780, 16'd11801, 16'd32833, 16'd32224, 16'd12206, 16'd13309, 16'd35623, 16'd32663, 16'd41588, 16'd3767, 16'd52264, 16'd57699, 16'd51353, 16'd45078, 16'd17954, 16'd62739, 16'd53587, 16'd15606, 16'd59053, 16'd25570, 16'd24371, 16'd17716, 16'd26389, 16'd10104, 16'd50041, 16'd56397});
	test_expansion(128'h30a02c7c67e487e6511c42f5cc85d226, {16'd53665, 16'd39407, 16'd35466, 16'd3357, 16'd42162, 16'd37064, 16'd56508, 16'd16105, 16'd30940, 16'd11972, 16'd9587, 16'd63248, 16'd45249, 16'd45823, 16'd29423, 16'd51482, 16'd33822, 16'd64479, 16'd11986, 16'd41651, 16'd43819, 16'd59700, 16'd8220, 16'd19301, 16'd4540, 16'd51529});
	test_expansion(128'hc0ec308c1960e5532d90208d99dd172c, {16'd43399, 16'd4624, 16'd3724, 16'd21831, 16'd9017, 16'd14533, 16'd1631, 16'd16014, 16'd24416, 16'd4401, 16'd13815, 16'd62821, 16'd5053, 16'd5872, 16'd51303, 16'd38836, 16'd56975, 16'd46606, 16'd15036, 16'd21899, 16'd60937, 16'd39109, 16'd62826, 16'd62916, 16'd57529, 16'd41739});
	test_expansion(128'h21223869f988709793ce05d610322000, {16'd55581, 16'd32539, 16'd62027, 16'd60759, 16'd2947, 16'd44104, 16'd6953, 16'd54905, 16'd16728, 16'd50285, 16'd49891, 16'd35754, 16'd31934, 16'd34217, 16'd31865, 16'd40842, 16'd25646, 16'd35631, 16'd9346, 16'd50016, 16'd60160, 16'd1126, 16'd57440, 16'd50599, 16'd46778, 16'd56632});
	test_expansion(128'h4c768061c69ccb9cbbd7f7afe76541bf, {16'd237, 16'd48346, 16'd63385, 16'd48446, 16'd36968, 16'd150, 16'd34607, 16'd15252, 16'd64864, 16'd62406, 16'd33243, 16'd63078, 16'd24811, 16'd34152, 16'd2659, 16'd46246, 16'd10225, 16'd41747, 16'd11498, 16'd19542, 16'd43671, 16'd11003, 16'd41939, 16'd29886, 16'd45164, 16'd18834});
	test_expansion(128'hc0f08febc242036c44bb887684b5dbd3, {16'd27248, 16'd17803, 16'd48652, 16'd59676, 16'd19951, 16'd16842, 16'd58572, 16'd37488, 16'd50062, 16'd39597, 16'd12805, 16'd38359, 16'd18460, 16'd38551, 16'd64554, 16'd24851, 16'd33572, 16'd16254, 16'd57435, 16'd29801, 16'd26182, 16'd23354, 16'd46645, 16'd49530, 16'd23011, 16'd11937});
	test_expansion(128'ha8c12c680ab4b25c4f020bf8912b3c19, {16'd55077, 16'd27797, 16'd22070, 16'd10030, 16'd19355, 16'd47012, 16'd49597, 16'd63829, 16'd27504, 16'd27068, 16'd24788, 16'd46188, 16'd42332, 16'd60174, 16'd60197, 16'd35167, 16'd14212, 16'd55354, 16'd36951, 16'd48663, 16'd8693, 16'd28172, 16'd44373, 16'd22304, 16'd44801, 16'd29763});
	test_expansion(128'h524af8c2c47c8524a22d087ae2cf8a21, {16'd50627, 16'd21800, 16'd28021, 16'd18071, 16'd5423, 16'd46115, 16'd29147, 16'd12362, 16'd51122, 16'd31138, 16'd52976, 16'd17168, 16'd42763, 16'd17169, 16'd46699, 16'd54828, 16'd10453, 16'd23603, 16'd56373, 16'd40015, 16'd30644, 16'd16306, 16'd39006, 16'd16429, 16'd26168, 16'd58510});
	test_expansion(128'h20b8dd6a3da15eddb879c74abe2239d7, {16'd16721, 16'd65092, 16'd60994, 16'd27504, 16'd56272, 16'd56087, 16'd59543, 16'd58811, 16'd19615, 16'd8713, 16'd4492, 16'd14753, 16'd49368, 16'd21319, 16'd17971, 16'd48600, 16'd28783, 16'd28195, 16'd32345, 16'd54128, 16'd39092, 16'd16150, 16'd63258, 16'd930, 16'd15234, 16'd60938});
	test_expansion(128'hb346e678888d47201b65b54e794008a4, {16'd54823, 16'd43361, 16'd61256, 16'd32191, 16'd52500, 16'd8186, 16'd5330, 16'd53471, 16'd25712, 16'd13986, 16'd47515, 16'd7981, 16'd26108, 16'd46371, 16'd51980, 16'd2031, 16'd57817, 16'd63760, 16'd42186, 16'd15575, 16'd3561, 16'd42603, 16'd35968, 16'd44366, 16'd44484, 16'd63457});
	test_expansion(128'h6ef5808b129f4fef018653123ca3e7b1, {16'd20472, 16'd41762, 16'd48991, 16'd42593, 16'd62371, 16'd48232, 16'd59929, 16'd15602, 16'd32158, 16'd16376, 16'd24987, 16'd61616, 16'd50989, 16'd40047, 16'd27628, 16'd62141, 16'd21876, 16'd64736, 16'd37028, 16'd48974, 16'd49885, 16'd65444, 16'd15088, 16'd60492, 16'd24462, 16'd64754});
	test_expansion(128'he086b61476ce7fce0dbecf895cdeeb2f, {16'd29201, 16'd1895, 16'd35143, 16'd41281, 16'd43567, 16'd52183, 16'd45875, 16'd17264, 16'd32322, 16'd29602, 16'd1855, 16'd20419, 16'd42880, 16'd6735, 16'd34543, 16'd15990, 16'd15545, 16'd11966, 16'd214, 16'd41377, 16'd60689, 16'd15348, 16'd480, 16'd37901, 16'd45153, 16'd6413});
	test_expansion(128'h33a8f0870a79bb506af4422911244776, {16'd58531, 16'd59864, 16'd52179, 16'd20993, 16'd23991, 16'd6482, 16'd51291, 16'd23714, 16'd54789, 16'd12150, 16'd51507, 16'd3441, 16'd4091, 16'd59532, 16'd39937, 16'd47623, 16'd2524, 16'd33627, 16'd43803, 16'd50793, 16'd51052, 16'd30921, 16'd5878, 16'd10902, 16'd3666, 16'd22297});
	test_expansion(128'h7fd37ccb4f72ebbf9c4ec5e1b5b2d863, {16'd41272, 16'd6383, 16'd49149, 16'd54575, 16'd54656, 16'd31548, 16'd48171, 16'd26038, 16'd16402, 16'd5844, 16'd53451, 16'd42253, 16'd45911, 16'd47650, 16'd12070, 16'd6152, 16'd34311, 16'd41162, 16'd17092, 16'd24089, 16'd26978, 16'd26062, 16'd41051, 16'd5058, 16'd47481, 16'd25429});
	test_expansion(128'h160affddd658e5183ceb4001d7dfc85a, {16'd459, 16'd14784, 16'd392, 16'd15828, 16'd4037, 16'd50112, 16'd6129, 16'd63737, 16'd14800, 16'd8093, 16'd9654, 16'd16811, 16'd21955, 16'd18714, 16'd20645, 16'd11845, 16'd11539, 16'd35488, 16'd30322, 16'd36459, 16'd27175, 16'd37521, 16'd56797, 16'd11758, 16'd228, 16'd54753});
	test_expansion(128'h74c53aff5e76d946033ff3db12869f0c, {16'd5463, 16'd62904, 16'd40353, 16'd21873, 16'd28944, 16'd44916, 16'd13080, 16'd38627, 16'd34563, 16'd10358, 16'd44081, 16'd46434, 16'd23858, 16'd49087, 16'd57506, 16'd64932, 16'd37619, 16'd58252, 16'd10514, 16'd45896, 16'd12743, 16'd30569, 16'd12357, 16'd12996, 16'd17479, 16'd45739});
	test_expansion(128'h9918c2f2b0cfa36ffa85f560e68179da, {16'd30442, 16'd38236, 16'd19599, 16'd55544, 16'd59882, 16'd58614, 16'd56591, 16'd23712, 16'd678, 16'd38597, 16'd12483, 16'd20346, 16'd58025, 16'd62187, 16'd63550, 16'd35907, 16'd6511, 16'd37752, 16'd56974, 16'd5879, 16'd7826, 16'd31947, 16'd63781, 16'd21353, 16'd42775, 16'd64568});
	test_expansion(128'hd736bb6e322fbc80b4dda6ff9fcf30ae, {16'd47635, 16'd50569, 16'd50758, 16'd60195, 16'd57802, 16'd34664, 16'd64986, 16'd36719, 16'd4075, 16'd65145, 16'd59036, 16'd3651, 16'd55075, 16'd26915, 16'd21149, 16'd54487, 16'd61975, 16'd34983, 16'd6275, 16'd22379, 16'd47796, 16'd1859, 16'd12839, 16'd44211, 16'd57121, 16'd29011});
	test_expansion(128'h184a9e70dd2291969b8a3d959b31015f, {16'd16829, 16'd49953, 16'd52910, 16'd35658, 16'd26591, 16'd36799, 16'd44717, 16'd1355, 16'd20422, 16'd4172, 16'd23590, 16'd27751, 16'd43049, 16'd44426, 16'd48878, 16'd49635, 16'd50257, 16'd64897, 16'd28832, 16'd50243, 16'd33107, 16'd32707, 16'd39070, 16'd27544, 16'd15848, 16'd11914});
	test_expansion(128'hd212270434ce945f2f8fb54b761145e8, {16'd59952, 16'd3726, 16'd35401, 16'd39324, 16'd34971, 16'd10926, 16'd25936, 16'd25137, 16'd37167, 16'd5317, 16'd53509, 16'd51038, 16'd44727, 16'd4469, 16'd16319, 16'd14054, 16'd51886, 16'd44391, 16'd2174, 16'd37638, 16'd33156, 16'd12001, 16'd19343, 16'd10131, 16'd7248, 16'd44353});
	test_expansion(128'hb64cd4dd85b2b6776a7eedf7fb4666a8, {16'd26166, 16'd28478, 16'd15668, 16'd43454, 16'd24449, 16'd60433, 16'd34101, 16'd4608, 16'd15007, 16'd24274, 16'd27162, 16'd15705, 16'd23933, 16'd50046, 16'd22783, 16'd48314, 16'd27269, 16'd34712, 16'd41421, 16'd44266, 16'd1432, 16'd54842, 16'd22620, 16'd61933, 16'd19134, 16'd38616});
	test_expansion(128'hcf278f1e0185b5c1f3c1104942d3cc3e, {16'd54398, 16'd60970, 16'd52645, 16'd15130, 16'd52560, 16'd53308, 16'd10480, 16'd8080, 16'd60912, 16'd49650, 16'd18002, 16'd49628, 16'd34154, 16'd24704, 16'd30218, 16'd50536, 16'd48766, 16'd65392, 16'd3699, 16'd64443, 16'd6985, 16'd6099, 16'd26386, 16'd48375, 16'd24548, 16'd30301});
	test_expansion(128'h1be3dc797c39d64b0456a1e686d19fb5, {16'd60600, 16'd20086, 16'd30494, 16'd59973, 16'd352, 16'd25885, 16'd59256, 16'd20749, 16'd4388, 16'd61104, 16'd44053, 16'd62289, 16'd2933, 16'd4609, 16'd7391, 16'd16432, 16'd53798, 16'd31673, 16'd61956, 16'd46039, 16'd50227, 16'd19884, 16'd44415, 16'd55916, 16'd57037, 16'd4265});
	test_expansion(128'hd345c35959157c82ffcc0cbde6b78e9f, {16'd18532, 16'd9545, 16'd38006, 16'd21574, 16'd46704, 16'd54519, 16'd32812, 16'd38245, 16'd19061, 16'd49973, 16'd3017, 16'd1338, 16'd50880, 16'd34712, 16'd31289, 16'd41566, 16'd17518, 16'd61671, 16'd15962, 16'd16044, 16'd52496, 16'd14688, 16'd29242, 16'd38106, 16'd53332, 16'd62943});
	test_expansion(128'h7a3967da3a6baadae482d85863ccac8d, {16'd8897, 16'd12689, 16'd13339, 16'd16173, 16'd40919, 16'd62137, 16'd19708, 16'd29422, 16'd19331, 16'd55250, 16'd31219, 16'd45253, 16'd27281, 16'd61652, 16'd52293, 16'd4019, 16'd46590, 16'd40629, 16'd25415, 16'd27975, 16'd40650, 16'd35117, 16'd17002, 16'd4036, 16'd34273, 16'd20188});
	test_expansion(128'h20fc7f4ce598beb654574d9109799588, {16'd12669, 16'd24295, 16'd29102, 16'd27147, 16'd57658, 16'd53944, 16'd50833, 16'd8093, 16'd22520, 16'd29749, 16'd11232, 16'd22367, 16'd44534, 16'd2192, 16'd50075, 16'd50970, 16'd49538, 16'd46818, 16'd36914, 16'd5255, 16'd18685, 16'd9189, 16'd26981, 16'd13072, 16'd40904, 16'd18850});
	test_expansion(128'h45c353a1951ae17a16b047d850054756, {16'd19016, 16'd11972, 16'd36235, 16'd53783, 16'd50136, 16'd61789, 16'd11741, 16'd20289, 16'd25217, 16'd38124, 16'd24485, 16'd39234, 16'd55590, 16'd22723, 16'd22264, 16'd10422, 16'd17143, 16'd731, 16'd55889, 16'd48744, 16'd65092, 16'd33513, 16'd2250, 16'd22371, 16'd6900, 16'd4481});
	test_expansion(128'hde559076217218c779b0a705328d8a16, {16'd1284, 16'd63327, 16'd36847, 16'd30745, 16'd25982, 16'd6904, 16'd41714, 16'd27601, 16'd2558, 16'd34269, 16'd25811, 16'd36713, 16'd2804, 16'd709, 16'd55582, 16'd53657, 16'd12797, 16'd20467, 16'd43564, 16'd51877, 16'd59058, 16'd21436, 16'd50681, 16'd9288, 16'd63008, 16'd1739});
	test_expansion(128'hc87eec59d8a100efdc0c5d3b41d7b854, {16'd37564, 16'd15113, 16'd47902, 16'd37258, 16'd55246, 16'd20485, 16'd39185, 16'd33170, 16'd44292, 16'd10997, 16'd57203, 16'd65438, 16'd42555, 16'd16845, 16'd27199, 16'd4201, 16'd21342, 16'd59365, 16'd33285, 16'd38354, 16'd48167, 16'd40683, 16'd16422, 16'd6563, 16'd31593, 16'd40613});
	test_expansion(128'h31dfa38ab2bfde89323beeb2363b9271, {16'd4697, 16'd16849, 16'd7564, 16'd33357, 16'd22891, 16'd17263, 16'd26721, 16'd17431, 16'd37227, 16'd60849, 16'd7484, 16'd28117, 16'd18884, 16'd9293, 16'd31447, 16'd2924, 16'd26473, 16'd24938, 16'd12053, 16'd49777, 16'd49241, 16'd7426, 16'd12776, 16'd22567, 16'd11862, 16'd59185});
	test_expansion(128'hcdab8ebcef9d26854889c1e9b07caaf5, {16'd29238, 16'd33833, 16'd11071, 16'd52708, 16'd60443, 16'd20062, 16'd3533, 16'd49577, 16'd47785, 16'd45854, 16'd18932, 16'd18585, 16'd63902, 16'd28807, 16'd2873, 16'd59680, 16'd62451, 16'd3104, 16'd25438, 16'd14421, 16'd45173, 16'd1747, 16'd47267, 16'd52945, 16'd45461, 16'd32442});
	test_expansion(128'hcc10a6a8bdc4b1ee0c03fadb5fa5406f, {16'd6102, 16'd49822, 16'd21467, 16'd7987, 16'd38454, 16'd33542, 16'd49312, 16'd11493, 16'd47031, 16'd42235, 16'd9476, 16'd17152, 16'd57201, 16'd56890, 16'd12129, 16'd39713, 16'd57355, 16'd45583, 16'd56134, 16'd3594, 16'd37522, 16'd7285, 16'd8343, 16'd1859, 16'd2833, 16'd5324});
	test_expansion(128'h03cbd5b9e2a330f572b4d30e8de38100, {16'd7089, 16'd49314, 16'd15614, 16'd61648, 16'd55458, 16'd21507, 16'd17527, 16'd891, 16'd34226, 16'd2546, 16'd53637, 16'd974, 16'd20369, 16'd31304, 16'd35467, 16'd3590, 16'd17244, 16'd4930, 16'd49002, 16'd22004, 16'd44355, 16'd1848, 16'd61213, 16'd24472, 16'd54297, 16'd55302});
	test_expansion(128'h2211ef86cf6a565f1d44e860858b0b9c, {16'd36643, 16'd18130, 16'd31714, 16'd8635, 16'd833, 16'd284, 16'd25977, 16'd57474, 16'd13447, 16'd57103, 16'd41904, 16'd42368, 16'd55304, 16'd64588, 16'd29949, 16'd27560, 16'd1800, 16'd2860, 16'd22696, 16'd56253, 16'd41533, 16'd59634, 16'd37599, 16'd19468, 16'd57945, 16'd65201});
	test_expansion(128'h8dbaf9e12851527f31d435d317e59128, {16'd47721, 16'd36642, 16'd9191, 16'd20005, 16'd19969, 16'd28654, 16'd47631, 16'd61653, 16'd23057, 16'd23914, 16'd12945, 16'd19833, 16'd7032, 16'd48046, 16'd42405, 16'd8862, 16'd5440, 16'd31024, 16'd58512, 16'd36990, 16'd52453, 16'd26805, 16'd24040, 16'd46494, 16'd2371, 16'd64060});
	test_expansion(128'hafbfa958ea52406ab5dbe25b3049a58e, {16'd21079, 16'd55849, 16'd1383, 16'd58222, 16'd55646, 16'd24687, 16'd19081, 16'd1831, 16'd2930, 16'd56680, 16'd6124, 16'd49634, 16'd36913, 16'd2232, 16'd49045, 16'd48336, 16'd38600, 16'd5991, 16'd64968, 16'd55179, 16'd45126, 16'd60066, 16'd22201, 16'd31782, 16'd13300, 16'd22085});
	test_expansion(128'h8ccf3c4a4d7596f7ff414bd51f36488d, {16'd48721, 16'd35185, 16'd10967, 16'd11842, 16'd38423, 16'd22175, 16'd61590, 16'd33852, 16'd20880, 16'd61591, 16'd32029, 16'd44239, 16'd27098, 16'd61669, 16'd55457, 16'd33628, 16'd38490, 16'd10610, 16'd31939, 16'd13848, 16'd4189, 16'd65354, 16'd24103, 16'd14417, 16'd12125, 16'd60452});
	test_expansion(128'h9f33ca9ccefd90f28010954cda7d5f39, {16'd46566, 16'd52986, 16'd38306, 16'd41599, 16'd29195, 16'd43395, 16'd10544, 16'd29497, 16'd59934, 16'd3965, 16'd21596, 16'd4837, 16'd2038, 16'd33954, 16'd29921, 16'd14387, 16'd19536, 16'd30489, 16'd37746, 16'd9290, 16'd55954, 16'd1066, 16'd46241, 16'd14707, 16'd27200, 16'd5111});
	test_expansion(128'h5cca438bc9581e72b14173695f6ed200, {16'd35956, 16'd40977, 16'd9680, 16'd54957, 16'd5061, 16'd5637, 16'd23619, 16'd10850, 16'd34416, 16'd23013, 16'd5520, 16'd23273, 16'd45416, 16'd25331, 16'd17951, 16'd7421, 16'd38661, 16'd65053, 16'd49724, 16'd32614, 16'd41035, 16'd721, 16'd48141, 16'd29543, 16'd46451, 16'd23505});
	test_expansion(128'h2d4aed5447b0c67560d9179638e8faeb, {16'd36176, 16'd17515, 16'd691, 16'd61117, 16'd20661, 16'd7824, 16'd56600, 16'd31708, 16'd28030, 16'd65493, 16'd32091, 16'd20801, 16'd54116, 16'd18312, 16'd1290, 16'd10185, 16'd40084, 16'd48472, 16'd39009, 16'd41795, 16'd47228, 16'd53152, 16'd4368, 16'd37261, 16'd18343, 16'd3305});
	test_expansion(128'h546ffdb79a9c18bc649bc16effb8da40, {16'd29612, 16'd44784, 16'd12054, 16'd33422, 16'd15570, 16'd52132, 16'd26066, 16'd50710, 16'd38526, 16'd48116, 16'd32320, 16'd12404, 16'd16226, 16'd23561, 16'd28787, 16'd56408, 16'd29489, 16'd5797, 16'd1546, 16'd60009, 16'd21737, 16'd16551, 16'd20011, 16'd40741, 16'd41360, 16'd3853});
	test_expansion(128'hb645834ed07c3b11bd8cd640f91f22a9, {16'd10369, 16'd59602, 16'd37561, 16'd44704, 16'd24259, 16'd52241, 16'd9297, 16'd24383, 16'd39699, 16'd11341, 16'd7186, 16'd14391, 16'd63098, 16'd46702, 16'd19645, 16'd65329, 16'd43881, 16'd903, 16'd9748, 16'd57065, 16'd49987, 16'd31464, 16'd29569, 16'd530, 16'd64605, 16'd40934});
	test_expansion(128'h53f9a9aaed0084d91fd8524b383630ef, {16'd16537, 16'd60208, 16'd32632, 16'd4662, 16'd30045, 16'd49665, 16'd60490, 16'd16345, 16'd21505, 16'd12327, 16'd32448, 16'd59332, 16'd7204, 16'd50241, 16'd27624, 16'd30889, 16'd46298, 16'd18402, 16'd27643, 16'd22117, 16'd60583, 16'd35414, 16'd46447, 16'd18357, 16'd22904, 16'd31950});
	test_expansion(128'h585cf26513c49edfbc4cb3f5307ecc2b, {16'd24925, 16'd49922, 16'd41189, 16'd10241, 16'd40655, 16'd39445, 16'd35660, 16'd63740, 16'd18974, 16'd56694, 16'd5579, 16'd32970, 16'd22588, 16'd30278, 16'd16389, 16'd9816, 16'd12402, 16'd41476, 16'd35234, 16'd18069, 16'd45158, 16'd10109, 16'd14418, 16'd15187, 16'd22549, 16'd59165});
	test_expansion(128'h4eaf1c538b7d072c3bd6cf9e3741028f, {16'd35405, 16'd59975, 16'd7954, 16'd41864, 16'd55154, 16'd52954, 16'd8126, 16'd8766, 16'd35991, 16'd51474, 16'd6597, 16'd17399, 16'd64915, 16'd65231, 16'd21525, 16'd48178, 16'd16272, 16'd7926, 16'd12955, 16'd44966, 16'd12595, 16'd46044, 16'd36848, 16'd65455, 16'd63067, 16'd31700});
	test_expansion(128'h4e96fdd7b30a54a7a2a9be8b531f84c3, {16'd41998, 16'd45581, 16'd58155, 16'd24477, 16'd41410, 16'd65391, 16'd19999, 16'd48135, 16'd20330, 16'd41376, 16'd17457, 16'd32956, 16'd52780, 16'd36147, 16'd58933, 16'd7078, 16'd1440, 16'd16793, 16'd60725, 16'd61038, 16'd14496, 16'd61137, 16'd55710, 16'd38493, 16'd1890, 16'd38457});
	test_expansion(128'h61b5621c3173018b11b6d46bf07fa5cd, {16'd8508, 16'd28285, 16'd54649, 16'd61047, 16'd26627, 16'd58858, 16'd4246, 16'd32416, 16'd48084, 16'd41318, 16'd56533, 16'd4261, 16'd15309, 16'd329, 16'd20035, 16'd16265, 16'd2506, 16'd2416, 16'd16709, 16'd30987, 16'd11624, 16'd4177, 16'd25408, 16'd25250, 16'd804, 16'd743});
	test_expansion(128'hc967e2a382dc73de619bd17f63be6d95, {16'd11865, 16'd46501, 16'd9936, 16'd53804, 16'd31708, 16'd11756, 16'd27622, 16'd48985, 16'd7498, 16'd994, 16'd65091, 16'd1921, 16'd14753, 16'd61345, 16'd59614, 16'd27392, 16'd31265, 16'd31362, 16'd41439, 16'd31033, 16'd28797, 16'd9967, 16'd50839, 16'd2164, 16'd15519, 16'd3403});
	test_expansion(128'h6ed95574aa983c79faaa567105541b98, {16'd53765, 16'd60333, 16'd16268, 16'd26573, 16'd59210, 16'd14145, 16'd45951, 16'd42919, 16'd9727, 16'd20367, 16'd48022, 16'd48183, 16'd57300, 16'd29190, 16'd9287, 16'd51816, 16'd62276, 16'd38509, 16'd42370, 16'd7401, 16'd64831, 16'd33890, 16'd16141, 16'd23028, 16'd64551, 16'd23869});
	test_expansion(128'h55fcb4f468bb30b62333bc9d1e1e528f, {16'd29434, 16'd31698, 16'd13471, 16'd5781, 16'd56869, 16'd60468, 16'd59438, 16'd16640, 16'd26681, 16'd56454, 16'd53864, 16'd38086, 16'd38146, 16'd62362, 16'd45389, 16'd4623, 16'd44473, 16'd6689, 16'd23562, 16'd57013, 16'd51661, 16'd8697, 16'd55222, 16'd42024, 16'd16446, 16'd3444});
	test_expansion(128'h8bbe651828d32e265b869b3c85162797, {16'd24804, 16'd65083, 16'd38995, 16'd59849, 16'd8965, 16'd20244, 16'd5570, 16'd60467, 16'd60501, 16'd57014, 16'd49076, 16'd30341, 16'd20869, 16'd60058, 16'd53263, 16'd25311, 16'd39649, 16'd53971, 16'd34676, 16'd20476, 16'd7268, 16'd14926, 16'd18582, 16'd44206, 16'd57860, 16'd41682});
	test_expansion(128'hb3c2699468bd538ef7b1dc84b28cfaf6, {16'd56413, 16'd9645, 16'd53084, 16'd42224, 16'd50432, 16'd12303, 16'd61399, 16'd393, 16'd24232, 16'd31129, 16'd38644, 16'd58187, 16'd982, 16'd33948, 16'd52703, 16'd12813, 16'd7617, 16'd14860, 16'd62894, 16'd60117, 16'd3678, 16'd60110, 16'd45754, 16'd13872, 16'd13334, 16'd6093});
	test_expansion(128'h661863471d19ff6d1408d75fc4a4aa08, {16'd39276, 16'd571, 16'd14622, 16'd30443, 16'd5530, 16'd22158, 16'd14446, 16'd20766, 16'd49545, 16'd24455, 16'd10344, 16'd54706, 16'd4502, 16'd13947, 16'd11108, 16'd3727, 16'd28430, 16'd47248, 16'd60684, 16'd46783, 16'd51558, 16'd39325, 16'd19903, 16'd34888, 16'd60972, 16'd22889});
	test_expansion(128'h50d53e4daa7878d4b4984764aaba0298, {16'd21226, 16'd55966, 16'd27562, 16'd11062, 16'd50964, 16'd48840, 16'd25451, 16'd10052, 16'd21544, 16'd31774, 16'd2939, 16'd16099, 16'd40105, 16'd24152, 16'd9900, 16'd11222, 16'd48383, 16'd2330, 16'd51932, 16'd14896, 16'd53000, 16'd60139, 16'd48253, 16'd63742, 16'd15384, 16'd41663});
	test_expansion(128'h78e7b3c21198e544c142d82ecd1c0d60, {16'd52829, 16'd52132, 16'd6626, 16'd27205, 16'd62105, 16'd17268, 16'd40863, 16'd55069, 16'd29910, 16'd41875, 16'd17883, 16'd54336, 16'd62182, 16'd11894, 16'd9879, 16'd48970, 16'd59654, 16'd51319, 16'd18980, 16'd29898, 16'd63248, 16'd13668, 16'd50184, 16'd53887, 16'd40119, 16'd15042});
	test_expansion(128'h66fec6a8f185d318d0deac5f5544b85a, {16'd35606, 16'd11983, 16'd39688, 16'd45726, 16'd55521, 16'd3292, 16'd12833, 16'd60096, 16'd62848, 16'd31854, 16'd37975, 16'd52778, 16'd51734, 16'd30831, 16'd33047, 16'd63644, 16'd5596, 16'd36685, 16'd30014, 16'd44079, 16'd43702, 16'd64540, 16'd273, 16'd25740, 16'd61320, 16'd56251});
	test_expansion(128'h835abbf0c9808b643452dd5892257e4d, {16'd29724, 16'd36063, 16'd33132, 16'd51630, 16'd37124, 16'd20594, 16'd19755, 16'd3876, 16'd41074, 16'd32192, 16'd56448, 16'd5952, 16'd5645, 16'd36069, 16'd42337, 16'd26768, 16'd5847, 16'd4478, 16'd9755, 16'd18955, 16'd30270, 16'd31610, 16'd7088, 16'd44513, 16'd22722, 16'd5147});
	test_expansion(128'h61d0d90b665d1d99e966fd850332c62d, {16'd38766, 16'd5813, 16'd52688, 16'd26259, 16'd44641, 16'd5295, 16'd58506, 16'd1975, 16'd40640, 16'd19184, 16'd32174, 16'd53076, 16'd46283, 16'd8064, 16'd23265, 16'd4955, 16'd58328, 16'd40035, 16'd39156, 16'd35230, 16'd22237, 16'd44592, 16'd36442, 16'd51146, 16'd51442, 16'd31922});
	test_expansion(128'h945d5a2e79da0ab77a898bb1cb4710a7, {16'd5193, 16'd51239, 16'd10805, 16'd38520, 16'd242, 16'd34626, 16'd23605, 16'd36522, 16'd40136, 16'd44818, 16'd28355, 16'd32931, 16'd58752, 16'd51977, 16'd21990, 16'd16945, 16'd33185, 16'd46210, 16'd21813, 16'd53683, 16'd63762, 16'd48366, 16'd37246, 16'd12497, 16'd19751, 16'd3469});
	test_expansion(128'h9a7b54f53456f84385a8144a6046418e, {16'd58771, 16'd39277, 16'd50606, 16'd60353, 16'd1134, 16'd52198, 16'd6156, 16'd3290, 16'd44117, 16'd46514, 16'd57557, 16'd31520, 16'd44515, 16'd11397, 16'd36704, 16'd46733, 16'd21509, 16'd37701, 16'd33260, 16'd23178, 16'd55378, 16'd29776, 16'd62188, 16'd46387, 16'd15210, 16'd49157});
	test_expansion(128'ha14a03c705d1050c12cd832a7079d522, {16'd54468, 16'd4696, 16'd15136, 16'd25354, 16'd3331, 16'd16152, 16'd63175, 16'd24705, 16'd58738, 16'd64500, 16'd27120, 16'd24217, 16'd14155, 16'd61766, 16'd26815, 16'd63045, 16'd36183, 16'd28262, 16'd31409, 16'd45482, 16'd18083, 16'd14477, 16'd8386, 16'd38521, 16'd11819, 16'd61217});
	test_expansion(128'hda574433681d4337ee6f4d7bbf0dba8e, {16'd20018, 16'd52472, 16'd30021, 16'd63697, 16'd4670, 16'd61795, 16'd15301, 16'd45302, 16'd10072, 16'd41630, 16'd57123, 16'd28100, 16'd62950, 16'd43031, 16'd29585, 16'd46571, 16'd62945, 16'd29799, 16'd49607, 16'd11544, 16'd59801, 16'd34240, 16'd5505, 16'd56405, 16'd14938, 16'd13043});
	test_expansion(128'ha1178df6c79e96fc7666614f4c9454c9, {16'd63016, 16'd44915, 16'd34269, 16'd62204, 16'd21342, 16'd22707, 16'd26431, 16'd46494, 16'd58405, 16'd29442, 16'd6985, 16'd37110, 16'd52705, 16'd65242, 16'd14125, 16'd39179, 16'd55525, 16'd26743, 16'd33921, 16'd10987, 16'd63886, 16'd2629, 16'd60998, 16'd28607, 16'd35138, 16'd23438});
	test_expansion(128'hdb52bdfc69ba77bd24e1e855b438557e, {16'd10873, 16'd5358, 16'd26735, 16'd594, 16'd22084, 16'd725, 16'd42275, 16'd1100, 16'd60461, 16'd24086, 16'd61251, 16'd38664, 16'd1587, 16'd58171, 16'd59490, 16'd52631, 16'd4510, 16'd44737, 16'd15795, 16'd9247, 16'd40356, 16'd38384, 16'd23682, 16'd1351, 16'd31121, 16'd42570});
	test_expansion(128'h0582b0ebe79ed96b7089ecd4e36d5bae, {16'd11484, 16'd39126, 16'd46386, 16'd1186, 16'd38051, 16'd37145, 16'd62905, 16'd52059, 16'd48813, 16'd10747, 16'd63326, 16'd42550, 16'd14389, 16'd2932, 16'd8484, 16'd42297, 16'd15447, 16'd52610, 16'd1636, 16'd55308, 16'd62604, 16'd9221, 16'd27939, 16'd5213, 16'd51492, 16'd54889});
	test_expansion(128'had08f2f7902e3fb082248092960295bc, {16'd15587, 16'd22703, 16'd11586, 16'd24522, 16'd31244, 16'd6690, 16'd56627, 16'd43076, 16'd37983, 16'd33704, 16'd27546, 16'd12054, 16'd64383, 16'd15023, 16'd34690, 16'd14807, 16'd37164, 16'd37433, 16'd33, 16'd32862, 16'd26916, 16'd29092, 16'd31894, 16'd37732, 16'd7850, 16'd29443});
	test_expansion(128'he151e66b92d8157240774d63c82222ff, {16'd1542, 16'd28889, 16'd34207, 16'd45936, 16'd53021, 16'd64357, 16'd44187, 16'd23005, 16'd63362, 16'd64627, 16'd27601, 16'd62066, 16'd37958, 16'd59453, 16'd8938, 16'd472, 16'd14640, 16'd12791, 16'd51509, 16'd40118, 16'd50395, 16'd44810, 16'd20892, 16'd158, 16'd51379, 16'd58810});
	test_expansion(128'ha2af5b6e0e9f95cb4661e615e78ed2f8, {16'd1798, 16'd23052, 16'd28412, 16'd49571, 16'd40606, 16'd26269, 16'd2965, 16'd58314, 16'd30827, 16'd62055, 16'd64528, 16'd13168, 16'd52933, 16'd6918, 16'd24833, 16'd5330, 16'd84, 16'd35023, 16'd31430, 16'd25608, 16'd53617, 16'd46629, 16'd48398, 16'd44173, 16'd4463, 16'd7111});
	test_expansion(128'h1ed415d36f10436af8efa00c12b5e8fe, {16'd32895, 16'd33845, 16'd64151, 16'd29631, 16'd4605, 16'd50587, 16'd26306, 16'd52275, 16'd65533, 16'd42835, 16'd63587, 16'd35771, 16'd64948, 16'd43535, 16'd17630, 16'd63930, 16'd8357, 16'd59524, 16'd60217, 16'd61377, 16'd20513, 16'd25701, 16'd59276, 16'd26256, 16'd8948, 16'd30135});
	test_expansion(128'h743680791e4f41d4c8636f1b1d023b96, {16'd58163, 16'd43389, 16'd31686, 16'd10857, 16'd37942, 16'd27596, 16'd24179, 16'd35193, 16'd54465, 16'd21668, 16'd55492, 16'd2724, 16'd3298, 16'd59230, 16'd7273, 16'd27322, 16'd64958, 16'd50141, 16'd56516, 16'd47844, 16'd9167, 16'd27317, 16'd64552, 16'd13037, 16'd49879, 16'd27065});
	test_expansion(128'hedf41135878a723220c77ca3d72802a2, {16'd57828, 16'd37826, 16'd60058, 16'd29537, 16'd55199, 16'd67, 16'd15039, 16'd4287, 16'd32834, 16'd11559, 16'd1282, 16'd40153, 16'd7416, 16'd26722, 16'd8138, 16'd57214, 16'd12632, 16'd61573, 16'd12494, 16'd59240, 16'd42503, 16'd49281, 16'd25059, 16'd54437, 16'd15888, 16'd6338});
	test_expansion(128'h66d8692027f5a484532967cf57afb1c1, {16'd46760, 16'd24473, 16'd40290, 16'd17248, 16'd51787, 16'd1691, 16'd22950, 16'd3866, 16'd55043, 16'd40094, 16'd54508, 16'd53807, 16'd36444, 16'd50271, 16'd64339, 16'd56962, 16'd46061, 16'd17222, 16'd62013, 16'd64934, 16'd22358, 16'd49019, 16'd59979, 16'd34425, 16'd17381, 16'd19663});
	test_expansion(128'h9be7ea7881cd251ce12ed702cd1411cb, {16'd65213, 16'd15833, 16'd64657, 16'd40866, 16'd32163, 16'd6097, 16'd46266, 16'd6061, 16'd55350, 16'd15297, 16'd48803, 16'd2954, 16'd65175, 16'd21840, 16'd40096, 16'd23861, 16'd56700, 16'd38460, 16'd43897, 16'd6121, 16'd50182, 16'd35527, 16'd20124, 16'd1713, 16'd54394, 16'd42500});
	test_expansion(128'hd4cd8dfc6e3ffb541d02fa0d2c9ebf96, {16'd21697, 16'd17088, 16'd8052, 16'd55959, 16'd62770, 16'd46755, 16'd61145, 16'd64607, 16'd12653, 16'd39052, 16'd13116, 16'd15754, 16'd46620, 16'd54967, 16'd31507, 16'd43148, 16'd40704, 16'd39350, 16'd27954, 16'd51298, 16'd62022, 16'd4532, 16'd23151, 16'd22248, 16'd28267, 16'd36478});
	test_expansion(128'h657903785cc5c7fdfdaca9bc498cd254, {16'd7481, 16'd26350, 16'd5950, 16'd34316, 16'd53939, 16'd47412, 16'd47461, 16'd42052, 16'd62779, 16'd47438, 16'd38089, 16'd12715, 16'd21098, 16'd39184, 16'd59491, 16'd2720, 16'd54052, 16'd17014, 16'd28924, 16'd34090, 16'd6000, 16'd3502, 16'd11578, 16'd28038, 16'd52527, 16'd57110});
	test_expansion(128'h1088cfcd892b3af203d7ddcfd3da9d1e, {16'd52698, 16'd35366, 16'd52801, 16'd61992, 16'd61086, 16'd48815, 16'd49038, 16'd51788, 16'd61075, 16'd9739, 16'd24494, 16'd39811, 16'd56355, 16'd37823, 16'd38312, 16'd55850, 16'd44757, 16'd52261, 16'd56841, 16'd63186, 16'd32832, 16'd51040, 16'd39755, 16'd52889, 16'd1281, 16'd16476});
	test_expansion(128'h0f24595142ea406d2d87ef2f3fbd42bc, {16'd61168, 16'd30751, 16'd22962, 16'd11999, 16'd59263, 16'd30395, 16'd48059, 16'd60345, 16'd14842, 16'd58392, 16'd17321, 16'd56782, 16'd26229, 16'd24890, 16'd59870, 16'd53966, 16'd19990, 16'd41128, 16'd54439, 16'd29983, 16'd39448, 16'd44232, 16'd20216, 16'd60090, 16'd51549, 16'd16938});
	test_expansion(128'h233e4090984e434d0d0efd951d09af2b, {16'd47014, 16'd13314, 16'd10825, 16'd37376, 16'd1889, 16'd49322, 16'd52151, 16'd6205, 16'd62012, 16'd47621, 16'd46577, 16'd39616, 16'd53691, 16'd65039, 16'd29321, 16'd65495, 16'd52909, 16'd41886, 16'd27935, 16'd33077, 16'd27494, 16'd63916, 16'd19580, 16'd21325, 16'd40244, 16'd26260});
	test_expansion(128'h37d0088df26ec76f733aa0b7be4013c6, {16'd19922, 16'd61134, 16'd58666, 16'd4712, 16'd7395, 16'd61294, 16'd31666, 16'd28722, 16'd18603, 16'd44004, 16'd21646, 16'd60019, 16'd37273, 16'd3875, 16'd45430, 16'd18510, 16'd49818, 16'd50449, 16'd18423, 16'd53314, 16'd30573, 16'd28064, 16'd36675, 16'd53516, 16'd14410, 16'd13979});
	test_expansion(128'h02869177c8ebda94211a0092750a5571, {16'd49919, 16'd38458, 16'd21382, 16'd13629, 16'd29462, 16'd57120, 16'd51350, 16'd53368, 16'd60361, 16'd29070, 16'd36449, 16'd60966, 16'd26050, 16'd27677, 16'd17322, 16'd64179, 16'd32389, 16'd40843, 16'd65371, 16'd21627, 16'd179, 16'd55666, 16'd51679, 16'd14450, 16'd41187, 16'd39753});
	test_expansion(128'hb87ae1b57e941c5f39721b3381cd1878, {16'd15941, 16'd7724, 16'd55980, 16'd2426, 16'd62088, 16'd24919, 16'd2322, 16'd50551, 16'd15952, 16'd12570, 16'd51228, 16'd10500, 16'd9151, 16'd49518, 16'd871, 16'd10351, 16'd22895, 16'd61167, 16'd47361, 16'd36341, 16'd6490, 16'd41336, 16'd10700, 16'd8032, 16'd44729, 16'd43795});
	test_expansion(128'hb3ca1e26494227787fbaba65654b7115, {16'd2924, 16'd55809, 16'd15949, 16'd20931, 16'd8325, 16'd22415, 16'd23794, 16'd14063, 16'd5566, 16'd7069, 16'd37976, 16'd57069, 16'd29785, 16'd25341, 16'd50218, 16'd49528, 16'd44450, 16'd62098, 16'd17982, 16'd55250, 16'd28400, 16'd59247, 16'd18944, 16'd25475, 16'd18583, 16'd15313});
	test_expansion(128'ha3972c615dc035539115fe52d79b6bfd, {16'd12343, 16'd51075, 16'd26970, 16'd48712, 16'd51436, 16'd991, 16'd59596, 16'd33565, 16'd6690, 16'd50031, 16'd53641, 16'd25704, 16'd47942, 16'd19142, 16'd43642, 16'd46951, 16'd20982, 16'd31268, 16'd46734, 16'd20934, 16'd52344, 16'd2797, 16'd4004, 16'd59603, 16'd28274, 16'd47607});
	test_expansion(128'h3d661bb1eaaf1b06e21d9677c98bf8a5, {16'd57570, 16'd43382, 16'd40811, 16'd46686, 16'd33057, 16'd64733, 16'd819, 16'd29173, 16'd1910, 16'd63305, 16'd16340, 16'd43205, 16'd57949, 16'd27223, 16'd44500, 16'd11186, 16'd7265, 16'd31309, 16'd520, 16'd52136, 16'd2063, 16'd39271, 16'd15980, 16'd15983, 16'd1844, 16'd22509});
	test_expansion(128'ha3a5567f370a454f8b32b2a4420c8c4f, {16'd64799, 16'd9536, 16'd7732, 16'd21335, 16'd1232, 16'd31506, 16'd4004, 16'd33837, 16'd23136, 16'd52551, 16'd47053, 16'd4901, 16'd54710, 16'd50354, 16'd34661, 16'd8933, 16'd26694, 16'd32101, 16'd64071, 16'd44265, 16'd25171, 16'd27788, 16'd14641, 16'd53699, 16'd34780, 16'd52486});
	test_expansion(128'ha52c51bc9d21b773656c32266ef5aa9a, {16'd57430, 16'd9959, 16'd31036, 16'd31346, 16'd40806, 16'd41100, 16'd21536, 16'd37563, 16'd38764, 16'd26062, 16'd30024, 16'd21325, 16'd21, 16'd26513, 16'd22973, 16'd11424, 16'd23810, 16'd64788, 16'd33958, 16'd12302, 16'd17034, 16'd48794, 16'd50265, 16'd59720, 16'd64930, 16'd55121});
	test_expansion(128'h02626d9550e11089eb89cf765cdbdaed, {16'd56600, 16'd48148, 16'd64438, 16'd61933, 16'd14399, 16'd18571, 16'd56875, 16'd30661, 16'd36440, 16'd41244, 16'd41592, 16'd31986, 16'd61872, 16'd9512, 16'd39322, 16'd27719, 16'd13006, 16'd57310, 16'd46113, 16'd47000, 16'd57989, 16'd30586, 16'd37600, 16'd24101, 16'd60151, 16'd52961});
	test_expansion(128'h48d61e864d9908b7d7bff533ba76348f, {16'd9754, 16'd58102, 16'd14516, 16'd50488, 16'd27990, 16'd15539, 16'd4752, 16'd32279, 16'd5683, 16'd16056, 16'd2065, 16'd26917, 16'd20160, 16'd8067, 16'd47492, 16'd59225, 16'd23366, 16'd19740, 16'd21350, 16'd58429, 16'd3183, 16'd29436, 16'd42543, 16'd28192, 16'd20221, 16'd41211});
	test_expansion(128'h7a127f4da31a2fd66f1d0d226c0f9beb, {16'd34293, 16'd52941, 16'd3519, 16'd50161, 16'd37875, 16'd28330, 16'd572, 16'd28252, 16'd5814, 16'd44343, 16'd27713, 16'd63595, 16'd34403, 16'd26743, 16'd55627, 16'd10236, 16'd51413, 16'd55905, 16'd13972, 16'd48181, 16'd24679, 16'd7502, 16'd35203, 16'd57908, 16'd58668, 16'd31049});
	test_expansion(128'hf320cf8df3762c3e30e7a47d2a76a5af, {16'd15701, 16'd39339, 16'd40451, 16'd3468, 16'd43210, 16'd44009, 16'd45978, 16'd15544, 16'd18293, 16'd37633, 16'd47594, 16'd27901, 16'd20260, 16'd38575, 16'd38654, 16'd32016, 16'd23131, 16'd30017, 16'd46336, 16'd9669, 16'd12357, 16'd17899, 16'd16010, 16'd13066, 16'd35674, 16'd4100});
	test_expansion(128'ha60874d29f7745f1701cbbeea28166b5, {16'd35529, 16'd6514, 16'd34336, 16'd26732, 16'd21178, 16'd63602, 16'd28414, 16'd42506, 16'd3411, 16'd61802, 16'd24860, 16'd62017, 16'd19735, 16'd52658, 16'd64565, 16'd17875, 16'd58246, 16'd33775, 16'd32114, 16'd8565, 16'd62310, 16'd18605, 16'd26779, 16'd31801, 16'd47533, 16'd37180});
	test_expansion(128'h756163f4b0bf2adbff5975bebfe341ea, {16'd55209, 16'd60548, 16'd33614, 16'd58258, 16'd18263, 16'd14474, 16'd34126, 16'd392, 16'd24816, 16'd28453, 16'd479, 16'd38876, 16'd17855, 16'd11639, 16'd10776, 16'd62474, 16'd30886, 16'd53980, 16'd24571, 16'd17385, 16'd42356, 16'd26407, 16'd49303, 16'd36704, 16'd60951, 16'd10702});
	test_expansion(128'ha1806bda2f5cbe442b5914acf2ad2f53, {16'd55128, 16'd63674, 16'd2817, 16'd28896, 16'd36745, 16'd62762, 16'd10524, 16'd62732, 16'd58799, 16'd36640, 16'd26360, 16'd47559, 16'd2894, 16'd57651, 16'd55542, 16'd42287, 16'd19962, 16'd51563, 16'd49420, 16'd56573, 16'd17857, 16'd33086, 16'd43444, 16'd9425, 16'd50799, 16'd46502});
	test_expansion(128'he0c947879e735956f43f4607c33b6026, {16'd36391, 16'd17805, 16'd47051, 16'd9757, 16'd1889, 16'd36759, 16'd41113, 16'd36634, 16'd49314, 16'd624, 16'd35549, 16'd32575, 16'd23875, 16'd50284, 16'd25659, 16'd26132, 16'd53610, 16'd861, 16'd5340, 16'd14359, 16'd47813, 16'd34139, 16'd29925, 16'd1089, 16'd34269, 16'd33342});
	test_expansion(128'h7118a5e8caac6d7709502b1f3c5526c3, {16'd16914, 16'd44110, 16'd8680, 16'd30904, 16'd52553, 16'd47542, 16'd61498, 16'd61934, 16'd65035, 16'd5161, 16'd36241, 16'd6858, 16'd46507, 16'd30185, 16'd65522, 16'd43816, 16'd27756, 16'd54039, 16'd26365, 16'd30522, 16'd25825, 16'd56006, 16'd46138, 16'd3001, 16'd61674, 16'd31568});
	test_expansion(128'h6b5e6be3f0f4b30963d99c17a7018e35, {16'd56033, 16'd60187, 16'd12006, 16'd30130, 16'd17019, 16'd58019, 16'd22277, 16'd23712, 16'd60744, 16'd64307, 16'd10284, 16'd44858, 16'd1578, 16'd32693, 16'd64690, 16'd10190, 16'd35752, 16'd1105, 16'd59728, 16'd65329, 16'd6770, 16'd20357, 16'd342, 16'd410, 16'd15503, 16'd55513});
	test_expansion(128'hc8db3b563ca7d1a4e2a7189a1b5dde13, {16'd2152, 16'd47515, 16'd29665, 16'd49353, 16'd15484, 16'd24135, 16'd54813, 16'd9596, 16'd6497, 16'd29672, 16'd8336, 16'd13832, 16'd51697, 16'd45758, 16'd53019, 16'd53050, 16'd45714, 16'd49887, 16'd59945, 16'd53314, 16'd58582, 16'd17902, 16'd29198, 16'd21589, 16'd44555, 16'd22561});
	test_expansion(128'h6f028a37d530118df108feba01e01857, {16'd29093, 16'd24913, 16'd9145, 16'd12075, 16'd38490, 16'd51539, 16'd20991, 16'd16888, 16'd37833, 16'd41145, 16'd15594, 16'd60123, 16'd37423, 16'd40118, 16'd17075, 16'd47004, 16'd15094, 16'd13460, 16'd24951, 16'd62046, 16'd12155, 16'd41233, 16'd18513, 16'd24588, 16'd27590, 16'd53374});
	test_expansion(128'he19e492548f1283735c4a25133b0b869, {16'd20462, 16'd51806, 16'd6552, 16'd51402, 16'd45108, 16'd54345, 16'd54060, 16'd40206, 16'd23382, 16'd65226, 16'd50286, 16'd728, 16'd47770, 16'd13761, 16'd44121, 16'd44205, 16'd43298, 16'd51136, 16'd13754, 16'd28270, 16'd27777, 16'd56683, 16'd32679, 16'd48769, 16'd44856, 16'd1338});
	test_expansion(128'hf336aabed9902d045e73880342422085, {16'd50199, 16'd28393, 16'd15285, 16'd8283, 16'd23913, 16'd57552, 16'd1228, 16'd7847, 16'd51943, 16'd41196, 16'd35251, 16'd53917, 16'd51024, 16'd45073, 16'd60303, 16'd33790, 16'd58638, 16'd44123, 16'd30742, 16'd43817, 16'd35366, 16'd15491, 16'd2752, 16'd57948, 16'd50939, 16'd13340});
	test_expansion(128'ha5335b58a817408cec8dde7df78bbe11, {16'd13083, 16'd22461, 16'd31696, 16'd55527, 16'd39903, 16'd62984, 16'd5205, 16'd37441, 16'd40473, 16'd20821, 16'd34318, 16'd35526, 16'd43749, 16'd28357, 16'd56441, 16'd54260, 16'd4795, 16'd25651, 16'd44556, 16'd55228, 16'd52974, 16'd16863, 16'd49768, 16'd59251, 16'd7404, 16'd20971});
	test_expansion(128'h867b5a5b782d2a18fde2ffbcd491dfb5, {16'd9925, 16'd41698, 16'd47098, 16'd2844, 16'd47502, 16'd30439, 16'd42875, 16'd57928, 16'd13060, 16'd46423, 16'd34416, 16'd59741, 16'd50046, 16'd31566, 16'd65406, 16'd45865, 16'd51760, 16'd27943, 16'd44539, 16'd55981, 16'd17656, 16'd33195, 16'd10671, 16'd24070, 16'd3700, 16'd37702});
	test_expansion(128'h7cdcde91536f47a5294294e7b060daec, {16'd20469, 16'd52298, 16'd10804, 16'd56224, 16'd31907, 16'd15948, 16'd29778, 16'd36152, 16'd57281, 16'd6526, 16'd57095, 16'd59127, 16'd10761, 16'd56459, 16'd39506, 16'd15480, 16'd43869, 16'd65281, 16'd11324, 16'd5131, 16'd39991, 16'd25375, 16'd45608, 16'd6270, 16'd54513, 16'd3149});
	test_expansion(128'he00a35486d5a949e1a53610a06de2588, {16'd47216, 16'd46264, 16'd34037, 16'd44155, 16'd39718, 16'd32491, 16'd58305, 16'd4145, 16'd40423, 16'd44487, 16'd32407, 16'd38106, 16'd12089, 16'd12781, 16'd60599, 16'd9071, 16'd47143, 16'd7278, 16'd33648, 16'd34698, 16'd52906, 16'd26808, 16'd30111, 16'd8184, 16'd18745, 16'd13306});
	test_expansion(128'h64b8f1bec2b6708e1eb2beed7283f9b3, {16'd2067, 16'd51421, 16'd32615, 16'd61094, 16'd64695, 16'd52413, 16'd62867, 16'd19197, 16'd42451, 16'd51360, 16'd9381, 16'd24476, 16'd2203, 16'd27921, 16'd25813, 16'd7563, 16'd32063, 16'd64679, 16'd36675, 16'd41960, 16'd38348, 16'd45033, 16'd53694, 16'd3243, 16'd11410, 16'd43020});
	test_expansion(128'h7cdbcfd0cdc1c0cc482c73cdd0ee20ca, {16'd53122, 16'd32156, 16'd42931, 16'd60214, 16'd41352, 16'd56408, 16'd46413, 16'd15979, 16'd23035, 16'd57497, 16'd19173, 16'd18523, 16'd16415, 16'd46202, 16'd9916, 16'd19361, 16'd60279, 16'd62296, 16'd56722, 16'd28687, 16'd4196, 16'd25648, 16'd8842, 16'd61721, 16'd15541, 16'd51235});
	test_expansion(128'h96547f7224475da05eee9f5021c514f4, {16'd7759, 16'd13145, 16'd38238, 16'd48777, 16'd39779, 16'd25617, 16'd57454, 16'd37495, 16'd18473, 16'd39111, 16'd45112, 16'd63604, 16'd4908, 16'd55001, 16'd62849, 16'd7604, 16'd64650, 16'd45910, 16'd9690, 16'd46753, 16'd62100, 16'd20407, 16'd55542, 16'd44994, 16'd2959, 16'd10507});
	test_expansion(128'hf3a84641f866fbef4c521ba4c3a0798b, {16'd43755, 16'd65217, 16'd24731, 16'd28541, 16'd10996, 16'd53373, 16'd43394, 16'd44131, 16'd42607, 16'd6984, 16'd63039, 16'd1444, 16'd58061, 16'd45747, 16'd39089, 16'd63826, 16'd39365, 16'd42931, 16'd39967, 16'd25664, 16'd20317, 16'd7020, 16'd54041, 16'd53238, 16'd22414, 16'd2136});
	test_expansion(128'h7d95973eae0e9774d513f6cf3455f852, {16'd47503, 16'd13977, 16'd15106, 16'd49233, 16'd63852, 16'd48997, 16'd52066, 16'd31989, 16'd43356, 16'd45506, 16'd58217, 16'd45357, 16'd34460, 16'd6586, 16'd46937, 16'd30344, 16'd55752, 16'd11338, 16'd1450, 16'd13194, 16'd38776, 16'd10785, 16'd46035, 16'd8899, 16'd53037, 16'd36669});
	test_expansion(128'he35cf5200fc651bbdb4656482f28c969, {16'd4036, 16'd61621, 16'd42775, 16'd43045, 16'd31393, 16'd46420, 16'd6268, 16'd47000, 16'd3290, 16'd35281, 16'd26464, 16'd21641, 16'd28344, 16'd60324, 16'd34846, 16'd64407, 16'd31833, 16'd13658, 16'd49254, 16'd32826, 16'd38688, 16'd6138, 16'd15732, 16'd4064, 16'd46022, 16'd25710});
	test_expansion(128'h7901fe59ada7316a9948fe4b51abd550, {16'd13484, 16'd27058, 16'd35489, 16'd30556, 16'd24399, 16'd22213, 16'd44292, 16'd54274, 16'd53145, 16'd40118, 16'd27243, 16'd41603, 16'd4620, 16'd62874, 16'd45724, 16'd16883, 16'd43506, 16'd9998, 16'd20559, 16'd64331, 16'd19641, 16'd9914, 16'd40572, 16'd62339, 16'd11830, 16'd43752});
	test_expansion(128'h3f0e74e6f8e4cf23424916f84a448397, {16'd58371, 16'd51947, 16'd31477, 16'd14272, 16'd31622, 16'd52880, 16'd15766, 16'd56356, 16'd58076, 16'd63611, 16'd57252, 16'd17645, 16'd61353, 16'd5604, 16'd31297, 16'd24798, 16'd39977, 16'd2410, 16'd22394, 16'd10996, 16'd24878, 16'd21361, 16'd21509, 16'd23134, 16'd50199, 16'd39945});
	test_expansion(128'h3783b411b5ad710adc45feb6b709b9b8, {16'd59364, 16'd57217, 16'd61885, 16'd846, 16'd44716, 16'd37770, 16'd31852, 16'd58330, 16'd2885, 16'd45941, 16'd61045, 16'd16814, 16'd20828, 16'd3139, 16'd43424, 16'd34880, 16'd34329, 16'd20413, 16'd815, 16'd49352, 16'd25438, 16'd10919, 16'd10938, 16'd10324, 16'd18885, 16'd38242});
	test_expansion(128'h25ac2d010fb34699cd13c652d28fc994, {16'd62940, 16'd7930, 16'd52139, 16'd11480, 16'd42198, 16'd27824, 16'd23965, 16'd58512, 16'd9891, 16'd5268, 16'd39601, 16'd3087, 16'd48470, 16'd65027, 16'd16254, 16'd61312, 16'd21997, 16'd24068, 16'd41957, 16'd28997, 16'd31601, 16'd22644, 16'd63816, 16'd56622, 16'd65513, 16'd40481});
	test_expansion(128'h4e3725132d30758f4a191a75ce9af03c, {16'd12084, 16'd33450, 16'd17664, 16'd11424, 16'd39588, 16'd5997, 16'd5430, 16'd26947, 16'd28957, 16'd51395, 16'd19033, 16'd25081, 16'd38813, 16'd32648, 16'd25314, 16'd61963, 16'd5954, 16'd45475, 16'd17389, 16'd36849, 16'd40960, 16'd62574, 16'd51871, 16'd57524, 16'd21167, 16'd21698});
	test_expansion(128'h6d92ac08bce037e962188b8c0b569a39, {16'd24149, 16'd15326, 16'd62908, 16'd32787, 16'd51148, 16'd21846, 16'd8720, 16'd16849, 16'd30170, 16'd19130, 16'd12801, 16'd55988, 16'd21215, 16'd52086, 16'd41846, 16'd33879, 16'd24026, 16'd36113, 16'd45804, 16'd48116, 16'd24118, 16'd31635, 16'd46758, 16'd58841, 16'd25242, 16'd24310});
	test_expansion(128'h7344e32cc475de0451facf693c91346d, {16'd49677, 16'd48942, 16'd42652, 16'd11060, 16'd8155, 16'd41563, 16'd38643, 16'd28475, 16'd28273, 16'd36807, 16'd42080, 16'd49864, 16'd24289, 16'd56541, 16'd15274, 16'd7484, 16'd16920, 16'd5897, 16'd38317, 16'd25025, 16'd12290, 16'd27784, 16'd5618, 16'd50758, 16'd25435, 16'd58993});
	test_expansion(128'hbe48443fb4eb644a975404ea4a76b381, {16'd45530, 16'd61349, 16'd4558, 16'd13778, 16'd55170, 16'd8079, 16'd46311, 16'd9847, 16'd6543, 16'd7766, 16'd48535, 16'd33284, 16'd43660, 16'd56, 16'd52816, 16'd20514, 16'd57702, 16'd61172, 16'd61450, 16'd37530, 16'd20067, 16'd62123, 16'd42119, 16'd45689, 16'd61631, 16'd51557});
	test_expansion(128'h610a60163d5356eb8e2b61bd85695ad7, {16'd40571, 16'd18786, 16'd19427, 16'd27533, 16'd10194, 16'd958, 16'd40162, 16'd43397, 16'd65174, 16'd19847, 16'd35369, 16'd33854, 16'd21015, 16'd32834, 16'd5771, 16'd10020, 16'd15695, 16'd54263, 16'd40173, 16'd52245, 16'd57419, 16'd38456, 16'd65046, 16'd19326, 16'd7560, 16'd12224});
	test_expansion(128'h245067e94f35808a4e6f3b08fa0e3112, {16'd29707, 16'd49004, 16'd23303, 16'd9259, 16'd34457, 16'd37735, 16'd56304, 16'd18765, 16'd33713, 16'd29212, 16'd31167, 16'd51167, 16'd35174, 16'd24122, 16'd61806, 16'd6794, 16'd27242, 16'd12852, 16'd184, 16'd3049, 16'd21427, 16'd24627, 16'd34958, 16'd23358, 16'd60662, 16'd54802});
	test_expansion(128'hb82f42bb5eca8d92af81399ceb832767, {16'd23230, 16'd46556, 16'd52955, 16'd288, 16'd53741, 16'd41752, 16'd62619, 16'd56592, 16'd45317, 16'd29300, 16'd34507, 16'd15386, 16'd27014, 16'd20358, 16'd1820, 16'd6197, 16'd60988, 16'd37288, 16'd64793, 16'd17466, 16'd27050, 16'd25605, 16'd34002, 16'd51798, 16'd13464, 16'd8727});
	test_expansion(128'h1fd56b7f9f2178b8907acb7dccc8af0e, {16'd55580, 16'd56819, 16'd38175, 16'd63815, 16'd23671, 16'd31433, 16'd29745, 16'd33853, 16'd63284, 16'd31859, 16'd30858, 16'd57522, 16'd46971, 16'd29614, 16'd8628, 16'd62544, 16'd32236, 16'd29035, 16'd5929, 16'd47257, 16'd27100, 16'd2103, 16'd63992, 16'd39268, 16'd15247, 16'd46244});
	test_expansion(128'h277d377a1100d862dda85b80943e8eec, {16'd48012, 16'd6066, 16'd6824, 16'd24158, 16'd58194, 16'd25112, 16'd10131, 16'd2543, 16'd40176, 16'd39648, 16'd61268, 16'd17208, 16'd24543, 16'd15894, 16'd30481, 16'd32449, 16'd19590, 16'd1878, 16'd42274, 16'd61090, 16'd26093, 16'd13225, 16'd52987, 16'd32024, 16'd3762, 16'd40588});
	test_expansion(128'h5fef44a4a4deaf78c8978e2dbd65b69e, {16'd18901, 16'd32776, 16'd46645, 16'd51945, 16'd60308, 16'd42872, 16'd34008, 16'd34988, 16'd31810, 16'd52865, 16'd41984, 16'd20277, 16'd12776, 16'd56958, 16'd14966, 16'd6141, 16'd36988, 16'd1736, 16'd28198, 16'd34028, 16'd26163, 16'd40346, 16'd27771, 16'd42482, 16'd42747, 16'd21336});
	test_expansion(128'h67a50a4b4a6d3dd97c54809cabe44302, {16'd55853, 16'd61056, 16'd11411, 16'd51924, 16'd45341, 16'd34292, 16'd42591, 16'd21348, 16'd45961, 16'd57651, 16'd32873, 16'd4324, 16'd41394, 16'd23910, 16'd7912, 16'd18704, 16'd48080, 16'd51151, 16'd3652, 16'd58703, 16'd2570, 16'd35066, 16'd18423, 16'd36988, 16'd48186, 16'd56442});
	test_expansion(128'h7d666bdb0790743539b16e3f0b8b7e9a, {16'd21133, 16'd7811, 16'd36761, 16'd65168, 16'd25316, 16'd27694, 16'd62452, 16'd13948, 16'd41879, 16'd35455, 16'd56058, 16'd1201, 16'd41005, 16'd57872, 16'd50416, 16'd42346, 16'd3933, 16'd64503, 16'd8471, 16'd46770, 16'd64249, 16'd1870, 16'd16265, 16'd4700, 16'd3118, 16'd18302});
	test_expansion(128'h6a55b3bd8cfb46583b558e6aa627a833, {16'd38511, 16'd42403, 16'd60131, 16'd45021, 16'd49446, 16'd58565, 16'd25280, 16'd38997, 16'd7406, 16'd35286, 16'd25808, 16'd43463, 16'd38664, 16'd38293, 16'd56368, 16'd41542, 16'd47079, 16'd40378, 16'd39175, 16'd49112, 16'd46989, 16'd41209, 16'd59840, 16'd58710, 16'd13427, 16'd31930});
	test_expansion(128'h661ad49b241fd4ef67e2127c0c7025ab, {16'd9603, 16'd62176, 16'd36116, 16'd62752, 16'd998, 16'd62634, 16'd46200, 16'd6052, 16'd48804, 16'd38378, 16'd48938, 16'd45771, 16'd20401, 16'd31454, 16'd20091, 16'd42964, 16'd48450, 16'd36573, 16'd65011, 16'd55539, 16'd34274, 16'd38527, 16'd10610, 16'd21720, 16'd12548, 16'd56529});
	test_expansion(128'hea8c56ccde8be49ef781698a97328a94, {16'd42615, 16'd62475, 16'd39429, 16'd42879, 16'd49136, 16'd26340, 16'd53813, 16'd17634, 16'd23418, 16'd46059, 16'd56582, 16'd48236, 16'd12043, 16'd53845, 16'd773, 16'd52437, 16'd44021, 16'd50082, 16'd56818, 16'd31809, 16'd43311, 16'd64804, 16'd10323, 16'd14412, 16'd46584, 16'd5000});
	test_expansion(128'hbf496a708c8ab963f97fcc6771e75d79, {16'd39641, 16'd63917, 16'd44623, 16'd47021, 16'd9719, 16'd44013, 16'd44069, 16'd44571, 16'd48621, 16'd35590, 16'd61617, 16'd61661, 16'd50846, 16'd26289, 16'd56492, 16'd6656, 16'd30842, 16'd29414, 16'd29601, 16'd2442, 16'd589, 16'd13789, 16'd24365, 16'd12785, 16'd16617, 16'd36384});
	test_expansion(128'h539f46187948d7e0147ab25689a342bf, {16'd64987, 16'd65196, 16'd50837, 16'd15445, 16'd49001, 16'd16714, 16'd40138, 16'd61585, 16'd38088, 16'd63960, 16'd63599, 16'd41324, 16'd24263, 16'd27891, 16'd52407, 16'd54305, 16'd50251, 16'd54438, 16'd56556, 16'd33908, 16'd51527, 16'd46362, 16'd6655, 16'd11675, 16'd50214, 16'd1697});
	test_expansion(128'hc6b684ebe75a73e6268515efbdeea727, {16'd63256, 16'd27641, 16'd57669, 16'd44540, 16'd49693, 16'd51550, 16'd6252, 16'd51635, 16'd53782, 16'd6595, 16'd50370, 16'd12033, 16'd18924, 16'd37954, 16'd3854, 16'd5052, 16'd9453, 16'd41372, 16'd25202, 16'd51211, 16'd52714, 16'd9298, 16'd30617, 16'd47483, 16'd42600, 16'd7549});
	test_expansion(128'heeac72d31c0aa315b1cd98e3b4aefe27, {16'd54092, 16'd52987, 16'd17727, 16'd54647, 16'd29169, 16'd60200, 16'd29257, 16'd46426, 16'd4173, 16'd11234, 16'd7962, 16'd11948, 16'd23684, 16'd48097, 16'd15673, 16'd18405, 16'd33897, 16'd31846, 16'd40797, 16'd168, 16'd45502, 16'd62748, 16'd11765, 16'd38092, 16'd32027, 16'd31092});
	test_expansion(128'ha136b3fdf3d0956b3cb4ac356bfaeffc, {16'd46211, 16'd23989, 16'd56932, 16'd17034, 16'd1318, 16'd1403, 16'd59781, 16'd46439, 16'd5230, 16'd12963, 16'd9813, 16'd51446, 16'd17088, 16'd16007, 16'd61024, 16'd4172, 16'd11994, 16'd20299, 16'd37390, 16'd9377, 16'd40842, 16'd9668, 16'd15114, 16'd27630, 16'd36289, 16'd12537});
	test_expansion(128'he28bd90e543e2e4c0efd1903ba9d6fd8, {16'd20879, 16'd35981, 16'd52228, 16'd25577, 16'd51563, 16'd8811, 16'd17141, 16'd33718, 16'd10335, 16'd7166, 16'd13671, 16'd53843, 16'd22454, 16'd48631, 16'd22597, 16'd34560, 16'd19183, 16'd17876, 16'd11872, 16'd34978, 16'd63941, 16'd42847, 16'd3862, 16'd40737, 16'd57093, 16'd51810});
	test_expansion(128'h9bd9b1239c5fecd33fee494eb544e575, {16'd25399, 16'd17632, 16'd59902, 16'd12886, 16'd4660, 16'd2180, 16'd61878, 16'd50222, 16'd46113, 16'd28950, 16'd35421, 16'd57620, 16'd33590, 16'd15327, 16'd65487, 16'd39985, 16'd57872, 16'd55654, 16'd43133, 16'd23610, 16'd23933, 16'd61272, 16'd45909, 16'd33953, 16'd17293, 16'd60116});
	test_expansion(128'hecc2452eeb681a59b02a1d93aee699e1, {16'd58182, 16'd64920, 16'd34650, 16'd15570, 16'd32797, 16'd53308, 16'd42813, 16'd51249, 16'd32000, 16'd30755, 16'd63933, 16'd12177, 16'd53791, 16'd53589, 16'd53454, 16'd32856, 16'd13653, 16'd39609, 16'd63859, 16'd12365, 16'd32524, 16'd43942, 16'd62029, 16'd5171, 16'd3391, 16'd17234});
	test_expansion(128'hf21b733fd0132f776fb0460598e5fcdd, {16'd48401, 16'd12884, 16'd51414, 16'd17644, 16'd9247, 16'd49925, 16'd59871, 16'd64599, 16'd2676, 16'd51591, 16'd57881, 16'd46398, 16'd43151, 16'd14577, 16'd30567, 16'd61069, 16'd16455, 16'd57711, 16'd45519, 16'd46164, 16'd18781, 16'd41701, 16'd44142, 16'd41487, 16'd34288, 16'd55464});
	test_expansion(128'h339e88c7e7253e53fafb74a4ec654571, {16'd26531, 16'd15809, 16'd39729, 16'd3506, 16'd58727, 16'd14740, 16'd38851, 16'd59793, 16'd28578, 16'd8141, 16'd46797, 16'd24194, 16'd40540, 16'd24474, 16'd57634, 16'd50218, 16'd6705, 16'd29714, 16'd47991, 16'd64534, 16'd20454, 16'd53332, 16'd57805, 16'd10346, 16'd59555, 16'd58435});
	test_expansion(128'h93944d0a8c2f0f5511bd6dc54068bb31, {16'd51963, 16'd3481, 16'd4171, 16'd31433, 16'd42065, 16'd50674, 16'd49173, 16'd7240, 16'd56718, 16'd38268, 16'd63620, 16'd28682, 16'd58094, 16'd7219, 16'd62493, 16'd41750, 16'd43256, 16'd27825, 16'd21195, 16'd23773, 16'd59772, 16'd39341, 16'd12598, 16'd4070, 16'd25042, 16'd1955});
	test_expansion(128'h317d049d577908a81202a29113ec4d04, {16'd58393, 16'd34046, 16'd230, 16'd21754, 16'd36691, 16'd64193, 16'd22428, 16'd47628, 16'd50441, 16'd63126, 16'd54969, 16'd3469, 16'd24051, 16'd63557, 16'd58428, 16'd33387, 16'd46262, 16'd45028, 16'd7940, 16'd26709, 16'd1736, 16'd52393, 16'd35590, 16'd20877, 16'd47372, 16'd23004});
	test_expansion(128'h935564ec09d11df4680ffaefe23af537, {16'd45257, 16'd16971, 16'd38979, 16'd40261, 16'd14928, 16'd24873, 16'd28792, 16'd49246, 16'd53595, 16'd42871, 16'd44759, 16'd31078, 16'd12636, 16'd11051, 16'd60022, 16'd24119, 16'd58048, 16'd29747, 16'd25520, 16'd31204, 16'd2762, 16'd52606, 16'd4585, 16'd45036, 16'd45869, 16'd61601});
	test_expansion(128'h9ae562b241516aa8785564b6fa6d2137, {16'd59093, 16'd44243, 16'd12163, 16'd40478, 16'd58142, 16'd53226, 16'd2999, 16'd39254, 16'd23980, 16'd28960, 16'd40054, 16'd18193, 16'd17952, 16'd62150, 16'd43654, 16'd24212, 16'd17053, 16'd42846, 16'd37818, 16'd63482, 16'd23623, 16'd26063, 16'd44185, 16'd44007, 16'd364, 16'd9385});
	test_expansion(128'h5a3ac109a2720f4be011e2a8271e09a1, {16'd37981, 16'd2055, 16'd60205, 16'd10214, 16'd7349, 16'd931, 16'd52362, 16'd51562, 16'd35718, 16'd11831, 16'd45801, 16'd15952, 16'd56997, 16'd34746, 16'd27923, 16'd53487, 16'd41799, 16'd40256, 16'd2183, 16'd36674, 16'd2300, 16'd63581, 16'd6236, 16'd7849, 16'd13649, 16'd61650});
	test_expansion(128'h7d0b2b165f7639375307850fa719d31e, {16'd19254, 16'd49632, 16'd31076, 16'd63907, 16'd9490, 16'd44251, 16'd54031, 16'd27748, 16'd23219, 16'd11266, 16'd21180, 16'd61120, 16'd15987, 16'd3517, 16'd11851, 16'd18840, 16'd65288, 16'd58441, 16'd23877, 16'd10323, 16'd41932, 16'd40155, 16'd41154, 16'd3130, 16'd36485, 16'd59357});
	test_expansion(128'hc4fddb278390d2f0ba93273a100cede2, {16'd23651, 16'd44412, 16'd44933, 16'd33328, 16'd37078, 16'd23406, 16'd33122, 16'd18066, 16'd20995, 16'd58745, 16'd8329, 16'd25192, 16'd51278, 16'd57297, 16'd39906, 16'd18559, 16'd38476, 16'd5599, 16'd1405, 16'd62004, 16'd49973, 16'd13222, 16'd33875, 16'd16016, 16'd41694, 16'd18452});
	test_expansion(128'h0a6a946e3122df7c978f97f1562979d2, {16'd16040, 16'd26901, 16'd53145, 16'd52484, 16'd63984, 16'd12396, 16'd51855, 16'd56758, 16'd13295, 16'd8895, 16'd13483, 16'd12109, 16'd964, 16'd48172, 16'd9134, 16'd50980, 16'd14479, 16'd48016, 16'd40381, 16'd34067, 16'd46857, 16'd10697, 16'd27798, 16'd14534, 16'd19177, 16'd40612});
	test_expansion(128'ha412e5943f2fcd18a5163dbb68e7acfd, {16'd3222, 16'd64498, 16'd46099, 16'd62003, 16'd10169, 16'd46779, 16'd44105, 16'd1691, 16'd62004, 16'd62806, 16'd33709, 16'd41117, 16'd8544, 16'd8026, 16'd44475, 16'd28638, 16'd12906, 16'd13796, 16'd33068, 16'd13072, 16'd27229, 16'd64523, 16'd7682, 16'd49287, 16'd24343, 16'd19626});
	test_expansion(128'h7a93fdbd7de32f692f28a25fa67e2848, {16'd21025, 16'd31510, 16'd9267, 16'd38261, 16'd54965, 16'd31187, 16'd8280, 16'd8508, 16'd5632, 16'd38517, 16'd15727, 16'd4093, 16'd28372, 16'd21134, 16'd56293, 16'd52691, 16'd33861, 16'd11147, 16'd43886, 16'd36821, 16'd259, 16'd55729, 16'd32316, 16'd31498, 16'd7933, 16'd55148});
	test_expansion(128'hc7a52e8aa6bd57f11a4a4ed970a09dbe, {16'd60303, 16'd3157, 16'd53338, 16'd33177, 16'd54389, 16'd52604, 16'd41196, 16'd36984, 16'd2708, 16'd16123, 16'd36857, 16'd28905, 16'd54952, 16'd43838, 16'd13968, 16'd58618, 16'd11325, 16'd58131, 16'd26957, 16'd39110, 16'd37226, 16'd16314, 16'd6435, 16'd64330, 16'd26774, 16'd8158});
	test_expansion(128'h945ff6bd465574e08d45b5fff3df3631, {16'd5138, 16'd36862, 16'd56296, 16'd13682, 16'd50460, 16'd11669, 16'd49165, 16'd8037, 16'd12986, 16'd10542, 16'd18342, 16'd28059, 16'd40230, 16'd52634, 16'd14144, 16'd44550, 16'd11947, 16'd48035, 16'd21601, 16'd30617, 16'd27526, 16'd9006, 16'd33182, 16'd41217, 16'd17800, 16'd25806});
	test_expansion(128'hd5d8e168f156de29c49303e18dbbb60b, {16'd49467, 16'd19216, 16'd50201, 16'd23190, 16'd13045, 16'd39921, 16'd23298, 16'd15926, 16'd41336, 16'd50968, 16'd26567, 16'd29554, 16'd8910, 16'd22139, 16'd53701, 16'd14068, 16'd65362, 16'd60754, 16'd23961, 16'd22008, 16'd47409, 16'd28070, 16'd37142, 16'd47748, 16'd36091, 16'd48515});
	test_expansion(128'hbbb21b8b2cd1ec0feaafdf2a3e76fa6d, {16'd11311, 16'd54262, 16'd11060, 16'd40986, 16'd58487, 16'd54161, 16'd34552, 16'd35390, 16'd18353, 16'd13908, 16'd1246, 16'd13249, 16'd59641, 16'd12534, 16'd13975, 16'd63670, 16'd48757, 16'd18133, 16'd35105, 16'd61647, 16'd4603, 16'd16667, 16'd8319, 16'd11022, 16'd57082, 16'd25941});
	test_expansion(128'hc09082084347405a32126288bc472bea, {16'd49404, 16'd55337, 16'd38926, 16'd964, 16'd44532, 16'd36969, 16'd25692, 16'd2368, 16'd18381, 16'd43488, 16'd38855, 16'd19428, 16'd4163, 16'd18993, 16'd53494, 16'd60510, 16'd21565, 16'd52507, 16'd3215, 16'd49137, 16'd64859, 16'd51111, 16'd16249, 16'd37437, 16'd13167, 16'd19834});
	test_expansion(128'h61ee32a9417d66e3bd2dfcf0fad2770c, {16'd57202, 16'd42104, 16'd41899, 16'd64032, 16'd11785, 16'd16476, 16'd34878, 16'd37772, 16'd1467, 16'd10882, 16'd63546, 16'd2998, 16'd22734, 16'd46879, 16'd49155, 16'd64571, 16'd17907, 16'd50767, 16'd37488, 16'd4198, 16'd64529, 16'd52047, 16'd60941, 16'd27114, 16'd24663, 16'd53509});
	test_expansion(128'h06c1a9c82fdb092828729b2de5c8ada1, {16'd22047, 16'd57426, 16'd23848, 16'd43092, 16'd62044, 16'd54220, 16'd47879, 16'd60008, 16'd20098, 16'd324, 16'd26352, 16'd55388, 16'd35039, 16'd64928, 16'd29253, 16'd34876, 16'd33235, 16'd15482, 16'd43351, 16'd32120, 16'd14600, 16'd32890, 16'd51128, 16'd50741, 16'd39971, 16'd9661});
	test_expansion(128'h40e9bb22d5d2acf7021be0f9ed81ec80, {16'd62623, 16'd9668, 16'd21584, 16'd18928, 16'd15537, 16'd4959, 16'd10910, 16'd59734, 16'd34163, 16'd53047, 16'd14828, 16'd31015, 16'd21830, 16'd41704, 16'd16474, 16'd62563, 16'd16585, 16'd47794, 16'd12492, 16'd40186, 16'd9544, 16'd3914, 16'd56776, 16'd28327, 16'd30032, 16'd63989});
	test_expansion(128'h7d0ca42bb53234b22edbc9283e9212f6, {16'd20703, 16'd55824, 16'd1715, 16'd61132, 16'd13088, 16'd51076, 16'd59125, 16'd59313, 16'd8189, 16'd8660, 16'd49312, 16'd27237, 16'd5832, 16'd51652, 16'd12060, 16'd61789, 16'd43806, 16'd38475, 16'd31821, 16'd11174, 16'd38215, 16'd31534, 16'd50653, 16'd26495, 16'd62393, 16'd18776});
	test_expansion(128'h5565ceb273e57b01069efa0a6916b8bf, {16'd4019, 16'd10131, 16'd50002, 16'd328, 16'd13889, 16'd50368, 16'd20476, 16'd42991, 16'd63636, 16'd24723, 16'd59767, 16'd58612, 16'd37167, 16'd38653, 16'd49958, 16'd26830, 16'd9962, 16'd31979, 16'd2298, 16'd25018, 16'd19914, 16'd36653, 16'd31289, 16'd37294, 16'd39841, 16'd34232});
	test_expansion(128'h3434959036f20fbc9e6629a6b2eee662, {16'd62642, 16'd11951, 16'd57910, 16'd40386, 16'd55002, 16'd45318, 16'd57228, 16'd48559, 16'd27076, 16'd51641, 16'd51955, 16'd37991, 16'd13888, 16'd4731, 16'd39390, 16'd2760, 16'd37127, 16'd58292, 16'd58563, 16'd48636, 16'd24713, 16'd29319, 16'd14378, 16'd30001, 16'd35622, 16'd57774});
	test_expansion(128'h90adb9956ac08aad3e23574440de1549, {16'd38908, 16'd59201, 16'd55308, 16'd64399, 16'd60156, 16'd9749, 16'd38419, 16'd4280, 16'd626, 16'd29334, 16'd21816, 16'd50862, 16'd33413, 16'd2945, 16'd16395, 16'd54362, 16'd7377, 16'd391, 16'd62682, 16'd40134, 16'd2278, 16'd22341, 16'd49338, 16'd43274, 16'd41291, 16'd8975});
	test_expansion(128'h0895f0f7d4bee8b9faf19917f4f6e808, {16'd38807, 16'd31241, 16'd51426, 16'd58784, 16'd24273, 16'd49576, 16'd31917, 16'd11266, 16'd24881, 16'd3813, 16'd50803, 16'd49495, 16'd63790, 16'd51349, 16'd41990, 16'd14506, 16'd55114, 16'd38845, 16'd19468, 16'd56183, 16'd45752, 16'd25419, 16'd63311, 16'd19566, 16'd57291, 16'd38335});
	test_expansion(128'h46481f8988f9f5e705f92ee30a8ce2a3, {16'd13644, 16'd8838, 16'd56613, 16'd56547, 16'd6713, 16'd31709, 16'd46936, 16'd56194, 16'd47950, 16'd12406, 16'd43230, 16'd48206, 16'd51115, 16'd21110, 16'd9449, 16'd10752, 16'd54814, 16'd17393, 16'd31283, 16'd24738, 16'd1244, 16'd43633, 16'd60840, 16'd58030, 16'd7076, 16'd16272});
	test_expansion(128'h76bca071fd3cfabd851be8eaac0975b3, {16'd34626, 16'd15493, 16'd16006, 16'd51295, 16'd41038, 16'd58047, 16'd12705, 16'd24327, 16'd57516, 16'd10092, 16'd20861, 16'd25544, 16'd37737, 16'd33238, 16'd9275, 16'd8699, 16'd20375, 16'd32715, 16'd22591, 16'd39008, 16'd50305, 16'd39968, 16'd54440, 16'd29392, 16'd64441, 16'd48253});
	test_expansion(128'h1df0666cfe845e2cd95a736acc0d6a89, {16'd44339, 16'd21726, 16'd46158, 16'd51256, 16'd42561, 16'd2286, 16'd2514, 16'd9526, 16'd33027, 16'd54010, 16'd10803, 16'd16821, 16'd38985, 16'd13426, 16'd44004, 16'd16047, 16'd41224, 16'd17798, 16'd57479, 16'd4996, 16'd64712, 16'd33295, 16'd54181, 16'd55462, 16'd46821, 16'd46052});
	test_expansion(128'h1172c779c8bb16778e23e760835380b0, {16'd31009, 16'd42882, 16'd46498, 16'd16105, 16'd27135, 16'd2954, 16'd55177, 16'd48813, 16'd56190, 16'd23428, 16'd28688, 16'd7613, 16'd52868, 16'd26960, 16'd38813, 16'd33073, 16'd43163, 16'd1663, 16'd28075, 16'd12839, 16'd50502, 16'd51066, 16'd8417, 16'd33000, 16'd1932, 16'd28479});
	test_expansion(128'h278cc8d143fbcf0bceeb3a34777c5a6b, {16'd64753, 16'd18530, 16'd35749, 16'd34717, 16'd11465, 16'd28387, 16'd11792, 16'd36548, 16'd2574, 16'd62012, 16'd31997, 16'd22115, 16'd33868, 16'd57125, 16'd58875, 16'd7886, 16'd56439, 16'd51878, 16'd41404, 16'd3571, 16'd62941, 16'd3874, 16'd50777, 16'd31942, 16'd43442, 16'd17346});
	test_expansion(128'h50788ccb0431c1bbfa34c013d1a9b438, {16'd39402, 16'd28006, 16'd41765, 16'd26660, 16'd1432, 16'd52229, 16'd27533, 16'd31169, 16'd39900, 16'd48776, 16'd87, 16'd22225, 16'd36653, 16'd55525, 16'd65143, 16'd32962, 16'd46845, 16'd35797, 16'd3224, 16'd64716, 16'd28706, 16'd56077, 16'd58343, 16'd23440, 16'd39771, 16'd36476});
	test_expansion(128'ha3b42e183030b4aefc71462adc02408d, {16'd53386, 16'd24480, 16'd53143, 16'd62833, 16'd6746, 16'd25574, 16'd57046, 16'd27979, 16'd12339, 16'd10640, 16'd42054, 16'd22219, 16'd5537, 16'd24618, 16'd5865, 16'd19203, 16'd333, 16'd64795, 16'd45409, 16'd37719, 16'd29677, 16'd39307, 16'd17665, 16'd53109, 16'd15116, 16'd3258});
	test_expansion(128'hba667b0eea91f83e070c87c56c182c7f, {16'd203, 16'd41229, 16'd41205, 16'd42682, 16'd25131, 16'd8513, 16'd56184, 16'd238, 16'd46659, 16'd502, 16'd47249, 16'd35651, 16'd6534, 16'd4573, 16'd283, 16'd44353, 16'd50049, 16'd55020, 16'd19738, 16'd58904, 16'd38211, 16'd40437, 16'd5442, 16'd55207, 16'd30437, 16'd15404});
	test_expansion(128'h191b48e6d6098444c1a87b623a698813, {16'd30236, 16'd2828, 16'd19031, 16'd51993, 16'd58998, 16'd15820, 16'd37288, 16'd58715, 16'd52598, 16'd37601, 16'd12348, 16'd48945, 16'd46547, 16'd24408, 16'd35358, 16'd23248, 16'd32842, 16'd13450, 16'd50875, 16'd20924, 16'd61225, 16'd64275, 16'd46593, 16'd26523, 16'd18432, 16'd53277});
	test_expansion(128'h62e9433cdee53df041a847f484e2e34f, {16'd36265, 16'd20431, 16'd60737, 16'd18319, 16'd45655, 16'd13718, 16'd32776, 16'd39053, 16'd34133, 16'd46108, 16'd56527, 16'd33249, 16'd4295, 16'd43271, 16'd51492, 16'd54845, 16'd57278, 16'd42745, 16'd32399, 16'd60776, 16'd19597, 16'd48550, 16'd12252, 16'd34710, 16'd16775, 16'd54967});
	test_expansion(128'h2c95a435dec4e9dbe68b9990abe2829a, {16'd38451, 16'd2277, 16'd11414, 16'd6363, 16'd11519, 16'd2642, 16'd17786, 16'd45897, 16'd45086, 16'd62580, 16'd29419, 16'd41392, 16'd24358, 16'd1311, 16'd49332, 16'd37444, 16'd17903, 16'd29287, 16'd55807, 16'd50541, 16'd24446, 16'd55105, 16'd29423, 16'd21922, 16'd23809, 16'd29127});
	test_expansion(128'h9d31da58157e4576e962a65edeba44ab, {16'd22615, 16'd50672, 16'd9946, 16'd59887, 16'd43929, 16'd44615, 16'd54304, 16'd43568, 16'd10841, 16'd49397, 16'd61703, 16'd521, 16'd24941, 16'd38243, 16'd38715, 16'd65317, 16'd10068, 16'd37820, 16'd43794, 16'd56146, 16'd454, 16'd6842, 16'd29739, 16'd6397, 16'd42811, 16'd2592});
	test_expansion(128'hd80f017251159b5c7b4bdb971e9a9f61, {16'd31298, 16'd6245, 16'd33954, 16'd32615, 16'd28752, 16'd29224, 16'd45646, 16'd35960, 16'd2996, 16'd35347, 16'd53666, 16'd8790, 16'd38895, 16'd1744, 16'd43741, 16'd32101, 16'd13697, 16'd22442, 16'd20803, 16'd48719, 16'd14992, 16'd23153, 16'd7561, 16'd31233, 16'd40134, 16'd43534});
	test_expansion(128'h4eb91cf99a9aa738a41277c4ef55729b, {16'd50965, 16'd24722, 16'd36169, 16'd19688, 16'd22614, 16'd50790, 16'd59723, 16'd64588, 16'd9908, 16'd51327, 16'd54006, 16'd20661, 16'd19822, 16'd41247, 16'd11632, 16'd24849, 16'd34963, 16'd43960, 16'd57330, 16'd33002, 16'd63758, 16'd17674, 16'd40817, 16'd52717, 16'd61771, 16'd48310});
	test_expansion(128'hef54cff3e9f8b41a77d1b72a2e5d2ee6, {16'd23781, 16'd9574, 16'd17056, 16'd60910, 16'd25109, 16'd10125, 16'd43689, 16'd5967, 16'd58338, 16'd22112, 16'd21663, 16'd41390, 16'd48025, 16'd57603, 16'd42483, 16'd41605, 16'd6379, 16'd37924, 16'd33346, 16'd53975, 16'd47119, 16'd46444, 16'd34589, 16'd27066, 16'd18807, 16'd38739});
	test_expansion(128'h89043228d301da0b91bcfac4ecd919ad, {16'd18441, 16'd44189, 16'd46249, 16'd928, 16'd48201, 16'd35301, 16'd31808, 16'd44575, 16'd20575, 16'd15164, 16'd4623, 16'd60534, 16'd58151, 16'd42166, 16'd58676, 16'd3916, 16'd37773, 16'd2599, 16'd15269, 16'd54556, 16'd61963, 16'd344, 16'd55315, 16'd23963, 16'd22610, 16'd1057});
	test_expansion(128'hf7fa3a584741d2d9d19c0b36259918ff, {16'd38638, 16'd27784, 16'd31974, 16'd46251, 16'd64678, 16'd18497, 16'd14703, 16'd64544, 16'd60356, 16'd16526, 16'd63745, 16'd22661, 16'd34679, 16'd58325, 16'd29910, 16'd47210, 16'd62175, 16'd23240, 16'd56846, 16'd52568, 16'd56517, 16'd7309, 16'd22846, 16'd39592, 16'd16386, 16'd58545});
	test_expansion(128'hadd668d7cfa0fe6016fbdc25acee2486, {16'd56608, 16'd41297, 16'd25181, 16'd27181, 16'd30018, 16'd18555, 16'd43610, 16'd54538, 16'd63790, 16'd15863, 16'd20049, 16'd4472, 16'd52956, 16'd23508, 16'd6328, 16'd6306, 16'd56894, 16'd41508, 16'd14139, 16'd21680, 16'd1342, 16'd22852, 16'd24223, 16'd5108, 16'd33073, 16'd7849});
	test_expansion(128'h850d075c576e28f8e497aba7359896b6, {16'd30110, 16'd9112, 16'd46113, 16'd20402, 16'd18573, 16'd6026, 16'd44132, 16'd20972, 16'd28326, 16'd57507, 16'd50673, 16'd32669, 16'd22943, 16'd31256, 16'd65449, 16'd2572, 16'd44413, 16'd17690, 16'd4298, 16'd24092, 16'd1814, 16'd64507, 16'd21063, 16'd38211, 16'd15564, 16'd16766});
	test_expansion(128'hd7e066a365be500dcc9c161134f76e20, {16'd20145, 16'd59457, 16'd19454, 16'd7208, 16'd9160, 16'd64965, 16'd49641, 16'd51668, 16'd25647, 16'd2442, 16'd40001, 16'd61293, 16'd8688, 16'd50577, 16'd29611, 16'd3890, 16'd6901, 16'd37044, 16'd36894, 16'd20452, 16'd56988, 16'd30369, 16'd64019, 16'd6857, 16'd44610, 16'd53029});
	test_expansion(128'h1234a7ffbe0b6ff87ab840569b2a30e3, {16'd9842, 16'd43979, 16'd52106, 16'd6299, 16'd19266, 16'd61241, 16'd40336, 16'd19581, 16'd18913, 16'd54278, 16'd54869, 16'd47416, 16'd56451, 16'd4007, 16'd42582, 16'd34828, 16'd25474, 16'd16402, 16'd21142, 16'd47509, 16'd9015, 16'd7785, 16'd17061, 16'd60368, 16'd16651, 16'd44993});
	test_expansion(128'h28e8c1fabd69d0dbfe5514a0dfe921c5, {16'd49361, 16'd36850, 16'd45878, 16'd20910, 16'd16014, 16'd8140, 16'd12400, 16'd62668, 16'd15291, 16'd1667, 16'd56595, 16'd5443, 16'd6904, 16'd33019, 16'd54586, 16'd24334, 16'd53493, 16'd19435, 16'd45412, 16'd60701, 16'd53990, 16'd36906, 16'd40051, 16'd6753, 16'd62829, 16'd53924});
	test_expansion(128'h591c06f98caf269fb650f38b94a5a717, {16'd19352, 16'd42997, 16'd20831, 16'd31254, 16'd2357, 16'd35998, 16'd19160, 16'd48593, 16'd35774, 16'd60506, 16'd30143, 16'd18669, 16'd19125, 16'd17267, 16'd27124, 16'd64374, 16'd25871, 16'd49075, 16'd22924, 16'd26063, 16'd28998, 16'd35943, 16'd26395, 16'd61656, 16'd48033, 16'd952});
	test_expansion(128'h64a7771c37618216bd07836bb10392e7, {16'd33002, 16'd44984, 16'd35070, 16'd61117, 16'd15995, 16'd55584, 16'd25220, 16'd37574, 16'd57138, 16'd12047, 16'd3564, 16'd16680, 16'd8274, 16'd4611, 16'd48735, 16'd7515, 16'd28309, 16'd41174, 16'd1769, 16'd38581, 16'd7632, 16'd3604, 16'd37654, 16'd12810, 16'd16976, 16'd61863});
	test_expansion(128'h401ba8c49cdb84b8d4a41eb37129feb9, {16'd37598, 16'd35288, 16'd5325, 16'd28043, 16'd60425, 16'd42469, 16'd42840, 16'd48741, 16'd54476, 16'd19481, 16'd64184, 16'd48341, 16'd53357, 16'd61234, 16'd6425, 16'd45537, 16'd36408, 16'd9239, 16'd14052, 16'd51338, 16'd9198, 16'd37793, 16'd44326, 16'd34674, 16'd48514, 16'd36706});
	test_expansion(128'h547f6af7fa7d39d2437542732cab4b6d, {16'd1074, 16'd51429, 16'd3474, 16'd9450, 16'd59681, 16'd54947, 16'd33981, 16'd45510, 16'd61152, 16'd55940, 16'd56367, 16'd9371, 16'd11736, 16'd30358, 16'd773, 16'd31849, 16'd40665, 16'd29369, 16'd65006, 16'd53138, 16'd56365, 16'd30291, 16'd9243, 16'd20468, 16'd4342, 16'd40320});
	test_expansion(128'hc9f0b6654fee09981ac59057ab817e01, {16'd22287, 16'd41610, 16'd56028, 16'd14745, 16'd5838, 16'd45245, 16'd7433, 16'd21515, 16'd16539, 16'd47291, 16'd10259, 16'd63952, 16'd52236, 16'd53316, 16'd751, 16'd20753, 16'd11862, 16'd2378, 16'd46545, 16'd28899, 16'd17457, 16'd34947, 16'd3452, 16'd54462, 16'd16738, 16'd41873});
	test_expansion(128'h68f7f2418eb3eacdbb6b3dca18b82a7e, {16'd36981, 16'd62078, 16'd36892, 16'd10304, 16'd21077, 16'd22358, 16'd29818, 16'd41595, 16'd37499, 16'd32545, 16'd44364, 16'd1100, 16'd9611, 16'd38505, 16'd11283, 16'd61411, 16'd58946, 16'd64835, 16'd16441, 16'd30904, 16'd56415, 16'd28247, 16'd44140, 16'd18563, 16'd3727, 16'd4871});
	test_expansion(128'h94a86d7e1d29d0a7ecbab31c454fb306, {16'd47849, 16'd29969, 16'd34047, 16'd45073, 16'd37651, 16'd6261, 16'd50504, 16'd8776, 16'd45307, 16'd23364, 16'd39710, 16'd61822, 16'd28016, 16'd14743, 16'd52515, 16'd9045, 16'd38034, 16'd5431, 16'd34034, 16'd53220, 16'd34100, 16'd48781, 16'd39165, 16'd14899, 16'd33416, 16'd44896});
	test_expansion(128'hd46a37a6e9be83594a4784b39eb9fbe5, {16'd27768, 16'd51900, 16'd9622, 16'd17225, 16'd47218, 16'd36911, 16'd64359, 16'd20640, 16'd5042, 16'd29932, 16'd46353, 16'd2415, 16'd61078, 16'd49850, 16'd1848, 16'd18274, 16'd9633, 16'd17625, 16'd46933, 16'd39785, 16'd5666, 16'd56506, 16'd27253, 16'd63787, 16'd34406, 16'd18540});
	test_expansion(128'h9a15895c8a13784ca0767fd925a64b14, {16'd52756, 16'd56031, 16'd29187, 16'd54989, 16'd4740, 16'd17683, 16'd43599, 16'd6691, 16'd54505, 16'd13747, 16'd19636, 16'd21669, 16'd33439, 16'd56164, 16'd10862, 16'd40270, 16'd34762, 16'd20775, 16'd18336, 16'd13963, 16'd22414, 16'd14340, 16'd65187, 16'd36623, 16'd18099, 16'd60429});
	test_expansion(128'h0dbb8c0e45d2f7b4fbbc7e8851688472, {16'd5863, 16'd27246, 16'd61171, 16'd57583, 16'd19599, 16'd58454, 16'd28356, 16'd42997, 16'd52241, 16'd18991, 16'd42878, 16'd28220, 16'd52977, 16'd44879, 16'd27835, 16'd40858, 16'd62051, 16'd43114, 16'd58416, 16'd33612, 16'd28957, 16'd57250, 16'd21056, 16'd56393, 16'd56168, 16'd19932});
	test_expansion(128'hdd1fc7b52e58b64685a2bfed7e7e02b1, {16'd51635, 16'd38921, 16'd2302, 16'd45570, 16'd1030, 16'd52735, 16'd7921, 16'd35055, 16'd24303, 16'd47768, 16'd42441, 16'd6280, 16'd54026, 16'd52515, 16'd2872, 16'd51760, 16'd64539, 16'd48887, 16'd25456, 16'd32724, 16'd9209, 16'd48565, 16'd14230, 16'd1557, 16'd6611, 16'd30485});
	test_expansion(128'h13e62066f41b0fe3c18eba32a6196630, {16'd19783, 16'd28612, 16'd19054, 16'd50338, 16'd53722, 16'd54544, 16'd5204, 16'd51564, 16'd61771, 16'd41553, 16'd48326, 16'd58263, 16'd59124, 16'd11274, 16'd26523, 16'd28644, 16'd8935, 16'd64578, 16'd46252, 16'd27329, 16'd45584, 16'd4648, 16'd9417, 16'd3588, 16'd22636, 16'd56749});
	test_expansion(128'h90a334c31acae100d5dea958571d21e2, {16'd20561, 16'd34513, 16'd5193, 16'd16062, 16'd5148, 16'd47508, 16'd14259, 16'd39767, 16'd59563, 16'd54654, 16'd10696, 16'd39689, 16'd35155, 16'd58680, 16'd39559, 16'd12293, 16'd14270, 16'd904, 16'd4907, 16'd43551, 16'd408, 16'd5886, 16'd18464, 16'd20654, 16'd26396, 16'd29876});
	test_expansion(128'h8a8ede420e3ddeda57ad08bb87de5f0f, {16'd31627, 16'd17304, 16'd28031, 16'd62731, 16'd14195, 16'd16593, 16'd51239, 16'd31488, 16'd7359, 16'd21724, 16'd24763, 16'd1731, 16'd24833, 16'd41301, 16'd21038, 16'd52862, 16'd31046, 16'd44647, 16'd46704, 16'd60597, 16'd12486, 16'd47801, 16'd25787, 16'd24235, 16'd10733, 16'd15378});
	test_expansion(128'h604f25596ac067d7b5e09dd71f9bf3a8, {16'd41939, 16'd49798, 16'd58439, 16'd54157, 16'd65195, 16'd10463, 16'd62605, 16'd10684, 16'd3398, 16'd11241, 16'd6464, 16'd16441, 16'd46086, 16'd44677, 16'd3468, 16'd27657, 16'd49811, 16'd24194, 16'd41437, 16'd15838, 16'd54758, 16'd15380, 16'd20939, 16'd63083, 16'd10484, 16'd40789});
	test_expansion(128'h1da8964f7e5183958906e0390db608cc, {16'd60760, 16'd59566, 16'd14805, 16'd23058, 16'd37565, 16'd19738, 16'd25141, 16'd16303, 16'd28640, 16'd47169, 16'd9698, 16'd58937, 16'd55875, 16'd21896, 16'd42972, 16'd21443, 16'd24122, 16'd5800, 16'd60552, 16'd48201, 16'd7923, 16'd59662, 16'd60961, 16'd18876, 16'd2636, 16'd23737});
	test_expansion(128'h7f6339a37d5a3b703720b0d2febec38d, {16'd41011, 16'd28313, 16'd15209, 16'd27465, 16'd59878, 16'd41822, 16'd49800, 16'd32264, 16'd60649, 16'd55965, 16'd3009, 16'd35387, 16'd12824, 16'd43608, 16'd40186, 16'd5134, 16'd45221, 16'd5364, 16'd47531, 16'd12850, 16'd20272, 16'd13554, 16'd19928, 16'd32150, 16'd5845, 16'd6341});
	test_expansion(128'hd26c0dc8dcbb4f05d4476432fc05d720, {16'd45478, 16'd60813, 16'd8969, 16'd14409, 16'd50444, 16'd20074, 16'd27112, 16'd49653, 16'd28977, 16'd48315, 16'd48924, 16'd51870, 16'd49974, 16'd30722, 16'd53178, 16'd60286, 16'd27078, 16'd26175, 16'd28720, 16'd58603, 16'd15846, 16'd56090, 16'd35003, 16'd20064, 16'd31397, 16'd10816});
	test_expansion(128'hf53bd577b3ce297e0c5b900908cfb822, {16'd49619, 16'd43426, 16'd33364, 16'd19311, 16'd51657, 16'd41246, 16'd52336, 16'd58557, 16'd22716, 16'd210, 16'd28166, 16'd62989, 16'd57072, 16'd35645, 16'd12604, 16'd7737, 16'd22663, 16'd27870, 16'd53374, 16'd24594, 16'd50653, 16'd46822, 16'd24678, 16'd34515, 16'd63617, 16'd35715});
	test_expansion(128'h4198dea4996bb813867ddd72b3ab54b2, {16'd44722, 16'd65470, 16'd51584, 16'd51638, 16'd29112, 16'd36340, 16'd42361, 16'd61982, 16'd16581, 16'd1434, 16'd23271, 16'd32455, 16'd8205, 16'd32555, 16'd6822, 16'd22466, 16'd35945, 16'd65207, 16'd43477, 16'd58594, 16'd50544, 16'd65175, 16'd21636, 16'd31870, 16'd26790, 16'd64293});
	test_expansion(128'hf4fdb38a8aa26bab3fdbdb3cacab0d53, {16'd43010, 16'd65224, 16'd29739, 16'd38319, 16'd43438, 16'd36795, 16'd43366, 16'd55635, 16'd9448, 16'd2515, 16'd44878, 16'd5971, 16'd27604, 16'd44351, 16'd32401, 16'd20187, 16'd49424, 16'd30533, 16'd50713, 16'd46663, 16'd46003, 16'd23960, 16'd48377, 16'd26276, 16'd61907, 16'd36333});
	test_expansion(128'h8c775a3ceddcc04aca413e5c13df6f9c, {16'd23234, 16'd37793, 16'd14282, 16'd21346, 16'd1816, 16'd28927, 16'd64359, 16'd434, 16'd57244, 16'd55954, 16'd41848, 16'd45972, 16'd37337, 16'd53636, 16'd16634, 16'd63071, 16'd25906, 16'd44276, 16'd32272, 16'd16689, 16'd30391, 16'd20886, 16'd18861, 16'd546, 16'd52730, 16'd35837});
	test_expansion(128'hc71aa9811380393cc264575053deacc7, {16'd29463, 16'd34260, 16'd56716, 16'd10151, 16'd25926, 16'd60057, 16'd64818, 16'd38409, 16'd58642, 16'd35546, 16'd7948, 16'd27442, 16'd29228, 16'd17961, 16'd18016, 16'd53749, 16'd37802, 16'd5949, 16'd5545, 16'd20846, 16'd2523, 16'd3589, 16'd16488, 16'd7773, 16'd17822, 16'd62683});
	test_expansion(128'h9038446ac130b3b07e4cb97bad8f9dff, {16'd6642, 16'd2478, 16'd27177, 16'd35428, 16'd14565, 16'd13606, 16'd28935, 16'd7765, 16'd44356, 16'd43622, 16'd4598, 16'd25623, 16'd36433, 16'd15439, 16'd26959, 16'd33324, 16'd55178, 16'd42345, 16'd24994, 16'd52444, 16'd38739, 16'd28635, 16'd39160, 16'd2183, 16'd23993, 16'd53223});
	test_expansion(128'hcfa29118835b8b5a4b5ffaa0952d929f, {16'd55291, 16'd52684, 16'd9622, 16'd55361, 16'd33414, 16'd3151, 16'd641, 16'd20797, 16'd33406, 16'd38821, 16'd11270, 16'd21959, 16'd49886, 16'd48302, 16'd29622, 16'd64187, 16'd19133, 16'd50883, 16'd51522, 16'd14382, 16'd42568, 16'd33291, 16'd23836, 16'd20650, 16'd34230, 16'd20309});
	test_expansion(128'hb9c9408339efcbb1194e6b7f46725eaa, {16'd35515, 16'd5004, 16'd38806, 16'd13798, 16'd193, 16'd62473, 16'd35892, 16'd50404, 16'd57653, 16'd22759, 16'd30660, 16'd17606, 16'd24578, 16'd35072, 16'd38983, 16'd1923, 16'd45503, 16'd50660, 16'd42877, 16'd25955, 16'd41517, 16'd11398, 16'd37124, 16'd38596, 16'd41101, 16'd43084});
	test_expansion(128'hb6f5de180893ff782d4af59b29c8907d, {16'd28585, 16'd29913, 16'd20945, 16'd54995, 16'd7969, 16'd52451, 16'd2985, 16'd39799, 16'd18333, 16'd47907, 16'd24066, 16'd63056, 16'd32398, 16'd7947, 16'd53275, 16'd51826, 16'd29825, 16'd59788, 16'd14110, 16'd1875, 16'd32500, 16'd12484, 16'd38770, 16'd42461, 16'd26659, 16'd6382});
	test_expansion(128'h13f81910ce1eae4ee6ac2266db08ff4c, {16'd52585, 16'd16841, 16'd46495, 16'd60586, 16'd6320, 16'd17044, 16'd44975, 16'd10379, 16'd11783, 16'd2655, 16'd25076, 16'd9110, 16'd13744, 16'd12758, 16'd9719, 16'd7679, 16'd59139, 16'd15235, 16'd28019, 16'd59115, 16'd3366, 16'd19495, 16'd44976, 16'd26369, 16'd44053, 16'd65064});
	test_expansion(128'h4a7faf6d50d078e1d2a73a025e2b2a18, {16'd23726, 16'd51071, 16'd41749, 16'd22011, 16'd52226, 16'd11523, 16'd31882, 16'd8545, 16'd29801, 16'd34714, 16'd52864, 16'd56703, 16'd65520, 16'd57088, 16'd25236, 16'd47742, 16'd9318, 16'd2172, 16'd40409, 16'd833, 16'd59201, 16'd42641, 16'd18506, 16'd65260, 16'd14807, 16'd37218});
	test_expansion(128'h0c0db62f9493ab2e9b1ebd821e0194c1, {16'd50094, 16'd22020, 16'd10990, 16'd26404, 16'd28918, 16'd18239, 16'd9774, 16'd10936, 16'd11247, 16'd13820, 16'd6215, 16'd16468, 16'd35174, 16'd9024, 16'd2262, 16'd30609, 16'd30631, 16'd59714, 16'd65109, 16'd35551, 16'd6385, 16'd56625, 16'd3631, 16'd47343, 16'd2287, 16'd8174});
	test_expansion(128'ha59bc98fb73b7866e024663326f133c6, {16'd16954, 16'd26627, 16'd11392, 16'd16631, 16'd46601, 16'd21019, 16'd38746, 16'd19486, 16'd48195, 16'd44735, 16'd32075, 16'd164, 16'd11714, 16'd20396, 16'd45616, 16'd17640, 16'd31163, 16'd46744, 16'd1762, 16'd55215, 16'd4219, 16'd41933, 16'd23342, 16'd3411, 16'd43630, 16'd9734});
	test_expansion(128'hfb6398cffb9c18fd14f8651da7a124f9, {16'd52953, 16'd63986, 16'd11936, 16'd63112, 16'd14928, 16'd50837, 16'd37338, 16'd4251, 16'd23174, 16'd65397, 16'd43818, 16'd44414, 16'd25162, 16'd1821, 16'd8042, 16'd56364, 16'd64064, 16'd27688, 16'd5900, 16'd24673, 16'd26964, 16'd10460, 16'd53651, 16'd3550, 16'd37152, 16'd1653});
	test_expansion(128'hccc9afe91c62edfa3267216816a751c5, {16'd51454, 16'd35452, 16'd26269, 16'd38739, 16'd46793, 16'd56656, 16'd13800, 16'd48482, 16'd58731, 16'd44452, 16'd19736, 16'd3291, 16'd65227, 16'd4214, 16'd25023, 16'd43724, 16'd35592, 16'd1825, 16'd927, 16'd15683, 16'd21096, 16'd40464, 16'd47505, 16'd54890, 16'd54139, 16'd40964});
	test_expansion(128'hb0d561c23e4820079667b7d07e391618, {16'd32762, 16'd8369, 16'd51344, 16'd62447, 16'd47927, 16'd60322, 16'd42886, 16'd42299, 16'd30017, 16'd59529, 16'd48592, 16'd51756, 16'd20142, 16'd9364, 16'd52847, 16'd38032, 16'd6913, 16'd47189, 16'd47684, 16'd41192, 16'd29044, 16'd8026, 16'd41587, 16'd57609, 16'd12493, 16'd27753});
	test_expansion(128'ha7da7ba2ba6e780048c351134673f8c4, {16'd28533, 16'd20637, 16'd34870, 16'd63258, 16'd28677, 16'd35916, 16'd27252, 16'd61421, 16'd50438, 16'd15087, 16'd61895, 16'd24548, 16'd30789, 16'd25070, 16'd27507, 16'd22587, 16'd34951, 16'd22820, 16'd15502, 16'd52617, 16'd195, 16'd1551, 16'd16895, 16'd34821, 16'd24975, 16'd54712});
	test_expansion(128'h6e85b1f97a1b759ab70343539d2fb4ae, {16'd40159, 16'd20362, 16'd21991, 16'd24318, 16'd35726, 16'd7775, 16'd6603, 16'd26649, 16'd27285, 16'd60784, 16'd33386, 16'd5070, 16'd29476, 16'd38060, 16'd46526, 16'd3347, 16'd12951, 16'd47834, 16'd15475, 16'd8423, 16'd12565, 16'd30619, 16'd48803, 16'd26706, 16'd14765, 16'd22889});
	test_expansion(128'h52b05fec741fb32635a614bc0fdcef31, {16'd12538, 16'd117, 16'd58018, 16'd51704, 16'd24438, 16'd9627, 16'd21223, 16'd59928, 16'd4501, 16'd57407, 16'd39451, 16'd56921, 16'd46054, 16'd33501, 16'd28399, 16'd35110, 16'd37173, 16'd29877, 16'd17989, 16'd3598, 16'd27730, 16'd20703, 16'd49446, 16'd51946, 16'd36635, 16'd42430});
	test_expansion(128'h2fa150e2b196ddf4fe9d672a5bcc78b3, {16'd17735, 16'd41846, 16'd15799, 16'd30559, 16'd62021, 16'd42223, 16'd7810, 16'd21463, 16'd23805, 16'd12205, 16'd61505, 16'd43155, 16'd64844, 16'd31436, 16'd52734, 16'd44800, 16'd46906, 16'd4359, 16'd21750, 16'd47988, 16'd52217, 16'd47879, 16'd37178, 16'd4765, 16'd29892, 16'd54157});
	test_expansion(128'h177481fc3bd64806c51db545150a9a74, {16'd4533, 16'd5702, 16'd46551, 16'd52990, 16'd6306, 16'd13773, 16'd17076, 16'd7291, 16'd17273, 16'd14983, 16'd3275, 16'd38692, 16'd15062, 16'd22004, 16'd15437, 16'd11763, 16'd22623, 16'd28645, 16'd45598, 16'd62794, 16'd54449, 16'd29160, 16'd2380, 16'd36645, 16'd9329, 16'd52986});
	test_expansion(128'hfd3489c905813e93086be59338e7cf63, {16'd33983, 16'd48848, 16'd22344, 16'd50695, 16'd44034, 16'd1810, 16'd63519, 16'd27194, 16'd7998, 16'd16045, 16'd51080, 16'd16536, 16'd1359, 16'd11469, 16'd34057, 16'd1895, 16'd26339, 16'd58077, 16'd18275, 16'd3852, 16'd45951, 16'd30083, 16'd1917, 16'd63606, 16'd36001, 16'd57752});
	test_expansion(128'hf886829db746202ee8d8e91f8ec88a2b, {16'd17564, 16'd46353, 16'd15482, 16'd53989, 16'd21369, 16'd26430, 16'd30237, 16'd34092, 16'd65318, 16'd13116, 16'd48739, 16'd53256, 16'd52123, 16'd13701, 16'd16118, 16'd47727, 16'd57837, 16'd45784, 16'd54836, 16'd35497, 16'd34785, 16'd19886, 16'd60313, 16'd5150, 16'd3556, 16'd30857});
	test_expansion(128'h9d579f8065a670d2cff6c5b390476474, {16'd19971, 16'd54099, 16'd64699, 16'd29607, 16'd42307, 16'd38142, 16'd15508, 16'd954, 16'd28679, 16'd52851, 16'd23477, 16'd17499, 16'd22145, 16'd50077, 16'd52377, 16'd13639, 16'd13772, 16'd7634, 16'd16160, 16'd55610, 16'd22682, 16'd5202, 16'd54296, 16'd63387, 16'd3719, 16'd12541});
	test_expansion(128'h7931af086cf01edb66b7684c11bd21bb, {16'd17168, 16'd16124, 16'd7976, 16'd49402, 16'd8843, 16'd41389, 16'd8466, 16'd22227, 16'd54997, 16'd1987, 16'd38031, 16'd56283, 16'd38467, 16'd51254, 16'd57716, 16'd25522, 16'd52291, 16'd49321, 16'd59022, 16'd2688, 16'd46435, 16'd56947, 16'd58295, 16'd28844, 16'd53724, 16'd37115});
	test_expansion(128'h10caf07816f11f22feacef1bacad3130, {16'd65312, 16'd19687, 16'd55911, 16'd39575, 16'd4922, 16'd34420, 16'd11193, 16'd9722, 16'd50507, 16'd56752, 16'd4483, 16'd55869, 16'd16034, 16'd14134, 16'd43527, 16'd41662, 16'd47081, 16'd555, 16'd37209, 16'd38503, 16'd28794, 16'd23978, 16'd17412, 16'd13073, 16'd9492, 16'd3098});
	test_expansion(128'h9b2534b1d277e104001f77f434d091b3, {16'd29914, 16'd34106, 16'd35228, 16'd48117, 16'd61849, 16'd15149, 16'd38108, 16'd56310, 16'd64859, 16'd46114, 16'd9204, 16'd264, 16'd10089, 16'd52800, 16'd14839, 16'd49907, 16'd42401, 16'd22435, 16'd42601, 16'd6859, 16'd28147, 16'd57925, 16'd40320, 16'd52299, 16'd59962, 16'd1387});
	test_expansion(128'h2113a20a697ba4a4e87d7c3917623993, {16'd44549, 16'd23676, 16'd6209, 16'd27500, 16'd41964, 16'd20137, 16'd17626, 16'd42649, 16'd36058, 16'd53392, 16'd38522, 16'd25529, 16'd12959, 16'd21785, 16'd41539, 16'd40708, 16'd7141, 16'd48044, 16'd59070, 16'd40724, 16'd15327, 16'd64285, 16'd12289, 16'd29379, 16'd59138, 16'd31928});
	test_expansion(128'h098bb99b31b2e17f53491c70af464a1e, {16'd19767, 16'd51404, 16'd1365, 16'd25335, 16'd18158, 16'd29168, 16'd40352, 16'd41429, 16'd9933, 16'd12934, 16'd51366, 16'd64049, 16'd12199, 16'd42026, 16'd18333, 16'd18778, 16'd13745, 16'd5834, 16'd49320, 16'd5958, 16'd2753, 16'd48861, 16'd414, 16'd37716, 16'd7943, 16'd23793});
	test_expansion(128'h362981c21c6f5ceba6d40488e12ea202, {16'd34579, 16'd43655, 16'd63249, 16'd40394, 16'd38379, 16'd27851, 16'd22873, 16'd35011, 16'd8939, 16'd38376, 16'd57639, 16'd9341, 16'd42252, 16'd61512, 16'd58744, 16'd20888, 16'd17809, 16'd32749, 16'd51382, 16'd49542, 16'd11453, 16'd10153, 16'd6373, 16'd10823, 16'd30745, 16'd34631});
	test_expansion(128'h5c8afe8f4d39d2f7fd4a6e7e0dbd0629, {16'd17378, 16'd30946, 16'd1984, 16'd64107, 16'd60596, 16'd5943, 16'd57100, 16'd11975, 16'd61334, 16'd5038, 16'd56300, 16'd9876, 16'd8259, 16'd34335, 16'd6899, 16'd54551, 16'd7301, 16'd51868, 16'd39503, 16'd44808, 16'd49606, 16'd186, 16'd38159, 16'd4195, 16'd22473, 16'd4186});
	test_expansion(128'haf1ef975202432529b528ff7e3f16ef2, {16'd13627, 16'd31990, 16'd35806, 16'd62895, 16'd2470, 16'd33291, 16'd42759, 16'd63597, 16'd59710, 16'd39410, 16'd58242, 16'd48863, 16'd29406, 16'd4955, 16'd21056, 16'd10154, 16'd36159, 16'd57232, 16'd63983, 16'd39115, 16'd7124, 16'd61412, 16'd45755, 16'd60283, 16'd38677, 16'd47901});
	test_expansion(128'h1799ad136474c9f76de71edb8cb43761, {16'd62733, 16'd21706, 16'd49594, 16'd52331, 16'd17878, 16'd50195, 16'd39027, 16'd27043, 16'd2736, 16'd56328, 16'd41994, 16'd23229, 16'd37174, 16'd17376, 16'd36716, 16'd45823, 16'd45132, 16'd40197, 16'd57300, 16'd10817, 16'd12097, 16'd19368, 16'd2090, 16'd22455, 16'd24618, 16'd30240});
	test_expansion(128'h74f0e0cdef7e5f4c44fec54f95e9b476, {16'd46675, 16'd56894, 16'd21479, 16'd30454, 16'd40301, 16'd19072, 16'd60987, 16'd36787, 16'd49173, 16'd53720, 16'd3397, 16'd23609, 16'd65057, 16'd46609, 16'd4898, 16'd62848, 16'd48523, 16'd36818, 16'd30176, 16'd36398, 16'd13917, 16'd57722, 16'd56615, 16'd62527, 16'd47561, 16'd57131});
	test_expansion(128'hed75ffcc7e7073065d7142f17dc6b043, {16'd26081, 16'd64505, 16'd27519, 16'd60657, 16'd14175, 16'd5026, 16'd49396, 16'd34705, 16'd36681, 16'd62000, 16'd11884, 16'd65497, 16'd64487, 16'd27611, 16'd50694, 16'd27822, 16'd12472, 16'd50348, 16'd22551, 16'd23682, 16'd15604, 16'd33930, 16'd34722, 16'd57519, 16'd47952, 16'd64317});
	test_expansion(128'hac25a796088260ccfe602093ab4478e2, {16'd56426, 16'd30528, 16'd27978, 16'd53052, 16'd64536, 16'd51843, 16'd16364, 16'd2668, 16'd55713, 16'd52447, 16'd3277, 16'd52284, 16'd38656, 16'd27514, 16'd31673, 16'd12272, 16'd60086, 16'd34347, 16'd52669, 16'd46128, 16'd6796, 16'd51684, 16'd54891, 16'd36379, 16'd40078, 16'd9270});
	test_expansion(128'h478c30be7576491c92d995ba1bbc30d8, {16'd41057, 16'd23019, 16'd24787, 16'd46791, 16'd64712, 16'd50527, 16'd34728, 16'd8968, 16'd46194, 16'd29933, 16'd62176, 16'd11759, 16'd42984, 16'd64417, 16'd30224, 16'd4281, 16'd61835, 16'd61412, 16'd9068, 16'd63913, 16'd63207, 16'd27245, 16'd5048, 16'd30454, 16'd51033, 16'd47722});
	test_expansion(128'heaad72491da9caa4f76766522d2cc4bd, {16'd2385, 16'd28154, 16'd46442, 16'd30050, 16'd4473, 16'd34673, 16'd51634, 16'd17267, 16'd50509, 16'd32963, 16'd27513, 16'd1431, 16'd13594, 16'd8915, 16'd43607, 16'd4959, 16'd3402, 16'd6784, 16'd16632, 16'd46603, 16'd16144, 16'd28252, 16'd26178, 16'd19717, 16'd58714, 16'd8594});
	test_expansion(128'h2dbd28017ef011e28671fe24b3b57a49, {16'd38822, 16'd215, 16'd27262, 16'd33368, 16'd7798, 16'd4801, 16'd13357, 16'd53289, 16'd50463, 16'd61402, 16'd15582, 16'd4766, 16'd43800, 16'd64032, 16'd49276, 16'd34988, 16'd50717, 16'd26014, 16'd12608, 16'd48069, 16'd50346, 16'd44539, 16'd35863, 16'd41098, 16'd11414, 16'd8190});
	test_expansion(128'h9d26382290be7ee1560738dc6a14b411, {16'd53151, 16'd26581, 16'd27443, 16'd24129, 16'd29030, 16'd34549, 16'd2093, 16'd26351, 16'd4520, 16'd27415, 16'd63001, 16'd19962, 16'd48647, 16'd27986, 16'd10146, 16'd53302, 16'd6042, 16'd38855, 16'd1251, 16'd40591, 16'd17613, 16'd9037, 16'd59473, 16'd42856, 16'd39096, 16'd18134});
	test_expansion(128'hc10ffa5bea253d91f5583c79f1d36aaf, {16'd8819, 16'd2643, 16'd22502, 16'd8041, 16'd45922, 16'd5660, 16'd34496, 16'd22508, 16'd51875, 16'd39656, 16'd61796, 16'd15615, 16'd3350, 16'd32844, 16'd27710, 16'd55867, 16'd8983, 16'd23068, 16'd26688, 16'd29553, 16'd19367, 16'd24785, 16'd61451, 16'd3053, 16'd42066, 16'd25729});
	test_expansion(128'hae40870ce3b662bb54081084dfadc0e4, {16'd32558, 16'd49201, 16'd15121, 16'd53406, 16'd60149, 16'd36395, 16'd21069, 16'd10199, 16'd36918, 16'd21270, 16'd32100, 16'd40847, 16'd36532, 16'd52861, 16'd17868, 16'd15599, 16'd6544, 16'd63630, 16'd59512, 16'd46342, 16'd48397, 16'd25910, 16'd701, 16'd22797, 16'd25644, 16'd35696});
	test_expansion(128'h3c1d8a489e7c371c987cab78c441ec4f, {16'd31078, 16'd28631, 16'd39357, 16'd62943, 16'd44011, 16'd62181, 16'd53910, 16'd49080, 16'd26925, 16'd27514, 16'd61380, 16'd28415, 16'd18018, 16'd52270, 16'd13237, 16'd41003, 16'd63353, 16'd15021, 16'd60216, 16'd1711, 16'd37159, 16'd10453, 16'd27858, 16'd65175, 16'd6268, 16'd2692});
	test_expansion(128'hc1777807398d384f57993673cc219961, {16'd42592, 16'd1435, 16'd60320, 16'd6060, 16'd42189, 16'd34862, 16'd47555, 16'd59889, 16'd17853, 16'd17666, 16'd56665, 16'd41517, 16'd10673, 16'd38115, 16'd25648, 16'd62628, 16'd26953, 16'd12829, 16'd25821, 16'd22695, 16'd47733, 16'd14227, 16'd23002, 16'd52549, 16'd32231, 16'd25196});
	test_expansion(128'h99348dba29bf5a89aee00d692f3552fa, {16'd27871, 16'd55608, 16'd54550, 16'd17313, 16'd57458, 16'd48438, 16'd23025, 16'd34091, 16'd7215, 16'd35042, 16'd34563, 16'd34334, 16'd63622, 16'd32290, 16'd29966, 16'd52798, 16'd24571, 16'd17464, 16'd45452, 16'd63053, 16'd32411, 16'd2645, 16'd13846, 16'd64305, 16'd17178, 16'd12910});
	test_expansion(128'h1fdcfc91b55ec996f3cca4a999a7c449, {16'd14084, 16'd61942, 16'd16864, 16'd59529, 16'd27020, 16'd59958, 16'd39933, 16'd11990, 16'd3127, 16'd49079, 16'd1611, 16'd15257, 16'd28431, 16'd56307, 16'd63348, 16'd61000, 16'd18163, 16'd13214, 16'd50674, 16'd63144, 16'd11206, 16'd45074, 16'd55965, 16'd47706, 16'd44956, 16'd59760});
	test_expansion(128'h28f035a0bdbc6d2f3e575b03dfd86758, {16'd28111, 16'd44889, 16'd56932, 16'd18925, 16'd2314, 16'd33560, 16'd43811, 16'd62367, 16'd43279, 16'd60743, 16'd57485, 16'd38641, 16'd19761, 16'd63477, 16'd23193, 16'd9999, 16'd270, 16'd28536, 16'd40215, 16'd10112, 16'd13874, 16'd8076, 16'd39639, 16'd46689, 16'd32259, 16'd65274});
	test_expansion(128'hc4c66a61d6869d7718e1608cdd02a2a6, {16'd38175, 16'd25278, 16'd44260, 16'd25302, 16'd22949, 16'd60689, 16'd16581, 16'd42554, 16'd50961, 16'd61951, 16'd12576, 16'd58426, 16'd51428, 16'd51743, 16'd49466, 16'd21139, 16'd7948, 16'd54134, 16'd23746, 16'd21366, 16'd17359, 16'd23082, 16'd63370, 16'd14992, 16'd45758, 16'd19450});
	test_expansion(128'hd0ef91a9f5c46d794a1c3fe127048348, {16'd26446, 16'd39834, 16'd3364, 16'd1887, 16'd19833, 16'd1381, 16'd12141, 16'd55296, 16'd40048, 16'd31419, 16'd1008, 16'd32306, 16'd36523, 16'd10022, 16'd27797, 16'd12280, 16'd38650, 16'd5218, 16'd20764, 16'd58888, 16'd28407, 16'd57532, 16'd1200, 16'd43331, 16'd53256, 16'd49627});
	test_expansion(128'hbeb76b9ef325e7085213f2a8ea6ee4c3, {16'd47548, 16'd34179, 16'd4456, 16'd38684, 16'd24319, 16'd5005, 16'd52748, 16'd34341, 16'd1655, 16'd15331, 16'd63961, 16'd60620, 16'd40559, 16'd32438, 16'd2574, 16'd42010, 16'd39845, 16'd39475, 16'd28939, 16'd27576, 16'd5928, 16'd10634, 16'd65364, 16'd55816, 16'd40046, 16'd15906});
	test_expansion(128'hc656eaf0d3a4630caa84fb415d8d57f7, {16'd28707, 16'd36330, 16'd24026, 16'd26567, 16'd24632, 16'd56209, 16'd12829, 16'd5613, 16'd52847, 16'd60479, 16'd29262, 16'd51346, 16'd63800, 16'd62530, 16'd19302, 16'd35747, 16'd55493, 16'd9242, 16'd20947, 16'd39513, 16'd36728, 16'd56394, 16'd59319, 16'd61419, 16'd11549, 16'd61774});
	test_expansion(128'ha14c46ff8d469d4d1adad39f507f1609, {16'd52342, 16'd24880, 16'd35225, 16'd8362, 16'd37499, 16'd34626, 16'd52619, 16'd57994, 16'd18506, 16'd61680, 16'd57328, 16'd37282, 16'd20777, 16'd19026, 16'd2649, 16'd49473, 16'd6470, 16'd19396, 16'd11157, 16'd17582, 16'd1685, 16'd34407, 16'd39308, 16'd46151, 16'd29833, 16'd47328});
	test_expansion(128'h38bc84d7d8e395954432ff82b04d7b01, {16'd42601, 16'd9865, 16'd15508, 16'd8488, 16'd41704, 16'd46554, 16'd30563, 16'd10710, 16'd55392, 16'd6351, 16'd4880, 16'd987, 16'd11314, 16'd5516, 16'd7848, 16'd6720, 16'd49263, 16'd48531, 16'd1589, 16'd18697, 16'd52727, 16'd33481, 16'd45656, 16'd42367, 16'd32246, 16'd63902});
	test_expansion(128'hdda2e5a8badae50d874aa170dcd77ecc, {16'd30404, 16'd29609, 16'd17484, 16'd17518, 16'd49620, 16'd56722, 16'd25583, 16'd25506, 16'd23503, 16'd52788, 16'd7107, 16'd28882, 16'd14002, 16'd8691, 16'd14432, 16'd24726, 16'd11182, 16'd42878, 16'd64865, 16'd19841, 16'd6645, 16'd11195, 16'd62984, 16'd52822, 16'd60588, 16'd59653});
	test_expansion(128'hde9383ae702dab6dee4baca2df3b7a76, {16'd8863, 16'd14206, 16'd39696, 16'd56038, 16'd26820, 16'd10449, 16'd26676, 16'd45707, 16'd45439, 16'd28340, 16'd63502, 16'd39988, 16'd9154, 16'd16284, 16'd12306, 16'd9037, 16'd53418, 16'd41455, 16'd39036, 16'd46884, 16'd38246, 16'd40670, 16'd43616, 16'd35642, 16'd31889, 16'd34880});
	test_expansion(128'hdac594e5928dae7e5f9f4332e548c3f8, {16'd31352, 16'd44661, 16'd33770, 16'd48275, 16'd62496, 16'd8400, 16'd6115, 16'd19872, 16'd27412, 16'd1602, 16'd40995, 16'd37073, 16'd56306, 16'd48182, 16'd20910, 16'd17697, 16'd643, 16'd39480, 16'd30032, 16'd36311, 16'd53178, 16'd53132, 16'd36632, 16'd14372, 16'd13438, 16'd2656});
	test_expansion(128'h336efcee2c79014a41619981b1acaeea, {16'd40231, 16'd33248, 16'd2413, 16'd24678, 16'd47725, 16'd53610, 16'd34723, 16'd62239, 16'd33298, 16'd49885, 16'd2441, 16'd34989, 16'd8534, 16'd9339, 16'd64431, 16'd11351, 16'd12010, 16'd56649, 16'd12838, 16'd16774, 16'd32442, 16'd14272, 16'd24302, 16'd38401, 16'd26831, 16'd21877});
	test_expansion(128'hc7d431aa74212b9b9804989cc98ba30a, {16'd34142, 16'd37037, 16'd46074, 16'd61278, 16'd34633, 16'd52283, 16'd31684, 16'd21081, 16'd46856, 16'd41788, 16'd45926, 16'd15603, 16'd37644, 16'd20414, 16'd18444, 16'd11014, 16'd36584, 16'd18243, 16'd8473, 16'd27652, 16'd59379, 16'd3695, 16'd64657, 16'd37154, 16'd7230, 16'd9018});
	test_expansion(128'h56bf24a5475eb2647eca7b762284233f, {16'd51122, 16'd63035, 16'd61253, 16'd31844, 16'd20149, 16'd56415, 16'd54082, 16'd20100, 16'd38271, 16'd65444, 16'd50500, 16'd19035, 16'd28035, 16'd57187, 16'd26036, 16'd16822, 16'd61400, 16'd23822, 16'd47166, 16'd21637, 16'd47184, 16'd47221, 16'd24060, 16'd17073, 16'd10373, 16'd1747});
	test_expansion(128'h9ad4b401ed95568f716d4df26f9a6dd7, {16'd12330, 16'd36996, 16'd51645, 16'd5851, 16'd48621, 16'd18170, 16'd50257, 16'd63257, 16'd23326, 16'd45070, 16'd32861, 16'd35350, 16'd8668, 16'd43619, 16'd1181, 16'd54222, 16'd59415, 16'd46797, 16'd13588, 16'd50202, 16'd35449, 16'd23196, 16'd46209, 16'd64930, 16'd47073, 16'd43037});
	test_expansion(128'h42da8ee74f9891380cdafc34b4fc0f49, {16'd44003, 16'd23729, 16'd56822, 16'd26390, 16'd39967, 16'd60443, 16'd25340, 16'd46538, 16'd62745, 16'd42944, 16'd34464, 16'd30870, 16'd12239, 16'd33778, 16'd11353, 16'd34160, 16'd33262, 16'd32762, 16'd63538, 16'd46611, 16'd38578, 16'd17825, 16'd39484, 16'd58499, 16'd21077, 16'd60290});
	test_expansion(128'h2068d9f19d8c5f269f6e719a69988550, {16'd27065, 16'd21376, 16'd3995, 16'd16913, 16'd42936, 16'd59430, 16'd55845, 16'd37948, 16'd1732, 16'd47982, 16'd44485, 16'd27570, 16'd40123, 16'd59839, 16'd23935, 16'd8119, 16'd12183, 16'd24066, 16'd33924, 16'd34142, 16'd36393, 16'd59799, 16'd41223, 16'd7442, 16'd33499, 16'd2197});
	test_expansion(128'h460b8bc12c161f9a4fcde4391a337091, {16'd2577, 16'd19321, 16'd11178, 16'd40744, 16'd36761, 16'd58389, 16'd4644, 16'd2864, 16'd61681, 16'd50855, 16'd1661, 16'd10275, 16'd51818, 16'd34318, 16'd27580, 16'd6034, 16'd56888, 16'd26707, 16'd23782, 16'd1372, 16'd22685, 16'd2493, 16'd50919, 16'd41022, 16'd60346, 16'd25552});
	test_expansion(128'hfadebe1450b68c8e2b15bcadbb973542, {16'd32729, 16'd52898, 16'd61144, 16'd3245, 16'd29974, 16'd32798, 16'd28756, 16'd31002, 16'd54985, 16'd49363, 16'd50236, 16'd48336, 16'd33082, 16'd14610, 16'd14878, 16'd3229, 16'd26618, 16'd58768, 16'd48330, 16'd50865, 16'd18621, 16'd31601, 16'd37979, 16'd17999, 16'd36286, 16'd57950});
	test_expansion(128'h0a7e46bb0bc1146988dfb92ddc98a924, {16'd30284, 16'd17744, 16'd28686, 16'd45954, 16'd57340, 16'd29145, 16'd36109, 16'd2661, 16'd8214, 16'd46719, 16'd39033, 16'd46203, 16'd27848, 16'd25511, 16'd21871, 16'd49076, 16'd15756, 16'd38496, 16'd19919, 16'd61530, 16'd55427, 16'd4350, 16'd35812, 16'd5957, 16'd60005, 16'd49032});
	test_expansion(128'h43a2a48d495046cd748334284f17f6be, {16'd50014, 16'd53881, 16'd50981, 16'd61473, 16'd19354, 16'd28048, 16'd64529, 16'd53790, 16'd51055, 16'd22429, 16'd23156, 16'd18291, 16'd14684, 16'd53367, 16'd11590, 16'd6985, 16'd39993, 16'd25543, 16'd50361, 16'd28784, 16'd46692, 16'd16790, 16'd64116, 16'd59936, 16'd47231, 16'd22743});
	test_expansion(128'hbeab4caaa241efa5a591d45d5643c09f, {16'd46630, 16'd1180, 16'd18261, 16'd9942, 16'd47618, 16'd5484, 16'd36087, 16'd5270, 16'd11606, 16'd55114, 16'd41126, 16'd10099, 16'd25397, 16'd62601, 16'd9249, 16'd48076, 16'd57261, 16'd51266, 16'd54938, 16'd38298, 16'd3315, 16'd19097, 16'd50602, 16'd29370, 16'd46809, 16'd23805});
	test_expansion(128'h9de862a1463cb4a720debcedfb007ac8, {16'd5197, 16'd50829, 16'd14441, 16'd19583, 16'd38976, 16'd34849, 16'd45731, 16'd18075, 16'd39073, 16'd13393, 16'd16090, 16'd8503, 16'd6542, 16'd18043, 16'd9369, 16'd31028, 16'd2508, 16'd16074, 16'd5023, 16'd25087, 16'd31824, 16'd43625, 16'd60348, 16'd11204, 16'd31440, 16'd45690});
	test_expansion(128'h21bae9b564b3ba253c4bc5a5bfc6d914, {16'd64317, 16'd52035, 16'd42466, 16'd16501, 16'd15455, 16'd15676, 16'd57909, 16'd33448, 16'd52896, 16'd36246, 16'd11902, 16'd58100, 16'd62888, 16'd58749, 16'd53202, 16'd8960, 16'd42725, 16'd4718, 16'd23423, 16'd56033, 16'd46605, 16'd40175, 16'd19022, 16'd28922, 16'd20284, 16'd40949});
	test_expansion(128'hc0c75c9291a10156ec6388b35ac79685, {16'd27088, 16'd40231, 16'd31521, 16'd10804, 16'd55824, 16'd40287, 16'd17952, 16'd28641, 16'd3470, 16'd30721, 16'd58571, 16'd60088, 16'd17984, 16'd42960, 16'd63632, 16'd18622, 16'd62172, 16'd59794, 16'd16242, 16'd17, 16'd3359, 16'd1563, 16'd34988, 16'd18440, 16'd54628, 16'd8740});
	test_expansion(128'h37196a8858ffbdbd8a7a98c74e26e1a6, {16'd49902, 16'd15057, 16'd11556, 16'd27215, 16'd48819, 16'd15690, 16'd47787, 16'd62580, 16'd9623, 16'd9461, 16'd43764, 16'd1454, 16'd43143, 16'd32336, 16'd47144, 16'd58683, 16'd57699, 16'd39103, 16'd3376, 16'd53319, 16'd11886, 16'd26153, 16'd41374, 16'd30900, 16'd38324, 16'd58193});
	test_expansion(128'ha83d75e21b73767601f30d08f2a0dd9e, {16'd56428, 16'd26298, 16'd16924, 16'd13740, 16'd36334, 16'd10619, 16'd59429, 16'd55477, 16'd45580, 16'd7796, 16'd41354, 16'd5227, 16'd17622, 16'd34425, 16'd6338, 16'd55485, 16'd45767, 16'd30662, 16'd20655, 16'd35412, 16'd7006, 16'd22946, 16'd29841, 16'd44745, 16'd57090, 16'd60277});
	test_expansion(128'hd1d2410cbb8a7659fbaa695d0d12e6b5, {16'd34673, 16'd37034, 16'd21125, 16'd62942, 16'd18633, 16'd12997, 16'd60728, 16'd1042, 16'd48797, 16'd29289, 16'd44450, 16'd60999, 16'd42538, 16'd36782, 16'd64837, 16'd52312, 16'd32556, 16'd34839, 16'd1933, 16'd11999, 16'd59371, 16'd42624, 16'd56501, 16'd39082, 16'd7582, 16'd22796});
	test_expansion(128'hf73142f5d82fe14e9ed45badb3fb9319, {16'd20262, 16'd59990, 16'd36885, 16'd64621, 16'd25349, 16'd32241, 16'd44852, 16'd3421, 16'd28303, 16'd52551, 16'd44351, 16'd3972, 16'd46139, 16'd15497, 16'd20276, 16'd14732, 16'd32007, 16'd58843, 16'd65224, 16'd33959, 16'd14863, 16'd29419, 16'd65518, 16'd50752, 16'd26145, 16'd40015});
	test_expansion(128'h5fdb17d2302ce952885e6f73c33ac19d, {16'd19183, 16'd52078, 16'd8369, 16'd38364, 16'd46092, 16'd30502, 16'd7709, 16'd28267, 16'd40067, 16'd27349, 16'd6687, 16'd16679, 16'd61733, 16'd11819, 16'd27068, 16'd48472, 16'd28640, 16'd56863, 16'd23117, 16'd22194, 16'd11503, 16'd41815, 16'd9300, 16'd30236, 16'd47352, 16'd41757});
	test_expansion(128'h5fc2a49d68bec439e3f961d7aa05fd89, {16'd64931, 16'd673, 16'd19511, 16'd16540, 16'd1107, 16'd20052, 16'd4658, 16'd27590, 16'd56388, 16'd44524, 16'd7277, 16'd62902, 16'd13534, 16'd16706, 16'd22298, 16'd25055, 16'd11878, 16'd8989, 16'd21877, 16'd6458, 16'd64406, 16'd32174, 16'd27573, 16'd43739, 16'd6547, 16'd18269});
	test_expansion(128'h42b740c8492eb10b38f43d1cdef84442, {16'd28045, 16'd24356, 16'd18043, 16'd31280, 16'd9178, 16'd8038, 16'd997, 16'd8490, 16'd38703, 16'd50014, 16'd35505, 16'd40703, 16'd60444, 16'd14178, 16'd38722, 16'd44560, 16'd25814, 16'd54480, 16'd40931, 16'd17462, 16'd55744, 16'd9940, 16'd10787, 16'd5161, 16'd15837, 16'd40390});
	test_expansion(128'he4b7a98b9839d6bff9f4ed379fccba3f, {16'd39100, 16'd17491, 16'd53158, 16'd8464, 16'd21061, 16'd24490, 16'd35371, 16'd48437, 16'd5294, 16'd11579, 16'd10112, 16'd15374, 16'd38742, 16'd48189, 16'd2659, 16'd5428, 16'd30583, 16'd9909, 16'd36126, 16'd50798, 16'd59043, 16'd30495, 16'd30614, 16'd5676, 16'd8713, 16'd16105});
	test_expansion(128'hcf617c9d19ffb662617755cf34446069, {16'd12426, 16'd19268, 16'd62079, 16'd59589, 16'd52515, 16'd26702, 16'd53503, 16'd65500, 16'd21185, 16'd58977, 16'd40124, 16'd53681, 16'd49509, 16'd31804, 16'd43008, 16'd49172, 16'd35843, 16'd57030, 16'd28822, 16'd42118, 16'd16458, 16'd52559, 16'd40452, 16'd15612, 16'd23874, 16'd1879});
	test_expansion(128'hcaf4952348bafe8dcb3fbc4fcf49c6db, {16'd34823, 16'd10369, 16'd42761, 16'd63161, 16'd14385, 16'd13885, 16'd45007, 16'd57433, 16'd1698, 16'd8202, 16'd4843, 16'd63369, 16'd1886, 16'd39192, 16'd41402, 16'd2613, 16'd42869, 16'd1602, 16'd42435, 16'd21985, 16'd30376, 16'd32756, 16'd37818, 16'd60292, 16'd50590, 16'd155});
	test_expansion(128'h862224f7eeaa8fdd8352cd623c7ec14c, {16'd55173, 16'd43780, 16'd26045, 16'd48489, 16'd6570, 16'd28004, 16'd47383, 16'd21903, 16'd37194, 16'd8761, 16'd18602, 16'd61885, 16'd38825, 16'd52607, 16'd58861, 16'd38537, 16'd18748, 16'd57401, 16'd42048, 16'd30487, 16'd32890, 16'd54422, 16'd5388, 16'd47331, 16'd32652, 16'd25952});
	test_expansion(128'hbbc935862aad03e76d2a51d20045a171, {16'd45098, 16'd34312, 16'd45600, 16'd47529, 16'd59826, 16'd46272, 16'd5277, 16'd63687, 16'd32773, 16'd51411, 16'd58674, 16'd25478, 16'd33124, 16'd19192, 16'd4519, 16'd4222, 16'd47429, 16'd53749, 16'd26976, 16'd18577, 16'd63060, 16'd13820, 16'd47270, 16'd29734, 16'd4045, 16'd40640});
	test_expansion(128'h75bd8293caee245252ce7ed4dcfbf294, {16'd41511, 16'd28814, 16'd53303, 16'd1313, 16'd50233, 16'd44702, 16'd39972, 16'd63371, 16'd14481, 16'd20109, 16'd16508, 16'd58845, 16'd25893, 16'd41983, 16'd47574, 16'd19984, 16'd46169, 16'd18755, 16'd50765, 16'd15613, 16'd35858, 16'd13309, 16'd59718, 16'd5858, 16'd48877, 16'd33521});
	test_expansion(128'h287ab53ba0ba6e640af4cbd3b3770765, {16'd55585, 16'd23017, 16'd3380, 16'd47041, 16'd17583, 16'd49823, 16'd37107, 16'd3839, 16'd52680, 16'd27935, 16'd28019, 16'd36102, 16'd5348, 16'd30909, 16'd1574, 16'd25632, 16'd1734, 16'd36542, 16'd22925, 16'd43345, 16'd35441, 16'd11724, 16'd54270, 16'd7433, 16'd28068, 16'd49558});
	test_expansion(128'ha06e3ff679dfb7d10612eeee13561190, {16'd33862, 16'd63899, 16'd58836, 16'd25280, 16'd19681, 16'd43335, 16'd19646, 16'd38690, 16'd43149, 16'd50540, 16'd45865, 16'd34545, 16'd49144, 16'd39640, 16'd22470, 16'd33863, 16'd32651, 16'd30335, 16'd49596, 16'd58378, 16'd47685, 16'd55261, 16'd12631, 16'd12103, 16'd46658, 16'd28051});
	test_expansion(128'h84b4ea1c3f793467ac4f2c640502e838, {16'd28978, 16'd19907, 16'd28526, 16'd49026, 16'd34435, 16'd5234, 16'd49268, 16'd49200, 16'd16133, 16'd14772, 16'd39705, 16'd47540, 16'd31885, 16'd50616, 16'd26106, 16'd14706, 16'd31575, 16'd11898, 16'd56236, 16'd54926, 16'd18691, 16'd58078, 16'd61484, 16'd61227, 16'd50299, 16'd55859});
	test_expansion(128'h18ace7a2d71772f14cd40e4648adfd25, {16'd27716, 16'd38905, 16'd56565, 16'd42353, 16'd25312, 16'd51048, 16'd9928, 16'd49458, 16'd6504, 16'd21045, 16'd61597, 16'd1086, 16'd21898, 16'd59840, 16'd29287, 16'd52146, 16'd8573, 16'd8492, 16'd53101, 16'd35406, 16'd56159, 16'd54966, 16'd57535, 16'd45416, 16'd34799, 16'd25524});
	test_expansion(128'hfda6668408a8fcc33da65c212a638856, {16'd59098, 16'd63456, 16'd7267, 16'd30573, 16'd42756, 16'd4843, 16'd22552, 16'd61015, 16'd34916, 16'd46322, 16'd65348, 16'd49438, 16'd55103, 16'd34667, 16'd43144, 16'd29107, 16'd61249, 16'd41542, 16'd25961, 16'd44440, 16'd43469, 16'd34642, 16'd44058, 16'd54009, 16'd65206, 16'd57332});
	test_expansion(128'h6a104e4a71e9275f828174a782cea3e0, {16'd25922, 16'd65091, 16'd33866, 16'd57392, 16'd20635, 16'd53012, 16'd27190, 16'd64897, 16'd6866, 16'd41252, 16'd58912, 16'd23625, 16'd15929, 16'd17459, 16'd30763, 16'd7057, 16'd7551, 16'd61395, 16'd19232, 16'd2917, 16'd56442, 16'd50654, 16'd48589, 16'd37684, 16'd37947, 16'd59067});
	test_expansion(128'hdeab31b44e9453283e4cfa430f9ccca4, {16'd64646, 16'd22803, 16'd34678, 16'd56270, 16'd57730, 16'd21496, 16'd62406, 16'd24251, 16'd58231, 16'd13568, 16'd47431, 16'd48600, 16'd5702, 16'd34567, 16'd40462, 16'd41757, 16'd45638, 16'd39539, 16'd1694, 16'd22740, 16'd39186, 16'd19165, 16'd29721, 16'd26979, 16'd27905, 16'd40217});
	test_expansion(128'hdc58d800d8982163febf533f20557ad6, {16'd44955, 16'd55623, 16'd8991, 16'd1548, 16'd4250, 16'd6532, 16'd59196, 16'd52980, 16'd13223, 16'd58884, 16'd49162, 16'd58637, 16'd57704, 16'd12984, 16'd55018, 16'd55444, 16'd47509, 16'd23413, 16'd19341, 16'd3936, 16'd18690, 16'd6646, 16'd1441, 16'd11518, 16'd7851, 16'd43970});
	test_expansion(128'hb5a4a93bb090d2ee362a70bc2b8f9d7c, {16'd18609, 16'd22166, 16'd62483, 16'd33900, 16'd34289, 16'd32880, 16'd41658, 16'd39863, 16'd58464, 16'd8893, 16'd62210, 16'd46318, 16'd55537, 16'd34117, 16'd32818, 16'd53734, 16'd58554, 16'd61133, 16'd9261, 16'd32979, 16'd31448, 16'd2491, 16'd47463, 16'd32261, 16'd3128, 16'd57140});
	test_expansion(128'he42b5e515797c61b8255a38df6efba54, {16'd30785, 16'd2426, 16'd7969, 16'd43510, 16'd39464, 16'd52267, 16'd37656, 16'd20801, 16'd34754, 16'd18775, 16'd48163, 16'd31826, 16'd21753, 16'd17590, 16'd55143, 16'd23528, 16'd45182, 16'd41117, 16'd41006, 16'd19150, 16'd22954, 16'd8288, 16'd13408, 16'd29641, 16'd24339, 16'd7595});
	test_expansion(128'hd71c764a8838f652c0b1dc4b69284b0f, {16'd35802, 16'd51550, 16'd56815, 16'd63072, 16'd50397, 16'd43447, 16'd35266, 16'd30181, 16'd43286, 16'd61358, 16'd18718, 16'd41168, 16'd14746, 16'd57716, 16'd10317, 16'd43672, 16'd62560, 16'd9799, 16'd23076, 16'd42148, 16'd23807, 16'd25643, 16'd37381, 16'd42760, 16'd53673, 16'd48222});
	test_expansion(128'hb6eb48fd07b7f14565d3394f23b0eade, {16'd38500, 16'd34199, 16'd12748, 16'd26684, 16'd1937, 16'd14269, 16'd64781, 16'd33406, 16'd9563, 16'd27130, 16'd31379, 16'd53331, 16'd51871, 16'd13756, 16'd29029, 16'd6619, 16'd47105, 16'd41840, 16'd7309, 16'd23904, 16'd2154, 16'd53795, 16'd61368, 16'd48929, 16'd19693, 16'd17859});
	test_expansion(128'h71404db1bf324abb0da58f319717fd2b, {16'd46212, 16'd52803, 16'd20407, 16'd61322, 16'd59812, 16'd50233, 16'd45429, 16'd11476, 16'd60481, 16'd16968, 16'd40579, 16'd24495, 16'd31749, 16'd39474, 16'd37953, 16'd28252, 16'd3059, 16'd64235, 16'd54438, 16'd35599, 16'd57557, 16'd22099, 16'd26870, 16'd36133, 16'd16491, 16'd1186});
	test_expansion(128'hf46cd45f10220225b60f670a9bae7c21, {16'd34892, 16'd61903, 16'd36625, 16'd29417, 16'd36496, 16'd29195, 16'd29757, 16'd49197, 16'd10812, 16'd28807, 16'd62205, 16'd46218, 16'd12360, 16'd63149, 16'd12126, 16'd47672, 16'd44237, 16'd61259, 16'd55970, 16'd43120, 16'd2730, 16'd64944, 16'd3210, 16'd41400, 16'd14704, 16'd31497});
	test_expansion(128'h24129d1dcd6434fcf3a6e241f77bdae3, {16'd14574, 16'd61420, 16'd21032, 16'd4999, 16'd49411, 16'd52619, 16'd46208, 16'd56360, 16'd17385, 16'd64436, 16'd4599, 16'd25860, 16'd60479, 16'd18949, 16'd1950, 16'd6041, 16'd5904, 16'd2290, 16'd56984, 16'd776, 16'd8597, 16'd1679, 16'd29640, 16'd21854, 16'd29239, 16'd6578});
	test_expansion(128'h0c73665c615e62bc06d4dcffb8aa7bc6, {16'd54519, 16'd28864, 16'd49230, 16'd3400, 16'd12087, 16'd14655, 16'd49266, 16'd52375, 16'd56994, 16'd65312, 16'd44222, 16'd30359, 16'd32549, 16'd24311, 16'd17102, 16'd5203, 16'd28024, 16'd30386, 16'd36554, 16'd62197, 16'd55085, 16'd13869, 16'd58058, 16'd38172, 16'd34314, 16'd56291});
	test_expansion(128'he1175b04ee0034d95b5c78cfd1e07584, {16'd23775, 16'd45754, 16'd51056, 16'd55610, 16'd50309, 16'd44546, 16'd33685, 16'd56792, 16'd3192, 16'd35908, 16'd43547, 16'd11729, 16'd35298, 16'd18104, 16'd9604, 16'd27218, 16'd34589, 16'd5421, 16'd6948, 16'd47994, 16'd57969, 16'd3898, 16'd49432, 16'd51516, 16'd28851, 16'd20091});
	test_expansion(128'h43bef641d3aa2fd0aa59bebbea3f0f59, {16'd49978, 16'd47453, 16'd49196, 16'd30133, 16'd27802, 16'd5843, 16'd3750, 16'd58100, 16'd23120, 16'd46499, 16'd33556, 16'd28201, 16'd1006, 16'd19138, 16'd65214, 16'd16447, 16'd18891, 16'd39176, 16'd45469, 16'd43877, 16'd41825, 16'd36616, 16'd9032, 16'd17118, 16'd17172, 16'd61458});
	test_expansion(128'ha248ebd1f31a5c836a18146d94670021, {16'd30038, 16'd3984, 16'd10349, 16'd64491, 16'd41031, 16'd65016, 16'd9872, 16'd7036, 16'd57552, 16'd11690, 16'd52020, 16'd31138, 16'd14925, 16'd60711, 16'd19370, 16'd2616, 16'd37261, 16'd16644, 16'd20272, 16'd25397, 16'd15165, 16'd29180, 16'd20013, 16'd45422, 16'd6101, 16'd46071});
	test_expansion(128'he49964489533952927144dd12e106f90, {16'd16101, 16'd47371, 16'd54433, 16'd52284, 16'd25682, 16'd29490, 16'd62085, 16'd57775, 16'd31434, 16'd9815, 16'd12959, 16'd51782, 16'd15729, 16'd24261, 16'd12095, 16'd58828, 16'd52801, 16'd3201, 16'd13498, 16'd48648, 16'd27840, 16'd42288, 16'd6097, 16'd44798, 16'd62045, 16'd11778});
	test_expansion(128'h2eda30314ece87e8590c38400c90be53, {16'd25060, 16'd12009, 16'd35707, 16'd13743, 16'd57793, 16'd172, 16'd44728, 16'd24627, 16'd61623, 16'd60888, 16'd53684, 16'd13189, 16'd14245, 16'd27644, 16'd34595, 16'd35053, 16'd53055, 16'd65041, 16'd34295, 16'd47094, 16'd31019, 16'd34464, 16'd11815, 16'd4901, 16'd21238, 16'd35534});
	test_expansion(128'hf8ce43daf8d22d39b007b0b5a53307e6, {16'd51810, 16'd19194, 16'd36611, 16'd31168, 16'd37178, 16'd666, 16'd52751, 16'd11327, 16'd37361, 16'd2600, 16'd4058, 16'd61672, 16'd33065, 16'd4685, 16'd11872, 16'd50333, 16'd44370, 16'd13614, 16'd3890, 16'd13372, 16'd44538, 16'd48588, 16'd24772, 16'd26013, 16'd2370, 16'd38274});
	test_expansion(128'h51e27493d5399e1d4ae10f7270ec5497, {16'd59469, 16'd28871, 16'd42051, 16'd34280, 16'd10408, 16'd7191, 16'd8674, 16'd8050, 16'd56969, 16'd4181, 16'd23481, 16'd8473, 16'd8332, 16'd9551, 16'd30664, 16'd40293, 16'd1779, 16'd46845, 16'd20849, 16'd3181, 16'd14913, 16'd32855, 16'd55326, 16'd51170, 16'd57157, 16'd29987});
	test_expansion(128'ha42d742d88ade5e67499f922fd171010, {16'd7304, 16'd37438, 16'd48721, 16'd55471, 16'd36631, 16'd26885, 16'd61346, 16'd3600, 16'd61269, 16'd60641, 16'd26300, 16'd24400, 16'd1937, 16'd59147, 16'd36994, 16'd48323, 16'd3260, 16'd43477, 16'd12918, 16'd20101, 16'd54523, 16'd36860, 16'd22934, 16'd15126, 16'd63050, 16'd46091});
	test_expansion(128'h7b959081a002ff505e6eedbc38e5e47f, {16'd64314, 16'd15821, 16'd28072, 16'd13378, 16'd42360, 16'd23817, 16'd45827, 16'd43643, 16'd62206, 16'd59244, 16'd58889, 16'd25291, 16'd4170, 16'd27849, 16'd61237, 16'd51449, 16'd11546, 16'd9950, 16'd63097, 16'd52701, 16'd48009, 16'd16968, 16'd48420, 16'd53845, 16'd921, 16'd41041});
	test_expansion(128'ha8e751f9519ff61d35c0545c447df45b, {16'd29450, 16'd8483, 16'd814, 16'd65328, 16'd63793, 16'd53429, 16'd15523, 16'd15268, 16'd24105, 16'd22414, 16'd26215, 16'd29566, 16'd40287, 16'd33526, 16'd42385, 16'd41315, 16'd47153, 16'd64340, 16'd52496, 16'd29578, 16'd63441, 16'd22037, 16'd50558, 16'd27772, 16'd58786, 16'd35858});
	test_expansion(128'h4daaa1f7c8e2f5185e9441282814df1b, {16'd62748, 16'd4700, 16'd29578, 16'd10553, 16'd49042, 16'd19227, 16'd43015, 16'd64983, 16'd59092, 16'd51193, 16'd507, 16'd63892, 16'd40238, 16'd9188, 16'd56637, 16'd64504, 16'd46719, 16'd36410, 16'd50631, 16'd44804, 16'd46578, 16'd39669, 16'd5744, 16'd44454, 16'd24726, 16'd44302});
	test_expansion(128'hb4c9aae88aec03bf2cfc9e982518d447, {16'd22560, 16'd20407, 16'd11257, 16'd17436, 16'd60428, 16'd4533, 16'd29647, 16'd6884, 16'd18965, 16'd59889, 16'd59067, 16'd19574, 16'd8672, 16'd54533, 16'd9447, 16'd35750, 16'd7037, 16'd64856, 16'd7414, 16'd9117, 16'd18048, 16'd32986, 16'd45542, 16'd45652, 16'd64701, 16'd42648});
	test_expansion(128'hf8ac9096587c3133ffc1e8858ba3dfdf, {16'd8363, 16'd43550, 16'd43833, 16'd41228, 16'd9584, 16'd47427, 16'd25036, 16'd37314, 16'd52102, 16'd51221, 16'd4404, 16'd33439, 16'd44984, 16'd7752, 16'd8098, 16'd20586, 16'd49569, 16'd16041, 16'd56401, 16'd38702, 16'd22818, 16'd29512, 16'd24348, 16'd47171, 16'd62483, 16'd47706});
	test_expansion(128'hf9bd6e57366973f0255e5820737c4eda, {16'd51104, 16'd2093, 16'd63484, 16'd58468, 16'd36329, 16'd7793, 16'd27950, 16'd44509, 16'd16261, 16'd36884, 16'd41446, 16'd12049, 16'd60068, 16'd13013, 16'd64394, 16'd37886, 16'd43761, 16'd29763, 16'd19211, 16'd16438, 16'd17918, 16'd30269, 16'd53689, 16'd33456, 16'd28435, 16'd14980});
	test_expansion(128'haaab59e0c60dc45b4dda2ce9cab9d797, {16'd16308, 16'd738, 16'd42635, 16'd11702, 16'd32996, 16'd10448, 16'd65094, 16'd9910, 16'd10251, 16'd43739, 16'd31246, 16'd64557, 16'd47302, 16'd23467, 16'd8429, 16'd11158, 16'd9089, 16'd60692, 16'd34471, 16'd51060, 16'd1916, 16'd41241, 16'd34456, 16'd6542, 16'd15358, 16'd52204});
	test_expansion(128'h780ac146964cbd5f136a5eb8d7120261, {16'd23528, 16'd57345, 16'd27835, 16'd48203, 16'd14662, 16'd39728, 16'd39242, 16'd28725, 16'd28549, 16'd9890, 16'd25376, 16'd49455, 16'd30062, 16'd3580, 16'd54702, 16'd50606, 16'd36599, 16'd4984, 16'd3416, 16'd62640, 16'd1078, 16'd50289, 16'd40776, 16'd17890, 16'd6606, 16'd5691});
	test_expansion(128'h8a91595b5f22abbc5bdedad1361e7c76, {16'd4878, 16'd43789, 16'd24063, 16'd30117, 16'd36537, 16'd24098, 16'd58032, 16'd51018, 16'd47135, 16'd37439, 16'd14198, 16'd8356, 16'd41802, 16'd29027, 16'd55696, 16'd47121, 16'd55120, 16'd18077, 16'd37382, 16'd63322, 16'd64864, 16'd57260, 16'd21343, 16'd52997, 16'd17544, 16'd30087});
	test_expansion(128'he5ad55f89b38a753211e2feaf65d2574, {16'd4984, 16'd12968, 16'd13779, 16'd34210, 16'd43280, 16'd27678, 16'd40119, 16'd63512, 16'd9022, 16'd652, 16'd60958, 16'd55044, 16'd40412, 16'd61549, 16'd24262, 16'd42305, 16'd20326, 16'd53113, 16'd26904, 16'd36750, 16'd22083, 16'd31106, 16'd51684, 16'd32011, 16'd31567, 16'd17765});
	test_expansion(128'h7b7f3e64d01111d1e89c94f58316e97b, {16'd56745, 16'd60581, 16'd43379, 16'd43517, 16'd11975, 16'd51244, 16'd42771, 16'd23408, 16'd20746, 16'd50327, 16'd45719, 16'd20612, 16'd8943, 16'd3226, 16'd42908, 16'd43979, 16'd22404, 16'd41058, 16'd36419, 16'd26808, 16'd39054, 16'd36494, 16'd20543, 16'd49393, 16'd61882, 16'd35777});
	test_expansion(128'h882810cfd5af5af72d0c0c4dda52a7b9, {16'd18797, 16'd50807, 16'd1294, 16'd45585, 16'd52863, 16'd27602, 16'd58867, 16'd32774, 16'd56128, 16'd64226, 16'd63663, 16'd1332, 16'd22937, 16'd9892, 16'd53507, 16'd12020, 16'd52542, 16'd37366, 16'd46800, 16'd51236, 16'd17054, 16'd51981, 16'd2491, 16'd14701, 16'd30889, 16'd461});
	test_expansion(128'hfc7ad426e300bbe9fab4877033bfb839, {16'd37963, 16'd11890, 16'd15391, 16'd56147, 16'd58557, 16'd53219, 16'd54313, 16'd48376, 16'd6844, 16'd32791, 16'd11874, 16'd5965, 16'd27649, 16'd55476, 16'd11877, 16'd921, 16'd48847, 16'd49871, 16'd4792, 16'd24733, 16'd1793, 16'd56739, 16'd49021, 16'd57314, 16'd18681, 16'd45855});
	test_expansion(128'hea797fda6cba3d528b8aeaadc3f28f4c, {16'd42996, 16'd41548, 16'd17521, 16'd21289, 16'd34556, 16'd53230, 16'd9470, 16'd43990, 16'd59690, 16'd61377, 16'd50509, 16'd44661, 16'd34226, 16'd9411, 16'd49521, 16'd1121, 16'd13430, 16'd14326, 16'd57477, 16'd6323, 16'd4216, 16'd29370, 16'd9184, 16'd18321, 16'd19708, 16'd33016});
	test_expansion(128'h8a161add77908d884ca67478d95be9ee, {16'd11525, 16'd32311, 16'd26439, 16'd44918, 16'd18638, 16'd31598, 16'd53667, 16'd64202, 16'd32225, 16'd42289, 16'd245, 16'd2959, 16'd36809, 16'd26881, 16'd12262, 16'd7516, 16'd59631, 16'd34257, 16'd47758, 16'd9646, 16'd10865, 16'd46287, 16'd54812, 16'd23876, 16'd25295, 16'd27676});
	test_expansion(128'h5b26a3f5feb58e2842e00e25519eb711, {16'd54180, 16'd44736, 16'd6262, 16'd2661, 16'd5889, 16'd48282, 16'd18149, 16'd18917, 16'd45374, 16'd49265, 16'd16308, 16'd61834, 16'd9742, 16'd23964, 16'd24423, 16'd50286, 16'd33960, 16'd9244, 16'd49250, 16'd118, 16'd19740, 16'd5252, 16'd28680, 16'd1377, 16'd40539, 16'd55179});
	test_expansion(128'hd5f4c14cc56412bb0b2ee9fd00930210, {16'd38110, 16'd1713, 16'd2354, 16'd10715, 16'd39183, 16'd4494, 16'd33821, 16'd56889, 16'd36009, 16'd52679, 16'd30165, 16'd5119, 16'd17488, 16'd39797, 16'd41441, 16'd27329, 16'd37665, 16'd3528, 16'd27399, 16'd65076, 16'd8295, 16'd41610, 16'd44161, 16'd33249, 16'd45198, 16'd34205});
	test_expansion(128'haf4e7171a5239bfc9e2d608a38909932, {16'd6705, 16'd43783, 16'd6557, 16'd59810, 16'd59174, 16'd20784, 16'd43071, 16'd51436, 16'd29907, 16'd26521, 16'd2969, 16'd49432, 16'd19301, 16'd13958, 16'd56040, 16'd35873, 16'd13998, 16'd10434, 16'd7929, 16'd30277, 16'd26874, 16'd50884, 16'd21773, 16'd25305, 16'd57004, 16'd18897});
	test_expansion(128'h0b47711d42846073aaa38fa660fc24d6, {16'd21806, 16'd24011, 16'd17053, 16'd59870, 16'd61791, 16'd49876, 16'd53165, 16'd23020, 16'd44769, 16'd27836, 16'd1166, 16'd45082, 16'd13442, 16'd6568, 16'd49653, 16'd40561, 16'd14590, 16'd60926, 16'd7878, 16'd45568, 16'd44284, 16'd11444, 16'd26714, 16'd62187, 16'd26492, 16'd61983});
	test_expansion(128'hf72b67db98ea4119fcc8f3748aa909c1, {16'd26000, 16'd17325, 16'd30570, 16'd29960, 16'd49472, 16'd49911, 16'd31545, 16'd63589, 16'd23429, 16'd16190, 16'd30342, 16'd51539, 16'd45615, 16'd14014, 16'd2035, 16'd40450, 16'd28624, 16'd20971, 16'd25391, 16'd20700, 16'd51903, 16'd25765, 16'd11738, 16'd53090, 16'd12782, 16'd50119});
	test_expansion(128'h4656215ff3fda9b5d81bca9f1f455f27, {16'd14242, 16'd6966, 16'd56580, 16'd43594, 16'd40432, 16'd56279, 16'd38988, 16'd9383, 16'd28870, 16'd14204, 16'd30671, 16'd42349, 16'd65031, 16'd6850, 16'd63434, 16'd38855, 16'd35014, 16'd8436, 16'd36105, 16'd36461, 16'd28678, 16'd7816, 16'd32977, 16'd1864, 16'd1649, 16'd24523});
	test_expansion(128'hc3a51a035c4be2c1cf33c770b9b0ba6b, {16'd15680, 16'd17860, 16'd36653, 16'd53722, 16'd59658, 16'd52628, 16'd31768, 16'd43226, 16'd30543, 16'd7326, 16'd61761, 16'd61318, 16'd24644, 16'd53752, 16'd58618, 16'd20268, 16'd1625, 16'd24117, 16'd19942, 16'd55203, 16'd19743, 16'd47730, 16'd21530, 16'd5906, 16'd39831, 16'd18838});
	test_expansion(128'h89a221122e85d7b58a8a8dc56ebab4e1, {16'd6605, 16'd41431, 16'd15105, 16'd40360, 16'd34141, 16'd39033, 16'd15554, 16'd1180, 16'd12411, 16'd35314, 16'd64159, 16'd56670, 16'd63504, 16'd39189, 16'd6037, 16'd54481, 16'd49792, 16'd40831, 16'd24934, 16'd46223, 16'd22605, 16'd62192, 16'd12670, 16'd13980, 16'd60321, 16'd7535});
	test_expansion(128'hdbf2461e8815ce4c8b6fefdbcf36cb54, {16'd690, 16'd3079, 16'd53034, 16'd32818, 16'd51272, 16'd23811, 16'd21925, 16'd60194, 16'd27221, 16'd50587, 16'd20474, 16'd50336, 16'd37016, 16'd56761, 16'd3779, 16'd28429, 16'd27363, 16'd21781, 16'd65437, 16'd5940, 16'd54650, 16'd15416, 16'd51070, 16'd61651, 16'd52330, 16'd6319});
	test_expansion(128'h60602ba74049e634ab40edc25c1ca4cb, {16'd4195, 16'd31084, 16'd28430, 16'd34765, 16'd41843, 16'd32515, 16'd15105, 16'd42431, 16'd3311, 16'd8150, 16'd12987, 16'd25737, 16'd31759, 16'd15001, 16'd25709, 16'd20879, 16'd27821, 16'd30022, 16'd37042, 16'd23751, 16'd44425, 16'd48405, 16'd53579, 16'd58481, 16'd28030, 16'd13911});
	test_expansion(128'h256162dd6c743833646ebd2b40fecad1, {16'd27694, 16'd4152, 16'd44365, 16'd19897, 16'd53091, 16'd53875, 16'd48654, 16'd38820, 16'd3611, 16'd55678, 16'd25726, 16'd36879, 16'd11659, 16'd33544, 16'd35009, 16'd34297, 16'd33511, 16'd12852, 16'd39133, 16'd7235, 16'd52064, 16'd34115, 16'd43340, 16'd37307, 16'd58006, 16'd40081});
	test_expansion(128'he9e883472f0c98e049fe0be5850492a3, {16'd25438, 16'd56338, 16'd38037, 16'd51260, 16'd29445, 16'd57806, 16'd37427, 16'd48587, 16'd23577, 16'd908, 16'd33679, 16'd34965, 16'd10736, 16'd38612, 16'd47961, 16'd31183, 16'd17627, 16'd30604, 16'd44207, 16'd47371, 16'd17877, 16'd39229, 16'd45736, 16'd10402, 16'd51646, 16'd24837});
	test_expansion(128'h7e78774728fabedc0c3c024eba6fff9c, {16'd37934, 16'd55225, 16'd17894, 16'd48904, 16'd16439, 16'd49164, 16'd4195, 16'd14486, 16'd42870, 16'd37232, 16'd45552, 16'd18308, 16'd56802, 16'd31267, 16'd45742, 16'd31131, 16'd26227, 16'd53609, 16'd3449, 16'd38409, 16'd62890, 16'd35315, 16'd35539, 16'd63847, 16'd31127, 16'd13130});
	test_expansion(128'hebf563a6e75e84cd3f8ed03b21b1ff65, {16'd8956, 16'd51438, 16'd46247, 16'd30581, 16'd56147, 16'd13017, 16'd52395, 16'd32073, 16'd54030, 16'd63567, 16'd48556, 16'd8813, 16'd12165, 16'd60552, 16'd684, 16'd57767, 16'd59041, 16'd20950, 16'd21614, 16'd4872, 16'd16763, 16'd928, 16'd45163, 16'd50679, 16'd13110, 16'd55439});
	test_expansion(128'h436ff4fcd3671a0ece89f1c3af700d15, {16'd57766, 16'd23841, 16'd65129, 16'd34247, 16'd47380, 16'd50711, 16'd20623, 16'd18731, 16'd28522, 16'd19494, 16'd13072, 16'd47689, 16'd10619, 16'd50085, 16'd26425, 16'd63851, 16'd48598, 16'd16071, 16'd62866, 16'd13583, 16'd33004, 16'd60258, 16'd20523, 16'd46300, 16'd52134, 16'd8556});
	test_expansion(128'h95d5cc8b133bc68913f13974c8bdb8e3, {16'd9525, 16'd46380, 16'd55992, 16'd51629, 16'd6818, 16'd11765, 16'd31122, 16'd45662, 16'd46000, 16'd45497, 16'd45446, 16'd29514, 16'd47728, 16'd23674, 16'd63296, 16'd51252, 16'd14872, 16'd53657, 16'd60985, 16'd12271, 16'd45102, 16'd23838, 16'd30789, 16'd43298, 16'd62671, 16'd26636});
	test_expansion(128'h7d54274ce47b6b94b0776aee7d97d795, {16'd25434, 16'd26380, 16'd50725, 16'd11605, 16'd20643, 16'd9743, 16'd50397, 16'd63852, 16'd41986, 16'd3310, 16'd7685, 16'd53352, 16'd34938, 16'd49791, 16'd36970, 16'd10854, 16'd6369, 16'd51972, 16'd65118, 16'd41798, 16'd36394, 16'd28348, 16'd17532, 16'd43989, 16'd50494, 16'd43438});
	test_expansion(128'hd18264554be8f939e3b2b57ecdfc5145, {16'd61545, 16'd35818, 16'd49651, 16'd63231, 16'd47685, 16'd56049, 16'd49080, 16'd18874, 16'd36312, 16'd15437, 16'd60712, 16'd40143, 16'd23533, 16'd63395, 16'd39657, 16'd44922, 16'd44068, 16'd12246, 16'd30308, 16'd37207, 16'd56089, 16'd7949, 16'd63003, 16'd28158, 16'd49353, 16'd13630});
	test_expansion(128'hae3e8d62144b8a4601508d8e233d04f0, {16'd30095, 16'd38870, 16'd17213, 16'd9976, 16'd40694, 16'd2574, 16'd57921, 16'd54631, 16'd33831, 16'd15244, 16'd54093, 16'd52500, 16'd2743, 16'd13334, 16'd31993, 16'd32948, 16'd47077, 16'd8479, 16'd31148, 16'd47539, 16'd49860, 16'd11867, 16'd24881, 16'd24651, 16'd5409, 16'd32079});
	test_expansion(128'h2e79af2c0c8bd5c9d20672ffe88766bc, {16'd64279, 16'd48086, 16'd35567, 16'd20919, 16'd15942, 16'd56735, 16'd48428, 16'd51128, 16'd62191, 16'd28008, 16'd61657, 16'd2752, 16'd56581, 16'd20959, 16'd9089, 16'd583, 16'd36282, 16'd32692, 16'd55423, 16'd3304, 16'd33101, 16'd61804, 16'd37253, 16'd8671, 16'd15729, 16'd39984});
	test_expansion(128'hf4c59d8f28ffcb1d2ac04723121434eb, {16'd33948, 16'd43488, 16'd34764, 16'd56498, 16'd23916, 16'd16077, 16'd1777, 16'd17735, 16'd9954, 16'd831, 16'd54399, 16'd46265, 16'd16802, 16'd30573, 16'd58489, 16'd28512, 16'd24920, 16'd63172, 16'd20798, 16'd561, 16'd36133, 16'd45972, 16'd60919, 16'd6608, 16'd18317, 16'd32931});
	test_expansion(128'h93672ec2b39224086dc05f6dbcc7dc50, {16'd55007, 16'd25045, 16'd21114, 16'd29417, 16'd30077, 16'd25722, 16'd51331, 16'd30457, 16'd43531, 16'd33011, 16'd8536, 16'd56671, 16'd5272, 16'd60842, 16'd5812, 16'd23594, 16'd47853, 16'd19518, 16'd7545, 16'd46518, 16'd46409, 16'd63015, 16'd41321, 16'd58359, 16'd40450, 16'd13883});
	test_expansion(128'ha7dac9be5345e1756fc55a1a8cfff9a9, {16'd16278, 16'd34420, 16'd18191, 16'd53759, 16'd40341, 16'd43834, 16'd24019, 16'd44282, 16'd22383, 16'd29269, 16'd59098, 16'd12450, 16'd32383, 16'd22350, 16'd21303, 16'd55957, 16'd22600, 16'd40463, 16'd7462, 16'd32697, 16'd26681, 16'd18143, 16'd1157, 16'd13661, 16'd21748, 16'd42171});
	test_expansion(128'he95742bf6ca82a3a9cca98cb599fc15d, {16'd53355, 16'd18752, 16'd14144, 16'd43165, 16'd39468, 16'd12290, 16'd53533, 16'd22359, 16'd55676, 16'd51121, 16'd16193, 16'd473, 16'd54011, 16'd10540, 16'd27612, 16'd7820, 16'd43636, 16'd60124, 16'd22420, 16'd14278, 16'd60917, 16'd25953, 16'd44078, 16'd27021, 16'd60091, 16'd52216});
	test_expansion(128'hbffc1657544233f39550c163ebacd0bb, {16'd44441, 16'd17096, 16'd34385, 16'd5824, 16'd33850, 16'd42402, 16'd43878, 16'd8521, 16'd37150, 16'd55039, 16'd12873, 16'd14255, 16'd36458, 16'd34677, 16'd35862, 16'd22596, 16'd62408, 16'd39518, 16'd25023, 16'd63592, 16'd53480, 16'd59799, 16'd54874, 16'd43234, 16'd54426, 16'd62845});
	test_expansion(128'h1e8ea2a9edc1e7a104cf55f0579709fe, {16'd14330, 16'd10980, 16'd8289, 16'd63950, 16'd1650, 16'd9744, 16'd19971, 16'd40504, 16'd60335, 16'd34179, 16'd16971, 16'd39185, 16'd21509, 16'd51403, 16'd20626, 16'd30738, 16'd43955, 16'd61497, 16'd9861, 16'd63205, 16'd40682, 16'd4347, 16'd57922, 16'd13922, 16'd28676, 16'd35663});
	test_expansion(128'h0afed7f266e98b47a5f9df4b7bc4850f, {16'd38913, 16'd38407, 16'd60292, 16'd26966, 16'd35950, 16'd32858, 16'd20068, 16'd19685, 16'd52901, 16'd64707, 16'd33532, 16'd36254, 16'd3808, 16'd16385, 16'd600, 16'd22580, 16'd5085, 16'd32673, 16'd34952, 16'd11908, 16'd16267, 16'd47559, 16'd46956, 16'd19657, 16'd186, 16'd64097});
	test_expansion(128'hfa02c47fa4a54ea6cfbf52f948ee82d3, {16'd22476, 16'd38146, 16'd61546, 16'd23936, 16'd53479, 16'd17805, 16'd49979, 16'd25334, 16'd7438, 16'd31361, 16'd19665, 16'd31767, 16'd8114, 16'd36834, 16'd44086, 16'd27522, 16'd61074, 16'd61991, 16'd20914, 16'd38469, 16'd4528, 16'd61394, 16'd44166, 16'd18867, 16'd36563, 16'd26840});
	test_expansion(128'h8df3f174fa187b08034f9fb0bb40b307, {16'd7843, 16'd41960, 16'd32980, 16'd62103, 16'd14239, 16'd11706, 16'd51906, 16'd19050, 16'd24197, 16'd47462, 16'd55613, 16'd27116, 16'd11580, 16'd46070, 16'd43437, 16'd11207, 16'd12149, 16'd49556, 16'd47567, 16'd30338, 16'd57399, 16'd24049, 16'd65193, 16'd35247, 16'd45863, 16'd17422});
	test_expansion(128'h12d1f607102e2827bdf33e505d400733, {16'd46790, 16'd8415, 16'd33306, 16'd61108, 16'd6380, 16'd32470, 16'd55516, 16'd61575, 16'd820, 16'd40289, 16'd29910, 16'd13307, 16'd11075, 16'd54336, 16'd49237, 16'd47288, 16'd40893, 16'd45475, 16'd3095, 16'd20543, 16'd39647, 16'd57174, 16'd48934, 16'd4073, 16'd13129, 16'd20445});
	test_expansion(128'hdac8cb4a580bdaca045f31925824436e, {16'd41350, 16'd25610, 16'd29020, 16'd1453, 16'd16172, 16'd36710, 16'd8509, 16'd60920, 16'd35264, 16'd62136, 16'd12570, 16'd21882, 16'd37446, 16'd45374, 16'd8798, 16'd60675, 16'd33341, 16'd41828, 16'd37426, 16'd18035, 16'd35540, 16'd60070, 16'd56444, 16'd13267, 16'd23887, 16'd41299});
	test_expansion(128'hf3fc019b3890cc85a3313cb684b06c9d, {16'd5585, 16'd55284, 16'd523, 16'd53805, 16'd29319, 16'd52441, 16'd62814, 16'd56537, 16'd46864, 16'd15861, 16'd60966, 16'd2571, 16'd23405, 16'd8499, 16'd43923, 16'd65270, 16'd47573, 16'd9288, 16'd56252, 16'd28829, 16'd688, 16'd46755, 16'd48170, 16'd21588, 16'd7051, 16'd14856});
	test_expansion(128'h29aad0fb4cf9255045de2819308e7aef, {16'd60501, 16'd17328, 16'd28354, 16'd19212, 16'd39146, 16'd63458, 16'd944, 16'd58703, 16'd4303, 16'd22326, 16'd41064, 16'd33175, 16'd53513, 16'd34930, 16'd37436, 16'd23245, 16'd58420, 16'd52507, 16'd10875, 16'd20141, 16'd30521, 16'd37964, 16'd34632, 16'd48169, 16'd47008, 16'd49720});
	test_expansion(128'hba8f2e9692eae738da5148bc2c5ba208, {16'd39133, 16'd20525, 16'd47919, 16'd8810, 16'd36509, 16'd30397, 16'd62490, 16'd42867, 16'd41932, 16'd63673, 16'd4287, 16'd25957, 16'd19762, 16'd19350, 16'd43839, 16'd50237, 16'd58442, 16'd28452, 16'd46075, 16'd59125, 16'd34958, 16'd62314, 16'd6809, 16'd15204, 16'd44716, 16'd41122});
	test_expansion(128'h85d92407ed38cefb41f8ac95cfb8263e, {16'd18497, 16'd22074, 16'd828, 16'd61615, 16'd29940, 16'd30228, 16'd63110, 16'd3810, 16'd20580, 16'd60923, 16'd6575, 16'd21900, 16'd27924, 16'd43595, 16'd21375, 16'd24302, 16'd12224, 16'd22818, 16'd53756, 16'd49921, 16'd15383, 16'd38504, 16'd14027, 16'd57741, 16'd60690, 16'd16945});
	test_expansion(128'h4b75464248d61a3f3079a9743c355c22, {16'd2814, 16'd57740, 16'd53324, 16'd5321, 16'd27536, 16'd24997, 16'd56517, 16'd27907, 16'd45498, 16'd29670, 16'd28601, 16'd41226, 16'd31266, 16'd21993, 16'd25271, 16'd21523, 16'd44453, 16'd58442, 16'd53494, 16'd12791, 16'd21116, 16'd47658, 16'd45315, 16'd49025, 16'd15275, 16'd27795});
	test_expansion(128'h0b9a206d81b8b484fe64a76ed24225fe, {16'd40422, 16'd51044, 16'd31291, 16'd61836, 16'd11142, 16'd19742, 16'd59275, 16'd25796, 16'd16433, 16'd488, 16'd61037, 16'd22091, 16'd60231, 16'd35589, 16'd60245, 16'd44405, 16'd8212, 16'd53339, 16'd263, 16'd22370, 16'd36565, 16'd50323, 16'd18372, 16'd33913, 16'd2715, 16'd57265});
	test_expansion(128'ha3ddca761ad17fe0c591ea7da8d8eab3, {16'd21583, 16'd47216, 16'd10161, 16'd28347, 16'd45658, 16'd56090, 16'd762, 16'd44449, 16'd58194, 16'd13423, 16'd60079, 16'd22591, 16'd29639, 16'd64045, 16'd23003, 16'd482, 16'd12663, 16'd11435, 16'd3081, 16'd27339, 16'd25819, 16'd28490, 16'd48906, 16'd60335, 16'd29981, 16'd49235});
	test_expansion(128'h74d80154970d6231bfaa543ba7aabdb1, {16'd13010, 16'd32661, 16'd33407, 16'd3630, 16'd1352, 16'd46663, 16'd45128, 16'd60064, 16'd4548, 16'd51616, 16'd17229, 16'd49779, 16'd59687, 16'd9867, 16'd3883, 16'd22199, 16'd61429, 16'd49197, 16'd43182, 16'd6038, 16'd56025, 16'd44186, 16'd4736, 16'd34162, 16'd22847, 16'd15734});
	test_expansion(128'hb04eb0c2802e068f50df54930fda1bb7, {16'd32952, 16'd1303, 16'd47276, 16'd56045, 16'd60935, 16'd2422, 16'd12331, 16'd18699, 16'd26176, 16'd19764, 16'd39657, 16'd37559, 16'd54787, 16'd16045, 16'd26830, 16'd62492, 16'd49922, 16'd59787, 16'd54844, 16'd60489, 16'd13155, 16'd54530, 16'd60779, 16'd44245, 16'd29825, 16'd29569});
	test_expansion(128'haf1314fc26fcc23c81c5dcf40f04da40, {16'd16475, 16'd58898, 16'd19399, 16'd44445, 16'd16658, 16'd18355, 16'd45699, 16'd36982, 16'd36965, 16'd37036, 16'd573, 16'd9039, 16'd4729, 16'd49175, 16'd23391, 16'd9585, 16'd11248, 16'd42137, 16'd9970, 16'd13163, 16'd45187, 16'd39201, 16'd23781, 16'd44280, 16'd15225, 16'd27788});
	test_expansion(128'h5c17fd41b8c77f2bd09fe45f10a150ae, {16'd14098, 16'd32168, 16'd23895, 16'd53878, 16'd54372, 16'd6943, 16'd37328, 16'd39531, 16'd19504, 16'd29779, 16'd14191, 16'd46473, 16'd44721, 16'd37494, 16'd10799, 16'd49662, 16'd38543, 16'd50789, 16'd28004, 16'd44016, 16'd53511, 16'd28145, 16'd37151, 16'd6863, 16'd993, 16'd3514});
	test_expansion(128'hec38ddafc22fb98ad59bf35868d77fd6, {16'd10018, 16'd44358, 16'd55937, 16'd57712, 16'd16423, 16'd36010, 16'd4103, 16'd19391, 16'd25759, 16'd51806, 16'd43774, 16'd31253, 16'd26184, 16'd13778, 16'd1197, 16'd16856, 16'd51381, 16'd43039, 16'd11743, 16'd15376, 16'd39772, 16'd28574, 16'd50615, 16'd45021, 16'd43666, 16'd49549});
	test_expansion(128'h9cbb45335038d00d2b3055c551a726cb, {16'd18294, 16'd36708, 16'd14286, 16'd36610, 16'd8341, 16'd37119, 16'd55534, 16'd12, 16'd55779, 16'd48996, 16'd25873, 16'd19577, 16'd20998, 16'd9415, 16'd17995, 16'd20358, 16'd57472, 16'd48585, 16'd57244, 16'd57671, 16'd10717, 16'd57234, 16'd25252, 16'd55878, 16'd58852, 16'd59436});
	test_expansion(128'hbce81b5c39f68c163ebae482e99f40f3, {16'd39176, 16'd26159, 16'd47889, 16'd29837, 16'd31995, 16'd18699, 16'd64512, 16'd9135, 16'd6408, 16'd32736, 16'd15224, 16'd31729, 16'd23844, 16'd47544, 16'd2423, 16'd7347, 16'd34013, 16'd5417, 16'd50219, 16'd35603, 16'd10682, 16'd43709, 16'd31413, 16'd29576, 16'd62557, 16'd63704});
	test_expansion(128'h7a8311fc28dc0689ae389cd42ef499ef, {16'd27664, 16'd21522, 16'd28873, 16'd63440, 16'd3467, 16'd37024, 16'd40317, 16'd48602, 16'd14488, 16'd62030, 16'd7942, 16'd50829, 16'd5265, 16'd65102, 16'd62756, 16'd6485, 16'd5729, 16'd47933, 16'd16798, 16'd19743, 16'd1590, 16'd12880, 16'd64326, 16'd195, 16'd11950, 16'd56532});
	test_expansion(128'hae9b183b6b156eb423b25e26150d540d, {16'd32793, 16'd1132, 16'd56463, 16'd22196, 16'd41909, 16'd59597, 16'd47608, 16'd62054, 16'd18293, 16'd17033, 16'd27579, 16'd27151, 16'd15164, 16'd39535, 16'd9101, 16'd49947, 16'd31871, 16'd46388, 16'd35925, 16'd8077, 16'd41632, 16'd47078, 16'd43542, 16'd38895, 16'd45777, 16'd47280});
	test_expansion(128'h4fd4d1627b3291fe5cd0552573637785, {16'd25923, 16'd25723, 16'd7851, 16'd8531, 16'd19004, 16'd49374, 16'd57663, 16'd44146, 16'd53037, 16'd57547, 16'd57019, 16'd37167, 16'd39425, 16'd20209, 16'd17536, 16'd6972, 16'd15307, 16'd60615, 16'd46520, 16'd47174, 16'd41017, 16'd1026, 16'd18373, 16'd43315, 16'd13388, 16'd39749});
	test_expansion(128'h474c1d66a6e495e88fc1977922832705, {16'd37233, 16'd40269, 16'd50972, 16'd11110, 16'd37079, 16'd50198, 16'd6974, 16'd16620, 16'd11088, 16'd911, 16'd53773, 16'd24836, 16'd7194, 16'd18453, 16'd30259, 16'd26094, 16'd40943, 16'd38647, 16'd23247, 16'd19806, 16'd24073, 16'd24083, 16'd49810, 16'd22982, 16'd40704, 16'd506});
	test_expansion(128'h90b8aff8006c1050d291b2ac4cd2a344, {16'd34796, 16'd18541, 16'd4580, 16'd39783, 16'd21294, 16'd59655, 16'd49068, 16'd1244, 16'd46318, 16'd43284, 16'd6213, 16'd41765, 16'd57852, 16'd12196, 16'd6290, 16'd32784, 16'd36125, 16'd11292, 16'd59935, 16'd57718, 16'd55005, 16'd57637, 16'd59231, 16'd39764, 16'd61611, 16'd34558});
	test_expansion(128'h769613864b1e947441aeb029f9f95800, {16'd26081, 16'd8325, 16'd37543, 16'd64219, 16'd9514, 16'd31667, 16'd1356, 16'd15612, 16'd53335, 16'd42487, 16'd48059, 16'd18354, 16'd45375, 16'd7483, 16'd57732, 16'd33468, 16'd30415, 16'd20348, 16'd572, 16'd61573, 16'd63787, 16'd13906, 16'd28746, 16'd35897, 16'd26251, 16'd35549});
	test_expansion(128'h25e85cdc419e193f341b0de9e0ac31da, {16'd659, 16'd22121, 16'd24197, 16'd16396, 16'd62497, 16'd57716, 16'd56801, 16'd26171, 16'd15107, 16'd28289, 16'd54590, 16'd49071, 16'd16743, 16'd52260, 16'd11432, 16'd22102, 16'd65492, 16'd59122, 16'd4320, 16'd16542, 16'd58952, 16'd22762, 16'd13633, 16'd15872, 16'd20059, 16'd32292});
	test_expansion(128'h85c8be272286b9e7986c2afc976a3ffb, {16'd30507, 16'd57138, 16'd18581, 16'd14031, 16'd31124, 16'd57572, 16'd15373, 16'd41906, 16'd29760, 16'd24217, 16'd56379, 16'd25757, 16'd19304, 16'd3772, 16'd4265, 16'd41864, 16'd59743, 16'd32926, 16'd37754, 16'd26302, 16'd11555, 16'd18312, 16'd4578, 16'd33848, 16'd1742, 16'd24305});
	test_expansion(128'hb56ada3114206b819969278cda931682, {16'd14527, 16'd32140, 16'd24806, 16'd19401, 16'd12446, 16'd54092, 16'd25491, 16'd42004, 16'd55499, 16'd47247, 16'd46471, 16'd62179, 16'd45452, 16'd33519, 16'd37236, 16'd22449, 16'd28552, 16'd46751, 16'd1563, 16'd45409, 16'd15018, 16'd30089, 16'd41338, 16'd49530, 16'd53843, 16'd33340});
	test_expansion(128'h19af29e1467de3e289712c149337556f, {16'd62563, 16'd16772, 16'd17847, 16'd59872, 16'd36605, 16'd32246, 16'd23429, 16'd57504, 16'd31197, 16'd44516, 16'd1755, 16'd13386, 16'd12355, 16'd5882, 16'd4005, 16'd39321, 16'd50560, 16'd22122, 16'd31053, 16'd56204, 16'd12603, 16'd46681, 16'd29636, 16'd61851, 16'd52254, 16'd35383});
	test_expansion(128'hfdd240e24e0bd801195d6730041147d7, {16'd52514, 16'd29679, 16'd32818, 16'd46000, 16'd6450, 16'd47426, 16'd16779, 16'd19022, 16'd37662, 16'd23434, 16'd26642, 16'd7609, 16'd22072, 16'd6387, 16'd49146, 16'd43934, 16'd33624, 16'd5554, 16'd10956, 16'd14172, 16'd10471, 16'd2371, 16'd23958, 16'd36017, 16'd52000, 16'd48729});
	test_expansion(128'he409bf9578f7dd98b02ff0784e37ea7c, {16'd7758, 16'd15892, 16'd20371, 16'd10000, 16'd43241, 16'd60031, 16'd14341, 16'd53397, 16'd23410, 16'd46303, 16'd63811, 16'd32513, 16'd53583, 16'd6761, 16'd18125, 16'd33352, 16'd59014, 16'd25584, 16'd33025, 16'd62666, 16'd20599, 16'd7306, 16'd6677, 16'd51079, 16'd50444, 16'd52290});
	test_expansion(128'hf6bb75afb96e5f6807696a7deeadd6a1, {16'd37961, 16'd50220, 16'd64915, 16'd22536, 16'd7972, 16'd24059, 16'd65375, 16'd60718, 16'd17662, 16'd6690, 16'd39873, 16'd22881, 16'd64205, 16'd32841, 16'd56197, 16'd22440, 16'd40028, 16'd53975, 16'd42260, 16'd36558, 16'd56948, 16'd25341, 16'd36505, 16'd40538, 16'd17590, 16'd59798});
	test_expansion(128'h8f16e949c749a9b89e7f8b2391b865dd, {16'd32587, 16'd27710, 16'd64336, 16'd54353, 16'd65009, 16'd42836, 16'd8897, 16'd40953, 16'd30962, 16'd58899, 16'd11448, 16'd43656, 16'd30564, 16'd15285, 16'd47115, 16'd20143, 16'd13840, 16'd14091, 16'd61008, 16'd60083, 16'd60851, 16'd11755, 16'd36276, 16'd65507, 16'd49786, 16'd9928});
	test_expansion(128'he1d0e468fab1bd1240149d81ff429d37, {16'd59293, 16'd11999, 16'd14181, 16'd8330, 16'd60244, 16'd3466, 16'd6421, 16'd54258, 16'd1607, 16'd62251, 16'd57450, 16'd45377, 16'd18362, 16'd38854, 16'd58298, 16'd41402, 16'd56436, 16'd32184, 16'd63085, 16'd6783, 16'd37389, 16'd47209, 16'd37418, 16'd49667, 16'd46500, 16'd55715});
	test_expansion(128'h39f5c2427a2fb30fca6d7dbe72734f13, {16'd28797, 16'd21109, 16'd9710, 16'd46375, 16'd50485, 16'd46361, 16'd26342, 16'd41456, 16'd4768, 16'd17658, 16'd25880, 16'd18736, 16'd22635, 16'd13340, 16'd11620, 16'd5184, 16'd47414, 16'd48933, 16'd8141, 16'd61170, 16'd24866, 16'd23696, 16'd19751, 16'd841, 16'd63988, 16'd20250});
	test_expansion(128'h129d4de8c12d56641fd38dbc5860ec0a, {16'd63371, 16'd3828, 16'd379, 16'd8573, 16'd17655, 16'd45991, 16'd9889, 16'd12808, 16'd35513, 16'd40705, 16'd41751, 16'd9927, 16'd18714, 16'd17105, 16'd58171, 16'd32120, 16'd21513, 16'd59279, 16'd13984, 16'd20330, 16'd9959, 16'd13370, 16'd7003, 16'd36410, 16'd14057, 16'd7713});
	test_expansion(128'hbc5a833f561e814fe64d3f2df4ae05f5, {16'd11201, 16'd36509, 16'd3659, 16'd25386, 16'd17455, 16'd31285, 16'd21115, 16'd25218, 16'd5939, 16'd16657, 16'd46410, 16'd49349, 16'd44436, 16'd6862, 16'd4, 16'd7010, 16'd62265, 16'd21991, 16'd30276, 16'd52378, 16'd19815, 16'd19596, 16'd18503, 16'd329, 16'd60438, 16'd21720});
	test_expansion(128'h2ba01222b101d717f3bce8cfdd59c1c9, {16'd13083, 16'd20013, 16'd33470, 16'd55007, 16'd12152, 16'd13666, 16'd39075, 16'd32854, 16'd63678, 16'd2027, 16'd52012, 16'd31160, 16'd25457, 16'd8124, 16'd19396, 16'd20054, 16'd12914, 16'd30249, 16'd59304, 16'd8873, 16'd26268, 16'd35324, 16'd40041, 16'd19876, 16'd56103, 16'd18845});
	test_expansion(128'h6ef69b3c77f947cde16dc5ecd7841098, {16'd54743, 16'd52682, 16'd39298, 16'd35207, 16'd63578, 16'd6028, 16'd2164, 16'd64927, 16'd10114, 16'd30233, 16'd40959, 16'd48252, 16'd3952, 16'd17851, 16'd42187, 16'd341, 16'd46800, 16'd24321, 16'd52073, 16'd44257, 16'd59586, 16'd44702, 16'd17719, 16'd50148, 16'd8325, 16'd20162});
	test_expansion(128'hf085883f8858d2fa0baa4c78f6207598, {16'd21084, 16'd35281, 16'd7383, 16'd13292, 16'd22219, 16'd6337, 16'd8672, 16'd11458, 16'd65378, 16'd672, 16'd12085, 16'd6846, 16'd37184, 16'd33599, 16'd14937, 16'd27488, 16'd60662, 16'd27271, 16'd19086, 16'd62083, 16'd29097, 16'd26348, 16'd48987, 16'd21014, 16'd34106, 16'd49669});
	test_expansion(128'h0966a22a25aede2c03309878093e258e, {16'd8932, 16'd57798, 16'd26195, 16'd39339, 16'd19905, 16'd5691, 16'd42640, 16'd25950, 16'd18876, 16'd765, 16'd26394, 16'd29132, 16'd61403, 16'd38648, 16'd36417, 16'd5193, 16'd34594, 16'd8784, 16'd32864, 16'd42646, 16'd7230, 16'd59317, 16'd14861, 16'd53402, 16'd15703, 16'd52509});
	test_expansion(128'hddc7132135f0d289c7e7c38da853f243, {16'd48022, 16'd3605, 16'd4195, 16'd62545, 16'd53150, 16'd19345, 16'd52730, 16'd27236, 16'd39440, 16'd33939, 16'd24219, 16'd60402, 16'd30719, 16'd8832, 16'd51258, 16'd25336, 16'd26622, 16'd8173, 16'd61571, 16'd38003, 16'd2045, 16'd27285, 16'd59973, 16'd37543, 16'd43588, 16'd49760});
	test_expansion(128'hb8b02d3ab898c4defa27087ff2c15488, {16'd42721, 16'd64320, 16'd33825, 16'd48475, 16'd35125, 16'd61212, 16'd12027, 16'd54139, 16'd17847, 16'd14455, 16'd52684, 16'd46285, 16'd9076, 16'd8102, 16'd48972, 16'd27832, 16'd33958, 16'd3346, 16'd2971, 16'd23922, 16'd43895, 16'd15111, 16'd33420, 16'd23318, 16'd47877, 16'd14850});
	test_expansion(128'h0074a336560071b62626c702770130b3, {16'd45754, 16'd23985, 16'd59219, 16'd33005, 16'd11237, 16'd8360, 16'd39207, 16'd49396, 16'd23534, 16'd17401, 16'd48054, 16'd24916, 16'd11359, 16'd2659, 16'd4962, 16'd50405, 16'd35104, 16'd62849, 16'd63636, 16'd24128, 16'd40671, 16'd9165, 16'd41712, 16'd34332, 16'd61088, 16'd15449});
	test_expansion(128'hab76598b080796d4c3c947fc574d59a9, {16'd29086, 16'd37005, 16'd53034, 16'd11313, 16'd13599, 16'd60197, 16'd12462, 16'd311, 16'd12578, 16'd46408, 16'd17017, 16'd47803, 16'd8923, 16'd29596, 16'd33434, 16'd24317, 16'd29036, 16'd64562, 16'd22276, 16'd19840, 16'd18328, 16'd26489, 16'd25826, 16'd56292, 16'd55766, 16'd38739});
	test_expansion(128'h758dbcf4d5f6c0bb39a3cbf236425f66, {16'd11818, 16'd6107, 16'd40701, 16'd42775, 16'd34370, 16'd50326, 16'd9851, 16'd34634, 16'd20767, 16'd604, 16'd38158, 16'd29554, 16'd23376, 16'd34995, 16'd12511, 16'd57390, 16'd30346, 16'd39113, 16'd8317, 16'd53422, 16'd55799, 16'd40641, 16'd10724, 16'd40672, 16'd46224, 16'd8059});
	test_expansion(128'h775b048d626deabde1164aba5c68cd0d, {16'd59558, 16'd42054, 16'd57549, 16'd1782, 16'd4556, 16'd30844, 16'd38178, 16'd58642, 16'd59176, 16'd4507, 16'd37534, 16'd26565, 16'd10576, 16'd46491, 16'd38200, 16'd37878, 16'd48691, 16'd55939, 16'd57290, 16'd46224, 16'd36996, 16'd23350, 16'd57935, 16'd13854, 16'd33322, 16'd42359});
	test_expansion(128'h9dc96e140979324a46336b5d9fcc8d50, {16'd17710, 16'd39171, 16'd17176, 16'd21959, 16'd50468, 16'd47365, 16'd9786, 16'd3997, 16'd29531, 16'd56516, 16'd4291, 16'd54759, 16'd35339, 16'd17879, 16'd42319, 16'd43000, 16'd5226, 16'd43265, 16'd35670, 16'd64174, 16'd55400, 16'd48985, 16'd44712, 16'd28622, 16'd51422, 16'd8263});
	test_expansion(128'h65a42d4f6b8a2fe656daf9edb82fe29e, {16'd42189, 16'd44321, 16'd18047, 16'd14374, 16'd38523, 16'd2281, 16'd24785, 16'd57447, 16'd5748, 16'd40336, 16'd28835, 16'd15276, 16'd33055, 16'd46023, 16'd40713, 16'd5096, 16'd17063, 16'd63684, 16'd8355, 16'd60872, 16'd59793, 16'd12867, 16'd46729, 16'd24992, 16'd11382, 16'd54849});
	test_expansion(128'hfc67e8076a21e2b4bee18cbab687fdcb, {16'd46119, 16'd53052, 16'd1584, 16'd26598, 16'd24891, 16'd19760, 16'd30908, 16'd36589, 16'd26198, 16'd14206, 16'd32689, 16'd33131, 16'd55651, 16'd61977, 16'd17781, 16'd29293, 16'd63361, 16'd23043, 16'd43440, 16'd58744, 16'd4252, 16'd46067, 16'd37705, 16'd16160, 16'd12506, 16'd1940});
	test_expansion(128'hd03ac4bd08f555be2cc8a0f6caf144ae, {16'd37293, 16'd33257, 16'd13819, 16'd7280, 16'd30363, 16'd14094, 16'd35216, 16'd25787, 16'd40701, 16'd15487, 16'd13806, 16'd5850, 16'd65321, 16'd35005, 16'd41800, 16'd30917, 16'd61386, 16'd6859, 16'd59058, 16'd20421, 16'd319, 16'd52216, 16'd60149, 16'd62195, 16'd54560, 16'd31864});
	test_expansion(128'hb1f050f541aeb72fa9c5060f5cdfb328, {16'd19105, 16'd31077, 16'd47598, 16'd28666, 16'd60804, 16'd31326, 16'd34324, 16'd3141, 16'd34094, 16'd39128, 16'd46732, 16'd64031, 16'd61076, 16'd39130, 16'd46789, 16'd15946, 16'd6728, 16'd34650, 16'd52296, 16'd45384, 16'd63423, 16'd48312, 16'd48646, 16'd55883, 16'd45366, 16'd21078});
	test_expansion(128'ha45adf967b48083a642b860b978adff8, {16'd50220, 16'd16130, 16'd36192, 16'd2313, 16'd22522, 16'd35766, 16'd54475, 16'd17595, 16'd34, 16'd7869, 16'd15672, 16'd32763, 16'd38758, 16'd60362, 16'd59880, 16'd60303, 16'd63114, 16'd39554, 16'd46668, 16'd45596, 16'd35275, 16'd1102, 16'd13528, 16'd24779, 16'd50521, 16'd44171});
	test_expansion(128'h45325f48c43e0f3d04d29aadde024c96, {16'd53544, 16'd23513, 16'd56822, 16'd30144, 16'd23945, 16'd33143, 16'd6958, 16'd53484, 16'd33037, 16'd33980, 16'd25910, 16'd43668, 16'd53328, 16'd62560, 16'd2496, 16'd2901, 16'd11146, 16'd2076, 16'd63319, 16'd14255, 16'd14201, 16'd63355, 16'd41814, 16'd35998, 16'd21264, 16'd56323});
	test_expansion(128'h758d92ee5b0d9ff9352d7945cba0c3b7, {16'd1402, 16'd3784, 16'd8212, 16'd63541, 16'd51198, 16'd53449, 16'd39271, 16'd37974, 16'd49065, 16'd60348, 16'd35372, 16'd21846, 16'd887, 16'd13337, 16'd27038, 16'd64722, 16'd32385, 16'd5531, 16'd49522, 16'd54282, 16'd7292, 16'd6263, 16'd35852, 16'd49856, 16'd60822, 16'd48057});
	test_expansion(128'habdc5d79ae30e5cdc714c690f55e086f, {16'd24118, 16'd14000, 16'd44868, 16'd38710, 16'd186, 16'd8523, 16'd52404, 16'd49646, 16'd62263, 16'd7540, 16'd44060, 16'd6861, 16'd28354, 16'd6205, 16'd63335, 16'd25039, 16'd12282, 16'd10597, 16'd8503, 16'd8763, 16'd35998, 16'd40785, 16'd25698, 16'd22679, 16'd9755, 16'd61402});
	test_expansion(128'h0a83dc25d8f19570121d4d521c620bf6, {16'd37937, 16'd46625, 16'd28259, 16'd13166, 16'd18006, 16'd30252, 16'd51954, 16'd20083, 16'd29084, 16'd37088, 16'd52403, 16'd2844, 16'd8967, 16'd24174, 16'd21972, 16'd53196, 16'd62388, 16'd32222, 16'd21907, 16'd23457, 16'd64893, 16'd59273, 16'd3106, 16'd5653, 16'd58706, 16'd9718});
	test_expansion(128'h0114a9a0e9c6686e7dc64cb9a575264e, {16'd55212, 16'd22331, 16'd62047, 16'd24634, 16'd32574, 16'd50256, 16'd64422, 16'd30579, 16'd18623, 16'd48831, 16'd46151, 16'd33654, 16'd361, 16'd22021, 16'd57685, 16'd46750, 16'd14814, 16'd23001, 16'd49186, 16'd46343, 16'd39213, 16'd53421, 16'd9754, 16'd2741, 16'd57526, 16'd23985});
	test_expansion(128'hfe90a4db69208c74f80744dddf976dcb, {16'd46617, 16'd46951, 16'd11808, 16'd11052, 16'd47294, 16'd2726, 16'd52253, 16'd51340, 16'd56797, 16'd58687, 16'd11741, 16'd33942, 16'd54470, 16'd29989, 16'd6053, 16'd65415, 16'd65439, 16'd40257, 16'd53481, 16'd45684, 16'd46071, 16'd28821, 16'd58061, 16'd56496, 16'd42993, 16'd49110});
	test_expansion(128'h0b3339031c7e49ff36b55388299a16aa, {16'd800, 16'd62223, 16'd8924, 16'd41225, 16'd2321, 16'd23343, 16'd57985, 16'd1178, 16'd27997, 16'd49514, 16'd173, 16'd48351, 16'd23519, 16'd40685, 16'd12567, 16'd38210, 16'd28787, 16'd13648, 16'd36616, 16'd61159, 16'd10817, 16'd14929, 16'd3185, 16'd12417, 16'd54498, 16'd55614});
	test_expansion(128'hdedec62402a9e372da7c36dc5d733e9e, {16'd56510, 16'd21703, 16'd20968, 16'd16949, 16'd48820, 16'd18755, 16'd9769, 16'd6988, 16'd15108, 16'd48487, 16'd63490, 16'd48777, 16'd10137, 16'd17282, 16'd16874, 16'd17493, 16'd4560, 16'd31624, 16'd49328, 16'd12024, 16'd2054, 16'd55967, 16'd60553, 16'd59276, 16'd44665, 16'd64069});
	test_expansion(128'h895417073374216fc57f766b2c962b6e, {16'd55291, 16'd6357, 16'd25994, 16'd42547, 16'd48490, 16'd81, 16'd4038, 16'd31360, 16'd10114, 16'd17601, 16'd64192, 16'd58582, 16'd59470, 16'd49122, 16'd37642, 16'd29733, 16'd54174, 16'd38785, 16'd54869, 16'd38117, 16'd65439, 16'd52577, 16'd28107, 16'd13351, 16'd46964, 16'd36833});
	test_expansion(128'hc3e1bf3c219a6f422130f2a3785a0ed6, {16'd9686, 16'd2206, 16'd52233, 16'd51197, 16'd42666, 16'd718, 16'd34932, 16'd19599, 16'd30386, 16'd48118, 16'd16185, 16'd61397, 16'd1841, 16'd4466, 16'd41564, 16'd19672, 16'd58986, 16'd41395, 16'd17027, 16'd13508, 16'd47899, 16'd42810, 16'd1387, 16'd51770, 16'd15004, 16'd38659});
	test_expansion(128'hd3982b8b434cc386d6dfe4af94da7be8, {16'd6205, 16'd684, 16'd4237, 16'd39269, 16'd26105, 16'd6608, 16'd1669, 16'd21485, 16'd25279, 16'd41155, 16'd35087, 16'd1431, 16'd63719, 16'd1456, 16'd55544, 16'd14723, 16'd39046, 16'd280, 16'd45931, 16'd14312, 16'd46909, 16'd29988, 16'd59082, 16'd20587, 16'd41064, 16'd2586});
	test_expansion(128'h689c40f66941f0a9fe18c8333c0ff08a, {16'd8056, 16'd54869, 16'd61462, 16'd44668, 16'd2535, 16'd60696, 16'd24050, 16'd4535, 16'd33729, 16'd25835, 16'd48997, 16'd37875, 16'd26598, 16'd33133, 16'd20362, 16'd27221, 16'd20950, 16'd57796, 16'd32582, 16'd54507, 16'd24283, 16'd1809, 16'd37, 16'd51017, 16'd16228, 16'd30309});
	test_expansion(128'haa8b71011b0c39d6f36a01d748744f4f, {16'd3220, 16'd63115, 16'd2705, 16'd29962, 16'd30247, 16'd28876, 16'd29472, 16'd60435, 16'd32820, 16'd18219, 16'd40011, 16'd41420, 16'd32059, 16'd55188, 16'd18819, 16'd62938, 16'd47706, 16'd26812, 16'd57818, 16'd4652, 16'd24884, 16'd29693, 16'd9322, 16'd47052, 16'd51309, 16'd6148});
	test_expansion(128'h44dac21dc5720feec447397418038485, {16'd63653, 16'd36389, 16'd37524, 16'd45602, 16'd5640, 16'd40067, 16'd54492, 16'd50540, 16'd57967, 16'd52124, 16'd48346, 16'd26456, 16'd49719, 16'd59251, 16'd11997, 16'd19233, 16'd35109, 16'd36802, 16'd20321, 16'd57204, 16'd56467, 16'd28736, 16'd54293, 16'd59122, 16'd2673, 16'd7816});
	test_expansion(128'h51f4f69cbe2d13f163ad8bc1c1a089a6, {16'd55057, 16'd61962, 16'd23038, 16'd40209, 16'd11415, 16'd56167, 16'd59987, 16'd17407, 16'd48908, 16'd39643, 16'd32312, 16'd35740, 16'd930, 16'd60087, 16'd58258, 16'd19287, 16'd16881, 16'd44151, 16'd4006, 16'd10085, 16'd9768, 16'd52232, 16'd38206, 16'd12300, 16'd54305, 16'd52050});
	test_expansion(128'hdc8606b30793f5b88367ccd4197dc1b6, {16'd33713, 16'd17753, 16'd18574, 16'd8968, 16'd59364, 16'd36212, 16'd59170, 16'd39496, 16'd21936, 16'd45531, 16'd63753, 16'd62354, 16'd20452, 16'd61712, 16'd19649, 16'd32739, 16'd47855, 16'd19507, 16'd34420, 16'd12894, 16'd14434, 16'd21726, 16'd20666, 16'd53042, 16'd3256, 16'd29779});
	test_expansion(128'hbc05294175417d2e07a05d2650476997, {16'd27326, 16'd31695, 16'd38075, 16'd1399, 16'd30363, 16'd58067, 16'd51280, 16'd8289, 16'd34167, 16'd50711, 16'd31508, 16'd48744, 16'd62369, 16'd53309, 16'd12147, 16'd51162, 16'd49169, 16'd29459, 16'd58840, 16'd1438, 16'd63433, 16'd48028, 16'd63346, 16'd9282, 16'd48913, 16'd60346});
	test_expansion(128'h3f9264feba23fb1ee1a3ae28f8f39c4a, {16'd26295, 16'd23128, 16'd45873, 16'd45740, 16'd24335, 16'd35230, 16'd18790, 16'd55357, 16'd52373, 16'd57956, 16'd56637, 16'd12501, 16'd53466, 16'd15695, 16'd12590, 16'd61561, 16'd13412, 16'd59559, 16'd21285, 16'd55408, 16'd53048, 16'd8015, 16'd64388, 16'd11400, 16'd2703, 16'd51092});
	test_expansion(128'h15eabf553f7781b05ebfcbabdb4f1cd6, {16'd36038, 16'd2521, 16'd36727, 16'd60079, 16'd45652, 16'd10973, 16'd29490, 16'd11189, 16'd36533, 16'd47730, 16'd28143, 16'd8703, 16'd17610, 16'd7030, 16'd56718, 16'd36787, 16'd414, 16'd30804, 16'd4440, 16'd50128, 16'd53587, 16'd37553, 16'd55187, 16'd63212, 16'd49060, 16'd13556});
	test_expansion(128'hec29eef9d2fad42c4390e29093072c24, {16'd42659, 16'd51132, 16'd55924, 16'd18285, 16'd45187, 16'd15943, 16'd11801, 16'd22997, 16'd5904, 16'd4113, 16'd12045, 16'd44942, 16'd48460, 16'd21645, 16'd26645, 16'd11889, 16'd9883, 16'd44513, 16'd4728, 16'd4084, 16'd55092, 16'd4429, 16'd8833, 16'd54918, 16'd44502, 16'd36762});
	test_expansion(128'h5f3c41778b6225198e609970159b81f2, {16'd2929, 16'd8020, 16'd22859, 16'd21711, 16'd47748, 16'd6002, 16'd40235, 16'd42594, 16'd14810, 16'd53732, 16'd351, 16'd24753, 16'd8140, 16'd56716, 16'd61991, 16'd57808, 16'd58179, 16'd31303, 16'd43679, 16'd16472, 16'd38600, 16'd27624, 16'd34168, 16'd17951, 16'd26618, 16'd27387});
	test_expansion(128'h5c2472b2736830f18a513b8b52547554, {16'd58832, 16'd24664, 16'd3090, 16'd60255, 16'd8097, 16'd20354, 16'd28657, 16'd47441, 16'd36370, 16'd55914, 16'd2515, 16'd39759, 16'd3162, 16'd54573, 16'd51198, 16'd20246, 16'd20296, 16'd19433, 16'd40415, 16'd50743, 16'd46340, 16'd6035, 16'd14360, 16'd4602, 16'd57598, 16'd27463});
	test_expansion(128'hbc739f3c4cd5564fd75a2bafa986a844, {16'd11497, 16'd13368, 16'd46730, 16'd50110, 16'd5727, 16'd38939, 16'd53127, 16'd14368, 16'd39802, 16'd31669, 16'd19303, 16'd58614, 16'd1942, 16'd20645, 16'd53370, 16'd905, 16'd22140, 16'd22977, 16'd58776, 16'd14601, 16'd30765, 16'd9228, 16'd57124, 16'd14986, 16'd57544, 16'd39125});
	test_expansion(128'h3469b1ecace4a362a43bb8fcd5bc0e17, {16'd49654, 16'd37989, 16'd26745, 16'd21474, 16'd2665, 16'd33585, 16'd14812, 16'd1343, 16'd62832, 16'd29919, 16'd58361, 16'd24071, 16'd2839, 16'd36271, 16'd28800, 16'd32682, 16'd20260, 16'd48625, 16'd43922, 16'd50689, 16'd38352, 16'd50810, 16'd20705, 16'd19882, 16'd3363, 16'd46960});
	test_expansion(128'h2af01593c00d1b89b17ec7749292563c, {16'd28959, 16'd8791, 16'd51077, 16'd33970, 16'd63219, 16'd20957, 16'd63838, 16'd11998, 16'd35019, 16'd30094, 16'd38231, 16'd37250, 16'd65518, 16'd943, 16'd45813, 16'd47616, 16'd32138, 16'd55944, 16'd44875, 16'd19586, 16'd27951, 16'd45994, 16'd2301, 16'd58190, 16'd16562, 16'd5251});
	test_expansion(128'hdd59183a144a9246ece20baf8dd5547a, {16'd45290, 16'd22263, 16'd6545, 16'd49147, 16'd34134, 16'd23459, 16'd48687, 16'd12364, 16'd27595, 16'd49952, 16'd36028, 16'd65165, 16'd28314, 16'd46379, 16'd48828, 16'd32768, 16'd49980, 16'd12310, 16'd54784, 16'd31518, 16'd44789, 16'd8902, 16'd1653, 16'd55518, 16'd19586, 16'd38499});
	test_expansion(128'hb116ac092c5bbaa5cfef36d6633ce3de, {16'd40082, 16'd6474, 16'd31596, 16'd25784, 16'd49008, 16'd37711, 16'd15367, 16'd5574, 16'd3244, 16'd13434, 16'd11905, 16'd32843, 16'd52507, 16'd36325, 16'd63090, 16'd9557, 16'd6576, 16'd41378, 16'd48295, 16'd15848, 16'd57055, 16'd44784, 16'd29361, 16'd10257, 16'd30621, 16'd23086});
	test_expansion(128'hf38ceb942ef566b5dcd07dfc8767e991, {16'd58736, 16'd55551, 16'd40835, 16'd4082, 16'd5027, 16'd5572, 16'd47751, 16'd6255, 16'd51934, 16'd36969, 16'd57694, 16'd4373, 16'd50655, 16'd36664, 16'd53981, 16'd47039, 16'd12595, 16'd49457, 16'd57898, 16'd52151, 16'd36299, 16'd17046, 16'd30861, 16'd57196, 16'd58955, 16'd28813});
	test_expansion(128'h92d57b71f928933cc8d529a17096aa7d, {16'd35795, 16'd54461, 16'd53144, 16'd12308, 16'd42559, 16'd7022, 16'd51253, 16'd9427, 16'd20930, 16'd45138, 16'd20654, 16'd50097, 16'd62731, 16'd29157, 16'd29589, 16'd46878, 16'd55351, 16'd28337, 16'd18126, 16'd49448, 16'd51708, 16'd55253, 16'd30875, 16'd1908, 16'd7666, 16'd12466});
	test_expansion(128'h31f7dbec406656278c76bdcfe9e93333, {16'd23780, 16'd12418, 16'd7465, 16'd30331, 16'd57181, 16'd35297, 16'd6916, 16'd50670, 16'd60582, 16'd24322, 16'd40528, 16'd21840, 16'd49623, 16'd12944, 16'd36524, 16'd45813, 16'd16603, 16'd46485, 16'd64426, 16'd40158, 16'd22743, 16'd37150, 16'd51183, 16'd51903, 16'd64076, 16'd38466});
	test_expansion(128'h95b1356e2e8bab7d2c5be37923c11adf, {16'd55284, 16'd9490, 16'd33011, 16'd3600, 16'd11581, 16'd7321, 16'd6245, 16'd27150, 16'd8641, 16'd28081, 16'd1620, 16'd24544, 16'd29527, 16'd61702, 16'd17157, 16'd51375, 16'd62730, 16'd56850, 16'd58371, 16'd17270, 16'd40089, 16'd65412, 16'd50530, 16'd21210, 16'd35441, 16'd36022});
	test_expansion(128'hd069b01e9a9077cdb90dbf4e9fcbc687, {16'd39574, 16'd6581, 16'd49291, 16'd14793, 16'd16679, 16'd40221, 16'd55856, 16'd65490, 16'd47138, 16'd42821, 16'd63423, 16'd5499, 16'd21744, 16'd13139, 16'd21596, 16'd4816, 16'd61808, 16'd1478, 16'd29390, 16'd56640, 16'd50261, 16'd41599, 16'd15825, 16'd48793, 16'd6330, 16'd18681});
	test_expansion(128'h8e0a4363cd4d8103d9959a5be9f6748f, {16'd29449, 16'd16860, 16'd58564, 16'd13634, 16'd13073, 16'd63323, 16'd59806, 16'd895, 16'd5733, 16'd55416, 16'd41570, 16'd49433, 16'd39288, 16'd63606, 16'd58505, 16'd32394, 16'd50598, 16'd43698, 16'd1623, 16'd11372, 16'd5127, 16'd33618, 16'd19408, 16'd4323, 16'd7904, 16'd9778});
	test_expansion(128'h05789870d130d59cdb301cfa5d5a47bd, {16'd34380, 16'd15619, 16'd57371, 16'd49410, 16'd57699, 16'd42889, 16'd6586, 16'd9987, 16'd63664, 16'd65191, 16'd33374, 16'd26123, 16'd23337, 16'd8532, 16'd45634, 16'd59437, 16'd47748, 16'd59205, 16'd11610, 16'd65330, 16'd10333, 16'd16959, 16'd30640, 16'd24785, 16'd58872, 16'd24306});
	test_expansion(128'h61a84574b6741050c0fc1253a7fd77aa, {16'd5092, 16'd30691, 16'd6522, 16'd39930, 16'd4842, 16'd58210, 16'd55448, 16'd32661, 16'd28634, 16'd18305, 16'd35511, 16'd47484, 16'd22050, 16'd49467, 16'd2905, 16'd22441, 16'd44443, 16'd47138, 16'd47376, 16'd46101, 16'd7171, 16'd55853, 16'd5792, 16'd61311, 16'd41140, 16'd20621});
	test_expansion(128'h6e69c1cf8bfaada36417d5a82c095754, {16'd53761, 16'd44758, 16'd44563, 16'd38271, 16'd20967, 16'd51562, 16'd49375, 16'd2811, 16'd50345, 16'd3513, 16'd39029, 16'd42562, 16'd54100, 16'd20306, 16'd25971, 16'd28614, 16'd50835, 16'd21994, 16'd40130, 16'd37698, 16'd37171, 16'd11943, 16'd7353, 16'd59285, 16'd55330, 16'd44240});
	test_expansion(128'he87154db80050933042d0d39bdda3aef, {16'd25155, 16'd35841, 16'd53872, 16'd50256, 16'd21240, 16'd61799, 16'd15988, 16'd47243, 16'd28565, 16'd23668, 16'd3406, 16'd5371, 16'd36539, 16'd3081, 16'd35022, 16'd11239, 16'd30279, 16'd57982, 16'd28533, 16'd22278, 16'd34172, 16'd51289, 16'd35804, 16'd44423, 16'd23815, 16'd44834});
	test_expansion(128'hbd455254e42d5d3e393eb75320f7ad7e, {16'd11145, 16'd17625, 16'd55432, 16'd21971, 16'd64107, 16'd36055, 16'd3245, 16'd50214, 16'd59804, 16'd46042, 16'd50324, 16'd29923, 16'd57003, 16'd866, 16'd37177, 16'd18717, 16'd13695, 16'd60029, 16'd24316, 16'd1894, 16'd60746, 16'd16211, 16'd58993, 16'd21532, 16'd1579, 16'd40657});
	test_expansion(128'h0e70109c5161c837ed12729dea960b16, {16'd6391, 16'd57215, 16'd41854, 16'd39439, 16'd58636, 16'd1419, 16'd5890, 16'd10279, 16'd12687, 16'd6282, 16'd16670, 16'd10159, 16'd36688, 16'd57294, 16'd34970, 16'd19201, 16'd51857, 16'd8737, 16'd29888, 16'd5072, 16'd45667, 16'd9926, 16'd25506, 16'd57425, 16'd18781, 16'd58200});
	test_expansion(128'hf3ccd87de8bc15aa7e255b42b3828025, {16'd28246, 16'd3773, 16'd3212, 16'd25202, 16'd19055, 16'd16575, 16'd54133, 16'd32012, 16'd2154, 16'd29862, 16'd20890, 16'd5899, 16'd27113, 16'd57900, 16'd12049, 16'd22995, 16'd64852, 16'd33151, 16'd63656, 16'd6283, 16'd24939, 16'd27764, 16'd18335, 16'd8504, 16'd14756, 16'd22464});
	test_expansion(128'h5a15919d23de144126e53174411c872b, {16'd18439, 16'd65255, 16'd51257, 16'd18532, 16'd4576, 16'd52714, 16'd7605, 16'd55014, 16'd55103, 16'd18533, 16'd33850, 16'd22305, 16'd28678, 16'd19871, 16'd28467, 16'd23447, 16'd39197, 16'd28686, 16'd35902, 16'd47428, 16'd12062, 16'd4518, 16'd8010, 16'd46450, 16'd53800, 16'd64741});
	test_expansion(128'hc9673b3c4bb89c970fb1c22f3f6b5a33, {16'd43109, 16'd33378, 16'd20908, 16'd23139, 16'd63711, 16'd12513, 16'd39763, 16'd55740, 16'd57148, 16'd25100, 16'd36029, 16'd63220, 16'd52592, 16'd61716, 16'd21463, 16'd58613, 16'd30825, 16'd10578, 16'd29087, 16'd44058, 16'd63513, 16'd12853, 16'd9656, 16'd52153, 16'd49911, 16'd29172});
	test_expansion(128'hbc2cfc249cfac3472aa71c5610015a7b, {16'd8902, 16'd53700, 16'd21800, 16'd47404, 16'd44357, 16'd21814, 16'd24528, 16'd21549, 16'd25485, 16'd61826, 16'd20581, 16'd32827, 16'd52199, 16'd7046, 16'd64428, 16'd18155, 16'd16640, 16'd61237, 16'd26942, 16'd648, 16'd50290, 16'd34258, 16'd29970, 16'd36293, 16'd10022, 16'd64731});
	test_expansion(128'h16baeca0380c23a54cacee197c0f0c4b, {16'd47111, 16'd19126, 16'd40879, 16'd2196, 16'd53706, 16'd49282, 16'd3669, 16'd45779, 16'd45234, 16'd58419, 16'd11773, 16'd789, 16'd41669, 16'd39116, 16'd64465, 16'd3233, 16'd13542, 16'd32727, 16'd36496, 16'd1827, 16'd44128, 16'd9006, 16'd6823, 16'd7259, 16'd60373, 16'd117});
	test_expansion(128'h71f6c370ac07eec14e4dfe6b012ac254, {16'd36922, 16'd54203, 16'd51400, 16'd4715, 16'd11063, 16'd26778, 16'd9087, 16'd39293, 16'd59203, 16'd30636, 16'd44794, 16'd39315, 16'd62974, 16'd47614, 16'd65442, 16'd9142, 16'd43840, 16'd61186, 16'd47354, 16'd10252, 16'd33234, 16'd45116, 16'd10942, 16'd48913, 16'd51118, 16'd26597});
	test_expansion(128'h19edba651486e096dd951986997132f5, {16'd42130, 16'd28463, 16'd53647, 16'd10109, 16'd7939, 16'd24258, 16'd20496, 16'd29082, 16'd21829, 16'd57279, 16'd37418, 16'd2058, 16'd55556, 16'd5804, 16'd28404, 16'd4772, 16'd58251, 16'd22406, 16'd50013, 16'd20516, 16'd47202, 16'd32403, 16'd58376, 16'd59664, 16'd15502, 16'd6932});
	test_expansion(128'h18970abc76dbe28d38d4608a06f596e5, {16'd33093, 16'd62340, 16'd45365, 16'd54029, 16'd55127, 16'd42400, 16'd34090, 16'd28923, 16'd50775, 16'd54041, 16'd8361, 16'd3143, 16'd20281, 16'd46818, 16'd33137, 16'd3193, 16'd39956, 16'd12774, 16'd23425, 16'd39251, 16'd53931, 16'd50672, 16'd58785, 16'd37524, 16'd31981, 16'd55939});
	test_expansion(128'h35b209b4f623110236441e76b6fa8ae3, {16'd22710, 16'd65179, 16'd25991, 16'd58944, 16'd10806, 16'd4962, 16'd60660, 16'd59864, 16'd4950, 16'd48990, 16'd47590, 16'd33834, 16'd36472, 16'd58626, 16'd55418, 16'd48763, 16'd12341, 16'd2427, 16'd21631, 16'd44336, 16'd43263, 16'd595, 16'd39372, 16'd28224, 16'd64867, 16'd10155});
	test_expansion(128'h72806eb5d37379c1b1964cfd340b3a4d, {16'd49396, 16'd10775, 16'd805, 16'd37310, 16'd6720, 16'd16428, 16'd52982, 16'd29672, 16'd61622, 16'd30344, 16'd48784, 16'd56622, 16'd29090, 16'd12303, 16'd36558, 16'd21328, 16'd25377, 16'd14622, 16'd30413, 16'd9694, 16'd10203, 16'd3605, 16'd38912, 16'd24369, 16'd38557, 16'd49761});
	test_expansion(128'hc4f5bf32fc4d9cde8491aa99d1455041, {16'd29919, 16'd25473, 16'd19715, 16'd9868, 16'd1740, 16'd22276, 16'd8592, 16'd10854, 16'd21985, 16'd22587, 16'd43627, 16'd26985, 16'd41758, 16'd13127, 16'd44986, 16'd37828, 16'd61954, 16'd29871, 16'd361, 16'd28009, 16'd31097, 16'd53927, 16'd45790, 16'd14871, 16'd17758, 16'd48013});
	test_expansion(128'h77b7afc3a726d82e30f31aa1f431dece, {16'd34785, 16'd49984, 16'd18596, 16'd38472, 16'd6955, 16'd41894, 16'd30266, 16'd28756, 16'd48382, 16'd4633, 16'd50921, 16'd35696, 16'd17537, 16'd14026, 16'd8474, 16'd61532, 16'd34159, 16'd7115, 16'd34495, 16'd27442, 16'd62008, 16'd21325, 16'd40669, 16'd64047, 16'd32197, 16'd40876});
	test_expansion(128'h7dd2c96b0a6a25c529578a1379867ff6, {16'd61916, 16'd49970, 16'd21823, 16'd13326, 16'd46215, 16'd12142, 16'd44270, 16'd61125, 16'd29978, 16'd23433, 16'd56656, 16'd3591, 16'd27935, 16'd20117, 16'd19363, 16'd32970, 16'd38487, 16'd42495, 16'd27006, 16'd55224, 16'd17664, 16'd29469, 16'd44868, 16'd19620, 16'd34421, 16'd56350});
	test_expansion(128'h55550918d61ea30fe1f862651180e588, {16'd43792, 16'd30989, 16'd15881, 16'd8683, 16'd31338, 16'd13214, 16'd46349, 16'd63478, 16'd23241, 16'd17866, 16'd912, 16'd33863, 16'd52771, 16'd41658, 16'd17186, 16'd61238, 16'd44751, 16'd50766, 16'd17261, 16'd37711, 16'd24356, 16'd21836, 16'd2734, 16'd29893, 16'd30823, 16'd22133});
	test_expansion(128'h404b8a47f761623c712282fb29208996, {16'd32548, 16'd60785, 16'd61682, 16'd24731, 16'd5736, 16'd52504, 16'd64657, 16'd20329, 16'd39046, 16'd21931, 16'd46792, 16'd62247, 16'd16998, 16'd23921, 16'd45257, 16'd65023, 16'd5051, 16'd8822, 16'd29515, 16'd51350, 16'd65075, 16'd30218, 16'd6092, 16'd9314, 16'd30922, 16'd54484});
	test_expansion(128'h8855c98556f80e3b1e00f3b0b1c20f23, {16'd17965, 16'd43223, 16'd65278, 16'd50459, 16'd34941, 16'd65469, 16'd18847, 16'd46145, 16'd32878, 16'd44266, 16'd52947, 16'd32036, 16'd16424, 16'd19629, 16'd50823, 16'd3324, 16'd21338, 16'd1347, 16'd35875, 16'd12560, 16'd19117, 16'd58392, 16'd57464, 16'd5064, 16'd11627, 16'd36771});
	test_expansion(128'hdcd1cb97e5a4728e0b43de602afe708a, {16'd54793, 16'd1329, 16'd49781, 16'd33511, 16'd60374, 16'd47398, 16'd22854, 16'd43684, 16'd46029, 16'd34947, 16'd57676, 16'd8298, 16'd37761, 16'd54706, 16'd20170, 16'd61965, 16'd23593, 16'd5004, 16'd4374, 16'd8670, 16'd60185, 16'd6435, 16'd29614, 16'd65164, 16'd52518, 16'd44279});
	test_expansion(128'h10847bb58fbc437f8fba6dd9c865b64d, {16'd5025, 16'd51027, 16'd64410, 16'd17203, 16'd20527, 16'd21776, 16'd60652, 16'd64528, 16'd41969, 16'd41659, 16'd4166, 16'd64554, 16'd7609, 16'd30557, 16'd51146, 16'd62082, 16'd2795, 16'd43802, 16'd3329, 16'd22197, 16'd35058, 16'd53200, 16'd36497, 16'd38317, 16'd1286, 16'd1641});
	test_expansion(128'h49cd6c494f03fca110fa9e3e1d91d242, {16'd21180, 16'd56938, 16'd57099, 16'd53122, 16'd11569, 16'd20067, 16'd61195, 16'd51609, 16'd62949, 16'd64172, 16'd39350, 16'd24307, 16'd52837, 16'd34289, 16'd54798, 16'd54158, 16'd661, 16'd26118, 16'd47524, 16'd36044, 16'd60018, 16'd20155, 16'd15909, 16'd12988, 16'd4359, 16'd12905});
	test_expansion(128'h1a734f6eda54c855ec66dfb1fcfb293e, {16'd20296, 16'd31792, 16'd32712, 16'd10253, 16'd7274, 16'd57924, 16'd37253, 16'd14398, 16'd12589, 16'd46658, 16'd49678, 16'd36882, 16'd14079, 16'd20505, 16'd41332, 16'd37187, 16'd59741, 16'd48972, 16'd59144, 16'd43655, 16'd38933, 16'd20374, 16'd45298, 16'd56699, 16'd55567, 16'd24072});
	test_expansion(128'habe5e367e28d9fb4bde9e6f7a7d535aa, {16'd15055, 16'd18623, 16'd23707, 16'd60879, 16'd3725, 16'd5836, 16'd5400, 16'd21424, 16'd55044, 16'd61340, 16'd3665, 16'd34136, 16'd33617, 16'd50811, 16'd59822, 16'd46960, 16'd60301, 16'd22216, 16'd49271, 16'd18730, 16'd35216, 16'd18693, 16'd53306, 16'd50725, 16'd14909, 16'd23939});
	test_expansion(128'hcdff51389aac0af0ed9b91ee26723a20, {16'd59179, 16'd27571, 16'd55363, 16'd17618, 16'd1292, 16'd55314, 16'd63508, 16'd58728, 16'd20487, 16'd49209, 16'd5149, 16'd56315, 16'd12522, 16'd19394, 16'd38820, 16'd24217, 16'd53458, 16'd41614, 16'd1688, 16'd28035, 16'd27249, 16'd50342, 16'd1811, 16'd40251, 16'd40337, 16'd2650});
	test_expansion(128'h3619065de782272ebfa07fdaeee692c5, {16'd207, 16'd17172, 16'd23565, 16'd61832, 16'd31584, 16'd57394, 16'd35251, 16'd64070, 16'd42126, 16'd47272, 16'd52338, 16'd11586, 16'd57860, 16'd47141, 16'd52240, 16'd25816, 16'd18772, 16'd64617, 16'd29442, 16'd5489, 16'd11231, 16'd32211, 16'd18327, 16'd50721, 16'd40205, 16'd32998});
	test_expansion(128'hd46e71d9f18f418742e7b7cd28a803d5, {16'd41619, 16'd35511, 16'd37336, 16'd53045, 16'd25680, 16'd47834, 16'd15512, 16'd18780, 16'd36623, 16'd59425, 16'd62363, 16'd40822, 16'd39572, 16'd21589, 16'd31528, 16'd24183, 16'd58995, 16'd52027, 16'd45072, 16'd22186, 16'd3510, 16'd19918, 16'd62583, 16'd45943, 16'd18194, 16'd3049});
	test_expansion(128'h3c458a28fc2c22b12190ca7a467c0442, {16'd24651, 16'd810, 16'd18998, 16'd370, 16'd20018, 16'd40018, 16'd42922, 16'd37909, 16'd30268, 16'd24986, 16'd36936, 16'd24865, 16'd14153, 16'd5892, 16'd17203, 16'd57558, 16'd7165, 16'd42092, 16'd65454, 16'd27890, 16'd64266, 16'd7053, 16'd33994, 16'd29528, 16'd1788, 16'd55500});
	test_expansion(128'h37a0db8e6a8d4f6b41bb059d05ded95b, {16'd44133, 16'd42788, 16'd65433, 16'd6454, 16'd54364, 16'd27030, 16'd33600, 16'd65237, 16'd2400, 16'd29083, 16'd7495, 16'd34376, 16'd42907, 16'd6206, 16'd5330, 16'd7053, 16'd32640, 16'd31314, 16'd27986, 16'd55193, 16'd39154, 16'd10429, 16'd20153, 16'd9612, 16'd21812, 16'd41402});
	test_expansion(128'hf91fde3de2ef46e62bae7a946300daa6, {16'd26375, 16'd30639, 16'd62438, 16'd38537, 16'd1994, 16'd62454, 16'd19663, 16'd61577, 16'd17666, 16'd29934, 16'd9214, 16'd2144, 16'd63227, 16'd56419, 16'd50400, 16'd64114, 16'd52308, 16'd29665, 16'd23710, 16'd57914, 16'd36317, 16'd36909, 16'd24236, 16'd19148, 16'd41494, 16'd54424});
	test_expansion(128'hc2e5b3b73ef8ecf49e431c7efabb4a3e, {16'd3154, 16'd37493, 16'd48160, 16'd54479, 16'd36938, 16'd5681, 16'd61623, 16'd1293, 16'd58943, 16'd3394, 16'd43520, 16'd15920, 16'd51990, 16'd33170, 16'd4250, 16'd42428, 16'd33387, 16'd38734, 16'd7125, 16'd52666, 16'd29927, 16'd51816, 16'd32333, 16'd27437, 16'd28391, 16'd31423});
	test_expansion(128'h541c019a2533a21ba3c6e4f927993ff8, {16'd58262, 16'd29831, 16'd30666, 16'd22082, 16'd18069, 16'd64806, 16'd41529, 16'd21817, 16'd42866, 16'd50357, 16'd30973, 16'd39791, 16'd37960, 16'd36, 16'd19978, 16'd5672, 16'd41637, 16'd54563, 16'd48823, 16'd26273, 16'd19295, 16'd48658, 16'd46414, 16'd14009, 16'd44823, 16'd12945});
	test_expansion(128'h5344088d14489748f1891a49dce45f81, {16'd54457, 16'd52800, 16'd11949, 16'd26860, 16'd45149, 16'd38462, 16'd1033, 16'd23669, 16'd42687, 16'd37664, 16'd37198, 16'd28487, 16'd27028, 16'd45177, 16'd3555, 16'd47647, 16'd63907, 16'd2190, 16'd3394, 16'd27255, 16'd58601, 16'd21726, 16'd14637, 16'd19488, 16'd7863, 16'd13733});
	test_expansion(128'h4bdb9564f0d7b651ae57f67964d394fa, {16'd7302, 16'd20111, 16'd60339, 16'd4576, 16'd5297, 16'd8892, 16'd65492, 16'd26486, 16'd28723, 16'd8209, 16'd63393, 16'd23809, 16'd29287, 16'd17134, 16'd15309, 16'd54218, 16'd27163, 16'd23550, 16'd15265, 16'd56112, 16'd29460, 16'd21314, 16'd32927, 16'd56831, 16'd60338, 16'd3727});
	test_expansion(128'ha9a656acbe06611da37481c358fba00c, {16'd35307, 16'd2555, 16'd16314, 16'd64586, 16'd4357, 16'd16361, 16'd33063, 16'd28958, 16'd3600, 16'd9310, 16'd45342, 16'd56391, 16'd19565, 16'd54071, 16'd6840, 16'd32501, 16'd41552, 16'd13111, 16'd18886, 16'd59640, 16'd49903, 16'd13532, 16'd1173, 16'd46678, 16'd50512, 16'd3412});
	test_expansion(128'he0792b3f4cd4647ba574ee1b4713c241, {16'd18639, 16'd8177, 16'd28842, 16'd483, 16'd10702, 16'd25021, 16'd42236, 16'd18078, 16'd4988, 16'd8689, 16'd25226, 16'd5186, 16'd5744, 16'd48326, 16'd24527, 16'd2628, 16'd25121, 16'd924, 16'd35548, 16'd4969, 16'd6678, 16'd115, 16'd3864, 16'd54661, 16'd18776, 16'd12165});
	test_expansion(128'h98b9a9144ea65f126375667d81a17836, {16'd1674, 16'd31091, 16'd14004, 16'd27432, 16'd3549, 16'd14440, 16'd29268, 16'd39982, 16'd53420, 16'd14043, 16'd10678, 16'd24789, 16'd53417, 16'd7069, 16'd28990, 16'd38053, 16'd25115, 16'd55856, 16'd17816, 16'd35817, 16'd2596, 16'd60617, 16'd36580, 16'd65454, 16'd29659, 16'd57483});
	test_expansion(128'h2aa3d6b1200d38fd9f5afff0044a4a43, {16'd4594, 16'd13017, 16'd5926, 16'd47938, 16'd19711, 16'd37805, 16'd42866, 16'd31998, 16'd51276, 16'd33134, 16'd55605, 16'd49855, 16'd56430, 16'd36982, 16'd20379, 16'd37321, 16'd61567, 16'd21813, 16'd42145, 16'd60059, 16'd33717, 16'd22510, 16'd41594, 16'd29648, 16'd59415, 16'd54462});
	test_expansion(128'h8d5d6ef10939d178511ba110b58b2de8, {16'd44597, 16'd36366, 16'd37365, 16'd24188, 16'd41329, 16'd48383, 16'd57258, 16'd6204, 16'd63909, 16'd45264, 16'd57263, 16'd20540, 16'd44463, 16'd22749, 16'd11554, 16'd37871, 16'd31416, 16'd26419, 16'd897, 16'd9203, 16'd2695, 16'd49363, 16'd19515, 16'd33456, 16'd2584, 16'd22327});
	test_expansion(128'h07820cbfc72d28ad8f0d068807dff66c, {16'd44458, 16'd19311, 16'd64900, 16'd39152, 16'd60010, 16'd18601, 16'd27909, 16'd3974, 16'd34193, 16'd11654, 16'd33567, 16'd6211, 16'd12073, 16'd51155, 16'd33057, 16'd7642, 16'd11615, 16'd20395, 16'd7594, 16'd53865, 16'd23083, 16'd60226, 16'd31756, 16'd40455, 16'd13650, 16'd1557});
	test_expansion(128'h1022d3e40981feadc9c6db59d69adae1, {16'd60743, 16'd50315, 16'd24959, 16'd17216, 16'd63890, 16'd46877, 16'd54402, 16'd18335, 16'd38189, 16'd80, 16'd48428, 16'd25140, 16'd61636, 16'd49218, 16'd37168, 16'd10269, 16'd16007, 16'd26058, 16'd492, 16'd2099, 16'd44968, 16'd15829, 16'd22419, 16'd43653, 16'd65171, 16'd41150});
	test_expansion(128'h3e7322353e5935e15b9e83fd811c5328, {16'd44292, 16'd37499, 16'd23065, 16'd61768, 16'd10272, 16'd22597, 16'd10356, 16'd59380, 16'd55040, 16'd16529, 16'd49420, 16'd29110, 16'd872, 16'd55409, 16'd50221, 16'd1601, 16'd39020, 16'd50862, 16'd5576, 16'd684, 16'd13068, 16'd41042, 16'd15025, 16'd12897, 16'd1273, 16'd18364});
	test_expansion(128'h902125a84c3475b7056e832a52497d6a, {16'd54715, 16'd40215, 16'd5655, 16'd42622, 16'd51630, 16'd24237, 16'd60209, 16'd208, 16'd5717, 16'd34492, 16'd53876, 16'd822, 16'd52992, 16'd52918, 16'd46080, 16'd17627, 16'd26015, 16'd12225, 16'd44504, 16'd29400, 16'd8141, 16'd48557, 16'd44736, 16'd24753, 16'd12762, 16'd40788});
	test_expansion(128'h07307dbb895c5899f85a3711703b55b4, {16'd15721, 16'd26939, 16'd48387, 16'd15009, 16'd44095, 16'd2424, 16'd54527, 16'd46277, 16'd4886, 16'd32087, 16'd62234, 16'd47761, 16'd25029, 16'd62164, 16'd61128, 16'd18181, 16'd19916, 16'd51923, 16'd11243, 16'd24854, 16'd7127, 16'd39551, 16'd52680, 16'd1151, 16'd14437, 16'd48861});
	test_expansion(128'h6cb7abe60855be21bfa025dffea8463f, {16'd12180, 16'd2151, 16'd44557, 16'd50797, 16'd50832, 16'd33292, 16'd41151, 16'd31947, 16'd8184, 16'd5648, 16'd26240, 16'd470, 16'd8116, 16'd30112, 16'd48709, 16'd47046, 16'd45230, 16'd59665, 16'd54006, 16'd51323, 16'd30048, 16'd23628, 16'd8929, 16'd57537, 16'd24407, 16'd26305});
	test_expansion(128'hdd2c967e0d9b931c580652eb296e7f94, {16'd59963, 16'd42574, 16'd30509, 16'd42574, 16'd50424, 16'd3050, 16'd37577, 16'd42460, 16'd50005, 16'd47516, 16'd22824, 16'd65238, 16'd18857, 16'd9472, 16'd27689, 16'd58167, 16'd64287, 16'd34265, 16'd21243, 16'd55772, 16'd35029, 16'd54300, 16'd29305, 16'd25219, 16'd61034, 16'd12266});
	test_expansion(128'h549c6b5db83ccffc6fd54b9db5fea62b, {16'd21773, 16'd43259, 16'd23022, 16'd52299, 16'd27337, 16'd26085, 16'd2186, 16'd38038, 16'd7224, 16'd62072, 16'd19855, 16'd41271, 16'd60825, 16'd55266, 16'd42211, 16'd33396, 16'd17380, 16'd25398, 16'd36303, 16'd15564, 16'd18111, 16'd4034, 16'd60086, 16'd10266, 16'd13907, 16'd18504});
	test_expansion(128'h3264523cc8d816335ecc855c3d9f6a77, {16'd28070, 16'd29703, 16'd5555, 16'd58147, 16'd30247, 16'd37668, 16'd29043, 16'd50830, 16'd13304, 16'd58811, 16'd37026, 16'd24424, 16'd53395, 16'd3933, 16'd45111, 16'd8119, 16'd19659, 16'd41764, 16'd13005, 16'd44965, 16'd14028, 16'd35169, 16'd37908, 16'd1309, 16'd16346, 16'd46127});
	test_expansion(128'hf2c7b957d17a2dc5f277473712753333, {16'd8631, 16'd45884, 16'd5082, 16'd16682, 16'd24353, 16'd33555, 16'd53394, 16'd61542, 16'd62773, 16'd38427, 16'd17243, 16'd6321, 16'd59151, 16'd19593, 16'd19003, 16'd28959, 16'd25061, 16'd19812, 16'd52550, 16'd52689, 16'd19200, 16'd56983, 16'd57352, 16'd63830, 16'd18562, 16'd33390});
	test_expansion(128'h44f01fdb3efc46e2d3da303af162f0cc, {16'd36049, 16'd37489, 16'd51069, 16'd50605, 16'd22180, 16'd45709, 16'd10162, 16'd20843, 16'd24012, 16'd41740, 16'd37066, 16'd52726, 16'd19529, 16'd35861, 16'd54967, 16'd48833, 16'd10999, 16'd51065, 16'd62768, 16'd8893, 16'd19315, 16'd54606, 16'd37891, 16'd31458, 16'd1339, 16'd61534});
	test_expansion(128'h90da7b51b10e0b7cb6b09b0e91122625, {16'd8314, 16'd25833, 16'd57452, 16'd49438, 16'd3662, 16'd37776, 16'd57914, 16'd58586, 16'd27892, 16'd60656, 16'd20875, 16'd22158, 16'd16484, 16'd47330, 16'd48841, 16'd38590, 16'd38462, 16'd53716, 16'd20529, 16'd40201, 16'd23389, 16'd64452, 16'd44900, 16'd51659, 16'd62011, 16'd1531});
	test_expansion(128'hde630d042c50483ea1df0e2001ca58ac, {16'd61375, 16'd25989, 16'd57690, 16'd59489, 16'd8114, 16'd9830, 16'd575, 16'd9396, 16'd19133, 16'd53732, 16'd35629, 16'd17523, 16'd1631, 16'd30472, 16'd43208, 16'd63312, 16'd41745, 16'd10204, 16'd53362, 16'd56982, 16'd51118, 16'd6460, 16'd36021, 16'd36377, 16'd12590, 16'd33849});
	test_expansion(128'h9a3c7e1b0e93364a541628af97b475d5, {16'd29365, 16'd47594, 16'd34244, 16'd63061, 16'd23449, 16'd3652, 16'd51093, 16'd39074, 16'd3329, 16'd45079, 16'd40797, 16'd5648, 16'd52200, 16'd40592, 16'd48672, 16'd37965, 16'd41611, 16'd64678, 16'd5409, 16'd35380, 16'd45884, 16'd62282, 16'd17039, 16'd8315, 16'd27, 16'd6061});
	test_expansion(128'ha5f4290cfde959099dbb70d4a5b23179, {16'd30376, 16'd30843, 16'd63438, 16'd40226, 16'd49419, 16'd58794, 16'd26910, 16'd4093, 16'd26210, 16'd58516, 16'd25785, 16'd50516, 16'd61323, 16'd14951, 16'd6026, 16'd38001, 16'd65364, 16'd29662, 16'd8079, 16'd27167, 16'd53518, 16'd62665, 16'd25789, 16'd19572, 16'd49834, 16'd51205});
	test_expansion(128'h27fb833dd185c8d20e1d280fce95f2a2, {16'd9046, 16'd58968, 16'd21536, 16'd54307, 16'd7742, 16'd15282, 16'd18407, 16'd32655, 16'd49767, 16'd49961, 16'd13390, 16'd8885, 16'd24291, 16'd30848, 16'd2243, 16'd56787, 16'd61241, 16'd57942, 16'd11003, 16'd39160, 16'd44279, 16'd35719, 16'd24066, 16'd25449, 16'd46406, 16'd8308});
	test_expansion(128'h05fe1e030799d1b6f517935166f04808, {16'd15895, 16'd61291, 16'd54172, 16'd28900, 16'd22545, 16'd25178, 16'd57284, 16'd14916, 16'd56519, 16'd27539, 16'd44489, 16'd35597, 16'd58333, 16'd19696, 16'd55844, 16'd58330, 16'd3470, 16'd46938, 16'd30996, 16'd65411, 16'd9089, 16'd37078, 16'd24922, 16'd60205, 16'd61310, 16'd45934});
	test_expansion(128'he34189f88764e8d199be3d157fe824a3, {16'd64116, 16'd32565, 16'd47623, 16'd28413, 16'd3722, 16'd47406, 16'd6992, 16'd41913, 16'd32176, 16'd51854, 16'd57847, 16'd64063, 16'd10440, 16'd65025, 16'd20670, 16'd53498, 16'd13473, 16'd12046, 16'd42658, 16'd35874, 16'd58862, 16'd57339, 16'd20042, 16'd51438, 16'd25714, 16'd62409});
	test_expansion(128'h9782254f57d1e0d47bf3749ba873ff06, {16'd49535, 16'd58628, 16'd20881, 16'd4827, 16'd43608, 16'd54968, 16'd34404, 16'd45140, 16'd55807, 16'd25337, 16'd35146, 16'd13539, 16'd37162, 16'd62767, 16'd47173, 16'd46853, 16'd9454, 16'd45865, 16'd9353, 16'd49026, 16'd6326, 16'd19068, 16'd34166, 16'd43821, 16'd34086, 16'd46704});
	test_expansion(128'hb75d7c006e2d6c2f50c22d4b19ed5e7a, {16'd42934, 16'd2459, 16'd28354, 16'd21748, 16'd59801, 16'd41774, 16'd7299, 16'd16580, 16'd16493, 16'd43817, 16'd62245, 16'd60266, 16'd12169, 16'd24187, 16'd24993, 16'd17590, 16'd55590, 16'd54467, 16'd59184, 16'd26368, 16'd25623, 16'd62067, 16'd30380, 16'd17671, 16'd55756, 16'd12968});
	test_expansion(128'h4fb295d06e3aebfa554361e2e476fd25, {16'd53026, 16'd39931, 16'd28421, 16'd15688, 16'd53220, 16'd11464, 16'd254, 16'd21307, 16'd56416, 16'd48718, 16'd54460, 16'd58833, 16'd16255, 16'd29128, 16'd8995, 16'd27061, 16'd42720, 16'd36074, 16'd58977, 16'd60491, 16'd49146, 16'd49737, 16'd23352, 16'd8053, 16'd37631, 16'd59532});
	test_expansion(128'h05c445f856685a7b386743ba6c70fc39, {16'd32849, 16'd37731, 16'd53709, 16'd17517, 16'd38092, 16'd65003, 16'd14328, 16'd865, 16'd25439, 16'd52149, 16'd7037, 16'd59347, 16'd5173, 16'd13472, 16'd52564, 16'd12018, 16'd25443, 16'd21938, 16'd13918, 16'd58898, 16'd61958, 16'd13706, 16'd44216, 16'd23223, 16'd13324, 16'd39231});
	test_expansion(128'h848e8d7c191b7d070b8bdd148380084a, {16'd25238, 16'd64319, 16'd54372, 16'd55465, 16'd21360, 16'd59541, 16'd50898, 16'd6135, 16'd41389, 16'd46079, 16'd19345, 16'd59992, 16'd63992, 16'd38333, 16'd17715, 16'd11448, 16'd46050, 16'd63268, 16'd51794, 16'd59139, 16'd23749, 16'd18652, 16'd60187, 16'd28615, 16'd42125, 16'd44595});
	test_expansion(128'h566b50e4a0c2da51c81c5c5fbc517aab, {16'd9987, 16'd37936, 16'd52143, 16'd61055, 16'd22249, 16'd40625, 16'd35658, 16'd11758, 16'd43864, 16'd20024, 16'd8261, 16'd43564, 16'd64057, 16'd13248, 16'd36289, 16'd44515, 16'd45195, 16'd16381, 16'd62424, 16'd39607, 16'd16019, 16'd18082, 16'd42929, 16'd58502, 16'd3026, 16'd53890});
	test_expansion(128'hae893a5122242a387616a7fedc215e44, {16'd21984, 16'd29214, 16'd64250, 16'd29657, 16'd1574, 16'd35316, 16'd10153, 16'd18899, 16'd31207, 16'd65357, 16'd31963, 16'd61081, 16'd32541, 16'd61475, 16'd16548, 16'd55494, 16'd29233, 16'd14541, 16'd13917, 16'd12873, 16'd14037, 16'd1045, 16'd56148, 16'd49048, 16'd47597, 16'd34564});
	test_expansion(128'h1c9304560bd10d185f6f657415eae15c, {16'd23915, 16'd20161, 16'd10797, 16'd5977, 16'd26137, 16'd56781, 16'd52480, 16'd10958, 16'd8337, 16'd48885, 16'd25355, 16'd49799, 16'd63098, 16'd10585, 16'd15396, 16'd58866, 16'd6259, 16'd58472, 16'd35214, 16'd17764, 16'd32502, 16'd36463, 16'd60365, 16'd19367, 16'd30762, 16'd58353});
	test_expansion(128'h96e5ca34b9256ff049d40e91e3715cf5, {16'd16904, 16'd39316, 16'd24781, 16'd52133, 16'd38702, 16'd57396, 16'd36157, 16'd30711, 16'd49209, 16'd36832, 16'd42691, 16'd62670, 16'd1554, 16'd5980, 16'd49395, 16'd28154, 16'd43295, 16'd16075, 16'd21582, 16'd32292, 16'd64826, 16'd11591, 16'd13208, 16'd9976, 16'd26656, 16'd45861});
	test_expansion(128'h084e1816d559e8e481972f3c77d1a716, {16'd24751, 16'd39835, 16'd8750, 16'd48481, 16'd1618, 16'd3604, 16'd43747, 16'd44136, 16'd6279, 16'd35041, 16'd61172, 16'd25464, 16'd13284, 16'd6878, 16'd53053, 16'd46817, 16'd39530, 16'd42864, 16'd53603, 16'd34970, 16'd27693, 16'd41702, 16'd42097, 16'd55221, 16'd30994, 16'd9447});
	test_expansion(128'hbaeca3534445121c0e4cf38caf38bb18, {16'd47151, 16'd53265, 16'd46825, 16'd38943, 16'd44959, 16'd58124, 16'd50998, 16'd15273, 16'd44230, 16'd62357, 16'd40909, 16'd2032, 16'd35399, 16'd51764, 16'd12792, 16'd26779, 16'd52648, 16'd11520, 16'd50306, 16'd17803, 16'd61896, 16'd13981, 16'd9247, 16'd51336, 16'd45536, 16'd54948});
	test_expansion(128'h911db24497442430cd0fafd663aca9ea, {16'd22379, 16'd56585, 16'd43966, 16'd55532, 16'd48341, 16'd28608, 16'd22278, 16'd54803, 16'd13499, 16'd14111, 16'd64028, 16'd60514, 16'd30964, 16'd57290, 16'd7042, 16'd57346, 16'd46425, 16'd9090, 16'd1826, 16'd60000, 16'd41933, 16'd51504, 16'd56246, 16'd15762, 16'd1119, 16'd37377});
	test_expansion(128'ha741d716ade97a4d257e3810458d2ccc, {16'd52107, 16'd25863, 16'd57779, 16'd3079, 16'd65091, 16'd29108, 16'd56248, 16'd31291, 16'd9628, 16'd21543, 16'd23005, 16'd704, 16'd19676, 16'd913, 16'd34757, 16'd45622, 16'd25492, 16'd65080, 16'd37016, 16'd34830, 16'd38047, 16'd40942, 16'd4955, 16'd26254, 16'd60497, 16'd46441});
	test_expansion(128'hf372f012b6a08a556738637654eca55f, {16'd50624, 16'd49993, 16'd27553, 16'd45170, 16'd27516, 16'd8615, 16'd11369, 16'd58734, 16'd16022, 16'd34235, 16'd5859, 16'd12332, 16'd47192, 16'd25931, 16'd61688, 16'd33366, 16'd48649, 16'd13394, 16'd50196, 16'd15237, 16'd7293, 16'd23323, 16'd42969, 16'd30255, 16'd21881, 16'd59160});
	test_expansion(128'hb83984428948c1cd576679cac668297d, {16'd35570, 16'd61539, 16'd16478, 16'd59083, 16'd41491, 16'd57012, 16'd48041, 16'd62949, 16'd14435, 16'd52771, 16'd42649, 16'd18236, 16'd32682, 16'd49546, 16'd22855, 16'd60190, 16'd28094, 16'd64126, 16'd1137, 16'd10668, 16'd42326, 16'd41261, 16'd11631, 16'd22997, 16'd56804, 16'd1595});
	test_expansion(128'h98e14fed9377c0841c40467b312b5936, {16'd4591, 16'd64889, 16'd47583, 16'd52308, 16'd4200, 16'd25889, 16'd36811, 16'd9292, 16'd30507, 16'd2985, 16'd60656, 16'd27585, 16'd34129, 16'd20660, 16'd34592, 16'd21293, 16'd61920, 16'd28111, 16'd3009, 16'd24289, 16'd35703, 16'd49427, 16'd3215, 16'd10299, 16'd37116, 16'd271});
	test_expansion(128'hc285edcc6cb73e23add2d4c602062aef, {16'd29700, 16'd52839, 16'd44599, 16'd37447, 16'd30297, 16'd46717, 16'd32041, 16'd15417, 16'd20653, 16'd39247, 16'd27725, 16'd18218, 16'd45515, 16'd42338, 16'd12127, 16'd1974, 16'd45578, 16'd2657, 16'd62777, 16'd52973, 16'd25779, 16'd50336, 16'd19341, 16'd25460, 16'd42550, 16'd42023});
	test_expansion(128'h55361d8dfeb7b60adf752dff7e2f8759, {16'd1763, 16'd31182, 16'd4307, 16'd3650, 16'd6856, 16'd55681, 16'd13084, 16'd17564, 16'd8118, 16'd58600, 16'd10068, 16'd43207, 16'd57649, 16'd65060, 16'd2377, 16'd42209, 16'd8251, 16'd22130, 16'd40861, 16'd26205, 16'd43791, 16'd51400, 16'd28809, 16'd18320, 16'd15113, 16'd54632});
	test_expansion(128'hbdc87303dcf7fbab7eb7d8ac17cc685b, {16'd54988, 16'd31525, 16'd61236, 16'd52964, 16'd10173, 16'd24753, 16'd464, 16'd5855, 16'd17330, 16'd533, 16'd24379, 16'd23269, 16'd31412, 16'd30891, 16'd55780, 16'd31395, 16'd4973, 16'd22188, 16'd43592, 16'd50, 16'd7012, 16'd20444, 16'd5806, 16'd63375, 16'd36869, 16'd26623});
	test_expansion(128'h418e797b2c228d2cc7e19b42b43e43b7, {16'd10998, 16'd2941, 16'd51082, 16'd55462, 16'd38718, 16'd51905, 16'd28538, 16'd31292, 16'd63662, 16'd45234, 16'd33137, 16'd51551, 16'd57194, 16'd61727, 16'd42286, 16'd41361, 16'd12104, 16'd62217, 16'd44273, 16'd11947, 16'd28430, 16'd18849, 16'd62362, 16'd55752, 16'd50479, 16'd41001});
	test_expansion(128'h5a64594aa78cc031bc8715c9bb4faa9e, {16'd38101, 16'd53833, 16'd60853, 16'd20442, 16'd45499, 16'd12416, 16'd792, 16'd51050, 16'd48521, 16'd28725, 16'd39815, 16'd43798, 16'd49968, 16'd40590, 16'd1310, 16'd62458, 16'd55238, 16'd13179, 16'd50789, 16'd50630, 16'd20132, 16'd9805, 16'd61404, 16'd64986, 16'd50809, 16'd26814});
	test_expansion(128'ha43e1a23b53095d8edc75134cc0ef260, {16'd4949, 16'd64254, 16'd55046, 16'd27381, 16'd65363, 16'd43362, 16'd35089, 16'd30554, 16'd19160, 16'd40167, 16'd59032, 16'd37601, 16'd53500, 16'd52927, 16'd1114, 16'd23204, 16'd8731, 16'd57381, 16'd51758, 16'd9374, 16'd33567, 16'd37358, 16'd17117, 16'd56941, 16'd21429, 16'd63724});
	test_expansion(128'h12a1052777e9dcbe84668ee9569943af, {16'd63490, 16'd13848, 16'd12878, 16'd30283, 16'd64364, 16'd4547, 16'd51706, 16'd30325, 16'd22572, 16'd37299, 16'd33384, 16'd1837, 16'd15387, 16'd7851, 16'd12226, 16'd16487, 16'd19651, 16'd37308, 16'd42376, 16'd17689, 16'd29160, 16'd11009, 16'd49424, 16'd21689, 16'd11689, 16'd7275});
	test_expansion(128'h76541b94a7ab5f078bf7d5761a6a0f3f, {16'd19045, 16'd30154, 16'd30292, 16'd39504, 16'd11838, 16'd12026, 16'd25851, 16'd39822, 16'd49748, 16'd16491, 16'd2023, 16'd49136, 16'd9199, 16'd14079, 16'd49147, 16'd5184, 16'd32405, 16'd3156, 16'd10276, 16'd16591, 16'd44829, 16'd38088, 16'd12788, 16'd26742, 16'd2735, 16'd48374});
	test_expansion(128'hae705845d9c4189cde37e37927b2dcb4, {16'd43145, 16'd64414, 16'd33256, 16'd27297, 16'd35040, 16'd42712, 16'd64968, 16'd32165, 16'd26952, 16'd7716, 16'd22011, 16'd39878, 16'd5420, 16'd12868, 16'd22771, 16'd30709, 16'd78, 16'd7227, 16'd4172, 16'd13356, 16'd7599, 16'd29994, 16'd40808, 16'd15670, 16'd62626, 16'd34712});
	test_expansion(128'h0400e1d06b6330c53fb378d3496d48fb, {16'd16273, 16'd50977, 16'd7771, 16'd53304, 16'd18700, 16'd30324, 16'd47325, 16'd31253, 16'd45618, 16'd64010, 16'd44822, 16'd54233, 16'd15904, 16'd42504, 16'd53576, 16'd22087, 16'd41274, 16'd16273, 16'd30808, 16'd42222, 16'd10299, 16'd58169, 16'd29193, 16'd21308, 16'd46814, 16'd54126});
	test_expansion(128'h81213d280ddc3ad79f8b5e20897c46cf, {16'd7222, 16'd405, 16'd44092, 16'd52588, 16'd64755, 16'd15114, 16'd40876, 16'd59277, 16'd44023, 16'd5147, 16'd54311, 16'd52866, 16'd40021, 16'd43463, 16'd25498, 16'd20225, 16'd28790, 16'd31717, 16'd17121, 16'd22058, 16'd48634, 16'd449, 16'd15744, 16'd15052, 16'd58290, 16'd19784});
	test_expansion(128'h2c7139aa72bb40b14018066eeb496571, {16'd23800, 16'd17412, 16'd60564, 16'd22311, 16'd41448, 16'd24068, 16'd3880, 16'd20795, 16'd12195, 16'd57727, 16'd15672, 16'd32003, 16'd42166, 16'd48929, 16'd50700, 16'd46274, 16'd46787, 16'd50642, 16'd18162, 16'd54265, 16'd4890, 16'd58548, 16'd39698, 16'd28879, 16'd54363, 16'd36850});
	test_expansion(128'h024890abee94922748f7cb8a75933d4b, {16'd21762, 16'd945, 16'd30070, 16'd331, 16'd47254, 16'd38117, 16'd38828, 16'd34445, 16'd60873, 16'd26402, 16'd26729, 16'd7324, 16'd26630, 16'd34803, 16'd60069, 16'd28716, 16'd65474, 16'd61675, 16'd60668, 16'd8568, 16'd7894, 16'd17266, 16'd45642, 16'd6313, 16'd15294, 16'd34491});
	test_expansion(128'hf79eac0fa2a2980c248328d899134ab3, {16'd12404, 16'd5274, 16'd22531, 16'd1278, 16'd50754, 16'd31308, 16'd43690, 16'd64575, 16'd53709, 16'd28454, 16'd37200, 16'd28116, 16'd2541, 16'd31676, 16'd51356, 16'd5925, 16'd3490, 16'd33033, 16'd57574, 16'd49242, 16'd28006, 16'd22536, 16'd45999, 16'd61933, 16'd6467, 16'd53535});
	test_expansion(128'h664c2ab7014c26528e921b45d01124ad, {16'd64259, 16'd28562, 16'd49410, 16'd43656, 16'd11386, 16'd57264, 16'd20902, 16'd55736, 16'd12622, 16'd48499, 16'd20603, 16'd54359, 16'd43510, 16'd11036, 16'd52108, 16'd34106, 16'd55168, 16'd37750, 16'd23430, 16'd22171, 16'd41394, 16'd51612, 16'd62982, 16'd21153, 16'd38636, 16'd63630});
	test_expansion(128'hb7dfdb8040a08e2fb6b048762a38ca14, {16'd11813, 16'd63822, 16'd32221, 16'd18960, 16'd63965, 16'd11943, 16'd12535, 16'd3964, 16'd27538, 16'd39958, 16'd44487, 16'd49192, 16'd13229, 16'd23657, 16'd2549, 16'd50520, 16'd63739, 16'd45966, 16'd43255, 16'd25010, 16'd20880, 16'd21116, 16'd64091, 16'd18314, 16'd25118, 16'd31126});
	test_expansion(128'h50ee00364b831a1ab9309478a9979b91, {16'd22129, 16'd21378, 16'd55389, 16'd32436, 16'd634, 16'd18539, 16'd10549, 16'd64028, 16'd61902, 16'd51872, 16'd62675, 16'd39248, 16'd32816, 16'd36002, 16'd34941, 16'd42897, 16'd61942, 16'd32638, 16'd64065, 16'd63814, 16'd8629, 16'd16651, 16'd11782, 16'd16093, 16'd28516, 16'd45163});
	test_expansion(128'h9928435ba4fc35bcad7c27402341b40a, {16'd42770, 16'd28789, 16'd52953, 16'd58319, 16'd3210, 16'd46093, 16'd36855, 16'd24101, 16'd23166, 16'd30375, 16'd33430, 16'd12795, 16'd63407, 16'd26245, 16'd6697, 16'd42490, 16'd40727, 16'd43920, 16'd60350, 16'd31026, 16'd18174, 16'd34270, 16'd39706, 16'd58189, 16'd5167, 16'd16126});
	test_expansion(128'hdbd76045c243161adfbd647b7a349f92, {16'd15886, 16'd17256, 16'd23856, 16'd60808, 16'd64613, 16'd25991, 16'd58123, 16'd24182, 16'd9991, 16'd65068, 16'd5569, 16'd36155, 16'd37021, 16'd58335, 16'd43262, 16'd47415, 16'd25943, 16'd61372, 16'd50159, 16'd15911, 16'd6730, 16'd34548, 16'd43673, 16'd30741, 16'd38521, 16'd19568});
	test_expansion(128'h1d12873e067f48b15c7cf4213a10953e, {16'd8264, 16'd59749, 16'd32997, 16'd16961, 16'd11000, 16'd56926, 16'd58980, 16'd29740, 16'd27172, 16'd9090, 16'd6559, 16'd50721, 16'd61757, 16'd49852, 16'd14585, 16'd60835, 16'd54117, 16'd17583, 16'd35262, 16'd63939, 16'd48504, 16'd20197, 16'd58510, 16'd28149, 16'd40428, 16'd11508});
	test_expansion(128'h70ade449c97cad905a79a2be0fe2105b, {16'd40554, 16'd26038, 16'd64133, 16'd64024, 16'd12422, 16'd21175, 16'd5514, 16'd38236, 16'd25349, 16'd37333, 16'd32806, 16'd35633, 16'd40286, 16'd57157, 16'd22709, 16'd39712, 16'd53282, 16'd61615, 16'd27124, 16'd10177, 16'd12853, 16'd56862, 16'd30147, 16'd8125, 16'd40912, 16'd51929});
	test_expansion(128'h5a156459aa16f27aa23981c05c511b78, {16'd61319, 16'd40990, 16'd51363, 16'd58063, 16'd39438, 16'd59978, 16'd16359, 16'd15207, 16'd60547, 16'd60542, 16'd3576, 16'd47890, 16'd19984, 16'd13211, 16'd30258, 16'd48045, 16'd65377, 16'd24056, 16'd4119, 16'd25892, 16'd23038, 16'd11634, 16'd54727, 16'd3470, 16'd30068, 16'd24429});
	test_expansion(128'hc397a8637c568384c7fa2166b39ffc29, {16'd5858, 16'd58272, 16'd22068, 16'd27935, 16'd29897, 16'd28404, 16'd40975, 16'd23844, 16'd53113, 16'd30289, 16'd24136, 16'd61851, 16'd51280, 16'd9927, 16'd42848, 16'd26183, 16'd20779, 16'd15609, 16'd32029, 16'd19268, 16'd23162, 16'd45179, 16'd34444, 16'd54401, 16'd28982, 16'd10052});
	test_expansion(128'h609dbedd295aed6e3a5ac187131d21d6, {16'd33698, 16'd61722, 16'd3199, 16'd47406, 16'd48775, 16'd50123, 16'd34015, 16'd4111, 16'd53245, 16'd62892, 16'd894, 16'd60680, 16'd51405, 16'd55490, 16'd39379, 16'd30735, 16'd2724, 16'd39371, 16'd29063, 16'd10503, 16'd10659, 16'd43879, 16'd37673, 16'd5586, 16'd22724, 16'd58064});
	test_expansion(128'h8598e6d41ef4514e956ef6ed9e30015c, {16'd2047, 16'd31075, 16'd38718, 16'd36626, 16'd64571, 16'd11035, 16'd16439, 16'd27621, 16'd21339, 16'd5207, 16'd28040, 16'd1985, 16'd40759, 16'd54924, 16'd33625, 16'd54124, 16'd29732, 16'd61275, 16'd39917, 16'd25698, 16'd16684, 16'd33737, 16'd49738, 16'd54242, 16'd49006, 16'd7532});
	test_expansion(128'h67209199a3a95de69444b1feaf565fff, {16'd8651, 16'd4425, 16'd39376, 16'd49940, 16'd19454, 16'd1459, 16'd41053, 16'd20275, 16'd37311, 16'd56886, 16'd54649, 16'd55064, 16'd11970, 16'd40107, 16'd45337, 16'd52745, 16'd36385, 16'd22347, 16'd11147, 16'd32845, 16'd44270, 16'd42983, 16'd63334, 16'd61720, 16'd47583, 16'd34112});
	test_expansion(128'h0215266809cbf7f6dbdb18ecc2b5cf61, {16'd63780, 16'd4202, 16'd57548, 16'd36241, 16'd20639, 16'd14781, 16'd45213, 16'd16563, 16'd29738, 16'd25275, 16'd34544, 16'd37979, 16'd9691, 16'd37263, 16'd64794, 16'd43768, 16'd9583, 16'd35863, 16'd8379, 16'd34612, 16'd22872, 16'd14081, 16'd7368, 16'd1780, 16'd62391, 16'd17481});
	test_expansion(128'hd3886ef485763e376d3b8843fb11307f, {16'd57193, 16'd60074, 16'd40352, 16'd65343, 16'd25047, 16'd39926, 16'd5070, 16'd36749, 16'd3419, 16'd33366, 16'd42457, 16'd20398, 16'd64475, 16'd27316, 16'd24641, 16'd23974, 16'd44834, 16'd20549, 16'd11686, 16'd25116, 16'd64599, 16'd33423, 16'd42114, 16'd14579, 16'd10046, 16'd19539});
	test_expansion(128'h54b68b91518c0e21ec85e7da47e80c8f, {16'd27916, 16'd902, 16'd27691, 16'd2842, 16'd19939, 16'd11151, 16'd60905, 16'd34248, 16'd18202, 16'd61507, 16'd51610, 16'd41540, 16'd11549, 16'd33666, 16'd14982, 16'd35092, 16'd57465, 16'd5418, 16'd34863, 16'd32470, 16'd57741, 16'd61765, 16'd8553, 16'd63816, 16'd19770, 16'd42840});
	test_expansion(128'h072cdbcc089cc26ccbf6681403ee82a1, {16'd9810, 16'd57789, 16'd53907, 16'd24054, 16'd64470, 16'd53214, 16'd56832, 16'd40811, 16'd42647, 16'd22368, 16'd47442, 16'd17798, 16'd31770, 16'd61216, 16'd10479, 16'd47783, 16'd16641, 16'd4446, 16'd36645, 16'd6743, 16'd41098, 16'd46936, 16'd41913, 16'd61176, 16'd9183, 16'd25463});
	test_expansion(128'h02d3ac7e1dacb0a88f9d998283ca5b85, {16'd58196, 16'd56015, 16'd22302, 16'd58511, 16'd27039, 16'd22532, 16'd44996, 16'd30205, 16'd64420, 16'd3526, 16'd27572, 16'd19369, 16'd58916, 16'd1127, 16'd49345, 16'd49112, 16'd9037, 16'd48577, 16'd22203, 16'd5975, 16'd17145, 16'd31192, 16'd40271, 16'd41109, 16'd26387, 16'd6912});
	test_expansion(128'hdf8dabf42964f1b8e9f2bb024be1841e, {16'd51981, 16'd43518, 16'd56016, 16'd19143, 16'd22302, 16'd46269, 16'd53642, 16'd58969, 16'd58176, 16'd63830, 16'd46456, 16'd53759, 16'd45596, 16'd53587, 16'd10445, 16'd53440, 16'd51429, 16'd12817, 16'd37070, 16'd31359, 16'd13919, 16'd54211, 16'd60930, 16'd36953, 16'd57691, 16'd36764});
	test_expansion(128'h2f461dcdf39b9ba2fb774cae27f9f850, {16'd42891, 16'd64098, 16'd59015, 16'd6299, 16'd7582, 16'd40572, 16'd52590, 16'd10670, 16'd12712, 16'd25371, 16'd44961, 16'd60488, 16'd19133, 16'd5262, 16'd43785, 16'd59207, 16'd33498, 16'd27812, 16'd3048, 16'd52226, 16'd31408, 16'd13874, 16'd57542, 16'd53892, 16'd51890, 16'd40966});
	test_expansion(128'h27f9c52fdc444de6d5961a4934d705d8, {16'd28115, 16'd39844, 16'd12617, 16'd37150, 16'd8043, 16'd57590, 16'd45536, 16'd6048, 16'd53038, 16'd11882, 16'd23989, 16'd64805, 16'd33898, 16'd54689, 16'd30089, 16'd52917, 16'd26864, 16'd3268, 16'd21612, 16'd59067, 16'd52253, 16'd63765, 16'd60640, 16'd16043, 16'd50668, 16'd49831});
	test_expansion(128'h4317a3ea3470a98b972bd361cc7bca22, {16'd4720, 16'd60042, 16'd32092, 16'd14962, 16'd9049, 16'd7, 16'd45414, 16'd60410, 16'd32413, 16'd63018, 16'd33278, 16'd13284, 16'd12660, 16'd56571, 16'd38675, 16'd53077, 16'd46841, 16'd27542, 16'd37697, 16'd40205, 16'd10744, 16'd21122, 16'd61605, 16'd24320, 16'd668, 16'd16037});
	test_expansion(128'hc30bf0c9579fb35e32d8d304e69479a7, {16'd48669, 16'd18256, 16'd22400, 16'd50179, 16'd18251, 16'd16489, 16'd5685, 16'd515, 16'd28139, 16'd38275, 16'd50762, 16'd32150, 16'd2880, 16'd4069, 16'd23441, 16'd9161, 16'd28283, 16'd1993, 16'd31831, 16'd26617, 16'd15834, 16'd34096, 16'd64668, 16'd43708, 16'd63920, 16'd31344});
	test_expansion(128'h4783e423a46d42ff630706c78ebbe9d5, {16'd21752, 16'd50149, 16'd6144, 16'd12331, 16'd60419, 16'd3886, 16'd62585, 16'd3922, 16'd64224, 16'd14292, 16'd56929, 16'd8946, 16'd17753, 16'd53681, 16'd31560, 16'd12159, 16'd55328, 16'd37014, 16'd46334, 16'd45671, 16'd51084, 16'd19451, 16'd54354, 16'd7291, 16'd61111, 16'd63079});
	test_expansion(128'he6c93cd0e3c41e077cc501ecb0531e27, {16'd53691, 16'd723, 16'd37443, 16'd64600, 16'd41441, 16'd8038, 16'd43768, 16'd56804, 16'd34409, 16'd45768, 16'd29856, 16'd60880, 16'd55800, 16'd12618, 16'd37400, 16'd6365, 16'd14575, 16'd33313, 16'd52150, 16'd7592, 16'd32481, 16'd44327, 16'd34434, 16'd29037, 16'd10789, 16'd21247});
	test_expansion(128'h6f565b92df013d26fbda155b84002370, {16'd13498, 16'd43278, 16'd44843, 16'd45081, 16'd45366, 16'd42708, 16'd10965, 16'd58125, 16'd13587, 16'd42892, 16'd18976, 16'd13062, 16'd20826, 16'd20479, 16'd53412, 16'd51651, 16'd16819, 16'd20496, 16'd35282, 16'd42740, 16'd8255, 16'd36707, 16'd9259, 16'd37178, 16'd46103, 16'd511});
	test_expansion(128'h582fa0298a0ea0e5e234a57583d078bb, {16'd49809, 16'd37337, 16'd21924, 16'd62284, 16'd7747, 16'd6106, 16'd39900, 16'd33460, 16'd28868, 16'd57861, 16'd25783, 16'd24698, 16'd62998, 16'd47646, 16'd36675, 16'd59833, 16'd8253, 16'd3012, 16'd39987, 16'd6021, 16'd5885, 16'd54546, 16'd3256, 16'd53455, 16'd3141, 16'd35223});
	test_expansion(128'h3a0805702f3d7a029a92239eaf0c6dd0, {16'd20100, 16'd6763, 16'd30190, 16'd55896, 16'd59368, 16'd23848, 16'd49361, 16'd41784, 16'd12218, 16'd51594, 16'd5108, 16'd19668, 16'd18156, 16'd63025, 16'd24116, 16'd40275, 16'd45120, 16'd30144, 16'd54361, 16'd52001, 16'd17319, 16'd37555, 16'd17537, 16'd1002, 16'd54045, 16'd49859});
	test_expansion(128'h4e8168bfcda85a2eb5bd836130359230, {16'd31638, 16'd6633, 16'd46320, 16'd47240, 16'd48320, 16'd42548, 16'd1380, 16'd25161, 16'd26024, 16'd2839, 16'd28503, 16'd62499, 16'd58586, 16'd46149, 16'd20347, 16'd55363, 16'd20180, 16'd26032, 16'd34715, 16'd40339, 16'd53256, 16'd8881, 16'd49599, 16'd60914, 16'd4606, 16'd33482});
	test_expansion(128'h7aaff58e1105d1fa62fd5cfe23dabccc, {16'd7947, 16'd43600, 16'd5251, 16'd12697, 16'd50779, 16'd52301, 16'd1168, 16'd10856, 16'd21500, 16'd49650, 16'd275, 16'd605, 16'd46446, 16'd55211, 16'd43666, 16'd6984, 16'd56521, 16'd10661, 16'd4888, 16'd52260, 16'd50167, 16'd21002, 16'd49709, 16'd58039, 16'd10244, 16'd41129});
	test_expansion(128'hd013aa61098bc9ad1f53f92263c85eb6, {16'd40024, 16'd50858, 16'd63598, 16'd61909, 16'd38980, 16'd53609, 16'd18805, 16'd19547, 16'd11088, 16'd33953, 16'd60931, 16'd42689, 16'd14115, 16'd7381, 16'd26498, 16'd39495, 16'd1282, 16'd39137, 16'd53803, 16'd37559, 16'd23072, 16'd17733, 16'd24115, 16'd35313, 16'd59399, 16'd10454});
	test_expansion(128'h8589a657e82b4a63770ffeb0e8ba758c, {16'd53079, 16'd28160, 16'd9630, 16'd7051, 16'd64307, 16'd11056, 16'd19310, 16'd33477, 16'd8680, 16'd25799, 16'd20056, 16'd5405, 16'd49234, 16'd17444, 16'd43283, 16'd2597, 16'd54040, 16'd59022, 16'd22424, 16'd1833, 16'd44602, 16'd23430, 16'd32604, 16'd11169, 16'd12991, 16'd63476});
	test_expansion(128'h1dbab5d2eb5c2b39120a9b4847f91027, {16'd71, 16'd12338, 16'd10027, 16'd14093, 16'd11913, 16'd31073, 16'd45234, 16'd36199, 16'd30587, 16'd34772, 16'd59504, 16'd36260, 16'd43654, 16'd15358, 16'd45809, 16'd15721, 16'd43162, 16'd50206, 16'd6574, 16'd56723, 16'd39272, 16'd50448, 16'd20158, 16'd23942, 16'd10860, 16'd65501});
	test_expansion(128'h171ceb837b8b64f821f3bba75a79c957, {16'd2438, 16'd22900, 16'd3532, 16'd63232, 16'd20934, 16'd29074, 16'd31768, 16'd18391, 16'd58776, 16'd2393, 16'd10915, 16'd56084, 16'd7486, 16'd38783, 16'd16782, 16'd25671, 16'd41922, 16'd27167, 16'd29565, 16'd24821, 16'd21102, 16'd38690, 16'd30144, 16'd54192, 16'd50673, 16'd7966});
	test_expansion(128'h5e44ca0844344edbd37b7eaca0a86ab2, {16'd8061, 16'd39407, 16'd35058, 16'd5206, 16'd14705, 16'd61204, 16'd27474, 16'd61916, 16'd55827, 16'd35622, 16'd25555, 16'd4184, 16'd63532, 16'd40237, 16'd16533, 16'd9398, 16'd51415, 16'd42440, 16'd64683, 16'd56159, 16'd8882, 16'd17360, 16'd37073, 16'd9459, 16'd18776, 16'd41801});
	test_expansion(128'hfe76f06760545fc554e4402e57f116fd, {16'd54544, 16'd29034, 16'd59274, 16'd42091, 16'd36763, 16'd62500, 16'd5973, 16'd15839, 16'd58138, 16'd37437, 16'd5594, 16'd54632, 16'd41907, 16'd41642, 16'd33856, 16'd1666, 16'd59930, 16'd46846, 16'd62295, 16'd46322, 16'd37800, 16'd39931, 16'd53349, 16'd16369, 16'd53165, 16'd1009});
	test_expansion(128'he530cf4bc93573d0a523fad68ee94a6f, {16'd58618, 16'd41358, 16'd46428, 16'd62962, 16'd48784, 16'd10738, 16'd34884, 16'd60817, 16'd40323, 16'd4741, 16'd48054, 16'd43337, 16'd26831, 16'd14457, 16'd63174, 16'd36601, 16'd14903, 16'd42176, 16'd4883, 16'd62985, 16'd26281, 16'd29601, 16'd18533, 16'd54760, 16'd61583, 16'd15804});
	test_expansion(128'hb1c963e4eeecd051bcdff0b7e79f099b, {16'd57003, 16'd36679, 16'd64314, 16'd1060, 16'd43538, 16'd3872, 16'd62094, 16'd58111, 16'd19201, 16'd6167, 16'd54626, 16'd8572, 16'd15422, 16'd39858, 16'd31617, 16'd29501, 16'd60599, 16'd35933, 16'd7598, 16'd13768, 16'd54629, 16'd19304, 16'd23325, 16'd38748, 16'd58049, 16'd1093});
	test_expansion(128'h922b947ce127ee2de0d5611997d7c764, {16'd36025, 16'd3030, 16'd23711, 16'd63662, 16'd29317, 16'd33773, 16'd23162, 16'd54863, 16'd38868, 16'd16618, 16'd27949, 16'd35102, 16'd32909, 16'd1164, 16'd1327, 16'd51509, 16'd33578, 16'd51110, 16'd26865, 16'd36780, 16'd54392, 16'd43841, 16'd51180, 16'd65316, 16'd20268, 16'd410});
	test_expansion(128'ha2c9408d41ff52ae413d0de2f284038e, {16'd49648, 16'd43839, 16'd33749, 16'd10533, 16'd52305, 16'd10848, 16'd28732, 16'd34063, 16'd58703, 16'd1673, 16'd33519, 16'd3361, 16'd7415, 16'd14528, 16'd19014, 16'd65504, 16'd6307, 16'd5375, 16'd50401, 16'd7846, 16'd15017, 16'd48183, 16'd34806, 16'd55328, 16'd25540, 16'd15192});
	test_expansion(128'hf41b7f305a9b4db2b88012bf98766a4c, {16'd31456, 16'd63554, 16'd35912, 16'd8970, 16'd3691, 16'd43231, 16'd36386, 16'd63246, 16'd57904, 16'd25932, 16'd22578, 16'd40241, 16'd20064, 16'd13985, 16'd45613, 16'd6591, 16'd53699, 16'd29972, 16'd27140, 16'd35883, 16'd18668, 16'd30484, 16'd4188, 16'd54852, 16'd15202, 16'd58490});
	test_expansion(128'h15b8349a9d5f475893894398ebab8ab9, {16'd52209, 16'd63268, 16'd46921, 16'd42626, 16'd60133, 16'd63108, 16'd38776, 16'd31870, 16'd44106, 16'd57758, 16'd54585, 16'd55002, 16'd43012, 16'd52088, 16'd60614, 16'd46524, 16'd58510, 16'd23059, 16'd44702, 16'd50099, 16'd58423, 16'd945, 16'd54196, 16'd11596, 16'd2010, 16'd51774});
	test_expansion(128'hdc80a50bb81c5951baddf2d1bbf653f6, {16'd32397, 16'd10659, 16'd33728, 16'd2322, 16'd41793, 16'd14270, 16'd26390, 16'd3398, 16'd26077, 16'd15489, 16'd65352, 16'd14635, 16'd59840, 16'd697, 16'd33509, 16'd26682, 16'd56146, 16'd28617, 16'd17511, 16'd40723, 16'd36668, 16'd54626, 16'd8890, 16'd32744, 16'd32742, 16'd10369});
	test_expansion(128'h824069f932aa484c8f3b7e8b11a0b520, {16'd30883, 16'd59255, 16'd45139, 16'd5858, 16'd39467, 16'd39222, 16'd24453, 16'd56520, 16'd33379, 16'd29587, 16'd34969, 16'd42901, 16'd63873, 16'd12174, 16'd54196, 16'd46949, 16'd29236, 16'd24589, 16'd30118, 16'd56405, 16'd3779, 16'd29924, 16'd33199, 16'd61672, 16'd61499, 16'd51410});
	test_expansion(128'h31f00ee5867688aa2550901be7f2afd1, {16'd23869, 16'd45936, 16'd4508, 16'd23744, 16'd63266, 16'd9596, 16'd20288, 16'd62111, 16'd4161, 16'd15546, 16'd16324, 16'd56657, 16'd25249, 16'd34705, 16'd9360, 16'd4325, 16'd48251, 16'd7557, 16'd35221, 16'd51877, 16'd39236, 16'd38508, 16'd12537, 16'd62172, 16'd15030, 16'd58497});
	test_expansion(128'hbd3d0db0ec3a753df26fe1ce3a4d800b, {16'd28576, 16'd42197, 16'd20548, 16'd10544, 16'd23399, 16'd44154, 16'd19615, 16'd56943, 16'd45063, 16'd62209, 16'd35796, 16'd62117, 16'd49408, 16'd33743, 16'd52540, 16'd25819, 16'd37353, 16'd58835, 16'd54247, 16'd55812, 16'd7294, 16'd15429, 16'd5500, 16'd1577, 16'd17297, 16'd59108});
	test_expansion(128'hf4aae9ba9203e0314cc942dfa9e9da85, {16'd54064, 16'd53140, 16'd19180, 16'd47774, 16'd16126, 16'd61135, 16'd11269, 16'd48301, 16'd42169, 16'd9624, 16'd24510, 16'd34349, 16'd1915, 16'd64878, 16'd47854, 16'd63360, 16'd65051, 16'd2001, 16'd17186, 16'd10706, 16'd32872, 16'd35334, 16'd34009, 16'd39833, 16'd52848, 16'd31141});
	test_expansion(128'h35e45167152bcb00a671f30989344a34, {16'd6178, 16'd63564, 16'd31332, 16'd48028, 16'd48597, 16'd27589, 16'd10366, 16'd14859, 16'd39255, 16'd5095, 16'd52917, 16'd27672, 16'd7583, 16'd36203, 16'd60513, 16'd9396, 16'd51856, 16'd40284, 16'd16496, 16'd24847, 16'd60143, 16'd60998, 16'd36321, 16'd39658, 16'd52691, 16'd23182});
	test_expansion(128'hafabc02e488a6cf377ace17c1080c33e, {16'd12011, 16'd10604, 16'd16216, 16'd53227, 16'd64023, 16'd22551, 16'd2048, 16'd27829, 16'd11511, 16'd15846, 16'd61065, 16'd11276, 16'd31505, 16'd39200, 16'd60601, 16'd54388, 16'd46832, 16'd27585, 16'd14622, 16'd62478, 16'd51940, 16'd24938, 16'd11470, 16'd45224, 16'd13838, 16'd10453});
	test_expansion(128'h1eba674f1d33844b80ebe7973bb345f5, {16'd59500, 16'd10949, 16'd31767, 16'd1886, 16'd51537, 16'd43847, 16'd62328, 16'd64615, 16'd41609, 16'd10796, 16'd1098, 16'd58451, 16'd8856, 16'd5377, 16'd12782, 16'd3091, 16'd15593, 16'd23299, 16'd19526, 16'd8533, 16'd10013, 16'd17191, 16'd56891, 16'd47302, 16'd20528, 16'd16050});
	test_expansion(128'hdf54205fe8c7e5d653cd4272601a7341, {16'd27256, 16'd25224, 16'd55629, 16'd43241, 16'd3154, 16'd42970, 16'd7837, 16'd1525, 16'd23692, 16'd61333, 16'd18876, 16'd25143, 16'd15698, 16'd39577, 16'd35257, 16'd58292, 16'd52236, 16'd9447, 16'd60867, 16'd59728, 16'd54652, 16'd43645, 16'd44396, 16'd60253, 16'd6333, 16'd48559});
	test_expansion(128'hd8afdd246931600e4448e8af3d8db8ef, {16'd21172, 16'd27259, 16'd12842, 16'd47037, 16'd7995, 16'd32075, 16'd4342, 16'd9762, 16'd64956, 16'd16758, 16'd41274, 16'd30598, 16'd12642, 16'd15432, 16'd49325, 16'd12008, 16'd5064, 16'd1033, 16'd61230, 16'd8740, 16'd671, 16'd49952, 16'd18685, 16'd30533, 16'd58447, 16'd25228});
	test_expansion(128'hf740e217b8ddb88f50faf3aab866dcfc, {16'd48054, 16'd9957, 16'd24425, 16'd64115, 16'd7054, 16'd24951, 16'd35896, 16'd63307, 16'd50833, 16'd32591, 16'd23490, 16'd1350, 16'd29486, 16'd64432, 16'd27830, 16'd2591, 16'd49041, 16'd6824, 16'd30400, 16'd12104, 16'd29324, 16'd55037, 16'd19620, 16'd30662, 16'd13661, 16'd59297});
	test_expansion(128'h62dc58c4e998757dbf667ed8a391f37f, {16'd12870, 16'd12157, 16'd36527, 16'd42579, 16'd51406, 16'd59537, 16'd34617, 16'd62758, 16'd46379, 16'd49788, 16'd58058, 16'd46791, 16'd63318, 16'd24288, 16'd19155, 16'd20144, 16'd6418, 16'd14919, 16'd53651, 16'd41416, 16'd20674, 16'd64382, 16'd16458, 16'd40135, 16'd29750, 16'd62939});
	test_expansion(128'hde583885b86b46d6fa3ea238beb2cb59, {16'd63790, 16'd61251, 16'd53262, 16'd58596, 16'd772, 16'd33276, 16'd60365, 16'd12910, 16'd89, 16'd43627, 16'd57825, 16'd56648, 16'd25709, 16'd8159, 16'd5975, 16'd27442, 16'd60634, 16'd10281, 16'd24817, 16'd3085, 16'd5005, 16'd64568, 16'd50325, 16'd42284, 16'd60113, 16'd57164});
	test_expansion(128'hc0d81db848ff3d637d24c0aad5e36770, {16'd8515, 16'd54978, 16'd45277, 16'd34443, 16'd30270, 16'd7746, 16'd2961, 16'd16079, 16'd38588, 16'd33250, 16'd61813, 16'd25675, 16'd154, 16'd14845, 16'd64807, 16'd33455, 16'd30592, 16'd38111, 16'd56640, 16'd49512, 16'd23196, 16'd35925, 16'd56608, 16'd44757, 16'd31335, 16'd20660});
	test_expansion(128'hcdd853366e6cf63bbf4d4e8fe45cb107, {16'd5106, 16'd52233, 16'd3011, 16'd24488, 16'd43201, 16'd60527, 16'd45789, 16'd60582, 16'd41699, 16'd47607, 16'd7590, 16'd47771, 16'd62267, 16'd5646, 16'd51768, 16'd12316, 16'd20171, 16'd18001, 16'd61905, 16'd26932, 16'd27519, 16'd8521, 16'd25329, 16'd30749, 16'd47051, 16'd12299});
	test_expansion(128'hf87fc8a9cdf80ad0c4d5cad407bab478, {16'd8491, 16'd26260, 16'd64152, 16'd43237, 16'd39238, 16'd12023, 16'd22895, 16'd30585, 16'd39667, 16'd6484, 16'd32584, 16'd3038, 16'd64610, 16'd12729, 16'd12868, 16'd37433, 16'd32496, 16'd54439, 16'd53430, 16'd62953, 16'd30890, 16'd31947, 16'd55759, 16'd46858, 16'd15913, 16'd13147});
	test_expansion(128'h697bfa16353fb568980704d5c0fdfb1b, {16'd46556, 16'd24014, 16'd4921, 16'd37039, 16'd27942, 16'd37929, 16'd49914, 16'd6056, 16'd32555, 16'd59030, 16'd60688, 16'd15514, 16'd48737, 16'd9708, 16'd46954, 16'd12380, 16'd20705, 16'd2478, 16'd41555, 16'd36327, 16'd3704, 16'd36407, 16'd15241, 16'd33228, 16'd38768, 16'd3064});
	test_expansion(128'h4f92615fefce1841ecf685c4fb758608, {16'd6325, 16'd213, 16'd21296, 16'd46337, 16'd28173, 16'd25433, 16'd30298, 16'd15459, 16'd23856, 16'd22527, 16'd5813, 16'd51834, 16'd27224, 16'd36781, 16'd18684, 16'd59535, 16'd3663, 16'd8950, 16'd15592, 16'd3453, 16'd53865, 16'd48913, 16'd49724, 16'd23518, 16'd10782, 16'd35897});
	test_expansion(128'h87a74b968c3c40cfd185ac5c8a596236, {16'd53988, 16'd5649, 16'd5478, 16'd14941, 16'd5731, 16'd18057, 16'd62574, 16'd28202, 16'd62973, 16'd14976, 16'd63848, 16'd36579, 16'd47264, 16'd10827, 16'd5568, 16'd12199, 16'd39070, 16'd54715, 16'd62061, 16'd39973, 16'd63157, 16'd23983, 16'd39792, 16'd14655, 16'd55486, 16'd1723});
	test_expansion(128'h148ef3449ee87a1fdecf8852b0e7b56f, {16'd43454, 16'd34419, 16'd62903, 16'd10167, 16'd19923, 16'd63297, 16'd23314, 16'd45526, 16'd26812, 16'd45100, 16'd21372, 16'd65516, 16'd28647, 16'd11124, 16'd48852, 16'd30290, 16'd38001, 16'd23391, 16'd16291, 16'd4411, 16'd1027, 16'd3886, 16'd24001, 16'd19251, 16'd13974, 16'd38330});
	test_expansion(128'h45e040f4930588356ab1424698997053, {16'd26256, 16'd21125, 16'd41259, 16'd27642, 16'd19098, 16'd62114, 16'd63362, 16'd44051, 16'd4671, 16'd46408, 16'd44546, 16'd45230, 16'd17919, 16'd13729, 16'd56404, 16'd18373, 16'd43093, 16'd50480, 16'd59769, 16'd45829, 16'd12882, 16'd45128, 16'd31822, 16'd12856, 16'd18668, 16'd37366});
	test_expansion(128'hffc7736efa2ffb15603a8591d93e64ee, {16'd55518, 16'd65381, 16'd42329, 16'd18913, 16'd50266, 16'd38058, 16'd34915, 16'd42968, 16'd33740, 16'd63327, 16'd6191, 16'd5719, 16'd35796, 16'd31340, 16'd61528, 16'd56298, 16'd9446, 16'd11560, 16'd57218, 16'd37909, 16'd246, 16'd45731, 16'd50924, 16'd48749, 16'd4581, 16'd28722});
	test_expansion(128'ha088a1f42314cc2dab382a162f820a23, {16'd14414, 16'd5310, 16'd55665, 16'd48729, 16'd11888, 16'd26412, 16'd14937, 16'd21317, 16'd31201, 16'd14267, 16'd17614, 16'd40794, 16'd9281, 16'd31525, 16'd44828, 16'd23511, 16'd6669, 16'd2058, 16'd28538, 16'd59314, 16'd54926, 16'd52211, 16'd1387, 16'd47338, 16'd6076, 16'd58315});
	test_expansion(128'h5f96c2c240e61a0b3786d91f3e1a0820, {16'd60031, 16'd2304, 16'd59930, 16'd64113, 16'd38286, 16'd46755, 16'd619, 16'd29398, 16'd7712, 16'd23632, 16'd55909, 16'd20529, 16'd2614, 16'd29926, 16'd63619, 16'd27759, 16'd4546, 16'd19974, 16'd913, 16'd21771, 16'd37017, 16'd56971, 16'd27616, 16'd17406, 16'd19446, 16'd23486});
	test_expansion(128'hfc31afcdfb15e1a35a7f1717da1678c2, {16'd40609, 16'd24492, 16'd22104, 16'd65132, 16'd57286, 16'd35801, 16'd41415, 16'd1166, 16'd19483, 16'd43225, 16'd4289, 16'd36908, 16'd62008, 16'd6652, 16'd26404, 16'd38254, 16'd34327, 16'd60788, 16'd4329, 16'd3330, 16'd1540, 16'd3170, 16'd17258, 16'd16465, 16'd13819, 16'd7409});
	test_expansion(128'hf861ed070d95aa04b232ca5168733eb4, {16'd39997, 16'd56056, 16'd11677, 16'd21264, 16'd45817, 16'd16664, 16'd18928, 16'd58247, 16'd18507, 16'd58424, 16'd27605, 16'd13660, 16'd60269, 16'd42216, 16'd33933, 16'd50070, 16'd23616, 16'd16278, 16'd15434, 16'd39188, 16'd16067, 16'd40434, 16'd61709, 16'd28748, 16'd31225, 16'd39286});
	test_expansion(128'hda197d6660585b4a45e4163e337c23c0, {16'd59795, 16'd57357, 16'd23593, 16'd7575, 16'd41346, 16'd59606, 16'd64838, 16'd32293, 16'd29229, 16'd53449, 16'd21215, 16'd46842, 16'd8015, 16'd60623, 16'd52644, 16'd47871, 16'd49354, 16'd28665, 16'd6135, 16'd4997, 16'd24577, 16'd26171, 16'd35628, 16'd47682, 16'd16887, 16'd29873});
	test_expansion(128'h2e90fcfd630a484bffd82bd954bf0a7f, {16'd52267, 16'd33039, 16'd49147, 16'd3312, 16'd12243, 16'd46690, 16'd29635, 16'd12387, 16'd35041, 16'd14137, 16'd21041, 16'd29033, 16'd41307, 16'd13971, 16'd4943, 16'd58968, 16'd37040, 16'd6855, 16'd12169, 16'd16879, 16'd11467, 16'd14977, 16'd38274, 16'd5702, 16'd39232, 16'd63912});
	test_expansion(128'hc1298934c706ad948ee375c7ae13e5e0, {16'd17350, 16'd30708, 16'd56028, 16'd22726, 16'd22819, 16'd5581, 16'd43353, 16'd49311, 16'd46110, 16'd26953, 16'd28356, 16'd9672, 16'd55586, 16'd18883, 16'd33132, 16'd7924, 16'd52186, 16'd63823, 16'd7769, 16'd62259, 16'd54187, 16'd34506, 16'd62001, 16'd20599, 16'd2681, 16'd59269});
	test_expansion(128'hd8cac3917cdb1bfd8c9813ddb54b0813, {16'd44292, 16'd2324, 16'd43226, 16'd18991, 16'd57376, 16'd65383, 16'd60116, 16'd42258, 16'd9260, 16'd18522, 16'd40604, 16'd39528, 16'd12991, 16'd48724, 16'd28465, 16'd45268, 16'd64841, 16'd11910, 16'd30474, 16'd60051, 16'd23318, 16'd26132, 16'd11506, 16'd4104, 16'd2098, 16'd57366});
	test_expansion(128'h68dc4f5bb63fd41df8f2ddc1717613cc, {16'd14763, 16'd45348, 16'd38692, 16'd41854, 16'd50865, 16'd21337, 16'd25865, 16'd26143, 16'd14621, 16'd59362, 16'd60106, 16'd52530, 16'd48648, 16'd27435, 16'd39352, 16'd27878, 16'd25383, 16'd45946, 16'd7199, 16'd19362, 16'd34171, 16'd26822, 16'd57306, 16'd6775, 16'd17616, 16'd25202});
	test_expansion(128'h79ab8ece0bba7d6cca6b8f394a406be5, {16'd25837, 16'd52913, 16'd14447, 16'd17091, 16'd27628, 16'd52421, 16'd9552, 16'd61821, 16'd54054, 16'd47545, 16'd40605, 16'd11444, 16'd24852, 16'd57263, 16'd20494, 16'd63187, 16'd57943, 16'd52247, 16'd22109, 16'd10763, 16'd51951, 16'd29396, 16'd28987, 16'd42337, 16'd7351, 16'd21372});
	test_expansion(128'h36d2a1a2699dd77c45903061d9b046f7, {16'd10728, 16'd10996, 16'd61344, 16'd34413, 16'd21813, 16'd10727, 16'd40213, 16'd3654, 16'd18336, 16'd18723, 16'd19422, 16'd58681, 16'd24738, 16'd40288, 16'd25493, 16'd26408, 16'd50740, 16'd64386, 16'd20290, 16'd17386, 16'd22230, 16'd45231, 16'd37038, 16'd2691, 16'd60260, 16'd59021});
	test_expansion(128'h88a861baac70aa6b2f86fdaf61494443, {16'd49674, 16'd5425, 16'd28702, 16'd31524, 16'd60901, 16'd58892, 16'd36063, 16'd14073, 16'd50006, 16'd28153, 16'd46252, 16'd23683, 16'd25989, 16'd58792, 16'd9247, 16'd39679, 16'd43824, 16'd50978, 16'd31903, 16'd40997, 16'd23388, 16'd15922, 16'd20487, 16'd34443, 16'd16747, 16'd6979});
	test_expansion(128'heb260e0ea7f3768461bd5c2423118999, {16'd12587, 16'd31245, 16'd55331, 16'd17178, 16'd58681, 16'd30636, 16'd3640, 16'd37083, 16'd47823, 16'd24278, 16'd40710, 16'd25535, 16'd29008, 16'd30340, 16'd22937, 16'd39524, 16'd44466, 16'd53992, 16'd24251, 16'd50309, 16'd39580, 16'd30659, 16'd709, 16'd3430, 16'd7347, 16'd44754});
	test_expansion(128'h9dd909fef03c36bf40d574e7002aac51, {16'd4096, 16'd8243, 16'd4342, 16'd13744, 16'd32066, 16'd24404, 16'd58068, 16'd10498, 16'd36453, 16'd15753, 16'd64374, 16'd19297, 16'd8089, 16'd48969, 16'd46886, 16'd19084, 16'd27519, 16'd11082, 16'd51826, 16'd890, 16'd41993, 16'd31918, 16'd54565, 16'd13581, 16'd63724, 16'd55240});
	test_expansion(128'h09090b5975b3e5eab02c4f7b05ab9d88, {16'd42264, 16'd1373, 16'd26863, 16'd25791, 16'd1988, 16'd36312, 16'd1630, 16'd55822, 16'd3613, 16'd3942, 16'd41414, 16'd52107, 16'd18612, 16'd31013, 16'd53567, 16'd27534, 16'd23929, 16'd40827, 16'd49027, 16'd62679, 16'd25001, 16'd15656, 16'd56653, 16'd15808, 16'd47510, 16'd61436});
	test_expansion(128'h4f1b38153e835436ca074ada6392e6b8, {16'd65397, 16'd8711, 16'd10318, 16'd32075, 16'd47627, 16'd24302, 16'd23370, 16'd50211, 16'd29650, 16'd35237, 16'd40583, 16'd63396, 16'd2254, 16'd40029, 16'd6137, 16'd17202, 16'd9911, 16'd31432, 16'd48485, 16'd47948, 16'd8995, 16'd24145, 16'd44034, 16'd30469, 16'd56042, 16'd45677});
	test_expansion(128'h533643de797e5eb08af756eaf1f2ecd1, {16'd37424, 16'd31633, 16'd15117, 16'd25774, 16'd49018, 16'd24949, 16'd11816, 16'd21091, 16'd36854, 16'd19870, 16'd54321, 16'd15930, 16'd1027, 16'd48286, 16'd32821, 16'd47720, 16'd47012, 16'd27928, 16'd3763, 16'd42745, 16'd43484, 16'd8167, 16'd34645, 16'd13067, 16'd58545, 16'd4676});
	test_expansion(128'hefac9242183757e94579194e65a14dc1, {16'd46554, 16'd18892, 16'd55335, 16'd45400, 16'd32294, 16'd28121, 16'd483, 16'd45681, 16'd8352, 16'd9768, 16'd59123, 16'd39483, 16'd52977, 16'd6904, 16'd10864, 16'd40646, 16'd35491, 16'd14983, 16'd19815, 16'd58687, 16'd46777, 16'd39687, 16'd28887, 16'd54472, 16'd18705, 16'd37699});
	test_expansion(128'h9625c37d5e44311ba2f933755514dd8a, {16'd29116, 16'd27054, 16'd12789, 16'd49575, 16'd15558, 16'd9792, 16'd1361, 16'd61994, 16'd22658, 16'd28811, 16'd50021, 16'd58530, 16'd14396, 16'd41824, 16'd42804, 16'd20913, 16'd65282, 16'd7609, 16'd772, 16'd49879, 16'd52792, 16'd37430, 16'd28155, 16'd52844, 16'd31194, 16'd580});
	test_expansion(128'he111e2716a708d2246ac7900c52a5a2f, {16'd34228, 16'd57320, 16'd3855, 16'd40110, 16'd8559, 16'd22802, 16'd42615, 16'd14526, 16'd35386, 16'd29032, 16'd5054, 16'd31569, 16'd22298, 16'd29486, 16'd28371, 16'd33167, 16'd51644, 16'd38177, 16'd21061, 16'd48347, 16'd55591, 16'd44953, 16'd53119, 16'd33357, 16'd36412, 16'd17342});
	test_expansion(128'haad8cc04245227612155560b530e500d, {16'd35778, 16'd7428, 16'd24664, 16'd43042, 16'd61919, 16'd51488, 16'd5697, 16'd22433, 16'd5974, 16'd1283, 16'd27058, 16'd24249, 16'd24737, 16'd5593, 16'd58216, 16'd28906, 16'd56334, 16'd52677, 16'd4827, 16'd59333, 16'd51306, 16'd41137, 16'd24918, 16'd22242, 16'd20878, 16'd27766});
	test_expansion(128'he398ef477ad7fc5efc2fc1a4e118b288, {16'd58600, 16'd49681, 16'd61979, 16'd41885, 16'd56907, 16'd65287, 16'd34832, 16'd28187, 16'd47484, 16'd57999, 16'd63885, 16'd33205, 16'd16978, 16'd10896, 16'd54304, 16'd22162, 16'd44140, 16'd14831, 16'd45157, 16'd12860, 16'd10097, 16'd58733, 16'd5031, 16'd7347, 16'd30681, 16'd35011});
	test_expansion(128'h93e2f7abb669f87659bae6ac9dcfbeba, {16'd16478, 16'd431, 16'd46108, 16'd41057, 16'd63915, 16'd30491, 16'd51931, 16'd43447, 16'd5207, 16'd36038, 16'd65501, 16'd38046, 16'd29355, 16'd54706, 16'd41590, 16'd60037, 16'd6098, 16'd43774, 16'd18883, 16'd46781, 16'd7544, 16'd23320, 16'd16316, 16'd27297, 16'd32528, 16'd7827});
	test_expansion(128'hdacffe294b78e15a9d7fb4f7a992324f, {16'd62101, 16'd53606, 16'd26026, 16'd2163, 16'd14030, 16'd20675, 16'd24897, 16'd40516, 16'd17859, 16'd31173, 16'd43827, 16'd41642, 16'd15529, 16'd5698, 16'd54880, 16'd4254, 16'd62346, 16'd49480, 16'd33696, 16'd50744, 16'd47257, 16'd29229, 16'd45514, 16'd33287, 16'd1375, 16'd30817});
	test_expansion(128'hecc981c333d2e089da658b9e8c9dde6e, {16'd23788, 16'd22275, 16'd71, 16'd873, 16'd4158, 16'd51206, 16'd43761, 16'd14357, 16'd46133, 16'd4638, 16'd47195, 16'd10216, 16'd24287, 16'd4368, 16'd46114, 16'd34355, 16'd25677, 16'd35001, 16'd11980, 16'd32720, 16'd32246, 16'd12702, 16'd19734, 16'd33440, 16'd53953, 16'd46475});
	test_expansion(128'h91f5b51d7d09f0a8d0e13a7d3ad98ca7, {16'd47096, 16'd56197, 16'd62120, 16'd14070, 16'd19173, 16'd53542, 16'd56631, 16'd19451, 16'd24224, 16'd48715, 16'd47369, 16'd53735, 16'd23664, 16'd10352, 16'd40466, 16'd49692, 16'd14833, 16'd37555, 16'd24593, 16'd40330, 16'd38927, 16'd25802, 16'd23420, 16'd52212, 16'd30919, 16'd31026});
	test_expansion(128'h8be3eeea35f6e48dc55eb9e27afbf373, {16'd40386, 16'd30413, 16'd50732, 16'd33108, 16'd2305, 16'd12985, 16'd12053, 16'd21891, 16'd20719, 16'd23832, 16'd26740, 16'd46381, 16'd14223, 16'd5098, 16'd56075, 16'd33192, 16'd16140, 16'd39985, 16'd50367, 16'd46712, 16'd30469, 16'd35652, 16'd25616, 16'd50700, 16'd34178, 16'd54938});
	test_expansion(128'h53c1ed40b4586442bff4deb804b5fb6c, {16'd48600, 16'd9117, 16'd2829, 16'd21171, 16'd7847, 16'd59091, 16'd8403, 16'd2773, 16'd63490, 16'd64695, 16'd19103, 16'd14326, 16'd4977, 16'd18247, 16'd26445, 16'd14767, 16'd29188, 16'd49007, 16'd25219, 16'd62025, 16'd53977, 16'd21030, 16'd11562, 16'd48046, 16'd47704, 16'd40645});
	test_expansion(128'h19b00c4d1162bef4dbc83a9882f7602c, {16'd62604, 16'd31891, 16'd9945, 16'd47568, 16'd8506, 16'd21686, 16'd52135, 16'd33219, 16'd22641, 16'd3903, 16'd6534, 16'd63465, 16'd37181, 16'd15675, 16'd19110, 16'd32196, 16'd26, 16'd13987, 16'd20829, 16'd62459, 16'd51773, 16'd55614, 16'd58763, 16'd43607, 16'd5546, 16'd61184});
	test_expansion(128'h7c284456fcbefd869b29306fb2987096, {16'd58483, 16'd26243, 16'd36414, 16'd18971, 16'd54241, 16'd20437, 16'd32763, 16'd20867, 16'd58185, 16'd1423, 16'd61946, 16'd14749, 16'd15188, 16'd63354, 16'd13432, 16'd60152, 16'd58598, 16'd22083, 16'd33260, 16'd40217, 16'd8062, 16'd54373, 16'd33966, 16'd20146, 16'd56419, 16'd54465});
	test_expansion(128'h93aaf04a9ee2c6b6ffe81871e685443d, {16'd7957, 16'd70, 16'd56554, 16'd19899, 16'd42136, 16'd29870, 16'd11471, 16'd14097, 16'd60472, 16'd40481, 16'd49277, 16'd21598, 16'd3180, 16'd38526, 16'd9395, 16'd36080, 16'd22909, 16'd4226, 16'd39742, 16'd22569, 16'd62679, 16'd15163, 16'd8091, 16'd46532, 16'd63154, 16'd49320});
	test_expansion(128'hf939be0189b947d2e5a969fb00062d21, {16'd46877, 16'd26747, 16'd51198, 16'd45274, 16'd61340, 16'd18078, 16'd24550, 16'd65525, 16'd44312, 16'd33875, 16'd53076, 16'd2222, 16'd21365, 16'd59275, 16'd21462, 16'd35284, 16'd4075, 16'd44530, 16'd53012, 16'd40012, 16'd15158, 16'd58781, 16'd55046, 16'd625, 16'd23093, 16'd53289});
	test_expansion(128'h799e19eb893e355534bbbb631a2dc4ac, {16'd5718, 16'd39782, 16'd58212, 16'd49868, 16'd45775, 16'd15481, 16'd53696, 16'd53339, 16'd14079, 16'd59509, 16'd43725, 16'd27416, 16'd64643, 16'd51733, 16'd9652, 16'd59703, 16'd55738, 16'd33620, 16'd30667, 16'd15688, 16'd56356, 16'd48480, 16'd1874, 16'd27700, 16'd63026, 16'd22137});
	test_expansion(128'hb5cc005f99ec5aeaaf68a00a11674d80, {16'd39192, 16'd55596, 16'd5341, 16'd35672, 16'd12006, 16'd27618, 16'd10633, 16'd10180, 16'd48486, 16'd15304, 16'd31821, 16'd22671, 16'd36136, 16'd52338, 16'd3042, 16'd54258, 16'd35770, 16'd31991, 16'd1776, 16'd6, 16'd44259, 16'd13911, 16'd28168, 16'd58689, 16'd34310, 16'd35450});
	test_expansion(128'hb6afd0b93606d3cb7c49a09bbd67ea62, {16'd20109, 16'd43448, 16'd32692, 16'd20846, 16'd11456, 16'd18119, 16'd994, 16'd6060, 16'd59792, 16'd29657, 16'd51348, 16'd27412, 16'd26729, 16'd37939, 16'd6910, 16'd44363, 16'd42759, 16'd31060, 16'd25050, 16'd62008, 16'd63753, 16'd4178, 16'd25146, 16'd34598, 16'd52981, 16'd27410});
	test_expansion(128'h0e72cb543435fb209ca2bdc55ae55d0f, {16'd52002, 16'd59519, 16'd5937, 16'd10928, 16'd13069, 16'd45630, 16'd28735, 16'd40409, 16'd17907, 16'd13098, 16'd32095, 16'd61268, 16'd58939, 16'd47586, 16'd20195, 16'd14154, 16'd29680, 16'd18453, 16'd15526, 16'd31947, 16'd60818, 16'd13155, 16'd64947, 16'd15199, 16'd27710, 16'd18100});
	test_expansion(128'h8a699767aca679c8a720e53bfb2e15f7, {16'd48198, 16'd14490, 16'd61005, 16'd57006, 16'd20313, 16'd36, 16'd59743, 16'd51045, 16'd58438, 16'd54938, 16'd17069, 16'd11246, 16'd47206, 16'd35403, 16'd58306, 16'd56966, 16'd1974, 16'd34314, 16'd63752, 16'd31517, 16'd9185, 16'd46361, 16'd42232, 16'd27575, 16'd14084, 16'd20823});
	test_expansion(128'haf01714c358a413cf13143378a3bea27, {16'd23519, 16'd52956, 16'd43835, 16'd63800, 16'd22397, 16'd43463, 16'd63765, 16'd56516, 16'd40023, 16'd40201, 16'd47749, 16'd2299, 16'd47197, 16'd61508, 16'd48301, 16'd50288, 16'd4264, 16'd14064, 16'd1584, 16'd20688, 16'd3894, 16'd23842, 16'd15042, 16'd56870, 16'd53705, 16'd41562});
	test_expansion(128'h38165c8a165243da50693bf35691b44a, {16'd41623, 16'd13549, 16'd60684, 16'd305, 16'd13192, 16'd19371, 16'd52264, 16'd42965, 16'd44381, 16'd57004, 16'd42317, 16'd1110, 16'd5407, 16'd13653, 16'd30190, 16'd16033, 16'd53358, 16'd12554, 16'd11028, 16'd16422, 16'd45380, 16'd40022, 16'd29212, 16'd14809, 16'd25620, 16'd1350});
	test_expansion(128'hb7b2e4753738a4d10dce5f6b47144c84, {16'd30597, 16'd6760, 16'd56716, 16'd2991, 16'd33710, 16'd62817, 16'd58061, 16'd53507, 16'd1218, 16'd51195, 16'd57954, 16'd56492, 16'd32418, 16'd27311, 16'd29756, 16'd41797, 16'd4193, 16'd24017, 16'd40165, 16'd5959, 16'd9386, 16'd36686, 16'd48266, 16'd5944, 16'd57684, 16'd28597});
	test_expansion(128'h8a636d1058aded038cc198e689fd2d8c, {16'd63317, 16'd37595, 16'd30554, 16'd30561, 16'd53666, 16'd32862, 16'd48327, 16'd36055, 16'd1446, 16'd36397, 16'd6546, 16'd60645, 16'd21642, 16'd30476, 16'd6298, 16'd40316, 16'd13455, 16'd8545, 16'd49261, 16'd31491, 16'd56408, 16'd43275, 16'd48541, 16'd49670, 16'd42618, 16'd44951});
	test_expansion(128'hdb6ad882530a3a71deb17714dc8f4f4c, {16'd30018, 16'd45106, 16'd45584, 16'd55344, 16'd63501, 16'd58417, 16'd2329, 16'd25682, 16'd43807, 16'd18048, 16'd26399, 16'd15785, 16'd62653, 16'd47900, 16'd29614, 16'd59228, 16'd46364, 16'd2409, 16'd11154, 16'd38513, 16'd56655, 16'd47369, 16'd44851, 16'd54818, 16'd22591, 16'd10770});
	test_expansion(128'h66d95a95f09df04a6017bf491a413f03, {16'd37099, 16'd57947, 16'd17193, 16'd46190, 16'd5926, 16'd14716, 16'd43609, 16'd719, 16'd41038, 16'd32528, 16'd39880, 16'd24233, 16'd707, 16'd12074, 16'd40707, 16'd61962, 16'd28783, 16'd19205, 16'd51328, 16'd17030, 16'd39623, 16'd18185, 16'd61264, 16'd48227, 16'd13325, 16'd5940});
	test_expansion(128'h94b9cd821f1c1a28404003fdcbc9605c, {16'd35449, 16'd31664, 16'd22121, 16'd4615, 16'd59476, 16'd1266, 16'd1572, 16'd52430, 16'd58318, 16'd4133, 16'd10205, 16'd245, 16'd60109, 16'd15913, 16'd2091, 16'd41438, 16'd36292, 16'd13125, 16'd25049, 16'd42422, 16'd9859, 16'd30123, 16'd32920, 16'd51869, 16'd46802, 16'd58807});
	test_expansion(128'hdaadbe877dad5ae35c67621423b95358, {16'd30624, 16'd50631, 16'd42344, 16'd44321, 16'd53235, 16'd39394, 16'd54946, 16'd12924, 16'd50238, 16'd55846, 16'd25515, 16'd45832, 16'd26087, 16'd16013, 16'd43714, 16'd4211, 16'd18238, 16'd29940, 16'd14884, 16'd40730, 16'd14927, 16'd34745, 16'd40956, 16'd57158, 16'd13560, 16'd35809});
	test_expansion(128'hdab5ec4a3ebb3d6bf0c2a24151b60831, {16'd28699, 16'd45235, 16'd15037, 16'd44654, 16'd43539, 16'd29612, 16'd60778, 16'd608, 16'd36949, 16'd16057, 16'd20395, 16'd11790, 16'd46914, 16'd56981, 16'd19749, 16'd55245, 16'd14578, 16'd63291, 16'd9513, 16'd34820, 16'd57170, 16'd50995, 16'd1195, 16'd58372, 16'd11108, 16'd651});
	test_expansion(128'h4600629b7f4a3c0ccdd17ac338a07d40, {16'd33814, 16'd4164, 16'd48752, 16'd61914, 16'd11484, 16'd17133, 16'd48487, 16'd22541, 16'd44910, 16'd52118, 16'd42572, 16'd25324, 16'd52065, 16'd48631, 16'd55021, 16'd12639, 16'd34194, 16'd27052, 16'd19563, 16'd47022, 16'd4053, 16'd16619, 16'd44097, 16'd54490, 16'd4007, 16'd44475});
	test_expansion(128'hf5b72c02098955e66ce9de8c29a2fa56, {16'd9688, 16'd39514, 16'd56403, 16'd2334, 16'd1057, 16'd11687, 16'd42522, 16'd35126, 16'd474, 16'd35746, 16'd18162, 16'd20766, 16'd7467, 16'd50440, 16'd24391, 16'd10568, 16'd39325, 16'd6529, 16'd26624, 16'd32920, 16'd3527, 16'd17130, 16'd44798, 16'd15094, 16'd31098, 16'd53490});
	test_expansion(128'hda35461a7befd42afa2bf1318dca6dc8, {16'd47617, 16'd64241, 16'd50045, 16'd55776, 16'd15414, 16'd2246, 16'd35557, 16'd38641, 16'd12782, 16'd6233, 16'd55978, 16'd28347, 16'd37762, 16'd8008, 16'd24959, 16'd41661, 16'd23783, 16'd32555, 16'd22570, 16'd49938, 16'd37782, 16'd49553, 16'd33603, 16'd28025, 16'd26551, 16'd2983});
	test_expansion(128'h4f7805406c3ed224c2f5580cab1a1656, {16'd34280, 16'd26388, 16'd15730, 16'd47812, 16'd18387, 16'd3917, 16'd40955, 16'd2520, 16'd24769, 16'd61341, 16'd58535, 16'd58610, 16'd15998, 16'd16215, 16'd40371, 16'd61470, 16'd29404, 16'd54235, 16'd59850, 16'd25940, 16'd33833, 16'd19872, 16'd63268, 16'd45548, 16'd41318, 16'd48257});
	test_expansion(128'h13a27ec563234f8ecab722785303ed8f, {16'd37904, 16'd14200, 16'd12269, 16'd37699, 16'd43734, 16'd13423, 16'd1962, 16'd3953, 16'd37123, 16'd43129, 16'd64124, 16'd50303, 16'd14394, 16'd21388, 16'd40572, 16'd31280, 16'd6364, 16'd6814, 16'd33016, 16'd10769, 16'd5039, 16'd23947, 16'd41307, 16'd22835, 16'd19181, 16'd38266});
	test_expansion(128'h4c7b7d1a8ccacc9919f1a42e8ac588a5, {16'd28703, 16'd9173, 16'd57169, 16'd56050, 16'd60632, 16'd30761, 16'd34418, 16'd36779, 16'd41635, 16'd28032, 16'd56347, 16'd31109, 16'd28749, 16'd60619, 16'd46404, 16'd33381, 16'd56288, 16'd25298, 16'd27909, 16'd43842, 16'd27109, 16'd41501, 16'd34925, 16'd25947, 16'd2141, 16'd9508});
	test_expansion(128'h65563e0a6511eb16c1c0ecd3e2ea2521, {16'd45914, 16'd60529, 16'd32369, 16'd20446, 16'd57726, 16'd43713, 16'd5890, 16'd54826, 16'd45486, 16'd24988, 16'd41641, 16'd4336, 16'd31950, 16'd2381, 16'd36989, 16'd46963, 16'd8488, 16'd7254, 16'd43970, 16'd37305, 16'd4593, 16'd41346, 16'd41023, 16'd50465, 16'd18335, 16'd11388});
	test_expansion(128'hc99db4ccad5a07af6275faeb563f3ce8, {16'd52883, 16'd45523, 16'd4379, 16'd24044, 16'd28761, 16'd64524, 16'd34509, 16'd25014, 16'd12234, 16'd23191, 16'd31732, 16'd31874, 16'd50765, 16'd60498, 16'd2378, 16'd7086, 16'd707, 16'd59551, 16'd3894, 16'd21143, 16'd23023, 16'd60919, 16'd46571, 16'd46482, 16'd53927, 16'd12528});
	test_expansion(128'ha81ed5b51eac57df17172b3bba361d65, {16'd51312, 16'd65293, 16'd44213, 16'd5941, 16'd11993, 16'd26107, 16'd29308, 16'd43741, 16'd9172, 16'd33101, 16'd54117, 16'd62718, 16'd40213, 16'd30332, 16'd32173, 16'd16791, 16'd62915, 16'd18480, 16'd29971, 16'd8397, 16'd61083, 16'd5528, 16'd39085, 16'd53142, 16'd18493, 16'd31060});
	test_expansion(128'hcab6d6f9e115a9bb9d02eafdc10acb54, {16'd43605, 16'd35331, 16'd21779, 16'd349, 16'd12587, 16'd26234, 16'd37844, 16'd15933, 16'd12212, 16'd222, 16'd51778, 16'd5306, 16'd16101, 16'd57429, 16'd23162, 16'd50993, 16'd6997, 16'd11968, 16'd9834, 16'd56199, 16'd44697, 16'd28349, 16'd38783, 16'd45299, 16'd63022, 16'd34749});
	test_expansion(128'h3d81a6a472a8af46674757bf93cd517d, {16'd62639, 16'd34986, 16'd20183, 16'd50575, 16'd39370, 16'd27116, 16'd37131, 16'd38295, 16'd7750, 16'd21845, 16'd3618, 16'd62642, 16'd48603, 16'd54803, 16'd17103, 16'd44885, 16'd64947, 16'd165, 16'd6103, 16'd12992, 16'd3659, 16'd17487, 16'd64749, 16'd7710, 16'd28114, 16'd42339});
	test_expansion(128'hc14b901980e641cefddb77f03fe20488, {16'd46366, 16'd9747, 16'd25237, 16'd17002, 16'd663, 16'd45947, 16'd56292, 16'd40026, 16'd34259, 16'd37961, 16'd23369, 16'd19204, 16'd15214, 16'd20555, 16'd62109, 16'd29365, 16'd25536, 16'd17042, 16'd19451, 16'd51868, 16'd29680, 16'd24424, 16'd35950, 16'd39258, 16'd5036, 16'd15775});
	test_expansion(128'hfaed2efa360e828f607a6d83dfea4901, {16'd55167, 16'd36842, 16'd53602, 16'd58577, 16'd5617, 16'd8035, 16'd42572, 16'd3511, 16'd65048, 16'd52505, 16'd51127, 16'd61284, 16'd43035, 16'd24538, 16'd18938, 16'd49612, 16'd7907, 16'd12991, 16'd6312, 16'd4470, 16'd63783, 16'd43693, 16'd40292, 16'd52830, 16'd10668, 16'd17176});
	test_expansion(128'h584007b564b549986c9aea57216b2c3e, {16'd40473, 16'd62372, 16'd13036, 16'd59388, 16'd43573, 16'd12695, 16'd14136, 16'd61633, 16'd40379, 16'd4398, 16'd3265, 16'd12670, 16'd49044, 16'd4279, 16'd14687, 16'd64405, 16'd14533, 16'd11160, 16'd8128, 16'd22832, 16'd56564, 16'd34907, 16'd55597, 16'd22672, 16'd35852, 16'd25135});
	test_expansion(128'h3b19b12a2650e30558f2c576aaabe710, {16'd57585, 16'd4599, 16'd93, 16'd24638, 16'd6589, 16'd27655, 16'd15801, 16'd33257, 16'd28938, 16'd57489, 16'd58667, 16'd41382, 16'd2911, 16'd11513, 16'd11663, 16'd56510, 16'd30939, 16'd4419, 16'd52844, 16'd44736, 16'd36520, 16'd57107, 16'd33390, 16'd29365, 16'd7557, 16'd8111});
	test_expansion(128'heac4eac8bf5ed4538ac9034e4b5375c4, {16'd19845, 16'd27578, 16'd57634, 16'd28535, 16'd11489, 16'd45067, 16'd9386, 16'd3801, 16'd28873, 16'd63829, 16'd58706, 16'd46129, 16'd27288, 16'd40865, 16'd65030, 16'd62477, 16'd36271, 16'd16620, 16'd23346, 16'd33166, 16'd9013, 16'd14521, 16'd44804, 16'd22609, 16'd37074, 16'd55921});
	test_expansion(128'hf7c0790e1a2f798934e66590ba91cbba, {16'd37582, 16'd11414, 16'd24891, 16'd20325, 16'd51981, 16'd39463, 16'd50068, 16'd48173, 16'd38972, 16'd11425, 16'd60511, 16'd18473, 16'd21754, 16'd40967, 16'd39598, 16'd40816, 16'd21886, 16'd45045, 16'd45648, 16'd8439, 16'd41290, 16'd2583, 16'd31874, 16'd20317, 16'd2847, 16'd14148});
	test_expansion(128'h88caedc6781d10fe60878106b5d3614c, {16'd28129, 16'd24494, 16'd53038, 16'd13325, 16'd62502, 16'd40103, 16'd25482, 16'd16304, 16'd31620, 16'd21670, 16'd64774, 16'd47265, 16'd43217, 16'd34636, 16'd39986, 16'd54845, 16'd20119, 16'd9729, 16'd63824, 16'd60802, 16'd59483, 16'd2766, 16'd28112, 16'd35875, 16'd46391, 16'd10089});
	test_expansion(128'h85a83205a9876a665697a45d8a78c315, {16'd63392, 16'd54793, 16'd31469, 16'd31588, 16'd31692, 16'd13775, 16'd47678, 16'd27026, 16'd19510, 16'd55127, 16'd5010, 16'd35771, 16'd4454, 16'd43909, 16'd33457, 16'd54277, 16'd54316, 16'd23528, 16'd35349, 16'd37042, 16'd44332, 16'd39167, 16'd1420, 16'd57617, 16'd51874, 16'd53213});
	test_expansion(128'h7b61b0d85f8c0268be54e333b9173b7b, {16'd44607, 16'd48607, 16'd61359, 16'd6335, 16'd15964, 16'd56371, 16'd41965, 16'd43367, 16'd3311, 16'd29309, 16'd14226, 16'd39566, 16'd18036, 16'd53357, 16'd33581, 16'd21811, 16'd45071, 16'd16108, 16'd6396, 16'd62025, 16'd37559, 16'd22106, 16'd42583, 16'd31610, 16'd63298, 16'd52801});
	test_expansion(128'h2d0e4e2295fa67b4ec655bf68cb56a9d, {16'd18146, 16'd28635, 16'd48805, 16'd40210, 16'd18773, 16'd12373, 16'd5839, 16'd20948, 16'd23038, 16'd22347, 16'd16564, 16'd40023, 16'd48805, 16'd17697, 16'd29224, 16'd44096, 16'd65042, 16'd35661, 16'd25752, 16'd17553, 16'd22568, 16'd48088, 16'd56327, 16'd58248, 16'd24737, 16'd47891});
	test_expansion(128'h4ab8d6fdfe2a058f3f3053edef388006, {16'd32750, 16'd31908, 16'd30403, 16'd37641, 16'd5950, 16'd27448, 16'd45096, 16'd57012, 16'd37817, 16'd43542, 16'd57581, 16'd31997, 16'd31045, 16'd33141, 16'd12301, 16'd37322, 16'd33878, 16'd20136, 16'd47851, 16'd57035, 16'd24207, 16'd4312, 16'd44772, 16'd29321, 16'd11824, 16'd20814});
	test_expansion(128'hbf2efa272d2164e36258505d7f4d5b0d, {16'd7755, 16'd52519, 16'd3622, 16'd10062, 16'd8668, 16'd42561, 16'd9759, 16'd58412, 16'd12309, 16'd37890, 16'd24791, 16'd3367, 16'd18962, 16'd41206, 16'd60167, 16'd33061, 16'd54014, 16'd46677, 16'd33777, 16'd58353, 16'd17469, 16'd18592, 16'd59958, 16'd8505, 16'd26235, 16'd55849});
	test_expansion(128'h163afbe22f357e749ca4cc91c5072ad4, {16'd28251, 16'd46295, 16'd41391, 16'd46797, 16'd8819, 16'd9428, 16'd12983, 16'd28361, 16'd21143, 16'd53786, 16'd11801, 16'd1158, 16'd44697, 16'd42374, 16'd36499, 16'd2753, 16'd36120, 16'd5166, 16'd47750, 16'd40848, 16'd12992, 16'd57367, 16'd55412, 16'd25104, 16'd16127, 16'd3350});
	test_expansion(128'h79f5d0b452b020cf46c9110ae625b83e, {16'd46850, 16'd38339, 16'd57831, 16'd11992, 16'd9149, 16'd64606, 16'd64036, 16'd21549, 16'd26906, 16'd65252, 16'd6289, 16'd63713, 16'd7780, 16'd62004, 16'd8225, 16'd15082, 16'd8240, 16'd38195, 16'd61712, 16'd32372, 16'd37132, 16'd54447, 16'd13459, 16'd61342, 16'd11481, 16'd20571});
	test_expansion(128'h62de226456ee436871d49e7eecb8a5a3, {16'd35662, 16'd759, 16'd29083, 16'd64314, 16'd12061, 16'd7691, 16'd29349, 16'd50680, 16'd13325, 16'd61580, 16'd64860, 16'd47788, 16'd55437, 16'd34062, 16'd62012, 16'd47544, 16'd22030, 16'd35458, 16'd51554, 16'd15786, 16'd57383, 16'd64192, 16'd16212, 16'd59105, 16'd59211, 16'd7797});
	test_expansion(128'ha9482049b121574a23d884df24c7bc12, {16'd1800, 16'd13860, 16'd59811, 16'd39219, 16'd25023, 16'd9428, 16'd57515, 16'd29236, 16'd10023, 16'd50831, 16'd58534, 16'd13341, 16'd49431, 16'd36129, 16'd61927, 16'd60016, 16'd26295, 16'd59496, 16'd28254, 16'd12575, 16'd50933, 16'd4612, 16'd8129, 16'd56506, 16'd49401, 16'd20487});
	test_expansion(128'h62737c1ecbc26f17c912d8e5274e1088, {16'd26704, 16'd9944, 16'd27426, 16'd2932, 16'd59185, 16'd28502, 16'd57484, 16'd49839, 16'd37949, 16'd26197, 16'd34397, 16'd24815, 16'd8436, 16'd29753, 16'd36984, 16'd4800, 16'd56200, 16'd11024, 16'd49558, 16'd52025, 16'd5676, 16'd27957, 16'd32262, 16'd34762, 16'd63671, 16'd57504});
	test_expansion(128'hfe78303022d127387c0d659bd69a8617, {16'd15622, 16'd29640, 16'd31485, 16'd2151, 16'd49888, 16'd43315, 16'd40366, 16'd26623, 16'd50249, 16'd57737, 16'd15037, 16'd8690, 16'd3099, 16'd10276, 16'd21420, 16'd40654, 16'd38696, 16'd62273, 16'd5480, 16'd35131, 16'd57170, 16'd60901, 16'd43116, 16'd8293, 16'd59471, 16'd64024});
	test_expansion(128'hc723d0341e0b86bddfb255d93c09c3eb, {16'd60130, 16'd2930, 16'd38811, 16'd38833, 16'd51746, 16'd61929, 16'd62264, 16'd1708, 16'd42341, 16'd65197, 16'd62475, 16'd6468, 16'd20070, 16'd52787, 16'd43439, 16'd19962, 16'd9260, 16'd63066, 16'd56043, 16'd21468, 16'd21068, 16'd34723, 16'd12511, 16'd46156, 16'd54965, 16'd42054});
	test_expansion(128'hdbb31d34889973f9a019a533206d7de2, {16'd8525, 16'd24760, 16'd64909, 16'd40715, 16'd48222, 16'd23338, 16'd56998, 16'd26254, 16'd29069, 16'd13085, 16'd32170, 16'd44179, 16'd36744, 16'd39631, 16'd50156, 16'd26047, 16'd27871, 16'd44945, 16'd12031, 16'd55861, 16'd57394, 16'd50757, 16'd27625, 16'd31116, 16'd3858, 16'd64053});
	test_expansion(128'hd4b4edbc32397005a5322b9ba4ff5598, {16'd4809, 16'd4706, 16'd9389, 16'd5680, 16'd57218, 16'd16798, 16'd15033, 16'd5792, 16'd56182, 16'd20348, 16'd3767, 16'd63674, 16'd45000, 16'd56820, 16'd15444, 16'd46407, 16'd6031, 16'd9020, 16'd40136, 16'd1243, 16'd47715, 16'd40912, 16'd55154, 16'd31779, 16'd55292, 16'd47521});
	test_expansion(128'hd46da062c0a41bd24b6a1bef34290303, {16'd60167, 16'd12953, 16'd55531, 16'd34466, 16'd52726, 16'd32587, 16'd26247, 16'd9089, 16'd25834, 16'd31208, 16'd20949, 16'd4731, 16'd35200, 16'd21950, 16'd41463, 16'd4594, 16'd46325, 16'd9887, 16'd59909, 16'd51239, 16'd9564, 16'd9977, 16'd63237, 16'd45962, 16'd12977, 16'd13609});
	test_expansion(128'hd06b3689e404bd97520244683771692b, {16'd26054, 16'd7630, 16'd48323, 16'd11002, 16'd7505, 16'd7984, 16'd18552, 16'd36093, 16'd48707, 16'd12963, 16'd19985, 16'd25756, 16'd35437, 16'd25213, 16'd5372, 16'd25741, 16'd26736, 16'd24675, 16'd62397, 16'd27195, 16'd11648, 16'd59703, 16'd37588, 16'd5664, 16'd41759, 16'd51294});
	test_expansion(128'hc231a962eb5677bb6def5dc723d33565, {16'd573, 16'd56684, 16'd60975, 16'd44009, 16'd61718, 16'd17965, 16'd20176, 16'd21888, 16'd39385, 16'd11171, 16'd30673, 16'd13865, 16'd15732, 16'd62115, 16'd25525, 16'd17437, 16'd33297, 16'd17691, 16'd4361, 16'd3417, 16'd47374, 16'd15534, 16'd61654, 16'd28547, 16'd40654, 16'd11757});
	test_expansion(128'h49289c0dbcc157f5f265c2d69d2cb923, {16'd16313, 16'd4017, 16'd28673, 16'd20561, 16'd55368, 16'd43953, 16'd34182, 16'd62024, 16'd61467, 16'd5853, 16'd46797, 16'd43511, 16'd20153, 16'd45481, 16'd18835, 16'd17466, 16'd46914, 16'd21157, 16'd34223, 16'd24615, 16'd36643, 16'd15870, 16'd26488, 16'd5743, 16'd46017, 16'd36770});
	test_expansion(128'h6a10a856e3f73f6cce9ab24cfab0c060, {16'd8385, 16'd31294, 16'd42153, 16'd22628, 16'd59268, 16'd4963, 16'd23075, 16'd11219, 16'd53627, 16'd9, 16'd48586, 16'd30145, 16'd47865, 16'd36064, 16'd34005, 16'd37130, 16'd64090, 16'd54398, 16'd41582, 16'd50887, 16'd21066, 16'd55364, 16'd43954, 16'd51751, 16'd60686, 16'd49398});
	test_expansion(128'hae12f3cd1afdbbd233da4dbc646004f5, {16'd39537, 16'd2038, 16'd8049, 16'd37412, 16'd7936, 16'd21666, 16'd53406, 16'd64944, 16'd40515, 16'd55586, 16'd452, 16'd36716, 16'd51559, 16'd52941, 16'd52160, 16'd51154, 16'd59773, 16'd43212, 16'd58840, 16'd42517, 16'd53558, 16'd60861, 16'd94, 16'd14096, 16'd12139, 16'd19530});
	test_expansion(128'h03a3ba614f6241c52a826c4311c43aec, {16'd51627, 16'd31198, 16'd22565, 16'd28680, 16'd15698, 16'd44595, 16'd61135, 16'd56906, 16'd62594, 16'd37572, 16'd47784, 16'd63595, 16'd51416, 16'd17331, 16'd9168, 16'd11569, 16'd15729, 16'd57863, 16'd59031, 16'd44371, 16'd40935, 16'd52819, 16'd10477, 16'd42584, 16'd3046, 16'd29067});
	test_expansion(128'h7f78b48e8afe4baff49faa01ceec34e6, {16'd55694, 16'd19448, 16'd27883, 16'd61425, 16'd45343, 16'd18713, 16'd57212, 16'd27165, 16'd43745, 16'd33838, 16'd59980, 16'd59060, 16'd28480, 16'd61641, 16'd56257, 16'd38453, 16'd49103, 16'd43786, 16'd2637, 16'd36080, 16'd54026, 16'd34499, 16'd59308, 16'd24973, 16'd30650, 16'd51913});
	test_expansion(128'h8ea8219a32ccef2b65bdb3c5d32e00a7, {16'd56674, 16'd58718, 16'd29127, 16'd65108, 16'd56639, 16'd24024, 16'd1383, 16'd42436, 16'd20225, 16'd65519, 16'd58079, 16'd64731, 16'd824, 16'd32150, 16'd41657, 16'd23374, 16'd51443, 16'd1721, 16'd63856, 16'd56914, 16'd34038, 16'd33330, 16'd13101, 16'd29761, 16'd2866, 16'd13798});
	test_expansion(128'h16a06dc1ba9f1100251745c4a1db54b7, {16'd15045, 16'd45062, 16'd13738, 16'd28833, 16'd23380, 16'd17943, 16'd31809, 16'd45580, 16'd6815, 16'd28530, 16'd5275, 16'd43431, 16'd35009, 16'd44634, 16'd3332, 16'd26156, 16'd10378, 16'd40533, 16'd2404, 16'd57596, 16'd22340, 16'd30941, 16'd36018, 16'd59538, 16'd43416, 16'd54442});
	test_expansion(128'h02c455e944a4cde1430ea1b44c081c62, {16'd3118, 16'd43690, 16'd38524, 16'd57240, 16'd59067, 16'd4971, 16'd48239, 16'd55358, 16'd26436, 16'd13937, 16'd55140, 16'd11325, 16'd51184, 16'd54178, 16'd59316, 16'd49825, 16'd19506, 16'd19695, 16'd16319, 16'd44279, 16'd41143, 16'd49000, 16'd46001, 16'd1918, 16'd2320, 16'd27392});
	test_expansion(128'habc8dafbe96d3ce317548bad21cd555e, {16'd55798, 16'd39314, 16'd63870, 16'd931, 16'd37701, 16'd34728, 16'd23330, 16'd1614, 16'd52840, 16'd289, 16'd50277, 16'd48840, 16'd60357, 16'd32656, 16'd59923, 16'd63375, 16'd5320, 16'd31273, 16'd25971, 16'd41936, 16'd53433, 16'd34099, 16'd60367, 16'd49825, 16'd52231, 16'd31646});
	test_expansion(128'h82f01824062c5e77091df73c340592f6, {16'd54679, 16'd8295, 16'd23984, 16'd8584, 16'd50926, 16'd8729, 16'd26692, 16'd55313, 16'd48452, 16'd11473, 16'd55720, 16'd12922, 16'd35810, 16'd8784, 16'd53196, 16'd12595, 16'd55958, 16'd54900, 16'd15519, 16'd29867, 16'd19802, 16'd15161, 16'd8914, 16'd59342, 16'd33923, 16'd52571});
	test_expansion(128'hd6b156257dbdf85353d69e66832ab473, {16'd39721, 16'd12743, 16'd63633, 16'd16554, 16'd46722, 16'd60367, 16'd24889, 16'd26526, 16'd22618, 16'd7515, 16'd61049, 16'd38106, 16'd37406, 16'd15396, 16'd46489, 16'd64285, 16'd36930, 16'd22788, 16'd64227, 16'd42273, 16'd47928, 16'd43813, 16'd8594, 16'd38810, 16'd3460, 16'd26132});
	test_expansion(128'he9e073331f6e1955520b2d54a5296f5f, {16'd32189, 16'd8869, 16'd50777, 16'd50510, 16'd44959, 16'd49554, 16'd23851, 16'd22739, 16'd23087, 16'd64754, 16'd24203, 16'd60883, 16'd62596, 16'd44028, 16'd6399, 16'd44915, 16'd25688, 16'd25522, 16'd31535, 16'd63580, 16'd5984, 16'd44716, 16'd46497, 16'd45374, 16'd37195, 16'd38475});
	test_expansion(128'hbe3560fb4492ea85a51ec8c4831b1f15, {16'd3358, 16'd5784, 16'd52682, 16'd2291, 16'd15291, 16'd36664, 16'd4571, 16'd58848, 16'd51522, 16'd60063, 16'd40437, 16'd49541, 16'd219, 16'd28088, 16'd25904, 16'd9063, 16'd43277, 16'd23809, 16'd37124, 16'd50605, 16'd8750, 16'd29626, 16'd15941, 16'd132, 16'd17023, 16'd32153});
	test_expansion(128'hd476c5c4c672039ded4897f627d13f36, {16'd41609, 16'd29849, 16'd59618, 16'd25287, 16'd58859, 16'd4426, 16'd44911, 16'd36878, 16'd44560, 16'd2141, 16'd5887, 16'd53700, 16'd24397, 16'd25718, 16'd55755, 16'd11036, 16'd26307, 16'd10795, 16'd20658, 16'd50238, 16'd7988, 16'd33685, 16'd45994, 16'd22159, 16'd13529, 16'd11149});
	test_expansion(128'h2c7e0019a1834983b6e23a4c4812a3d7, {16'd52603, 16'd12344, 16'd36781, 16'd2757, 16'd52516, 16'd48520, 16'd17216, 16'd43995, 16'd57042, 16'd54059, 16'd41552, 16'd16053, 16'd6584, 16'd19695, 16'd14624, 16'd54613, 16'd35098, 16'd61537, 16'd43783, 16'd58350, 16'd3316, 16'd41534, 16'd9406, 16'd21309, 16'd15756, 16'd4344});
	test_expansion(128'h452d0e3b32588ef930a82577ad7462c2, {16'd23366, 16'd13105, 16'd5662, 16'd2964, 16'd49403, 16'd21990, 16'd39887, 16'd33906, 16'd21531, 16'd12585, 16'd21565, 16'd52535, 16'd61577, 16'd9947, 16'd16230, 16'd1972, 16'd30494, 16'd55812, 16'd53828, 16'd54850, 16'd25044, 16'd17895, 16'd1248, 16'd22244, 16'd37125, 16'd41059});
	test_expansion(128'h00d172b12c573e7cb0c52279e5e9c36a, {16'd56988, 16'd62278, 16'd58562, 16'd44507, 16'd36275, 16'd47505, 16'd49259, 16'd40913, 16'd54688, 16'd27482, 16'd40544, 16'd53670, 16'd31435, 16'd32511, 16'd31284, 16'd8545, 16'd63128, 16'd34761, 16'd16117, 16'd46479, 16'd18922, 16'd25574, 16'd48246, 16'd64614, 16'd62882, 16'd7927});
	test_expansion(128'he33ad9410be1c5ef9cdc953404b94744, {16'd37413, 16'd13539, 16'd44588, 16'd30279, 16'd3378, 16'd40522, 16'd19372, 16'd3015, 16'd38428, 16'd40667, 16'd264, 16'd27520, 16'd50221, 16'd30384, 16'd7092, 16'd275, 16'd15105, 16'd1397, 16'd31744, 16'd61188, 16'd56485, 16'd19063, 16'd16414, 16'd50793, 16'd37632, 16'd8587});
	test_expansion(128'hb7562fba913af9dddbf68e9d38711d5b, {16'd34294, 16'd32089, 16'd20592, 16'd21582, 16'd38077, 16'd27862, 16'd8488, 16'd59170, 16'd10808, 16'd12070, 16'd36304, 16'd55155, 16'd51443, 16'd5142, 16'd2817, 16'd61285, 16'd40021, 16'd58302, 16'd62504, 16'd33225, 16'd55891, 16'd16466, 16'd39603, 16'd50730, 16'd30809, 16'd60106});
	test_expansion(128'h82435087b81cc2374d6e08603175149d, {16'd15903, 16'd46618, 16'd50237, 16'd15500, 16'd17794, 16'd60058, 16'd60810, 16'd21966, 16'd7707, 16'd50627, 16'd43495, 16'd55795, 16'd56573, 16'd8584, 16'd23252, 16'd11103, 16'd50332, 16'd24305, 16'd4510, 16'd10593, 16'd50645, 16'd64293, 16'd2919, 16'd46214, 16'd29754, 16'd30369});
	test_expansion(128'ha5d82b791691262d01f340730c869f27, {16'd13638, 16'd29152, 16'd65391, 16'd8193, 16'd36956, 16'd50212, 16'd45101, 16'd15666, 16'd10, 16'd60822, 16'd23420, 16'd3711, 16'd29329, 16'd27615, 16'd4914, 16'd8413, 16'd37959, 16'd32693, 16'd34900, 16'd27281, 16'd2791, 16'd17084, 16'd9257, 16'd26165, 16'd53052, 16'd54424});
	test_expansion(128'hb5b37b73bdbb42be955b49de11b3addc, {16'd1011, 16'd23418, 16'd62783, 16'd55943, 16'd27547, 16'd6924, 16'd43547, 16'd14228, 16'd11640, 16'd60017, 16'd31238, 16'd30199, 16'd17590, 16'd42200, 16'd50089, 16'd37711, 16'd63516, 16'd40138, 16'd47855, 16'd31974, 16'd57290, 16'd20329, 16'd22430, 16'd32082, 16'd59917, 16'd25579});
	test_expansion(128'h0dd340b549db463e3694c39246843e6f, {16'd60036, 16'd48531, 16'd50223, 16'd57719, 16'd41867, 16'd46585, 16'd11894, 16'd25984, 16'd64865, 16'd8916, 16'd17263, 16'd60590, 16'd2619, 16'd48269, 16'd23728, 16'd8489, 16'd33086, 16'd53861, 16'd29447, 16'd26253, 16'd63687, 16'd53423, 16'd51466, 16'd9662, 16'd61776, 16'd43252});
	test_expansion(128'h11551c41ce6d8e82e93e127258dab29f, {16'd49356, 16'd20762, 16'd63115, 16'd1800, 16'd14495, 16'd31107, 16'd54034, 16'd59360, 16'd6409, 16'd50225, 16'd38886, 16'd3199, 16'd28197, 16'd46565, 16'd26556, 16'd24453, 16'd38347, 16'd28265, 16'd34361, 16'd55165, 16'd53450, 16'd48519, 16'd20888, 16'd17388, 16'd17054, 16'd26117});
	test_expansion(128'h128dc2827bb567ddfc338b07a8ababc4, {16'd39229, 16'd43623, 16'd16201, 16'd33530, 16'd7665, 16'd31049, 16'd52013, 16'd15522, 16'd544, 16'd38662, 16'd23565, 16'd61106, 16'd26926, 16'd57567, 16'd55092, 16'd36255, 16'd61556, 16'd35856, 16'd20372, 16'd35335, 16'd2910, 16'd11485, 16'd8993, 16'd12755, 16'd20736, 16'd23086});
	test_expansion(128'hbcdf98538665a6cbf48718a5a11e1c9d, {16'd1187, 16'd62135, 16'd9758, 16'd36314, 16'd13473, 16'd28291, 16'd35058, 16'd7493, 16'd44807, 16'd15970, 16'd23872, 16'd21999, 16'd19786, 16'd49666, 16'd19713, 16'd12738, 16'd55032, 16'd37706, 16'd38021, 16'd30080, 16'd61001, 16'd49534, 16'd23302, 16'd31662, 16'd57536, 16'd33335});
	test_expansion(128'h4599a77771261ae74cd6f6d6b98b8134, {16'd58270, 16'd55150, 16'd42992, 16'd38712, 16'd7120, 16'd17404, 16'd65303, 16'd12363, 16'd31117, 16'd29499, 16'd33662, 16'd23357, 16'd1169, 16'd29777, 16'd8932, 16'd59936, 16'd10543, 16'd65102, 16'd31725, 16'd55398, 16'd47085, 16'd17662, 16'd27033, 16'd33835, 16'd23691, 16'd13010});
	test_expansion(128'h6cd43dc18f6f697500ef811136bafdb0, {16'd2575, 16'd29155, 16'd36589, 16'd27056, 16'd24336, 16'd31873, 16'd36541, 16'd33545, 16'd52216, 16'd13582, 16'd2544, 16'd15033, 16'd2429, 16'd13910, 16'd34371, 16'd7978, 16'd14523, 16'd18221, 16'd64673, 16'd56842, 16'd29787, 16'd55774, 16'd41781, 16'd8379, 16'd635, 16'd65158});
	test_expansion(128'h6d28c9816180bdaf140266a08a0d78d0, {16'd62949, 16'd12416, 16'd62394, 16'd38364, 16'd15456, 16'd46486, 16'd45497, 16'd8000, 16'd19551, 16'd42386, 16'd4089, 16'd51075, 16'd9390, 16'd50449, 16'd57884, 16'd30810, 16'd3234, 16'd16905, 16'd6408, 16'd6002, 16'd33014, 16'd33461, 16'd20187, 16'd9779, 16'd49078, 16'd59449});
	test_expansion(128'hc13b81f768017e93822eb83447b076dc, {16'd36387, 16'd49808, 16'd30927, 16'd9900, 16'd46864, 16'd521, 16'd60549, 16'd58707, 16'd47222, 16'd45453, 16'd27244, 16'd30643, 16'd60343, 16'd40877, 16'd64835, 16'd31385, 16'd14326, 16'd30895, 16'd26552, 16'd51942, 16'd30202, 16'd38209, 16'd58413, 16'd49156, 16'd4768, 16'd53864});
	test_expansion(128'h4956f29330b75a44bdee0d40a628a998, {16'd18456, 16'd30132, 16'd14460, 16'd49811, 16'd14483, 16'd60435, 16'd17258, 16'd25202, 16'd35209, 16'd18630, 16'd12128, 16'd32482, 16'd41480, 16'd47207, 16'd62017, 16'd44618, 16'd2643, 16'd12202, 16'd7888, 16'd48138, 16'd32504, 16'd53360, 16'd14903, 16'd7693, 16'd34569, 16'd19018});
	test_expansion(128'hd287976f41c0b2d44aef68daab07de77, {16'd12363, 16'd46573, 16'd63323, 16'd15871, 16'd12778, 16'd16551, 16'd39162, 16'd9067, 16'd20847, 16'd22326, 16'd64784, 16'd30190, 16'd61077, 16'd39767, 16'd28288, 16'd32853, 16'd33788, 16'd55801, 16'd44692, 16'd35797, 16'd48965, 16'd28742, 16'd56389, 16'd33996, 16'd13250, 16'd21267});
	test_expansion(128'he68f69165e9b4b7731e2286b22387a17, {16'd37314, 16'd33613, 16'd54287, 16'd26409, 16'd16461, 16'd6202, 16'd30494, 16'd21801, 16'd10047, 16'd18528, 16'd33076, 16'd3479, 16'd29851, 16'd43040, 16'd7825, 16'd49802, 16'd33275, 16'd46690, 16'd777, 16'd37967, 16'd57609, 16'd12580, 16'd10226, 16'd20793, 16'd44770, 16'd47527});
	test_expansion(128'hb15b1902e9df2eb61b06184420aea9e9, {16'd10574, 16'd15994, 16'd59308, 16'd20977, 16'd63379, 16'd43223, 16'd54563, 16'd36468, 16'd60534, 16'd54981, 16'd60240, 16'd23460, 16'd57064, 16'd19239, 16'd64376, 16'd8512, 16'd8038, 16'd45695, 16'd41820, 16'd10146, 16'd42904, 16'd6642, 16'd25096, 16'd10622, 16'd7097, 16'd5737});
	test_expansion(128'hf6d679b251f1e4849192b4a8deffc1b9, {16'd5512, 16'd36990, 16'd16768, 16'd65014, 16'd38888, 16'd45989, 16'd1170, 16'd23939, 16'd1503, 16'd57206, 16'd35897, 16'd34344, 16'd29974, 16'd26203, 16'd11820, 16'd50466, 16'd44014, 16'd28938, 16'd27366, 16'd49184, 16'd2658, 16'd43158, 16'd43372, 16'd36059, 16'd46960, 16'd3494});
	test_expansion(128'hb25b98a9071201202d148d60e51946aa, {16'd20041, 16'd35909, 16'd50185, 16'd39012, 16'd43081, 16'd31777, 16'd25650, 16'd7062, 16'd60434, 16'd32336, 16'd58852, 16'd16449, 16'd4748, 16'd20889, 16'd32919, 16'd28236, 16'd24285, 16'd64585, 16'd29215, 16'd27553, 16'd64141, 16'd41048, 16'd42258, 16'd31629, 16'd33166, 16'd46661});
	test_expansion(128'hb39a59f1af9072d3d4d899be2fb010ef, {16'd49673, 16'd57924, 16'd29657, 16'd59247, 16'd38826, 16'd23308, 16'd53499, 16'd38299, 16'd20293, 16'd19088, 16'd61516, 16'd26846, 16'd8322, 16'd60623, 16'd5055, 16'd10822, 16'd30049, 16'd39292, 16'd15674, 16'd17203, 16'd29746, 16'd374, 16'd21227, 16'd32517, 16'd42925, 16'd8643});
	test_expansion(128'h0b74345cf1da4d6244413f028e1dca6e, {16'd64517, 16'd52539, 16'd42786, 16'd648, 16'd42332, 16'd2456, 16'd35887, 16'd26118, 16'd23025, 16'd19467, 16'd2362, 16'd22875, 16'd6219, 16'd57410, 16'd52568, 16'd19174, 16'd62964, 16'd42473, 16'd17915, 16'd33620, 16'd42862, 16'd11773, 16'd30693, 16'd18348, 16'd16839, 16'd7919});
	test_expansion(128'h686a5bf3789ae292f0821479399475a9, {16'd8176, 16'd42047, 16'd35638, 16'd39654, 16'd149, 16'd24457, 16'd64902, 16'd34021, 16'd39159, 16'd36297, 16'd43365, 16'd36074, 16'd17239, 16'd63364, 16'd5939, 16'd15816, 16'd50636, 16'd23945, 16'd46679, 16'd23423, 16'd48933, 16'd21153, 16'd35496, 16'd64136, 16'd41835, 16'd4955});
	test_expansion(128'haafcb2db107216d645d8f40ab3e86ab3, {16'd50091, 16'd61824, 16'd3530, 16'd22463, 16'd22168, 16'd12002, 16'd60351, 16'd4231, 16'd38055, 16'd5203, 16'd36514, 16'd27239, 16'd48987, 16'd52575, 16'd10620, 16'd43278, 16'd45663, 16'd4105, 16'd9910, 16'd56726, 16'd44499, 16'd26206, 16'd58310, 16'd37468, 16'd30837, 16'd48175});
	test_expansion(128'h0d8a2e790332dcb5d95a2017c7902aae, {16'd24219, 16'd14527, 16'd53884, 16'd40120, 16'd23175, 16'd32006, 16'd54641, 16'd42527, 16'd28907, 16'd25188, 16'd51173, 16'd60589, 16'd13308, 16'd20889, 16'd23815, 16'd26599, 16'd45843, 16'd47218, 16'd47369, 16'd29979, 16'd52410, 16'd24646, 16'd2008, 16'd52972, 16'd51164, 16'd5848});
	test_expansion(128'h7c15821a6a39575cb6b6a87fe04028e0, {16'd42483, 16'd11444, 16'd32280, 16'd34844, 16'd48016, 16'd58168, 16'd45014, 16'd50837, 16'd55940, 16'd4465, 16'd60820, 16'd42263, 16'd59923, 16'd13516, 16'd47274, 16'd31627, 16'd64202, 16'd20483, 16'd54664, 16'd61055, 16'd24650, 16'd19556, 16'd11801, 16'd47423, 16'd30380, 16'd55832});
	test_expansion(128'h4320d4a23eadf8860498693424c54bca, {16'd9759, 16'd10890, 16'd21063, 16'd55573, 16'd50200, 16'd64450, 16'd61189, 16'd51604, 16'd12786, 16'd55568, 16'd38087, 16'd41320, 16'd48330, 16'd10542, 16'd770, 16'd37923, 16'd25517, 16'd46751, 16'd56265, 16'd43244, 16'd22026, 16'd20765, 16'd40730, 16'd12702, 16'd50521, 16'd18651});
	test_expansion(128'h495056cb8121bb605ec063ea884d80ce, {16'd38751, 16'd64997, 16'd33527, 16'd12642, 16'd20024, 16'd30008, 16'd33992, 16'd56728, 16'd35702, 16'd30616, 16'd32689, 16'd4836, 16'd3562, 16'd59146, 16'd4976, 16'd29768, 16'd63455, 16'd9450, 16'd18190, 16'd46400, 16'd19257, 16'd45142, 16'd4538, 16'd12355, 16'd60429, 16'd41267});
	test_expansion(128'h190e3f5bcb364e5a56dafe428b9307fa, {16'd56512, 16'd14886, 16'd14228, 16'd29609, 16'd39662, 16'd35588, 16'd16396, 16'd20299, 16'd40732, 16'd53867, 16'd49175, 16'd28246, 16'd5993, 16'd64494, 16'd7750, 16'd1221, 16'd48186, 16'd3148, 16'd14421, 16'd18959, 16'd3328, 16'd50475, 16'd16062, 16'd53133, 16'd63214, 16'd2307});
	test_expansion(128'h20ccec0cb65766b74329a52b638f56aa, {16'd25763, 16'd31848, 16'd25637, 16'd17586, 16'd35519, 16'd53394, 16'd1678, 16'd14300, 16'd37022, 16'd63813, 16'd7810, 16'd28850, 16'd33484, 16'd54108, 16'd51725, 16'd22765, 16'd32624, 16'd40540, 16'd61624, 16'd47348, 16'd34093, 16'd24598, 16'd33957, 16'd8351, 16'd27485, 16'd13236});
	test_expansion(128'h55fe32954c8eedf4ecd210006e9b1e2f, {16'd41138, 16'd36520, 16'd18665, 16'd54310, 16'd14013, 16'd15948, 16'd32224, 16'd59444, 16'd17531, 16'd2184, 16'd36153, 16'd34151, 16'd61236, 16'd1757, 16'd50718, 16'd53557, 16'd20919, 16'd57672, 16'd47897, 16'd58226, 16'd24805, 16'd40506, 16'd11436, 16'd52855, 16'd54207, 16'd44587});
	test_expansion(128'h7a033c717f0733f1dcda96a9828d5ea0, {16'd6315, 16'd45527, 16'd12914, 16'd18613, 16'd13792, 16'd39422, 16'd49913, 16'd20838, 16'd48523, 16'd6780, 16'd54434, 16'd19999, 16'd21802, 16'd7099, 16'd62613, 16'd54009, 16'd56915, 16'd55269, 16'd16336, 16'd47066, 16'd29214, 16'd42650, 16'd52778, 16'd23451, 16'd43751, 16'd43533});
	test_expansion(128'hde0268c522032ed76188133d59fe128b, {16'd54132, 16'd50476, 16'd11960, 16'd16530, 16'd27081, 16'd22397, 16'd9207, 16'd32133, 16'd50318, 16'd33732, 16'd261, 16'd7868, 16'd46161, 16'd61231, 16'd28357, 16'd45591, 16'd50710, 16'd41305, 16'd61210, 16'd32824, 16'd37672, 16'd55050, 16'd58612, 16'd17967, 16'd16491, 16'd42769});
	test_expansion(128'h0261074ea87262db93252e9b3c17e7de, {16'd51185, 16'd32764, 16'd40889, 16'd11058, 16'd47622, 16'd46565, 16'd12824, 16'd29496, 16'd32547, 16'd13216, 16'd40033, 16'd46624, 16'd4334, 16'd33090, 16'd26142, 16'd46137, 16'd49062, 16'd41196, 16'd52471, 16'd28480, 16'd28319, 16'd57304, 16'd46623, 16'd54822, 16'd26457, 16'd60738});
	test_expansion(128'h1abaa9f11505ad34e6a17dcb240285c3, {16'd16216, 16'd45947, 16'd28309, 16'd45971, 16'd16, 16'd17621, 16'd15725, 16'd21218, 16'd44827, 16'd52402, 16'd23190, 16'd53079, 16'd10483, 16'd24531, 16'd39548, 16'd42869, 16'd3469, 16'd52575, 16'd52757, 16'd54416, 16'd484, 16'd48474, 16'd668, 16'd24234, 16'd27391, 16'd31203});
	test_expansion(128'hd2c1df47292f1a4cb67e1069e0791e30, {16'd22129, 16'd58533, 16'd63889, 16'd26812, 16'd14052, 16'd17416, 16'd35333, 16'd32946, 16'd37945, 16'd36334, 16'd21131, 16'd4979, 16'd46049, 16'd23708, 16'd400, 16'd13267, 16'd40650, 16'd3600, 16'd2898, 16'd2341, 16'd42102, 16'd59750, 16'd39210, 16'd34495, 16'd14372, 16'd54295});
	test_expansion(128'hda6f2f9df621fdf447a466123a678e66, {16'd16997, 16'd61174, 16'd36607, 16'd10603, 16'd42281, 16'd33052, 16'd15439, 16'd23034, 16'd46802, 16'd33369, 16'd34916, 16'd57200, 16'd4321, 16'd27724, 16'd57608, 16'd31318, 16'd41930, 16'd7161, 16'd21924, 16'd11733, 16'd57645, 16'd51529, 16'd12547, 16'd843, 16'd27381, 16'd26910});
	test_expansion(128'h4e60abbe475ca0d0760ff0a9c21f0c3b, {16'd46792, 16'd35826, 16'd39317, 16'd49579, 16'd32328, 16'd46793, 16'd34492, 16'd15490, 16'd61866, 16'd49597, 16'd33398, 16'd14725, 16'd28386, 16'd59654, 16'd35643, 16'd26701, 16'd33639, 16'd22376, 16'd36875, 16'd62201, 16'd23923, 16'd65425, 16'd16882, 16'd56570, 16'd59383, 16'd40775});
	test_expansion(128'h258d3827ffe2dc12388e573ae2e32d68, {16'd25453, 16'd18522, 16'd42716, 16'd21505, 16'd8198, 16'd65424, 16'd37548, 16'd54719, 16'd24592, 16'd35486, 16'd20342, 16'd51714, 16'd49726, 16'd60345, 16'd57304, 16'd21406, 16'd61809, 16'd8854, 16'd38627, 16'd1692, 16'd10137, 16'd35115, 16'd9858, 16'd8545, 16'd49383, 16'd61952});
	test_expansion(128'h572b6946c09f00e46bd20ed9c517d6d7, {16'd56878, 16'd51959, 16'd1678, 16'd10250, 16'd19733, 16'd43437, 16'd25130, 16'd26351, 16'd63651, 16'd12370, 16'd28401, 16'd21454, 16'd26570, 16'd56631, 16'd47390, 16'd33383, 16'd41130, 16'd60002, 16'd28278, 16'd52934, 16'd48682, 16'd25423, 16'd51028, 16'd40559, 16'd50654, 16'd39602});
	test_expansion(128'h58ee9140734376886b37f3219e653ebc, {16'd12826, 16'd57152, 16'd7683, 16'd17329, 16'd3198, 16'd51837, 16'd45447, 16'd32458, 16'd11024, 16'd63742, 16'd21320, 16'd922, 16'd22258, 16'd50191, 16'd48902, 16'd9264, 16'd57145, 16'd50943, 16'd38630, 16'd10439, 16'd49824, 16'd14503, 16'd12268, 16'd5915, 16'd56885, 16'd55253});
	test_expansion(128'h6b983a6341055132dfc78d36a54432e7, {16'd44922, 16'd21849, 16'd48301, 16'd19139, 16'd2494, 16'd29831, 16'd7992, 16'd30003, 16'd12786, 16'd12549, 16'd29813, 16'd13269, 16'd15598, 16'd43856, 16'd4148, 16'd56116, 16'd28407, 16'd5178, 16'd15598, 16'd38155, 16'd26061, 16'd6891, 16'd64510, 16'd4063, 16'd17704, 16'd55861});
	test_expansion(128'hbe4435446d9ec43b55649d5cc73bccc1, {16'd1515, 16'd63930, 16'd23610, 16'd26910, 16'd61366, 16'd24147, 16'd53184, 16'd9277, 16'd52463, 16'd44804, 16'd63055, 16'd8039, 16'd63227, 16'd51900, 16'd65210, 16'd11013, 16'd8118, 16'd615, 16'd27627, 16'd36430, 16'd30353, 16'd8365, 16'd45302, 16'd32765, 16'd33180, 16'd25618});
	test_expansion(128'h8ac0b3b8314aa9dc20906640f73737d9, {16'd38543, 16'd2743, 16'd62871, 16'd60664, 16'd1838, 16'd19692, 16'd18119, 16'd7588, 16'd64550, 16'd9388, 16'd62442, 16'd19701, 16'd56889, 16'd17658, 16'd34206, 16'd53661, 16'd21725, 16'd42454, 16'd20736, 16'd36566, 16'd53308, 16'd9011, 16'd64020, 16'd49695, 16'd44289, 16'd37996});
	test_expansion(128'he0cd9303216ceee967a60977f692ee94, {16'd17184, 16'd44220, 16'd32742, 16'd35318, 16'd17391, 16'd21092, 16'd64885, 16'd30077, 16'd39103, 16'd27402, 16'd15398, 16'd15455, 16'd42785, 16'd31190, 16'd59115, 16'd44300, 16'd63130, 16'd46041, 16'd5053, 16'd47524, 16'd30822, 16'd16737, 16'd58744, 16'd16415, 16'd51116, 16'd15102});
	test_expansion(128'hc74b43c7f5530609ddc07b9dbb8b8fec, {16'd34734, 16'd12620, 16'd21822, 16'd10339, 16'd51901, 16'd8177, 16'd22644, 16'd2912, 16'd33643, 16'd54166, 16'd4585, 16'd4468, 16'd13624, 16'd41320, 16'd58750, 16'd14291, 16'd32366, 16'd42437, 16'd35756, 16'd32602, 16'd36516, 16'd32950, 16'd52498, 16'd47312, 16'd15763, 16'd46476});
	test_expansion(128'h499adc31b3214cda8dc55fac9c402811, {16'd40648, 16'd62609, 16'd42757, 16'd46836, 16'd63284, 16'd33555, 16'd15634, 16'd61800, 16'd26686, 16'd57745, 16'd5484, 16'd33193, 16'd60535, 16'd34679, 16'd6024, 16'd64561, 16'd43409, 16'd56804, 16'd57959, 16'd16396, 16'd12519, 16'd13199, 16'd50649, 16'd28853, 16'd13522, 16'd51163});
	test_expansion(128'hf980ab77b57e3b770523bc8916e53247, {16'd41559, 16'd42386, 16'd27910, 16'd56434, 16'd52686, 16'd22778, 16'd26307, 16'd1789, 16'd50184, 16'd34747, 16'd7219, 16'd52776, 16'd39457, 16'd36510, 16'd11402, 16'd10198, 16'd13330, 16'd63024, 16'd44957, 16'd20882, 16'd60911, 16'd53351, 16'd33618, 16'd36445, 16'd38058, 16'd43003});
	test_expansion(128'hfdc17cd2336747a6b3bfc3d1c84dae37, {16'd4298, 16'd38406, 16'd47196, 16'd25097, 16'd4185, 16'd17771, 16'd33531, 16'd11175, 16'd32768, 16'd18621, 16'd23953, 16'd36964, 16'd13113, 16'd22657, 16'd62529, 16'd56861, 16'd18432, 16'd4697, 16'd49587, 16'd25245, 16'd20566, 16'd39275, 16'd47209, 16'd17148, 16'd38176, 16'd54922});
	test_expansion(128'h73f10b34e88e7eab5fb6bb7d39feaac2, {16'd41818, 16'd35021, 16'd62824, 16'd45641, 16'd33308, 16'd63124, 16'd655, 16'd49641, 16'd8966, 16'd5784, 16'd32692, 16'd19090, 16'd43618, 16'd50849, 16'd6945, 16'd61873, 16'd14281, 16'd58114, 16'd16780, 16'd50310, 16'd10541, 16'd28543, 16'd22314, 16'd43263, 16'd48675, 16'd45067});
	test_expansion(128'h7bcff058a5ba91458764470314c252e0, {16'd52345, 16'd20620, 16'd16142, 16'd50376, 16'd50342, 16'd19337, 16'd8944, 16'd13110, 16'd1334, 16'd35935, 16'd25139, 16'd62145, 16'd19805, 16'd17126, 16'd24300, 16'd28787, 16'd40206, 16'd61582, 16'd11206, 16'd48873, 16'd65146, 16'd12301, 16'd13135, 16'd51701, 16'd29170, 16'd38841});
	test_expansion(128'h094dcaedc6085890ac2f756910475986, {16'd47134, 16'd52558, 16'd30309, 16'd36013, 16'd7578, 16'd52442, 16'd46125, 16'd10662, 16'd40407, 16'd61703, 16'd45945, 16'd453, 16'd4133, 16'd5718, 16'd56214, 16'd44860, 16'd57598, 16'd55883, 16'd35086, 16'd38373, 16'd27556, 16'd29203, 16'd63337, 16'd21541, 16'd23254, 16'd7025});
	test_expansion(128'he91154efef4d5dccb12c04092576d43b, {16'd45197, 16'd42896, 16'd7369, 16'd10961, 16'd53279, 16'd57633, 16'd56602, 16'd62609, 16'd7320, 16'd2461, 16'd46244, 16'd9859, 16'd4657, 16'd19155, 16'd48079, 16'd16183, 16'd22022, 16'd33893, 16'd50553, 16'd35557, 16'd3385, 16'd58739, 16'd27309, 16'd22115, 16'd21241, 16'd62330});
	test_expansion(128'h3d3c44451622299c6029f33135448985, {16'd63637, 16'd18179, 16'd31406, 16'd27106, 16'd49619, 16'd16766, 16'd21871, 16'd49191, 16'd37491, 16'd64837, 16'd45821, 16'd38896, 16'd22757, 16'd31879, 16'd3389, 16'd51527, 16'd10723, 16'd57144, 16'd21554, 16'd45151, 16'd56354, 16'd10229, 16'd51267, 16'd8765, 16'd61698, 16'd55965});
	test_expansion(128'h0f4ecd0d6b429821fd8e3bfccc42eb9a, {16'd51515, 16'd32415, 16'd17361, 16'd22042, 16'd32673, 16'd23866, 16'd39528, 16'd45019, 16'd34263, 16'd29208, 16'd20551, 16'd26057, 16'd12687, 16'd21027, 16'd55896, 16'd30803, 16'd57424, 16'd10484, 16'd41360, 16'd37055, 16'd53411, 16'd4192, 16'd25890, 16'd27752, 16'd9279, 16'd23801});
	test_expansion(128'h2d0f5bd05750fc5d1724592061945d61, {16'd24404, 16'd55601, 16'd40013, 16'd40119, 16'd55877, 16'd41860, 16'd23615, 16'd26934, 16'd48793, 16'd18055, 16'd18824, 16'd65250, 16'd14962, 16'd38253, 16'd17140, 16'd48911, 16'd5086, 16'd9464, 16'd11667, 16'd19956, 16'd2521, 16'd7588, 16'd39694, 16'd21417, 16'd14507, 16'd22806});
	test_expansion(128'h63aa9329f86656ad2e0e0079e0181976, {16'd3616, 16'd46660, 16'd20271, 16'd9571, 16'd16680, 16'd52514, 16'd26725, 16'd42279, 16'd19683, 16'd19750, 16'd31362, 16'd21608, 16'd64593, 16'd64895, 16'd37005, 16'd29052, 16'd9211, 16'd27966, 16'd19922, 16'd38786, 16'd59791, 16'd64638, 16'd6486, 16'd2660, 16'd55679, 16'd57318});
	test_expansion(128'h9da31d45250803d1d03ae821cfca1947, {16'd56206, 16'd14220, 16'd58383, 16'd25017, 16'd22818, 16'd35585, 16'd39561, 16'd25245, 16'd8300, 16'd47875, 16'd55534, 16'd15101, 16'd40859, 16'd38457, 16'd47641, 16'd3272, 16'd48465, 16'd42417, 16'd42913, 16'd8132, 16'd38376, 16'd19018, 16'd65185, 16'd52127, 16'd20908, 16'd38816});
	test_expansion(128'h2022bb66d2f36a695a0f1166fb3d7e70, {16'd26341, 16'd16255, 16'd58130, 16'd59537, 16'd6260, 16'd44256, 16'd45845, 16'd62906, 16'd63351, 16'd9188, 16'd41663, 16'd24287, 16'd1629, 16'd48113, 16'd1725, 16'd35936, 16'd47146, 16'd2619, 16'd59753, 16'd32891, 16'd49782, 16'd38708, 16'd53489, 16'd9490, 16'd33668, 16'd4206});
	test_expansion(128'h4a3a524566f848eaedb8c4e08e2419f9, {16'd63429, 16'd51354, 16'd47776, 16'd42239, 16'd8508, 16'd39865, 16'd44868, 16'd37751, 16'd17449, 16'd12365, 16'd8829, 16'd29497, 16'd32091, 16'd59090, 16'd24829, 16'd36952, 16'd43452, 16'd14789, 16'd58015, 16'd36926, 16'd35411, 16'd12210, 16'd18220, 16'd16937, 16'd23404, 16'd16638});
	test_expansion(128'h45394f56950612f46246a5ca2d2cf81e, {16'd23629, 16'd61005, 16'd2364, 16'd6293, 16'd63298, 16'd60568, 16'd35986, 16'd32925, 16'd9455, 16'd63250, 16'd45233, 16'd46387, 16'd14937, 16'd64478, 16'd5319, 16'd32439, 16'd33270, 16'd51772, 16'd25159, 16'd8057, 16'd22205, 16'd35236, 16'd51127, 16'd35934, 16'd51942, 16'd11770});
	test_expansion(128'hd7dfb9f8869508d93a8bca287d30587b, {16'd39041, 16'd8857, 16'd46262, 16'd50356, 16'd22403, 16'd17730, 16'd32085, 16'd24888, 16'd21501, 16'd29073, 16'd17794, 16'd26639, 16'd54043, 16'd33627, 16'd465, 16'd41795, 16'd65400, 16'd46189, 16'd56568, 16'd36481, 16'd7172, 16'd5389, 16'd56448, 16'd2769, 16'd18046, 16'd31301});
	test_expansion(128'h2dc3a241af508fcc7fbf79eeaeda06ee, {16'd8832, 16'd27324, 16'd63182, 16'd18033, 16'd42636, 16'd10882, 16'd25397, 16'd216, 16'd61103, 16'd3242, 16'd11701, 16'd39404, 16'd32635, 16'd28890, 16'd40226, 16'd32297, 16'd16881, 16'd42296, 16'd33565, 16'd10189, 16'd37080, 16'd32323, 16'd7693, 16'd22469, 16'd23189, 16'd48579});
	test_expansion(128'ha8842c2ed7d330217eabf6ce94717996, {16'd13797, 16'd6477, 16'd5724, 16'd25378, 16'd11923, 16'd33316, 16'd10239, 16'd47644, 16'd39562, 16'd14650, 16'd64442, 16'd35873, 16'd15936, 16'd26807, 16'd1737, 16'd510, 16'd15759, 16'd15785, 16'd32921, 16'd32691, 16'd867, 16'd54379, 16'd40975, 16'd15332, 16'd5442, 16'd25147});
	test_expansion(128'hff38fd4977691ade691816170fe477b0, {16'd18840, 16'd21618, 16'd1479, 16'd26529, 16'd45731, 16'd11518, 16'd10081, 16'd18175, 16'd45829, 16'd51012, 16'd43457, 16'd64136, 16'd34026, 16'd57617, 16'd1510, 16'd23223, 16'd57, 16'd30593, 16'd55561, 16'd43855, 16'd8658, 16'd60678, 16'd37261, 16'd42864, 16'd5979, 16'd29148});
	test_expansion(128'h77eba9dbbac61dbe4d0ca2a711590478, {16'd56400, 16'd52400, 16'd14053, 16'd12689, 16'd47281, 16'd29528, 16'd33788, 16'd21313, 16'd1413, 16'd7252, 16'd6163, 16'd11717, 16'd10573, 16'd45357, 16'd31710, 16'd9063, 16'd53365, 16'd58217, 16'd53150, 16'd46485, 16'd23661, 16'd53134, 16'd37734, 16'd545, 16'd5617, 16'd65469});
	test_expansion(128'hed475b790f549e04f9e9ca2295d4898d, {16'd52388, 16'd7606, 16'd41952, 16'd16829, 16'd55388, 16'd31876, 16'd14470, 16'd35721, 16'd62178, 16'd22451, 16'd61751, 16'd19860, 16'd30339, 16'd52109, 16'd18259, 16'd25125, 16'd44863, 16'd653, 16'd41535, 16'd15945, 16'd18324, 16'd21013, 16'd33130, 16'd29164, 16'd42636, 16'd38107});
	test_expansion(128'h4acc52e6b44ec68352a16c6a120a6776, {16'd23760, 16'd21675, 16'd15888, 16'd36854, 16'd62847, 16'd37512, 16'd24976, 16'd4709, 16'd41535, 16'd40194, 16'd40559, 16'd20542, 16'd41027, 16'd4169, 16'd55948, 16'd41674, 16'd55113, 16'd64236, 16'd56511, 16'd54576, 16'd12488, 16'd62090, 16'd52124, 16'd23851, 16'd11279, 16'd37175});
	test_expansion(128'hbaf5dd6c83ba5da213d242015acacd32, {16'd42337, 16'd17613, 16'd39214, 16'd35031, 16'd29664, 16'd43474, 16'd17401, 16'd26349, 16'd50596, 16'd18728, 16'd35433, 16'd13967, 16'd48580, 16'd52381, 16'd42939, 16'd13259, 16'd44874, 16'd8114, 16'd3763, 16'd47705, 16'd42526, 16'd26875, 16'd53423, 16'd4484, 16'd41862, 16'd38704});
	test_expansion(128'h12c7f861de780727a5256af09607edef, {16'd39452, 16'd25506, 16'd4297, 16'd21063, 16'd23545, 16'd63360, 16'd25993, 16'd11604, 16'd21265, 16'd6453, 16'd61725, 16'd24844, 16'd55005, 16'd40943, 16'd28676, 16'd28595, 16'd11930, 16'd25752, 16'd38789, 16'd48454, 16'd16201, 16'd33913, 16'd26194, 16'd45218, 16'd16500, 16'd63811});
	test_expansion(128'he514e67aa5115beee0204d51642f1375, {16'd24605, 16'd32912, 16'd6490, 16'd53199, 16'd3471, 16'd31377, 16'd16926, 16'd15014, 16'd19968, 16'd23889, 16'd65422, 16'd50793, 16'd44066, 16'd21449, 16'd6183, 16'd20229, 16'd37920, 16'd31725, 16'd37901, 16'd64643, 16'd29747, 16'd25295, 16'd64468, 16'd2949, 16'd52222, 16'd5555});
	test_expansion(128'hd83e4b511c32d6121dd152f59317d5f0, {16'd908, 16'd21104, 16'd54328, 16'd38103, 16'd50764, 16'd41638, 16'd24440, 16'd17604, 16'd23887, 16'd12223, 16'd2000, 16'd1858, 16'd4977, 16'd41497, 16'd1160, 16'd966, 16'd57973, 16'd14736, 16'd46577, 16'd13066, 16'd42965, 16'd28457, 16'd43000, 16'd39604, 16'd48328, 16'd26646});
	test_expansion(128'h3d5aa39433abfa6abe5c8e8bd1d15b4a, {16'd5305, 16'd31300, 16'd42421, 16'd12975, 16'd41283, 16'd57404, 16'd2579, 16'd31744, 16'd18840, 16'd27844, 16'd55310, 16'd55487, 16'd44742, 16'd37089, 16'd8599, 16'd23085, 16'd8036, 16'd62422, 16'd49664, 16'd46004, 16'd46176, 16'd24634, 16'd31702, 16'd55980, 16'd42496, 16'd2081});
	test_expansion(128'h7de56d1725ab119def9088f7818d83a9, {16'd5071, 16'd14531, 16'd59052, 16'd46446, 16'd34330, 16'd47065, 16'd32425, 16'd60332, 16'd41858, 16'd44906, 16'd11399, 16'd29782, 16'd2503, 16'd3033, 16'd42418, 16'd35207, 16'd54876, 16'd12938, 16'd13799, 16'd29740, 16'd47259, 16'd2964, 16'd31522, 16'd63599, 16'd40142, 16'd58103});
	test_expansion(128'h194d9538a57e86d4ab870ae30847a147, {16'd49650, 16'd27979, 16'd63600, 16'd26792, 16'd53510, 16'd56238, 16'd31151, 16'd51796, 16'd47917, 16'd27009, 16'd27473, 16'd39030, 16'd26619, 16'd29435, 16'd31819, 16'd55080, 16'd34008, 16'd33214, 16'd44045, 16'd962, 16'd21749, 16'd40857, 16'd19799, 16'd35761, 16'd61411, 16'd4345});
	test_expansion(128'hc3f5445c024250f99a997609dc0d08f0, {16'd51093, 16'd60479, 16'd2145, 16'd40884, 16'd16715, 16'd4558, 16'd18029, 16'd24408, 16'd32183, 16'd34017, 16'd56889, 16'd26152, 16'd35204, 16'd26799, 16'd37986, 16'd39848, 16'd53320, 16'd57632, 16'd34219, 16'd9459, 16'd54917, 16'd39717, 16'd44155, 16'd29930, 16'd32328, 16'd65094});
	test_expansion(128'hb57df04181bf7829e140574232d35b64, {16'd18961, 16'd30435, 16'd28895, 16'd14208, 16'd15875, 16'd56243, 16'd59503, 16'd57893, 16'd1231, 16'd3547, 16'd34538, 16'd64457, 16'd46216, 16'd23509, 16'd48297, 16'd16033, 16'd30466, 16'd6308, 16'd15275, 16'd5364, 16'd6224, 16'd60414, 16'd3192, 16'd30111, 16'd37710, 16'd51371});
	test_expansion(128'hb3689578b2b53acebd08b356670c3319, {16'd39189, 16'd65270, 16'd38875, 16'd4765, 16'd58921, 16'd27779, 16'd45189, 16'd2835, 16'd28855, 16'd36296, 16'd12445, 16'd58783, 16'd6627, 16'd30273, 16'd21515, 16'd21818, 16'd50497, 16'd4535, 16'd8762, 16'd15436, 16'd64125, 16'd26102, 16'd22076, 16'd58817, 16'd52858, 16'd28597});
	test_expansion(128'h8d2f9271b3a71f19e090770594d4d5fe, {16'd41561, 16'd46602, 16'd62381, 16'd42580, 16'd1661, 16'd16159, 16'd39853, 16'd55148, 16'd30533, 16'd60759, 16'd41563, 16'd13924, 16'd52409, 16'd41010, 16'd59187, 16'd32600, 16'd56526, 16'd57500, 16'd36066, 16'd10082, 16'd4189, 16'd61464, 16'd27846, 16'd45254, 16'd11158, 16'd39579});
	test_expansion(128'ha0b769cb923dd81970356658d886a963, {16'd57606, 16'd20075, 16'd3257, 16'd62494, 16'd27904, 16'd1551, 16'd60735, 16'd35018, 16'd45275, 16'd14134, 16'd20372, 16'd55431, 16'd21423, 16'd1101, 16'd17544, 16'd28185, 16'd41835, 16'd2637, 16'd20451, 16'd57445, 16'd20399, 16'd24002, 16'd32312, 16'd43148, 16'd10426, 16'd24005});
	test_expansion(128'hc05be77859cdb1147c714a2b3350c3b8, {16'd1138, 16'd11987, 16'd48300, 16'd4524, 16'd47341, 16'd32033, 16'd19837, 16'd64872, 16'd65233, 16'd45223, 16'd62518, 16'd54936, 16'd4500, 16'd39256, 16'd50933, 16'd24666, 16'd55320, 16'd13303, 16'd65323, 16'd4277, 16'd28339, 16'd21333, 16'd62326, 16'd50678, 16'd40593, 16'd12856});
	test_expansion(128'h2cc11a8b7826e3f93aa06405a2997a47, {16'd55871, 16'd14818, 16'd49448, 16'd28493, 16'd45690, 16'd53071, 16'd58884, 16'd36358, 16'd61815, 16'd32732, 16'd28526, 16'd51676, 16'd56414, 16'd7864, 16'd41067, 16'd3441, 16'd43102, 16'd40460, 16'd60939, 16'd304, 16'd3033, 16'd34539, 16'd254, 16'd9253, 16'd19638, 16'd31852});
	test_expansion(128'h6f6e3a68d8c04b1edee6491ecd9e7674, {16'd63625, 16'd15975, 16'd24137, 16'd14378, 16'd57638, 16'd29186, 16'd49956, 16'd56033, 16'd21619, 16'd63641, 16'd15770, 16'd42094, 16'd33965, 16'd39583, 16'd34110, 16'd20799, 16'd36785, 16'd38121, 16'd41465, 16'd52538, 16'd49265, 16'd49939, 16'd24147, 16'd4011, 16'd20937, 16'd40902});
	test_expansion(128'hebf2051ff3e92eb6506ffae5c9d6ebdd, {16'd6035, 16'd19838, 16'd26670, 16'd61667, 16'd213, 16'd22529, 16'd58124, 16'd48595, 16'd1670, 16'd47012, 16'd40242, 16'd49358, 16'd20411, 16'd59218, 16'd20750, 16'd41581, 16'd30108, 16'd33086, 16'd41579, 16'd41001, 16'd18140, 16'd7209, 16'd64545, 16'd55419, 16'd1239, 16'd11964});
	test_expansion(128'h4ea766bb3bd7a73f039e390bc3831e73, {16'd45462, 16'd45195, 16'd56429, 16'd1540, 16'd6603, 16'd1203, 16'd37898, 16'd28862, 16'd40538, 16'd60035, 16'd34028, 16'd16928, 16'd42446, 16'd13961, 16'd957, 16'd28534, 16'd40487, 16'd23834, 16'd13609, 16'd61911, 16'd63331, 16'd58044, 16'd29992, 16'd49115, 16'd44918, 16'd44680});
	test_expansion(128'h23347317268936f64dd7421ba639f3cf, {16'd22751, 16'd39158, 16'd28706, 16'd5801, 16'd54057, 16'd17054, 16'd45013, 16'd53800, 16'd9613, 16'd23018, 16'd16581, 16'd31908, 16'd26973, 16'd49409, 16'd62132, 16'd38574, 16'd61585, 16'd62094, 16'd28538, 16'd19867, 16'd60826, 16'd44750, 16'd43622, 16'd61404, 16'd58325, 16'd24683});
	test_expansion(128'had17df66d1a60735ca336925e43db188, {16'd40130, 16'd41212, 16'd48049, 16'd16837, 16'd24747, 16'd22030, 16'd15704, 16'd23049, 16'd16848, 16'd34070, 16'd63404, 16'd57734, 16'd57592, 16'd42366, 16'd25241, 16'd35301, 16'd37424, 16'd28444, 16'd25400, 16'd11161, 16'd11648, 16'd51551, 16'd35118, 16'd15804, 16'd59824, 16'd8876});
	test_expansion(128'he8a7d3edd7a75e2216be0cf2299f3a47, {16'd32444, 16'd12024, 16'd24909, 16'd46802, 16'd20866, 16'd28504, 16'd48226, 16'd42201, 16'd10944, 16'd34130, 16'd64976, 16'd3624, 16'd30681, 16'd42255, 16'd4317, 16'd908, 16'd266, 16'd56425, 16'd51392, 16'd45735, 16'd23100, 16'd33642, 16'd47255, 16'd24736, 16'd63532, 16'd40111});
	test_expansion(128'hac438774f079341e85d72e07e1344766, {16'd62814, 16'd65199, 16'd12523, 16'd15575, 16'd40402, 16'd4940, 16'd10855, 16'd24912, 16'd58896, 16'd33866, 16'd26101, 16'd9888, 16'd56442, 16'd49124, 16'd45238, 16'd31933, 16'd9972, 16'd12493, 16'd63429, 16'd14891, 16'd46203, 16'd58786, 16'd4286, 16'd1629, 16'd13106, 16'd36532});
	test_expansion(128'hd2d842772d33716ae36b8ccfd5bfcc5b, {16'd7009, 16'd29601, 16'd2362, 16'd41316, 16'd34357, 16'd32662, 16'd13454, 16'd52269, 16'd30171, 16'd10751, 16'd40953, 16'd2772, 16'd27346, 16'd38556, 16'd47098, 16'd52944, 16'd45946, 16'd19538, 16'd44398, 16'd50167, 16'd10275, 16'd48240, 16'd32227, 16'd47746, 16'd39177, 16'd42814});
	test_expansion(128'h2843f184e88644900421a98f4238cb99, {16'd22164, 16'd36281, 16'd7264, 16'd26861, 16'd9839, 16'd23003, 16'd3979, 16'd45064, 16'd40373, 16'd9020, 16'd51623, 16'd61971, 16'd3200, 16'd42469, 16'd2103, 16'd30509, 16'd47348, 16'd46147, 16'd1143, 16'd23320, 16'd9444, 16'd51326, 16'd55494, 16'd17894, 16'd19729, 16'd50324});
	test_expansion(128'h27e9ee9f6a1cb58a168c4f6488c9b617, {16'd21527, 16'd5999, 16'd1402, 16'd15012, 16'd6855, 16'd41338, 16'd46856, 16'd65049, 16'd8719, 16'd21998, 16'd63734, 16'd10299, 16'd45914, 16'd20436, 16'd21076, 16'd5058, 16'd46289, 16'd43680, 16'd18386, 16'd21609, 16'd25142, 16'd52061, 16'd6702, 16'd64022, 16'd35163, 16'd283});
	test_expansion(128'h8917bf90be133980faf10ebe4a8f2024, {16'd51452, 16'd42973, 16'd43094, 16'd22839, 16'd15937, 16'd11908, 16'd56176, 16'd38379, 16'd40868, 16'd10160, 16'd46857, 16'd12145, 16'd13153, 16'd10833, 16'd13681, 16'd21162, 16'd29675, 16'd53487, 16'd761, 16'd57508, 16'd39424, 16'd25090, 16'd31084, 16'd52664, 16'd39636, 16'd3621});
	test_expansion(128'h0989f2589387bea2aab5733804dfaf3a, {16'd34892, 16'd62659, 16'd52407, 16'd3919, 16'd10878, 16'd62090, 16'd43989, 16'd41197, 16'd35625, 16'd39214, 16'd39332, 16'd26838, 16'd14409, 16'd65305, 16'd34475, 16'd1344, 16'd11872, 16'd60834, 16'd22045, 16'd51385, 16'd22759, 16'd46740, 16'd2275, 16'd54772, 16'd16180, 16'd60129});
	test_expansion(128'hbb9514ceef2de7b7c9e2840fad4f0492, {16'd11325, 16'd65037, 16'd55740, 16'd6905, 16'd47650, 16'd14009, 16'd29387, 16'd61889, 16'd45153, 16'd34545, 16'd29695, 16'd44459, 16'd1471, 16'd11249, 16'd9937, 16'd7267, 16'd17573, 16'd3532, 16'd28657, 16'd6212, 16'd18161, 16'd15056, 16'd30657, 16'd49871, 16'd23645, 16'd47228});
	test_expansion(128'h7ccc0c4c559ddccd802403ff6faef41f, {16'd60743, 16'd62680, 16'd63671, 16'd12095, 16'd35486, 16'd2216, 16'd24679, 16'd56619, 16'd18231, 16'd49850, 16'd39663, 16'd35196, 16'd51628, 16'd54334, 16'd3471, 16'd27390, 16'd19628, 16'd27658, 16'd61305, 16'd22692, 16'd31429, 16'd58209, 16'd61272, 16'd4217, 16'd11731, 16'd8658});
	test_expansion(128'h2573d55eb029a64ff58b0fb490600613, {16'd36889, 16'd57683, 16'd23406, 16'd2410, 16'd57297, 16'd26511, 16'd38817, 16'd29813, 16'd33894, 16'd45363, 16'd16125, 16'd20269, 16'd41871, 16'd64113, 16'd5414, 16'd61057, 16'd26620, 16'd36457, 16'd34007, 16'd36194, 16'd18014, 16'd64990, 16'd732, 16'd37518, 16'd22383, 16'd5622});
	test_expansion(128'hdc11872f3ba218b4c97fb715fbc76994, {16'd18923, 16'd63070, 16'd57275, 16'd11614, 16'd50621, 16'd26621, 16'd61510, 16'd36550, 16'd39372, 16'd16107, 16'd4139, 16'd59998, 16'd37782, 16'd64643, 16'd19205, 16'd22024, 16'd29638, 16'd51202, 16'd39544, 16'd23741, 16'd6547, 16'd38984, 16'd52762, 16'd4096, 16'd26140, 16'd57871});
	test_expansion(128'h4c0591aa1203dc1becac47159f037c98, {16'd17064, 16'd50679, 16'd37239, 16'd31795, 16'd55008, 16'd36307, 16'd23383, 16'd814, 16'd27601, 16'd15471, 16'd9633, 16'd11399, 16'd55718, 16'd3773, 16'd59677, 16'd22976, 16'd64851, 16'd5390, 16'd15960, 16'd14055, 16'd50369, 16'd22867, 16'd8582, 16'd16950, 16'd2254, 16'd40529});
	test_expansion(128'h0267d0d227f915f8a178f9a650e622a6, {16'd56947, 16'd5485, 16'd45792, 16'd3879, 16'd59125, 16'd51619, 16'd50367, 16'd34385, 16'd15747, 16'd16182, 16'd25142, 16'd4233, 16'd33867, 16'd57826, 16'd40439, 16'd29122, 16'd63068, 16'd28926, 16'd62708, 16'd25351, 16'd52973, 16'd60741, 16'd61646, 16'd38324, 16'd19023, 16'd11712});
	test_expansion(128'h3fc4c9e69d76b00f48c65b7cb6fba42c, {16'd59877, 16'd13943, 16'd57155, 16'd51509, 16'd39796, 16'd7220, 16'd29191, 16'd2244, 16'd3102, 16'd21157, 16'd46820, 16'd53830, 16'd5720, 16'd38813, 16'd13869, 16'd236, 16'd9578, 16'd18529, 16'd64362, 16'd47147, 16'd50048, 16'd35696, 16'd28668, 16'd36985, 16'd35739, 16'd44019});
	test_expansion(128'hf91045436bae8662092f53d228df77bc, {16'd19970, 16'd53792, 16'd40550, 16'd20912, 16'd4940, 16'd34807, 16'd13282, 16'd31244, 16'd6592, 16'd26896, 16'd11710, 16'd13225, 16'd38307, 16'd56583, 16'd14239, 16'd17091, 16'd37409, 16'd21094, 16'd33097, 16'd12424, 16'd30763, 16'd63957, 16'd45738, 16'd30129, 16'd44287, 16'd46970});
	test_expansion(128'h7ce4cf24a2f098080a716a3896d74aa0, {16'd32275, 16'd44548, 16'd64056, 16'd44785, 16'd39984, 16'd14126, 16'd4065, 16'd33891, 16'd34773, 16'd50432, 16'd59178, 16'd42074, 16'd17631, 16'd557, 16'd42445, 16'd16330, 16'd8479, 16'd44866, 16'd39740, 16'd9408, 16'd7791, 16'd1325, 16'd31932, 16'd41465, 16'd25670, 16'd25339});
	test_expansion(128'h0ad82b65bba8e46cff15713b4ec29ade, {16'd46979, 16'd43546, 16'd44153, 16'd49263, 16'd49895, 16'd32033, 16'd9067, 16'd43754, 16'd62924, 16'd5393, 16'd31135, 16'd58331, 16'd46814, 16'd11637, 16'd24888, 16'd5108, 16'd7398, 16'd54818, 16'd22208, 16'd1723, 16'd3034, 16'd43175, 16'd44911, 16'd6410, 16'd31896, 16'd54220});
	test_expansion(128'h527c612d556a1e6f88c0fa5286eb3fe4, {16'd62381, 16'd59559, 16'd1564, 16'd15492, 16'd22230, 16'd63917, 16'd17867, 16'd8440, 16'd47142, 16'd19477, 16'd52466, 16'd4729, 16'd574, 16'd41853, 16'd27009, 16'd44907, 16'd21537, 16'd33675, 16'd9334, 16'd12721, 16'd51627, 16'd14480, 16'd25599, 16'd16315, 16'd16146, 16'd64138});
	test_expansion(128'h8b0132931006d09455a42ba49110e5e4, {16'd43249, 16'd41421, 16'd58427, 16'd60596, 16'd15970, 16'd43308, 16'd15660, 16'd65336, 16'd44455, 16'd17143, 16'd45091, 16'd32524, 16'd37968, 16'd21738, 16'd15394, 16'd39584, 16'd45937, 16'd21098, 16'd20412, 16'd38607, 16'd62392, 16'd38168, 16'd37508, 16'd51670, 16'd37403, 16'd2696});
	test_expansion(128'h4e7a0adc3c2620e254c0b09fd62534c6, {16'd15185, 16'd12286, 16'd58260, 16'd24854, 16'd54969, 16'd46888, 16'd54345, 16'd35226, 16'd19883, 16'd60678, 16'd40136, 16'd21846, 16'd8467, 16'd43540, 16'd20311, 16'd5968, 16'd29239, 16'd49682, 16'd45153, 16'd41900, 16'd56270, 16'd21673, 16'd28876, 16'd40130, 16'd55720, 16'd49640});
	test_expansion(128'ha6ed9e70efb83f0ca87758a3037dd67b, {16'd40629, 16'd49502, 16'd20499, 16'd46802, 16'd42302, 16'd62977, 16'd4623, 16'd13442, 16'd48867, 16'd21218, 16'd28728, 16'd25458, 16'd28924, 16'd65435, 16'd11828, 16'd57991, 16'd51923, 16'd21059, 16'd55455, 16'd26826, 16'd29447, 16'd42863, 16'd1919, 16'd7610, 16'd50645, 16'd39546});
	test_expansion(128'h39c971d99597c5ddf83de841a3bce70e, {16'd18821, 16'd42182, 16'd5027, 16'd23167, 16'd29732, 16'd39649, 16'd18696, 16'd16040, 16'd41156, 16'd35153, 16'd41175, 16'd11682, 16'd30642, 16'd20902, 16'd14247, 16'd10914, 16'd10368, 16'd21953, 16'd3729, 16'd4884, 16'd45967, 16'd1595, 16'd45787, 16'd11307, 16'd52423, 16'd63456});
	test_expansion(128'h103f8ac7617aba669dbdf9af9a5d3845, {16'd28790, 16'd14030, 16'd61172, 16'd65277, 16'd803, 16'd62176, 16'd45793, 16'd1530, 16'd33796, 16'd57089, 16'd48335, 16'd9864, 16'd59473, 16'd30689, 16'd44459, 16'd62271, 16'd53111, 16'd1671, 16'd18884, 16'd62202, 16'd9110, 16'd55171, 16'd27976, 16'd32937, 16'd27337, 16'd37268});
	test_expansion(128'h23155360ed4318cf65c10a04e547faf8, {16'd42857, 16'd43457, 16'd11944, 16'd36043, 16'd47060, 16'd1522, 16'd65090, 16'd50270, 16'd32606, 16'd52023, 16'd18029, 16'd45099, 16'd1396, 16'd5991, 16'd6959, 16'd6391, 16'd31250, 16'd8493, 16'd20427, 16'd61361, 16'd10698, 16'd1475, 16'd17880, 16'd48971, 16'd28914, 16'd43599});
	test_expansion(128'h01d61653002f6e3c549749c6210b34f2, {16'd13741, 16'd56360, 16'd645, 16'd13962, 16'd38892, 16'd55999, 16'd49750, 16'd3867, 16'd13440, 16'd7089, 16'd53276, 16'd64022, 16'd43336, 16'd60028, 16'd51712, 16'd12750, 16'd25974, 16'd60751, 16'd15070, 16'd64692, 16'd57446, 16'd58670, 16'd37039, 16'd43564, 16'd62014, 16'd1483});
	test_expansion(128'h4a713d3e49307dd42ade0f07e520983f, {16'd53416, 16'd41657, 16'd8193, 16'd40347, 16'd29970, 16'd38654, 16'd43366, 16'd50385, 16'd62227, 16'd54729, 16'd25497, 16'd19545, 16'd3719, 16'd4557, 16'd48938, 16'd39102, 16'd45419, 16'd20821, 16'd35343, 16'd16866, 16'd1920, 16'd17550, 16'd4219, 16'd669, 16'd7323, 16'd40302});
	test_expansion(128'h168fbcccbb393b8ba0cc61577145cb52, {16'd44713, 16'd18343, 16'd39211, 16'd15647, 16'd48533, 16'd11420, 16'd50987, 16'd45492, 16'd60255, 16'd18092, 16'd51225, 16'd51246, 16'd35045, 16'd61291, 16'd11917, 16'd60918, 16'd12884, 16'd26873, 16'd34438, 16'd33156, 16'd48550, 16'd3941, 16'd23725, 16'd6147, 16'd63998, 16'd5234});
	test_expansion(128'h00e5582e620443c40895bfcf2c4458ec, {16'd45028, 16'd50738, 16'd4261, 16'd4538, 16'd45726, 16'd29075, 16'd29885, 16'd58711, 16'd61767, 16'd62520, 16'd9319, 16'd55652, 16'd5660, 16'd31859, 16'd60413, 16'd48792, 16'd36040, 16'd52992, 16'd57164, 16'd46772, 16'd19916, 16'd5269, 16'd58838, 16'd18013, 16'd35273, 16'd56124});
	test_expansion(128'h5bb0fe6add5d922a7b3212b7f33c5c62, {16'd48908, 16'd46677, 16'd40953, 16'd46473, 16'd38288, 16'd5958, 16'd20379, 16'd14903, 16'd14781, 16'd6377, 16'd28929, 16'd42490, 16'd41379, 16'd45623, 16'd56249, 16'd40758, 16'd42751, 16'd64284, 16'd23034, 16'd57168, 16'd34578, 16'd38431, 16'd43266, 16'd63435, 16'd12677, 16'd54154});
	test_expansion(128'h0de582dae28002dae55d0e658b18eea1, {16'd12872, 16'd41589, 16'd22931, 16'd47587, 16'd33167, 16'd20734, 16'd13500, 16'd40168, 16'd40928, 16'd12699, 16'd20355, 16'd64675, 16'd15331, 16'd23669, 16'd54042, 16'd22530, 16'd9283, 16'd43108, 16'd30527, 16'd7231, 16'd60076, 16'd22637, 16'd58719, 16'd52506, 16'd64577, 16'd19704});
	test_expansion(128'had67aced39d80ba077be18d019aa18bc, {16'd29350, 16'd149, 16'd45783, 16'd11813, 16'd54324, 16'd65248, 16'd64955, 16'd37827, 16'd63295, 16'd42719, 16'd63214, 16'd51617, 16'd16023, 16'd35975, 16'd565, 16'd828, 16'd40956, 16'd56180, 16'd56309, 16'd55587, 16'd52707, 16'd18822, 16'd39439, 16'd39715, 16'd39067, 16'd27295});
	test_expansion(128'h9046e3003acb7ec154c425d051869ac7, {16'd53007, 16'd36924, 16'd34581, 16'd59687, 16'd2678, 16'd46847, 16'd16945, 16'd58653, 16'd38868, 16'd45708, 16'd31400, 16'd53318, 16'd52443, 16'd13272, 16'd12249, 16'd35605, 16'd3059, 16'd15790, 16'd31302, 16'd24178, 16'd7847, 16'd55084, 16'd46876, 16'd31996, 16'd21586, 16'd49480});
	test_expansion(128'h672963a06d39f679175e81e6592995ad, {16'd32561, 16'd16392, 16'd732, 16'd23221, 16'd6263, 16'd53131, 16'd38334, 16'd55664, 16'd64597, 16'd52046, 16'd35069, 16'd55211, 16'd17050, 16'd36104, 16'd54963, 16'd3343, 16'd24350, 16'd29206, 16'd60211, 16'd39515, 16'd30954, 16'd16306, 16'd61201, 16'd12369, 16'd61371, 16'd13241});
	test_expansion(128'hd5a6f571cd75f62ccc251099c4595240, {16'd35613, 16'd36121, 16'd51102, 16'd52963, 16'd12038, 16'd54581, 16'd41688, 16'd36738, 16'd24546, 16'd58571, 16'd47437, 16'd4842, 16'd59840, 16'd47548, 16'd7631, 16'd1509, 16'd62078, 16'd31440, 16'd7167, 16'd20207, 16'd34675, 16'd32736, 16'd62285, 16'd32122, 16'd46292, 16'd54761});
	test_expansion(128'hd85b680e378b87ad4f61d8500e70dd0e, {16'd53964, 16'd34988, 16'd18814, 16'd27741, 16'd19065, 16'd18604, 16'd20389, 16'd49955, 16'd12121, 16'd20567, 16'd2545, 16'd39891, 16'd52599, 16'd64048, 16'd16262, 16'd25302, 16'd34646, 16'd15574, 16'd10037, 16'd5153, 16'd57881, 16'd57485, 16'd53168, 16'd38110, 16'd20618, 16'd39573});
	test_expansion(128'h337fd7aa727a9c2226ebe34f57884e5e, {16'd58654, 16'd40301, 16'd26806, 16'd51208, 16'd54204, 16'd65532, 16'd49346, 16'd60320, 16'd55311, 16'd33367, 16'd53568, 16'd11247, 16'd20833, 16'd44433, 16'd58368, 16'd15153, 16'd27137, 16'd28436, 16'd55206, 16'd24878, 16'd29073, 16'd57356, 16'd6824, 16'd32096, 16'd23838, 16'd23458});
	test_expansion(128'hc00eee05f4d075cba5d4cbda66d3d635, {16'd34227, 16'd13711, 16'd49738, 16'd54149, 16'd11118, 16'd55211, 16'd15311, 16'd60042, 16'd5711, 16'd33696, 16'd30849, 16'd37540, 16'd18480, 16'd64822, 16'd61883, 16'd42927, 16'd3531, 16'd19191, 16'd55766, 16'd39801, 16'd44025, 16'd28186, 16'd50516, 16'd3488, 16'd18540, 16'd54314});
	test_expansion(128'h4cc1be6b519c77bbe207bfa2be8f1a5d, {16'd62004, 16'd39529, 16'd63398, 16'd10353, 16'd57875, 16'd61153, 16'd9817, 16'd42385, 16'd51274, 16'd39241, 16'd18000, 16'd46272, 16'd37335, 16'd12262, 16'd41528, 16'd3828, 16'd17234, 16'd43851, 16'd37964, 16'd54481, 16'd31502, 16'd9057, 16'd42330, 16'd59511, 16'd58585, 16'd61647});
	test_expansion(128'hb86d027358d261b7f6bf8d46f4121dcb, {16'd23926, 16'd39977, 16'd31667, 16'd36079, 16'd17221, 16'd1182, 16'd63632, 16'd60388, 16'd4067, 16'd16507, 16'd58442, 16'd64296, 16'd11829, 16'd3177, 16'd62192, 16'd22972, 16'd1586, 16'd3366, 16'd34813, 16'd40292, 16'd37453, 16'd49300, 16'd39465, 16'd8864, 16'd23947, 16'd214});
	test_expansion(128'h8709e7aaf211679494f48f797c8111a0, {16'd31090, 16'd62911, 16'd31778, 16'd30705, 16'd30733, 16'd12105, 16'd48980, 16'd46882, 16'd40651, 16'd35362, 16'd59729, 16'd29908, 16'd55316, 16'd53790, 16'd6891, 16'd3297, 16'd37695, 16'd9694, 16'd8689, 16'd23558, 16'd45053, 16'd25215, 16'd12482, 16'd52332, 16'd50978, 16'd30554});
	test_expansion(128'hff346262db19421e6cacbbe2de87dc2b, {16'd3708, 16'd29454, 16'd4895, 16'd63391, 16'd52636, 16'd60151, 16'd41757, 16'd35613, 16'd24133, 16'd2688, 16'd41642, 16'd13977, 16'd5393, 16'd37920, 16'd53565, 16'd34557, 16'd57441, 16'd58656, 16'd30449, 16'd28478, 16'd2849, 16'd33575, 16'd46563, 16'd64910, 16'd25045, 16'd50926});
	test_expansion(128'h3f6b695b7b8fce6fc961eaad890de2a6, {16'd32752, 16'd40517, 16'd55943, 16'd4104, 16'd10852, 16'd30051, 16'd10396, 16'd30889, 16'd52434, 16'd45823, 16'd37869, 16'd31036, 16'd40666, 16'd62796, 16'd46006, 16'd53085, 16'd53051, 16'd43301, 16'd60542, 16'd55665, 16'd37982, 16'd26159, 16'd39152, 16'd16565, 16'd53913, 16'd9741});
	test_expansion(128'h89546fcae92cef9f188208da724ce6b4, {16'd54702, 16'd41631, 16'd52501, 16'd70, 16'd43835, 16'd26061, 16'd15974, 16'd7608, 16'd7573, 16'd6768, 16'd1128, 16'd46405, 16'd29398, 16'd32546, 16'd40945, 16'd48419, 16'd61386, 16'd38853, 16'd56464, 16'd49687, 16'd29782, 16'd61386, 16'd64864, 16'd47855, 16'd29265, 16'd21475});
	test_expansion(128'h735c65db5577e0bba6a10da6657036c6, {16'd46571, 16'd13022, 16'd30133, 16'd51786, 16'd35893, 16'd27663, 16'd14084, 16'd59031, 16'd53197, 16'd6141, 16'd51282, 16'd23161, 16'd23357, 16'd60997, 16'd56521, 16'd33383, 16'd25734, 16'd43275, 16'd41436, 16'd46523, 16'd48752, 16'd12657, 16'd19088, 16'd15349, 16'd16520, 16'd41408});
	test_expansion(128'h36e5de59f0209ec887d08b15acb44aed, {16'd15575, 16'd7092, 16'd19082, 16'd10997, 16'd48252, 16'd55174, 16'd15481, 16'd56058, 16'd33461, 16'd34498, 16'd53658, 16'd31190, 16'd18945, 16'd59914, 16'd37296, 16'd37760, 16'd335, 16'd43593, 16'd5765, 16'd18949, 16'd24774, 16'd59570, 16'd27593, 16'd57192, 16'd39753, 16'd65297});
	test_expansion(128'h09a194eb28c2c07a2cdaf18d6ab36b92, {16'd2299, 16'd35675, 16'd10617, 16'd64132, 16'd29779, 16'd46371, 16'd43516, 16'd4598, 16'd43977, 16'd45712, 16'd64479, 16'd24678, 16'd21934, 16'd8573, 16'd42326, 16'd58101, 16'd2287, 16'd53175, 16'd7770, 16'd369, 16'd25231, 16'd16781, 16'd11701, 16'd18681, 16'd17643, 16'd3650});
	test_expansion(128'hd0f6f35131385770bade5fd02515c133, {16'd6142, 16'd48902, 16'd44909, 16'd64281, 16'd58257, 16'd34521, 16'd48622, 16'd28033, 16'd60946, 16'd52289, 16'd43737, 16'd32101, 16'd10463, 16'd44408, 16'd43223, 16'd64590, 16'd29744, 16'd7083, 16'd8061, 16'd14120, 16'd27069, 16'd44843, 16'd61519, 16'd16559, 16'd54795, 16'd9626});
	test_expansion(128'h64378930231b4a85713ef6dd40fbeb81, {16'd20250, 16'd11721, 16'd60636, 16'd52155, 16'd21651, 16'd8199, 16'd60159, 16'd20186, 16'd41390, 16'd36912, 16'd35356, 16'd32397, 16'd63315, 16'd45586, 16'd748, 16'd56501, 16'd40688, 16'd56223, 16'd21588, 16'd19061, 16'd29721, 16'd49710, 16'd33030, 16'd11881, 16'd27142, 16'd25351});
	test_expansion(128'hc392cee28988ef113376df01194f4ee9, {16'd24695, 16'd22020, 16'd44188, 16'd16445, 16'd40664, 16'd43653, 16'd63872, 16'd1782, 16'd14975, 16'd8420, 16'd47432, 16'd8703, 16'd1053, 16'd40562, 16'd64648, 16'd55551, 16'd59830, 16'd25626, 16'd55240, 16'd58686, 16'd35980, 16'd32973, 16'd40725, 16'd44885, 16'd35297, 16'd27667});
	test_expansion(128'h024b71684ac47025bd25d09919d692b9, {16'd12421, 16'd8598, 16'd50281, 16'd18051, 16'd31246, 16'd60829, 16'd32878, 16'd62336, 16'd45382, 16'd17999, 16'd44484, 16'd19024, 16'd41439, 16'd438, 16'd21637, 16'd53327, 16'd13389, 16'd5133, 16'd9197, 16'd41363, 16'd6684, 16'd29956, 16'd24697, 16'd202, 16'd45108, 16'd13544});
	test_expansion(128'h463e148e80a69d39df58829895c3475e, {16'd23275, 16'd50170, 16'd22675, 16'd20959, 16'd61091, 16'd17377, 16'd20361, 16'd24628, 16'd17093, 16'd48048, 16'd39280, 16'd37658, 16'd61379, 16'd31097, 16'd12637, 16'd23263, 16'd29962, 16'd32148, 16'd51159, 16'd61294, 16'd61420, 16'd49670, 16'd54340, 16'd40076, 16'd3050, 16'd51230});
	test_expansion(128'had378732103db60704a793ef923b2d00, {16'd1223, 16'd12499, 16'd15181, 16'd11430, 16'd2401, 16'd59771, 16'd5293, 16'd65237, 16'd26707, 16'd56628, 16'd59372, 16'd45395, 16'd49919, 16'd16310, 16'd3870, 16'd59277, 16'd2249, 16'd36832, 16'd46575, 16'd65407, 16'd32459, 16'd34885, 16'd5993, 16'd38227, 16'd10700, 16'd3050});
	test_expansion(128'h5df4855cf2d4e6e2180c11b6fb56826a, {16'd31149, 16'd55614, 16'd51850, 16'd43640, 16'd42705, 16'd17171, 16'd33322, 16'd59099, 16'd12125, 16'd47014, 16'd25716, 16'd4352, 16'd51567, 16'd45350, 16'd6745, 16'd9080, 16'd22261, 16'd30615, 16'd39994, 16'd56607, 16'd44645, 16'd41602, 16'd51242, 16'd36261, 16'd2833, 16'd20210});
	test_expansion(128'h3b77792912c77a54f069e4dac8347c99, {16'd36020, 16'd3967, 16'd58993, 16'd38623, 16'd2674, 16'd42063, 16'd21190, 16'd4159, 16'd45529, 16'd7447, 16'd9757, 16'd29047, 16'd47784, 16'd7835, 16'd60156, 16'd33819, 16'd849, 16'd43299, 16'd31799, 16'd42352, 16'd28902, 16'd16862, 16'd36209, 16'd12344, 16'd8025, 16'd59691});
	test_expansion(128'hb1fbf17bedc97f61a7d7bcc580513c94, {16'd6617, 16'd17324, 16'd8507, 16'd44054, 16'd41839, 16'd62286, 16'd39456, 16'd56710, 16'd44800, 16'd34700, 16'd39133, 16'd40875, 16'd60591, 16'd31067, 16'd12505, 16'd4523, 16'd15143, 16'd2887, 16'd3808, 16'd56068, 16'd62995, 16'd20110, 16'd34425, 16'd53683, 16'd41056, 16'd26446});
	test_expansion(128'hab7e8d015f01e5e721ba185fc308b4fb, {16'd661, 16'd10283, 16'd32530, 16'd52837, 16'd30233, 16'd1911, 16'd8514, 16'd53106, 16'd20001, 16'd58069, 16'd50038, 16'd45902, 16'd23725, 16'd34121, 16'd51068, 16'd56289, 16'd27944, 16'd7054, 16'd23414, 16'd7919, 16'd59155, 16'd42173, 16'd43517, 16'd3496, 16'd9893, 16'd62057});
	test_expansion(128'h378b6ddd21952b38cf1d5174ece38307, {16'd52735, 16'd9590, 16'd57461, 16'd37463, 16'd13101, 16'd64754, 16'd38266, 16'd12288, 16'd54022, 16'd52456, 16'd12940, 16'd32706, 16'd40037, 16'd24126, 16'd842, 16'd6863, 16'd44919, 16'd61106, 16'd54010, 16'd45345, 16'd15991, 16'd6143, 16'd22278, 16'd7058, 16'd57799, 16'd9986});
	test_expansion(128'h38ef5717ce7d6c3918eb52ec68126579, {16'd5269, 16'd40985, 16'd47564, 16'd30988, 16'd57085, 16'd20377, 16'd42803, 16'd20844, 16'd22491, 16'd46983, 16'd36890, 16'd4995, 16'd4049, 16'd1253, 16'd10252, 16'd47214, 16'd8896, 16'd38845, 16'd61166, 16'd28884, 16'd9402, 16'd29139, 16'd14223, 16'd46462, 16'd34009, 16'd8837});
	test_expansion(128'hf3533e5efeef81ec932a514752d63755, {16'd64590, 16'd29739, 16'd60781, 16'd9512, 16'd44841, 16'd2006, 16'd26375, 16'd13198, 16'd20785, 16'd26309, 16'd38377, 16'd22382, 16'd61053, 16'd3757, 16'd57132, 16'd58966, 16'd16769, 16'd44463, 16'd22078, 16'd40393, 16'd1978, 16'd45421, 16'd34007, 16'd40460, 16'd40596, 16'd49825});
	test_expansion(128'h6b7990d775b843e28c91dffd3c01be3b, {16'd58462, 16'd36620, 16'd31256, 16'd46756, 16'd52952, 16'd9856, 16'd24154, 16'd10519, 16'd18805, 16'd54194, 16'd32900, 16'd38112, 16'd20869, 16'd38833, 16'd14431, 16'd46006, 16'd45782, 16'd32988, 16'd13359, 16'd51826, 16'd21237, 16'd46801, 16'd59827, 16'd34692, 16'd12148, 16'd23182});
	test_expansion(128'he7b990c1a0678988747001bca8fdc81d, {16'd47466, 16'd3827, 16'd35814, 16'd13469, 16'd21163, 16'd4329, 16'd50401, 16'd37167, 16'd57153, 16'd57607, 16'd54615, 16'd37492, 16'd19260, 16'd56874, 16'd57160, 16'd13207, 16'd11864, 16'd45527, 16'd12074, 16'd54284, 16'd45787, 16'd50156, 16'd63765, 16'd54963, 16'd480, 16'd1442});
	test_expansion(128'hdfbc5546f117500e24560bd7d0aaee11, {16'd42857, 16'd22496, 16'd8231, 16'd15629, 16'd42760, 16'd4426, 16'd40269, 16'd46296, 16'd27518, 16'd15591, 16'd27697, 16'd46212, 16'd33577, 16'd1745, 16'd3976, 16'd42603, 16'd36757, 16'd46087, 16'd30361, 16'd64434, 16'd28631, 16'd41517, 16'd54355, 16'd61819, 16'd53476, 16'd27868});
	test_expansion(128'h7f4872756bef743c607265626f06827b, {16'd16195, 16'd38913, 16'd62987, 16'd22380, 16'd28524, 16'd24713, 16'd2919, 16'd46793, 16'd58578, 16'd16382, 16'd46530, 16'd983, 16'd56921, 16'd28683, 16'd59142, 16'd49356, 16'd36972, 16'd791, 16'd53733, 16'd9572, 16'd17299, 16'd46336, 16'd25717, 16'd47010, 16'd7529, 16'd24142});
	test_expansion(128'hb3412ade19d0afc7f303cc9fdd56f6d0, {16'd11547, 16'd17883, 16'd11869, 16'd30986, 16'd32363, 16'd22841, 16'd48251, 16'd31488, 16'd48441, 16'd40432, 16'd36088, 16'd64849, 16'd48663, 16'd62956, 16'd4646, 16'd59811, 16'd39340, 16'd31394, 16'd2698, 16'd5914, 16'd62523, 16'd33096, 16'd40819, 16'd33679, 16'd64601, 16'd45802});
	test_expansion(128'h5e20590ce375d567624068f6e7978a7d, {16'd24752, 16'd31252, 16'd64646, 16'd13809, 16'd39858, 16'd44885, 16'd56461, 16'd45744, 16'd35060, 16'd31508, 16'd29708, 16'd14455, 16'd98, 16'd3871, 16'd11044, 16'd38381, 16'd44157, 16'd18755, 16'd58700, 16'd5066, 16'd4822, 16'd21571, 16'd61973, 16'd36408, 16'd18803, 16'd50224});
	test_expansion(128'h1eb23e8fdeb7851bfda9bd21000deb6a, {16'd19044, 16'd6838, 16'd24043, 16'd60449, 16'd6341, 16'd59384, 16'd38615, 16'd30770, 16'd35104, 16'd57881, 16'd27542, 16'd59702, 16'd64988, 16'd52862, 16'd14785, 16'd42170, 16'd41171, 16'd10068, 16'd14925, 16'd42286, 16'd40404, 16'd39604, 16'd50678, 16'd25042, 16'd39609, 16'd24091});
	test_expansion(128'h894ff62f3b72639fa52151cf28db9f13, {16'd37843, 16'd36825, 16'd61914, 16'd52357, 16'd198, 16'd39477, 16'd5628, 16'd26855, 16'd9136, 16'd42982, 16'd57292, 16'd63315, 16'd45022, 16'd60528, 16'd51902, 16'd23468, 16'd8460, 16'd25620, 16'd22300, 16'd48399, 16'd60590, 16'd37543, 16'd34338, 16'd25824, 16'd4275, 16'd62030});
	test_expansion(128'hbf444857883d4be897c77990015a6d67, {16'd37474, 16'd27995, 16'd59297, 16'd54898, 16'd52547, 16'd42292, 16'd50042, 16'd33073, 16'd41108, 16'd54664, 16'd8366, 16'd54331, 16'd3404, 16'd33354, 16'd62992, 16'd9097, 16'd44278, 16'd7781, 16'd7460, 16'd13493, 16'd19079, 16'd47731, 16'd11386, 16'd5261, 16'd10918, 16'd60425});
	test_expansion(128'h7c45396699b5caf61f73680fc533378f, {16'd43192, 16'd33110, 16'd50295, 16'd64621, 16'd49904, 16'd46973, 16'd2417, 16'd38396, 16'd30050, 16'd14167, 16'd52154, 16'd16199, 16'd999, 16'd18064, 16'd27607, 16'd49455, 16'd47495, 16'd9933, 16'd20597, 16'd6529, 16'd17735, 16'd23387, 16'd41712, 16'd37339, 16'd21548, 16'd38319});
	test_expansion(128'h643dc2709b41246ab575e5da9ca8a85b, {16'd39990, 16'd14187, 16'd16396, 16'd1333, 16'd20500, 16'd46520, 16'd38035, 16'd8031, 16'd14921, 16'd19719, 16'd24065, 16'd54727, 16'd22645, 16'd17773, 16'd59793, 16'd63114, 16'd21513, 16'd29415, 16'd18811, 16'd4120, 16'd9275, 16'd14215, 16'd9964, 16'd59293, 16'd63656, 16'd53513});
	test_expansion(128'h811bf662db03ae7d49162626ea2fa425, {16'd34345, 16'd59090, 16'd19264, 16'd4053, 16'd10325, 16'd26162, 16'd1022, 16'd19890, 16'd42008, 16'd61225, 16'd31371, 16'd25390, 16'd54949, 16'd20042, 16'd11326, 16'd19655, 16'd51306, 16'd63103, 16'd12390, 16'd55584, 16'd57222, 16'd46104, 16'd18928, 16'd26403, 16'd3422, 16'd29822});
	test_expansion(128'hd8cb2fd61957c7e48262b8d1bd2c4ce8, {16'd43323, 16'd57104, 16'd46800, 16'd192, 16'd12746, 16'd21653, 16'd42164, 16'd45872, 16'd41518, 16'd26861, 16'd56550, 16'd6451, 16'd49431, 16'd23970, 16'd1674, 16'd8341, 16'd25298, 16'd61499, 16'd52328, 16'd29502, 16'd10584, 16'd27886, 16'd58520, 16'd46583, 16'd57883, 16'd24440});
	test_expansion(128'hbd060fcc249ba05e15d59b0e5d946c7d, {16'd58081, 16'd46596, 16'd38361, 16'd36519, 16'd45186, 16'd47051, 16'd32168, 16'd30365, 16'd10438, 16'd13917, 16'd36800, 16'd53393, 16'd55579, 16'd2601, 16'd59708, 16'd38237, 16'd24034, 16'd43371, 16'd38266, 16'd4213, 16'd12398, 16'd31012, 16'd51581, 16'd26023, 16'd34351, 16'd27088});
	test_expansion(128'h0f5f9db4a45fa3881f90e5698237df42, {16'd31082, 16'd49815, 16'd9942, 16'd11477, 16'd57911, 16'd20076, 16'd32879, 16'd46015, 16'd29127, 16'd60195, 16'd14028, 16'd11240, 16'd23172, 16'd35599, 16'd56519, 16'd19664, 16'd10702, 16'd35902, 16'd36968, 16'd19268, 16'd60384, 16'd37672, 16'd13592, 16'd5969, 16'd30059, 16'd20563});
	test_expansion(128'h2cec5a690238aca7fe207012a58d4904, {16'd6669, 16'd39234, 16'd58334, 16'd48136, 16'd28579, 16'd40133, 16'd25677, 16'd31599, 16'd4020, 16'd14886, 16'd15974, 16'd36319, 16'd16582, 16'd40738, 16'd51806, 16'd11988, 16'd1813, 16'd5151, 16'd56847, 16'd32614, 16'd40541, 16'd37003, 16'd38209, 16'd1000, 16'd33824, 16'd21430});
	test_expansion(128'h735ab5b04ca501888291816fa8e9aad9, {16'd46280, 16'd46464, 16'd5915, 16'd3325, 16'd29776, 16'd9179, 16'd38967, 16'd57751, 16'd46961, 16'd40397, 16'd34538, 16'd3817, 16'd916, 16'd12381, 16'd35380, 16'd18751, 16'd60748, 16'd39256, 16'd49742, 16'd4896, 16'd26106, 16'd3370, 16'd25194, 16'd31980, 16'd44050, 16'd21015});
	test_expansion(128'h399c33c94b56a953d57139714808d8d9, {16'd56097, 16'd36542, 16'd43903, 16'd8190, 16'd2577, 16'd23023, 16'd44741, 16'd37978, 16'd35571, 16'd1260, 16'd123, 16'd64093, 16'd57958, 16'd2385, 16'd64033, 16'd41785, 16'd2165, 16'd40097, 16'd16425, 16'd42046, 16'd40159, 16'd26131, 16'd13995, 16'd6251, 16'd23931, 16'd35848});
	test_expansion(128'h93fc4073fddc660efb6591fbefbd8298, {16'd17627, 16'd33605, 16'd36645, 16'd62902, 16'd19328, 16'd3074, 16'd50146, 16'd60860, 16'd45612, 16'd7183, 16'd16698, 16'd36490, 16'd64813, 16'd52126, 16'd13849, 16'd11487, 16'd46246, 16'd30436, 16'd58003, 16'd65045, 16'd42824, 16'd36272, 16'd20567, 16'd53411, 16'd52013, 16'd48486});
	test_expansion(128'h0d7988d01c64b94cc20b563c04510969, {16'd60638, 16'd3802, 16'd41000, 16'd62588, 16'd11831, 16'd46875, 16'd36930, 16'd24637, 16'd36045, 16'd54920, 16'd29523, 16'd47328, 16'd10116, 16'd9024, 16'd3876, 16'd5656, 16'd30901, 16'd25274, 16'd54702, 16'd10951, 16'd37849, 16'd32187, 16'd27167, 16'd33435, 16'd8042, 16'd41081});
	test_expansion(128'hc7525db6a8764cf7e1a71e963c5596fd, {16'd33464, 16'd8377, 16'd15439, 16'd12431, 16'd49665, 16'd19564, 16'd56670, 16'd16310, 16'd46471, 16'd39510, 16'd44152, 16'd59388, 16'd3506, 16'd3321, 16'd62654, 16'd57531, 16'd34708, 16'd40876, 16'd50876, 16'd60833, 16'd32103, 16'd28106, 16'd62434, 16'd44335, 16'd18696, 16'd37484});
	test_expansion(128'hc84213bae8c37fabf12a0506b072ef40, {16'd63757, 16'd38890, 16'd2029, 16'd64363, 16'd58636, 16'd7620, 16'd50611, 16'd44987, 16'd65106, 16'd12849, 16'd50022, 16'd56172, 16'd33306, 16'd32995, 16'd12022, 16'd17099, 16'd9548, 16'd3018, 16'd27363, 16'd29640, 16'd12502, 16'd23849, 16'd37035, 16'd35903, 16'd15701, 16'd58766});
	test_expansion(128'h06e2455bd9f0a15957397f7baa91d00a, {16'd2055, 16'd410, 16'd37251, 16'd47637, 16'd53203, 16'd44992, 16'd58676, 16'd50462, 16'd50359, 16'd51364, 16'd28345, 16'd28024, 16'd46998, 16'd34825, 16'd35031, 16'd501, 16'd62529, 16'd28347, 16'd40804, 16'd51372, 16'd4630, 16'd7277, 16'd23381, 16'd2236, 16'd6289, 16'd61567});
	test_expansion(128'h2997e81ac6ee24d1e0fae6f8fe074beb, {16'd540, 16'd58647, 16'd37005, 16'd29079, 16'd64133, 16'd39244, 16'd25498, 16'd48727, 16'd4463, 16'd52854, 16'd64280, 16'd34375, 16'd29992, 16'd2005, 16'd48996, 16'd43446, 16'd312, 16'd63401, 16'd58001, 16'd2805, 16'd2742, 16'd56398, 16'd15443, 16'd51292, 16'd27547, 16'd56478});
	test_expansion(128'h4aa957e75944b1ba3f7556d1d29f9779, {16'd56504, 16'd40513, 16'd63042, 16'd45227, 16'd60787, 16'd17969, 16'd23453, 16'd15703, 16'd46073, 16'd33013, 16'd62961, 16'd45330, 16'd64487, 16'd19433, 16'd51655, 16'd11289, 16'd19608, 16'd43141, 16'd58035, 16'd44208, 16'd46457, 16'd40315, 16'd61061, 16'd57619, 16'd63668, 16'd25451});
	test_expansion(128'h663832c7164e62a07d9f1427129fddc2, {16'd23650, 16'd34271, 16'd46679, 16'd39983, 16'd2642, 16'd49005, 16'd49516, 16'd52275, 16'd18952, 16'd51675, 16'd33543, 16'd4927, 16'd20544, 16'd24901, 16'd30183, 16'd13798, 16'd50779, 16'd48202, 16'd5951, 16'd45935, 16'd12285, 16'd22053, 16'd16697, 16'd64021, 16'd10828, 16'd13842});
	test_expansion(128'hd5f528ddfa0f1b3988991c1c6f7bfe95, {16'd61330, 16'd18822, 16'd44350, 16'd40955, 16'd18862, 16'd37006, 16'd3782, 16'd30079, 16'd62897, 16'd25680, 16'd56491, 16'd12593, 16'd16089, 16'd27651, 16'd63348, 16'd22360, 16'd36147, 16'd3978, 16'd43423, 16'd27695, 16'd45147, 16'd37925, 16'd45669, 16'd45718, 16'd52460, 16'd54483});
	test_expansion(128'hf6f065c8ce9b32689aa82ac16b9f0410, {16'd55221, 16'd30887, 16'd47503, 16'd64170, 16'd35805, 16'd46024, 16'd41281, 16'd23952, 16'd61775, 16'd7231, 16'd52971, 16'd2152, 16'd57543, 16'd2380, 16'd35542, 16'd40470, 16'd40885, 16'd20797, 16'd16943, 16'd42742, 16'd12829, 16'd59272, 16'd31446, 16'd45453, 16'd47928, 16'd46355});
	test_expansion(128'h020997ab7914021a0cf77b69e5bc9433, {16'd58840, 16'd20579, 16'd35584, 16'd59658, 16'd46496, 16'd3321, 16'd51774, 16'd29772, 16'd27055, 16'd3405, 16'd25523, 16'd4031, 16'd26703, 16'd13763, 16'd6927, 16'd36386, 16'd57144, 16'd47186, 16'd10938, 16'd15232, 16'd29791, 16'd56799, 16'd52538, 16'd61101, 16'd45068, 16'd39150});
	test_expansion(128'h690f0d9985be24681f0fb532870f4a4d, {16'd30665, 16'd26954, 16'd2167, 16'd32291, 16'd46677, 16'd35222, 16'd14223, 16'd52060, 16'd39389, 16'd15064, 16'd48183, 16'd34244, 16'd13322, 16'd2026, 16'd24052, 16'd52737, 16'd17012, 16'd47715, 16'd16335, 16'd11877, 16'd9944, 16'd27825, 16'd27923, 16'd10195, 16'd52648, 16'd47567});
	test_expansion(128'h5f887734a9fab8a05a3949241cae37de, {16'd63252, 16'd40879, 16'd13919, 16'd40202, 16'd25644, 16'd36790, 16'd14830, 16'd851, 16'd3024, 16'd28334, 16'd22895, 16'd44544, 16'd45916, 16'd35072, 16'd60434, 16'd24891, 16'd8196, 16'd39558, 16'd38348, 16'd32225, 16'd19310, 16'd46015, 16'd59403, 16'd14594, 16'd3730, 16'd2705});
	test_expansion(128'heb2a6ae11e3ea58d292a7296ab241700, {16'd22543, 16'd42056, 16'd4451, 16'd9405, 16'd2259, 16'd25614, 16'd34198, 16'd34095, 16'd6713, 16'd3736, 16'd9495, 16'd43631, 16'd31883, 16'd50203, 16'd41678, 16'd56205, 16'd13612, 16'd14948, 16'd18909, 16'd50821, 16'd34180, 16'd58922, 16'd19084, 16'd22832, 16'd23372, 16'd9289});
	test_expansion(128'hfcc676a28acb4a033694641140e92ea5, {16'd62261, 16'd1193, 16'd9222, 16'd20807, 16'd28440, 16'd31481, 16'd43129, 16'd39018, 16'd238, 16'd20623, 16'd37124, 16'd34681, 16'd30589, 16'd23518, 16'd27182, 16'd1151, 16'd4796, 16'd61788, 16'd24047, 16'd28832, 16'd55367, 16'd30522, 16'd41286, 16'd19787, 16'd28495, 16'd17446});
	test_expansion(128'hf7c2aeb83f658cdb54d2935ae74a191b, {16'd62495, 16'd63488, 16'd16229, 16'd63934, 16'd34078, 16'd38385, 16'd14171, 16'd18626, 16'd34899, 16'd9656, 16'd11400, 16'd24799, 16'd40404, 16'd42719, 16'd49050, 16'd51423, 16'd15535, 16'd14987, 16'd3317, 16'd58463, 16'd43510, 16'd51251, 16'd33121, 16'd32963, 16'd13026, 16'd56902});
	test_expansion(128'hfe05df12bd687ef6476f25215c5f71bd, {16'd11430, 16'd33612, 16'd40358, 16'd7655, 16'd16718, 16'd49757, 16'd48080, 16'd9383, 16'd30670, 16'd1999, 16'd15745, 16'd34164, 16'd301, 16'd56086, 16'd20389, 16'd43563, 16'd56879, 16'd52768, 16'd30073, 16'd61982, 16'd22386, 16'd11464, 16'd14050, 16'd18367, 16'd25033, 16'd41812});
	test_expansion(128'h402260f3c1b78f8b0073a2c1e0b1b929, {16'd30441, 16'd59814, 16'd13477, 16'd5146, 16'd59109, 16'd63757, 16'd23516, 16'd17082, 16'd28283, 16'd55219, 16'd13224, 16'd21884, 16'd40002, 16'd39981, 16'd41065, 16'd24350, 16'd187, 16'd21899, 16'd51095, 16'd45650, 16'd10910, 16'd51122, 16'd32276, 16'd25134, 16'd58809, 16'd18702});
	test_expansion(128'h80738f960c8f51e1186b5795f70824b4, {16'd2915, 16'd12329, 16'd55864, 16'd34806, 16'd64080, 16'd41511, 16'd842, 16'd4781, 16'd30658, 16'd55532, 16'd2578, 16'd28752, 16'd14700, 16'd29836, 16'd17251, 16'd10656, 16'd43871, 16'd1016, 16'd59852, 16'd51665, 16'd44426, 16'd44228, 16'd61840, 16'd5161, 16'd53533, 16'd11880});
	test_expansion(128'heb3e118f78bccd178cef1bd4e61cb006, {16'd23358, 16'd31716, 16'd40917, 16'd32187, 16'd9487, 16'd20645, 16'd52674, 16'd16887, 16'd21521, 16'd759, 16'd63971, 16'd18555, 16'd5301, 16'd11814, 16'd33984, 16'd6068, 16'd51194, 16'd27893, 16'd50198, 16'd26798, 16'd25307, 16'd51760, 16'd2760, 16'd1714, 16'd30231, 16'd18072});
	test_expansion(128'hf09bbb48eb4cfbd39afe4cceea8ccf2f, {16'd53752, 16'd20460, 16'd60906, 16'd19212, 16'd9149, 16'd46888, 16'd1646, 16'd24631, 16'd24479, 16'd245, 16'd3648, 16'd7935, 16'd55302, 16'd53231, 16'd36916, 16'd9060, 16'd29086, 16'd38955, 16'd22856, 16'd5653, 16'd22352, 16'd2190, 16'd40657, 16'd64561, 16'd52735, 16'd23074});
	test_expansion(128'h6cab5c776cc95803179efa032e7ae615, {16'd63168, 16'd12316, 16'd13628, 16'd64101, 16'd49276, 16'd36304, 16'd50901, 16'd39419, 16'd53616, 16'd1758, 16'd44231, 16'd30171, 16'd56739, 16'd14934, 16'd22926, 16'd43619, 16'd369, 16'd27320, 16'd59027, 16'd48784, 16'd30522, 16'd36368, 16'd42356, 16'd30450, 16'd13386, 16'd40402});
	test_expansion(128'h76f355d0aae3c672892b641351c5e169, {16'd46665, 16'd39476, 16'd21988, 16'd64260, 16'd42027, 16'd45478, 16'd60322, 16'd55622, 16'd44277, 16'd6675, 16'd16525, 16'd65193, 16'd57695, 16'd53908, 16'd17472, 16'd17312, 16'd40035, 16'd53956, 16'd2179, 16'd12302, 16'd54646, 16'd28917, 16'd44028, 16'd13545, 16'd19551, 16'd4721});
	test_expansion(128'h0728a0bb369f3fe67acfc0d91fc6bda9, {16'd2995, 16'd55985, 16'd19056, 16'd59539, 16'd20219, 16'd40644, 16'd61855, 16'd3039, 16'd26996, 16'd64683, 16'd10655, 16'd34452, 16'd29365, 16'd40496, 16'd65147, 16'd3029, 16'd13979, 16'd13956, 16'd1197, 16'd51283, 16'd29174, 16'd13196, 16'd55689, 16'd64182, 16'd36756, 16'd33902});
	test_expansion(128'hfb1f192b4de19752be1c44c5a95c248e, {16'd60803, 16'd26430, 16'd51066, 16'd1905, 16'd62203, 16'd64599, 16'd17863, 16'd58476, 16'd50972, 16'd29927, 16'd32917, 16'd9410, 16'd41546, 16'd10277, 16'd10450, 16'd13626, 16'd25900, 16'd65504, 16'd17665, 16'd46352, 16'd64458, 16'd41011, 16'd8565, 16'd46301, 16'd46573, 16'd58468});
	test_expansion(128'h554c97d102690b5aaa22f93d3ba8bb68, {16'd64766, 16'd7499, 16'd40166, 16'd18681, 16'd37022, 16'd3879, 16'd17369, 16'd20708, 16'd63479, 16'd51571, 16'd12195, 16'd46058, 16'd2626, 16'd43376, 16'd1102, 16'd11474, 16'd7394, 16'd25241, 16'd62653, 16'd54398, 16'd59247, 16'd35246, 16'd14663, 16'd24851, 16'd4354, 16'd1639});
	test_expansion(128'h2468df4a12ec1af32a6c749319e77d76, {16'd16315, 16'd26546, 16'd2345, 16'd48188, 16'd20018, 16'd26607, 16'd31484, 16'd44549, 16'd6355, 16'd12502, 16'd26965, 16'd45828, 16'd27142, 16'd21720, 16'd6759, 16'd59697, 16'd51224, 16'd32723, 16'd44536, 16'd56695, 16'd20267, 16'd430, 16'd44187, 16'd11253, 16'd32194, 16'd29923});
	test_expansion(128'h2665a338b5c86ded5287480f2cb45fcb, {16'd59856, 16'd41209, 16'd57771, 16'd46291, 16'd8210, 16'd6211, 16'd2930, 16'd49706, 16'd29869, 16'd11307, 16'd44904, 16'd2295, 16'd36912, 16'd23610, 16'd12418, 16'd26968, 16'd55859, 16'd30739, 16'd33104, 16'd13001, 16'd62950, 16'd47327, 16'd919, 16'd21365, 16'd17047, 16'd20104});
	test_expansion(128'h0986f9c8dd95353e8e490599152fb679, {16'd29901, 16'd58257, 16'd53392, 16'd30686, 16'd40645, 16'd26702, 16'd17261, 16'd23109, 16'd38168, 16'd44977, 16'd57373, 16'd24890, 16'd39950, 16'd15681, 16'd10284, 16'd25905, 16'd2761, 16'd60273, 16'd57902, 16'd31514, 16'd2340, 16'd39961, 16'd41574, 16'd26654, 16'd26380, 16'd1489});
	test_expansion(128'hc6fad3fc5210d3dc680ab3952839df45, {16'd14667, 16'd30900, 16'd15177, 16'd45685, 16'd22239, 16'd44768, 16'd2859, 16'd57587, 16'd46238, 16'd24612, 16'd41994, 16'd45908, 16'd45767, 16'd60536, 16'd35130, 16'd566, 16'd9116, 16'd61132, 16'd10296, 16'd61456, 16'd24528, 16'd48812, 16'd44649, 16'd46484, 16'd20235, 16'd45688});
	test_expansion(128'h5e1c27224b60658fe8280f7602e1dcd2, {16'd60, 16'd1417, 16'd57992, 16'd22069, 16'd34019, 16'd58293, 16'd28212, 16'd43917, 16'd31529, 16'd48511, 16'd12465, 16'd36981, 16'd60801, 16'd5360, 16'd3450, 16'd39724, 16'd59412, 16'd34342, 16'd22961, 16'd16047, 16'd31094, 16'd46129, 16'd45816, 16'd37543, 16'd680, 16'd50764});
	test_expansion(128'h64f657c263659920cf4cca86bb1a2d70, {16'd9963, 16'd40170, 16'd27251, 16'd13945, 16'd42599, 16'd25417, 16'd47640, 16'd47188, 16'd9034, 16'd51163, 16'd12096, 16'd14247, 16'd17992, 16'd28082, 16'd58259, 16'd61091, 16'd52946, 16'd6747, 16'd28694, 16'd14712, 16'd43027, 16'd47671, 16'd33465, 16'd39279, 16'd57731, 16'd11230});
	test_expansion(128'h8a7b08088c7abfa67742a04d3b0f7ff1, {16'd34357, 16'd59600, 16'd23491, 16'd15225, 16'd39727, 16'd27972, 16'd3000, 16'd24769, 16'd31213, 16'd39336, 16'd9210, 16'd54929, 16'd34209, 16'd48677, 16'd48149, 16'd14817, 16'd3536, 16'd22430, 16'd32060, 16'd48702, 16'd9316, 16'd41397, 16'd19623, 16'd26891, 16'd18188, 16'd45294});
	test_expansion(128'h278109aecdd179d69ea804de4a4d86e5, {16'd3432, 16'd28094, 16'd20975, 16'd42545, 16'd46973, 16'd21587, 16'd33339, 16'd10046, 16'd8289, 16'd60800, 16'd45063, 16'd6552, 16'd30787, 16'd36840, 16'd23946, 16'd48951, 16'd58652, 16'd62497, 16'd37263, 16'd38626, 16'd48597, 16'd45308, 16'd18161, 16'd22099, 16'd18266, 16'd55998});
	test_expansion(128'hc96deff9db3d00d43cd8a4b100548960, {16'd28366, 16'd51135, 16'd41472, 16'd4047, 16'd49376, 16'd16626, 16'd43985, 16'd58316, 16'd54500, 16'd9842, 16'd48284, 16'd2937, 16'd12756, 16'd61995, 16'd42057, 16'd26472, 16'd44388, 16'd52866, 16'd43456, 16'd35407, 16'd56794, 16'd54623, 16'd62203, 16'd32651, 16'd43530, 16'd36917});
	test_expansion(128'h5f44dc9280975faf5b6ee7703802c241, {16'd4894, 16'd50407, 16'd36581, 16'd42306, 16'd18324, 16'd55782, 16'd15810, 16'd41175, 16'd18803, 16'd57717, 16'd37053, 16'd40638, 16'd40563, 16'd19071, 16'd33123, 16'd59915, 16'd18042, 16'd52963, 16'd20209, 16'd1021, 16'd23, 16'd30652, 16'd39113, 16'd29884, 16'd38072, 16'd24094});
	test_expansion(128'h6ae70cca3911d5d956a67d594a8de8ba, {16'd36247, 16'd1554, 16'd4848, 16'd25602, 16'd19664, 16'd30803, 16'd36515, 16'd14299, 16'd20175, 16'd92, 16'd60700, 16'd30656, 16'd4753, 16'd5201, 16'd29242, 16'd51932, 16'd60650, 16'd41295, 16'd18626, 16'd7771, 16'd50957, 16'd63472, 16'd47340, 16'd55290, 16'd29956, 16'd8512});
	test_expansion(128'h258e84d2a0e9d13708619fca721196d1, {16'd35920, 16'd24235, 16'd10188, 16'd62724, 16'd31589, 16'd35327, 16'd26332, 16'd59921, 16'd2501, 16'd37425, 16'd57828, 16'd36947, 16'd63862, 16'd38002, 16'd7757, 16'd10220, 16'd43005, 16'd1824, 16'd8902, 16'd11563, 16'd37082, 16'd51380, 16'd25496, 16'd17215, 16'd20864, 16'd51772});
	test_expansion(128'hd4d512e658473c6f313f224876fefbdc, {16'd27414, 16'd28713, 16'd37346, 16'd51732, 16'd24144, 16'd13329, 16'd12562, 16'd62420, 16'd57574, 16'd51912, 16'd58912, 16'd10025, 16'd31929, 16'd18046, 16'd2542, 16'd30505, 16'd20313, 16'd55893, 16'd8543, 16'd19914, 16'd11082, 16'd25615, 16'd63236, 16'd27312, 16'd2298, 16'd8748});
	test_expansion(128'h7d3d73330577e9742abf5849503ba679, {16'd41304, 16'd58468, 16'd46677, 16'd7950, 16'd50994, 16'd61983, 16'd28536, 16'd21312, 16'd9563, 16'd64932, 16'd15624, 16'd42870, 16'd25218, 16'd9261, 16'd25798, 16'd39257, 16'd36835, 16'd10448, 16'd34075, 16'd44184, 16'd51402, 16'd24023, 16'd44383, 16'd41506, 16'd49562, 16'd3814});
	test_expansion(128'h5450067e23763b75a2b0f23425617099, {16'd23366, 16'd18474, 16'd4070, 16'd35130, 16'd48702, 16'd51791, 16'd28715, 16'd44170, 16'd63038, 16'd13672, 16'd38061, 16'd61639, 16'd12335, 16'd52705, 16'd57460, 16'd6700, 16'd42972, 16'd8378, 16'd15354, 16'd4424, 16'd47294, 16'd56881, 16'd50764, 16'd26344, 16'd36639, 16'd25429});
	test_expansion(128'h7ea6480f6a1c5db62ca91a7b1c78b15a, {16'd26031, 16'd28689, 16'd61810, 16'd37192, 16'd40561, 16'd4123, 16'd52019, 16'd53774, 16'd6395, 16'd7785, 16'd14406, 16'd50490, 16'd52312, 16'd30846, 16'd27369, 16'd2903, 16'd58173, 16'd47058, 16'd54454, 16'd29038, 16'd44169, 16'd41585, 16'd18727, 16'd29431, 16'd19294, 16'd41300});
	test_expansion(128'h60ac298fcd840f2d45329fa1436311a9, {16'd37472, 16'd29179, 16'd40744, 16'd36269, 16'd43338, 16'd42698, 16'd27514, 16'd50458, 16'd22547, 16'd58727, 16'd57884, 16'd31142, 16'd34600, 16'd58324, 16'd269, 16'd17288, 16'd39036, 16'd36742, 16'd837, 16'd14680, 16'd12679, 16'd62640, 16'd17925, 16'd9075, 16'd18687, 16'd64784});
	test_expansion(128'h07172924933f3c607938dd68b0314c72, {16'd41580, 16'd3224, 16'd37450, 16'd16223, 16'd62311, 16'd15050, 16'd54608, 16'd52876, 16'd59942, 16'd5737, 16'd22757, 16'd27002, 16'd18904, 16'd37575, 16'd35834, 16'd57419, 16'd50347, 16'd2813, 16'd37957, 16'd34137, 16'd34750, 16'd1610, 16'd54995, 16'd52244, 16'd22042, 16'd16111});
	test_expansion(128'hb6eacaa2b7396703365cde129f9b2d8a, {16'd43234, 16'd34691, 16'd13529, 16'd26449, 16'd51163, 16'd49023, 16'd17328, 16'd53089, 16'd42725, 16'd48699, 16'd51943, 16'd19917, 16'd15172, 16'd1031, 16'd26863, 16'd5542, 16'd26013, 16'd1623, 16'd12197, 16'd17645, 16'd50238, 16'd35181, 16'd10578, 16'd1551, 16'd56394, 16'd55330});
	test_expansion(128'h9a01cceebc3b65afd0038c7667587837, {16'd41458, 16'd1083, 16'd32883, 16'd55563, 16'd31903, 16'd25552, 16'd14020, 16'd52467, 16'd21423, 16'd4190, 16'd51257, 16'd57280, 16'd23248, 16'd25795, 16'd32727, 16'd25826, 16'd23733, 16'd27129, 16'd54755, 16'd35909, 16'd25802, 16'd61687, 16'd41447, 16'd63523, 16'd43882, 16'd9717});
	test_expansion(128'h17bf896f672c1d6fa8ce0ed0fe5add70, {16'd52257, 16'd9530, 16'd37445, 16'd56410, 16'd55469, 16'd14091, 16'd48217, 16'd30940, 16'd432, 16'd52119, 16'd6192, 16'd8293, 16'd65253, 16'd28785, 16'd33143, 16'd9418, 16'd8615, 16'd50738, 16'd49498, 16'd36332, 16'd45412, 16'd41153, 16'd58272, 16'd49988, 16'd28608, 16'd8176});
	test_expansion(128'h736645b7b4c005c5179b03f1c0453b36, {16'd33649, 16'd59632, 16'd50121, 16'd47627, 16'd54773, 16'd31567, 16'd8163, 16'd33528, 16'd3718, 16'd45331, 16'd6337, 16'd42265, 16'd2837, 16'd59851, 16'd18951, 16'd56689, 16'd45265, 16'd32137, 16'd40399, 16'd42830, 16'd63907, 16'd40876, 16'd52420, 16'd9725, 16'd18072, 16'd28299});
	test_expansion(128'h502f2c407cfec8e163c5c90b37026c14, {16'd56005, 16'd34233, 16'd53544, 16'd10672, 16'd32097, 16'd59049, 16'd14802, 16'd55042, 16'd13427, 16'd34981, 16'd7798, 16'd34156, 16'd57378, 16'd43874, 16'd26417, 16'd5826, 16'd54068, 16'd59839, 16'd62925, 16'd47204, 16'd43802, 16'd2572, 16'd37305, 16'd12977, 16'd47726, 16'd44547});
	test_expansion(128'h8c73c39de262e7a0718306dac798882b, {16'd18082, 16'd29079, 16'd1458, 16'd33137, 16'd6123, 16'd54971, 16'd42344, 16'd16387, 16'd41391, 16'd57289, 16'd57341, 16'd44605, 16'd56122, 16'd1726, 16'd19595, 16'd64695, 16'd30904, 16'd25113, 16'd9766, 16'd13096, 16'd18743, 16'd45066, 16'd47374, 16'd20420, 16'd29880, 16'd11162});
	test_expansion(128'h6cae4c1444702d5af9b344587655ab5b, {16'd17134, 16'd9271, 16'd36643, 16'd36985, 16'd61366, 16'd48571, 16'd13469, 16'd17098, 16'd44663, 16'd3880, 16'd35045, 16'd40351, 16'd51907, 16'd15174, 16'd6649, 16'd42498, 16'd23789, 16'd25336, 16'd3867, 16'd5851, 16'd480, 16'd11426, 16'd46156, 16'd50211, 16'd41661, 16'd15972});
	test_expansion(128'ha97dc9a1941d8b3f8906ef2434b19fa1, {16'd50893, 16'd47335, 16'd54853, 16'd5215, 16'd47377, 16'd32355, 16'd50875, 16'd42140, 16'd54397, 16'd16056, 16'd65102, 16'd35547, 16'd32992, 16'd10765, 16'd44209, 16'd31804, 16'd56259, 16'd56039, 16'd31150, 16'd52439, 16'd64542, 16'd22212, 16'd51553, 16'd8149, 16'd18674, 16'd45148});
	test_expansion(128'h35769741978acc468f0a8ef527432225, {16'd61295, 16'd40077, 16'd62851, 16'd6642, 16'd14525, 16'd36132, 16'd22528, 16'd51613, 16'd57617, 16'd61473, 16'd34191, 16'd33051, 16'd45078, 16'd51642, 16'd61530, 16'd8523, 16'd63180, 16'd21364, 16'd61708, 16'd3300, 16'd35787, 16'd63788, 16'd39869, 16'd7367, 16'd4916, 16'd23583});
	test_expansion(128'hb5ba28cb6362503ffd95fd5b1e3aded3, {16'd49558, 16'd29618, 16'd40767, 16'd28798, 16'd32598, 16'd65499, 16'd49103, 16'd28571, 16'd57541, 16'd24537, 16'd14892, 16'd41002, 16'd27631, 16'd60042, 16'd63089, 16'd20777, 16'd40733, 16'd23905, 16'd30765, 16'd19016, 16'd22623, 16'd57099, 16'd56486, 16'd20966, 16'd13492, 16'd38135});
	test_expansion(128'h26a6bdc4e9b361a0aafb42ecde0be5e2, {16'd31489, 16'd17866, 16'd21604, 16'd36184, 16'd21868, 16'd47225, 16'd18662, 16'd3354, 16'd9257, 16'd8211, 16'd2089, 16'd63828, 16'd34024, 16'd13535, 16'd28783, 16'd39235, 16'd36506, 16'd34948, 16'd22790, 16'd53978, 16'd42005, 16'd38340, 16'd1069, 16'd57519, 16'd8217, 16'd23841});
	test_expansion(128'h62255ae877ed5160844e4d2bff77f941, {16'd1378, 16'd21120, 16'd33479, 16'd40003, 16'd6268, 16'd35498, 16'd37893, 16'd62454, 16'd6672, 16'd33215, 16'd22546, 16'd53783, 16'd1480, 16'd28737, 16'd34730, 16'd41650, 16'd16481, 16'd45526, 16'd38759, 16'd54538, 16'd13235, 16'd23961, 16'd51054, 16'd54244, 16'd15256, 16'd46569});
	test_expansion(128'h19cc4889f4c18760de39c53455cd49d3, {16'd24892, 16'd43252, 16'd54918, 16'd23953, 16'd58898, 16'd5045, 16'd10754, 16'd3794, 16'd59634, 16'd4215, 16'd4733, 16'd62551, 16'd3642, 16'd26368, 16'd43612, 16'd13249, 16'd45370, 16'd29712, 16'd15493, 16'd64073, 16'd7541, 16'd52769, 16'd55100, 16'd32724, 16'd35026, 16'd55807});
	test_expansion(128'h0eb86557711201b30305d91c8c253c59, {16'd43299, 16'd47781, 16'd7473, 16'd47716, 16'd59182, 16'd43708, 16'd35220, 16'd38495, 16'd48304, 16'd64352, 16'd27032, 16'd62100, 16'd28496, 16'd45437, 16'd30462, 16'd52326, 16'd63410, 16'd33396, 16'd44643, 16'd31333, 16'd4606, 16'd35447, 16'd26953, 16'd11774, 16'd32905, 16'd57695});
	test_expansion(128'hc202eba037a2c1820f8cc877837c33eb, {16'd60522, 16'd16365, 16'd62516, 16'd1595, 16'd52600, 16'd39096, 16'd36095, 16'd1509, 16'd22864, 16'd18199, 16'd38550, 16'd2050, 16'd61570, 16'd58260, 16'd11521, 16'd12956, 16'd13919, 16'd22497, 16'd12889, 16'd39175, 16'd18119, 16'd9217, 16'd36334, 16'd56838, 16'd22763, 16'd63499});
	test_expansion(128'h1b270db0e186d3156a4d542ed437e20d, {16'd63216, 16'd5149, 16'd48783, 16'd52867, 16'd42657, 16'd23825, 16'd27042, 16'd11876, 16'd61810, 16'd58962, 16'd25602, 16'd36275, 16'd29363, 16'd10575, 16'd1932, 16'd23573, 16'd13347, 16'd22776, 16'd28629, 16'd32569, 16'd61487, 16'd53899, 16'd54529, 16'd63956, 16'd14662, 16'd56952});
	test_expansion(128'h5616082ef352147a1ca72d8c9c257619, {16'd45538, 16'd21740, 16'd11785, 16'd11070, 16'd28326, 16'd50756, 16'd11893, 16'd11621, 16'd50331, 16'd18079, 16'd37498, 16'd26610, 16'd36787, 16'd49094, 16'd33342, 16'd61779, 16'd18080, 16'd3491, 16'd57988, 16'd22137, 16'd42942, 16'd53680, 16'd63154, 16'd33668, 16'd52415, 16'd32198});
	test_expansion(128'hcd94e27c53848b170e184cd92a8e07ea, {16'd18016, 16'd60666, 16'd52973, 16'd24691, 16'd8608, 16'd27555, 16'd61037, 16'd21242, 16'd21808, 16'd11418, 16'd39612, 16'd30051, 16'd44960, 16'd10166, 16'd40684, 16'd47509, 16'd6775, 16'd48640, 16'd11984, 16'd36545, 16'd9564, 16'd43285, 16'd25310, 16'd16601, 16'd63128, 16'd1979});
	test_expansion(128'h5e77810744068e0e2166dc7042ec3331, {16'd3375, 16'd42886, 16'd58504, 16'd59430, 16'd50812, 16'd60760, 16'd33456, 16'd62679, 16'd14435, 16'd44622, 16'd46386, 16'd61173, 16'd51232, 16'd56131, 16'd7562, 16'd59043, 16'd34978, 16'd56331, 16'd8924, 16'd3613, 16'd35332, 16'd58821, 16'd48686, 16'd33659, 16'd59931, 16'd57717});
	test_expansion(128'hb7c27e7612e467fa4fbfce6a3c26f1d8, {16'd17075, 16'd20764, 16'd23020, 16'd26757, 16'd20541, 16'd52726, 16'd13874, 16'd49484, 16'd36600, 16'd46207, 16'd23191, 16'd27496, 16'd41230, 16'd35705, 16'd13743, 16'd41180, 16'd38966, 16'd38824, 16'd5042, 16'd38898, 16'd49851, 16'd8365, 16'd25383, 16'd45201, 16'd30325, 16'd26130});
	test_expansion(128'h06729ea9d6f73d657b3694d14f40ac36, {16'd32814, 16'd17567, 16'd54456, 16'd36398, 16'd6351, 16'd16174, 16'd10225, 16'd1791, 16'd52982, 16'd25893, 16'd4272, 16'd277, 16'd36879, 16'd17209, 16'd44493, 16'd23951, 16'd8767, 16'd19927, 16'd21400, 16'd61039, 16'd32807, 16'd55688, 16'd39553, 16'd60923, 16'd2991, 16'd27843});
	test_expansion(128'h5ec9860adfa1563c59ad9f25f624ba14, {16'd37874, 16'd61157, 16'd53773, 16'd5125, 16'd13285, 16'd32457, 16'd64208, 16'd42578, 16'd35203, 16'd29640, 16'd44867, 16'd16585, 16'd48544, 16'd6539, 16'd48786, 16'd37193, 16'd17853, 16'd20321, 16'd40029, 16'd8642, 16'd53262, 16'd55288, 16'd259, 16'd52679, 16'd47910, 16'd65244});
	test_expansion(128'hdfb67fb4ba23fd98c5517411692c7a96, {16'd34556, 16'd64840, 16'd25556, 16'd38764, 16'd22935, 16'd38637, 16'd43037, 16'd58337, 16'd11752, 16'd39534, 16'd20550, 16'd6996, 16'd24353, 16'd7093, 16'd46687, 16'd29851, 16'd61548, 16'd5774, 16'd50015, 16'd16737, 16'd41173, 16'd31849, 16'd45804, 16'd54381, 16'd30868, 16'd59899});
	test_expansion(128'h4a30dec2d813bb66ffe97c38bd969f15, {16'd46000, 16'd18735, 16'd37201, 16'd39406, 16'd52089, 16'd40647, 16'd63839, 16'd15631, 16'd51074, 16'd39723, 16'd45562, 16'd37129, 16'd51326, 16'd37115, 16'd51489, 16'd37537, 16'd48326, 16'd55188, 16'd30031, 16'd61557, 16'd11310, 16'd6041, 16'd34779, 16'd30577, 16'd48428, 16'd5082});
	test_expansion(128'hd246c0a5b80e5c921420ab1ca6965508, {16'd9075, 16'd26642, 16'd61614, 16'd8603, 16'd40040, 16'd11090, 16'd7475, 16'd38950, 16'd51099, 16'd62497, 16'd18217, 16'd19584, 16'd35327, 16'd49685, 16'd8137, 16'd32061, 16'd13421, 16'd42063, 16'd15285, 16'd3830, 16'd42588, 16'd43147, 16'd22776, 16'd58409, 16'd35741, 16'd45668});
	test_expansion(128'ha3c39d3c14be613419f941d369962d25, {16'd5457, 16'd41548, 16'd47567, 16'd48552, 16'd57454, 16'd64887, 16'd51492, 16'd33516, 16'd7800, 16'd53917, 16'd36598, 16'd34943, 16'd61367, 16'd21138, 16'd40610, 16'd22179, 16'd5385, 16'd48411, 16'd1701, 16'd3744, 16'd54203, 16'd47139, 16'd26348, 16'd24885, 16'd9771, 16'd47053});
	test_expansion(128'h2494c3fbb0f4b99d0710577531638ec6, {16'd27726, 16'd41857, 16'd21602, 16'd65018, 16'd26208, 16'd13551, 16'd21571, 16'd62074, 16'd43451, 16'd19077, 16'd59965, 16'd35330, 16'd8883, 16'd30140, 16'd62331, 16'd16928, 16'd64544, 16'd20150, 16'd12784, 16'd60156, 16'd28188, 16'd4223, 16'd39294, 16'd44335, 16'd26766, 16'd22763});
	test_expansion(128'h6369f166fbb353d792079f296908d587, {16'd20303, 16'd41980, 16'd26742, 16'd37182, 16'd16331, 16'd40921, 16'd8003, 16'd42912, 16'd51643, 16'd37854, 16'd2725, 16'd2390, 16'd48846, 16'd33055, 16'd22285, 16'd10509, 16'd12088, 16'd13900, 16'd30257, 16'd46998, 16'd46795, 16'd30003, 16'd12097, 16'd17276, 16'd48601, 16'd34360});
	test_expansion(128'hd1ab2b82d807a48582c5ab9f9e12f1b9, {16'd24680, 16'd49587, 16'd27113, 16'd54242, 16'd40844, 16'd31125, 16'd63356, 16'd63427, 16'd60489, 16'd16931, 16'd47949, 16'd25668, 16'd60361, 16'd20849, 16'd61747, 16'd47547, 16'd54508, 16'd26848, 16'd4546, 16'd3719, 16'd50656, 16'd26640, 16'd5529, 16'd23765, 16'd2830, 16'd34336});
	test_expansion(128'h2dd27a256a59a4d2fb8a9871fe36b418, {16'd42348, 16'd39466, 16'd45038, 16'd29657, 16'd23226, 16'd33570, 16'd52398, 16'd12605, 16'd47017, 16'd55462, 16'd49137, 16'd33999, 16'd25212, 16'd54930, 16'd61499, 16'd17064, 16'd48103, 16'd9230, 16'd17755, 16'd23065, 16'd39290, 16'd8161, 16'd4516, 16'd26749, 16'd29808, 16'd37971});
	test_expansion(128'he967b679c197540d59e8cf32530003ed, {16'd23716, 16'd7321, 16'd16571, 16'd21084, 16'd59299, 16'd38893, 16'd50542, 16'd28067, 16'd41855, 16'd41831, 16'd21777, 16'd6575, 16'd2159, 16'd6149, 16'd47849, 16'd43032, 16'd6337, 16'd166, 16'd50518, 16'd39219, 16'd6218, 16'd18270, 16'd9160, 16'd4194, 16'd64054, 16'd28888});
	test_expansion(128'hf77e01bc8c8beeef9c4544cfb0cf88ba, {16'd60583, 16'd18520, 16'd47122, 16'd62380, 16'd24594, 16'd21636, 16'd7964, 16'd60475, 16'd48426, 16'd633, 16'd35386, 16'd28275, 16'd25937, 16'd34610, 16'd44692, 16'd43418, 16'd31247, 16'd64322, 16'd64080, 16'd4062, 16'd31592, 16'd4092, 16'd60214, 16'd15527, 16'd23483, 16'd389});
	test_expansion(128'hacf75d10ee75b32b223306c375bb7b41, {16'd8039, 16'd27861, 16'd55424, 16'd8707, 16'd13230, 16'd27287, 16'd49322, 16'd28530, 16'd55103, 16'd59537, 16'd53611, 16'd29012, 16'd64929, 16'd8737, 16'd51099, 16'd18737, 16'd36445, 16'd49888, 16'd41148, 16'd37298, 16'd41033, 16'd8875, 16'd23329, 16'd43297, 16'd45730, 16'd62301});
	test_expansion(128'hf89886a0d3a011df6fa82121fd8804b4, {16'd31892, 16'd48914, 16'd14621, 16'd56399, 16'd9737, 16'd4043, 16'd56819, 16'd45739, 16'd43897, 16'd10811, 16'd39049, 16'd43665, 16'd63191, 16'd64779, 16'd49525, 16'd20741, 16'd26259, 16'd12432, 16'd25827, 16'd18406, 16'd30956, 16'd15596, 16'd11292, 16'd22429, 16'd9128, 16'd27075});
	test_expansion(128'h25143b42fabfb7db5eed985a8cbb98d8, {16'd10490, 16'd3463, 16'd45986, 16'd41357, 16'd21454, 16'd23511, 16'd40174, 16'd28301, 16'd47604, 16'd62704, 16'd25283, 16'd43624, 16'd6412, 16'd34627, 16'd7197, 16'd10611, 16'd14802, 16'd3489, 16'd33869, 16'd36882, 16'd43824, 16'd47430, 16'd44733, 16'd18034, 16'd26313, 16'd30852});
	test_expansion(128'h55788c58902c41d1f6183f752aa893bb, {16'd23853, 16'd7317, 16'd23733, 16'd12533, 16'd29389, 16'd20775, 16'd8441, 16'd2810, 16'd60960, 16'd47785, 16'd7605, 16'd14330, 16'd65531, 16'd42149, 16'd15698, 16'd62214, 16'd19166, 16'd27436, 16'd26845, 16'd52017, 16'd10176, 16'd2076, 16'd61850, 16'd46239, 16'd29146, 16'd32173});
	test_expansion(128'h5b17ffee0853aeef9f48d10d1bc7a4b3, {16'd31137, 16'd46345, 16'd35630, 16'd1432, 16'd40122, 16'd21518, 16'd54023, 16'd13069, 16'd60729, 16'd50719, 16'd62120, 16'd7261, 16'd35007, 16'd1233, 16'd31569, 16'd34008, 16'd46287, 16'd46536, 16'd63472, 16'd43748, 16'd29716, 16'd31408, 16'd49188, 16'd8345, 16'd45711, 16'd37514});
	test_expansion(128'h8b31dd6e40586b3b321927303290a99a, {16'd24555, 16'd23687, 16'd30437, 16'd42806, 16'd4532, 16'd17581, 16'd18621, 16'd61933, 16'd53000, 16'd22002, 16'd7049, 16'd21836, 16'd3536, 16'd20247, 16'd64309, 16'd12096, 16'd14887, 16'd10576, 16'd25028, 16'd40018, 16'd47710, 16'd52029, 16'd54955, 16'd56372, 16'd42724, 16'd22129});
	test_expansion(128'h7382ab1583a259fea3ca2b545d715127, {16'd43033, 16'd19326, 16'd23393, 16'd56747, 16'd44839, 16'd39683, 16'd22473, 16'd20904, 16'd26335, 16'd44634, 16'd51787, 16'd24620, 16'd26079, 16'd18466, 16'd40123, 16'd33009, 16'd14569, 16'd2714, 16'd306, 16'd27573, 16'd26268, 16'd23861, 16'd4881, 16'd10248, 16'd60186, 16'd12241});
	test_expansion(128'h37e8877c05f8c9eaea1a8ee7ae39ca34, {16'd33078, 16'd63637, 16'd36936, 16'd52442, 16'd7813, 16'd53331, 16'd30560, 16'd19265, 16'd41595, 16'd25429, 16'd61836, 16'd24483, 16'd295, 16'd57296, 16'd26828, 16'd29071, 16'd38677, 16'd46639, 16'd24793, 16'd12574, 16'd21862, 16'd26977, 16'd40281, 16'd27047, 16'd13394, 16'd7455});
	test_expansion(128'hb071d7a1eeb1c6fe57485b889b383a34, {16'd3767, 16'd13580, 16'd55742, 16'd14539, 16'd57019, 16'd54600, 16'd36287, 16'd65161, 16'd38378, 16'd7436, 16'd51755, 16'd8143, 16'd39699, 16'd34306, 16'd10333, 16'd43514, 16'd28918, 16'd56952, 16'd43086, 16'd36162, 16'd10199, 16'd35563, 16'd47728, 16'd44518, 16'd51600, 16'd35013});
	test_expansion(128'h9ca71f88dcbfbe7c7e6da9e824c33a68, {16'd25438, 16'd46575, 16'd54874, 16'd49478, 16'd62653, 16'd27424, 16'd17354, 16'd7825, 16'd9655, 16'd5672, 16'd11865, 16'd24496, 16'd4301, 16'd49808, 16'd36063, 16'd64410, 16'd53410, 16'd18945, 16'd6319, 16'd32930, 16'd43904, 16'd9145, 16'd60573, 16'd26511, 16'd1474, 16'd17758});
	test_expansion(128'h0b91896f52a6d850a490d98407691c70, {16'd54826, 16'd34712, 16'd35980, 16'd22123, 16'd9684, 16'd29292, 16'd15315, 16'd41082, 16'd50747, 16'd48414, 16'd50239, 16'd11577, 16'd34688, 16'd28872, 16'd23093, 16'd7146, 16'd47504, 16'd23050, 16'd6682, 16'd58733, 16'd37266, 16'd17750, 16'd12933, 16'd57847, 16'd35793, 16'd38998});
	test_expansion(128'h0c69db51d484624258cfcdafe0dd5df4, {16'd57396, 16'd15833, 16'd31240, 16'd11019, 16'd28360, 16'd24457, 16'd52592, 16'd57538, 16'd34013, 16'd48592, 16'd53220, 16'd36820, 16'd31807, 16'd27580, 16'd32213, 16'd10885, 16'd10559, 16'd27188, 16'd43800, 16'd25493, 16'd38373, 16'd315, 16'd51258, 16'd5483, 16'd14725, 16'd31644});
	test_expansion(128'hae7589132196ef73120c7f97834759f4, {16'd59139, 16'd52562, 16'd47510, 16'd53928, 16'd2367, 16'd9393, 16'd45937, 16'd21348, 16'd25193, 16'd38520, 16'd48180, 16'd17515, 16'd25044, 16'd29137, 16'd47665, 16'd32593, 16'd62227, 16'd7308, 16'd11170, 16'd53111, 16'd58843, 16'd51711, 16'd8746, 16'd23271, 16'd10261, 16'd27547});
	test_expansion(128'h1a5a69a482ccc9491550b7d86a9f5579, {16'd35554, 16'd50783, 16'd50058, 16'd28665, 16'd31371, 16'd61334, 16'd10313, 16'd33105, 16'd56670, 16'd34701, 16'd49711, 16'd64793, 16'd6442, 16'd38430, 16'd44606, 16'd36347, 16'd63280, 16'd30923, 16'd19721, 16'd39928, 16'd22163, 16'd62636, 16'd44653, 16'd43564, 16'd8905, 16'd16228});
	test_expansion(128'h9c5f120aee348ed5b98f9defba590afd, {16'd31602, 16'd63504, 16'd38490, 16'd28373, 16'd4139, 16'd23094, 16'd24978, 16'd53516, 16'd19423, 16'd19160, 16'd42500, 16'd42476, 16'd60894, 16'd20487, 16'd35655, 16'd4020, 16'd30491, 16'd27475, 16'd32783, 16'd48715, 16'd15403, 16'd21425, 16'd40948, 16'd14882, 16'd31834, 16'd11993});
	test_expansion(128'hc482f3bb4fd81d476c395472cdefa167, {16'd56389, 16'd14905, 16'd14821, 16'd48135, 16'd55873, 16'd42572, 16'd45663, 16'd36085, 16'd42045, 16'd14487, 16'd29968, 16'd51318, 16'd54076, 16'd39000, 16'd65143, 16'd10249, 16'd10148, 16'd9743, 16'd64784, 16'd13220, 16'd42029, 16'd8588, 16'd45488, 16'd43459, 16'd38996, 16'd7043});
	test_expansion(128'hf3f8afb0d0f7cb33c1f5d7314c074c91, {16'd43144, 16'd4251, 16'd63772, 16'd51381, 16'd58571, 16'd48160, 16'd31209, 16'd10624, 16'd2737, 16'd8719, 16'd27779, 16'd31971, 16'd6138, 16'd30413, 16'd63602, 16'd11563, 16'd10174, 16'd20332, 16'd37395, 16'd36952, 16'd50074, 16'd29445, 16'd47058, 16'd62542, 16'd36369, 16'd20437});
	test_expansion(128'h5075f5a737ec9ab7f8ddc736f3a8eb40, {16'd50565, 16'd65249, 16'd24999, 16'd48219, 16'd20109, 16'd43721, 16'd63495, 16'd20963, 16'd54869, 16'd19417, 16'd1885, 16'd42352, 16'd7608, 16'd36372, 16'd9841, 16'd11276, 16'd58326, 16'd14179, 16'd27186, 16'd27166, 16'd54589, 16'd34094, 16'd59560, 16'd58647, 16'd33423, 16'd28391});
	test_expansion(128'h70300e80a4dd119caacc33ad5909fca6, {16'd62211, 16'd7748, 16'd50153, 16'd18666, 16'd48373, 16'd35892, 16'd43357, 16'd12721, 16'd32141, 16'd1945, 16'd64410, 16'd38813, 16'd23780, 16'd19424, 16'd35617, 16'd17844, 16'd26710, 16'd17513, 16'd26581, 16'd3054, 16'd49748, 16'd22282, 16'd44885, 16'd53291, 16'd64018, 16'd21446});
	test_expansion(128'h02d3f7e6a327e697186ff61df46c6ab0, {16'd16308, 16'd42481, 16'd24634, 16'd31198, 16'd26935, 16'd62535, 16'd46541, 16'd58216, 16'd36103, 16'd4372, 16'd22052, 16'd58390, 16'd33494, 16'd49774, 16'd64552, 16'd31590, 16'd49318, 16'd63475, 16'd14653, 16'd35146, 16'd44176, 16'd11751, 16'd24793, 16'd49047, 16'd46288, 16'd30801});
	test_expansion(128'hb1a148459649a1d0f12eba216fdac2b8, {16'd15021, 16'd54163, 16'd27666, 16'd57435, 16'd59376, 16'd7512, 16'd50856, 16'd36367, 16'd62179, 16'd27860, 16'd39443, 16'd57715, 16'd23847, 16'd7459, 16'd3051, 16'd50395, 16'd16490, 16'd52159, 16'd30174, 16'd15670, 16'd46477, 16'd2812, 16'd61815, 16'd42646, 16'd34590, 16'd52577});
	test_expansion(128'hca95b1b1a6a64f329e89fac998a81a67, {16'd891, 16'd29140, 16'd22982, 16'd21141, 16'd34074, 16'd40472, 16'd24034, 16'd52611, 16'd62390, 16'd13744, 16'd49485, 16'd10754, 16'd5381, 16'd63380, 16'd8576, 16'd45074, 16'd57371, 16'd18448, 16'd11557, 16'd42046, 16'd53234, 16'd21926, 16'd29416, 16'd16874, 16'd48329, 16'd46090});
	test_expansion(128'hc99f80aafd731a761d61a2cdcec5366a, {16'd52631, 16'd46102, 16'd10770, 16'd37858, 16'd65024, 16'd36201, 16'd13046, 16'd62811, 16'd36160, 16'd25788, 16'd11734, 16'd3142, 16'd15758, 16'd34470, 16'd35639, 16'd15089, 16'd20178, 16'd38632, 16'd4749, 16'd53936, 16'd57242, 16'd23304, 16'd9638, 16'd23742, 16'd51752, 16'd30889});
	test_expansion(128'he6fb0d54ad9ebfd9d6250560530f0c9d, {16'd34917, 16'd26194, 16'd9514, 16'd20777, 16'd37496, 16'd18199, 16'd40937, 16'd38005, 16'd16414, 16'd2786, 16'd61240, 16'd63858, 16'd2308, 16'd17017, 16'd64910, 16'd35509, 16'd34855, 16'd5137, 16'd17715, 16'd13508, 16'd32598, 16'd13928, 16'd42400, 16'd12971, 16'd21984, 16'd23385});
	test_expansion(128'h8f78515d88340c790a3c6ab014d75242, {16'd17854, 16'd63038, 16'd41503, 16'd43896, 16'd36183, 16'd16346, 16'd55538, 16'd20218, 16'd42997, 16'd2114, 16'd15314, 16'd43260, 16'd48920, 16'd64759, 16'd51412, 16'd47677, 16'd40335, 16'd56796, 16'd8561, 16'd29925, 16'd56266, 16'd41244, 16'd16517, 16'd16153, 16'd19248, 16'd19664});
	test_expansion(128'h201d87d6511ff51874575148f6816c85, {16'd24885, 16'd31151, 16'd7796, 16'd21341, 16'd6577, 16'd61482, 16'd50035, 16'd60196, 16'd5118, 16'd51486, 16'd5352, 16'd27708, 16'd58501, 16'd26776, 16'd45695, 16'd59277, 16'd21750, 16'd46154, 16'd62530, 16'd37454, 16'd58139, 16'd19799, 16'd29184, 16'd61272, 16'd27394, 16'd31278});
	test_expansion(128'h70b916eaeaf4678c13cf203fa41b44c0, {16'd22657, 16'd46872, 16'd6725, 16'd17627, 16'd53204, 16'd16423, 16'd37861, 16'd44752, 16'd59393, 16'd16429, 16'd28410, 16'd7652, 16'd34242, 16'd24615, 16'd65377, 16'd49593, 16'd49123, 16'd24499, 16'd64428, 16'd54453, 16'd17565, 16'd65132, 16'd31436, 16'd9742, 16'd15226, 16'd15326});
	test_expansion(128'h5343851a218c04b5c3cd31524ce537ff, {16'd53818, 16'd2795, 16'd31482, 16'd31861, 16'd37304, 16'd8056, 16'd48828, 16'd31314, 16'd34769, 16'd6536, 16'd2703, 16'd31988, 16'd50212, 16'd65226, 16'd46920, 16'd28903, 16'd48159, 16'd4260, 16'd27279, 16'd33520, 16'd2744, 16'd35960, 16'd58517, 16'd61142, 16'd43570, 16'd56171});
	test_expansion(128'he5e558296e266d5fcebd5a5c493a0f13, {16'd23704, 16'd7203, 16'd32524, 16'd27404, 16'd65442, 16'd37643, 16'd59744, 16'd9738, 16'd7060, 16'd40102, 16'd38301, 16'd45008, 16'd20865, 16'd58299, 16'd63175, 16'd31213, 16'd52673, 16'd16435, 16'd59642, 16'd16251, 16'd34025, 16'd54505, 16'd26473, 16'd45856, 16'd9948, 16'd15100});
	test_expansion(128'h406e2ea9cd9fc184649faf0db1119402, {16'd9038, 16'd9692, 16'd33609, 16'd19117, 16'd16037, 16'd30507, 16'd53498, 16'd56828, 16'd2668, 16'd56896, 16'd54422, 16'd57874, 16'd58837, 16'd58796, 16'd22773, 16'd9015, 16'd50901, 16'd14515, 16'd3951, 16'd36673, 16'd4906, 16'd60649, 16'd11418, 16'd50079, 16'd58940, 16'd14485});
	test_expansion(128'h5ecbfe3de873091e1b707519cfa9d378, {16'd30780, 16'd56728, 16'd22212, 16'd11681, 16'd32794, 16'd18568, 16'd42421, 16'd27058, 16'd42692, 16'd47888, 16'd52173, 16'd13116, 16'd46532, 16'd5950, 16'd20230, 16'd26179, 16'd37266, 16'd51174, 16'd36066, 16'd9524, 16'd44902, 16'd29100, 16'd212, 16'd34750, 16'd50785, 16'd59591});
	test_expansion(128'h0b4b8eb397e21fceaf51205003dea46c, {16'd40963, 16'd49810, 16'd9493, 16'd47683, 16'd7177, 16'd584, 16'd57568, 16'd52663, 16'd25303, 16'd53795, 16'd6363, 16'd5590, 16'd15280, 16'd38605, 16'd9102, 16'd36328, 16'd6061, 16'd60910, 16'd22194, 16'd38721, 16'd28201, 16'd35139, 16'd41359, 16'd21101, 16'd11079, 16'd19393});
	test_expansion(128'h8456af1d5913bcb3ac53ca54eee787c5, {16'd63032, 16'd59566, 16'd35150, 16'd18197, 16'd13141, 16'd63835, 16'd50126, 16'd3419, 16'd54984, 16'd15950, 16'd38851, 16'd34811, 16'd12979, 16'd49011, 16'd35989, 16'd55058, 16'd60194, 16'd6743, 16'd46204, 16'd61393, 16'd46046, 16'd28392, 16'd39916, 16'd43700, 16'd21240, 16'd16226});
	test_expansion(128'h1abc07121bb678ef062d96696205cefd, {16'd55558, 16'd10129, 16'd52979, 16'd17178, 16'd62580, 16'd50978, 16'd64679, 16'd38264, 16'd17106, 16'd27597, 16'd32752, 16'd47712, 16'd10170, 16'd3902, 16'd32273, 16'd13909, 16'd55234, 16'd26828, 16'd10649, 16'd52818, 16'd15105, 16'd54000, 16'd1961, 16'd36568, 16'd34861, 16'd45804});
	test_expansion(128'h6607b7951c93566f0cdd1929b95a7f55, {16'd62848, 16'd26075, 16'd45693, 16'd3377, 16'd42753, 16'd12545, 16'd24545, 16'd2333, 16'd56724, 16'd55017, 16'd48368, 16'd2599, 16'd15757, 16'd50099, 16'd4103, 16'd12709, 16'd28352, 16'd14668, 16'd7037, 16'd51640, 16'd51051, 16'd63715, 16'd57739, 16'd59411, 16'd51044, 16'd29760});
	test_expansion(128'h21fa8c76ad47ca02a09dd2a469327fd3, {16'd8925, 16'd42745, 16'd29872, 16'd65063, 16'd53462, 16'd19660, 16'd33737, 16'd11644, 16'd24442, 16'd7740, 16'd61265, 16'd5899, 16'd13983, 16'd62696, 16'd51499, 16'd63168, 16'd38641, 16'd53024, 16'd62595, 16'd8618, 16'd10703, 16'd6199, 16'd64582, 16'd37988, 16'd10860, 16'd22098});
	test_expansion(128'h136ffb30aba34b151ed15f52f4d9ecce, {16'd21908, 16'd30317, 16'd61540, 16'd64247, 16'd24794, 16'd46223, 16'd65316, 16'd36676, 16'd10839, 16'd56860, 16'd15752, 16'd57358, 16'd27115, 16'd45994, 16'd55461, 16'd24536, 16'd35543, 16'd3018, 16'd18593, 16'd21787, 16'd26942, 16'd63733, 16'd16833, 16'd46275, 16'd65041, 16'd64761});
	test_expansion(128'hc3e1456468bd4aae102b378e2a834106, {16'd3096, 16'd40047, 16'd36710, 16'd49813, 16'd58830, 16'd15461, 16'd48843, 16'd12920, 16'd36855, 16'd9078, 16'd6807, 16'd51695, 16'd41051, 16'd44435, 16'd29, 16'd53448, 16'd18182, 16'd52003, 16'd32281, 16'd20285, 16'd26757, 16'd27544, 16'd59204, 16'd4239, 16'd48113, 16'd2969});
	test_expansion(128'h3add44a19060159ac77a915bb5e42477, {16'd15300, 16'd40377, 16'd41528, 16'd30773, 16'd63115, 16'd637, 16'd37253, 16'd62963, 16'd62815, 16'd14761, 16'd17119, 16'd2533, 16'd21125, 16'd24142, 16'd44280, 16'd45857, 16'd1472, 16'd40633, 16'd25820, 16'd17152, 16'd25353, 16'd42171, 16'd39385, 16'd6951, 16'd20062, 16'd48303});
	test_expansion(128'hc54195d9f2ca5fe665c18548e972e1d8, {16'd63818, 16'd22098, 16'd9958, 16'd59320, 16'd21996, 16'd29710, 16'd12209, 16'd49259, 16'd13013, 16'd22226, 16'd38097, 16'd63142, 16'd17862, 16'd23178, 16'd55872, 16'd10408, 16'd40300, 16'd23610, 16'd48747, 16'd16354, 16'd46258, 16'd18915, 16'd44922, 16'd53472, 16'd60936, 16'd64703});
	test_expansion(128'h78f19d3940624d72b5ae6142220b74d2, {16'd18685, 16'd1140, 16'd44580, 16'd36789, 16'd31674, 16'd64533, 16'd50804, 16'd40872, 16'd8463, 16'd64602, 16'd43324, 16'd62205, 16'd44912, 16'd63208, 16'd24153, 16'd13953, 16'd58524, 16'd30171, 16'd12026, 16'd9321, 16'd44578, 16'd35415, 16'd60800, 16'd4891, 16'd17503, 16'd62287});
	test_expansion(128'h27f0935e4ce9068c4a83d061da91037e, {16'd39869, 16'd64954, 16'd41789, 16'd56895, 16'd8972, 16'd30650, 16'd45271, 16'd8825, 16'd63382, 16'd65475, 16'd35168, 16'd29382, 16'd36096, 16'd50279, 16'd3562, 16'd50856, 16'd11388, 16'd25694, 16'd16822, 16'd23014, 16'd34017, 16'd53283, 16'd21122, 16'd17479, 16'd43642, 16'd7074});
	test_expansion(128'hd87040f6a8f2a426206bb7a44c32913e, {16'd38310, 16'd50754, 16'd54977, 16'd40013, 16'd27390, 16'd34688, 16'd38581, 16'd55620, 16'd14913, 16'd4445, 16'd62095, 16'd64696, 16'd52670, 16'd43138, 16'd53506, 16'd39614, 16'd13818, 16'd7756, 16'd25888, 16'd49238, 16'd40028, 16'd23202, 16'd28785, 16'd24801, 16'd27113, 16'd3131});
	test_expansion(128'h7f112329ab5a2be99097b32c6af23a86, {16'd3348, 16'd10928, 16'd22844, 16'd33096, 16'd55592, 16'd65025, 16'd21251, 16'd17540, 16'd6913, 16'd42682, 16'd48071, 16'd41492, 16'd61434, 16'd35400, 16'd37603, 16'd38707, 16'd17130, 16'd2548, 16'd35013, 16'd42317, 16'd54316, 16'd14018, 16'd61217, 16'd15675, 16'd6227, 16'd33411});
	test_expansion(128'h34a09db4d5ce2b5093cfd7996eefceda, {16'd35686, 16'd21687, 16'd60895, 16'd23979, 16'd38446, 16'd6832, 16'd24941, 16'd61246, 16'd57627, 16'd18950, 16'd19264, 16'd41519, 16'd56349, 16'd33830, 16'd15644, 16'd29483, 16'd19183, 16'd22611, 16'd5971, 16'd22700, 16'd40163, 16'd49887, 16'd36497, 16'd7280, 16'd2079, 16'd2469});
	test_expansion(128'h4861d5470316c1e88451fe98a60ca8e2, {16'd14178, 16'd10894, 16'd7436, 16'd60059, 16'd35870, 16'd59164, 16'd23428, 16'd27263, 16'd63793, 16'd49048, 16'd2856, 16'd56117, 16'd56841, 16'd39801, 16'd64383, 16'd47398, 16'd3573, 16'd59932, 16'd58347, 16'd49240, 16'd35049, 16'd5495, 16'd65387, 16'd29243, 16'd51950, 16'd2181});
	test_expansion(128'h1302bc52ff7bbe1bbc4aa378464cee30, {16'd38855, 16'd4182, 16'd41591, 16'd18310, 16'd56028, 16'd2979, 16'd38036, 16'd8370, 16'd55083, 16'd6188, 16'd3206, 16'd61714, 16'd48738, 16'd59452, 16'd3358, 16'd14720, 16'd62341, 16'd54359, 16'd21033, 16'd19522, 16'd62787, 16'd53711, 16'd61289, 16'd19669, 16'd24984, 16'd41928});
	test_expansion(128'h3844df4be6e7faaa7be7dea8cf4a28bf, {16'd8914, 16'd27780, 16'd7950, 16'd38134, 16'd23021, 16'd37022, 16'd12503, 16'd19359, 16'd876, 16'd43017, 16'd4793, 16'd15049, 16'd18701, 16'd25465, 16'd53830, 16'd48003, 16'd39099, 16'd45473, 16'd55020, 16'd55112, 16'd4676, 16'd19598, 16'd15949, 16'd32856, 16'd34885, 16'd57658});
	test_expansion(128'he52861725d477c27dc6c67210cdb2067, {16'd63507, 16'd60591, 16'd26720, 16'd19402, 16'd29495, 16'd41857, 16'd37327, 16'd22435, 16'd15286, 16'd13687, 16'd23640, 16'd23081, 16'd35021, 16'd1819, 16'd6101, 16'd26905, 16'd41233, 16'd12215, 16'd11632, 16'd34851, 16'd57356, 16'd8858, 16'd7964, 16'd32348, 16'd1441, 16'd14412});
	test_expansion(128'h18af4a6bc6c6bbc5a47b7df0d354b8f1, {16'd37055, 16'd16956, 16'd3677, 16'd42763, 16'd32914, 16'd3858, 16'd55147, 16'd44735, 16'd5375, 16'd50628, 16'd31758, 16'd10959, 16'd9333, 16'd36235, 16'd6872, 16'd31550, 16'd56396, 16'd58207, 16'd52324, 16'd42905, 16'd4929, 16'd36224, 16'd63900, 16'd48663, 16'd3615, 16'd44547});
	test_expansion(128'h03b6458a4910df6077582995597a2b79, {16'd16129, 16'd5865, 16'd20017, 16'd38691, 16'd53743, 16'd10955, 16'd64868, 16'd35968, 16'd24097, 16'd16988, 16'd44047, 16'd6870, 16'd48885, 16'd14356, 16'd23915, 16'd36457, 16'd6021, 16'd59135, 16'd46789, 16'd48348, 16'd30735, 16'd8863, 16'd56083, 16'd20675, 16'd12287, 16'd8866});
	test_expansion(128'h891a68bd88963c05342691ade8bad1d8, {16'd48397, 16'd17680, 16'd24701, 16'd58049, 16'd27074, 16'd6454, 16'd61027, 16'd26619, 16'd59166, 16'd25935, 16'd20359, 16'd27839, 16'd5184, 16'd9926, 16'd40104, 16'd20564, 16'd9105, 16'd20371, 16'd43658, 16'd473, 16'd20045, 16'd32551, 16'd31223, 16'd4753, 16'd46550, 16'd10681});
	test_expansion(128'hf1fa24cc196a4e3f1135d671719dd4ca, {16'd55798, 16'd28885, 16'd1973, 16'd5997, 16'd44828, 16'd41803, 16'd56273, 16'd20544, 16'd62393, 16'd45997, 16'd55394, 16'd18900, 16'd25472, 16'd27788, 16'd26132, 16'd4924, 16'd22540, 16'd51312, 16'd25922, 16'd10247, 16'd42353, 16'd16003, 16'd64477, 16'd12230, 16'd7082, 16'd20149});
	test_expansion(128'h3bc4a3b8613811cdaf57eaa22fb4434d, {16'd4010, 16'd62717, 16'd38782, 16'd53504, 16'd14452, 16'd44940, 16'd18953, 16'd3680, 16'd30674, 16'd50449, 16'd63791, 16'd39086, 16'd24662, 16'd55980, 16'd63902, 16'd8048, 16'd39363, 16'd3690, 16'd23003, 16'd39850, 16'd61684, 16'd58403, 16'd46325, 16'd56847, 16'd56738, 16'd14881});
	test_expansion(128'h705104f0efce040237fd3ad4d7ce5ab4, {16'd46061, 16'd44893, 16'd19680, 16'd4184, 16'd15296, 16'd15970, 16'd62171, 16'd44636, 16'd64765, 16'd64382, 16'd47613, 16'd37075, 16'd9681, 16'd65056, 16'd54726, 16'd20855, 16'd62330, 16'd50315, 16'd26446, 16'd3381, 16'd24661, 16'd41964, 16'd37841, 16'd64303, 16'd25619, 16'd7429});
	test_expansion(128'h062db7f14d3c00275bb32b15b877c5f3, {16'd4904, 16'd48805, 16'd60024, 16'd22358, 16'd47286, 16'd17000, 16'd53980, 16'd16249, 16'd23939, 16'd29858, 16'd45248, 16'd57195, 16'd50134, 16'd10064, 16'd56607, 16'd41830, 16'd7741, 16'd36250, 16'd51114, 16'd26658, 16'd15476, 16'd7500, 16'd35037, 16'd48366, 16'd42104, 16'd49491});
	test_expansion(128'h498a81a9b3e66928065537224d3950f0, {16'd13076, 16'd2897, 16'd22569, 16'd38803, 16'd5764, 16'd50952, 16'd22241, 16'd24973, 16'd26910, 16'd33395, 16'd20207, 16'd44070, 16'd10746, 16'd49924, 16'd58284, 16'd61526, 16'd7839, 16'd29514, 16'd47157, 16'd28120, 16'd40813, 16'd19437, 16'd21708, 16'd48624, 16'd9141, 16'd34928});
	test_expansion(128'h6e67aaaf25ff1ae57dfc02974937a8ab, {16'd48020, 16'd25222, 16'd5904, 16'd19855, 16'd36611, 16'd57091, 16'd6447, 16'd21811, 16'd61438, 16'd38684, 16'd31835, 16'd56769, 16'd57034, 16'd36568, 16'd59548, 16'd2566, 16'd18313, 16'd58321, 16'd30863, 16'd37189, 16'd19836, 16'd14271, 16'd541, 16'd20742, 16'd22439, 16'd37766});
	test_expansion(128'hdd0f6534a80013a0fb7296531aacb7d6, {16'd37185, 16'd45695, 16'd24096, 16'd21713, 16'd46736, 16'd15598, 16'd6920, 16'd16687, 16'd4726, 16'd52585, 16'd57645, 16'd40859, 16'd14644, 16'd45296, 16'd2444, 16'd39820, 16'd32069, 16'd28809, 16'd3018, 16'd12163, 16'd14477, 16'd24956, 16'd4387, 16'd50274, 16'd64787, 16'd31047});
	test_expansion(128'hc8f914d4f870d4a80db4166b42e8ca14, {16'd9400, 16'd23306, 16'd51908, 16'd35582, 16'd21419, 16'd5712, 16'd42307, 16'd23846, 16'd7471, 16'd20275, 16'd4154, 16'd10191, 16'd54284, 16'd46379, 16'd51513, 16'd3427, 16'd13055, 16'd6608, 16'd62615, 16'd13511, 16'd56730, 16'd17064, 16'd8627, 16'd62949, 16'd19089, 16'd34705});
	test_expansion(128'ha234c315198253b532077542b32d62e7, {16'd978, 16'd55702, 16'd29672, 16'd45148, 16'd4131, 16'd58455, 16'd58938, 16'd57910, 16'd26930, 16'd17459, 16'd574, 16'd28192, 16'd4029, 16'd32837, 16'd24662, 16'd3916, 16'd53304, 16'd36150, 16'd18148, 16'd44936, 16'd34711, 16'd36732, 16'd47757, 16'd33450, 16'd7598, 16'd10364});
	test_expansion(128'h16f1855b0f60c8eeab38c5b2136f56e2, {16'd43216, 16'd15298, 16'd11490, 16'd40056, 16'd21367, 16'd23855, 16'd23578, 16'd32337, 16'd34694, 16'd43117, 16'd10620, 16'd20014, 16'd57652, 16'd39876, 16'd10131, 16'd29608, 16'd33738, 16'd40470, 16'd11275, 16'd10687, 16'd16819, 16'd18658, 16'd27390, 16'd9571, 16'd37174, 16'd6836});
	test_expansion(128'hb28dfea377c3343bc574bae5720eca2f, {16'd10933, 16'd40022, 16'd54287, 16'd50359, 16'd54806, 16'd63428, 16'd48295, 16'd44225, 16'd58964, 16'd57643, 16'd61458, 16'd1727, 16'd31237, 16'd57453, 16'd53285, 16'd57790, 16'd61858, 16'd54228, 16'd63770, 16'd23521, 16'd37846, 16'd61291, 16'd51819, 16'd3094, 16'd37874, 16'd58164});
	test_expansion(128'ha13628c23cc8241ecf0940e01866428a, {16'd40849, 16'd22077, 16'd2082, 16'd6866, 16'd26861, 16'd63989, 16'd57670, 16'd5347, 16'd38141, 16'd22446, 16'd26022, 16'd28538, 16'd10063, 16'd6831, 16'd28142, 16'd63051, 16'd63217, 16'd48426, 16'd62110, 16'd15831, 16'd23502, 16'd18274, 16'd43538, 16'd31547, 16'd56198, 16'd23051});
	test_expansion(128'h12e64fa80c65b4a4e58851a1af82b204, {16'd23940, 16'd52974, 16'd59403, 16'd35376, 16'd14120, 16'd16980, 16'd4796, 16'd59426, 16'd64055, 16'd23919, 16'd40360, 16'd46527, 16'd46700, 16'd57606, 16'd43730, 16'd3790, 16'd50141, 16'd190, 16'd45382, 16'd9116, 16'd63279, 16'd34871, 16'd3151, 16'd42044, 16'd8404, 16'd14337});
	test_expansion(128'h4f6a09032fc3cb10a23608828d16eb2b, {16'd11574, 16'd64409, 16'd23749, 16'd16223, 16'd32846, 16'd4548, 16'd20330, 16'd11466, 16'd64374, 16'd60181, 16'd24485, 16'd63251, 16'd54706, 16'd7596, 16'd2045, 16'd19447, 16'd31053, 16'd23934, 16'd36471, 16'd13233, 16'd24222, 16'd33905, 16'd31106, 16'd7164, 16'd20252, 16'd23530});
	test_expansion(128'hb17acb0aabb048bcbea915bdb7bf3f27, {16'd48392, 16'd11938, 16'd18977, 16'd35379, 16'd3690, 16'd62822, 16'd662, 16'd49795, 16'd51411, 16'd402, 16'd18381, 16'd49706, 16'd57890, 16'd33777, 16'd62836, 16'd23790, 16'd53425, 16'd53703, 16'd1199, 16'd50633, 16'd7814, 16'd5249, 16'd41059, 16'd11263, 16'd1876, 16'd4803});
	test_expansion(128'hbd160ba097d3619d5e9ffcfba9e68adf, {16'd49514, 16'd45173, 16'd47609, 16'd12034, 16'd43000, 16'd39691, 16'd61548, 16'd24999, 16'd38597, 16'd46117, 16'd31894, 16'd63358, 16'd64559, 16'd14745, 16'd47547, 16'd48898, 16'd62363, 16'd38395, 16'd52323, 16'd61887, 16'd23493, 16'd46806, 16'd19331, 16'd18044, 16'd25054, 16'd39928});
	test_expansion(128'h381715975de0cd7cb9bed905964b6f5c, {16'd4940, 16'd15704, 16'd14330, 16'd32601, 16'd6824, 16'd16739, 16'd23213, 16'd36179, 16'd26388, 16'd63691, 16'd33041, 16'd660, 16'd11567, 16'd63514, 16'd24316, 16'd24246, 16'd1039, 16'd29590, 16'd17337, 16'd39766, 16'd26365, 16'd3603, 16'd9092, 16'd27315, 16'd9787, 16'd4133});
	test_expansion(128'hea756e0f689c07c30a1701e6dc3c5ba0, {16'd52760, 16'd38993, 16'd60929, 16'd27147, 16'd40116, 16'd40813, 16'd57234, 16'd4471, 16'd33957, 16'd44714, 16'd14367, 16'd49584, 16'd5054, 16'd34047, 16'd9923, 16'd45527, 16'd2614, 16'd1369, 16'd2755, 16'd58410, 16'd3965, 16'd4480, 16'd21168, 16'd38182, 16'd34083, 16'd51823});
	test_expansion(128'hacd68bfc296bcfc98fa380bb07e1788b, {16'd30223, 16'd29940, 16'd60490, 16'd19616, 16'd47868, 16'd63009, 16'd51148, 16'd32636, 16'd31572, 16'd54753, 16'd61281, 16'd50053, 16'd9269, 16'd56437, 16'd11282, 16'd61907, 16'd54763, 16'd33716, 16'd65012, 16'd17491, 16'd55916, 16'd49490, 16'd17960, 16'd47619, 16'd60121, 16'd30291});
	test_expansion(128'h927559b9d1241e3dbf932d49a69311fe, {16'd25092, 16'd2117, 16'd26082, 16'd47256, 16'd6719, 16'd34262, 16'd23909, 16'd64071, 16'd4677, 16'd4878, 16'd54504, 16'd55264, 16'd19763, 16'd32441, 16'd44992, 16'd58789, 16'd33656, 16'd34306, 16'd14291, 16'd45701, 16'd59527, 16'd35433, 16'd63972, 16'd11452, 16'd31535, 16'd7385});
	test_expansion(128'h00f4d978f31f12a9b8c9231d6f9d232f, {16'd16857, 16'd5413, 16'd50269, 16'd40872, 16'd16069, 16'd53824, 16'd15136, 16'd64786, 16'd57045, 16'd2998, 16'd30516, 16'd13109, 16'd38962, 16'd49548, 16'd14422, 16'd40409, 16'd13881, 16'd34748, 16'd24796, 16'd63806, 16'd63908, 16'd28609, 16'd40829, 16'd578, 16'd55262, 16'd50511});
	test_expansion(128'h1140b6d53d06db65d7cd95ee2506b945, {16'd55222, 16'd38640, 16'd50920, 16'd56506, 16'd37546, 16'd2063, 16'd58624, 16'd151, 16'd26337, 16'd33039, 16'd33991, 16'd33348, 16'd14398, 16'd462, 16'd23419, 16'd37339, 16'd64704, 16'd52769, 16'd8305, 16'd64710, 16'd1175, 16'd41413, 16'd1977, 16'd64576, 16'd38666, 16'd40471});
	test_expansion(128'h9739e2aaa8ef4634dd56cdc80575a3b8, {16'd13246, 16'd59851, 16'd46506, 16'd37387, 16'd22126, 16'd58991, 16'd6649, 16'd31447, 16'd12881, 16'd35979, 16'd1637, 16'd35775, 16'd13469, 16'd33989, 16'd34288, 16'd45099, 16'd61742, 16'd24653, 16'd31598, 16'd34094, 16'd19973, 16'd44417, 16'd571, 16'd25275, 16'd39702, 16'd51800});
	test_expansion(128'hb3324d8ea2ab16edc09076c97f456ef2, {16'd30183, 16'd48660, 16'd9762, 16'd64778, 16'd17787, 16'd3572, 16'd50183, 16'd4020, 16'd39171, 16'd22644, 16'd42491, 16'd62712, 16'd17896, 16'd21712, 16'd58352, 16'd12966, 16'd12199, 16'd7896, 16'd14393, 16'd29144, 16'd44837, 16'd39283, 16'd60082, 16'd57784, 16'd20299, 16'd19959});
	test_expansion(128'hce57b8adfd1beefb1cf08331e88299c3, {16'd54731, 16'd24656, 16'd4768, 16'd13807, 16'd43340, 16'd9142, 16'd41178, 16'd6972, 16'd4700, 16'd10529, 16'd1006, 16'd29431, 16'd44842, 16'd3306, 16'd25360, 16'd15442, 16'd12828, 16'd2445, 16'd37706, 16'd33187, 16'd24056, 16'd41475, 16'd3857, 16'd7992, 16'd11764, 16'd42401});
	test_expansion(128'h12c0d819657cc1c9b930d16b2508f7ad, {16'd63784, 16'd28790, 16'd27973, 16'd28836, 16'd59594, 16'd51026, 16'd13608, 16'd20885, 16'd3542, 16'd10154, 16'd2647, 16'd59487, 16'd34964, 16'd39897, 16'd11080, 16'd49953, 16'd3678, 16'd41109, 16'd17963, 16'd56361, 16'd30562, 16'd18329, 16'd24375, 16'd48438, 16'd4383, 16'd48283});
	test_expansion(128'hacfa6cbbde60f89d5deebe6ba8e49c79, {16'd24113, 16'd11046, 16'd39123, 16'd21379, 16'd2354, 16'd20877, 16'd44672, 16'd4556, 16'd22131, 16'd25077, 16'd56947, 16'd15618, 16'd57081, 16'd15128, 16'd50222, 16'd40443, 16'd6619, 16'd62784, 16'd4357, 16'd60781, 16'd32209, 16'd60825, 16'd30929, 16'd49600, 16'd23557, 16'd46407});
	test_expansion(128'h46fc6b77427afc7d8b18b33d39ce9c13, {16'd43591, 16'd31091, 16'd7147, 16'd17631, 16'd44642, 16'd50787, 16'd20230, 16'd57, 16'd54466, 16'd54993, 16'd27199, 16'd4053, 16'd4960, 16'd59407, 16'd29900, 16'd10523, 16'd17276, 16'd45028, 16'd48500, 16'd64287, 16'd38284, 16'd15154, 16'd12787, 16'd6300, 16'd42295, 16'd1277});
	test_expansion(128'hb4dae336ffaa246c2110535b0390ee13, {16'd53579, 16'd36156, 16'd50308, 16'd33457, 16'd22390, 16'd4026, 16'd1123, 16'd9692, 16'd28004, 16'd31891, 16'd5526, 16'd5585, 16'd12230, 16'd25525, 16'd56119, 16'd51106, 16'd12924, 16'd26606, 16'd42941, 16'd20403, 16'd2267, 16'd31557, 16'd6710, 16'd43648, 16'd51021, 16'd36139});
	test_expansion(128'h2780271134799283e87e714162fd92e9, {16'd44315, 16'd16644, 16'd22819, 16'd20056, 16'd17814, 16'd30658, 16'd25645, 16'd36230, 16'd30670, 16'd58936, 16'd9519, 16'd16475, 16'd11924, 16'd61489, 16'd31095, 16'd5575, 16'd32352, 16'd2471, 16'd8664, 16'd2719, 16'd53592, 16'd31309, 16'd14600, 16'd46802, 16'd18185, 16'd57821});
	test_expansion(128'hb2d8e0aad05a373a7781219ee6b8a3ab, {16'd39545, 16'd7176, 16'd63787, 16'd20220, 16'd27238, 16'd53182, 16'd3750, 16'd19545, 16'd47938, 16'd47308, 16'd37041, 16'd16409, 16'd12516, 16'd25238, 16'd9596, 16'd31592, 16'd28629, 16'd55211, 16'd57340, 16'd7245, 16'd38246, 16'd36336, 16'd23869, 16'd40380, 16'd19601, 16'd44814});
	test_expansion(128'hbeeef56f70a6c2c32b779bd5b1e1c981, {16'd39361, 16'd44380, 16'd52176, 16'd29735, 16'd36430, 16'd12335, 16'd35194, 16'd51913, 16'd42726, 16'd34148, 16'd24904, 16'd3440, 16'd20638, 16'd17261, 16'd46568, 16'd18451, 16'd59118, 16'd24741, 16'd31386, 16'd60331, 16'd1098, 16'd45431, 16'd9095, 16'd60682, 16'd56146, 16'd54426});
	test_expansion(128'h3d168a83be9cad8338f3bf833cfbaffb, {16'd56462, 16'd22874, 16'd50854, 16'd36761, 16'd32397, 16'd18940, 16'd28249, 16'd56899, 16'd62847, 16'd29640, 16'd13187, 16'd57810, 16'd62690, 16'd25173, 16'd54598, 16'd62707, 16'd14397, 16'd18822, 16'd33169, 16'd52086, 16'd65027, 16'd26382, 16'd19052, 16'd29510, 16'd16345, 16'd1149});
	test_expansion(128'h886b9b59e1b8d53203af1c3cf8c0e37b, {16'd43204, 16'd12555, 16'd61677, 16'd5068, 16'd47857, 16'd36969, 16'd20077, 16'd41020, 16'd58407, 16'd57000, 16'd9010, 16'd39011, 16'd19161, 16'd1562, 16'd36602, 16'd28120, 16'd57268, 16'd59035, 16'd55809, 16'd36662, 16'd51979, 16'd57003, 16'd14078, 16'd38586, 16'd34334, 16'd30598});
	test_expansion(128'h73a7381b585d5f4cdffb683fb95dca84, {16'd28313, 16'd38866, 16'd13665, 16'd58308, 16'd46189, 16'd62501, 16'd8465, 16'd27499, 16'd55154, 16'd30794, 16'd29720, 16'd6445, 16'd44279, 16'd26767, 16'd40753, 16'd12369, 16'd59401, 16'd54698, 16'd56364, 16'd29383, 16'd46080, 16'd4676, 16'd877, 16'd7179, 16'd55507, 16'd62154});
	test_expansion(128'hf1b3a7f810f3818a5441169fb9126d34, {16'd38499, 16'd44257, 16'd57305, 16'd2253, 16'd8298, 16'd36004, 16'd64342, 16'd27135, 16'd4031, 16'd44785, 16'd61508, 16'd51682, 16'd13586, 16'd26537, 16'd2257, 16'd12881, 16'd13551, 16'd64445, 16'd6195, 16'd28178, 16'd1205, 16'd4381, 16'd9427, 16'd40347, 16'd60169, 16'd34622});
	test_expansion(128'hac6b942c090e9a0b7ece16882a6043c8, {16'd41948, 16'd42920, 16'd16214, 16'd14465, 16'd1945, 16'd15809, 16'd19713, 16'd4491, 16'd27417, 16'd45015, 16'd192, 16'd46170, 16'd64296, 16'd36678, 16'd36104, 16'd46246, 16'd49135, 16'd48396, 16'd11216, 16'd61770, 16'd64726, 16'd27895, 16'd23580, 16'd59428, 16'd49086, 16'd29463});
	test_expansion(128'ha9ba6de5343ed64c2b1402b3e71ff4ba, {16'd53803, 16'd42079, 16'd8134, 16'd30134, 16'd59713, 16'd624, 16'd19970, 16'd36560, 16'd11940, 16'd24304, 16'd29195, 16'd7219, 16'd7315, 16'd45297, 16'd12270, 16'd14827, 16'd60397, 16'd51853, 16'd36533, 16'd26329, 16'd20326, 16'd56989, 16'd58212, 16'd65198, 16'd20417, 16'd44682});
	test_expansion(128'hc8f0d5c028ea48feaaaa2f5f0ee18813, {16'd33485, 16'd2082, 16'd24334, 16'd39617, 16'd38217, 16'd5183, 16'd39385, 16'd60767, 16'd36320, 16'd25770, 16'd16086, 16'd63740, 16'd18199, 16'd44587, 16'd34026, 16'd9284, 16'd11137, 16'd470, 16'd10141, 16'd24425, 16'd52258, 16'd38527, 16'd11877, 16'd49457, 16'd62033, 16'd56219});
	test_expansion(128'h183f5291f33e78e4cc9a22e607882d7d, {16'd12343, 16'd19578, 16'd8205, 16'd64630, 16'd59986, 16'd10312, 16'd56901, 16'd36997, 16'd13635, 16'd38090, 16'd51690, 16'd44648, 16'd11170, 16'd20831, 16'd16097, 16'd30266, 16'd26528, 16'd15682, 16'd15755, 16'd47810, 16'd46526, 16'd12068, 16'd37784, 16'd9009, 16'd9869, 16'd57566});
	test_expansion(128'h19857bb835e43709bf844709f3306b24, {16'd10032, 16'd38354, 16'd4139, 16'd48267, 16'd21809, 16'd23505, 16'd4122, 16'd47669, 16'd33356, 16'd56935, 16'd10514, 16'd5632, 16'd32045, 16'd7268, 16'd19862, 16'd44233, 16'd64814, 16'd55675, 16'd23516, 16'd9905, 16'd11356, 16'd22496, 16'd30407, 16'd9155, 16'd58666, 16'd60236});
	test_expansion(128'h898b144fae89f617293c69387135225c, {16'd45633, 16'd3657, 16'd54206, 16'd65344, 16'd32487, 16'd35830, 16'd10776, 16'd131, 16'd15366, 16'd55651, 16'd4127, 16'd64820, 16'd10527, 16'd9316, 16'd38539, 16'd28084, 16'd18142, 16'd15117, 16'd5455, 16'd53493, 16'd57967, 16'd21868, 16'd17177, 16'd30683, 16'd29782, 16'd43388});
	test_expansion(128'h0bde5f5699382b89fcc94314c6cd8b28, {16'd15443, 16'd38959, 16'd11684, 16'd25832, 16'd42076, 16'd4375, 16'd64428, 16'd31139, 16'd2992, 16'd377, 16'd1354, 16'd54449, 16'd20121, 16'd48187, 16'd51938, 16'd64235, 16'd16951, 16'd40761, 16'd27151, 16'd57017, 16'd42701, 16'd15481, 16'd61341, 16'd6138, 16'd61337, 16'd4705});
	test_expansion(128'h75b78b24c7b57b0bbabd1a363644f3bf, {16'd1491, 16'd4334, 16'd27766, 16'd28048, 16'd26585, 16'd3319, 16'd10614, 16'd35144, 16'd16553, 16'd37106, 16'd37411, 16'd3944, 16'd30853, 16'd38483, 16'd37295, 16'd21982, 16'd37455, 16'd22918, 16'd61581, 16'd31057, 16'd59730, 16'd20205, 16'd38145, 16'd4851, 16'd54357, 16'd41235});
	test_expansion(128'hfcc9ba9e1e00516ab30e61dacb084551, {16'd55357, 16'd50495, 16'd54607, 16'd33901, 16'd4914, 16'd37690, 16'd43259, 16'd3557, 16'd12133, 16'd57375, 16'd15228, 16'd43523, 16'd55677, 16'd47680, 16'd22233, 16'd32924, 16'd37699, 16'd60409, 16'd27978, 16'd34643, 16'd28484, 16'd8813, 16'd52728, 16'd20082, 16'd30444, 16'd50186});
	test_expansion(128'hee62c20968e41501c42d86aae30b3cef, {16'd54848, 16'd63475, 16'd51731, 16'd25594, 16'd22603, 16'd26170, 16'd2860, 16'd26219, 16'd52282, 16'd18666, 16'd2912, 16'd28442, 16'd60493, 16'd22938, 16'd32452, 16'd12972, 16'd62904, 16'd2434, 16'd48798, 16'd39560, 16'd61506, 16'd3641, 16'd62365, 16'd8848, 16'd53054, 16'd63278});
	test_expansion(128'h1928716f85512678e5f066edcdc5e989, {16'd4476, 16'd23027, 16'd34135, 16'd24592, 16'd35002, 16'd24815, 16'd62294, 16'd53589, 16'd4842, 16'd26742, 16'd5057, 16'd26072, 16'd26489, 16'd3306, 16'd5797, 16'd38842, 16'd20882, 16'd26754, 16'd57586, 16'd52105, 16'd13965, 16'd15209, 16'd1556, 16'd37221, 16'd15792, 16'd56939});
	test_expansion(128'hf3bd9034afa584f99f02ad1aeef195a6, {16'd47679, 16'd5946, 16'd20596, 16'd41352, 16'd50732, 16'd34884, 16'd15881, 16'd26368, 16'd35630, 16'd60399, 16'd54881, 16'd33050, 16'd35718, 16'd52184, 16'd19904, 16'd29193, 16'd29290, 16'd25687, 16'd65512, 16'd39364, 16'd23526, 16'd18312, 16'd63913, 16'd42981, 16'd58118, 16'd49014});
	test_expansion(128'h7f49a0a8a7a2dd12a1f8454ef24ba924, {16'd16974, 16'd59176, 16'd30867, 16'd5415, 16'd64446, 16'd46803, 16'd24389, 16'd52959, 16'd23659, 16'd58608, 16'd48041, 16'd12321, 16'd56750, 16'd41997, 16'd36115, 16'd506, 16'd21915, 16'd32392, 16'd51229, 16'd18302, 16'd40147, 16'd46251, 16'd43194, 16'd33615, 16'd24862, 16'd59148});
	test_expansion(128'h01937b270ef21f1cfc0ac4a13d28a62d, {16'd36445, 16'd48437, 16'd37793, 16'd29182, 16'd10780, 16'd39559, 16'd2549, 16'd47541, 16'd52680, 16'd26761, 16'd51822, 16'd5052, 16'd62412, 16'd43158, 16'd29288, 16'd62390, 16'd46458, 16'd16180, 16'd36372, 16'd12339, 16'd36466, 16'd50620, 16'd48694, 16'd63352, 16'd59892, 16'd9170});
	test_expansion(128'h5fa45097d77182a213c07eac67ce2203, {16'd7682, 16'd62937, 16'd52991, 16'd57066, 16'd4922, 16'd12552, 16'd6412, 16'd57567, 16'd51000, 16'd26422, 16'd20401, 16'd52460, 16'd25348, 16'd40153, 16'd48435, 16'd1412, 16'd40902, 16'd38775, 16'd51003, 16'd44352, 16'd52961, 16'd326, 16'd41670, 16'd61770, 16'd57717, 16'd4053});
	test_expansion(128'h3ae334046fed7ffe6b60ea877a334841, {16'd56011, 16'd22414, 16'd3493, 16'd24887, 16'd25317, 16'd13320, 16'd20252, 16'd4487, 16'd22531, 16'd18171, 16'd45660, 16'd9599, 16'd15664, 16'd34742, 16'd59340, 16'd15796, 16'd49033, 16'd40942, 16'd65055, 16'd3569, 16'd59794, 16'd20748, 16'd14404, 16'd27482, 16'd54451, 16'd2757});
	test_expansion(128'h2740c8d4e1830ea551f5632cc8e0f4d7, {16'd22207, 16'd5329, 16'd23880, 16'd28539, 16'd28109, 16'd64205, 16'd50036, 16'd32502, 16'd32061, 16'd35623, 16'd42790, 16'd52532, 16'd9715, 16'd29317, 16'd34775, 16'd4385, 16'd59554, 16'd12750, 16'd21700, 16'd29621, 16'd35970, 16'd3253, 16'd18674, 16'd23896, 16'd628, 16'd12954});
	test_expansion(128'h32a4222b9ab9296ca3789c7e72c1ae5a, {16'd62383, 16'd28663, 16'd15665, 16'd11425, 16'd12619, 16'd12014, 16'd6083, 16'd14138, 16'd51372, 16'd17164, 16'd29656, 16'd10025, 16'd53506, 16'd54367, 16'd37523, 16'd63122, 16'd1041, 16'd41750, 16'd24888, 16'd17717, 16'd22246, 16'd302, 16'd1894, 16'd30342, 16'd50832, 16'd33999});
	test_expansion(128'h2067311e85797dd7655ace679a44fbef, {16'd42115, 16'd26764, 16'd36306, 16'd27029, 16'd42322, 16'd7594, 16'd41749, 16'd37550, 16'd40071, 16'd7625, 16'd33810, 16'd13672, 16'd35350, 16'd14956, 16'd55586, 16'd3323, 16'd12217, 16'd64191, 16'd380, 16'd37106, 16'd12717, 16'd65158, 16'd43459, 16'd56596, 16'd10115, 16'd6319});
	test_expansion(128'h5360ce1a4447b852d41c65ef4925f14c, {16'd35323, 16'd33999, 16'd12807, 16'd20955, 16'd13790, 16'd63989, 16'd42985, 16'd57212, 16'd39588, 16'd63517, 16'd56183, 16'd53124, 16'd31579, 16'd37831, 16'd6226, 16'd4963, 16'd12001, 16'd29970, 16'd36649, 16'd22504, 16'd61902, 16'd24781, 16'd61359, 16'd2117, 16'd34945, 16'd10731});
	test_expansion(128'h8d4176b0401f40fbadb3318d14896966, {16'd17989, 16'd32044, 16'd43839, 16'd13484, 16'd63408, 16'd34378, 16'd57019, 16'd26550, 16'd21521, 16'd36039, 16'd35661, 16'd56509, 16'd24753, 16'd24972, 16'd62636, 16'd36126, 16'd38892, 16'd28681, 16'd11217, 16'd8030, 16'd32143, 16'd7731, 16'd5761, 16'd18404, 16'd17826, 16'd13104});
	test_expansion(128'h55352c780eb8106ea06814dabe268f35, {16'd20575, 16'd16328, 16'd45106, 16'd618, 16'd52121, 16'd50862, 16'd8998, 16'd60023, 16'd11239, 16'd27581, 16'd23514, 16'd8151, 16'd62199, 16'd20245, 16'd20180, 16'd7315, 16'd47875, 16'd38818, 16'd5794, 16'd45383, 16'd33416, 16'd21396, 16'd32535, 16'd61322, 16'd13164, 16'd37334});
	test_expansion(128'h9e49237b4d35a7d95e478ba2e62d7363, {16'd18565, 16'd7749, 16'd53197, 16'd63845, 16'd54428, 16'd2872, 16'd17057, 16'd20994, 16'd30288, 16'd7187, 16'd60281, 16'd60234, 16'd12854, 16'd62010, 16'd29841, 16'd38748, 16'd32221, 16'd16163, 16'd8591, 16'd41852, 16'd56423, 16'd55107, 16'd36127, 16'd3132, 16'd43113, 16'd60855});
	test_expansion(128'h0a1a2d9c39658a35d6fad240dae702fb, {16'd10549, 16'd13840, 16'd49448, 16'd16184, 16'd6049, 16'd38474, 16'd43306, 16'd38056, 16'd40846, 16'd57302, 16'd11544, 16'd39022, 16'd60855, 16'd42270, 16'd36866, 16'd17199, 16'd36925, 16'd50810, 16'd8269, 16'd28574, 16'd58555, 16'd25747, 16'd60139, 16'd46430, 16'd7001, 16'd11703});
	test_expansion(128'hc855d664fbbfc22c56d8d04df6cbf21b, {16'd57255, 16'd13585, 16'd57936, 16'd55129, 16'd3779, 16'd29025, 16'd17194, 16'd62624, 16'd41553, 16'd62122, 16'd47961, 16'd26770, 16'd4437, 16'd6809, 16'd44073, 16'd7305, 16'd56707, 16'd23886, 16'd30073, 16'd40336, 16'd62267, 16'd29182, 16'd9717, 16'd62512, 16'd34702, 16'd16022});
	test_expansion(128'h7c48b059236ca52b0639fc2f1cc176a3, {16'd33396, 16'd17592, 16'd65485, 16'd49879, 16'd48446, 16'd47267, 16'd38445, 16'd26330, 16'd78, 16'd14614, 16'd64016, 16'd16373, 16'd17358, 16'd13810, 16'd61008, 16'd14016, 16'd27289, 16'd7707, 16'd61043, 16'd11302, 16'd22591, 16'd32138, 16'd44992, 16'd55536, 16'd44387, 16'd12484});
	test_expansion(128'h1d412f16a2546ada8ce9211a2e57aa71, {16'd44936, 16'd65512, 16'd60588, 16'd60740, 16'd45307, 16'd45963, 16'd40841, 16'd37935, 16'd44875, 16'd2363, 16'd48434, 16'd52106, 16'd22264, 16'd59050, 16'd40040, 16'd2138, 16'd57614, 16'd13462, 16'd15070, 16'd14328, 16'd62880, 16'd40963, 16'd3647, 16'd59165, 16'd17157, 16'd28550});
	test_expansion(128'h6ec5a2d65c6d5e199b15c4b1a98cc00b, {16'd26864, 16'd42078, 16'd56583, 16'd38258, 16'd19109, 16'd44783, 16'd37237, 16'd48710, 16'd10923, 16'd64476, 16'd5991, 16'd31779, 16'd1688, 16'd63618, 16'd28890, 16'd56688, 16'd19735, 16'd55260, 16'd60234, 16'd30479, 16'd19677, 16'd28817, 16'd10559, 16'd32397, 16'd23900, 16'd9508});
	test_expansion(128'h45dad449f66c17322a37bf5e2321eaf7, {16'd22431, 16'd7092, 16'd57343, 16'd25573, 16'd59765, 16'd599, 16'd39543, 16'd9638, 16'd23033, 16'd65198, 16'd3620, 16'd27398, 16'd33767, 16'd63346, 16'd4936, 16'd24641, 16'd27575, 16'd32668, 16'd30445, 16'd26388, 16'd62632, 16'd430, 16'd55769, 16'd59906, 16'd54806, 16'd8940});
	test_expansion(128'h07a6c133b910d723466b58f8cf4dd3ac, {16'd56261, 16'd32550, 16'd2877, 16'd27595, 16'd58736, 16'd39822, 16'd48580, 16'd50428, 16'd43235, 16'd25545, 16'd1242, 16'd30298, 16'd12989, 16'd35972, 16'd1950, 16'd40276, 16'd22848, 16'd57077, 16'd6760, 16'd15788, 16'd51863, 16'd59024, 16'd48973, 16'd4077, 16'd40748, 16'd35104});
	test_expansion(128'h60d8fe6623f9b15c4205b164478f5739, {16'd19890, 16'd9368, 16'd65000, 16'd39128, 16'd18876, 16'd21295, 16'd55972, 16'd16905, 16'd47953, 16'd19226, 16'd48993, 16'd58994, 16'd62177, 16'd33808, 16'd27214, 16'd61400, 16'd63157, 16'd20527, 16'd6841, 16'd61364, 16'd50480, 16'd19628, 16'd34216, 16'd22067, 16'd19907, 16'd51767});
	test_expansion(128'hf2a7d83f7201005a62d38189df1da460, {16'd50049, 16'd64655, 16'd59411, 16'd20080, 16'd29944, 16'd37446, 16'd31416, 16'd17377, 16'd41042, 16'd55251, 16'd29647, 16'd13188, 16'd20738, 16'd46774, 16'd47193, 16'd54350, 16'd1482, 16'd48115, 16'd11407, 16'd6265, 16'd42645, 16'd23756, 16'd27305, 16'd29228, 16'd64926, 16'd50237});
	test_expansion(128'h9052ac2d6a1555372472e928a2eb702c, {16'd31914, 16'd10297, 16'd15460, 16'd2610, 16'd63687, 16'd37717, 16'd24120, 16'd13843, 16'd38186, 16'd58764, 16'd59882, 16'd14137, 16'd61893, 16'd7277, 16'd1917, 16'd7874, 16'd29091, 16'd15928, 16'd5233, 16'd64012, 16'd33712, 16'd29206, 16'd58073, 16'd53363, 16'd31571, 16'd13085});
	test_expansion(128'h231e5f103250ce0359bb22cec73ab6fe, {16'd61527, 16'd20338, 16'd55834, 16'd55977, 16'd5186, 16'd50037, 16'd42411, 16'd51493, 16'd50137, 16'd34800, 16'd58726, 16'd34740, 16'd52255, 16'd19256, 16'd62490, 16'd60450, 16'd57954, 16'd15353, 16'd5632, 16'd13163, 16'd25906, 16'd40904, 16'd37389, 16'd27412, 16'd54746, 16'd47211});
	test_expansion(128'hc0f3f0adbd566ff7d336da8e86fe005d, {16'd38423, 16'd4381, 16'd21398, 16'd2609, 16'd63502, 16'd43090, 16'd3974, 16'd26769, 16'd63717, 16'd23460, 16'd55287, 16'd47338, 16'd39416, 16'd60854, 16'd1352, 16'd4221, 16'd54379, 16'd8862, 16'd14388, 16'd5264, 16'd10935, 16'd57388, 16'd2048, 16'd41494, 16'd26034, 16'd8322});
	test_expansion(128'hc6d654c18350af67275d371592232aa0, {16'd55708, 16'd11926, 16'd46483, 16'd50212, 16'd33292, 16'd30591, 16'd25386, 16'd18493, 16'd3746, 16'd33740, 16'd8970, 16'd64017, 16'd45548, 16'd48786, 16'd32827, 16'd29589, 16'd49276, 16'd60875, 16'd28171, 16'd10543, 16'd42362, 16'd20208, 16'd8590, 16'd25388, 16'd11077, 16'd52907});
	test_expansion(128'h9a0ef4eedacbcf9b89da493786cee45b, {16'd18299, 16'd23669, 16'd6450, 16'd55291, 16'd34257, 16'd30489, 16'd41450, 16'd51537, 16'd28737, 16'd27672, 16'd44224, 16'd20534, 16'd64891, 16'd32017, 16'd21898, 16'd26224, 16'd27499, 16'd3638, 16'd29533, 16'd13409, 16'd1101, 16'd32250, 16'd4587, 16'd36330, 16'd51599, 16'd31931});
	test_expansion(128'hf7c333b35d34ad6ba6e7076d86b61d4d, {16'd61079, 16'd48152, 16'd20510, 16'd30023, 16'd59519, 16'd16767, 16'd63468, 16'd35314, 16'd24383, 16'd12845, 16'd30174, 16'd20254, 16'd19175, 16'd28825, 16'd12892, 16'd58770, 16'd5480, 16'd42648, 16'd58493, 16'd36119, 16'd4448, 16'd56607, 16'd20624, 16'd10219, 16'd40465, 16'd45928});
	test_expansion(128'h9ce53c3394745f8c20c20b2e767c04a0, {16'd18949, 16'd12158, 16'd25471, 16'd22527, 16'd21492, 16'd42520, 16'd28893, 16'd11737, 16'd23724, 16'd52540, 16'd48558, 16'd53258, 16'd59764, 16'd27536, 16'd16510, 16'd64554, 16'd9395, 16'd52177, 16'd16314, 16'd46229, 16'd48304, 16'd2018, 16'd44101, 16'd13661, 16'd1635, 16'd60317});
	test_expansion(128'hf669b332e67adb07fcbacceae8acdf9b, {16'd15206, 16'd16341, 16'd57668, 16'd28008, 16'd44110, 16'd19574, 16'd34063, 16'd46480, 16'd18803, 16'd33820, 16'd22844, 16'd9565, 16'd31674, 16'd11934, 16'd3203, 16'd11687, 16'd64007, 16'd22488, 16'd45979, 16'd53908, 16'd130, 16'd64483, 16'd18928, 16'd37217, 16'd18641, 16'd21270});
	test_expansion(128'h0d985cb077126ca9222d9c9c5ad71adc, {16'd33456, 16'd63618, 16'd61139, 16'd21466, 16'd40062, 16'd22688, 16'd58715, 16'd63284, 16'd27498, 16'd9144, 16'd18117, 16'd53798, 16'd1971, 16'd52335, 16'd2449, 16'd8113, 16'd35105, 16'd38116, 16'd55172, 16'd18393, 16'd53789, 16'd58950, 16'd18785, 16'd57375, 16'd17611, 16'd10153});
	test_expansion(128'h2c2ff8267dadd8a0f7581b000a500468, {16'd18689, 16'd22717, 16'd37611, 16'd3823, 16'd30896, 16'd64543, 16'd11105, 16'd40892, 16'd65080, 16'd8097, 16'd41633, 16'd8684, 16'd29750, 16'd38361, 16'd2550, 16'd7448, 16'd21555, 16'd54491, 16'd39587, 16'd24919, 16'd24213, 16'd41603, 16'd9440, 16'd16699, 16'd33050, 16'd2066});
	test_expansion(128'h3cad57f5f0f59ff054710912fedf9f50, {16'd21880, 16'd522, 16'd41343, 16'd31375, 16'd52222, 16'd39203, 16'd43913, 16'd41342, 16'd51589, 16'd29315, 16'd44133, 16'd13595, 16'd31885, 16'd63057, 16'd43026, 16'd26329, 16'd9225, 16'd60870, 16'd53086, 16'd4033, 16'd27009, 16'd25391, 16'd21033, 16'd38384, 16'd22357, 16'd60494});
	test_expansion(128'h435d6083a1c4fff1539f7d1f09757ae5, {16'd34064, 16'd37620, 16'd24188, 16'd47688, 16'd42151, 16'd990, 16'd41567, 16'd28997, 16'd16147, 16'd32096, 16'd2568, 16'd24596, 16'd11341, 16'd12355, 16'd55479, 16'd39164, 16'd44678, 16'd1861, 16'd8877, 16'd660, 16'd51827, 16'd64997, 16'd56377, 16'd41080, 16'd62195, 16'd62766});
	test_expansion(128'h22180c51340056013bbbb5e695a20f91, {16'd58550, 16'd15435, 16'd26673, 16'd29313, 16'd32611, 16'd36467, 16'd57500, 16'd19037, 16'd4152, 16'd37082, 16'd20084, 16'd14213, 16'd53503, 16'd63463, 16'd14341, 16'd25765, 16'd49995, 16'd30220, 16'd3552, 16'd23955, 16'd41188, 16'd61118, 16'd21531, 16'd53807, 16'd48865, 16'd26896});
	test_expansion(128'h25bec1b3d5442df7d6fa249d92a1aee5, {16'd32224, 16'd56317, 16'd31080, 16'd26887, 16'd44486, 16'd29809, 16'd14407, 16'd34137, 16'd56104, 16'd63266, 16'd1739, 16'd14143, 16'd25229, 16'd22985, 16'd31860, 16'd28722, 16'd6407, 16'd54883, 16'd39668, 16'd21256, 16'd41261, 16'd20296, 16'd6446, 16'd19521, 16'd34473, 16'd64980});
	test_expansion(128'h8893a754817b18cd81a670eccef7e1a7, {16'd58580, 16'd17706, 16'd31567, 16'd30669, 16'd47908, 16'd10471, 16'd50919, 16'd17211, 16'd18485, 16'd41257, 16'd27630, 16'd49261, 16'd10489, 16'd11005, 16'd33762, 16'd29527, 16'd8045, 16'd26949, 16'd3895, 16'd13904, 16'd6746, 16'd7172, 16'd48353, 16'd32507, 16'd33214, 16'd15980});
	test_expansion(128'hf86310edaea7fefe146d509768dbafb6, {16'd4063, 16'd49606, 16'd8180, 16'd58071, 16'd1732, 16'd37406, 16'd40535, 16'd250, 16'd58728, 16'd40970, 16'd9920, 16'd22435, 16'd55798, 16'd978, 16'd4384, 16'd12115, 16'd61968, 16'd52587, 16'd25864, 16'd13511, 16'd32013, 16'd52399, 16'd55904, 16'd34827, 16'd61485, 16'd5366});
	test_expansion(128'h0bad0f0967cd05ba6338927c23bea1b4, {16'd4354, 16'd18959, 16'd50981, 16'd46637, 16'd1189, 16'd28403, 16'd52587, 16'd16833, 16'd62768, 16'd38507, 16'd16333, 16'd9711, 16'd27093, 16'd58619, 16'd30146, 16'd47587, 16'd32118, 16'd48258, 16'd10606, 16'd13035, 16'd13676, 16'd12531, 16'd26977, 16'd11316, 16'd50065, 16'd13215});
	test_expansion(128'hf4daeccd1c182799b970443ab79e90c6, {16'd19539, 16'd13679, 16'd4737, 16'd9484, 16'd45075, 16'd2151, 16'd27221, 16'd48597, 16'd23417, 16'd63771, 16'd20230, 16'd26848, 16'd59797, 16'd33677, 16'd41471, 16'd35501, 16'd38273, 16'd12422, 16'd22909, 16'd28299, 16'd9821, 16'd51357, 16'd38302, 16'd60024, 16'd53522, 16'd11293});
	test_expansion(128'hc2f04d1898341e4f01582a9f65e25887, {16'd64480, 16'd55817, 16'd53081, 16'd31336, 16'd14746, 16'd63347, 16'd59451, 16'd5274, 16'd5805, 16'd20768, 16'd64650, 16'd34576, 16'd39119, 16'd1569, 16'd23176, 16'd58757, 16'd35228, 16'd52996, 16'd26260, 16'd14331, 16'd46778, 16'd31573, 16'd55430, 16'd31580, 16'd19937, 16'd34329});
	test_expansion(128'hd5348735322c359fca3aabdab8cc8a77, {16'd61330, 16'd8486, 16'd6703, 16'd58382, 16'd498, 16'd57899, 16'd4193, 16'd58357, 16'd1144, 16'd20122, 16'd50933, 16'd25329, 16'd28095, 16'd45793, 16'd27581, 16'd29077, 16'd39929, 16'd35344, 16'd30719, 16'd46695, 16'd3854, 16'd27221, 16'd43249, 16'd48937, 16'd9713, 16'd35253});
	test_expansion(128'h9b6ca85462b1b3f40163cd86882eb95f, {16'd45715, 16'd37450, 16'd19903, 16'd60915, 16'd60521, 16'd209, 16'd34813, 16'd6910, 16'd54057, 16'd56200, 16'd56409, 16'd62753, 16'd58447, 16'd5657, 16'd30106, 16'd58177, 16'd41239, 16'd25891, 16'd9910, 16'd46101, 16'd46004, 16'd44989, 16'd49945, 16'd4854, 16'd52237, 16'd38090});
	test_expansion(128'hee77845d85576e8cfea559140789fb84, {16'd23495, 16'd30526, 16'd27435, 16'd59297, 16'd59377, 16'd31811, 16'd6696, 16'd46794, 16'd30170, 16'd65500, 16'd41785, 16'd45408, 16'd4506, 16'd59133, 16'd6733, 16'd62403, 16'd56985, 16'd30209, 16'd65503, 16'd11682, 16'd46772, 16'd6048, 16'd25973, 16'd1416, 16'd6619, 16'd30770});
	test_expansion(128'h2fd1b759cdab9c91b0247e231ca4caed, {16'd1433, 16'd18937, 16'd46495, 16'd5708, 16'd2908, 16'd63790, 16'd61073, 16'd15205, 16'd6909, 16'd2909, 16'd39702, 16'd9825, 16'd12883, 16'd35474, 16'd52288, 16'd7840, 16'd22400, 16'd43999, 16'd59653, 16'd6952, 16'd62418, 16'd64259, 16'd21404, 16'd36848, 16'd12213, 16'd26102});
	test_expansion(128'hf30d63c6b292995ac46fb87d9fec0a0f, {16'd13618, 16'd54322, 16'd10361, 16'd48687, 16'd12293, 16'd51695, 16'd4053, 16'd60454, 16'd22987, 16'd40029, 16'd35382, 16'd22395, 16'd19080, 16'd57246, 16'd41425, 16'd22101, 16'd26842, 16'd36786, 16'd31774, 16'd11121, 16'd23450, 16'd64022, 16'd43610, 16'd15180, 16'd33779, 16'd49442});
	test_expansion(128'h967c2cd1b44322a60ad9341a9fd7628a, {16'd22572, 16'd44251, 16'd38077, 16'd17158, 16'd18532, 16'd61287, 16'd45607, 16'd60695, 16'd1208, 16'd7150, 16'd9882, 16'd57096, 16'd39619, 16'd3223, 16'd58663, 16'd17301, 16'd59767, 16'd59391, 16'd15585, 16'd52614, 16'd13664, 16'd44705, 16'd30239, 16'd58850, 16'd40260, 16'd2845});
	test_expansion(128'hcdbd588285fc7630b8c67905fce5b81a, {16'd42771, 16'd58224, 16'd63178, 16'd42764, 16'd13942, 16'd21957, 16'd7910, 16'd55203, 16'd47329, 16'd41548, 16'd54887, 16'd24602, 16'd56462, 16'd52453, 16'd24374, 16'd53991, 16'd46191, 16'd61188, 16'd62004, 16'd49042, 16'd493, 16'd28734, 16'd62473, 16'd35911, 16'd56913, 16'd8508});
	test_expansion(128'h6ff7f6239c132e4faa4f99e1d26821de, {16'd57601, 16'd44197, 16'd42677, 16'd18332, 16'd59754, 16'd11239, 16'd59926, 16'd45064, 16'd56489, 16'd52226, 16'd40867, 16'd27616, 16'd34564, 16'd6336, 16'd44396, 16'd31368, 16'd52914, 16'd52336, 16'd41801, 16'd58405, 16'd45390, 16'd26283, 16'd59328, 16'd6641, 16'd55484, 16'd34922});
	test_expansion(128'h0354262af556fb5241f91a8c9af9d897, {16'd45210, 16'd23153, 16'd50108, 16'd60345, 16'd59839, 16'd50215, 16'd643, 16'd51540, 16'd33401, 16'd48325, 16'd21775, 16'd20164, 16'd58118, 16'd34756, 16'd27670, 16'd17716, 16'd47118, 16'd17309, 16'd19066, 16'd51249, 16'd41333, 16'd57899, 16'd40534, 16'd22595, 16'd45829, 16'd45050});
	test_expansion(128'ha6116a111e1a9c34b71957fcb226a420, {16'd19195, 16'd9959, 16'd21155, 16'd22036, 16'd53532, 16'd58252, 16'd29937, 16'd30673, 16'd50059, 16'd48219, 16'd26011, 16'd679, 16'd47895, 16'd56851, 16'd57390, 16'd26251, 16'd48948, 16'd41511, 16'd48524, 16'd45701, 16'd57391, 16'd4778, 16'd24193, 16'd53245, 16'd38454, 16'd1173});
	test_expansion(128'hc0210152d896232515bd72e1e6d9e94b, {16'd47624, 16'd59412, 16'd53938, 16'd44577, 16'd49641, 16'd35998, 16'd60169, 16'd61268, 16'd56381, 16'd8987, 16'd44196, 16'd29886, 16'd50514, 16'd3043, 16'd43146, 16'd57948, 16'd39226, 16'd62374, 16'd53430, 16'd43061, 16'd19207, 16'd39228, 16'd14628, 16'd49478, 16'd397, 16'd45955});
	test_expansion(128'h5f2b42a4bf1f4b053b1c14ea8e771b38, {16'd26952, 16'd22124, 16'd33758, 16'd38742, 16'd56340, 16'd20913, 16'd24069, 16'd39996, 16'd29649, 16'd51937, 16'd39253, 16'd60422, 16'd48655, 16'd38326, 16'd58992, 16'd13519, 16'd10554, 16'd24543, 16'd61120, 16'd57428, 16'd12271, 16'd61755, 16'd30706, 16'd3864, 16'd23408, 16'd24810});
	test_expansion(128'hafae244ddec5e3f47b3b411ac8fc12d8, {16'd47098, 16'd56652, 16'd35088, 16'd1501, 16'd37012, 16'd20961, 16'd15915, 16'd48906, 16'd14768, 16'd9841, 16'd26689, 16'd44551, 16'd9956, 16'd36240, 16'd35135, 16'd14012, 16'd2098, 16'd49621, 16'd58562, 16'd7844, 16'd40804, 16'd7415, 16'd5765, 16'd28418, 16'd62937, 16'd17164});
	test_expansion(128'hb872682c61c9dc04f356a2407ada1c20, {16'd19172, 16'd47100, 16'd31344, 16'd38335, 16'd43682, 16'd60640, 16'd30990, 16'd14799, 16'd805, 16'd24492, 16'd14928, 16'd6212, 16'd9733, 16'd1970, 16'd35576, 16'd17451, 16'd14776, 16'd53105, 16'd13391, 16'd26213, 16'd23140, 16'd25442, 16'd44277, 16'd8833, 16'd62909, 16'd30234});
	test_expansion(128'h5845c26a0a8de34ae45e04e80fd0ce3d, {16'd3164, 16'd22329, 16'd112, 16'd47439, 16'd42769, 16'd23615, 16'd48371, 16'd53612, 16'd57784, 16'd63192, 16'd13499, 16'd20634, 16'd60715, 16'd17716, 16'd58804, 16'd31689, 16'd55149, 16'd59572, 16'd19783, 16'd1371, 16'd15670, 16'd27446, 16'd478, 16'd53233, 16'd53132, 16'd26145});
	test_expansion(128'h3dd79a9f8979199a54bcf282405626b4, {16'd23189, 16'd47496, 16'd52466, 16'd58533, 16'd4836, 16'd36051, 16'd22438, 16'd48121, 16'd33334, 16'd49148, 16'd28130, 16'd4702, 16'd49245, 16'd29582, 16'd54524, 16'd2733, 16'd10550, 16'd35767, 16'd25222, 16'd40524, 16'd19789, 16'd44114, 16'd44099, 16'd62241, 16'd61948, 16'd11796});
	test_expansion(128'h089c999481b13484aadadf3d290f77c3, {16'd40534, 16'd42928, 16'd58241, 16'd25827, 16'd46608, 16'd51941, 16'd19201, 16'd47929, 16'd19144, 16'd35038, 16'd20485, 16'd12969, 16'd18033, 16'd30169, 16'd31236, 16'd33182, 16'd55902, 16'd47812, 16'd30043, 16'd21210, 16'd51935, 16'd30001, 16'd35432, 16'd11922, 16'd16332, 16'd57445});
	test_expansion(128'had6762caedc4bc95cfc9f9eb7dfaa41c, {16'd48707, 16'd33989, 16'd12802, 16'd4683, 16'd4238, 16'd12934, 16'd13259, 16'd38733, 16'd12968, 16'd35338, 16'd23463, 16'd31816, 16'd38579, 16'd55571, 16'd55789, 16'd63117, 16'd50578, 16'd11537, 16'd9825, 16'd27919, 16'd2318, 16'd1658, 16'd2474, 16'd50254, 16'd28607, 16'd42362});
	test_expansion(128'hc4be1e9d78ccbad8311d3b08f059fc96, {16'd61273, 16'd28328, 16'd23235, 16'd3077, 16'd42281, 16'd34984, 16'd49503, 16'd40757, 16'd60827, 16'd33437, 16'd9418, 16'd46547, 16'd44547, 16'd41505, 16'd45001, 16'd46321, 16'd48803, 16'd49833, 16'd40455, 16'd29620, 16'd43647, 16'd48925, 16'd51656, 16'd53371, 16'd5367, 16'd10597});
	test_expansion(128'h008b157b16e71a7e0dc8f36a18464f90, {16'd34273, 16'd32842, 16'd46458, 16'd21837, 16'd38149, 16'd54430, 16'd55434, 16'd41143, 16'd28414, 16'd32408, 16'd7169, 16'd10462, 16'd18185, 16'd11182, 16'd6816, 16'd48277, 16'd47368, 16'd42137, 16'd59344, 16'd36594, 16'd45989, 16'd27248, 16'd37944, 16'd42018, 16'd54409, 16'd46428});
	test_expansion(128'hf0574c3a3d4e53595446950488f186cc, {16'd65027, 16'd22147, 16'd22585, 16'd32577, 16'd17969, 16'd64850, 16'd47365, 16'd64098, 16'd39402, 16'd41993, 16'd17587, 16'd17096, 16'd19209, 16'd3818, 16'd64456, 16'd56480, 16'd34551, 16'd41421, 16'd11121, 16'd23430, 16'd17524, 16'd57285, 16'd53872, 16'd3445, 16'd22717, 16'd53924});
	test_expansion(128'ha1a9176ce634e98ff4b15244ec6ee791, {16'd43264, 16'd49377, 16'd9717, 16'd48950, 16'd25447, 16'd28358, 16'd40077, 16'd4219, 16'd44327, 16'd62871, 16'd15031, 16'd12606, 16'd29674, 16'd3008, 16'd28427, 16'd58081, 16'd34347, 16'd45682, 16'd13996, 16'd51080, 16'd38672, 16'd15175, 16'd51068, 16'd30254, 16'd40218, 16'd29655});
	test_expansion(128'h44025ff9d03ce1529099acbb7d5fd030, {16'd24911, 16'd12739, 16'd56567, 16'd32379, 16'd34075, 16'd40847, 16'd52306, 16'd19351, 16'd54550, 16'd15711, 16'd15304, 16'd47943, 16'd19569, 16'd44148, 16'd14324, 16'd29210, 16'd26570, 16'd18887, 16'd12746, 16'd315, 16'd7339, 16'd6360, 16'd12184, 16'd31282, 16'd37298, 16'd2459});
	test_expansion(128'hc25dc436de40e68d942fabd1a4a3e285, {16'd30057, 16'd34558, 16'd7853, 16'd53044, 16'd55922, 16'd17869, 16'd25246, 16'd25708, 16'd31450, 16'd30108, 16'd40056, 16'd43244, 16'd57597, 16'd51414, 16'd12716, 16'd47052, 16'd18639, 16'd64168, 16'd36780, 16'd56634, 16'd61515, 16'd26627, 16'd31194, 16'd6401, 16'd49881, 16'd18764});
	test_expansion(128'h31d65fdd2f5b902500ba6d2ef9a47309, {16'd13316, 16'd42046, 16'd15956, 16'd57260, 16'd25200, 16'd58239, 16'd4874, 16'd33212, 16'd33739, 16'd19705, 16'd4482, 16'd59701, 16'd58424, 16'd4082, 16'd32859, 16'd20475, 16'd12210, 16'd38267, 16'd47043, 16'd34317, 16'd64333, 16'd12924, 16'd59146, 16'd58746, 16'd41998, 16'd33582});
	test_expansion(128'hd3b97958956f63b2d54a6cffcb9261f8, {16'd17301, 16'd64996, 16'd14826, 16'd9481, 16'd38371, 16'd24984, 16'd54718, 16'd28629, 16'd27929, 16'd60594, 16'd17362, 16'd373, 16'd57876, 16'd12946, 16'd18422, 16'd42904, 16'd47866, 16'd34753, 16'd64776, 16'd14122, 16'd10240, 16'd9040, 16'd29491, 16'd2529, 16'd38323, 16'd58860});
	test_expansion(128'h9d1182e326eb1533db8671570ce31fc7, {16'd16062, 16'd21815, 16'd1965, 16'd34837, 16'd25438, 16'd23964, 16'd1370, 16'd14799, 16'd15517, 16'd40482, 16'd20842, 16'd1225, 16'd3394, 16'd37905, 16'd62030, 16'd9049, 16'd39284, 16'd17480, 16'd109, 16'd6005, 16'd63057, 16'd32911, 16'd19161, 16'd53044, 16'd34104, 16'd17543});
	test_expansion(128'h5b664d55b1c36921627ac10ae33db5b1, {16'd9164, 16'd33881, 16'd33838, 16'd1899, 16'd6047, 16'd38614, 16'd8474, 16'd43429, 16'd64825, 16'd29149, 16'd53494, 16'd60457, 16'd57220, 16'd44201, 16'd17541, 16'd52188, 16'd24140, 16'd30943, 16'd48460, 16'd40098, 16'd49985, 16'd32004, 16'd41348, 16'd59920, 16'd46933, 16'd40736});
	test_expansion(128'h60f61eca5d03ef604fe89abf381fd953, {16'd12015, 16'd50799, 16'd32451, 16'd54942, 16'd64056, 16'd1910, 16'd36874, 16'd49109, 16'd8837, 16'd58231, 16'd52994, 16'd15868, 16'd51964, 16'd56118, 16'd62549, 16'd52880, 16'd40584, 16'd2467, 16'd16059, 16'd37519, 16'd64463, 16'd11887, 16'd11897, 16'd16026, 16'd22327, 16'd34953});
	test_expansion(128'h0a2ac0f9d23dbcc3ec3082d99d8c258f, {16'd5198, 16'd40099, 16'd32613, 16'd803, 16'd30575, 16'd57393, 16'd52407, 16'd34096, 16'd10983, 16'd15466, 16'd35219, 16'd49281, 16'd58038, 16'd48604, 16'd2500, 16'd64885, 16'd43260, 16'd32700, 16'd6751, 16'd17250, 16'd61658, 16'd25519, 16'd5492, 16'd41268, 16'd38902, 16'd58044});
	test_expansion(128'hf7170f5d6c108d1ac4847d9d021d79bd, {16'd29116, 16'd49668, 16'd55498, 16'd40323, 16'd4220, 16'd498, 16'd28772, 16'd2886, 16'd20958, 16'd50897, 16'd12880, 16'd37049, 16'd55587, 16'd55839, 16'd31093, 16'd63611, 16'd46276, 16'd26553, 16'd39008, 16'd31087, 16'd36607, 16'd50654, 16'd59012, 16'd51912, 16'd19384, 16'd64480});
	test_expansion(128'h0415b05ea5168bf570326671518ecc88, {16'd19405, 16'd11475, 16'd52377, 16'd56798, 16'd61839, 16'd16327, 16'd46351, 16'd20824, 16'd3796, 16'd46280, 16'd14593, 16'd3129, 16'd56260, 16'd50405, 16'd10521, 16'd26079, 16'd24590, 16'd47379, 16'd43684, 16'd56566, 16'd45720, 16'd5052, 16'd60053, 16'd30958, 16'd23335, 16'd22396});
	test_expansion(128'h3e20f23a1b41144c0ec1d90abb4e30be, {16'd21690, 16'd44302, 16'd16824, 16'd34020, 16'd28877, 16'd64953, 16'd1038, 16'd23506, 16'd64390, 16'd42077, 16'd42612, 16'd17217, 16'd51361, 16'd13794, 16'd57946, 16'd65400, 16'd8680, 16'd43019, 16'd61325, 16'd32728, 16'd16874, 16'd13023, 16'd51030, 16'd45040, 16'd2102, 16'd24139});
	test_expansion(128'hf34b0c9a923de67237337f8497b2fb6a, {16'd17622, 16'd26408, 16'd36233, 16'd7931, 16'd25542, 16'd41677, 16'd49741, 16'd43939, 16'd6917, 16'd2393, 16'd3284, 16'd65380, 16'd50598, 16'd62120, 16'd55876, 16'd3118, 16'd50059, 16'd14599, 16'd54714, 16'd51745, 16'd24845, 16'd58676, 16'd40198, 16'd25203, 16'd20158, 16'd63155});
	test_expansion(128'h7f900c4c3f36c11652f8b30e91278fda, {16'd39694, 16'd52192, 16'd33508, 16'd24041, 16'd15478, 16'd59744, 16'd18126, 16'd48534, 16'd52978, 16'd45887, 16'd49892, 16'd50510, 16'd62133, 16'd40334, 16'd21234, 16'd52372, 16'd39274, 16'd16948, 16'd35211, 16'd60613, 16'd11796, 16'd15401, 16'd25651, 16'd58771, 16'd29711, 16'd55467});
	test_expansion(128'h9f97331b4d8def3b85bf037f969537bf, {16'd43948, 16'd20176, 16'd60119, 16'd49726, 16'd10311, 16'd21054, 16'd40550, 16'd53442, 16'd27619, 16'd34629, 16'd10378, 16'd32872, 16'd28027, 16'd48257, 16'd15383, 16'd34616, 16'd3104, 16'd48486, 16'd10892, 16'd9966, 16'd50784, 16'd36946, 16'd3923, 16'd36900, 16'd34558, 16'd23083});
	test_expansion(128'hd6f82d08f715e6143bd7fc00d9fef3b8, {16'd52761, 16'd7763, 16'd62709, 16'd45805, 16'd55218, 16'd33776, 16'd43764, 16'd17130, 16'd21812, 16'd41686, 16'd38568, 16'd29481, 16'd41962, 16'd36079, 16'd37898, 16'd31096, 16'd38731, 16'd60819, 16'd6121, 16'd42839, 16'd24524, 16'd9285, 16'd22986, 16'd64801, 16'd41730, 16'd20566});
	test_expansion(128'h791e1a82f22180dfec73f0f6fceb472e, {16'd44367, 16'd41414, 16'd28008, 16'd37454, 16'd36655, 16'd33968, 16'd6088, 16'd42366, 16'd42419, 16'd64306, 16'd54243, 16'd8140, 16'd54707, 16'd46349, 16'd23551, 16'd35507, 16'd21111, 16'd58080, 16'd18153, 16'd42735, 16'd1889, 16'd31086, 16'd49352, 16'd10423, 16'd54468, 16'd49996});
	test_expansion(128'h5207ed76cc63af2f49bc7c5b7ed5acbf, {16'd55756, 16'd29910, 16'd28354, 16'd54934, 16'd20416, 16'd61531, 16'd55709, 16'd31319, 16'd18944, 16'd50395, 16'd59453, 16'd36264, 16'd27363, 16'd24837, 16'd61748, 16'd64926, 16'd7323, 16'd59783, 16'd33561, 16'd56820, 16'd4164, 16'd30021, 16'd9373, 16'd6675, 16'd25683, 16'd24423});
	test_expansion(128'hb56ee6368b690d91ddcb9825e3dbec78, {16'd51617, 16'd9242, 16'd26951, 16'd45724, 16'd37659, 16'd46445, 16'd9219, 16'd43527, 16'd22552, 16'd30199, 16'd9834, 16'd24109, 16'd13299, 16'd42870, 16'd55901, 16'd17858, 16'd31847, 16'd39092, 16'd30032, 16'd18519, 16'd3771, 16'd32669, 16'd6149, 16'd2209, 16'd63567, 16'd64769});
	test_expansion(128'h8d08d4905ecdb9e39e5213dff51a67d8, {16'd32774, 16'd6092, 16'd20110, 16'd21656, 16'd55902, 16'd27408, 16'd64438, 16'd48754, 16'd37211, 16'd40468, 16'd8038, 16'd7951, 16'd49205, 16'd5954, 16'd31251, 16'd5087, 16'd28966, 16'd6841, 16'd45322, 16'd31773, 16'd16560, 16'd49467, 16'd48606, 16'd9131, 16'd44255, 16'd41667});
	test_expansion(128'h1882ebd16b663fd40b8829c13b0c3f94, {16'd58218, 16'd30252, 16'd45251, 16'd54515, 16'd35154, 16'd14512, 16'd23875, 16'd37496, 16'd5053, 16'd12695, 16'd46052, 16'd33669, 16'd950, 16'd30174, 16'd20229, 16'd25192, 16'd34757, 16'd10368, 16'd30726, 16'd2234, 16'd11039, 16'd17128, 16'd4707, 16'd55555, 16'd64324, 16'd22832});
	test_expansion(128'h9e5424249560129856f3e6b3c7cd264a, {16'd54131, 16'd12779, 16'd41018, 16'd46419, 16'd32931, 16'd12215, 16'd26992, 16'd30496, 16'd46778, 16'd18150, 16'd3853, 16'd32535, 16'd36724, 16'd40479, 16'd16317, 16'd45555, 16'd31586, 16'd46367, 16'd15166, 16'd26325, 16'd59924, 16'd34471, 16'd36170, 16'd34384, 16'd1511, 16'd40352});
	test_expansion(128'h7adce0de3ddec5334504ef0a2db2f4b3, {16'd47989, 16'd58331, 16'd9584, 16'd48514, 16'd6973, 16'd21477, 16'd19719, 16'd378, 16'd2065, 16'd58995, 16'd6364, 16'd19795, 16'd59686, 16'd38931, 16'd15189, 16'd15455, 16'd2134, 16'd15496, 16'd29559, 16'd50664, 16'd43446, 16'd19771, 16'd10995, 16'd33434, 16'd24813, 16'd14818});
	test_expansion(128'h2d56dee9b0f09833dba8da9001037f34, {16'd43518, 16'd25506, 16'd27976, 16'd18716, 16'd39847, 16'd3701, 16'd3103, 16'd36241, 16'd33101, 16'd10270, 16'd10303, 16'd18077, 16'd35855, 16'd39506, 16'd17889, 16'd27344, 16'd51574, 16'd5780, 16'd65164, 16'd3701, 16'd37581, 16'd26439, 16'd43726, 16'd9479, 16'd16020, 16'd46733});
	test_expansion(128'h9bee535f9bf675d40aff1424807e40a8, {16'd44802, 16'd20852, 16'd48687, 16'd30498, 16'd9825, 16'd9724, 16'd20901, 16'd34329, 16'd60311, 16'd48855, 16'd12279, 16'd34895, 16'd427, 16'd35504, 16'd8614, 16'd31502, 16'd63804, 16'd42793, 16'd12753, 16'd5518, 16'd38002, 16'd45063, 16'd65163, 16'd24201, 16'd34222, 16'd19849});
	test_expansion(128'ha4d2add2e32197304f410637375594f1, {16'd815, 16'd17838, 16'd19722, 16'd52623, 16'd56502, 16'd29254, 16'd51420, 16'd14441, 16'd61539, 16'd8248, 16'd48754, 16'd11925, 16'd7857, 16'd38442, 16'd26457, 16'd56142, 16'd57930, 16'd5531, 16'd61583, 16'd55435, 16'd7868, 16'd44010, 16'd23691, 16'd59330, 16'd8915, 16'd18417});
	test_expansion(128'h5bf5f4dbde4b6e4853e18c6069afbd3d, {16'd26684, 16'd49795, 16'd44471, 16'd21270, 16'd52396, 16'd27990, 16'd15344, 16'd1833, 16'd25848, 16'd31806, 16'd9450, 16'd12898, 16'd2341, 16'd29765, 16'd58088, 16'd60850, 16'd64936, 16'd43529, 16'd39677, 16'd59075, 16'd11631, 16'd31430, 16'd19443, 16'd7299, 16'd18072, 16'd39008});
	test_expansion(128'h3366f416cd6695d0e3a9d49a9af8a9aa, {16'd31963, 16'd11501, 16'd24127, 16'd13360, 16'd19265, 16'd12463, 16'd6449, 16'd49999, 16'd30713, 16'd9640, 16'd7723, 16'd55472, 16'd1679, 16'd32194, 16'd37896, 16'd27255, 16'd450, 16'd14426, 16'd45372, 16'd38654, 16'd15834, 16'd48233, 16'd22565, 16'd48001, 16'd45036, 16'd16845});
	test_expansion(128'h77a25ed180b5de091d8a744639abd81d, {16'd720, 16'd29052, 16'd16721, 16'd5886, 16'd46993, 16'd19114, 16'd31416, 16'd2309, 16'd31932, 16'd37650, 16'd37523, 16'd957, 16'd37021, 16'd53579, 16'd32358, 16'd16431, 16'd42833, 16'd36438, 16'd52331, 16'd39316, 16'd863, 16'd45758, 16'd21663, 16'd40229, 16'd35323, 16'd8982});
	test_expansion(128'h9735f55f8fd3a61de586cfcaa2e2c6bd, {16'd50884, 16'd42616, 16'd42760, 16'd13892, 16'd3721, 16'd2315, 16'd58357, 16'd7356, 16'd16798, 16'd55784, 16'd55451, 16'd33832, 16'd56766, 16'd19182, 16'd21255, 16'd58822, 16'd58733, 16'd30391, 16'd18257, 16'd16870, 16'd24151, 16'd24812, 16'd16510, 16'd27563, 16'd13541, 16'd31802});
	test_expansion(128'hf463e618e9c2e2395a1583cd5fe3a8eb, {16'd33507, 16'd3407, 16'd41661, 16'd1205, 16'd64603, 16'd44901, 16'd36117, 16'd33638, 16'd10624, 16'd11797, 16'd61730, 16'd62183, 16'd10844, 16'd18351, 16'd51547, 16'd37428, 16'd36762, 16'd46014, 16'd65532, 16'd5623, 16'd11310, 16'd64435, 16'd14106, 16'd34493, 16'd43315, 16'd1952});
	test_expansion(128'hbee13b3e85493a479812aec12d1f7a5a, {16'd9470, 16'd27090, 16'd57146, 16'd33206, 16'd7561, 16'd4051, 16'd34103, 16'd5947, 16'd38392, 16'd44004, 16'd48801, 16'd16567, 16'd41585, 16'd44380, 16'd18272, 16'd854, 16'd57235, 16'd9836, 16'd10372, 16'd37090, 16'd36250, 16'd1400, 16'd1348, 16'd54821, 16'd39284, 16'd34028});
	test_expansion(128'h0734b973a9304ba2e5e650b68c972ab6, {16'd14163, 16'd10484, 16'd44811, 16'd56401, 16'd2161, 16'd60329, 16'd41222, 16'd31641, 16'd35069, 16'd23703, 16'd27728, 16'd48581, 16'd20164, 16'd23857, 16'd53690, 16'd19307, 16'd42217, 16'd41135, 16'd20916, 16'd4636, 16'd40099, 16'd53895, 16'd40045, 16'd57327, 16'd2571, 16'd35148});
	test_expansion(128'hf4aaed0030ee9aac2e086cde6929c3d6, {16'd30960, 16'd7254, 16'd17566, 16'd44334, 16'd9398, 16'd63770, 16'd24149, 16'd29816, 16'd8382, 16'd25258, 16'd26820, 16'd39101, 16'd19491, 16'd2350, 16'd5357, 16'd22275, 16'd60786, 16'd54655, 16'd5540, 16'd5485, 16'd34500, 16'd40331, 16'd19697, 16'd25564, 16'd15339, 16'd29307});
	test_expansion(128'h538c197bb6c31227774b584e788257eb, {16'd33175, 16'd57821, 16'd31877, 16'd54794, 16'd63746, 16'd30884, 16'd13010, 16'd30432, 16'd55080, 16'd24546, 16'd30969, 16'd60012, 16'd38833, 16'd29131, 16'd53043, 16'd10469, 16'd59332, 16'd59103, 16'd18566, 16'd32596, 16'd8686, 16'd51073, 16'd40788, 16'd46657, 16'd39328, 16'd44133});
	test_expansion(128'h1879c5d5b81519879bff9b3af3e1d3ef, {16'd53260, 16'd7641, 16'd36700, 16'd37519, 16'd32758, 16'd42604, 16'd57076, 16'd3134, 16'd40391, 16'd58990, 16'd8274, 16'd55881, 16'd33186, 16'd57222, 16'd30733, 16'd65254, 16'd54482, 16'd62899, 16'd56934, 16'd58533, 16'd10375, 16'd63209, 16'd32175, 16'd29078, 16'd46840, 16'd42725});
	test_expansion(128'he8366c0ab026633cc84534dc4ea3ef88, {16'd34527, 16'd61543, 16'd15467, 16'd40259, 16'd38110, 16'd63680, 16'd8443, 16'd57229, 16'd891, 16'd62417, 16'd2694, 16'd12442, 16'd17225, 16'd64217, 16'd24327, 16'd49994, 16'd58562, 16'd27217, 16'd605, 16'd22549, 16'd55057, 16'd11956, 16'd37900, 16'd23245, 16'd27540, 16'd37293});
	test_expansion(128'hc7244533044ef6aaabbd07082c2232ec, {16'd9118, 16'd31880, 16'd58379, 16'd16849, 16'd27622, 16'd27446, 16'd40747, 16'd23636, 16'd44724, 16'd45447, 16'd11866, 16'd22291, 16'd4381, 16'd17228, 16'd29333, 16'd29204, 16'd22108, 16'd40866, 16'd56306, 16'd31784, 16'd41500, 16'd28329, 16'd32845, 16'd56955, 16'd31638, 16'd42559});
	test_expansion(128'h68b3c07d3a63c9fe4f787f4db4c15faf, {16'd5232, 16'd8496, 16'd3741, 16'd43767, 16'd32020, 16'd11643, 16'd10514, 16'd11083, 16'd55174, 16'd43650, 16'd63601, 16'd50409, 16'd35306, 16'd59724, 16'd34931, 16'd45810, 16'd12980, 16'd1036, 16'd38010, 16'd55448, 16'd38374, 16'd58466, 16'd65131, 16'd19185, 16'd33595, 16'd15088});
	test_expansion(128'h29d1e73ad8aae4edd5d012ba19c16a7c, {16'd28459, 16'd42061, 16'd36870, 16'd6768, 16'd42934, 16'd63022, 16'd14006, 16'd20795, 16'd3392, 16'd224, 16'd33329, 16'd52462, 16'd61326, 16'd12620, 16'd45672, 16'd30542, 16'd19352, 16'd60950, 16'd660, 16'd1419, 16'd61925, 16'd18694, 16'd33993, 16'd20836, 16'd49701, 16'd41895});
	test_expansion(128'h1e971bfcc05192c8015cf00da5aab781, {16'd14099, 16'd19143, 16'd34665, 16'd33916, 16'd58466, 16'd11167, 16'd8745, 16'd53795, 16'd47504, 16'd63000, 16'd59376, 16'd32408, 16'd35265, 16'd12727, 16'd63033, 16'd48840, 16'd5846, 16'd45745, 16'd65160, 16'd47821, 16'd35267, 16'd34081, 16'd53149, 16'd59705, 16'd30979, 16'd54268});
	test_expansion(128'hd8f1fe3f0ee70ffe79891523d21fb89f, {16'd55072, 16'd6015, 16'd21084, 16'd59267, 16'd34117, 16'd29685, 16'd56054, 16'd41342, 16'd15790, 16'd5865, 16'd63691, 16'd44973, 16'd54576, 16'd8045, 16'd53071, 16'd15274, 16'd41799, 16'd14895, 16'd19733, 16'd13246, 16'd48033, 16'd44599, 16'd50756, 16'd5325, 16'd13986, 16'd61040});
	test_expansion(128'hf1856075f5bf6eae560dd5abda0c8efb, {16'd42948, 16'd39514, 16'd33406, 16'd56732, 16'd25626, 16'd29195, 16'd19825, 16'd64187, 16'd39747, 16'd21510, 16'd55861, 16'd42779, 16'd25891, 16'd33360, 16'd11814, 16'd23902, 16'd42463, 16'd9293, 16'd44657, 16'd53923, 16'd45646, 16'd59929, 16'd35779, 16'd16160, 16'd53277, 16'd16626});
	test_expansion(128'h268d4bc41f3f97663fe6fb6f08810fef, {16'd50559, 16'd36960, 16'd42670, 16'd43226, 16'd41030, 16'd8277, 16'd49850, 16'd6678, 16'd34419, 16'd27977, 16'd20721, 16'd43171, 16'd54050, 16'd39279, 16'd2849, 16'd75, 16'd63752, 16'd46448, 16'd52166, 16'd55316, 16'd12837, 16'd50632, 16'd7950, 16'd2367, 16'd20874, 16'd22846});
	test_expansion(128'h0ed7a58859bdda315330e4ee95b01702, {16'd38595, 16'd53056, 16'd45887, 16'd24538, 16'd56766, 16'd62010, 16'd35937, 16'd9303, 16'd23072, 16'd29545, 16'd17995, 16'd22134, 16'd44028, 16'd31384, 16'd42212, 16'd22542, 16'd48055, 16'd15987, 16'd64701, 16'd56345, 16'd45409, 16'd124, 16'd2437, 16'd11897, 16'd4700, 16'd52790});
	test_expansion(128'had842d0d41852b53812a40a7e096e2c0, {16'd57505, 16'd32208, 16'd52585, 16'd28593, 16'd17204, 16'd55034, 16'd34987, 16'd63146, 16'd25361, 16'd58835, 16'd16658, 16'd2236, 16'd20274, 16'd56989, 16'd17846, 16'd54937, 16'd8286, 16'd5443, 16'd26331, 16'd34218, 16'd62572, 16'd54535, 16'd26046, 16'd1370, 16'd34605, 16'd45000});
	test_expansion(128'h92050098da0e5d0f1c3d2b101952bede, {16'd42655, 16'd17905, 16'd18015, 16'd48895, 16'd52432, 16'd38382, 16'd44531, 16'd2336, 16'd59001, 16'd56840, 16'd11292, 16'd1247, 16'd14264, 16'd22162, 16'd54355, 16'd43915, 16'd10940, 16'd18584, 16'd52387, 16'd34057, 16'd23309, 16'd20452, 16'd26103, 16'd47483, 16'd60432, 16'd6937});
	test_expansion(128'hd86c47c5ccebba22494401381d416324, {16'd63078, 16'd19183, 16'd49981, 16'd47008, 16'd42127, 16'd57975, 16'd54828, 16'd26283, 16'd5270, 16'd35281, 16'd44195, 16'd3667, 16'd32343, 16'd9401, 16'd52517, 16'd17250, 16'd33505, 16'd8435, 16'd58431, 16'd44791, 16'd21741, 16'd60486, 16'd28540, 16'd62042, 16'd29041, 16'd61363});
	test_expansion(128'h2a11db356b2f429e23b47301bebb1d98, {16'd21644, 16'd41884, 16'd16129, 16'd56955, 16'd4510, 16'd41358, 16'd11423, 16'd29142, 16'd25395, 16'd24535, 16'd55882, 16'd42953, 16'd24594, 16'd24808, 16'd42939, 16'd6410, 16'd48077, 16'd57510, 16'd29710, 16'd10120, 16'd23863, 16'd54519, 16'd6141, 16'd44504, 16'd54722, 16'd14445});
	test_expansion(128'h77c5ecf46266c88eb36adc8f7f50de24, {16'd17425, 16'd40470, 16'd49757, 16'd12618, 16'd55540, 16'd31414, 16'd21995, 16'd6525, 16'd24603, 16'd22072, 16'd58357, 16'd14221, 16'd59227, 16'd28178, 16'd28826, 16'd39460, 16'd23237, 16'd8885, 16'd44825, 16'd34214, 16'd26354, 16'd54215, 16'd10994, 16'd26805, 16'd54405, 16'd23197});
	test_expansion(128'h50a66f36c2864dee68cd7e3847e988da, {16'd51832, 16'd62780, 16'd62255, 16'd23662, 16'd11511, 16'd49715, 16'd52169, 16'd5172, 16'd28302, 16'd4405, 16'd29676, 16'd55789, 16'd46583, 16'd43310, 16'd9089, 16'd59332, 16'd29513, 16'd18809, 16'd22568, 16'd34412, 16'd18080, 16'd23420, 16'd49199, 16'd25557, 16'd52871, 16'd61390});
	test_expansion(128'hf725f8b0269a7535209e607b7836c8da, {16'd52231, 16'd17301, 16'd45628, 16'd33757, 16'd24185, 16'd14784, 16'd45233, 16'd15778, 16'd31781, 16'd24744, 16'd36998, 16'd36185, 16'd9174, 16'd13580, 16'd41854, 16'd43753, 16'd58105, 16'd2871, 16'd57390, 16'd53587, 16'd39536, 16'd43745, 16'd36759, 16'd11683, 16'd50242, 16'd14655});
	test_expansion(128'ha3e002f57ef3badcbf88f220cc1ca22a, {16'd20698, 16'd29195, 16'd23965, 16'd22956, 16'd34795, 16'd47130, 16'd18642, 16'd13761, 16'd9252, 16'd8328, 16'd28138, 16'd7131, 16'd39074, 16'd22510, 16'd38995, 16'd19038, 16'd62295, 16'd20214, 16'd51058, 16'd30432, 16'd49712, 16'd50082, 16'd64519, 16'd34660, 16'd35800, 16'd30381});
	test_expansion(128'hd971a8165146c12e343a541281906be2, {16'd20399, 16'd25355, 16'd10213, 16'd54558, 16'd16117, 16'd15628, 16'd23356, 16'd25133, 16'd40678, 16'd27865, 16'd44022, 16'd19291, 16'd14571, 16'd52004, 16'd23180, 16'd64895, 16'd16404, 16'd54386, 16'd30850, 16'd45839, 16'd26486, 16'd28550, 16'd16381, 16'd52061, 16'd36139, 16'd54066});
	test_expansion(128'h2c156a07bd6c26190e5c70b04ba27bca, {16'd40211, 16'd27369, 16'd26133, 16'd17434, 16'd58065, 16'd16820, 16'd48873, 16'd11382, 16'd26633, 16'd34429, 16'd32167, 16'd35354, 16'd20644, 16'd53378, 16'd5589, 16'd1280, 16'd40073, 16'd36953, 16'd33685, 16'd39731, 16'd16279, 16'd40976, 16'd19310, 16'd55932, 16'd24944, 16'd50854});
	test_expansion(128'h734d4583a6fa94b8efc5401de1d8c43f, {16'd6582, 16'd10672, 16'd19686, 16'd41508, 16'd59571, 16'd2523, 16'd58646, 16'd65500, 16'd45455, 16'd5895, 16'd51011, 16'd37671, 16'd46593, 16'd27896, 16'd39546, 16'd14695, 16'd37996, 16'd40587, 16'd24379, 16'd14671, 16'd3182, 16'd52977, 16'd55151, 16'd42, 16'd53433, 16'd56139});
	test_expansion(128'hf4b68d6d7e8c88cf9ccf4576be7a77be, {16'd11874, 16'd60317, 16'd21398, 16'd62754, 16'd61022, 16'd54488, 16'd54604, 16'd8552, 16'd41253, 16'd47577, 16'd34664, 16'd12113, 16'd35562, 16'd60962, 16'd7807, 16'd42383, 16'd5718, 16'd56875, 16'd56566, 16'd24335, 16'd54227, 16'd47473, 16'd9771, 16'd1644, 16'd45288, 16'd58578});
	test_expansion(128'h4d09bf7ef93fe934e9ae0077d54224c8, {16'd25850, 16'd14443, 16'd55879, 16'd16221, 16'd60583, 16'd51363, 16'd26511, 16'd19138, 16'd49635, 16'd50580, 16'd13468, 16'd10059, 16'd5900, 16'd53128, 16'd956, 16'd33989, 16'd56379, 16'd5808, 16'd60056, 16'd23616, 16'd45639, 16'd58698, 16'd40815, 16'd26381, 16'd10375, 16'd44405});
	test_expansion(128'hb450c34f610636ccb31464a864021796, {16'd3988, 16'd20909, 16'd1275, 16'd33178, 16'd29631, 16'd9793, 16'd51689, 16'd13157, 16'd15682, 16'd17405, 16'd37151, 16'd45850, 16'd17604, 16'd14026, 16'd2125, 16'd55144, 16'd51034, 16'd30899, 16'd23826, 16'd43136, 16'd3126, 16'd34553, 16'd50499, 16'd51462, 16'd43424, 16'd65386});
	test_expansion(128'hac0a15d270f0de7be81002eca283b69b, {16'd61245, 16'd61791, 16'd40658, 16'd62, 16'd2217, 16'd45086, 16'd11580, 16'd24784, 16'd39531, 16'd20496, 16'd45103, 16'd21233, 16'd37478, 16'd36599, 16'd370, 16'd29132, 16'd33465, 16'd13509, 16'd37502, 16'd35147, 16'd64936, 16'd17792, 16'd35922, 16'd64132, 16'd27655, 16'd24363});
	test_expansion(128'hf6444eece376fef81491c669317beb04, {16'd52953, 16'd40247, 16'd60784, 16'd42307, 16'd25816, 16'd34730, 16'd56402, 16'd50800, 16'd40443, 16'd25592, 16'd55175, 16'd28861, 16'd33853, 16'd10339, 16'd30097, 16'd22567, 16'd52705, 16'd44148, 16'd39296, 16'd60440, 16'd26323, 16'd47285, 16'd20155, 16'd62717, 16'd21724, 16'd50768});
	test_expansion(128'hf2bf47698669fd7ee6cca5b15a7ae21e, {16'd50838, 16'd24646, 16'd19625, 16'd3455, 16'd30873, 16'd22842, 16'd28685, 16'd7355, 16'd15469, 16'd53125, 16'd46604, 16'd24530, 16'd46198, 16'd7753, 16'd55597, 16'd39007, 16'd24725, 16'd5794, 16'd30109, 16'd42306, 16'd36504, 16'd60227, 16'd50863, 16'd43257, 16'd39037, 16'd48207});
	test_expansion(128'h72a3e7cce21f1a5b81eeae1ceed3c388, {16'd20906, 16'd53908, 16'd16989, 16'd12022, 16'd35394, 16'd23073, 16'd23047, 16'd1923, 16'd21443, 16'd24029, 16'd13322, 16'd2995, 16'd62779, 16'd53545, 16'd40503, 16'd24687, 16'd60890, 16'd33153, 16'd878, 16'd61886, 16'd2937, 16'd43209, 16'd44439, 16'd63209, 16'd10710, 16'd55092});
	test_expansion(128'h0dc3117f8fa58122f9e89aa538e886f9, {16'd31109, 16'd37298, 16'd12622, 16'd61170, 16'd62572, 16'd9849, 16'd6938, 16'd61594, 16'd46362, 16'd48071, 16'd48842, 16'd24986, 16'd34989, 16'd38347, 16'd49868, 16'd54121, 16'd56028, 16'd40680, 16'd61759, 16'd28701, 16'd38301, 16'd9685, 16'd25069, 16'd370, 16'd59615, 16'd24143});
	test_expansion(128'h6d7dbfb5da41b75c58acdea4e8438265, {16'd46830, 16'd18282, 16'd17820, 16'd54135, 16'd58950, 16'd16263, 16'd48564, 16'd4506, 16'd60744, 16'd28117, 16'd11110, 16'd19368, 16'd57666, 16'd26071, 16'd50825, 16'd30148, 16'd10923, 16'd62482, 16'd43486, 16'd15354, 16'd52943, 16'd61170, 16'd47470, 16'd58925, 16'd42380, 16'd321});
	test_expansion(128'hd68ff13199128b9f0bb2530d459be362, {16'd53883, 16'd32293, 16'd20362, 16'd62136, 16'd11939, 16'd64374, 16'd36107, 16'd54568, 16'd61941, 16'd6877, 16'd42372, 16'd27724, 16'd63355, 16'd54093, 16'd62384, 16'd53034, 16'd14706, 16'd27417, 16'd6800, 16'd51464, 16'd56065, 16'd31864, 16'd5088, 16'd24483, 16'd50024, 16'd21160});
	test_expansion(128'h7b92a382c2cf1090d75e5d005b41ad41, {16'd45679, 16'd12441, 16'd7194, 16'd21183, 16'd37452, 16'd35311, 16'd52079, 16'd37477, 16'd37700, 16'd36268, 16'd54673, 16'd41927, 16'd30259, 16'd26145, 16'd55519, 16'd4502, 16'd15793, 16'd33065, 16'd62799, 16'd58491, 16'd15375, 16'd32952, 16'd8135, 16'd37588, 16'd59812, 16'd19140});
	test_expansion(128'h5cd956a2253df5d2fc4caeaab74c3e8c, {16'd62183, 16'd38279, 16'd8004, 16'd22826, 16'd51728, 16'd22663, 16'd53655, 16'd2997, 16'd46432, 16'd39241, 16'd7006, 16'd26687, 16'd40, 16'd6398, 16'd62545, 16'd46252, 16'd39682, 16'd30841, 16'd378, 16'd25889, 16'd64124, 16'd12526, 16'd31240, 16'd12251, 16'd47005, 16'd6111});
	test_expansion(128'h4d0458acc6d6a2aabfd0643aa6bfcb89, {16'd44600, 16'd64775, 16'd59878, 16'd29690, 16'd48803, 16'd57478, 16'd44481, 16'd7644, 16'd811, 16'd15642, 16'd38450, 16'd51860, 16'd56124, 16'd46576, 16'd57183, 16'd31348, 16'd55468, 16'd37667, 16'd14874, 16'd11440, 16'd37811, 16'd56437, 16'd56565, 16'd7932, 16'd32405, 16'd52093});
	test_expansion(128'hbf6e61e8aec9c420641b36b1a867760d, {16'd26457, 16'd23194, 16'd44537, 16'd60337, 16'd35289, 16'd40181, 16'd20614, 16'd44531, 16'd32714, 16'd28962, 16'd3993, 16'd54442, 16'd46755, 16'd39426, 16'd24500, 16'd12921, 16'd940, 16'd30387, 16'd35617, 16'd13557, 16'd47195, 16'd1969, 16'd20891, 16'd6152, 16'd52534, 16'd56979});
	test_expansion(128'hfa9520f622d899085f5c87a518d0129c, {16'd63530, 16'd5803, 16'd26057, 16'd44309, 16'd45172, 16'd14078, 16'd24895, 16'd30416, 16'd61367, 16'd21874, 16'd1575, 16'd57671, 16'd19246, 16'd34669, 16'd5139, 16'd42684, 16'd11843, 16'd45792, 16'd17225, 16'd52953, 16'd57011, 16'd19212, 16'd50273, 16'd17160, 16'd19365, 16'd53194});
	test_expansion(128'ha7966711b85cecb04d79d256d3e60029, {16'd12277, 16'd59345, 16'd49367, 16'd38065, 16'd123, 16'd54922, 16'd28497, 16'd41553, 16'd39808, 16'd40361, 16'd46176, 16'd15460, 16'd10042, 16'd55382, 16'd43718, 16'd49659, 16'd29229, 16'd61904, 16'd39145, 16'd15370, 16'd41771, 16'd64787, 16'd52365, 16'd6564, 16'd33779, 16'd14733});
	test_expansion(128'ha7db07067e9b356d45bf9bfd4898ff73, {16'd56506, 16'd33244, 16'd16743, 16'd184, 16'd16246, 16'd42887, 16'd18307, 16'd12889, 16'd32140, 16'd58337, 16'd37070, 16'd64296, 16'd32219, 16'd64710, 16'd2985, 16'd52554, 16'd45680, 16'd57867, 16'd44352, 16'd43289, 16'd29614, 16'd10948, 16'd18872, 16'd58441, 16'd15513, 16'd40275});
	test_expansion(128'h6a5533d5a0c067dcc079bafc185b17b4, {16'd48522, 16'd44288, 16'd62634, 16'd48730, 16'd9555, 16'd18050, 16'd43394, 16'd53465, 16'd38809, 16'd23962, 16'd26559, 16'd61409, 16'd21656, 16'd47078, 16'd37077, 16'd50320, 16'd37158, 16'd56965, 16'd2087, 16'd54214, 16'd42359, 16'd29954, 16'd43914, 16'd988, 16'd37592, 16'd4490});
	test_expansion(128'h144bb71f17539f6b3a3d9398e5e3e53e, {16'd29329, 16'd59606, 16'd55941, 16'd49151, 16'd36689, 16'd17456, 16'd3219, 16'd5143, 16'd54932, 16'd34660, 16'd30222, 16'd14279, 16'd94, 16'd60665, 16'd57029, 16'd65157, 16'd49242, 16'd39689, 16'd347, 16'd59616, 16'd5367, 16'd21892, 16'd45935, 16'd32326, 16'd44868, 16'd8952});
	test_expansion(128'h115e28da999ba168313e2e4cf88565d5, {16'd48544, 16'd32591, 16'd3253, 16'd52991, 16'd13482, 16'd40882, 16'd36459, 16'd131, 16'd42972, 16'd31969, 16'd61358, 16'd16746, 16'd45933, 16'd51434, 16'd45290, 16'd4049, 16'd34807, 16'd60295, 16'd37458, 16'd45610, 16'd29405, 16'd40606, 16'd25352, 16'd23753, 16'd29401, 16'd16931});
	test_expansion(128'h202fc207210961939a7ddcdd7090578c, {16'd23505, 16'd363, 16'd11323, 16'd7920, 16'd7649, 16'd49545, 16'd19337, 16'd29548, 16'd27125, 16'd27102, 16'd3481, 16'd40074, 16'd54954, 16'd14939, 16'd31122, 16'd32727, 16'd58729, 16'd48401, 16'd61353, 16'd45565, 16'd22492, 16'd31297, 16'd37546, 16'd60237, 16'd38550, 16'd39476});
	test_expansion(128'h4c330a84145a75c98049a9f672107340, {16'd5924, 16'd27845, 16'd9392, 16'd27170, 16'd8403, 16'd36587, 16'd6693, 16'd35663, 16'd25641, 16'd56912, 16'd23715, 16'd64481, 16'd12056, 16'd5777, 16'd5672, 16'd10607, 16'd57002, 16'd49703, 16'd48825, 16'd18446, 16'd3359, 16'd42265, 16'd49946, 16'd3961, 16'd39618, 16'd35933});
	test_expansion(128'hf05af7f6af9adfe01f24fdf49fb6e5e6, {16'd55788, 16'd64703, 16'd9232, 16'd39628, 16'd25018, 16'd40605, 16'd3023, 16'd60628, 16'd46147, 16'd20228, 16'd31514, 16'd47492, 16'd58413, 16'd47867, 16'd44384, 16'd36039, 16'd17578, 16'd10705, 16'd13040, 16'd23301, 16'd39891, 16'd39847, 16'd1602, 16'd31070, 16'd4542, 16'd60828});
	test_expansion(128'heaf92828bef5d3fe4b64ad149111e9f8, {16'd16078, 16'd23855, 16'd4322, 16'd17886, 16'd18887, 16'd19444, 16'd5703, 16'd24404, 16'd25226, 16'd24984, 16'd57564, 16'd34083, 16'd40141, 16'd45147, 16'd4637, 16'd54340, 16'd44296, 16'd40588, 16'd32624, 16'd19600, 16'd44965, 16'd44191, 16'd49229, 16'd15912, 16'd56859, 16'd34097});
	test_expansion(128'h88af44b31915d042d095fc8bdb4c68f6, {16'd60539, 16'd45669, 16'd30388, 16'd30787, 16'd27772, 16'd1309, 16'd20925, 16'd47479, 16'd38593, 16'd46272, 16'd61850, 16'd29821, 16'd24026, 16'd18775, 16'd56033, 16'd27770, 16'd9300, 16'd21138, 16'd15887, 16'd18764, 16'd32435, 16'd2312, 16'd6212, 16'd10261, 16'd41326, 16'd55141});
	test_expansion(128'hc8f25d6775fbee3694fb602f9c79a50c, {16'd64946, 16'd26705, 16'd15229, 16'd38061, 16'd54073, 16'd12872, 16'd35342, 16'd19713, 16'd11444, 16'd47, 16'd64030, 16'd52254, 16'd39977, 16'd410, 16'd61209, 16'd60353, 16'd749, 16'd60148, 16'd11960, 16'd27471, 16'd20809, 16'd51986, 16'd21384, 16'd8110, 16'd40563, 16'd37434});
	test_expansion(128'h67220ed5a7de9f0c7761005732438b3a, {16'd17139, 16'd5884, 16'd46246, 16'd9237, 16'd400, 16'd18263, 16'd49181, 16'd18175, 16'd56569, 16'd51954, 16'd59230, 16'd29371, 16'd29268, 16'd23698, 16'd14200, 16'd876, 16'd59563, 16'd58347, 16'd32640, 16'd33454, 16'd14835, 16'd36326, 16'd10212, 16'd25302, 16'd61095, 16'd58120});
	test_expansion(128'hfab7618008dd0f2686b261588bbdf7fc, {16'd1202, 16'd16940, 16'd10144, 16'd5535, 16'd41243, 16'd25625, 16'd12663, 16'd39212, 16'd57625, 16'd1341, 16'd54490, 16'd1618, 16'd44705, 16'd55110, 16'd9411, 16'd2493, 16'd36742, 16'd18599, 16'd44403, 16'd7521, 16'd29806, 16'd44841, 16'd12264, 16'd16711, 16'd15466, 16'd34205});
	test_expansion(128'ha9e09c4b17bd27864c68636d7f2e3472, {16'd13501, 16'd51777, 16'd16247, 16'd6584, 16'd21338, 16'd45182, 16'd46701, 16'd57114, 16'd8377, 16'd20508, 16'd873, 16'd37848, 16'd61476, 16'd7210, 16'd45461, 16'd2477, 16'd49895, 16'd60284, 16'd4364, 16'd13573, 16'd8671, 16'd63024, 16'd60180, 16'd4423, 16'd12279, 16'd60675});
	test_expansion(128'ha72d483aa3bf6a689763727946d1a7cd, {16'd12934, 16'd64695, 16'd4676, 16'd56986, 16'd47950, 16'd50352, 16'd13628, 16'd36537, 16'd35683, 16'd37091, 16'd28015, 16'd734, 16'd23302, 16'd28501, 16'd13286, 16'd28030, 16'd37498, 16'd48717, 16'd51988, 16'd30827, 16'd42235, 16'd58315, 16'd24402, 16'd41449, 16'd8929, 16'd65276});
	test_expansion(128'hd98f7e14fe318ab67b81440b915f0510, {16'd39901, 16'd36851, 16'd43920, 16'd56190, 16'd57113, 16'd47884, 16'd14805, 16'd38340, 16'd61843, 16'd39011, 16'd5776, 16'd53117, 16'd6216, 16'd22179, 16'd24733, 16'd50401, 16'd60455, 16'd30567, 16'd11616, 16'd37058, 16'd37792, 16'd29721, 16'd57564, 16'd63577, 16'd3923, 16'd62400});
	test_expansion(128'hfab8e9439ee315d525bf5f84908fc511, {16'd31690, 16'd38887, 16'd28738, 16'd56782, 16'd22017, 16'd20025, 16'd64985, 16'd4310, 16'd47259, 16'd4034, 16'd23885, 16'd10659, 16'd35904, 16'd5509, 16'd20120, 16'd43225, 16'd17795, 16'd37163, 16'd50712, 16'd11024, 16'd24905, 16'd43526, 16'd40607, 16'd37265, 16'd37348, 16'd59257});
	test_expansion(128'haeccd1158280835fc27838084c6e6a38, {16'd16162, 16'd43030, 16'd55429, 16'd30686, 16'd49561, 16'd60125, 16'd19446, 16'd19798, 16'd60086, 16'd50926, 16'd7705, 16'd63955, 16'd24334, 16'd11041, 16'd35005, 16'd52439, 16'd64079, 16'd45885, 16'd16458, 16'd61056, 16'd34738, 16'd41772, 16'd19573, 16'd59424, 16'd16315, 16'd43587});
	test_expansion(128'hf06381a5c975cf388ce026433fb44b56, {16'd16730, 16'd24085, 16'd63494, 16'd44112, 16'd49710, 16'd4390, 16'd43496, 16'd16556, 16'd942, 16'd18165, 16'd11970, 16'd30632, 16'd60434, 16'd15348, 16'd2909, 16'd35422, 16'd44560, 16'd35373, 16'd57406, 16'd7314, 16'd6627, 16'd2665, 16'd12884, 16'd51458, 16'd34709, 16'd22106});
	test_expansion(128'h7b9847a2c102f0694b0c64563a38badf, {16'd54123, 16'd54211, 16'd46186, 16'd61681, 16'd55709, 16'd10880, 16'd29520, 16'd45587, 16'd24216, 16'd12634, 16'd10674, 16'd53524, 16'd26627, 16'd53196, 16'd51467, 16'd37333, 16'd14447, 16'd56233, 16'd39586, 16'd58516, 16'd11278, 16'd35095, 16'd61158, 16'd32203, 16'd46382, 16'd41858});
	test_expansion(128'h497daa47ccca422e58d86c8bc6c51dad, {16'd32798, 16'd31971, 16'd4401, 16'd56664, 16'd31962, 16'd24839, 16'd65218, 16'd30247, 16'd38091, 16'd1794, 16'd29686, 16'd35376, 16'd16471, 16'd5278, 16'd19738, 16'd46672, 16'd43311, 16'd17427, 16'd45780, 16'd53032, 16'd28298, 16'd17947, 16'd52975, 16'd27712, 16'd47036, 16'd46455});
	test_expansion(128'h19b8bd6ed9cabb1be9fc84a2730e7a79, {16'd45180, 16'd6163, 16'd10720, 16'd5372, 16'd10439, 16'd20607, 16'd62797, 16'd976, 16'd22581, 16'd2862, 16'd32635, 16'd10069, 16'd26464, 16'd40994, 16'd3998, 16'd48242, 16'd65160, 16'd50119, 16'd23893, 16'd56584, 16'd8190, 16'd8698, 16'd49209, 16'd35766, 16'd1393, 16'd15575});
	test_expansion(128'h1e192349c6810e077dfb59d33d350418, {16'd15058, 16'd54887, 16'd27402, 16'd48914, 16'd54880, 16'd32722, 16'd7666, 16'd8080, 16'd10455, 16'd47014, 16'd9284, 16'd46099, 16'd32651, 16'd37010, 16'd22079, 16'd42286, 16'd61169, 16'd60073, 16'd61730, 16'd21285, 16'd37124, 16'd51933, 16'd26254, 16'd8751, 16'd44622, 16'd21795});
	test_expansion(128'hfbe4fd14158036bee57f1ba3edf67242, {16'd21741, 16'd26168, 16'd59971, 16'd64461, 16'd39008, 16'd33932, 16'd32397, 16'd44542, 16'd32225, 16'd57563, 16'd380, 16'd3879, 16'd15091, 16'd49095, 16'd50144, 16'd22192, 16'd40365, 16'd30625, 16'd47708, 16'd56255, 16'd64634, 16'd683, 16'd47979, 16'd16582, 16'd10484, 16'd49000});
	test_expansion(128'hfaad77e40493d05995d280d2c5e1a1b8, {16'd35846, 16'd15003, 16'd359, 16'd57194, 16'd8357, 16'd19786, 16'd56231, 16'd63026, 16'd8020, 16'd28360, 16'd41491, 16'd47617, 16'd32120, 16'd28808, 16'd43315, 16'd36242, 16'd54616, 16'd12595, 16'd33762, 16'd39875, 16'd52905, 16'd58627, 16'd16320, 16'd56388, 16'd12471, 16'd22586});
	test_expansion(128'hf9409a5a9f226de4b0492cf39537d44f, {16'd24926, 16'd62089, 16'd4257, 16'd8790, 16'd45415, 16'd55521, 16'd61820, 16'd53944, 16'd1168, 16'd39763, 16'd31885, 16'd5172, 16'd59196, 16'd51691, 16'd64736, 16'd35381, 16'd47185, 16'd16082, 16'd36497, 16'd36148, 16'd50154, 16'd34605, 16'd15369, 16'd20905, 16'd8966, 16'd16745});
	test_expansion(128'hb8c675ef0128561e5281df243ff90caf, {16'd44862, 16'd9864, 16'd9548, 16'd12534, 16'd10905, 16'd28968, 16'd24578, 16'd2751, 16'd46158, 16'd12438, 16'd29324, 16'd18431, 16'd30583, 16'd3162, 16'd36623, 16'd37853, 16'd39504, 16'd56628, 16'd34751, 16'd63201, 16'd50456, 16'd14206, 16'd17355, 16'd41877, 16'd45337, 16'd1962});
	test_expansion(128'h1ed5f8cb8cb88d457a8f9bc350de31ce, {16'd59649, 16'd49650, 16'd869, 16'd35686, 16'd35571, 16'd64116, 16'd37128, 16'd29268, 16'd2165, 16'd22500, 16'd22572, 16'd20283, 16'd2670, 16'd46267, 16'd58429, 16'd53625, 16'd60969, 16'd40165, 16'd25914, 16'd64911, 16'd50503, 16'd5225, 16'd15878, 16'd12843, 16'd455, 16'd19483});
	test_expansion(128'he5f9cae06938fc6a5eddb7a7f238c59c, {16'd11546, 16'd38886, 16'd15204, 16'd8387, 16'd34806, 16'd2902, 16'd43130, 16'd14889, 16'd14115, 16'd8731, 16'd60731, 16'd54615, 16'd8597, 16'd58848, 16'd57240, 16'd7854, 16'd58814, 16'd32332, 16'd26096, 16'd12662, 16'd42715, 16'd57958, 16'd31272, 16'd26970, 16'd65305, 16'd13526});
	test_expansion(128'haa783d20c06ba18fe34a226174606047, {16'd29931, 16'd64871, 16'd9345, 16'd47147, 16'd11366, 16'd48170, 16'd4939, 16'd18044, 16'd11154, 16'd29482, 16'd42164, 16'd24309, 16'd28057, 16'd45473, 16'd43292, 16'd40488, 16'd33060, 16'd52610, 16'd8376, 16'd42362, 16'd29761, 16'd20629, 16'd20809, 16'd9415, 16'd57449, 16'd33321});
	test_expansion(128'hc8e0bc28dd4f63d24e94112ef10484fe, {16'd54561, 16'd20460, 16'd42441, 16'd16824, 16'd61774, 16'd43718, 16'd50, 16'd21677, 16'd37058, 16'd4454, 16'd52520, 16'd58642, 16'd5392, 16'd43425, 16'd55436, 16'd7652, 16'd27924, 16'd18023, 16'd36636, 16'd61471, 16'd50905, 16'd40299, 16'd1488, 16'd16661, 16'd30492, 16'd54152});
	test_expansion(128'h753fc994fda0994a4b6f2d43ff0f2858, {16'd29200, 16'd20745, 16'd45779, 16'd32983, 16'd34053, 16'd11881, 16'd5003, 16'd25103, 16'd3226, 16'd3618, 16'd49591, 16'd52941, 16'd64398, 16'd44591, 16'd62840, 16'd36013, 16'd45974, 16'd59305, 16'd16295, 16'd29793, 16'd63852, 16'd47031, 16'd44473, 16'd3327, 16'd38713, 16'd30194});
	test_expansion(128'h2ee8085ae97712110d6b0bcac9b94503, {16'd15403, 16'd52434, 16'd23168, 16'd10136, 16'd44981, 16'd14750, 16'd38606, 16'd24211, 16'd44342, 16'd45990, 16'd52563, 16'd34583, 16'd14738, 16'd50570, 16'd40666, 16'd60838, 16'd20444, 16'd18381, 16'd2350, 16'd43278, 16'd8263, 16'd54692, 16'd59151, 16'd13377, 16'd25253, 16'd49014});
	test_expansion(128'h3ed29c59c80cb2fcfb47378fbe5ed588, {16'd33691, 16'd64656, 16'd26354, 16'd26136, 16'd17480, 16'd15128, 16'd8357, 16'd57986, 16'd12190, 16'd58246, 16'd12404, 16'd3148, 16'd42501, 16'd5975, 16'd50852, 16'd53861, 16'd13509, 16'd47667, 16'd61330, 16'd36147, 16'd53377, 16'd42814, 16'd26220, 16'd10003, 16'd27803, 16'd31982});
	test_expansion(128'h62b5c08efbc0274d18b3cc203e61182c, {16'd9429, 16'd21868, 16'd1154, 16'd22580, 16'd18329, 16'd49352, 16'd29616, 16'd25033, 16'd835, 16'd26762, 16'd48857, 16'd24220, 16'd33276, 16'd51105, 16'd49964, 16'd61584, 16'd24894, 16'd17161, 16'd23214, 16'd12821, 16'd20872, 16'd9839, 16'd59539, 16'd14911, 16'd57957, 16'd37449});
	test_expansion(128'h6299c1ae7ccd610b5e576fe09ca1c25c, {16'd55906, 16'd18370, 16'd40930, 16'd27545, 16'd15401, 16'd56789, 16'd12173, 16'd60194, 16'd21313, 16'd43677, 16'd12722, 16'd17732, 16'd61629, 16'd12693, 16'd46126, 16'd9391, 16'd2223, 16'd6968, 16'd65230, 16'd55743, 16'd43210, 16'd15222, 16'd5468, 16'd64978, 16'd43448, 16'd33078});
	test_expansion(128'hca4a4785204e430d5250ec116a20a630, {16'd35157, 16'd61392, 16'd26601, 16'd30036, 16'd9215, 16'd59723, 16'd17857, 16'd15752, 16'd33706, 16'd3190, 16'd5836, 16'd30025, 16'd37440, 16'd35369, 16'd14737, 16'd43879, 16'd25746, 16'd36236, 16'd37877, 16'd16620, 16'd50136, 16'd37040, 16'd50309, 16'd43380, 16'd31122, 16'd6807});
	test_expansion(128'h30baed6893f550b4fa3ce7a69f2a3039, {16'd60509, 16'd9997, 16'd19489, 16'd27408, 16'd50608, 16'd15686, 16'd18400, 16'd33257, 16'd52114, 16'd3064, 16'd9866, 16'd55504, 16'd24988, 16'd49477, 16'd23144, 16'd43074, 16'd54555, 16'd39385, 16'd65155, 16'd50317, 16'd29350, 16'd10621, 16'd58886, 16'd42810, 16'd23527, 16'd38814});
	test_expansion(128'h4e136ed073c673e6d3509be966828d96, {16'd51122, 16'd965, 16'd17557, 16'd44692, 16'd26672, 16'd63942, 16'd43128, 16'd18488, 16'd3378, 16'd52228, 16'd4361, 16'd51642, 16'd63304, 16'd5859, 16'd26849, 16'd19035, 16'd10111, 16'd56632, 16'd33840, 16'd34934, 16'd39713, 16'd41359, 16'd8591, 16'd31494, 16'd54265, 16'd42159});
	test_expansion(128'hcb5ed240a7a8a6ed0e1bf273fe1ef5d4, {16'd20315, 16'd42551, 16'd58060, 16'd33489, 16'd51453, 16'd57177, 16'd32068, 16'd40893, 16'd50373, 16'd5253, 16'd29780, 16'd33273, 16'd35872, 16'd23028, 16'd55322, 16'd31469, 16'd30273, 16'd11703, 16'd36319, 16'd64546, 16'd52419, 16'd40085, 16'd13824, 16'd41247, 16'd32566, 16'd62623});
	test_expansion(128'h7daa9daeba887827f64c0f4ce0f9e27d, {16'd2221, 16'd8866, 16'd31879, 16'd30561, 16'd22565, 16'd15740, 16'd41805, 16'd42965, 16'd51175, 16'd32015, 16'd28139, 16'd34455, 16'd35925, 16'd17028, 16'd29542, 16'd12100, 16'd23525, 16'd59010, 16'd51572, 16'd43419, 16'd62787, 16'd41399, 16'd7833, 16'd38000, 16'd30462, 16'd55633});
	test_expansion(128'h197afe60fa221f48e85657f316a14b91, {16'd57786, 16'd41439, 16'd50517, 16'd50824, 16'd33727, 16'd61274, 16'd62335, 16'd43308, 16'd30953, 16'd149, 16'd57647, 16'd46734, 16'd22286, 16'd31844, 16'd5119, 16'd2961, 16'd30465, 16'd20911, 16'd30371, 16'd12199, 16'd28846, 16'd41983, 16'd20795, 16'd49209, 16'd9077, 16'd48338});
	test_expansion(128'h248a44c0ad270435a77619698026e157, {16'd49322, 16'd59544, 16'd8632, 16'd44996, 16'd28028, 16'd42371, 16'd54867, 16'd41174, 16'd42150, 16'd8612, 16'd12918, 16'd23695, 16'd42406, 16'd19263, 16'd17611, 16'd9567, 16'd48576, 16'd25998, 16'd40423, 16'd1751, 16'd16889, 16'd44734, 16'd65442, 16'd59856, 16'd12138, 16'd34622});
	test_expansion(128'h8ec6547f8e32f60e58058f2e201b303a, {16'd5421, 16'd766, 16'd18872, 16'd43307, 16'd60121, 16'd23339, 16'd25453, 16'd36268, 16'd23742, 16'd4552, 16'd20876, 16'd37148, 16'd65405, 16'd7982, 16'd575, 16'd61741, 16'd6164, 16'd7576, 16'd46769, 16'd37022, 16'd51362, 16'd23845, 16'd994, 16'd55443, 16'd40083, 16'd8564});
	test_expansion(128'h2878464a30c8865038b2905be686787b, {16'd50607, 16'd32224, 16'd11792, 16'd61092, 16'd42362, 16'd7578, 16'd25324, 16'd26571, 16'd33610, 16'd24956, 16'd32990, 16'd7739, 16'd51220, 16'd43617, 16'd65468, 16'd55925, 16'd53088, 16'd24375, 16'd22798, 16'd56428, 16'd34714, 16'd58301, 16'd36143, 16'd10741, 16'd16793, 16'd2866});
	test_expansion(128'hf60834a94af26b68e3457fba6a3533da, {16'd27526, 16'd22016, 16'd13621, 16'd42629, 16'd36426, 16'd18597, 16'd15980, 16'd225, 16'd39453, 16'd29974, 16'd37871, 16'd7323, 16'd30338, 16'd41490, 16'd62013, 16'd29012, 16'd43684, 16'd43528, 16'd22747, 16'd22837, 16'd14674, 16'd45347, 16'd15801, 16'd2679, 16'd54634, 16'd24642});
	test_expansion(128'h51294bc19490e85a392a6bd01e53f897, {16'd33378, 16'd44390, 16'd1386, 16'd46882, 16'd43818, 16'd43704, 16'd5477, 16'd1262, 16'd7583, 16'd34116, 16'd7231, 16'd29682, 16'd37527, 16'd58043, 16'd2686, 16'd60399, 16'd12569, 16'd8301, 16'd55035, 16'd53888, 16'd41548, 16'd29966, 16'd3575, 16'd64745, 16'd54140, 16'd61296});
	test_expansion(128'h25d0910c891421d318c77c784c34943d, {16'd37756, 16'd46208, 16'd46815, 16'd41420, 16'd17052, 16'd4195, 16'd63954, 16'd46516, 16'd40005, 16'd43560, 16'd7840, 16'd13595, 16'd32710, 16'd22539, 16'd35701, 16'd24910, 16'd14559, 16'd8170, 16'd51677, 16'd13011, 16'd46372, 16'd13451, 16'd35279, 16'd11006, 16'd21944, 16'd7945});
	test_expansion(128'h08e134883bf0f3d942827cddb884cf79, {16'd65457, 16'd52208, 16'd48242, 16'd52924, 16'd14896, 16'd37834, 16'd62407, 16'd14187, 16'd55955, 16'd23194, 16'd60716, 16'd35322, 16'd11372, 16'd14011, 16'd54309, 16'd26475, 16'd19479, 16'd18020, 16'd5843, 16'd23272, 16'd22164, 16'd9462, 16'd48542, 16'd47296, 16'd46527, 16'd62499});
	test_expansion(128'hfca3d1c65d198ddf532d6e18bb0b6e8d, {16'd55286, 16'd32768, 16'd63669, 16'd11340, 16'd41584, 16'd14363, 16'd2281, 16'd47921, 16'd7885, 16'd37879, 16'd34278, 16'd58498, 16'd59156, 16'd64028, 16'd44480, 16'd52640, 16'd10271, 16'd55952, 16'd62327, 16'd58299, 16'd11019, 16'd18423, 16'd37410, 16'd46317, 16'd29155, 16'd33818});
	test_expansion(128'h19945b72ea3e8068d839db04ee23e567, {16'd49487, 16'd39623, 16'd39373, 16'd38411, 16'd36895, 16'd24757, 16'd39810, 16'd59264, 16'd49189, 16'd56841, 16'd42858, 16'd8453, 16'd45699, 16'd31454, 16'd201, 16'd19795, 16'd34365, 16'd60091, 16'd46201, 16'd34539, 16'd38475, 16'd64205, 16'd6007, 16'd31321, 16'd51130, 16'd60249});
	test_expansion(128'ha7bfd4ff3c2183e5c01942097e112058, {16'd25272, 16'd20283, 16'd56781, 16'd64560, 16'd39981, 16'd44325, 16'd34209, 16'd59284, 16'd52937, 16'd15918, 16'd37635, 16'd5113, 16'd33970, 16'd27551, 16'd25159, 16'd22623, 16'd13693, 16'd1124, 16'd27953, 16'd50238, 16'd38297, 16'd55671, 16'd43824, 16'd7211, 16'd22331, 16'd44379});
	test_expansion(128'hf2ec3302a86c9d73846ebb805915a960, {16'd58261, 16'd64725, 16'd21041, 16'd42057, 16'd17772, 16'd21966, 16'd12692, 16'd7115, 16'd25045, 16'd16035, 16'd61219, 16'd13809, 16'd52491, 16'd22674, 16'd54479, 16'd22182, 16'd6931, 16'd5656, 16'd40482, 16'd57260, 16'd39775, 16'd42291, 16'd29710, 16'd29167, 16'd36747, 16'd59318});
	test_expansion(128'hb9303a3706fb8100349e81148bbed221, {16'd8664, 16'd26795, 16'd48857, 16'd56561, 16'd47378, 16'd56772, 16'd10432, 16'd42251, 16'd10022, 16'd55599, 16'd10592, 16'd23702, 16'd24117, 16'd53884, 16'd35932, 16'd56665, 16'd43558, 16'd7872, 16'd9128, 16'd6694, 16'd25272, 16'd30683, 16'd59108, 16'd16335, 16'd36908, 16'd8263});
	test_expansion(128'h036d01d582c07a2b718ca0c2dce36335, {16'd63354, 16'd30899, 16'd35787, 16'd50552, 16'd13166, 16'd21967, 16'd21507, 16'd7494, 16'd27146, 16'd50895, 16'd61363, 16'd34856, 16'd32418, 16'd60455, 16'd31147, 16'd18032, 16'd4632, 16'd44303, 16'd1796, 16'd15547, 16'd634, 16'd3260, 16'd14071, 16'd15173, 16'd7616, 16'd44497});
	test_expansion(128'h0ad502d4b4483b808dcbadb39630bbc8, {16'd51542, 16'd32177, 16'd33377, 16'd45525, 16'd8737, 16'd47283, 16'd7503, 16'd61835, 16'd46733, 16'd18183, 16'd56486, 16'd59068, 16'd15735, 16'd20684, 16'd54518, 16'd54771, 16'd9048, 16'd11228, 16'd24015, 16'd56079, 16'd55025, 16'd8919, 16'd37820, 16'd18798, 16'd46126, 16'd16999});
	test_expansion(128'h8e027ce1af3bfcc88171b4568a9945d5, {16'd56861, 16'd43474, 16'd51832, 16'd42048, 16'd13550, 16'd6980, 16'd14040, 16'd15035, 16'd47424, 16'd44129, 16'd32932, 16'd2151, 16'd33144, 16'd57199, 16'd62003, 16'd47607, 16'd7110, 16'd52386, 16'd54247, 16'd56091, 16'd53821, 16'd27073, 16'd29079, 16'd19035, 16'd33589, 16'd3812});
	test_expansion(128'hba11952fb2bcae644b77a5c12e2454de, {16'd33654, 16'd59747, 16'd57192, 16'd36089, 16'd55113, 16'd50767, 16'd35317, 16'd36768, 16'd3721, 16'd21059, 16'd61600, 16'd62831, 16'd55363, 16'd26443, 16'd35976, 16'd15247, 16'd36352, 16'd23119, 16'd9027, 16'd2570, 16'd44212, 16'd41174, 16'd11528, 16'd30206, 16'd43812, 16'd22924});
	test_expansion(128'h9e66423dcd44e8280248f3ba98a73424, {16'd21107, 16'd56083, 16'd56144, 16'd4374, 16'd11109, 16'd16778, 16'd14723, 16'd843, 16'd60595, 16'd45507, 16'd56853, 16'd41599, 16'd15268, 16'd26772, 16'd16426, 16'd19379, 16'd51023, 16'd36191, 16'd18299, 16'd31833, 16'd21115, 16'd48864, 16'd12815, 16'd29343, 16'd34883, 16'd48811});
	test_expansion(128'hc9a90730454c8ce407804c5b1c92df34, {16'd11022, 16'd14413, 16'd59417, 16'd39951, 16'd46606, 16'd4153, 16'd13370, 16'd17812, 16'd53420, 16'd39860, 16'd39989, 16'd52693, 16'd46930, 16'd10407, 16'd51992, 16'd21581, 16'd12894, 16'd44660, 16'd60577, 16'd34400, 16'd28671, 16'd64271, 16'd20413, 16'd25426, 16'd44793, 16'd15615});
	test_expansion(128'h3f6220eb20260b20895d83b11749381a, {16'd28394, 16'd58547, 16'd14397, 16'd63384, 16'd15021, 16'd12457, 16'd55132, 16'd56640, 16'd63090, 16'd19706, 16'd51357, 16'd47639, 16'd56743, 16'd18225, 16'd62665, 16'd16677, 16'd31907, 16'd27891, 16'd31802, 16'd33320, 16'd17639, 16'd57375, 16'd64004, 16'd42047, 16'd11583, 16'd59696});
	test_expansion(128'hd3c2a63c8a314c505c562e64ba6aa11c, {16'd48273, 16'd14491, 16'd12074, 16'd35524, 16'd29735, 16'd22429, 16'd13922, 16'd55234, 16'd37475, 16'd24689, 16'd48203, 16'd54909, 16'd64168, 16'd60914, 16'd18978, 16'd39769, 16'd3873, 16'd57592, 16'd17796, 16'd9530, 16'd53059, 16'd26206, 16'd1729, 16'd57103, 16'd14282, 16'd3395});
	test_expansion(128'ha7b935e462f577c0163c923f45a39a16, {16'd54888, 16'd29707, 16'd44028, 16'd20014, 16'd55570, 16'd30311, 16'd41728, 16'd28964, 16'd2851, 16'd38535, 16'd58136, 16'd34853, 16'd60008, 16'd21416, 16'd30037, 16'd32758, 16'd2725, 16'd10724, 16'd63458, 16'd20726, 16'd6731, 16'd26482, 16'd33872, 16'd14112, 16'd9063, 16'd51020});
	test_expansion(128'h5c3dda6a85fcb7e40d293223d66fc12e, {16'd4386, 16'd21285, 16'd51469, 16'd18757, 16'd20151, 16'd9809, 16'd24993, 16'd58444, 16'd30400, 16'd4975, 16'd3400, 16'd16083, 16'd48316, 16'd58012, 16'd44604, 16'd37784, 16'd6224, 16'd62269, 16'd49497, 16'd57832, 16'd5932, 16'd43052, 16'd14638, 16'd19363, 16'd12222, 16'd36714});
	test_expansion(128'h5cb9e2474ec708072734bf8ea1630a9d, {16'd59570, 16'd25734, 16'd17240, 16'd18876, 16'd20651, 16'd56234, 16'd62437, 16'd3188, 16'd40446, 16'd36743, 16'd10120, 16'd40893, 16'd62845, 16'd53103, 16'd12828, 16'd7703, 16'd47601, 16'd51690, 16'd58051, 16'd52121, 16'd49197, 16'd41338, 16'd4197, 16'd29277, 16'd17823, 16'd21897});
	test_expansion(128'h0604fea12ad07f5f490d8d015f408d5d, {16'd96, 16'd19016, 16'd52603, 16'd41590, 16'd34933, 16'd56395, 16'd30099, 16'd58750, 16'd47131, 16'd37668, 16'd35334, 16'd31676, 16'd44312, 16'd32347, 16'd25362, 16'd28838, 16'd46579, 16'd17045, 16'd50246, 16'd42463, 16'd63353, 16'd47684, 16'd55043, 16'd10410, 16'd44881, 16'd26239});
	test_expansion(128'h566551f84277710912b52896fd3a3dc2, {16'd50349, 16'd12943, 16'd61019, 16'd43643, 16'd36284, 16'd44342, 16'd27488, 16'd21081, 16'd48751, 16'd34109, 16'd11010, 16'd38054, 16'd58718, 16'd56536, 16'd39267, 16'd59860, 16'd46986, 16'd1932, 16'd58148, 16'd42608, 16'd57239, 16'd46234, 16'd32734, 16'd23295, 16'd33998, 16'd52091});
	test_expansion(128'hc2721218163298ddd726ad16580e24f5, {16'd34704, 16'd52951, 16'd285, 16'd2207, 16'd49969, 16'd18993, 16'd55652, 16'd26566, 16'd15715, 16'd14444, 16'd36956, 16'd34305, 16'd28508, 16'd38839, 16'd55342, 16'd32887, 16'd30086, 16'd56648, 16'd13814, 16'd55648, 16'd18778, 16'd51786, 16'd29417, 16'd46538, 16'd11028, 16'd25681});
	test_expansion(128'h4f679f71fbf309445053fd320184c4f6, {16'd64927, 16'd5390, 16'd50560, 16'd33549, 16'd11076, 16'd9829, 16'd6298, 16'd20673, 16'd49728, 16'd58582, 16'd30137, 16'd11194, 16'd26278, 16'd44543, 16'd31399, 16'd24821, 16'd1332, 16'd55711, 16'd54851, 16'd15954, 16'd20388, 16'd57147, 16'd64176, 16'd1162, 16'd64463, 16'd48702});
	test_expansion(128'h10a71f64dc4772a5b71a70618fea8002, {16'd54360, 16'd61224, 16'd39103, 16'd18078, 16'd31909, 16'd42305, 16'd24437, 16'd32959, 16'd59997, 16'd3891, 16'd20432, 16'd1119, 16'd60371, 16'd58511, 16'd41608, 16'd20986, 16'd63563, 16'd7832, 16'd33635, 16'd9686, 16'd60865, 16'd53982, 16'd21458, 16'd30603, 16'd14583, 16'd839});
	test_expansion(128'h52a1a47fca592f21645ac8e346915584, {16'd18770, 16'd34819, 16'd13264, 16'd38304, 16'd13936, 16'd5325, 16'd28128, 16'd25810, 16'd8740, 16'd19934, 16'd53251, 16'd49719, 16'd60386, 16'd33022, 16'd16385, 16'd55549, 16'd15883, 16'd48201, 16'd5180, 16'd4500, 16'd36515, 16'd39016, 16'd29424, 16'd3155, 16'd20584, 16'd56653});
	test_expansion(128'h236e5b9bc214287cd97bc7b335e311e4, {16'd21894, 16'd8793, 16'd31978, 16'd15359, 16'd44677, 16'd15692, 16'd27916, 16'd26549, 16'd33248, 16'd32894, 16'd58597, 16'd34961, 16'd62803, 16'd15413, 16'd60341, 16'd36023, 16'd37467, 16'd49254, 16'd51852, 16'd63602, 16'd28129, 16'd2999, 16'd54368, 16'd10824, 16'd23221, 16'd35231});
	test_expansion(128'h4353293612056bbf279131b2f27838a2, {16'd14675, 16'd25639, 16'd45429, 16'd34718, 16'd51963, 16'd37067, 16'd63885, 16'd39821, 16'd34758, 16'd41777, 16'd15988, 16'd56251, 16'd413, 16'd19452, 16'd2425, 16'd64695, 16'd16044, 16'd5215, 16'd34573, 16'd410, 16'd55365, 16'd50226, 16'd54095, 16'd4067, 16'd26405, 16'd30640});
	test_expansion(128'h87781242143928f71497a7bd95d59437, {16'd56717, 16'd7129, 16'd45277, 16'd34152, 16'd19368, 16'd40474, 16'd56830, 16'd38201, 16'd54223, 16'd42318, 16'd32724, 16'd46733, 16'd53571, 16'd64505, 16'd15048, 16'd4748, 16'd55256, 16'd16543, 16'd52626, 16'd64123, 16'd60199, 16'd29150, 16'd38157, 16'd5487, 16'd62175, 16'd22992});
	test_expansion(128'h3f55cecd6b84b87bab2e753f327b0644, {16'd16358, 16'd64420, 16'd36464, 16'd5778, 16'd57334, 16'd50674, 16'd22456, 16'd59103, 16'd3151, 16'd62049, 16'd24307, 16'd64010, 16'd8634, 16'd50898, 16'd46847, 16'd20144, 16'd11917, 16'd3601, 16'd62358, 16'd12584, 16'd25786, 16'd62454, 16'd30057, 16'd54064, 16'd45466, 16'd10130});
	test_expansion(128'h7d8e2dc8f140dd1faa744636b6223737, {16'd44902, 16'd23771, 16'd51864, 16'd36021, 16'd26281, 16'd35845, 16'd24453, 16'd57959, 16'd60716, 16'd33367, 16'd28719, 16'd11656, 16'd48893, 16'd27205, 16'd14938, 16'd27279, 16'd43797, 16'd39871, 16'd16513, 16'd8014, 16'd64566, 16'd42869, 16'd28600, 16'd25747, 16'd17630, 16'd39122});
	test_expansion(128'hb1b81f0fbc34c45a4f71ea1321a84f36, {16'd17658, 16'd53498, 16'd13714, 16'd21630, 16'd33684, 16'd21240, 16'd7063, 16'd12780, 16'd19284, 16'd50392, 16'd55729, 16'd46730, 16'd9187, 16'd54359, 16'd22103, 16'd17102, 16'd9212, 16'd7705, 16'd33608, 16'd49794, 16'd31884, 16'd37891, 16'd11180, 16'd34463, 16'd23213, 16'd61631});
	test_expansion(128'h85983c147d1e823cd676c2791c435ca7, {16'd27480, 16'd64648, 16'd42973, 16'd64056, 16'd26483, 16'd16652, 16'd45518, 16'd48092, 16'd16453, 16'd48674, 16'd44647, 16'd43976, 16'd38292, 16'd6211, 16'd51259, 16'd21409, 16'd12565, 16'd61563, 16'd10866, 16'd36598, 16'd12840, 16'd9348, 16'd60516, 16'd64935, 16'd53408, 16'd11567});
	test_expansion(128'hbba10044c039af31a96ba5009f596d0e, {16'd22884, 16'd24828, 16'd28418, 16'd10671, 16'd27405, 16'd42166, 16'd42790, 16'd26379, 16'd39000, 16'd37117, 16'd4633, 16'd8881, 16'd12193, 16'd46566, 16'd64189, 16'd16421, 16'd17353, 16'd51798, 16'd6620, 16'd54890, 16'd3378, 16'd2238, 16'd5668, 16'd30555, 16'd25587, 16'd33121});
	test_expansion(128'h120ad3f82e6498a40a22327f32635519, {16'd35323, 16'd51453, 16'd45366, 16'd19874, 16'd5371, 16'd25389, 16'd6475, 16'd56716, 16'd25593, 16'd18943, 16'd16584, 16'd7123, 16'd49928, 16'd220, 16'd35854, 16'd59746, 16'd631, 16'd9832, 16'd7289, 16'd14858, 16'd54717, 16'd28420, 16'd36691, 16'd36566, 16'd10178, 16'd36334});
	test_expansion(128'h4ee00d5f703b5610e47236028256f82e, {16'd8229, 16'd9586, 16'd3171, 16'd64697, 16'd4673, 16'd7212, 16'd28596, 16'd33717, 16'd45336, 16'd17938, 16'd41039, 16'd1872, 16'd7590, 16'd44071, 16'd53250, 16'd31917, 16'd61776, 16'd27929, 16'd32178, 16'd17564, 16'd28435, 16'd44706, 16'd45635, 16'd21683, 16'd25260, 16'd55333});
	test_expansion(128'h8582e9019309f5da29911de0cb514345, {16'd19618, 16'd60599, 16'd17604, 16'd9668, 16'd38852, 16'd20276, 16'd25417, 16'd32113, 16'd11814, 16'd46039, 16'd35015, 16'd58155, 16'd22914, 16'd51155, 16'd29446, 16'd33428, 16'd29510, 16'd8792, 16'd24763, 16'd38251, 16'd28221, 16'd21169, 16'd63454, 16'd55231, 16'd5539, 16'd45164});
	test_expansion(128'h6775efa9b700ec45638b0448f7054a70, {16'd64537, 16'd1402, 16'd49129, 16'd47132, 16'd9178, 16'd55749, 16'd15024, 16'd11039, 16'd9829, 16'd15046, 16'd23370, 16'd37717, 16'd19348, 16'd47108, 16'd57522, 16'd24901, 16'd51488, 16'd2742, 16'd25121, 16'd17949, 16'd45995, 16'd30318, 16'd45191, 16'd10875, 16'd28986, 16'd21168});
	test_expansion(128'h597108464e3a58497c0277c42fce2648, {16'd63370, 16'd35741, 16'd117, 16'd2500, 16'd39799, 16'd53005, 16'd25558, 16'd19947, 16'd52982, 16'd56846, 16'd39483, 16'd2523, 16'd56463, 16'd31464, 16'd33593, 16'd54181, 16'd46294, 16'd12974, 16'd8596, 16'd51198, 16'd54021, 16'd56184, 16'd5906, 16'd59532, 16'd40167, 16'd58700});
	test_expansion(128'hfe2619efbc994322762dffdde8803a76, {16'd21539, 16'd64480, 16'd62483, 16'd38257, 16'd9447, 16'd14644, 16'd4999, 16'd27617, 16'd410, 16'd2201, 16'd63566, 16'd5428, 16'd26546, 16'd20197, 16'd50344, 16'd39242, 16'd23991, 16'd54007, 16'd64084, 16'd54520, 16'd53305, 16'd31495, 16'd14392, 16'd53543, 16'd53541, 16'd39037});
	test_expansion(128'hf281073e52e663be497f7171223d0c82, {16'd38892, 16'd35754, 16'd46302, 16'd17899, 16'd62443, 16'd3289, 16'd55135, 16'd25585, 16'd35448, 16'd39446, 16'd24659, 16'd47919, 16'd58047, 16'd16475, 16'd8299, 16'd58743, 16'd33371, 16'd63267, 16'd1679, 16'd6017, 16'd27189, 16'd27146, 16'd53650, 16'd33573, 16'd60523, 16'd31633});
	test_expansion(128'hb32b8224a3025a9a5edddf7f8fe2504a, {16'd55310, 16'd36580, 16'd52650, 16'd45523, 16'd32971, 16'd63333, 16'd50119, 16'd43148, 16'd17572, 16'd44695, 16'd6559, 16'd14802, 16'd20843, 16'd60731, 16'd45035, 16'd38105, 16'd41005, 16'd60559, 16'd12360, 16'd44713, 16'd33478, 16'd23286, 16'd29900, 16'd28989, 16'd34881, 16'd13860});
	test_expansion(128'h199a2c50472a6b440ef6e924ca795071, {16'd46249, 16'd29350, 16'd41691, 16'd50080, 16'd13086, 16'd20197, 16'd4666, 16'd34152, 16'd40704, 16'd44623, 16'd17588, 16'd49534, 16'd2601, 16'd12836, 16'd23928, 16'd29433, 16'd6408, 16'd32850, 16'd39498, 16'd49058, 16'd37603, 16'd61886, 16'd11871, 16'd43493, 16'd57847, 16'd48296});
	test_expansion(128'h19cc04d7b2a790eb84e22f3fdb2e24d4, {16'd19198, 16'd39543, 16'd44891, 16'd5663, 16'd599, 16'd40155, 16'd7637, 16'd46070, 16'd57152, 16'd2260, 16'd42662, 16'd41830, 16'd58736, 16'd46983, 16'd46109, 16'd21565, 16'd16043, 16'd15312, 16'd17568, 16'd32075, 16'd2359, 16'd13182, 16'd62384, 16'd3618, 16'd5405, 16'd39114});
	test_expansion(128'h2f735ff5c83d225954c559996231c426, {16'd20031, 16'd59672, 16'd53479, 16'd39075, 16'd22426, 16'd40764, 16'd61521, 16'd6901, 16'd53333, 16'd22383, 16'd21313, 16'd15612, 16'd3, 16'd24031, 16'd44969, 16'd39108, 16'd12920, 16'd10446, 16'd57221, 16'd32177, 16'd7895, 16'd26068, 16'd56951, 16'd3657, 16'd47417, 16'd13320});
	test_expansion(128'h063a85ba1c313a7f994e64ae0ee498db, {16'd56844, 16'd49662, 16'd39133, 16'd40755, 16'd63820, 16'd60567, 16'd931, 16'd44247, 16'd57768, 16'd27093, 16'd50071, 16'd36856, 16'd32838, 16'd21598, 16'd7931, 16'd6638, 16'd58429, 16'd48714, 16'd27674, 16'd24353, 16'd29134, 16'd40325, 16'd47475, 16'd42149, 16'd3249, 16'd54916});
	test_expansion(128'hf4e568bda4a55214af5daf50dc2aaadd, {16'd28772, 16'd49757, 16'd43099, 16'd6376, 16'd28060, 16'd45292, 16'd36679, 16'd6906, 16'd32387, 16'd6361, 16'd39740, 16'd8286, 16'd47985, 16'd30836, 16'd33571, 16'd6664, 16'd54117, 16'd30926, 16'd11609, 16'd27082, 16'd4939, 16'd21249, 16'd15259, 16'd58809, 16'd5658, 16'd1279});
	test_expansion(128'h41e8048589c5b3a37a7e91ddc34d9010, {16'd58097, 16'd35508, 16'd9782, 16'd23941, 16'd4464, 16'd28052, 16'd42472, 16'd56742, 16'd17548, 16'd39484, 16'd26750, 16'd59122, 16'd4278, 16'd28334, 16'd22851, 16'd16096, 16'd62373, 16'd26075, 16'd15190, 16'd61824, 16'd64956, 16'd37057, 16'd18896, 16'd19525, 16'd11410, 16'd24102});
	test_expansion(128'h8fabfd76c0570faa39da106d0b12b4e4, {16'd28211, 16'd48883, 16'd56089, 16'd65113, 16'd59313, 16'd10638, 16'd23917, 16'd13675, 16'd16953, 16'd60489, 16'd54010, 16'd14216, 16'd18367, 16'd29782, 16'd29255, 16'd21149, 16'd15677, 16'd15626, 16'd33845, 16'd19049, 16'd4087, 16'd5667, 16'd15805, 16'd29579, 16'd30461, 16'd10638});
	test_expansion(128'h77b88228cc0e7be8485bf04f7b29ff1e, {16'd42379, 16'd15150, 16'd60668, 16'd34099, 16'd14523, 16'd32616, 16'd8293, 16'd11813, 16'd31560, 16'd13488, 16'd8872, 16'd34466, 16'd51828, 16'd2192, 16'd55943, 16'd24454, 16'd39369, 16'd30972, 16'd12334, 16'd36110, 16'd17454, 16'd35978, 16'd20732, 16'd45016, 16'd41856, 16'd51505});
	test_expansion(128'h96ff97768ce41fe6d7e3e0c23e7f4b73, {16'd51283, 16'd29811, 16'd8351, 16'd47359, 16'd61427, 16'd53347, 16'd47459, 16'd18572, 16'd35762, 16'd62315, 16'd60142, 16'd34345, 16'd34162, 16'd61323, 16'd49260, 16'd45286, 16'd10724, 16'd48741, 16'd57900, 16'd60950, 16'd54662, 16'd32146, 16'd31492, 16'd43745, 16'd31551, 16'd55118});
	test_expansion(128'h924dfdcada9079021a484e4619b65f96, {16'd23553, 16'd8160, 16'd52026, 16'd7250, 16'd60289, 16'd52255, 16'd19747, 16'd63819, 16'd37429, 16'd41835, 16'd40936, 16'd2220, 16'd41658, 16'd50359, 16'd7429, 16'd64802, 16'd49334, 16'd17658, 16'd64352, 16'd45013, 16'd50782, 16'd10458, 16'd45267, 16'd22132, 16'd35251, 16'd29454});
	test_expansion(128'ha6da7548bd55bd2cd6aad6968d869dc2, {16'd54489, 16'd54503, 16'd49544, 16'd46772, 16'd1310, 16'd21865, 16'd30573, 16'd3393, 16'd64179, 16'd36431, 16'd20919, 16'd6093, 16'd10958, 16'd51180, 16'd54510, 16'd37023, 16'd5696, 16'd27274, 16'd43487, 16'd47583, 16'd16185, 16'd16931, 16'd1430, 16'd49575, 16'd62389, 16'd48605});
	test_expansion(128'he4934ee9ab3b558567d9279e2beeccbc, {16'd54224, 16'd7857, 16'd42461, 16'd959, 16'd9047, 16'd1966, 16'd61044, 16'd60619, 16'd51200, 16'd43671, 16'd3092, 16'd58620, 16'd58770, 16'd62116, 16'd46585, 16'd9125, 16'd55876, 16'd17643, 16'd14183, 16'd25258, 16'd57738, 16'd25282, 16'd15547, 16'd1593, 16'd39753, 16'd51961});
	test_expansion(128'h14268d04aac6d5619c9d48b07e483b23, {16'd41911, 16'd18637, 16'd50467, 16'd62710, 16'd38054, 16'd1109, 16'd44049, 16'd893, 16'd48732, 16'd21384, 16'd27836, 16'd52470, 16'd24271, 16'd47869, 16'd18568, 16'd37369, 16'd58509, 16'd58825, 16'd29990, 16'd33550, 16'd64409, 16'd9814, 16'd28852, 16'd11176, 16'd11747, 16'd48969});
	test_expansion(128'h5a481ffb10bf452bcbe8eac98f8f7b8a, {16'd31233, 16'd10264, 16'd40228, 16'd28038, 16'd38575, 16'd20981, 16'd21845, 16'd62044, 16'd33332, 16'd24450, 16'd60474, 16'd47256, 16'd42265, 16'd45155, 16'd9428, 16'd23866, 16'd64888, 16'd27688, 16'd57626, 16'd49767, 16'd45176, 16'd51697, 16'd59251, 16'd52100, 16'd61684, 16'd20948});
	test_expansion(128'hdfdc886fd864c3648c003b09fc3dd2fe, {16'd41621, 16'd45226, 16'd43864, 16'd21256, 16'd34372, 16'd4291, 16'd35355, 16'd64102, 16'd28788, 16'd12506, 16'd8168, 16'd51692, 16'd41879, 16'd37220, 16'd27056, 16'd7738, 16'd9276, 16'd62376, 16'd30326, 16'd64717, 16'd37656, 16'd58914, 16'd55685, 16'd22752, 16'd56510, 16'd16971});
	test_expansion(128'h04eca3893c56c09cafa83e3aa6a42e0c, {16'd33546, 16'd34278, 16'd56038, 16'd50804, 16'd11296, 16'd58496, 16'd6998, 16'd19037, 16'd61930, 16'd24594, 16'd39636, 16'd9499, 16'd2049, 16'd52942, 16'd19619, 16'd36326, 16'd40968, 16'd54847, 16'd1628, 16'd44254, 16'd24416, 16'd36633, 16'd21709, 16'd14271, 16'd15513, 16'd18592});
	test_expansion(128'h07ffcf723ae12c0e678b6f17153f3fe5, {16'd29984, 16'd19433, 16'd37931, 16'd41222, 16'd15064, 16'd15967, 16'd63636, 16'd5041, 16'd3626, 16'd15295, 16'd37957, 16'd55782, 16'd33452, 16'd53765, 16'd45302, 16'd21220, 16'd30828, 16'd59564, 16'd42065, 16'd26896, 16'd62481, 16'd18300, 16'd12708, 16'd24624, 16'd47908, 16'd50718});
	test_expansion(128'hbcf068b4239ce60f89f8c4b368964f65, {16'd49728, 16'd14686, 16'd31371, 16'd21549, 16'd1783, 16'd62532, 16'd39411, 16'd53277, 16'd45544, 16'd48468, 16'd8422, 16'd55110, 16'd21884, 16'd1360, 16'd44078, 16'd30941, 16'd14635, 16'd3563, 16'd9170, 16'd62968, 16'd34320, 16'd44908, 16'd41975, 16'd26523, 16'd44148, 16'd24755});
	test_expansion(128'h51810f14acea8fe1ca9cb8368a4f75c9, {16'd32677, 16'd45706, 16'd13271, 16'd46244, 16'd5083, 16'd3321, 16'd34651, 16'd37838, 16'd30693, 16'd64374, 16'd42378, 16'd32197, 16'd4840, 16'd773, 16'd30945, 16'd1727, 16'd30223, 16'd56252, 16'd26974, 16'd65323, 16'd51127, 16'd34915, 16'd11402, 16'd65109, 16'd37290, 16'd11935});
	test_expansion(128'h3eec45489025e045786bdbb0dd15c12d, {16'd9740, 16'd4932, 16'd21981, 16'd39261, 16'd43991, 16'd35250, 16'd46739, 16'd27971, 16'd24475, 16'd25315, 16'd62897, 16'd26149, 16'd974, 16'd12881, 16'd60404, 16'd3228, 16'd19810, 16'd34883, 16'd28653, 16'd24130, 16'd44813, 16'd57808, 16'd2686, 16'd513, 16'd48885, 16'd3136});
	test_expansion(128'hd14a06412b38e3e948b645b52052f7e7, {16'd8123, 16'd21439, 16'd38344, 16'd56447, 16'd632, 16'd22266, 16'd2551, 16'd30616, 16'd17092, 16'd33133, 16'd17823, 16'd51579, 16'd20916, 16'd27830, 16'd34409, 16'd33359, 16'd49278, 16'd49994, 16'd35879, 16'd12004, 16'd53596, 16'd55026, 16'd40786, 16'd61141, 16'd37076, 16'd32560});
	test_expansion(128'h2ed85159772734e68a0b7720e7348abc, {16'd12542, 16'd11609, 16'd31762, 16'd60722, 16'd60544, 16'd22536, 16'd48472, 16'd45431, 16'd13246, 16'd25986, 16'd40385, 16'd36363, 16'd18876, 16'd28791, 16'd29044, 16'd63810, 16'd51982, 16'd3839, 16'd1794, 16'd25280, 16'd47383, 16'd54103, 16'd45134, 16'd50009, 16'd33625, 16'd39603});
	test_expansion(128'h6fc449bb2af4299b5b29b5cf38a07981, {16'd25626, 16'd51774, 16'd2929, 16'd41642, 16'd34692, 16'd42291, 16'd42051, 16'd5299, 16'd26876, 16'd4467, 16'd37653, 16'd13820, 16'd20408, 16'd54531, 16'd29681, 16'd19910, 16'd58428, 16'd55744, 16'd38199, 16'd43281, 16'd44910, 16'd46864, 16'd10407, 16'd26190, 16'd29931, 16'd58740});
	test_expansion(128'h270fed757c275869dbeba8c88634c8ba, {16'd61569, 16'd12267, 16'd54589, 16'd48373, 16'd29258, 16'd20030, 16'd51369, 16'd56028, 16'd38301, 16'd54083, 16'd17693, 16'd21801, 16'd60026, 16'd61512, 16'd42017, 16'd26928, 16'd33250, 16'd10732, 16'd3762, 16'd53255, 16'd38698, 16'd47251, 16'd29225, 16'd49645, 16'd19526, 16'd64856});
	test_expansion(128'hae258c68e16a3e9319be1535c3ef65b0, {16'd65231, 16'd55040, 16'd51143, 16'd23842, 16'd55713, 16'd8882, 16'd5178, 16'd65502, 16'd54882, 16'd31614, 16'd54822, 16'd59139, 16'd34167, 16'd41488, 16'd24462, 16'd11681, 16'd28847, 16'd52681, 16'd27347, 16'd44082, 16'd30441, 16'd7641, 16'd53718, 16'd3991, 16'd53676, 16'd32351});
	test_expansion(128'h86ee7282b1cc8ad33ba696b262d9c527, {16'd42129, 16'd48992, 16'd8383, 16'd14435, 16'd12527, 16'd33523, 16'd3184, 16'd54184, 16'd24099, 16'd27497, 16'd29401, 16'd52685, 16'd29865, 16'd40698, 16'd11556, 16'd31477, 16'd43454, 16'd39794, 16'd46497, 16'd36214, 16'd64545, 16'd7825, 16'd49708, 16'd54511, 16'd56605, 16'd30499});
	test_expansion(128'he6aae087fc128b06ade48ea2f004e6bd, {16'd29941, 16'd31645, 16'd37903, 16'd62998, 16'd16401, 16'd60282, 16'd47903, 16'd53164, 16'd34540, 16'd40912, 16'd21488, 16'd13928, 16'd38443, 16'd48677, 16'd20646, 16'd15256, 16'd31500, 16'd5461, 16'd56921, 16'd15842, 16'd53889, 16'd35795, 16'd22237, 16'd54126, 16'd26219, 16'd33367});
	test_expansion(128'hec6ce859d6753bc91abdbb0fe1c2c09e, {16'd53907, 16'd47981, 16'd8985, 16'd25101, 16'd31343, 16'd32655, 16'd58337, 16'd1515, 16'd39426, 16'd12893, 16'd44804, 16'd7387, 16'd10428, 16'd55262, 16'd30411, 16'd58459, 16'd27294, 16'd56719, 16'd4306, 16'd27243, 16'd32143, 16'd23831, 16'd9920, 16'd40771, 16'd13129, 16'd20216});
	test_expansion(128'h57637982d9c0c167de4b047582108e49, {16'd9419, 16'd26193, 16'd51348, 16'd39585, 16'd33763, 16'd16560, 16'd25620, 16'd51163, 16'd43643, 16'd52712, 16'd1567, 16'd59403, 16'd857, 16'd14817, 16'd7018, 16'd6596, 16'd44721, 16'd12750, 16'd62183, 16'd35876, 16'd62052, 16'd12165, 16'd60992, 16'd45106, 16'd57526, 16'd45450});
	test_expansion(128'h0fc21481962a72107e9abca98831e7b2, {16'd17508, 16'd45479, 16'd5328, 16'd35281, 16'd45297, 16'd7703, 16'd37942, 16'd64476, 16'd63576, 16'd30003, 16'd9848, 16'd28034, 16'd53755, 16'd27175, 16'd8572, 16'd44562, 16'd57798, 16'd57944, 16'd46935, 16'd30841, 16'd44461, 16'd30222, 16'd59147, 16'd42470, 16'd60377, 16'd54451});
	test_expansion(128'hc469154edd1bfba1fbe9285e39c2b580, {16'd17288, 16'd18317, 16'd65092, 16'd58943, 16'd31095, 16'd57166, 16'd41779, 16'd25588, 16'd15354, 16'd18690, 16'd3628, 16'd59651, 16'd50933, 16'd27569, 16'd32004, 16'd8261, 16'd42901, 16'd58039, 16'd52787, 16'd64167, 16'd14990, 16'd32158, 16'd618, 16'd34101, 16'd31504, 16'd3534});
	test_expansion(128'h3628c4728031594df06e72f65fe5c97d, {16'd30802, 16'd56565, 16'd8012, 16'd18450, 16'd3504, 16'd18016, 16'd4040, 16'd7601, 16'd20940, 16'd52344, 16'd56880, 16'd825, 16'd36057, 16'd30741, 16'd64648, 16'd31220, 16'd55546, 16'd38771, 16'd8507, 16'd30556, 16'd32362, 16'd22087, 16'd14371, 16'd24980, 16'd8509, 16'd20383});
	test_expansion(128'headb5ac679dbd693b7b61a8eebb3baa0, {16'd28153, 16'd57066, 16'd65300, 16'd30229, 16'd30721, 16'd60579, 16'd30287, 16'd44548, 16'd28513, 16'd55853, 16'd32536, 16'd40103, 16'd30944, 16'd54245, 16'd34297, 16'd19854, 16'd51063, 16'd40494, 16'd41923, 16'd44490, 16'd62416, 16'd7918, 16'd55299, 16'd37226, 16'd16723, 16'd62296});
	test_expansion(128'hdda110a16102b5801afe80528083b20f, {16'd28721, 16'd9591, 16'd42713, 16'd50547, 16'd32665, 16'd40082, 16'd31849, 16'd56191, 16'd48898, 16'd19308, 16'd33600, 16'd44746, 16'd22460, 16'd43343, 16'd49805, 16'd13269, 16'd13600, 16'd38698, 16'd37892, 16'd19592, 16'd11944, 16'd56154, 16'd44282, 16'd2312, 16'd54010, 16'd6812});
	test_expansion(128'h8d1c64a36306b7d330f214269a7216da, {16'd39950, 16'd42160, 16'd33170, 16'd14437, 16'd39863, 16'd242, 16'd63684, 16'd45594, 16'd10761, 16'd47420, 16'd51352, 16'd45729, 16'd58338, 16'd12265, 16'd40902, 16'd12653, 16'd47346, 16'd11433, 16'd49822, 16'd3096, 16'd16588, 16'd13049, 16'd15800, 16'd28122, 16'd30136, 16'd9530});
	test_expansion(128'h2cdecbd55f9199e5845cc7a14e50d880, {16'd25149, 16'd58666, 16'd39847, 16'd42290, 16'd14095, 16'd49229, 16'd28201, 16'd33636, 16'd12187, 16'd46721, 16'd58340, 16'd20555, 16'd60730, 16'd47011, 16'd18282, 16'd57377, 16'd16537, 16'd25769, 16'd60710, 16'd25724, 16'd12870, 16'd4215, 16'd37950, 16'd44340, 16'd58041, 16'd5257});
	test_expansion(128'h4e9fc8ea4eb8c835eae68f21a022ef72, {16'd39306, 16'd55313, 16'd59157, 16'd33349, 16'd61393, 16'd23897, 16'd48900, 16'd60565, 16'd45473, 16'd26519, 16'd6901, 16'd49838, 16'd63620, 16'd62873, 16'd13980, 16'd10621, 16'd37811, 16'd63318, 16'd9994, 16'd7798, 16'd59432, 16'd12003, 16'd17572, 16'd56308, 16'd47325, 16'd30144});
	test_expansion(128'h7c9c1dbf63e3f500b2d9c3cd974c5933, {16'd18623, 16'd54360, 16'd7069, 16'd49176, 16'd62098, 16'd52570, 16'd48342, 16'd36744, 16'd47216, 16'd1562, 16'd24422, 16'd21360, 16'd63897, 16'd12451, 16'd1613, 16'd21260, 16'd8420, 16'd3736, 16'd46115, 16'd21289, 16'd63335, 16'd65286, 16'd64305, 16'd46874, 16'd1745, 16'd44935});
	test_expansion(128'hb80da4fcb35ba767f8775925b885159e, {16'd42743, 16'd9505, 16'd13454, 16'd46741, 16'd29060, 16'd6140, 16'd28387, 16'd55127, 16'd61764, 16'd25632, 16'd4096, 16'd8353, 16'd12602, 16'd40875, 16'd22837, 16'd22020, 16'd36430, 16'd61194, 16'd54203, 16'd28161, 16'd17615, 16'd36995, 16'd8061, 16'd46891, 16'd27744, 16'd13319});
	test_expansion(128'ha23b03a22f209a76acaf0502bb2b9da3, {16'd63449, 16'd44699, 16'd63692, 16'd41496, 16'd52492, 16'd52792, 16'd44292, 16'd14923, 16'd19075, 16'd1819, 16'd3270, 16'd62694, 16'd17916, 16'd38184, 16'd51397, 16'd39580, 16'd47564, 16'd13458, 16'd5913, 16'd26538, 16'd33537, 16'd32899, 16'd26248, 16'd44961, 16'd34989, 16'd19453});
	test_expansion(128'h047656cfe1b289570c2bbe2af11ef088, {16'd11208, 16'd3632, 16'd64347, 16'd25095, 16'd12545, 16'd20733, 16'd7028, 16'd43712, 16'd46216, 16'd63026, 16'd11072, 16'd37276, 16'd32569, 16'd30678, 16'd58357, 16'd53346, 16'd47940, 16'd55142, 16'd28852, 16'd7693, 16'd20677, 16'd37885, 16'd24558, 16'd30706, 16'd28844, 16'd51788});
	test_expansion(128'h1bb875a40a1426f8933661370fe01826, {16'd1985, 16'd34323, 16'd61959, 16'd21240, 16'd15789, 16'd47380, 16'd14877, 16'd29227, 16'd32743, 16'd2759, 16'd25223, 16'd28688, 16'd34934, 16'd1302, 16'd54250, 16'd15431, 16'd26905, 16'd17372, 16'd43048, 16'd57381, 16'd60246, 16'd11994, 16'd41323, 16'd41907, 16'd63930, 16'd26128});
	test_expansion(128'h7a591f4ebcc6d61f54867d5ac6785111, {16'd27256, 16'd47156, 16'd61963, 16'd890, 16'd60297, 16'd43848, 16'd52263, 16'd33216, 16'd61904, 16'd21328, 16'd17463, 16'd43047, 16'd58183, 16'd41209, 16'd44016, 16'd36533, 16'd57561, 16'd50820, 16'd48891, 16'd10469, 16'd48112, 16'd48374, 16'd44095, 16'd8116, 16'd11192, 16'd40071});
	test_expansion(128'h825f668a265463995eb9d4ab6416e955, {16'd58355, 16'd45643, 16'd8980, 16'd34860, 16'd42284, 16'd43423, 16'd40910, 16'd34650, 16'd15018, 16'd51844, 16'd4350, 16'd23562, 16'd20253, 16'd2370, 16'd4452, 16'd39008, 16'd5113, 16'd50436, 16'd12621, 16'd17434, 16'd23493, 16'd59970, 16'd36309, 16'd13622, 16'd65055, 16'd54416});
	test_expansion(128'hf5fff09d0d927d03d5f24407967bd952, {16'd13307, 16'd35448, 16'd18944, 16'd58273, 16'd49843, 16'd40577, 16'd12843, 16'd29620, 16'd25843, 16'd62559, 16'd3351, 16'd32681, 16'd49693, 16'd36558, 16'd2020, 16'd13332, 16'd42457, 16'd8314, 16'd64710, 16'd62786, 16'd38932, 16'd39416, 16'd11279, 16'd25960, 16'd16834, 16'd52826});
	test_expansion(128'haf1c8c1f1543135b7ce3617e4cc80a83, {16'd17022, 16'd41477, 16'd51608, 16'd32689, 16'd52855, 16'd25415, 16'd31964, 16'd51258, 16'd34180, 16'd29314, 16'd58710, 16'd58375, 16'd62726, 16'd34860, 16'd34921, 16'd46293, 16'd39158, 16'd28560, 16'd50639, 16'd46252, 16'd96, 16'd32094, 16'd39532, 16'd44828, 16'd57150, 16'd4549});
	test_expansion(128'h1e2fdb665f2455385fbbfc8da085f99e, {16'd16962, 16'd57215, 16'd4536, 16'd63167, 16'd4240, 16'd4836, 16'd47855, 16'd27387, 16'd3730, 16'd39121, 16'd967, 16'd64836, 16'd27481, 16'd50720, 16'd34429, 16'd13497, 16'd41327, 16'd56007, 16'd11434, 16'd51420, 16'd31483, 16'd45413, 16'd10198, 16'd49268, 16'd55293, 16'd53259});
	test_expansion(128'he01c7fcf3faede096f0716b76ec97127, {16'd6306, 16'd44583, 16'd47393, 16'd42495, 16'd17070, 16'd28775, 16'd63566, 16'd25887, 16'd62473, 16'd14497, 16'd58141, 16'd64916, 16'd23206, 16'd64989, 16'd65092, 16'd8794, 16'd81, 16'd53868, 16'd8318, 16'd39894, 16'd43134, 16'd40417, 16'd43057, 16'd10930, 16'd63541, 16'd59080});
	test_expansion(128'h33c9c5545b09cfd809549bb0d08c095d, {16'd34920, 16'd42790, 16'd22111, 16'd52101, 16'd55124, 16'd45930, 16'd32635, 16'd16142, 16'd26248, 16'd60022, 16'd7604, 16'd62443, 16'd48887, 16'd13697, 16'd34058, 16'd36119, 16'd22488, 16'd26963, 16'd4567, 16'd24775, 16'd21354, 16'd49082, 16'd18741, 16'd60465, 16'd3120, 16'd51569});
	test_expansion(128'h05ff2e62a11e79e581823983357fa6fa, {16'd32839, 16'd6670, 16'd32684, 16'd13026, 16'd15338, 16'd4628, 16'd27686, 16'd52031, 16'd60895, 16'd52018, 16'd54946, 16'd25073, 16'd26518, 16'd19679, 16'd12648, 16'd33495, 16'd58257, 16'd49410, 16'd59469, 16'd29116, 16'd10713, 16'd26883, 16'd7214, 16'd59547, 16'd46409, 16'd26429});
	test_expansion(128'hb8275cfbefee5ae289a1530a95522573, {16'd22823, 16'd65448, 16'd31459, 16'd25828, 16'd23817, 16'd59913, 16'd44708, 16'd40799, 16'd122, 16'd12524, 16'd49102, 16'd21436, 16'd44650, 16'd17482, 16'd13280, 16'd52472, 16'd24999, 16'd16435, 16'd49989, 16'd56373, 16'd3097, 16'd14090, 16'd50922, 16'd22781, 16'd14569, 16'd12056});
	test_expansion(128'he4a2eb29dfa7b5091d00b1ca153f2be1, {16'd59269, 16'd34918, 16'd53015, 16'd33568, 16'd64002, 16'd8090, 16'd54007, 16'd52113, 16'd54292, 16'd62230, 16'd27046, 16'd59803, 16'd6997, 16'd44789, 16'd43511, 16'd676, 16'd16757, 16'd40348, 16'd41776, 16'd7320, 16'd60003, 16'd47168, 16'd2201, 16'd58060, 16'd22061, 16'd14367});
	test_expansion(128'he42a44c5e7105ea1653a430f372f621c, {16'd286, 16'd10278, 16'd65101, 16'd51095, 16'd63152, 16'd23245, 16'd41464, 16'd60288, 16'd61233, 16'd34551, 16'd9059, 16'd22028, 16'd11168, 16'd15692, 16'd18508, 16'd20091, 16'd9352, 16'd31273, 16'd51358, 16'd36148, 16'd23017, 16'd21832, 16'd55337, 16'd5878, 16'd61649, 16'd56159});
	test_expansion(128'h8f4ecc972066b01fd69b278ae19c312e, {16'd4415, 16'd3171, 16'd55493, 16'd53469, 16'd19834, 16'd39079, 16'd38512, 16'd63280, 16'd15780, 16'd2980, 16'd58859, 16'd28089, 16'd7653, 16'd49997, 16'd57721, 16'd58114, 16'd41318, 16'd15612, 16'd2656, 16'd7102, 16'd53144, 16'd27325, 16'd43022, 16'd18654, 16'd7186, 16'd32714});
	test_expansion(128'h7ff232a5c841f9e17bfe93155318f033, {16'd8993, 16'd50474, 16'd54298, 16'd64798, 16'd12506, 16'd14571, 16'd22014, 16'd24535, 16'd14015, 16'd55436, 16'd54338, 16'd63957, 16'd18986, 16'd35341, 16'd64494, 16'd62284, 16'd52484, 16'd19851, 16'd21751, 16'd62316, 16'd30552, 16'd57069, 16'd53650, 16'd542, 16'd520, 16'd14777});
	test_expansion(128'hfff3e49a3cab988fabebdd1122c30eb7, {16'd21610, 16'd32768, 16'd3081, 16'd23771, 16'd65510, 16'd14405, 16'd6726, 16'd56297, 16'd35584, 16'd48876, 16'd43267, 16'd41824, 16'd2226, 16'd14217, 16'd32422, 16'd52055, 16'd14150, 16'd31756, 16'd1373, 16'd29373, 16'd50777, 16'd1306, 16'd38062, 16'd31576, 16'd16852, 16'd3075});
	test_expansion(128'h4b1d4fbee1512aa546f48c84270ec888, {16'd14260, 16'd42664, 16'd16527, 16'd63544, 16'd14053, 16'd22568, 16'd57944, 16'd31272, 16'd48215, 16'd36649, 16'd49, 16'd4840, 16'd39412, 16'd3336, 16'd46913, 16'd10884, 16'd7081, 16'd27909, 16'd12262, 16'd3628, 16'd31662, 16'd7535, 16'd41142, 16'd58431, 16'd5565, 16'd33637});
	test_expansion(128'h4bfe94689d214eb9b6a33d94d5955646, {16'd12669, 16'd65407, 16'd8812, 16'd13902, 16'd31624, 16'd43255, 16'd41829, 16'd53086, 16'd6993, 16'd33354, 16'd39551, 16'd33011, 16'd817, 16'd64162, 16'd20424, 16'd17311, 16'd59671, 16'd34494, 16'd38463, 16'd61923, 16'd63323, 16'd63706, 16'd42893, 16'd24572, 16'd31806, 16'd53383});
	test_expansion(128'h5e5ea271a401da5b8d7747dc082822b2, {16'd64842, 16'd54958, 16'd4890, 16'd18927, 16'd17564, 16'd32805, 16'd38651, 16'd26701, 16'd55931, 16'd52809, 16'd31941, 16'd18277, 16'd38049, 16'd61212, 16'd49479, 16'd49277, 16'd30395, 16'd48607, 16'd39520, 16'd29389, 16'd15361, 16'd18640, 16'd59453, 16'd48569, 16'd39164, 16'd64366});
	test_expansion(128'h846c063c336e86b2eccf3ebf65cad307, {16'd39878, 16'd21940, 16'd38268, 16'd24532, 16'd12180, 16'd38525, 16'd62339, 16'd4986, 16'd54646, 16'd13962, 16'd16166, 16'd351, 16'd14969, 16'd48210, 16'd25747, 16'd611, 16'd444, 16'd42198, 16'd27293, 16'd1232, 16'd31072, 16'd10212, 16'd9066, 16'd40704, 16'd2240, 16'd1038});
	test_expansion(128'ha8a726a1004efce6285df2160997fbaf, {16'd39519, 16'd55633, 16'd46377, 16'd62692, 16'd980, 16'd4121, 16'd5069, 16'd34150, 16'd7658, 16'd4472, 16'd3022, 16'd29680, 16'd57352, 16'd36267, 16'd55453, 16'd65368, 16'd21010, 16'd17787, 16'd11626, 16'd49629, 16'd4299, 16'd35730, 16'd21756, 16'd2817, 16'd19943, 16'd40651});
	test_expansion(128'hc0e37a9ba9b091711217d3740f68c709, {16'd2406, 16'd20391, 16'd50267, 16'd52243, 16'd58749, 16'd48918, 16'd24601, 16'd52395, 16'd36896, 16'd46784, 16'd24861, 16'd20758, 16'd59070, 16'd10617, 16'd3656, 16'd15769, 16'd60257, 16'd34540, 16'd22734, 16'd19237, 16'd1891, 16'd9433, 16'd13052, 16'd16249, 16'd36198, 16'd51792});
	test_expansion(128'h7444599a2eb4933eba2ec9c354e779d4, {16'd864, 16'd7534, 16'd13132, 16'd544, 16'd39971, 16'd52575, 16'd35009, 16'd19907, 16'd61463, 16'd59851, 16'd52860, 16'd64492, 16'd23139, 16'd20649, 16'd17461, 16'd56268, 16'd41234, 16'd59216, 16'd1857, 16'd19413, 16'd51471, 16'd13072, 16'd63699, 16'd25883, 16'd31159, 16'd4261});
	test_expansion(128'h0a3fe808399e57f2718ef1de3abe4bde, {16'd55992, 16'd39364, 16'd43183, 16'd58722, 16'd16312, 16'd20182, 16'd48974, 16'd5933, 16'd26023, 16'd4300, 16'd53391, 16'd3340, 16'd51071, 16'd50946, 16'd10760, 16'd55353, 16'd61648, 16'd62586, 16'd50852, 16'd953, 16'd32548, 16'd48083, 16'd26297, 16'd20096, 16'd47093, 16'd18388});
	test_expansion(128'h6ba4ca7bb2067f314c3af6ed7758c1f4, {16'd37151, 16'd58118, 16'd15571, 16'd7397, 16'd3504, 16'd64300, 16'd100, 16'd64194, 16'd19081, 16'd14108, 16'd49798, 16'd10991, 16'd32247, 16'd21808, 16'd22967, 16'd63993, 16'd58113, 16'd52408, 16'd51613, 16'd17639, 16'd37357, 16'd60635, 16'd54625, 16'd38594, 16'd47264, 16'd7043});
	test_expansion(128'hacbe00d776a8faf3b613e35ba6c1e293, {16'd33413, 16'd29668, 16'd25701, 16'd14840, 16'd12965, 16'd19589, 16'd21596, 16'd55409, 16'd30314, 16'd62408, 16'd1959, 16'd43954, 16'd15607, 16'd33329, 16'd739, 16'd51348, 16'd43882, 16'd42278, 16'd39763, 16'd26012, 16'd46838, 16'd18102, 16'd46718, 16'd50588, 16'd21687, 16'd8547});
	test_expansion(128'h69e782b75f1cebcad9a205a5ac4d8694, {16'd1549, 16'd7732, 16'd40584, 16'd57473, 16'd1409, 16'd39132, 16'd39060, 16'd22159, 16'd34801, 16'd24801, 16'd60981, 16'd30162, 16'd51508, 16'd53065, 16'd29452, 16'd43510, 16'd32046, 16'd9761, 16'd64093, 16'd41037, 16'd8173, 16'd50489, 16'd34228, 16'd54917, 16'd31521, 16'd60203});
	test_expansion(128'h8167a6ea32837a30bce2612dd533ca55, {16'd19506, 16'd57176, 16'd20955, 16'd267, 16'd23619, 16'd24471, 16'd29551, 16'd34816, 16'd44330, 16'd50516, 16'd33725, 16'd27822, 16'd988, 16'd58476, 16'd50000, 16'd19053, 16'd59527, 16'd45989, 16'd6987, 16'd36368, 16'd65357, 16'd95, 16'd4335, 16'd38322, 16'd32790, 16'd18283});
	test_expansion(128'hc426d4d7e55adf990aafc8c8cef309d8, {16'd53325, 16'd65533, 16'd10574, 16'd13009, 16'd26809, 16'd56865, 16'd62830, 16'd57915, 16'd52384, 16'd39860, 16'd44186, 16'd18219, 16'd20803, 16'd2595, 16'd27633, 16'd60999, 16'd49296, 16'd64323, 16'd3676, 16'd47588, 16'd18784, 16'd11, 16'd11105, 16'd38838, 16'd20244, 16'd46149});
	test_expansion(128'hfa352f3d760302e80ef0d90420d6453a, {16'd22590, 16'd62713, 16'd24842, 16'd15043, 16'd60080, 16'd51770, 16'd62608, 16'd23859, 16'd20332, 16'd49112, 16'd11470, 16'd39929, 16'd26447, 16'd20602, 16'd31854, 16'd22734, 16'd65065, 16'd48600, 16'd2139, 16'd41214, 16'd11011, 16'd23188, 16'd49990, 16'd60801, 16'd44438, 16'd57311});
	test_expansion(128'he27c0167273a952eb939a364386f73f1, {16'd57422, 16'd33033, 16'd65102, 16'd8464, 16'd61689, 16'd21413, 16'd57613, 16'd743, 16'd1567, 16'd38625, 16'd39532, 16'd42642, 16'd29372, 16'd12874, 16'd40582, 16'd55050, 16'd2166, 16'd17265, 16'd60382, 16'd60756, 16'd32759, 16'd65366, 16'd50733, 16'd30761, 16'd710, 16'd27717});
	test_expansion(128'h4a90661e6316748ffe3191c89d5ca823, {16'd2420, 16'd46836, 16'd61895, 16'd58878, 16'd38141, 16'd39688, 16'd53748, 16'd28589, 16'd59336, 16'd57153, 16'd48630, 16'd45616, 16'd33906, 16'd27844, 16'd53581, 16'd27985, 16'd857, 16'd7820, 16'd50862, 16'd5783, 16'd53599, 16'd20858, 16'd33054, 16'd56673, 16'd45951, 16'd57573});
	test_expansion(128'hbaecea086a7a0662f278c79fe04bfdf4, {16'd57740, 16'd52341, 16'd30022, 16'd62236, 16'd10155, 16'd41294, 16'd31236, 16'd1279, 16'd46709, 16'd24707, 16'd29163, 16'd29688, 16'd20377, 16'd22678, 16'd60480, 16'd40528, 16'd11976, 16'd8768, 16'd10351, 16'd33622, 16'd48655, 16'd31973, 16'd36389, 16'd59448, 16'd48484, 16'd2200});
	test_expansion(128'he3fb2b0c67fb65e103ae8a07b22727c0, {16'd33385, 16'd59759, 16'd9338, 16'd12774, 16'd32242, 16'd7590, 16'd22743, 16'd7197, 16'd57086, 16'd48334, 16'd51573, 16'd49258, 16'd48383, 16'd40954, 16'd65517, 16'd57371, 16'd71, 16'd43720, 16'd9565, 16'd28957, 16'd65457, 16'd50542, 16'd2256, 16'd38831, 16'd13100, 16'd20092});
	test_expansion(128'h5a58d2a611aa45c5e9c832bcc718fbf3, {16'd6237, 16'd8813, 16'd44018, 16'd63099, 16'd25332, 16'd42463, 16'd57815, 16'd57115, 16'd16168, 16'd59776, 16'd57551, 16'd47395, 16'd7587, 16'd28268, 16'd53081, 16'd55813, 16'd25757, 16'd50881, 16'd41410, 16'd4359, 16'd30261, 16'd6021, 16'd46088, 16'd9667, 16'd11534, 16'd51490});
	test_expansion(128'h30192aa6f34c3ef43ec4848344279cab, {16'd45773, 16'd48131, 16'd13805, 16'd14213, 16'd61167, 16'd14028, 16'd39781, 16'd37599, 16'd28251, 16'd25569, 16'd24904, 16'd5205, 16'd15515, 16'd16684, 16'd36963, 16'd27891, 16'd39798, 16'd42106, 16'd11785, 16'd25015, 16'd14001, 16'd10600, 16'd22393, 16'd4588, 16'd18789, 16'd36622});
	test_expansion(128'hd4951c9ad825340cbf761b4b62fa33f5, {16'd50851, 16'd19904, 16'd54523, 16'd486, 16'd61940, 16'd43238, 16'd48008, 16'd20010, 16'd32964, 16'd48815, 16'd29740, 16'd29501, 16'd51260, 16'd18994, 16'd44545, 16'd3329, 16'd65393, 16'd3574, 16'd12157, 16'd18157, 16'd58823, 16'd10095, 16'd30813, 16'd57574, 16'd3913, 16'd15281});
	test_expansion(128'he1b1c034dfcd2b100dc6d6dcce8cf540, {16'd13271, 16'd6881, 16'd16897, 16'd17441, 16'd15536, 16'd29548, 16'd38701, 16'd63523, 16'd26780, 16'd11689, 16'd46716, 16'd62611, 16'd23886, 16'd54329, 16'd44341, 16'd22607, 16'd62137, 16'd9851, 16'd34768, 16'd1736, 16'd39109, 16'd40690, 16'd5945, 16'd36406, 16'd59400, 16'd56924});
	test_expansion(128'hc10e9f1de11253a539362e2710ea4b88, {16'd51781, 16'd47008, 16'd21863, 16'd24310, 16'd1894, 16'd63272, 16'd12928, 16'd51890, 16'd62122, 16'd59352, 16'd13411, 16'd59271, 16'd10774, 16'd38495, 16'd60474, 16'd16340, 16'd52844, 16'd3159, 16'd58258, 16'd29556, 16'd5775, 16'd22649, 16'd43026, 16'd3729, 16'd10963, 16'd9058});
	test_expansion(128'h1261159ac0cdab758c6153333fe062cc, {16'd48013, 16'd53849, 16'd8873, 16'd25837, 16'd6516, 16'd52392, 16'd17353, 16'd10787, 16'd56867, 16'd21565, 16'd26737, 16'd31484, 16'd44337, 16'd35180, 16'd650, 16'd43327, 16'd53567, 16'd24275, 16'd7357, 16'd56719, 16'd56761, 16'd42369, 16'd61146, 16'd43646, 16'd23324, 16'd11664});
	test_expansion(128'h8a3008b059607d0f26a484fa5e31e919, {16'd2987, 16'd2044, 16'd65276, 16'd36120, 16'd52035, 16'd6615, 16'd30920, 16'd31742, 16'd19168, 16'd20473, 16'd5300, 16'd9029, 16'd16778, 16'd23575, 16'd59356, 16'd16917, 16'd16688, 16'd523, 16'd60315, 16'd50738, 16'd29671, 16'd36930, 16'd32276, 16'd58797, 16'd51144, 16'd4855});
	test_expansion(128'h871135195aad2b5cf8038b6b4a9f7fbc, {16'd32990, 16'd37570, 16'd20315, 16'd16515, 16'd8305, 16'd45483, 16'd50669, 16'd31590, 16'd48993, 16'd17256, 16'd29178, 16'd53402, 16'd5234, 16'd65384, 16'd45168, 16'd35513, 16'd15657, 16'd61521, 16'd59890, 16'd2421, 16'd4118, 16'd46183, 16'd53259, 16'd27186, 16'd48397, 16'd8356});
	test_expansion(128'ha489f6b36b4a669c0859da4d3b1e451e, {16'd60552, 16'd20252, 16'd8660, 16'd11579, 16'd123, 16'd3697, 16'd25741, 16'd30131, 16'd16594, 16'd50176, 16'd64720, 16'd12988, 16'd50269, 16'd61505, 16'd18446, 16'd55967, 16'd4160, 16'd18970, 16'd47239, 16'd30473, 16'd7949, 16'd63491, 16'd28523, 16'd9271, 16'd56901, 16'd23877});
	test_expansion(128'h41b4f9a79bf2f2684573d0e70fdc090a, {16'd54830, 16'd48214, 16'd20153, 16'd5896, 16'd19903, 16'd32702, 16'd1429, 16'd55932, 16'd59932, 16'd29705, 16'd31022, 16'd59904, 16'd18746, 16'd61440, 16'd28605, 16'd1251, 16'd41807, 16'd6890, 16'd17181, 16'd27162, 16'd51990, 16'd27753, 16'd42903, 16'd3026, 16'd26750, 16'd28329});
	test_expansion(128'hdf560fbacc2efb5614b81e4b19c8c721, {16'd24198, 16'd39725, 16'd18444, 16'd4900, 16'd48045, 16'd27363, 16'd33655, 16'd25796, 16'd20306, 16'd14476, 16'd51825, 16'd62980, 16'd5206, 16'd49146, 16'd43563, 16'd21696, 16'd29807, 16'd22612, 16'd58852, 16'd31319, 16'd21289, 16'd48409, 16'd3126, 16'd54965, 16'd63619, 16'd59913});
	test_expansion(128'h0fe9a7fd243d98fb8ccf3d1a8c036a7d, {16'd7720, 16'd60354, 16'd33271, 16'd50687, 16'd30392, 16'd43634, 16'd50417, 16'd9877, 16'd32873, 16'd8888, 16'd52547, 16'd32186, 16'd45278, 16'd27078, 16'd41485, 16'd10297, 16'd49917, 16'd36749, 16'd7656, 16'd14368, 16'd42656, 16'd53108, 16'd4922, 16'd65379, 16'd62234, 16'd7772});
	test_expansion(128'h4a38bca8eeb23ada16a6266f8f8e89c5, {16'd3635, 16'd48641, 16'd2003, 16'd30210, 16'd49017, 16'd36065, 16'd58285, 16'd65297, 16'd26812, 16'd33175, 16'd15826, 16'd58634, 16'd59642, 16'd50422, 16'd20174, 16'd17855, 16'd20451, 16'd13158, 16'd47339, 16'd48258, 16'd46002, 16'd846, 16'd57142, 16'd2644, 16'd30426, 16'd54908});
	test_expansion(128'h5b91e7093e5f923d5c8d26f363309461, {16'd21855, 16'd33981, 16'd42530, 16'd31953, 16'd6942, 16'd35566, 16'd27192, 16'd11606, 16'd31023, 16'd55565, 16'd37800, 16'd31407, 16'd28407, 16'd17397, 16'd12598, 16'd58346, 16'd7767, 16'd44365, 16'd3864, 16'd43214, 16'd65478, 16'd49468, 16'd2519, 16'd29222, 16'd54409, 16'd44484});
	test_expansion(128'hfdfd44660d9974e56c8c608b97fecfbd, {16'd2238, 16'd34827, 16'd59765, 16'd28554, 16'd7717, 16'd47297, 16'd44431, 16'd6539, 16'd12623, 16'd7546, 16'd52789, 16'd4244, 16'd28274, 16'd10789, 16'd51644, 16'd5159, 16'd63372, 16'd58599, 16'd48435, 16'd55804, 16'd34675, 16'd45197, 16'd20088, 16'd9265, 16'd7214, 16'd30496});
	test_expansion(128'h04f4f9dbe3e80ad90f43e099ef276e46, {16'd44656, 16'd23388, 16'd14228, 16'd48389, 16'd34929, 16'd6359, 16'd2432, 16'd49192, 16'd55685, 16'd54728, 16'd54096, 16'd33319, 16'd63880, 16'd34449, 16'd31797, 16'd50957, 16'd13899, 16'd814, 16'd63359, 16'd4745, 16'd54704, 16'd31661, 16'd18039, 16'd3948, 16'd63405, 16'd43673});
	test_expansion(128'h489bdf0f486eabcd76faada04deb4a13, {16'd52674, 16'd65149, 16'd57682, 16'd54029, 16'd40192, 16'd7045, 16'd34141, 16'd56894, 16'd57732, 16'd56660, 16'd55133, 16'd36200, 16'd20058, 16'd17459, 16'd48028, 16'd3133, 16'd7729, 16'd30259, 16'd46384, 16'd6112, 16'd36471, 16'd63050, 16'd32829, 16'd24394, 16'd49924, 16'd38103});
	test_expansion(128'h22ec12ecd420fee4b5a8460212241b04, {16'd22360, 16'd4406, 16'd13524, 16'd53708, 16'd1757, 16'd6933, 16'd47873, 16'd9201, 16'd1824, 16'd63778, 16'd50201, 16'd57732, 16'd14997, 16'd59469, 16'd11585, 16'd6620, 16'd46579, 16'd19110, 16'd472, 16'd35479, 16'd17722, 16'd35084, 16'd22921, 16'd18414, 16'd20126, 16'd32954});
	test_expansion(128'hdd3c710528908e838e894a9f10c448dd, {16'd60874, 16'd62439, 16'd63748, 16'd42050, 16'd11655, 16'd41043, 16'd34713, 16'd24628, 16'd33573, 16'd44145, 16'd54333, 16'd64586, 16'd44523, 16'd63184, 16'd63574, 16'd55779, 16'd4763, 16'd42880, 16'd40432, 16'd24309, 16'd41094, 16'd29829, 16'd24331, 16'd64992, 16'd10715, 16'd51836});
	test_expansion(128'h4a5578819152e5e8991030c681501223, {16'd45496, 16'd27325, 16'd58519, 16'd8566, 16'd63791, 16'd46200, 16'd9646, 16'd47169, 16'd12695, 16'd35984, 16'd22838, 16'd33199, 16'd37236, 16'd44124, 16'd51528, 16'd60539, 16'd55355, 16'd25333, 16'd38440, 16'd5258, 16'd40761, 16'd1697, 16'd49430, 16'd11673, 16'd20561, 16'd44320});
	test_expansion(128'h3bd96cc809b1d52de077b3fb6621065c, {16'd56974, 16'd10664, 16'd32058, 16'd6577, 16'd22295, 16'd47824, 16'd36113, 16'd44822, 16'd19258, 16'd33180, 16'd49410, 16'd61067, 16'd45853, 16'd18242, 16'd59906, 16'd34178, 16'd53976, 16'd12958, 16'd22042, 16'd63521, 16'd47408, 16'd27510, 16'd39911, 16'd40724, 16'd39920, 16'd41288});
	test_expansion(128'hcffb801148eadad5eaa18fcdc5a952bf, {16'd40776, 16'd21887, 16'd21373, 16'd25605, 16'd28461, 16'd43411, 16'd43745, 16'd39777, 16'd53427, 16'd25792, 16'd11426, 16'd59003, 16'd46559, 16'd56308, 16'd2757, 16'd12202, 16'd2636, 16'd38495, 16'd21874, 16'd28724, 16'd5495, 16'd36754, 16'd21988, 16'd7667, 16'd27137, 16'd19029});
	test_expansion(128'h7964f406a418cd8f5a92cbfe6856b481, {16'd50061, 16'd9344, 16'd64929, 16'd45506, 16'd26337, 16'd31030, 16'd51972, 16'd55830, 16'd61682, 16'd36326, 16'd1602, 16'd39405, 16'd58559, 16'd52684, 16'd62336, 16'd11398, 16'd8600, 16'd49529, 16'd17816, 16'd1215, 16'd46014, 16'd11354, 16'd46008, 16'd43614, 16'd33402, 16'd22366});
	test_expansion(128'h9279ce554135f250996cebd0c9b70383, {16'd61828, 16'd55209, 16'd17234, 16'd23589, 16'd57059, 16'd54603, 16'd11096, 16'd28824, 16'd56885, 16'd24172, 16'd5237, 16'd55510, 16'd2355, 16'd617, 16'd28184, 16'd52501, 16'd14886, 16'd35538, 16'd51620, 16'd56114, 16'd11783, 16'd56093, 16'd49434, 16'd49684, 16'd58241, 16'd379});
	test_expansion(128'he3598403c2ef3fcb772d21492e050138, {16'd29680, 16'd14467, 16'd51806, 16'd45588, 16'd2364, 16'd20997, 16'd50000, 16'd60715, 16'd64106, 16'd1641, 16'd38936, 16'd12216, 16'd31353, 16'd18169, 16'd14176, 16'd19599, 16'd17246, 16'd60452, 16'd25006, 16'd14979, 16'd23615, 16'd19035, 16'd24462, 16'd33991, 16'd18714, 16'd39045});
	test_expansion(128'h925718386113743398fe19cec0386d09, {16'd52227, 16'd40405, 16'd55432, 16'd60400, 16'd25854, 16'd54083, 16'd47428, 16'd61570, 16'd40111, 16'd46659, 16'd1801, 16'd42232, 16'd20599, 16'd30679, 16'd36762, 16'd32178, 16'd22419, 16'd42042, 16'd41221, 16'd4892, 16'd28699, 16'd63534, 16'd6076, 16'd41659, 16'd52617, 16'd13318});
	test_expansion(128'h578d16e23784a7fd642e235c7cbd5fba, {16'd28306, 16'd8972, 16'd64029, 16'd35291, 16'd21217, 16'd56168, 16'd16945, 16'd54774, 16'd51632, 16'd7280, 16'd8210, 16'd63641, 16'd20552, 16'd20803, 16'd4646, 16'd13299, 16'd26946, 16'd18569, 16'd61327, 16'd4325, 16'd40099, 16'd29906, 16'd15970, 16'd13559, 16'd5840, 16'd35322});
	test_expansion(128'h6092254e627257b7d6707982f11ffcf7, {16'd25451, 16'd23752, 16'd30939, 16'd53236, 16'd9860, 16'd7042, 16'd57848, 16'd48109, 16'd53861, 16'd24628, 16'd7043, 16'd31929, 16'd21170, 16'd49167, 16'd49347, 16'd52821, 16'd38355, 16'd20210, 16'd29307, 16'd49069, 16'd63266, 16'd28783, 16'd7643, 16'd45342, 16'd47085, 16'd4003});
	test_expansion(128'hb4a7417e3a01020342b4e43f734218dc, {16'd12305, 16'd60628, 16'd34491, 16'd23401, 16'd48876, 16'd48306, 16'd64579, 16'd625, 16'd5512, 16'd61157, 16'd22594, 16'd58639, 16'd31250, 16'd14768, 16'd39077, 16'd46247, 16'd59085, 16'd44156, 16'd40866, 16'd17891, 16'd452, 16'd60799, 16'd56622, 16'd18295, 16'd35211, 16'd8718});
	test_expansion(128'hdf1d1af8480476bd99b6d633800e9cc5, {16'd4565, 16'd22351, 16'd61700, 16'd30553, 16'd21301, 16'd5526, 16'd61110, 16'd7444, 16'd62526, 16'd62496, 16'd56493, 16'd23810, 16'd57538, 16'd9128, 16'd4306, 16'd581, 16'd60290, 16'd26810, 16'd51187, 16'd12915, 16'd32604, 16'd8067, 16'd9723, 16'd46828, 16'd30640, 16'd64533});
	test_expansion(128'h6fd300ae207ba5b75b3527324d18c626, {16'd48974, 16'd55094, 16'd5746, 16'd53518, 16'd35587, 16'd9437, 16'd50304, 16'd20602, 16'd61371, 16'd5846, 16'd17860, 16'd49479, 16'd37026, 16'd5753, 16'd24079, 16'd1268, 16'd34899, 16'd35376, 16'd47887, 16'd18757, 16'd57683, 16'd6823, 16'd57812, 16'd28411, 16'd15608, 16'd27708});
	test_expansion(128'h73337b0f6e137c6f99cf60dff13fdb82, {16'd37953, 16'd11768, 16'd19772, 16'd48771, 16'd2399, 16'd55507, 16'd44914, 16'd40339, 16'd30805, 16'd12647, 16'd25228, 16'd54031, 16'd3541, 16'd45561, 16'd11829, 16'd52832, 16'd56934, 16'd11585, 16'd16892, 16'd41647, 16'd47785, 16'd25324, 16'd54247, 16'd23460, 16'd45487, 16'd56845});
	test_expansion(128'h96a03a857c4252354caa8a52378469fe, {16'd35595, 16'd65286, 16'd28884, 16'd57630, 16'd53411, 16'd18729, 16'd22843, 16'd12658, 16'd32597, 16'd51267, 16'd30336, 16'd19021, 16'd14407, 16'd6685, 16'd54610, 16'd23331, 16'd23922, 16'd24981, 16'd9136, 16'd617, 16'd27464, 16'd8658, 16'd15327, 16'd16304, 16'd45780, 16'd20383});
	test_expansion(128'hfd3548c511c94ea6bf0062c43470aa1e, {16'd43994, 16'd10035, 16'd12442, 16'd50497, 16'd54535, 16'd785, 16'd4880, 16'd1853, 16'd42519, 16'd48415, 16'd1364, 16'd12106, 16'd30262, 16'd52895, 16'd13572, 16'd10650, 16'd55012, 16'd6631, 16'd5319, 16'd64720, 16'd40591, 16'd43045, 16'd65092, 16'd62209, 16'd27547, 16'd33695});
	test_expansion(128'hacb146432688412161969c355b5c901f, {16'd62178, 16'd30741, 16'd62462, 16'd45848, 16'd62179, 16'd3296, 16'd42613, 16'd50534, 16'd48779, 16'd60307, 16'd1035, 16'd29525, 16'd63354, 16'd64586, 16'd35295, 16'd33842, 16'd28535, 16'd34514, 16'd33939, 16'd42845, 16'd13653, 16'd29815, 16'd63882, 16'd18489, 16'd27050, 16'd17626});
	test_expansion(128'h748d68c87541e299022db39f45315abe, {16'd22160, 16'd61085, 16'd15390, 16'd48280, 16'd19375, 16'd43455, 16'd60540, 16'd28293, 16'd5727, 16'd2429, 16'd1990, 16'd52639, 16'd8518, 16'd2117, 16'd34253, 16'd3905, 16'd32130, 16'd32083, 16'd32653, 16'd10566, 16'd52484, 16'd51569, 16'd61896, 16'd19980, 16'd5240, 16'd33578});
	test_expansion(128'hdf3572a7b33d1e9fa3ebf3f5fcbd9c9b, {16'd1324, 16'd7135, 16'd8562, 16'd1995, 16'd33755, 16'd40778, 16'd16871, 16'd49008, 16'd2451, 16'd15509, 16'd28333, 16'd39506, 16'd32450, 16'd30313, 16'd59854, 16'd41149, 16'd7661, 16'd23528, 16'd64655, 16'd35507, 16'd51433, 16'd33745, 16'd50536, 16'd56655, 16'd44701, 16'd43720});
	test_expansion(128'hbaacd04f071056b914030fd6bf5e8865, {16'd14812, 16'd59788, 16'd37027, 16'd37688, 16'd4684, 16'd37264, 16'd18691, 16'd15708, 16'd41390, 16'd4142, 16'd47482, 16'd48358, 16'd46165, 16'd52730, 16'd34498, 16'd43745, 16'd17654, 16'd13369, 16'd42721, 16'd48087, 16'd28590, 16'd34650, 16'd48413, 16'd20716, 16'd11669, 16'd50212});
	test_expansion(128'h16da52ef3fb561df6b1dd23ba7e9feef, {16'd17211, 16'd42152, 16'd25148, 16'd22295, 16'd25397, 16'd3397, 16'd34314, 16'd51940, 16'd9839, 16'd37650, 16'd62441, 16'd15282, 16'd35639, 16'd6857, 16'd19709, 16'd38311, 16'd50552, 16'd35586, 16'd11244, 16'd56884, 16'd14491, 16'd56121, 16'd14445, 16'd47643, 16'd38952, 16'd6413});
	test_expansion(128'ha59bc695c089b3955d53d72c45f5b7e8, {16'd56296, 16'd22884, 16'd31926, 16'd4813, 16'd31764, 16'd60526, 16'd5562, 16'd24565, 16'd6963, 16'd12772, 16'd38102, 16'd27397, 16'd46726, 16'd60293, 16'd40934, 16'd21977, 16'd46065, 16'd30266, 16'd34733, 16'd29473, 16'd19661, 16'd50289, 16'd38713, 16'd18074, 16'd33785, 16'd38871});
	test_expansion(128'h206c2f56ad9974e740dc4444ec9ad9ea, {16'd49270, 16'd22922, 16'd23415, 16'd64838, 16'd46274, 16'd23596, 16'd43058, 16'd20763, 16'd36603, 16'd52993, 16'd26419, 16'd54961, 16'd20519, 16'd51613, 16'd3982, 16'd18447, 16'd29834, 16'd51712, 16'd38863, 16'd14400, 16'd34427, 16'd64001, 16'd54322, 16'd21439, 16'd12851, 16'd16732});
	test_expansion(128'h110123c140fb7bac7b0998e0392b1158, {16'd9492, 16'd50961, 16'd3590, 16'd49346, 16'd13665, 16'd10632, 16'd28588, 16'd12669, 16'd23599, 16'd62207, 16'd55486, 16'd45118, 16'd30900, 16'd49971, 16'd5698, 16'd38931, 16'd17100, 16'd46688, 16'd53643, 16'd33026, 16'd22704, 16'd8576, 16'd24069, 16'd48180, 16'd34132, 16'd60271});
	test_expansion(128'h78e02009b8587702244f04a65c2085de, {16'd23187, 16'd1828, 16'd12716, 16'd47192, 16'd9188, 16'd56782, 16'd16367, 16'd62038, 16'd22490, 16'd65289, 16'd24310, 16'd32408, 16'd38353, 16'd37483, 16'd7627, 16'd38731, 16'd59048, 16'd52859, 16'd41816, 16'd3723, 16'd7371, 16'd16706, 16'd7553, 16'd11038, 16'd21594, 16'd54546});
	test_expansion(128'hf281e9280a8997799e0fea821faacb73, {16'd25738, 16'd31909, 16'd35864, 16'd10015, 16'd29416, 16'd17744, 16'd48568, 16'd4421, 16'd49767, 16'd33963, 16'd17725, 16'd58600, 16'd13341, 16'd8522, 16'd50940, 16'd62824, 16'd32231, 16'd32711, 16'd3023, 16'd27450, 16'd62472, 16'd5921, 16'd8152, 16'd20875, 16'd58131, 16'd52290});
	test_expansion(128'h309d64f8dfed895d873d8f47bbda7ebf, {16'd64670, 16'd6996, 16'd63098, 16'd14277, 16'd11231, 16'd8973, 16'd16517, 16'd10066, 16'd13713, 16'd62183, 16'd11663, 16'd58621, 16'd29075, 16'd3824, 16'd52071, 16'd51372, 16'd23778, 16'd1947, 16'd34976, 16'd33646, 16'd39463, 16'd32662, 16'd2140, 16'd43723, 16'd16842, 16'd14953});
	test_expansion(128'h501564ab27ede1879c991f003a350a65, {16'd50753, 16'd32972, 16'd55775, 16'd40806, 16'd16569, 16'd54114, 16'd40244, 16'd41098, 16'd11258, 16'd173, 16'd24848, 16'd20902, 16'd24684, 16'd55785, 16'd31927, 16'd47811, 16'd44785, 16'd56989, 16'd36211, 16'd43697, 16'd60207, 16'd3294, 16'd5302, 16'd6860, 16'd38503, 16'd60771});
	test_expansion(128'h9d6dd8d9ecee1d8618ba4c644cc7b42d, {16'd20189, 16'd12532, 16'd19509, 16'd29023, 16'd25536, 16'd41539, 16'd18203, 16'd6404, 16'd46039, 16'd13855, 16'd25838, 16'd53304, 16'd13020, 16'd40931, 16'd55722, 16'd51013, 16'd59650, 16'd2017, 16'd34016, 16'd60376, 16'd14766, 16'd4035, 16'd27891, 16'd63488, 16'd46731, 16'd37333});
	test_expansion(128'h9f68620785dc69d5b3f285f53196d743, {16'd50098, 16'd59441, 16'd7488, 16'd21901, 16'd16654, 16'd64892, 16'd10616, 16'd49895, 16'd53896, 16'd22302, 16'd50305, 16'd25676, 16'd47229, 16'd10073, 16'd62224, 16'd56918, 16'd58987, 16'd63238, 16'd61318, 16'd54467, 16'd9709, 16'd28654, 16'd30918, 16'd56191, 16'd58171, 16'd47120});
	test_expansion(128'h6f3e500ca4c4befe339d4ca573ca43c8, {16'd54936, 16'd37270, 16'd12428, 16'd59607, 16'd61311, 16'd9317, 16'd63897, 16'd31727, 16'd42129, 16'd46924, 16'd57923, 16'd33096, 16'd30692, 16'd58152, 16'd64738, 16'd37236, 16'd15055, 16'd35942, 16'd32136, 16'd46202, 16'd35545, 16'd14838, 16'd40632, 16'd3901, 16'd43438, 16'd14782});
	test_expansion(128'h8d870cfda94bd1c3e2110da9d0a7fbab, {16'd51858, 16'd23588, 16'd56845, 16'd21256, 16'd35700, 16'd14965, 16'd45774, 16'd3749, 16'd2149, 16'd39652, 16'd61459, 16'd42854, 16'd53851, 16'd15871, 16'd60182, 16'd23610, 16'd26830, 16'd38410, 16'd32789, 16'd30426, 16'd20244, 16'd49915, 16'd16187, 16'd3063, 16'd47976, 16'd1343});
	test_expansion(128'h00d62de710b5fc7e08064ae2756e95ce, {16'd13455, 16'd64280, 16'd37142, 16'd17033, 16'd283, 16'd35300, 16'd64271, 16'd49541, 16'd7821, 16'd36164, 16'd18068, 16'd20761, 16'd45443, 16'd25049, 16'd12977, 16'd41218, 16'd6310, 16'd57053, 16'd45049, 16'd11627, 16'd52492, 16'd10500, 16'd13460, 16'd17610, 16'd11715, 16'd51861});
	test_expansion(128'h5ca328748742b62cf2a6cf78517de556, {16'd47330, 16'd58067, 16'd8648, 16'd1637, 16'd38415, 16'd8201, 16'd2369, 16'd4833, 16'd28559, 16'd32064, 16'd44622, 16'd55078, 16'd35380, 16'd32216, 16'd21361, 16'd12843, 16'd47027, 16'd49692, 16'd10505, 16'd52198, 16'd45268, 16'd62225, 16'd36197, 16'd8704, 16'd27352, 16'd23955});
	test_expansion(128'he866114030cdc3362fa10ccafc1d8cc8, {16'd1611, 16'd48484, 16'd18836, 16'd9511, 16'd35791, 16'd50942, 16'd33097, 16'd46488, 16'd46903, 16'd22110, 16'd485, 16'd54074, 16'd52491, 16'd2378, 16'd56807, 16'd3300, 16'd47752, 16'd18454, 16'd13423, 16'd32232, 16'd42094, 16'd13779, 16'd45094, 16'd60513, 16'd6675, 16'd46743});
	test_expansion(128'h34432544a6d5dcfd64be4748b1271215, {16'd10506, 16'd55386, 16'd53742, 16'd56946, 16'd20507, 16'd47125, 16'd48272, 16'd49855, 16'd40974, 16'd58231, 16'd51530, 16'd5643, 16'd60783, 16'd14833, 16'd18640, 16'd19051, 16'd56378, 16'd24206, 16'd7934, 16'd7813, 16'd59521, 16'd13513, 16'd14833, 16'd48020, 16'd2674, 16'd65321});
	test_expansion(128'h0aa7fec1562daa6980c42528c3c8d01d, {16'd11358, 16'd40683, 16'd31443, 16'd29259, 16'd23547, 16'd65467, 16'd36829, 16'd33291, 16'd40968, 16'd22001, 16'd14494, 16'd50350, 16'd42253, 16'd41623, 16'd23796, 16'd30727, 16'd2617, 16'd18009, 16'd60465, 16'd28466, 16'd38248, 16'd251, 16'd2093, 16'd36515, 16'd27188, 16'd59921});
	test_expansion(128'ha26ab9c2d79962a3c412818d723614f0, {16'd3219, 16'd45000, 16'd56504, 16'd54258, 16'd12785, 16'd37908, 16'd59145, 16'd56856, 16'd59161, 16'd6833, 16'd44750, 16'd27680, 16'd52854, 16'd6517, 16'd32006, 16'd28256, 16'd35488, 16'd40260, 16'd37745, 16'd50573, 16'd22470, 16'd19564, 16'd62326, 16'd50544, 16'd15931, 16'd32010});
	test_expansion(128'h419bfc39808b3ffed277b569e60028c2, {16'd61790, 16'd56659, 16'd29807, 16'd9636, 16'd33826, 16'd33023, 16'd30395, 16'd61046, 16'd41557, 16'd6833, 16'd53286, 16'd37565, 16'd10088, 16'd17, 16'd4521, 16'd3364, 16'd3072, 16'd19231, 16'd41140, 16'd54439, 16'd16523, 16'd26545, 16'd45849, 16'd56140, 16'd1536, 16'd31118});
	test_expansion(128'h7a055741959331c5456aac7b030bf1b8, {16'd25075, 16'd37957, 16'd16385, 16'd42857, 16'd5623, 16'd33559, 16'd54194, 16'd42911, 16'd30371, 16'd30915, 16'd42353, 16'd25082, 16'd37021, 16'd58161, 16'd39986, 16'd40073, 16'd28320, 16'd43625, 16'd59093, 16'd4247, 16'd64137, 16'd12700, 16'd10368, 16'd53352, 16'd46, 16'd51033});
	test_expansion(128'h1f1684c44faf80eb654785ba2a4423d0, {16'd29616, 16'd52689, 16'd19765, 16'd46040, 16'd38878, 16'd27656, 16'd65264, 16'd33425, 16'd65311, 16'd17954, 16'd46176, 16'd14084, 16'd50160, 16'd45336, 16'd4511, 16'd18277, 16'd56162, 16'd10535, 16'd18941, 16'd50803, 16'd783, 16'd7201, 16'd50929, 16'd30831, 16'd47385, 16'd5951});
	test_expansion(128'h0698a0992821543730336578c858973b, {16'd60545, 16'd23311, 16'd42482, 16'd32428, 16'd46099, 16'd32454, 16'd53785, 16'd59297, 16'd40163, 16'd65189, 16'd9383, 16'd42353, 16'd64675, 16'd6341, 16'd50859, 16'd30692, 16'd13498, 16'd36865, 16'd44615, 16'd18541, 16'd10320, 16'd38710, 16'd62058, 16'd26159, 16'd39697, 16'd36089});
	test_expansion(128'h81ee0a85b13a7c0f9531ce1d3b811f55, {16'd42395, 16'd32477, 16'd25579, 16'd62223, 16'd40127, 16'd12942, 16'd14207, 16'd63971, 16'd17177, 16'd11864, 16'd39710, 16'd52697, 16'd19404, 16'd31099, 16'd29151, 16'd13175, 16'd8206, 16'd21305, 16'd41783, 16'd41262, 16'd6599, 16'd55497, 16'd19009, 16'd41656, 16'd23328, 16'd35748});
	test_expansion(128'ha79608ff3b41a3f12bef6844cfce55c4, {16'd51735, 16'd58382, 16'd49515, 16'd32264, 16'd29006, 16'd58440, 16'd60329, 16'd32565, 16'd62239, 16'd5815, 16'd35262, 16'd55806, 16'd58773, 16'd9445, 16'd13343, 16'd63224, 16'd28657, 16'd53050, 16'd9990, 16'd29872, 16'd17491, 16'd24288, 16'd62153, 16'd49910, 16'd31123, 16'd58612});
	test_expansion(128'he9710f42d435510b927121a6fb769b38, {16'd7441, 16'd11984, 16'd65172, 16'd12283, 16'd43689, 16'd29683, 16'd13521, 16'd60357, 16'd58448, 16'd51157, 16'd55234, 16'd25953, 16'd35071, 16'd53669, 16'd9010, 16'd59770, 16'd30674, 16'd44796, 16'd55187, 16'd31240, 16'd13533, 16'd4280, 16'd45464, 16'd56334, 16'd36550, 16'd4453});
	test_expansion(128'h7106c4896184af45bc3af18361ebfe81, {16'd10097, 16'd60469, 16'd47095, 16'd32139, 16'd50556, 16'd64929, 16'd22304, 16'd45912, 16'd61140, 16'd27546, 16'd21967, 16'd39584, 16'd35115, 16'd7284, 16'd12969, 16'd4348, 16'd24020, 16'd10765, 16'd51182, 16'd53383, 16'd7469, 16'd45207, 16'd20388, 16'd9710, 16'd56844, 16'd40176});
	test_expansion(128'h43e775369b4149682d0bb0249c2a093f, {16'd34177, 16'd44477, 16'd20618, 16'd58822, 16'd4068, 16'd32614, 16'd57125, 16'd59023, 16'd21609, 16'd1960, 16'd31799, 16'd40389, 16'd17502, 16'd7911, 16'd21815, 16'd36160, 16'd37996, 16'd41840, 16'd63975, 16'd21969, 16'd46886, 16'd54499, 16'd50086, 16'd15271, 16'd38781, 16'd55156});
	test_expansion(128'h7da307b417b5149d2b647945a52da7de, {16'd34763, 16'd33497, 16'd41653, 16'd47579, 16'd51982, 16'd61347, 16'd11536, 16'd60187, 16'd44153, 16'd26170, 16'd62294, 16'd62692, 16'd35551, 16'd4031, 16'd31469, 16'd32056, 16'd21773, 16'd2933, 16'd9524, 16'd52063, 16'd51146, 16'd48508, 16'd61889, 16'd26921, 16'd19706, 16'd34904});
	test_expansion(128'h45c5fccd7406ef47c24332b9f039ebf4, {16'd47212, 16'd62003, 16'd34962, 16'd60057, 16'd12069, 16'd19499, 16'd20590, 16'd21225, 16'd34509, 16'd26582, 16'd17105, 16'd13432, 16'd23821, 16'd19688, 16'd13819, 16'd14170, 16'd52378, 16'd64854, 16'd59688, 16'd45146, 16'd7919, 16'd45737, 16'd35604, 16'd18630, 16'd9867, 16'd33578});
	test_expansion(128'hf238e69e152d2d10a209fad3dfbe68a9, {16'd37937, 16'd29435, 16'd50193, 16'd45711, 16'd50201, 16'd39554, 16'd10086, 16'd2788, 16'd11611, 16'd57877, 16'd29533, 16'd64202, 16'd18258, 16'd59484, 16'd28027, 16'd52098, 16'd59324, 16'd6415, 16'd33370, 16'd11279, 16'd52626, 16'd60705, 16'd27083, 16'd42776, 16'd48276, 16'd11435});
	test_expansion(128'h4c071d11949ed48c5777957667b2b47e, {16'd48957, 16'd37991, 16'd18713, 16'd13206, 16'd55442, 16'd5458, 16'd29637, 16'd25384, 16'd21422, 16'd47529, 16'd26310, 16'd58677, 16'd445, 16'd41592, 16'd15802, 16'd46982, 16'd63803, 16'd21802, 16'd33485, 16'd16046, 16'd20777, 16'd52042, 16'd1163, 16'd15226, 16'd2367, 16'd7198});
	test_expansion(128'hf55bbef3b370456e57785c187691082b, {16'd53954, 16'd54350, 16'd25569, 16'd51502, 16'd21938, 16'd21803, 16'd28729, 16'd27183, 16'd9579, 16'd40406, 16'd36904, 16'd19834, 16'd49769, 16'd13667, 16'd15261, 16'd56003, 16'd31434, 16'd7321, 16'd41356, 16'd63858, 16'd16395, 16'd5363, 16'd31435, 16'd17423, 16'd2866, 16'd51076});
	test_expansion(128'h71655892eedf68254ec20ae49917ede1, {16'd4859, 16'd53057, 16'd48835, 16'd39834, 16'd38422, 16'd14247, 16'd57123, 16'd34185, 16'd47556, 16'd39988, 16'd37572, 16'd4658, 16'd42664, 16'd20032, 16'd9279, 16'd8698, 16'd35738, 16'd18907, 16'd59069, 16'd60463, 16'd7820, 16'd39906, 16'd21270, 16'd23297, 16'd30469, 16'd41567});
	test_expansion(128'hb4b29754984bcfb9fc0865c4c8c01fe3, {16'd22245, 16'd55807, 16'd850, 16'd63113, 16'd17813, 16'd56455, 16'd3932, 16'd44154, 16'd59272, 16'd13570, 16'd46701, 16'd10117, 16'd53376, 16'd3299, 16'd33677, 16'd16892, 16'd60621, 16'd27097, 16'd12820, 16'd46692, 16'd2367, 16'd42928, 16'd25323, 16'd11346, 16'd3572, 16'd16225});
	test_expansion(128'hc268648ab241bab5e3fee3af9c09c780, {16'd33189, 16'd60531, 16'd3465, 16'd1077, 16'd14720, 16'd47690, 16'd34673, 16'd43777, 16'd26064, 16'd32475, 16'd55302, 16'd15997, 16'd41052, 16'd27159, 16'd8960, 16'd24154, 16'd25696, 16'd17382, 16'd5471, 16'd30152, 16'd7796, 16'd43118, 16'd18945, 16'd46472, 16'd6214, 16'd830});
	test_expansion(128'h0c6f6a0a1818c8139b5744e1e087962c, {16'd178, 16'd2691, 16'd28217, 16'd60343, 16'd56942, 16'd51706, 16'd11987, 16'd59840, 16'd2274, 16'd57350, 16'd49385, 16'd22926, 16'd32898, 16'd51301, 16'd33316, 16'd14682, 16'd20146, 16'd44606, 16'd39537, 16'd49042, 16'd600, 16'd53462, 16'd59947, 16'd35937, 16'd44182, 16'd18259});
	test_expansion(128'h6eafa1d6deb865b80bfd260408b0ec40, {16'd659, 16'd14914, 16'd20375, 16'd4828, 16'd30465, 16'd65493, 16'd53348, 16'd13473, 16'd16461, 16'd20117, 16'd45389, 16'd13351, 16'd2702, 16'd3685, 16'd31858, 16'd46454, 16'd39453, 16'd19357, 16'd46064, 16'd55282, 16'd45348, 16'd8267, 16'd63776, 16'd15552, 16'd55734, 16'd49136});
	test_expansion(128'hac1bd935c0f988fde9eaacb0c702d60f, {16'd5225, 16'd21754, 16'd57289, 16'd17822, 16'd39686, 16'd35339, 16'd63157, 16'd16333, 16'd29671, 16'd61225, 16'd2535, 16'd39524, 16'd26632, 16'd57196, 16'd56062, 16'd55346, 16'd59221, 16'd6641, 16'd52693, 16'd44960, 16'd12339, 16'd46164, 16'd29073, 16'd17562, 16'd3346, 16'd57697});
	test_expansion(128'hb9e29699465bce612f5eb1d17e3d0ae0, {16'd32162, 16'd55043, 16'd25280, 16'd13244, 16'd28005, 16'd20314, 16'd32595, 16'd52678, 16'd39155, 16'd46849, 16'd24697, 16'd28885, 16'd27868, 16'd16161, 16'd14541, 16'd54617, 16'd32599, 16'd28993, 16'd38361, 16'd19098, 16'd2712, 16'd9194, 16'd55709, 16'd41379, 16'd31338, 16'd25487});
	test_expansion(128'hf39d0ed6b3cf9070bf7e1147914b8833, {16'd37925, 16'd2864, 16'd14332, 16'd8511, 16'd55724, 16'd32003, 16'd54236, 16'd48154, 16'd43159, 16'd8373, 16'd43509, 16'd54934, 16'd33097, 16'd47454, 16'd60912, 16'd45687, 16'd42244, 16'd17241, 16'd50356, 16'd53257, 16'd5231, 16'd57220, 16'd26151, 16'd43912, 16'd10705, 16'd26329});
	test_expansion(128'h676bf02c7da7e7d885280dbeb9338c99, {16'd37707, 16'd46117, 16'd25849, 16'd60880, 16'd17183, 16'd11407, 16'd50835, 16'd33271, 16'd42108, 16'd31970, 16'd15033, 16'd46701, 16'd42497, 16'd58813, 16'd45340, 16'd27640, 16'd5800, 16'd11486, 16'd62338, 16'd29714, 16'd33175, 16'd28687, 16'd13728, 16'd12978, 16'd104, 16'd37252});
	test_expansion(128'h54e22eaf0b9ecf1cb32c8dfc5b2282c9, {16'd29790, 16'd10989, 16'd10303, 16'd10606, 16'd9644, 16'd4550, 16'd29874, 16'd58402, 16'd25008, 16'd43776, 16'd21925, 16'd37517, 16'd14270, 16'd19515, 16'd38060, 16'd57942, 16'd725, 16'd33368, 16'd59121, 16'd44460, 16'd2563, 16'd55813, 16'd63807, 16'd19244, 16'd63703, 16'd41457});
	test_expansion(128'h8936431c868ba3186204d4b6924d32f1, {16'd59765, 16'd16831, 16'd50621, 16'd52936, 16'd16193, 16'd8623, 16'd21308, 16'd35360, 16'd56863, 16'd10186, 16'd24256, 16'd4176, 16'd45273, 16'd57707, 16'd44669, 16'd64916, 16'd62175, 16'd30653, 16'd5401, 16'd23361, 16'd64030, 16'd34083, 16'd49403, 16'd15423, 16'd53295, 16'd59603});
	test_expansion(128'h7cffd9bb4ea2978f09cfd8a199338756, {16'd36077, 16'd35795, 16'd3322, 16'd46670, 16'd46632, 16'd55910, 16'd54210, 16'd12485, 16'd65052, 16'd47134, 16'd55842, 16'd10081, 16'd60815, 16'd37523, 16'd22153, 16'd20270, 16'd26048, 16'd56253, 16'd25552, 16'd30036, 16'd11817, 16'd56677, 16'd9290, 16'd62121, 16'd60372, 16'd9680});
	test_expansion(128'hfc19e01c7a213119c207ca8bd388e7ee, {16'd65268, 16'd27776, 16'd5501, 16'd45907, 16'd38807, 16'd25002, 16'd7284, 16'd53508, 16'd29607, 16'd56062, 16'd60064, 16'd9077, 16'd9052, 16'd59519, 16'd1658, 16'd18470, 16'd35493, 16'd48782, 16'd28497, 16'd5162, 16'd37614, 16'd53386, 16'd64113, 16'd16869, 16'd6069, 16'd39806});
	test_expansion(128'h1e3ef7428c704cbe15f250ad62a2fa96, {16'd30332, 16'd28942, 16'd43501, 16'd6451, 16'd27345, 16'd19092, 16'd43818, 16'd35249, 16'd44687, 16'd39711, 16'd27322, 16'd1438, 16'd51615, 16'd62366, 16'd50009, 16'd43759, 16'd51206, 16'd7215, 16'd54855, 16'd21885, 16'd31822, 16'd20719, 16'd44836, 16'd32827, 16'd52869, 16'd37663});
	test_expansion(128'hfa135bf6c87ff158d2ab37dc2f69da89, {16'd31300, 16'd17008, 16'd64459, 16'd27118, 16'd43587, 16'd64292, 16'd1970, 16'd54559, 16'd15513, 16'd6842, 16'd47788, 16'd22555, 16'd32633, 16'd50760, 16'd16410, 16'd42839, 16'd12849, 16'd14122, 16'd10052, 16'd28836, 16'd22971, 16'd57045, 16'd13781, 16'd20220, 16'd55071, 16'd26955});
	test_expansion(128'he7974d646794e0fae7ad5e31c82be8fd, {16'd25480, 16'd34958, 16'd9726, 16'd17542, 16'd60940, 16'd24500, 16'd3015, 16'd34219, 16'd64220, 16'd35548, 16'd30742, 16'd48553, 16'd58245, 16'd44807, 16'd55083, 16'd29838, 16'd38830, 16'd38295, 16'd10686, 16'd27775, 16'd36962, 16'd40165, 16'd14064, 16'd50619, 16'd2043, 16'd42419});
	test_expansion(128'hfab262e6ef188bcae64293ccbf25ea1d, {16'd24771, 16'd27665, 16'd6896, 16'd31728, 16'd43356, 16'd52792, 16'd36329, 16'd47853, 16'd53830, 16'd7457, 16'd1081, 16'd12723, 16'd1560, 16'd50564, 16'd55707, 16'd15865, 16'd10041, 16'd41862, 16'd31302, 16'd53662, 16'd59409, 16'd60712, 16'd23367, 16'd2610, 16'd15656, 16'd62613});
	test_expansion(128'hb6c97d41ad39b4433c4e5265c4d930de, {16'd65347, 16'd209, 16'd24732, 16'd6215, 16'd21493, 16'd3308, 16'd26556, 16'd5648, 16'd43688, 16'd35653, 16'd39840, 16'd11900, 16'd52041, 16'd13528, 16'd20565, 16'd39781, 16'd16917, 16'd35547, 16'd58837, 16'd62692, 16'd2855, 16'd60111, 16'd699, 16'd48107, 16'd25312, 16'd20180});
	test_expansion(128'hf4616c311d87075e774b6c018040f7bc, {16'd19338, 16'd29829, 16'd49028, 16'd50727, 16'd32653, 16'd55262, 16'd41948, 16'd7336, 16'd2728, 16'd14536, 16'd9637, 16'd15505, 16'd37583, 16'd50316, 16'd22658, 16'd6533, 16'd35314, 16'd12053, 16'd38, 16'd3956, 16'd31136, 16'd25776, 16'd7850, 16'd29825, 16'd16506, 16'd43631});
	test_expansion(128'hf17e74204166974742ef2eaee0e3c93c, {16'd44300, 16'd2149, 16'd50240, 16'd14587, 16'd10592, 16'd19788, 16'd64983, 16'd15576, 16'd5774, 16'd62307, 16'd460, 16'd56185, 16'd34621, 16'd12454, 16'd18000, 16'd36430, 16'd7495, 16'd54934, 16'd15173, 16'd48864, 16'd21972, 16'd45920, 16'd25511, 16'd60895, 16'd29522, 16'd58348});
	test_expansion(128'h196bf94db086403e279e057d71fdd099, {16'd43391, 16'd27235, 16'd62320, 16'd951, 16'd77, 16'd15270, 16'd28514, 16'd42962, 16'd16845, 16'd16948, 16'd2420, 16'd20332, 16'd38299, 16'd9058, 16'd16208, 16'd36229, 16'd9681, 16'd13103, 16'd41620, 16'd63936, 16'd42997, 16'd5446, 16'd32881, 16'd44678, 16'd10976, 16'd63240});
	test_expansion(128'h29ddff00b8d91c6d45a4e02dba33971d, {16'd32920, 16'd64396, 16'd5744, 16'd21477, 16'd10616, 16'd21990, 16'd44389, 16'd53726, 16'd19641, 16'd18360, 16'd201, 16'd22675, 16'd62733, 16'd1569, 16'd7270, 16'd18097, 16'd50474, 16'd8022, 16'd32710, 16'd28420, 16'd16489, 16'd30266, 16'd11326, 16'd12052, 16'd30303, 16'd37090});
	test_expansion(128'h3dff376da78072f475ead75e79dad833, {16'd4659, 16'd22341, 16'd46580, 16'd15316, 16'd26171, 16'd15418, 16'd36229, 16'd47738, 16'd45511, 16'd43326, 16'd28335, 16'd4711, 16'd37869, 16'd50161, 16'd28677, 16'd24885, 16'd60999, 16'd18688, 16'd7950, 16'd9933, 16'd51305, 16'd29508, 16'd38401, 16'd32815, 16'd5874, 16'd61406});
	test_expansion(128'h66957d37842fbe25a44583bb882f6e75, {16'd16739, 16'd42207, 16'd38819, 16'd35023, 16'd57658, 16'd53956, 16'd58624, 16'd58735, 16'd2770, 16'd7703, 16'd684, 16'd46644, 16'd37790, 16'd21328, 16'd48154, 16'd53255, 16'd7001, 16'd5075, 16'd9369, 16'd39457, 16'd27341, 16'd32243, 16'd64770, 16'd40938, 16'd41507, 16'd5944});
	test_expansion(128'h7064eb460589e9dac583f2ec1b16df81, {16'd4312, 16'd52369, 16'd18999, 16'd25817, 16'd29374, 16'd46527, 16'd65470, 16'd3858, 16'd35151, 16'd21830, 16'd60205, 16'd33593, 16'd31690, 16'd39456, 16'd59505, 16'd17811, 16'd56735, 16'd18, 16'd3037, 16'd56048, 16'd39897, 16'd13244, 16'd30107, 16'd54025, 16'd54052, 16'd64129});
	test_expansion(128'hba28708ab82f6aa09f2a5c5c1ff10e62, {16'd39860, 16'd60120, 16'd26049, 16'd878, 16'd27386, 16'd63274, 16'd38675, 16'd8429, 16'd7835, 16'd1715, 16'd54773, 16'd14473, 16'd28127, 16'd63334, 16'd27042, 16'd8382, 16'd9220, 16'd45946, 16'd52694, 16'd33328, 16'd30993, 16'd28366, 16'd23747, 16'd42960, 16'd38359, 16'd60609});
	test_expansion(128'he8985f148953aab9a77a1d05b7e6309f, {16'd49852, 16'd10479, 16'd58172, 16'd48555, 16'd53898, 16'd26593, 16'd39280, 16'd40849, 16'd37439, 16'd32836, 16'd53408, 16'd24543, 16'd57307, 16'd51763, 16'd61301, 16'd8709, 16'd16822, 16'd49990, 16'd62816, 16'd9799, 16'd53264, 16'd14120, 16'd29893, 16'd1150, 16'd7710, 16'd46094});
	test_expansion(128'h2169fa08db2c05fd97a5660a58e283df, {16'd51420, 16'd34933, 16'd15113, 16'd11949, 16'd36354, 16'd4130, 16'd19833, 16'd59742, 16'd8200, 16'd32706, 16'd52926, 16'd59515, 16'd14568, 16'd33937, 16'd39823, 16'd9313, 16'd62507, 16'd50583, 16'd34906, 16'd31873, 16'd9153, 16'd63390, 16'd43097, 16'd63737, 16'd7665, 16'd27139});
	test_expansion(128'hc8645d19b78a7442a63249cb42fd4bd7, {16'd20495, 16'd48392, 16'd24990, 16'd22517, 16'd33398, 16'd7082, 16'd1077, 16'd27235, 16'd16660, 16'd43349, 16'd37180, 16'd20790, 16'd19515, 16'd38246, 16'd53656, 16'd46871, 16'd23542, 16'd27684, 16'd24252, 16'd30368, 16'd64329, 16'd10531, 16'd25978, 16'd61234, 16'd31841, 16'd15609});
	test_expansion(128'h9b3a25841553307bd38bb744827d1e9b, {16'd297, 16'd19964, 16'd62876, 16'd16319, 16'd60822, 16'd14278, 16'd29402, 16'd28548, 16'd5455, 16'd65196, 16'd26448, 16'd37787, 16'd46159, 16'd22912, 16'd27917, 16'd54119, 16'd7147, 16'd45900, 16'd55132, 16'd5813, 16'd56319, 16'd61801, 16'd19336, 16'd23885, 16'd65245, 16'd36875});
	test_expansion(128'hdd3d9e0231aa0e52683f4e29519449f5, {16'd61302, 16'd23128, 16'd52742, 16'd14069, 16'd5972, 16'd47009, 16'd21556, 16'd3334, 16'd21639, 16'd10261, 16'd543, 16'd28544, 16'd39354, 16'd15551, 16'd45737, 16'd24662, 16'd56783, 16'd14216, 16'd8252, 16'd60124, 16'd45771, 16'd61061, 16'd45792, 16'd84, 16'd7316, 16'd51487});
	test_expansion(128'h5f35694335aee5af5630b4fa44f5445a, {16'd16585, 16'd48832, 16'd44607, 16'd16188, 16'd28184, 16'd42775, 16'd23706, 16'd20429, 16'd30993, 16'd13335, 16'd12208, 16'd16135, 16'd65221, 16'd3903, 16'd59484, 16'd44271, 16'd48466, 16'd26759, 16'd459, 16'd40022, 16'd43218, 16'd12263, 16'd25545, 16'd60183, 16'd8849, 16'd2049});
	test_expansion(128'hc903b8d296f17224ec79b5b543a1e7fa, {16'd27314, 16'd26467, 16'd32978, 16'd16430, 16'd29461, 16'd46925, 16'd17541, 16'd3917, 16'd36026, 16'd9915, 16'd45627, 16'd37613, 16'd29113, 16'd45241, 16'd56185, 16'd24542, 16'd9282, 16'd24042, 16'd60030, 16'd53077, 16'd57015, 16'd6594, 16'd57906, 16'd27625, 16'd254, 16'd31933});
	test_expansion(128'h0e22e278aa1013d15d7b1a52d2cf2012, {16'd29697, 16'd20759, 16'd37912, 16'd12710, 16'd40441, 16'd20675, 16'd45532, 16'd38361, 16'd19893, 16'd49444, 16'd36372, 16'd9566, 16'd41874, 16'd38698, 16'd64075, 16'd44715, 16'd14777, 16'd8015, 16'd19727, 16'd57576, 16'd23094, 16'd33125, 16'd44533, 16'd42471, 16'd64647, 16'd24075});
	test_expansion(128'h6b793fecde904791da255bb70440ed8b, {16'd61223, 16'd63494, 16'd20550, 16'd58956, 16'd4535, 16'd2271, 16'd11274, 16'd51160, 16'd12132, 16'd35230, 16'd8036, 16'd56858, 16'd52230, 16'd52910, 16'd49150, 16'd15545, 16'd7224, 16'd20125, 16'd15817, 16'd15040, 16'd63528, 16'd4239, 16'd24183, 16'd64704, 16'd10530, 16'd57911});
	test_expansion(128'h10f2347d1626be2c68f22a1c23edf016, {16'd34411, 16'd46964, 16'd4296, 16'd35472, 16'd50029, 16'd61379, 16'd27207, 16'd58835, 16'd50188, 16'd32911, 16'd45807, 16'd36406, 16'd32403, 16'd4920, 16'd50074, 16'd58788, 16'd26669, 16'd52506, 16'd33798, 16'd12394, 16'd60697, 16'd20636, 16'd7460, 16'd26263, 16'd31987, 16'd7949});
	test_expansion(128'h41b1304e206513e9037af64d811d9bfe, {16'd19738, 16'd60712, 16'd43752, 16'd37083, 16'd61674, 16'd50418, 16'd24689, 16'd25949, 16'd56244, 16'd22790, 16'd8519, 16'd45092, 16'd43474, 16'd18052, 16'd38721, 16'd9508, 16'd53070, 16'd18462, 16'd18463, 16'd56140, 16'd41646, 16'd45130, 16'd52243, 16'd20349, 16'd10517, 16'd25427});
	test_expansion(128'hbd211713b0f28807c4a99a0949fa4916, {16'd31236, 16'd52868, 16'd5206, 16'd27238, 16'd49018, 16'd65148, 16'd18551, 16'd35402, 16'd23706, 16'd38115, 16'd42171, 16'd9133, 16'd58186, 16'd16526, 16'd50339, 16'd1597, 16'd41562, 16'd18990, 16'd4958, 16'd61575, 16'd56688, 16'd31320, 16'd16264, 16'd22903, 16'd43719, 16'd47072});
	test_expansion(128'h392b410bdf33b211ec98f82ee991e0f8, {16'd27206, 16'd60438, 16'd6061, 16'd8330, 16'd29471, 16'd45173, 16'd45991, 16'd32291, 16'd30659, 16'd13072, 16'd43436, 16'd10124, 16'd54116, 16'd28967, 16'd49338, 16'd41400, 16'd54379, 16'd20534, 16'd32727, 16'd12181, 16'd65229, 16'd64277, 16'd22106, 16'd16739, 16'd16789, 16'd63448});
	test_expansion(128'hb1cff008a55aba4612c3554f6cfd673f, {16'd61454, 16'd8523, 16'd60591, 16'd32788, 16'd15469, 16'd37028, 16'd54546, 16'd28687, 16'd46401, 16'd65316, 16'd28627, 16'd9981, 16'd36357, 16'd2937, 16'd31, 16'd5562, 16'd19816, 16'd28805, 16'd43747, 16'd14153, 16'd43754, 16'd7587, 16'd55340, 16'd1004, 16'd15147, 16'd33387});
	test_expansion(128'hfc9292b9862d2b65a9d31fbbc9f965b6, {16'd50124, 16'd18286, 16'd54948, 16'd8243, 16'd62115, 16'd27845, 16'd19344, 16'd9824, 16'd11235, 16'd1358, 16'd36963, 16'd8520, 16'd44571, 16'd14019, 16'd58859, 16'd47270, 16'd15475, 16'd7661, 16'd6729, 16'd13188, 16'd33777, 16'd6109, 16'd44866, 16'd58057, 16'd1064, 16'd27583});
	test_expansion(128'hd9d9046c4306f0b1066f1a5858ab2fd4, {16'd30677, 16'd54305, 16'd1297, 16'd51146, 16'd48121, 16'd29865, 16'd46578, 16'd65277, 16'd64942, 16'd22885, 16'd17061, 16'd64038, 16'd16507, 16'd15777, 16'd55536, 16'd56994, 16'd21485, 16'd46714, 16'd63831, 16'd2716, 16'd4512, 16'd48308, 16'd57833, 16'd29302, 16'd9712, 16'd13693});
	test_expansion(128'hf6a1b991741db7718e812705563c9f13, {16'd56960, 16'd43819, 16'd23565, 16'd21037, 16'd24435, 16'd14882, 16'd2939, 16'd35779, 16'd52919, 16'd20194, 16'd15953, 16'd53405, 16'd61735, 16'd12653, 16'd44948, 16'd38102, 16'd9196, 16'd48379, 16'd19856, 16'd11120, 16'd21491, 16'd36580, 16'd25620, 16'd57743, 16'd37035, 16'd50491});
	test_expansion(128'hb4c2deb1d37d88abf6e41b4cc8a21a2f, {16'd30490, 16'd16910, 16'd21555, 16'd61149, 16'd6697, 16'd104, 16'd5730, 16'd52333, 16'd21420, 16'd24448, 16'd742, 16'd15595, 16'd33644, 16'd1760, 16'd8440, 16'd19693, 16'd62180, 16'd16103, 16'd36913, 16'd18366, 16'd16876, 16'd28192, 16'd53656, 16'd8684, 16'd8273, 16'd26411});
	test_expansion(128'h16538b1225329b9329a97fd14e0fe684, {16'd47941, 16'd13359, 16'd7769, 16'd60639, 16'd31078, 16'd47251, 16'd57997, 16'd36690, 16'd41705, 16'd15893, 16'd17310, 16'd10603, 16'd42482, 16'd310, 16'd41384, 16'd48943, 16'd50632, 16'd37357, 16'd53553, 16'd16199, 16'd6294, 16'd20748, 16'd26825, 16'd56279, 16'd28916, 16'd40982});
	test_expansion(128'h5b302923d872c6efea33c18b5eb5ddc3, {16'd28721, 16'd9243, 16'd57874, 16'd64172, 16'd27705, 16'd33165, 16'd35899, 16'd4607, 16'd30312, 16'd51324, 16'd27332, 16'd59036, 16'd34669, 16'd21772, 16'd58587, 16'd3852, 16'd61181, 16'd18128, 16'd54755, 16'd17030, 16'd4178, 16'd13058, 16'd48616, 16'd29188, 16'd8920, 16'd14507});
	test_expansion(128'ha0f0db15fd33ce3ddd411994b3a577ed, {16'd53472, 16'd13599, 16'd26608, 16'd52207, 16'd59258, 16'd39430, 16'd61578, 16'd7477, 16'd24521, 16'd8570, 16'd37193, 16'd12915, 16'd24755, 16'd54357, 16'd41133, 16'd21691, 16'd56804, 16'd31289, 16'd50191, 16'd38188, 16'd48432, 16'd18219, 16'd62217, 16'd24294, 16'd30382, 16'd22755});
	test_expansion(128'hd27ca803694e1e824e5060891f150847, {16'd51662, 16'd52578, 16'd21497, 16'd24887, 16'd56186, 16'd37814, 16'd33319, 16'd785, 16'd1909, 16'd13148, 16'd56720, 16'd18661, 16'd47947, 16'd32490, 16'd61218, 16'd34311, 16'd29480, 16'd60245, 16'd10843, 16'd14735, 16'd48909, 16'd61194, 16'd53186, 16'd46647, 16'd11105, 16'd13159});
	test_expansion(128'h42c293e44a7a9ab38822ddb1a15599b5, {16'd22954, 16'd33216, 16'd16888, 16'd21436, 16'd35490, 16'd16076, 16'd15670, 16'd13662, 16'd12046, 16'd36664, 16'd38403, 16'd27282, 16'd33580, 16'd23190, 16'd27526, 16'd4990, 16'd30010, 16'd48191, 16'd51663, 16'd12723, 16'd38595, 16'd63342, 16'd24564, 16'd60631, 16'd17831, 16'd56351});
	test_expansion(128'h6e59ae5e6ac87b0f5587f799eaaf5f95, {16'd59257, 16'd47775, 16'd60976, 16'd42343, 16'd25415, 16'd56711, 16'd19726, 16'd63667, 16'd11628, 16'd41255, 16'd38924, 16'd32393, 16'd12859, 16'd65151, 16'd7622, 16'd63908, 16'd264, 16'd3106, 16'd56923, 16'd3545, 16'd5124, 16'd52103, 16'd48181, 16'd51574, 16'd20972, 16'd49982});
	test_expansion(128'h501fd0dea44097863b8ed999988aa5a5, {16'd36454, 16'd53917, 16'd64608, 16'd16923, 16'd35773, 16'd20178, 16'd25263, 16'd54900, 16'd16393, 16'd19016, 16'd53473, 16'd26733, 16'd10420, 16'd41477, 16'd4110, 16'd1548, 16'd44165, 16'd35874, 16'd20751, 16'd33218, 16'd32802, 16'd44563, 16'd5959, 16'd46289, 16'd45581, 16'd40991});
	test_expansion(128'h9d10b2405cb3cf601ac66d56d89e8810, {16'd4231, 16'd62532, 16'd2088, 16'd54569, 16'd67, 16'd1618, 16'd29475, 16'd57927, 16'd31194, 16'd27802, 16'd58881, 16'd39459, 16'd4358, 16'd54942, 16'd61640, 16'd29971, 16'd63758, 16'd28563, 16'd58375, 16'd57054, 16'd42633, 16'd15016, 16'd37892, 16'd19796, 16'd16405, 16'd101});
	test_expansion(128'hf1ac77c29e29c98178603b5992bda7a9, {16'd24353, 16'd37563, 16'd6372, 16'd49260, 16'd55510, 16'd30716, 16'd27410, 16'd6183, 16'd48248, 16'd40886, 16'd55590, 16'd20413, 16'd476, 16'd8474, 16'd7660, 16'd41249, 16'd12403, 16'd20152, 16'd12578, 16'd47690, 16'd37313, 16'd29798, 16'd58811, 16'd48611, 16'd64048, 16'd8401});
	test_expansion(128'h6364d1baef546183648aeab8a5a132ec, {16'd54092, 16'd17678, 16'd60392, 16'd29447, 16'd45811, 16'd30534, 16'd24097, 16'd21554, 16'd64896, 16'd55129, 16'd2994, 16'd38061, 16'd51847, 16'd23112, 16'd45154, 16'd28246, 16'd64352, 16'd57035, 16'd26697, 16'd10330, 16'd44129, 16'd63038, 16'd29400, 16'd57352, 16'd37016, 16'd49976});
	test_expansion(128'h92fce416f3b4192215545cde7378cc0d, {16'd39383, 16'd29343, 16'd59752, 16'd44040, 16'd55428, 16'd26801, 16'd864, 16'd47192, 16'd4956, 16'd4927, 16'd56458, 16'd59280, 16'd47206, 16'd5640, 16'd63966, 16'd25454, 16'd22925, 16'd11113, 16'd29910, 16'd30580, 16'd63210, 16'd28674, 16'd37992, 16'd2690, 16'd37030, 16'd38799});
	test_expansion(128'ha1e0a6bf957e6f37b8d440de8d82fec1, {16'd49990, 16'd34450, 16'd60528, 16'd39250, 16'd22724, 16'd4998, 16'd42291, 16'd29507, 16'd36338, 16'd55055, 16'd12907, 16'd26566, 16'd64891, 16'd5869, 16'd7575, 16'd5843, 16'd8249, 16'd30675, 16'd60235, 16'd28004, 16'd35343, 16'd12876, 16'd58401, 16'd57326, 16'd30626, 16'd10936});
	test_expansion(128'h8f837016c4687bb74613a132fa894ec7, {16'd46625, 16'd27691, 16'd48793, 16'd20588, 16'd30173, 16'd50172, 16'd7440, 16'd41441, 16'd13451, 16'd39965, 16'd18780, 16'd37481, 16'd25348, 16'd34953, 16'd2231, 16'd61085, 16'd59166, 16'd27532, 16'd45026, 16'd21019, 16'd22043, 16'd20910, 16'd54578, 16'd33890, 16'd10299, 16'd18679});
	test_expansion(128'h70f8c09d9131fee6574317030a22bfd0, {16'd39303, 16'd40551, 16'd3943, 16'd1980, 16'd49124, 16'd64552, 16'd64700, 16'd33582, 16'd40141, 16'd32320, 16'd64788, 16'd11106, 16'd54910, 16'd12817, 16'd5386, 16'd5432, 16'd9354, 16'd37053, 16'd19163, 16'd42217, 16'd58037, 16'd6132, 16'd24081, 16'd8699, 16'd38318, 16'd28819});
	test_expansion(128'hfa3749e87101c79016dae77e9287bfd9, {16'd28450, 16'd10504, 16'd4253, 16'd18877, 16'd50309, 16'd12220, 16'd13263, 16'd38452, 16'd11477, 16'd45821, 16'd41493, 16'd54142, 16'd64542, 16'd31109, 16'd64079, 16'd17481, 16'd64092, 16'd36360, 16'd38283, 16'd20409, 16'd34616, 16'd3364, 16'd45205, 16'd46188, 16'd23498, 16'd16773});
	test_expansion(128'h327cfff1fbde212c55019a6fbf5e287f, {16'd54810, 16'd44299, 16'd41945, 16'd35209, 16'd49161, 16'd61752, 16'd6697, 16'd42729, 16'd37598, 16'd43574, 16'd43422, 16'd39262, 16'd23491, 16'd56252, 16'd46311, 16'd42475, 16'd1949, 16'd15320, 16'd3536, 16'd43507, 16'd41492, 16'd33165, 16'd10697, 16'd42739, 16'd44883, 16'd47341});
	test_expansion(128'hf7e1b03e182168df2ba3217dadde7317, {16'd34987, 16'd7844, 16'd22438, 16'd59653, 16'd57762, 16'd58052, 16'd51725, 16'd14751, 16'd35036, 16'd3798, 16'd6994, 16'd23408, 16'd62101, 16'd38565, 16'd42236, 16'd19333, 16'd12195, 16'd58242, 16'd21663, 16'd850, 16'd6268, 16'd45198, 16'd14981, 16'd17053, 16'd23779, 16'd4345});
	test_expansion(128'h8e1eff63e5c88b5d2076e5f7d26554a0, {16'd20061, 16'd17811, 16'd24926, 16'd30874, 16'd25468, 16'd17147, 16'd46337, 16'd19513, 16'd49139, 16'd54936, 16'd56924, 16'd40264, 16'd1300, 16'd51417, 16'd55612, 16'd42851, 16'd12490, 16'd20209, 16'd21915, 16'd32718, 16'd36053, 16'd43008, 16'd52722, 16'd14704, 16'd57455, 16'd58285});
	test_expansion(128'h29846c6170b0cab5c98461c7295a841c, {16'd65292, 16'd24440, 16'd48460, 16'd36918, 16'd36835, 16'd25776, 16'd35746, 16'd41166, 16'd59648, 16'd33135, 16'd59760, 16'd21141, 16'd3363, 16'd52512, 16'd6204, 16'd32041, 16'd30291, 16'd46637, 16'd64200, 16'd34649, 16'd13451, 16'd52067, 16'd51981, 16'd5545, 16'd28289, 16'd3657});
	test_expansion(128'hd10aa3ad249ba4ef73110ca629560b40, {16'd25705, 16'd33173, 16'd26864, 16'd40436, 16'd62690, 16'd23112, 16'd17123, 16'd48194, 16'd43525, 16'd27240, 16'd7684, 16'd10352, 16'd10622, 16'd31350, 16'd35617, 16'd15414, 16'd51643, 16'd33502, 16'd16585, 16'd63774, 16'd7689, 16'd44537, 16'd46946, 16'd21144, 16'd31935, 16'd6496});
	test_expansion(128'he70fbde20a02884d8a87e80b4fed09f1, {16'd47518, 16'd61215, 16'd30947, 16'd52437, 16'd24198, 16'd59205, 16'd36161, 16'd62061, 16'd32199, 16'd34606, 16'd31089, 16'd29091, 16'd44886, 16'd33534, 16'd48312, 16'd45035, 16'd48146, 16'd6538, 16'd37034, 16'd27700, 16'd15532, 16'd10114, 16'd28478, 16'd58682, 16'd9265, 16'd28997});
	test_expansion(128'h1f1245ff86973e501ac990b93c771299, {16'd59757, 16'd45245, 16'd29714, 16'd59013, 16'd1156, 16'd16694, 16'd25532, 16'd5257, 16'd40301, 16'd20819, 16'd33442, 16'd11483, 16'd48730, 16'd57884, 16'd4812, 16'd20743, 16'd54985, 16'd41692, 16'd21622, 16'd57282, 16'd33548, 16'd13970, 16'd9206, 16'd4846, 16'd60138, 16'd24678});
	test_expansion(128'h767ce8d1a276101eb0399373cf431a9d, {16'd39806, 16'd27023, 16'd188, 16'd22161, 16'd53554, 16'd36494, 16'd28091, 16'd38865, 16'd61, 16'd8525, 16'd114, 16'd59683, 16'd43242, 16'd7886, 16'd23606, 16'd23759, 16'd10443, 16'd18540, 16'd6465, 16'd16631, 16'd6343, 16'd61850, 16'd51368, 16'd19886, 16'd848, 16'd3683});
	test_expansion(128'h3c88de1c8bd7e144acb913024913ffd7, {16'd56308, 16'd52704, 16'd18082, 16'd52574, 16'd24828, 16'd6192, 16'd30778, 16'd26416, 16'd65392, 16'd44256, 16'd59529, 16'd55906, 16'd50990, 16'd45324, 16'd464, 16'd21548, 16'd61733, 16'd53746, 16'd47591, 16'd41477, 16'd52569, 16'd26645, 16'd4478, 16'd38468, 16'd65412, 16'd8921});
	test_expansion(128'h76676f689eb4ef69c27261a34923e7a7, {16'd29479, 16'd45313, 16'd45191, 16'd5706, 16'd17839, 16'd2888, 16'd43224, 16'd10749, 16'd3783, 16'd31271, 16'd45911, 16'd15497, 16'd40397, 16'd58811, 16'd15459, 16'd4253, 16'd32838, 16'd47959, 16'd52424, 16'd57798, 16'd25124, 16'd17654, 16'd19486, 16'd39725, 16'd51214, 16'd53911});
	test_expansion(128'hc18fadfe6fe5842497ae2fc8e16dcd15, {16'd15326, 16'd22285, 16'd4770, 16'd57935, 16'd58995, 16'd33655, 16'd23957, 16'd28356, 16'd12013, 16'd1612, 16'd31743, 16'd40466, 16'd49686, 16'd19575, 16'd20331, 16'd42901, 16'd7490, 16'd6147, 16'd16698, 16'd56542, 16'd8667, 16'd26482, 16'd53631, 16'd59841, 16'd62396, 16'd57537});
	test_expansion(128'hfb4557cd807c143be4c6813efc9aaeda, {16'd62243, 16'd19129, 16'd32736, 16'd30405, 16'd36737, 16'd4134, 16'd33024, 16'd47185, 16'd45754, 16'd62735, 16'd7358, 16'd22285, 16'd65510, 16'd12167, 16'd45129, 16'd34866, 16'd56422, 16'd51338, 16'd42381, 16'd25280, 16'd23157, 16'd60475, 16'd49134, 16'd59439, 16'd1354, 16'd44728});
	test_expansion(128'h6080d9476f0b899bd54c0463edcc48b3, {16'd26619, 16'd23636, 16'd42608, 16'd3246, 16'd27357, 16'd15489, 16'd49999, 16'd61332, 16'd20510, 16'd3885, 16'd60002, 16'd54214, 16'd51338, 16'd8493, 16'd3771, 16'd53767, 16'd56740, 16'd58367, 16'd64714, 16'd19283, 16'd54168, 16'd53738, 16'd41625, 16'd25318, 16'd61472, 16'd50398});
	test_expansion(128'h7c79dc6a3c965a9944d193ea30cd77dd, {16'd63819, 16'd17050, 16'd14523, 16'd47141, 16'd64020, 16'd36496, 16'd8554, 16'd57238, 16'd39936, 16'd32109, 16'd34019, 16'd36446, 16'd23971, 16'd38578, 16'd43570, 16'd514, 16'd2031, 16'd52476, 16'd42099, 16'd36260, 16'd45963, 16'd58368, 16'd50716, 16'd12526, 16'd3344, 16'd41964});
	test_expansion(128'hf37e121a55247600811902c4e99c83f6, {16'd16486, 16'd49769, 16'd2341, 16'd31070, 16'd13198, 16'd59562, 16'd4784, 16'd121, 16'd53293, 16'd40156, 16'd19395, 16'd1983, 16'd56683, 16'd52567, 16'd63278, 16'd12602, 16'd1966, 16'd17602, 16'd3356, 16'd53847, 16'd31691, 16'd11471, 16'd22199, 16'd26683, 16'd22649, 16'd49510});
	test_expansion(128'he7e43225fd582425fd2c2e62c1506898, {16'd12351, 16'd49218, 16'd34786, 16'd22089, 16'd44432, 16'd62397, 16'd828, 16'd63371, 16'd52497, 16'd277, 16'd4756, 16'd30195, 16'd50768, 16'd45085, 16'd1785, 16'd14626, 16'd15143, 16'd51535, 16'd56581, 16'd39258, 16'd20720, 16'd64744, 16'd33159, 16'd40381, 16'd54978, 16'd57349});
	test_expansion(128'h1202fde6d4f00b483aab4c182109405d, {16'd25508, 16'd31783, 16'd28858, 16'd2476, 16'd16984, 16'd64893, 16'd59880, 16'd65527, 16'd14349, 16'd218, 16'd8814, 16'd53475, 16'd21632, 16'd27564, 16'd50068, 16'd38138, 16'd65298, 16'd4416, 16'd27490, 16'd15158, 16'd13394, 16'd192, 16'd8079, 16'd27739, 16'd5192, 16'd32286});
	test_expansion(128'h732739c52d1d38848cc888a06d48dd4c, {16'd33868, 16'd31419, 16'd58346, 16'd54162, 16'd12012, 16'd65361, 16'd21877, 16'd9303, 16'd10769, 16'd53639, 16'd25905, 16'd28320, 16'd7873, 16'd63395, 16'd9730, 16'd40002, 16'd58544, 16'd4818, 16'd30556, 16'd25732, 16'd1430, 16'd10774, 16'd22444, 16'd33961, 16'd39072, 16'd21463});
	test_expansion(128'hf58871e4195a452b89106b7a0ce1d095, {16'd60325, 16'd18959, 16'd22567, 16'd9763, 16'd27418, 16'd48828, 16'd32796, 16'd56840, 16'd58469, 16'd54043, 16'd62208, 16'd47594, 16'd42006, 16'd61575, 16'd6416, 16'd61621, 16'd25514, 16'd5531, 16'd33017, 16'd53501, 16'd40536, 16'd62743, 16'd19509, 16'd44106, 16'd8871, 16'd64689});
	test_expansion(128'h4680e78dd1eef2ce3ff75e73b8d6aa0e, {16'd59542, 16'd19194, 16'd38363, 16'd65152, 16'd7399, 16'd39339, 16'd6788, 16'd43077, 16'd22425, 16'd14327, 16'd26974, 16'd20392, 16'd20776, 16'd34531, 16'd50023, 16'd55154, 16'd25753, 16'd50037, 16'd55906, 16'd20781, 16'd56613, 16'd33273, 16'd36813, 16'd47774, 16'd11673, 16'd64041});
	test_expansion(128'hc93562c745f439b77ffeeb4f99e22908, {16'd59876, 16'd39743, 16'd41217, 16'd50164, 16'd60363, 16'd29836, 16'd58569, 16'd45772, 16'd48120, 16'd37223, 16'd54555, 16'd55789, 16'd6192, 16'd82, 16'd41708, 16'd21540, 16'd25565, 16'd18266, 16'd61737, 16'd8725, 16'd22269, 16'd23125, 16'd49795, 16'd58157, 16'd19846, 16'd1711});
	test_expansion(128'h3f9e44028ce14c90621f2b20e11285dc, {16'd31497, 16'd16776, 16'd33808, 16'd21359, 16'd36195, 16'd10484, 16'd54321, 16'd56100, 16'd11983, 16'd23016, 16'd4720, 16'd27777, 16'd34058, 16'd9868, 16'd23805, 16'd12568, 16'd28556, 16'd15834, 16'd30928, 16'd981, 16'd31567, 16'd61665, 16'd43384, 16'd5399, 16'd63759, 16'd64498});
	test_expansion(128'h8e00f1d766637a65a8e4c567c943f792, {16'd33315, 16'd3107, 16'd59912, 16'd19165, 16'd26825, 16'd4884, 16'd3411, 16'd10395, 16'd11508, 16'd52590, 16'd44669, 16'd35840, 16'd62755, 16'd65517, 16'd48155, 16'd39946, 16'd40106, 16'd65041, 16'd15477, 16'd48665, 16'd49901, 16'd33171, 16'd55123, 16'd60244, 16'd18424, 16'd17904});
	test_expansion(128'h1aade5d2c7abdd2705db80d0c8ba9413, {16'd41085, 16'd42650, 16'd1869, 16'd44634, 16'd48853, 16'd56249, 16'd33012, 16'd64100, 16'd25902, 16'd27316, 16'd41081, 16'd50171, 16'd27219, 16'd45131, 16'd2353, 16'd17883, 16'd16707, 16'd60047, 16'd27799, 16'd57939, 16'd66, 16'd51943, 16'd47947, 16'd48100, 16'd59821, 16'd3191});
	test_expansion(128'ha75be1c0791b335c5631a95121fdfdd8, {16'd63019, 16'd26373, 16'd23069, 16'd53811, 16'd49466, 16'd18131, 16'd23062, 16'd64409, 16'd41729, 16'd43635, 16'd58123, 16'd45434, 16'd42058, 16'd37419, 16'd30405, 16'd60234, 16'd4190, 16'd27757, 16'd47855, 16'd31480, 16'd51196, 16'd28187, 16'd58364, 16'd38335, 16'd29789, 16'd12539});
	test_expansion(128'hcfa5e126ca64d73832b77c6385118af0, {16'd12600, 16'd20898, 16'd16813, 16'd62679, 16'd25074, 16'd3025, 16'd4106, 16'd47977, 16'd15996, 16'd55558, 16'd20596, 16'd14965, 16'd58425, 16'd36366, 16'd19387, 16'd58927, 16'd35512, 16'd57678, 16'd44436, 16'd26944, 16'd19414, 16'd29393, 16'd4402, 16'd23233, 16'd25574, 16'd22962});
	test_expansion(128'h82a6553f581d0a9007d69a195f9ce147, {16'd35993, 16'd23106, 16'd33806, 16'd20684, 16'd5665, 16'd59094, 16'd43101, 16'd5977, 16'd59104, 16'd47555, 16'd4428, 16'd35655, 16'd44732, 16'd53969, 16'd10953, 16'd9513, 16'd51022, 16'd62760, 16'd25166, 16'd1908, 16'd9454, 16'd3250, 16'd35064, 16'd9893, 16'd7706, 16'd30673});
	test_expansion(128'hc6d1652affaf5418d1844ace3d06bb3e, {16'd11, 16'd37301, 16'd47713, 16'd4881, 16'd21410, 16'd33583, 16'd40105, 16'd1925, 16'd47238, 16'd33158, 16'd9568, 16'd25479, 16'd45001, 16'd40015, 16'd60302, 16'd44952, 16'd58314, 16'd21318, 16'd34861, 16'd29725, 16'd26926, 16'd8123, 16'd15244, 16'd3009, 16'd46733, 16'd51355});
	test_expansion(128'h4d775a319595068f04e31bfa48fbd286, {16'd52388, 16'd969, 16'd64451, 16'd31184, 16'd59093, 16'd21349, 16'd5805, 16'd18852, 16'd6193, 16'd21542, 16'd46501, 16'd26772, 16'd54255, 16'd55265, 16'd50066, 16'd6560, 16'd6637, 16'd58370, 16'd21145, 16'd820, 16'd56934, 16'd956, 16'd65169, 16'd8967, 16'd27613, 16'd17730});
	test_expansion(128'h1d928ab7b848d79dfa915ecd64bb900c, {16'd14371, 16'd31480, 16'd7972, 16'd44550, 16'd51349, 16'd44331, 16'd19759, 16'd16975, 16'd1097, 16'd37643, 16'd50082, 16'd20490, 16'd54509, 16'd60548, 16'd19045, 16'd39909, 16'd34218, 16'd62152, 16'd40993, 16'd18320, 16'd4523, 16'd53492, 16'd24247, 16'd32013, 16'd16398, 16'd39323});
	test_expansion(128'h0bd04ff284b2d9b096d4f97dad9ae044, {16'd40951, 16'd14508, 16'd13456, 16'd28948, 16'd25328, 16'd54128, 16'd10208, 16'd28218, 16'd20068, 16'd12829, 16'd9222, 16'd43657, 16'd28377, 16'd27494, 16'd55453, 16'd17788, 16'd38800, 16'd28969, 16'd58662, 16'd43443, 16'd45869, 16'd2663, 16'd53428, 16'd11551, 16'd3282, 16'd19846});
	test_expansion(128'he0810a2a6fd989acd7dc84398a6a47ab, {16'd8877, 16'd6394, 16'd58358, 16'd12417, 16'd7837, 16'd63845, 16'd60296, 16'd49551, 16'd64053, 16'd56681, 16'd15746, 16'd32065, 16'd50798, 16'd29820, 16'd30270, 16'd48801, 16'd7323, 16'd12616, 16'd58020, 16'd19049, 16'd64036, 16'd9599, 16'd45558, 16'd37024, 16'd63219, 16'd33774});
	test_expansion(128'h3efa571cf90baf4b737f607d31a22347, {16'd8866, 16'd341, 16'd12448, 16'd58550, 16'd63922, 16'd42305, 16'd34122, 16'd4529, 16'd7464, 16'd1299, 16'd54231, 16'd20748, 16'd58337, 16'd17187, 16'd8352, 16'd62860, 16'd32957, 16'd4610, 16'd1270, 16'd58861, 16'd38851, 16'd45490, 16'd27040, 16'd64606, 16'd61860, 16'd53140});
	test_expansion(128'h287d08b24b564f3c94d3ffe7e6b1d49c, {16'd56208, 16'd39424, 16'd52462, 16'd40046, 16'd51519, 16'd23227, 16'd64947, 16'd24926, 16'd32063, 16'd64101, 16'd27924, 16'd3820, 16'd45820, 16'd21159, 16'd56053, 16'd23208, 16'd25360, 16'd20639, 16'd29985, 16'd55889, 16'd207, 16'd29050, 16'd6261, 16'd35749, 16'd54427, 16'd38763});
	test_expansion(128'h54c7753b2f1102b7b4e1eb6c1f3c6830, {16'd27636, 16'd38812, 16'd44312, 16'd40625, 16'd7168, 16'd18881, 16'd34914, 16'd43601, 16'd55911, 16'd21047, 16'd61266, 16'd5762, 16'd54062, 16'd30153, 16'd16601, 16'd30069, 16'd37013, 16'd30836, 16'd65083, 16'd33713, 16'd49861, 16'd54987, 16'd30429, 16'd51331, 16'd32606, 16'd64122});
	test_expansion(128'hf381f2494090eaf9699ab4da064afbf4, {16'd54582, 16'd1034, 16'd57762, 16'd56387, 16'd29128, 16'd5951, 16'd53318, 16'd8111, 16'd4602, 16'd54452, 16'd28677, 16'd7482, 16'd25476, 16'd7147, 16'd47632, 16'd5182, 16'd15550, 16'd61314, 16'd13276, 16'd16844, 16'd33593, 16'd10106, 16'd8192, 16'd51225, 16'd35639, 16'd49886});
	test_expansion(128'hb5bf1bc1dd3402645a74f495436bf177, {16'd31429, 16'd3213, 16'd50113, 16'd10057, 16'd20731, 16'd37507, 16'd3677, 16'd25599, 16'd59274, 16'd10475, 16'd7870, 16'd38082, 16'd19320, 16'd36411, 16'd26311, 16'd65239, 16'd34603, 16'd50839, 16'd13026, 16'd49599, 16'd17307, 16'd36296, 16'd16630, 16'd34691, 16'd50744, 16'd4224});
	test_expansion(128'hed084f853da7920199f1411155ca7eb6, {16'd21931, 16'd16050, 16'd31, 16'd33179, 16'd16601, 16'd58983, 16'd43131, 16'd7743, 16'd53424, 16'd13185, 16'd53169, 16'd2605, 16'd42438, 16'd37105, 16'd28450, 16'd895, 16'd23659, 16'd48738, 16'd37073, 16'd11657, 16'd24248, 16'd9404, 16'd4325, 16'd15641, 16'd15317, 16'd45513});
	test_expansion(128'h45be98097c8705de421408f79dfd5b75, {16'd38927, 16'd6827, 16'd33244, 16'd22221, 16'd45783, 16'd11195, 16'd17376, 16'd29652, 16'd3343, 16'd33366, 16'd10686, 16'd19632, 16'd60031, 16'd58416, 16'd33590, 16'd63566, 16'd38819, 16'd4712, 16'd41580, 16'd524, 16'd11575, 16'd22758, 16'd38433, 16'd11033, 16'd26747, 16'd23947});
	test_expansion(128'he5275acb5d7bc49417f66f4e06cdc48d, {16'd51537, 16'd8499, 16'd34354, 16'd15421, 16'd54007, 16'd3083, 16'd26907, 16'd59461, 16'd23308, 16'd45317, 16'd10105, 16'd35298, 16'd50079, 16'd23288, 16'd45865, 16'd54782, 16'd54465, 16'd15883, 16'd4694, 16'd45881, 16'd14710, 16'd30961, 16'd53104, 16'd11489, 16'd31256, 16'd55761});
	test_expansion(128'hfb567ba44c83e8972fafd4e6a45d57e8, {16'd34695, 16'd35568, 16'd49367, 16'd37456, 16'd26052, 16'd17813, 16'd14793, 16'd65372, 16'd56616, 16'd36474, 16'd32778, 16'd65149, 16'd35331, 16'd40646, 16'd64632, 16'd20100, 16'd37342, 16'd46166, 16'd55697, 16'd25633, 16'd40332, 16'd53785, 16'd38900, 16'd57262, 16'd39511, 16'd47065});
	test_expansion(128'h3c5b44b73af29114ad68e5b7aafd5949, {16'd25937, 16'd30011, 16'd21638, 16'd61857, 16'd65433, 16'd46499, 16'd30505, 16'd50511, 16'd21813, 16'd22258, 16'd13285, 16'd32225, 16'd3485, 16'd30546, 16'd35899, 16'd47126, 16'd32061, 16'd6537, 16'd58309, 16'd59289, 16'd37183, 16'd60320, 16'd30165, 16'd18019, 16'd9679, 16'd1345});
	test_expansion(128'h1fb2615f677ad221e0d5de01e73734c9, {16'd54347, 16'd35343, 16'd45668, 16'd39604, 16'd18264, 16'd42255, 16'd60805, 16'd32225, 16'd54004, 16'd52174, 16'd22767, 16'd55753, 16'd36974, 16'd22096, 16'd43683, 16'd3813, 16'd8141, 16'd40810, 16'd51443, 16'd31856, 16'd59166, 16'd47721, 16'd35479, 16'd8324, 16'd63054, 16'd36195});
	test_expansion(128'he2cbc781524b227a5edba9c47397ceab, {16'd394, 16'd6900, 16'd5623, 16'd36874, 16'd47730, 16'd45483, 16'd3585, 16'd63236, 16'd13230, 16'd45607, 16'd45525, 16'd33417, 16'd59339, 16'd38991, 16'd59631, 16'd25536, 16'd34551, 16'd8503, 16'd1878, 16'd6638, 16'd47966, 16'd63883, 16'd39577, 16'd52170, 16'd43845, 16'd42794});
	test_expansion(128'he1a2a5515f0eb4d050982bdff4819506, {16'd14006, 16'd2085, 16'd15923, 16'd20915, 16'd51826, 16'd61756, 16'd24719, 16'd4785, 16'd55548, 16'd29630, 16'd19100, 16'd49908, 16'd38421, 16'd45848, 16'd46069, 16'd49248, 16'd25947, 16'd36956, 16'd65371, 16'd42257, 16'd29696, 16'd47452, 16'd14134, 16'd18212, 16'd18896, 16'd45112});
	test_expansion(128'h0ee87d140984a8e32a6d0c85c013d670, {16'd64527, 16'd33319, 16'd9245, 16'd40759, 16'd14180, 16'd32111, 16'd27092, 16'd22786, 16'd58273, 16'd52839, 16'd61271, 16'd7794, 16'd12875, 16'd41245, 16'd22775, 16'd15612, 16'd52529, 16'd61673, 16'd41678, 16'd36442, 16'd1037, 16'd18391, 16'd32742, 16'd33928, 16'd32216, 16'd47870});
	test_expansion(128'habb923ecee03d63a2dc13823a0ea98d3, {16'd28976, 16'd27733, 16'd1636, 16'd19579, 16'd35654, 16'd64095, 16'd23797, 16'd29015, 16'd23062, 16'd63690, 16'd53377, 16'd15886, 16'd41276, 16'd29586, 16'd30071, 16'd48013, 16'd59709, 16'd1543, 16'd13327, 16'd26209, 16'd37734, 16'd27856, 16'd6953, 16'd21653, 16'd34226, 16'd37424});
	test_expansion(128'hacda2bcb2d9c815bff8ec51b14a8744a, {16'd40288, 16'd14678, 16'd21887, 16'd22541, 16'd23924, 16'd41553, 16'd49131, 16'd10786, 16'd25352, 16'd58727, 16'd61722, 16'd39657, 16'd11813, 16'd49817, 16'd61570, 16'd27884, 16'd22512, 16'd63850, 16'd39645, 16'd45672, 16'd30759, 16'd48692, 16'd26062, 16'd29838, 16'd45113, 16'd46428});
	test_expansion(128'h967b6a6030f2bd041c749f124247543f, {16'd40608, 16'd45974, 16'd45655, 16'd6408, 16'd7370, 16'd2045, 16'd28791, 16'd14946, 16'd61414, 16'd16089, 16'd36502, 16'd15526, 16'd47286, 16'd30324, 16'd42150, 16'd58378, 16'd18632, 16'd41810, 16'd9658, 16'd50764, 16'd53045, 16'd20408, 16'd30847, 16'd46576, 16'd60474, 16'd24997});
	test_expansion(128'h983fce2aa244ea5c1cccca6acd3f2812, {16'd57572, 16'd43041, 16'd55657, 16'd45606, 16'd12300, 16'd59423, 16'd47999, 16'd39051, 16'd60123, 16'd40657, 16'd42922, 16'd51388, 16'd1120, 16'd60207, 16'd48312, 16'd23952, 16'd10554, 16'd8346, 16'd64498, 16'd19097, 16'd18207, 16'd31256, 16'd55086, 16'd36341, 16'd4104, 16'd53971});
	test_expansion(128'hfead1d5254b8c5debf9115da1dc35007, {16'd21064, 16'd12439, 16'd38453, 16'd10330, 16'd31437, 16'd25978, 16'd37916, 16'd36520, 16'd14913, 16'd32372, 16'd14925, 16'd43387, 16'd37600, 16'd24497, 16'd22944, 16'd42849, 16'd17050, 16'd65147, 16'd28458, 16'd14611, 16'd45623, 16'd27237, 16'd49676, 16'd15059, 16'd60176, 16'd5072});
	test_expansion(128'h34d0371b0584ff2ca0dc2dc8ebe44f2f, {16'd45665, 16'd26919, 16'd15725, 16'd36983, 16'd14515, 16'd29522, 16'd52873, 16'd17159, 16'd60326, 16'd31124, 16'd12640, 16'd62053, 16'd54722, 16'd3769, 16'd6100, 16'd22940, 16'd52909, 16'd1098, 16'd10269, 16'd6711, 16'd42057, 16'd1650, 16'd1623, 16'd56042, 16'd19244, 16'd39419});
	test_expansion(128'h5223a59f7e773fc50cdd6a26af2f1c84, {16'd21823, 16'd38222, 16'd58234, 16'd4405, 16'd14446, 16'd28939, 16'd62839, 16'd42969, 16'd55767, 16'd8672, 16'd17946, 16'd63746, 16'd26028, 16'd60592, 16'd20113, 16'd23885, 16'd24308, 16'd4883, 16'd44635, 16'd22322, 16'd56253, 16'd51358, 16'd38281, 16'd36823, 16'd15276, 16'd60557});
	test_expansion(128'h987e0792aae1deddcc0b389ffa9d4127, {16'd30405, 16'd28319, 16'd11192, 16'd62861, 16'd52579, 16'd24435, 16'd43431, 16'd9810, 16'd13541, 16'd58454, 16'd56195, 16'd46573, 16'd10368, 16'd1721, 16'd17352, 16'd57615, 16'd8191, 16'd13024, 16'd18641, 16'd62806, 16'd47288, 16'd53476, 16'd30846, 16'd8821, 16'd56975, 16'd11784});
	test_expansion(128'h34f4c0a9cad1f0fbef1d167be310eb55, {16'd52065, 16'd35400, 16'd44337, 16'd45611, 16'd8044, 16'd10240, 16'd31475, 16'd29661, 16'd9816, 16'd44224, 16'd41567, 16'd19255, 16'd20036, 16'd39908, 16'd49103, 16'd42373, 16'd23500, 16'd21917, 16'd35653, 16'd25478, 16'd37225, 16'd38874, 16'd27569, 16'd34707, 16'd63174, 16'd47886});
	test_expansion(128'hef4a8a001769a49b4bfa0eed927c0d0d, {16'd55676, 16'd35077, 16'd42364, 16'd31588, 16'd5444, 16'd65022, 16'd59661, 16'd30236, 16'd65035, 16'd53571, 16'd48226, 16'd59636, 16'd57742, 16'd6609, 16'd6070, 16'd3975, 16'd54896, 16'd44069, 16'd43323, 16'd3246, 16'd23690, 16'd6820, 16'd50169, 16'd20448, 16'd24807, 16'd21403});
	test_expansion(128'hcca556ada5162a1ef3abdfe521cef18c, {16'd49152, 16'd39484, 16'd61246, 16'd54928, 16'd50216, 16'd22708, 16'd46226, 16'd46912, 16'd16312, 16'd26005, 16'd37025, 16'd6528, 16'd8082, 16'd49998, 16'd52360, 16'd1559, 16'd41524, 16'd50670, 16'd28019, 16'd7788, 16'd64571, 16'd38094, 16'd58872, 16'd24388, 16'd19126, 16'd28330});
	test_expansion(128'h3460b1274826a61bedf8dc890717b73a, {16'd30849, 16'd61299, 16'd57876, 16'd48250, 16'd64542, 16'd58213, 16'd63151, 16'd12841, 16'd8149, 16'd9259, 16'd48061, 16'd7155, 16'd2567, 16'd12936, 16'd19094, 16'd37158, 16'd16811, 16'd3377, 16'd45103, 16'd56985, 16'd43397, 16'd49982, 16'd39848, 16'd55236, 16'd59715, 16'd17097});
	test_expansion(128'hf560e87f1d6f38a9e25a9cf365f422cc, {16'd14513, 16'd65026, 16'd33067, 16'd62675, 16'd48111, 16'd41021, 16'd51878, 16'd51745, 16'd16938, 16'd48364, 16'd42017, 16'd60503, 16'd22858, 16'd48740, 16'd61321, 16'd25850, 16'd8763, 16'd61907, 16'd63624, 16'd26772, 16'd64219, 16'd10804, 16'd54205, 16'd25907, 16'd33895, 16'd4565});
	test_expansion(128'h1ca2ce75540931a592a95dfe2b06e13f, {16'd19852, 16'd9297, 16'd33627, 16'd57079, 16'd51420, 16'd33505, 16'd61349, 16'd5671, 16'd30761, 16'd59620, 16'd3845, 16'd59234, 16'd24709, 16'd43728, 16'd43945, 16'd64517, 16'd9010, 16'd21777, 16'd26648, 16'd56147, 16'd16111, 16'd21481, 16'd19722, 16'd27241, 16'd28221, 16'd13454});
	test_expansion(128'h3dea69771af2378aad4cff53a7ca0f43, {16'd29210, 16'd42014, 16'd15758, 16'd24917, 16'd5039, 16'd56503, 16'd39142, 16'd22287, 16'd58169, 16'd0, 16'd36206, 16'd347, 16'd53817, 16'd25206, 16'd46479, 16'd34678, 16'd62036, 16'd65498, 16'd33047, 16'd49230, 16'd25466, 16'd23117, 16'd53220, 16'd23999, 16'd3649, 16'd35509});
	test_expansion(128'h7dd06b37b6465984220f17c59ab943cb, {16'd10252, 16'd34145, 16'd35540, 16'd9714, 16'd47075, 16'd64807, 16'd21819, 16'd54833, 16'd62454, 16'd26078, 16'd13523, 16'd10304, 16'd48663, 16'd2900, 16'd35885, 16'd41390, 16'd22802, 16'd21017, 16'd33088, 16'd64484, 16'd663, 16'd10629, 16'd3711, 16'd28415, 16'd24630, 16'd55950});
	test_expansion(128'h3616654ed6ad560079403ed90413fd12, {16'd63241, 16'd58150, 16'd21571, 16'd45011, 16'd17827, 16'd18044, 16'd48754, 16'd3999, 16'd34783, 16'd37406, 16'd64466, 16'd45089, 16'd26573, 16'd4613, 16'd55655, 16'd29030, 16'd58488, 16'd24676, 16'd5441, 16'd6853, 16'd34543, 16'd25005, 16'd36870, 16'd29008, 16'd6460, 16'd27087});
	test_expansion(128'h3bfc7a9cc53f6162768f20ac522a5480, {16'd59958, 16'd2565, 16'd16987, 16'd43035, 16'd61585, 16'd57945, 16'd62896, 16'd3088, 16'd468, 16'd62886, 16'd15705, 16'd61413, 16'd59699, 16'd31087, 16'd5552, 16'd25694, 16'd42699, 16'd54304, 16'd54250, 16'd8252, 16'd14745, 16'd19500, 16'd47685, 16'd42839, 16'd55974, 16'd55521});
	test_expansion(128'hab65db49807b0998f3b23914930fc734, {16'd43162, 16'd63007, 16'd9900, 16'd56285, 16'd891, 16'd4950, 16'd14657, 16'd23932, 16'd8044, 16'd43361, 16'd39095, 16'd28113, 16'd8553, 16'd28920, 16'd15505, 16'd22953, 16'd28594, 16'd63573, 16'd3287, 16'd60155, 16'd34935, 16'd5910, 16'd954, 16'd38599, 16'd32314, 16'd28918});
	test_expansion(128'h0a81a6c0fcd7ea9a05843764bb9f09fc, {16'd47619, 16'd12657, 16'd35469, 16'd31728, 16'd21643, 16'd13492, 16'd26000, 16'd24595, 16'd54847, 16'd16742, 16'd34752, 16'd47373, 16'd43210, 16'd4525, 16'd39082, 16'd62035, 16'd10454, 16'd34230, 16'd44828, 16'd5696, 16'd9362, 16'd12791, 16'd59634, 16'd1469, 16'd59983, 16'd6326});
	test_expansion(128'hd59c6e80bb8e20eacf462cf8e7ebd5f5, {16'd49438, 16'd37330, 16'd5492, 16'd5185, 16'd4647, 16'd49799, 16'd39902, 16'd51661, 16'd64785, 16'd24686, 16'd18326, 16'd34048, 16'd35368, 16'd31671, 16'd55883, 16'd32382, 16'd13413, 16'd57645, 16'd26443, 16'd55675, 16'd1856, 16'd65482, 16'd54836, 16'd53039, 16'd51579, 16'd3711});
	test_expansion(128'h5a0c456970cb787a2c59a7a29d97ea85, {16'd37169, 16'd61265, 16'd64150, 16'd18782, 16'd36016, 16'd11529, 16'd45701, 16'd37360, 16'd64850, 16'd25405, 16'd23235, 16'd63399, 16'd63813, 16'd15375, 16'd47924, 16'd28589, 16'd65516, 16'd58798, 16'd59084, 16'd20356, 16'd28826, 16'd61105, 16'd6509, 16'd13602, 16'd11033, 16'd25493});
	test_expansion(128'h268e818841bb07329c0515d9aec01766, {16'd13029, 16'd45174, 16'd11160, 16'd9016, 16'd47155, 16'd31109, 16'd2926, 16'd36979, 16'd4750, 16'd52469, 16'd33165, 16'd60804, 16'd38468, 16'd14292, 16'd46370, 16'd56859, 16'd6123, 16'd53193, 16'd22876, 16'd38423, 16'd9841, 16'd34338, 16'd33599, 16'd7236, 16'd43321, 16'd23166});
	test_expansion(128'hbc8bda7e9b2cc413a08e2ed4d6124427, {16'd21788, 16'd13767, 16'd53774, 16'd59101, 16'd24684, 16'd3371, 16'd21481, 16'd38865, 16'd4434, 16'd51617, 16'd22658, 16'd4600, 16'd30312, 16'd38732, 16'd27313, 16'd50526, 16'd46773, 16'd6632, 16'd27079, 16'd56315, 16'd40552, 16'd29714, 16'd17564, 16'd56263, 16'd38944, 16'd33928});
	test_expansion(128'hb258cb4208d8dd193bfadfa47da1d0d8, {16'd26206, 16'd38693, 16'd584, 16'd44807, 16'd529, 16'd14269, 16'd25062, 16'd24741, 16'd22544, 16'd59577, 16'd28066, 16'd64475, 16'd11760, 16'd143, 16'd20510, 16'd10374, 16'd57942, 16'd37287, 16'd11038, 16'd39704, 16'd56093, 16'd40981, 16'd19763, 16'd63913, 16'd46855, 16'd61868});
	test_expansion(128'hfb053e3f9b6bc7f9b9cea569b9df5f82, {16'd52943, 16'd47881, 16'd64823, 16'd64423, 16'd41069, 16'd27336, 16'd45544, 16'd10222, 16'd24335, 16'd50779, 16'd17665, 16'd20653, 16'd26728, 16'd43202, 16'd26898, 16'd48440, 16'd31244, 16'd14612, 16'd1937, 16'd59244, 16'd48464, 16'd11144, 16'd62118, 16'd39530, 16'd53334, 16'd56176});
	test_expansion(128'h3acbd423293091f8086daad10073c970, {16'd56689, 16'd46552, 16'd63090, 16'd55256, 16'd53960, 16'd10552, 16'd54765, 16'd63985, 16'd33872, 16'd11153, 16'd10910, 16'd7001, 16'd62978, 16'd2351, 16'd34937, 16'd8690, 16'd8165, 16'd42312, 16'd60770, 16'd24317, 16'd32294, 16'd3104, 16'd39723, 16'd39486, 16'd9459, 16'd19500});
	test_expansion(128'h94ff5913c76e428fb554c4cca8991f15, {16'd12374, 16'd24688, 16'd46751, 16'd62562, 16'd46274, 16'd9162, 16'd40192, 16'd27361, 16'd18067, 16'd32820, 16'd11227, 16'd26845, 16'd16986, 16'd47571, 16'd40174, 16'd31989, 16'd15670, 16'd42686, 16'd30230, 16'd54033, 16'd1687, 16'd31356, 16'd18853, 16'd35022, 16'd52359, 16'd19777});
	test_expansion(128'h0c6d2fa5bfc5bdb74a627b129ebd6eca, {16'd43654, 16'd13403, 16'd17513, 16'd21189, 16'd55784, 16'd38909, 16'd34793, 16'd1825, 16'd5015, 16'd62219, 16'd31527, 16'd29900, 16'd42489, 16'd34769, 16'd2372, 16'd37144, 16'd23403, 16'd63763, 16'd55056, 16'd65070, 16'd44829, 16'd41328, 16'd50092, 16'd48277, 16'd59295, 16'd40674});
	test_expansion(128'h7221a0ab51df0c0b39d308e9e87f2757, {16'd40812, 16'd31365, 16'd21997, 16'd11609, 16'd27868, 16'd30059, 16'd63627, 16'd55696, 16'd36708, 16'd48656, 16'd42813, 16'd46653, 16'd6482, 16'd36967, 16'd19152, 16'd52043, 16'd10154, 16'd8768, 16'd52435, 16'd4260, 16'd26492, 16'd55736, 16'd20199, 16'd26168, 16'd30804, 16'd16132});
	test_expansion(128'h84b0872828c83f294159ec084b0b52b2, {16'd9370, 16'd5931, 16'd19269, 16'd34781, 16'd34072, 16'd7137, 16'd35007, 16'd20229, 16'd14956, 16'd44891, 16'd12569, 16'd41766, 16'd47992, 16'd52752, 16'd18166, 16'd65150, 16'd18386, 16'd5300, 16'd57819, 16'd3655, 16'd49711, 16'd51588, 16'd6567, 16'd41799, 16'd18082, 16'd37030});
	test_expansion(128'h501cf2458edcb7e2f0e7ffcac705978a, {16'd59487, 16'd19288, 16'd46401, 16'd26499, 16'd28878, 16'd52229, 16'd29537, 16'd48703, 16'd50656, 16'd35518, 16'd14628, 16'd6382, 16'd32583, 16'd4326, 16'd12294, 16'd65215, 16'd27290, 16'd57230, 16'd2395, 16'd19790, 16'd29239, 16'd39528, 16'd54206, 16'd14968, 16'd11215, 16'd57464});
	test_expansion(128'h30f6da4b39dcdfddef8e5fbef84da41a, {16'd22636, 16'd43232, 16'd65425, 16'd19507, 16'd58587, 16'd43723, 16'd21395, 16'd58747, 16'd44880, 16'd25559, 16'd19193, 16'd54209, 16'd24933, 16'd53309, 16'd51472, 16'd63900, 16'd42477, 16'd264, 16'd64273, 16'd59446, 16'd10385, 16'd48200, 16'd28235, 16'd49310, 16'd54355, 16'd23289});
	test_expansion(128'h9efb61c7d2f207dfc811379fc343e857, {16'd19790, 16'd25348, 16'd1802, 16'd35505, 16'd39087, 16'd51567, 16'd17140, 16'd31756, 16'd63274, 16'd43920, 16'd1802, 16'd31052, 16'd26656, 16'd791, 16'd1138, 16'd42559, 16'd40166, 16'd3710, 16'd44871, 16'd58757, 16'd52717, 16'd5894, 16'd44077, 16'd13316, 16'd12112, 16'd36353});
	test_expansion(128'h38d5bfee52506e610f4ebc6d3fbd1680, {16'd7488, 16'd1618, 16'd64165, 16'd6204, 16'd51475, 16'd43238, 16'd23365, 16'd15332, 16'd55583, 16'd61707, 16'd49464, 16'd17258, 16'd32508, 16'd2436, 16'd54157, 16'd12931, 16'd1653, 16'd42158, 16'd43086, 16'd11800, 16'd23499, 16'd51576, 16'd23398, 16'd35362, 16'd1782, 16'd26817});
	test_expansion(128'hb56385e11bc4e8803b27f0ce39066c68, {16'd22599, 16'd40131, 16'd44884, 16'd15000, 16'd833, 16'd60922, 16'd59612, 16'd40187, 16'd16095, 16'd6034, 16'd24373, 16'd7321, 16'd49996, 16'd18306, 16'd24239, 16'd47148, 16'd48705, 16'd3414, 16'd9839, 16'd4977, 16'd18719, 16'd61592, 16'd57061, 16'd14587, 16'd9020, 16'd39512});
	test_expansion(128'h22e450b17bcdb2c9a19b9840c93e88e1, {16'd44646, 16'd31098, 16'd30598, 16'd21093, 16'd23698, 16'd16458, 16'd48201, 16'd6410, 16'd43055, 16'd24494, 16'd27241, 16'd13767, 16'd54011, 16'd42701, 16'd55138, 16'd55980, 16'd52664, 16'd56447, 16'd5130, 16'd1362, 16'd18918, 16'd48142, 16'd7286, 16'd8692, 16'd3742, 16'd12302});
	test_expansion(128'h9c8586bb1f3a1be8f4379125f6d71479, {16'd16311, 16'd3473, 16'd21592, 16'd59099, 16'd13302, 16'd65445, 16'd24632, 16'd58515, 16'd30294, 16'd10201, 16'd45491, 16'd42168, 16'd8886, 16'd36199, 16'd25158, 16'd10415, 16'd5952, 16'd26062, 16'd23505, 16'd2739, 16'd44985, 16'd54885, 16'd44604, 16'd23513, 16'd8231, 16'd9487});
	test_expansion(128'h5d9138d9556d953cc8a89247b095c5d2, {16'd51968, 16'd38503, 16'd17220, 16'd51288, 16'd43234, 16'd43721, 16'd57123, 16'd16549, 16'd60782, 16'd19685, 16'd37508, 16'd51480, 16'd25391, 16'd16095, 16'd30570, 16'd36902, 16'd925, 16'd44069, 16'd13097, 16'd46933, 16'd56238, 16'd58825, 16'd108, 16'd19656, 16'd54674, 16'd2997});
	test_expansion(128'h8cf412d091324af165d3c1c9d6a11ebe, {16'd10525, 16'd59868, 16'd44864, 16'd29440, 16'd53061, 16'd65449, 16'd58227, 16'd30648, 16'd31223, 16'd49333, 16'd54172, 16'd23382, 16'd54565, 16'd6076, 16'd31259, 16'd62285, 16'd19818, 16'd56298, 16'd64113, 16'd11902, 16'd3693, 16'd8533, 16'd56151, 16'd27190, 16'd44995, 16'd50766});
	test_expansion(128'h046b000a97c1d237846db5ec702b44bb, {16'd11659, 16'd11884, 16'd58484, 16'd42341, 16'd35043, 16'd63220, 16'd58343, 16'd55641, 16'd17438, 16'd63583, 16'd34807, 16'd43240, 16'd51315, 16'd42514, 16'd54586, 16'd63780, 16'd25963, 16'd1530, 16'd64945, 16'd20763, 16'd19865, 16'd3784, 16'd43623, 16'd45930, 16'd24837, 16'd23877});
	test_expansion(128'h3f3594e449312c79d435686c45c7a116, {16'd32871, 16'd51778, 16'd38354, 16'd33147, 16'd7588, 16'd7671, 16'd60452, 16'd62744, 16'd41684, 16'd4910, 16'd23428, 16'd52157, 16'd58871, 16'd22434, 16'd34977, 16'd26470, 16'd48206, 16'd62912, 16'd30979, 16'd26303, 16'd219, 16'd49932, 16'd42772, 16'd6873, 16'd55601, 16'd28965});
	test_expansion(128'h823f9e68cc82b59e07a8fcd4b5694c29, {16'd54805, 16'd59416, 16'd62734, 16'd26959, 16'd54016, 16'd21814, 16'd58942, 16'd15017, 16'd47323, 16'd8724, 16'd43722, 16'd21238, 16'd50854, 16'd36758, 16'd29615, 16'd63692, 16'd42965, 16'd38720, 16'd44796, 16'd22678, 16'd60006, 16'd12238, 16'd50148, 16'd48623, 16'd63658, 16'd27369});
	test_expansion(128'h1dc087d1d21898c38bb777cb3dae317a, {16'd39972, 16'd28280, 16'd21297, 16'd27317, 16'd19917, 16'd53582, 16'd13617, 16'd18712, 16'd41482, 16'd62205, 16'd33169, 16'd55528, 16'd47278, 16'd7026, 16'd2307, 16'd15903, 16'd46580, 16'd14579, 16'd18392, 16'd12285, 16'd49829, 16'd22764, 16'd57185, 16'd59846, 16'd61419, 16'd22907});
	test_expansion(128'hdc58106aef8ba965ee09e2833b6fc3e2, {16'd36587, 16'd11388, 16'd28519, 16'd37061, 16'd40648, 16'd54865, 16'd56174, 16'd48148, 16'd33116, 16'd20716, 16'd21009, 16'd12741, 16'd37265, 16'd59835, 16'd59704, 16'd17964, 16'd24774, 16'd30259, 16'd29677, 16'd49202, 16'd4797, 16'd9833, 16'd8288, 16'd14170, 16'd14474, 16'd56871});
	test_expansion(128'h07b48f136b1a72ba4bf5c9a7c22ded6e, {16'd61349, 16'd59224, 16'd46819, 16'd34700, 16'd54986, 16'd56570, 16'd65159, 16'd21835, 16'd49207, 16'd22337, 16'd43622, 16'd15668, 16'd46384, 16'd34287, 16'd14034, 16'd64958, 16'd4221, 16'd17481, 16'd40089, 16'd35596, 16'd18255, 16'd32108, 16'd34538, 16'd2662, 16'd48798, 16'd11535});
	test_expansion(128'h45858f64ecb273e3e36d9aad2c0174ea, {16'd13671, 16'd18922, 16'd3145, 16'd4382, 16'd704, 16'd61864, 16'd3975, 16'd25263, 16'd35714, 16'd46892, 16'd26151, 16'd16714, 16'd34510, 16'd31709, 16'd19382, 16'd16782, 16'd10222, 16'd22669, 16'd16938, 16'd58768, 16'd22196, 16'd51456, 16'd11686, 16'd24235, 16'd62275, 16'd52833});
	test_expansion(128'h8c0dd02fabc364a227bfbee254b36731, {16'd6732, 16'd6580, 16'd57110, 16'd17558, 16'd55383, 16'd51896, 16'd43501, 16'd407, 16'd41103, 16'd56378, 16'd50951, 16'd35336, 16'd16737, 16'd19768, 16'd25274, 16'd14495, 16'd232, 16'd11853, 16'd21466, 16'd44350, 16'd18784, 16'd1242, 16'd8613, 16'd30751, 16'd5432, 16'd26942});
	test_expansion(128'h58eef56cac5f0ff1a772f1e7a3511e91, {16'd62289, 16'd44830, 16'd10019, 16'd45091, 16'd20026, 16'd5412, 16'd29776, 16'd664, 16'd1608, 16'd33842, 16'd51953, 16'd1872, 16'd10831, 16'd12150, 16'd52072, 16'd21453, 16'd442, 16'd4563, 16'd61539, 16'd3824, 16'd58586, 16'd7147, 16'd32826, 16'd40069, 16'd44141, 16'd61164});
	test_expansion(128'h17b0a8e7f830bef0b5557625ba486ee4, {16'd63871, 16'd30672, 16'd45662, 16'd11299, 16'd38155, 16'd9220, 16'd1899, 16'd9574, 16'd11794, 16'd52332, 16'd353, 16'd6234, 16'd38730, 16'd62258, 16'd41276, 16'd51179, 16'd28182, 16'd13832, 16'd10925, 16'd4586, 16'd35107, 16'd50669, 16'd47713, 16'd55445, 16'd1542, 16'd14606});
	test_expansion(128'h6394f2e0da1b871b5cffcd8936905884, {16'd19224, 16'd45603, 16'd38683, 16'd59449, 16'd44099, 16'd57387, 16'd8766, 16'd24353, 16'd27996, 16'd5593, 16'd22360, 16'd23067, 16'd23641, 16'd30679, 16'd42514, 16'd23974, 16'd25715, 16'd36647, 16'd37751, 16'd7628, 16'd57279, 16'd5585, 16'd55702, 16'd37765, 16'd7904, 16'd32827});
	test_expansion(128'hd0e14cc2421de52bebe18ac08ec1bfc6, {16'd10685, 16'd1553, 16'd13892, 16'd44006, 16'd54251, 16'd11452, 16'd36487, 16'd9187, 16'd54298, 16'd41985, 16'd39680, 16'd40560, 16'd21842, 16'd52562, 16'd29781, 16'd23994, 16'd60419, 16'd51895, 16'd49908, 16'd62762, 16'd29084, 16'd30547, 16'd38596, 16'd10515, 16'd44591, 16'd58103});
	test_expansion(128'h678610ec8d64b75d2bdc304c6c0d7dd9, {16'd7053, 16'd18059, 16'd53972, 16'd4287, 16'd16741, 16'd49099, 16'd387, 16'd46965, 16'd11582, 16'd33980, 16'd1075, 16'd65116, 16'd9490, 16'd48110, 16'd36355, 16'd26729, 16'd22104, 16'd4957, 16'd19985, 16'd16509, 16'd14374, 16'd4140, 16'd64015, 16'd58634, 16'd50332, 16'd7363});
	test_expansion(128'h779405ce8cbc86a6acc66aa238d75bd9, {16'd18618, 16'd10460, 16'd4113, 16'd59310, 16'd17259, 16'd20237, 16'd59911, 16'd27494, 16'd2394, 16'd57638, 16'd30481, 16'd9763, 16'd14664, 16'd32665, 16'd46470, 16'd54842, 16'd55267, 16'd16548, 16'd62097, 16'd44025, 16'd27747, 16'd12054, 16'd55487, 16'd14736, 16'd4938, 16'd28199});
	test_expansion(128'ha3cc56210930210ba459ed970fb82b24, {16'd5797, 16'd32493, 16'd7386, 16'd13227, 16'd59203, 16'd25726, 16'd51008, 16'd22833, 16'd59318, 16'd34752, 16'd25230, 16'd9610, 16'd51058, 16'd19736, 16'd58827, 16'd34431, 16'd19755, 16'd25238, 16'd3271, 16'd31383, 16'd8242, 16'd37579, 16'd7416, 16'd28954, 16'd62841, 16'd57980});
	test_expansion(128'h2294a37a3235bc53564485fb77324114, {16'd57693, 16'd55127, 16'd64900, 16'd63621, 16'd5671, 16'd16769, 16'd6952, 16'd12363, 16'd15604, 16'd20990, 16'd55213, 16'd57097, 16'd48235, 16'd3338, 16'd21325, 16'd9294, 16'd33843, 16'd9615, 16'd36161, 16'd2299, 16'd16026, 16'd1740, 16'd7763, 16'd15281, 16'd37905, 16'd25885});
	test_expansion(128'h9b3c7cb2ff9bd55a30696aa30596ec5d, {16'd52370, 16'd24751, 16'd55748, 16'd13843, 16'd17742, 16'd45135, 16'd35914, 16'd58051, 16'd37375, 16'd36498, 16'd7314, 16'd29365, 16'd48495, 16'd64030, 16'd42262, 16'd45818, 16'd50083, 16'd28178, 16'd15939, 16'd445, 16'd15075, 16'd34392, 16'd9749, 16'd35528, 16'd61855, 16'd52024});
	test_expansion(128'h49e490f22b29be715a02bd7e80553caf, {16'd12486, 16'd4268, 16'd39228, 16'd1300, 16'd23438, 16'd60493, 16'd17603, 16'd36231, 16'd54608, 16'd46318, 16'd3379, 16'd14202, 16'd10618, 16'd37006, 16'd3556, 16'd15357, 16'd3685, 16'd44118, 16'd61326, 16'd38108, 16'd38679, 16'd11425, 16'd39236, 16'd55264, 16'd55760, 16'd57906});
	test_expansion(128'hb2a75a2a929417913c290459709a99eb, {16'd42415, 16'd33558, 16'd44822, 16'd44396, 16'd45144, 16'd3919, 16'd43931, 16'd11357, 16'd33550, 16'd26934, 16'd2046, 16'd11885, 16'd30464, 16'd55533, 16'd32924, 16'd45417, 16'd36169, 16'd2779, 16'd12821, 16'd17367, 16'd34699, 16'd29151, 16'd55115, 16'd30920, 16'd34855, 16'd55672});
	test_expansion(128'heeca6c0db2984cab7b165d90a524d58f, {16'd1391, 16'd43634, 16'd28603, 16'd31804, 16'd11457, 16'd36818, 16'd50711, 16'd45555, 16'd63699, 16'd50112, 16'd39960, 16'd16491, 16'd45913, 16'd22061, 16'd19407, 16'd17987, 16'd17772, 16'd24326, 16'd44461, 16'd34218, 16'd51985, 16'd25028, 16'd21210, 16'd58805, 16'd9111, 16'd52652});
	test_expansion(128'h7a614b2077c6c5565ceda1ec555ccd6d, {16'd41341, 16'd59673, 16'd3544, 16'd65464, 16'd10279, 16'd14378, 16'd57876, 16'd20498, 16'd28018, 16'd24628, 16'd40162, 16'd8868, 16'd23601, 16'd22042, 16'd26223, 16'd47107, 16'd26068, 16'd56410, 16'd34041, 16'd46279, 16'd1909, 16'd37412, 16'd39790, 16'd13040, 16'd6281, 16'd5711});
	test_expansion(128'h75a3e306b8dd92f5cb695e6b9296dccd, {16'd21808, 16'd49331, 16'd34828, 16'd33475, 16'd8968, 16'd12569, 16'd35385, 16'd18401, 16'd64886, 16'd39261, 16'd35614, 16'd44509, 16'd20055, 16'd31407, 16'd28006, 16'd7660, 16'd9147, 16'd5083, 16'd20715, 16'd41621, 16'd58517, 16'd62441, 16'd6447, 16'd17287, 16'd24882, 16'd14718});
	test_expansion(128'hdcd603ee533696b59780c115ff3f2ec3, {16'd63611, 16'd62423, 16'd62039, 16'd16506, 16'd20333, 16'd31022, 16'd47181, 16'd25262, 16'd20042, 16'd1270, 16'd27390, 16'd53313, 16'd4539, 16'd27618, 16'd60252, 16'd53296, 16'd59354, 16'd64959, 16'd41185, 16'd25938, 16'd28474, 16'd45006, 16'd42425, 16'd29457, 16'd52052, 16'd58326});
	test_expansion(128'h2a1d20b8deeba2d9739582d55fb6a303, {16'd14486, 16'd53032, 16'd52933, 16'd7811, 16'd23884, 16'd3460, 16'd828, 16'd13075, 16'd495, 16'd20551, 16'd13965, 16'd49910, 16'd478, 16'd57586, 16'd46180, 16'd9734, 16'd8547, 16'd17968, 16'd39642, 16'd46635, 16'd40719, 16'd23621, 16'd61897, 16'd19263, 16'd9111, 16'd58957});
	test_expansion(128'h17554ca1a4fb23f3e4aa12b94fa1e3d9, {16'd53438, 16'd53221, 16'd29069, 16'd31093, 16'd39357, 16'd49333, 16'd54192, 16'd51030, 16'd8479, 16'd48737, 16'd55861, 16'd4422, 16'd27118, 16'd47889, 16'd33566, 16'd26323, 16'd55236, 16'd22207, 16'd4640, 16'd8420, 16'd41797, 16'd4919, 16'd17904, 16'd16042, 16'd48170, 16'd49967});
	test_expansion(128'hed9c15c28889a95fc7a96f690337cabf, {16'd40674, 16'd32449, 16'd21431, 16'd65066, 16'd10165, 16'd59930, 16'd214, 16'd16659, 16'd58208, 16'd40849, 16'd55767, 16'd59790, 16'd61507, 16'd49854, 16'd41354, 16'd32097, 16'd16757, 16'd51071, 16'd62327, 16'd14902, 16'd17394, 16'd54317, 16'd53619, 16'd63650, 16'd1175, 16'd20589});
	test_expansion(128'h11b2a6bbd846b87ff9369074201cbe8d, {16'd9578, 16'd5081, 16'd50077, 16'd17059, 16'd36438, 16'd58843, 16'd35713, 16'd31092, 16'd45739, 16'd57844, 16'd27580, 16'd7951, 16'd52347, 16'd5585, 16'd61108, 16'd61325, 16'd10528, 16'd30987, 16'd15863, 16'd47267, 16'd18650, 16'd3033, 16'd55845, 16'd801, 16'd672, 16'd39278});
	test_expansion(128'h1a6b8bd2d12b62b1e43979db05cac734, {16'd19133, 16'd22564, 16'd785, 16'd43103, 16'd17220, 16'd62753, 16'd41988, 16'd56368, 16'd57931, 16'd11624, 16'd14725, 16'd61929, 16'd52813, 16'd47231, 16'd10761, 16'd18277, 16'd32066, 16'd50544, 16'd43725, 16'd43623, 16'd22791, 16'd984, 16'd42653, 16'd47807, 16'd21765, 16'd53013});
	test_expansion(128'hca76aec97bd2e33ed9174e2f806b08c0, {16'd15759, 16'd60897, 16'd36993, 16'd26265, 16'd52813, 16'd27767, 16'd36897, 16'd64176, 16'd44182, 16'd56391, 16'd52986, 16'd47234, 16'd13797, 16'd12326, 16'd56673, 16'd34045, 16'd12993, 16'd58519, 16'd30337, 16'd8739, 16'd22542, 16'd13909, 16'd26189, 16'd20439, 16'd19404, 16'd60332});
	test_expansion(128'hcb0694a63705f7a50cc8653b7f71b7c4, {16'd47106, 16'd23975, 16'd57666, 16'd18528, 16'd5530, 16'd45331, 16'd55386, 16'd59993, 16'd33384, 16'd59394, 16'd40970, 16'd64792, 16'd17244, 16'd34738, 16'd63321, 16'd12705, 16'd3428, 16'd2030, 16'd49739, 16'd4559, 16'd60342, 16'd46659, 16'd31553, 16'd37768, 16'd47874, 16'd9698});
	test_expansion(128'h47bb36d3f2a5beb114233a94ad475a10, {16'd7028, 16'd34176, 16'd38976, 16'd20983, 16'd5739, 16'd24989, 16'd9924, 16'd11362, 16'd26303, 16'd64593, 16'd57048, 16'd18189, 16'd48796, 16'd14008, 16'd25049, 16'd21950, 16'd17107, 16'd57366, 16'd29387, 16'd23137, 16'd54186, 16'd43074, 16'd63871, 16'd47318, 16'd58049, 16'd39120});
	test_expansion(128'h99949a2c0a751215232ae2b5e84aeabf, {16'd31552, 16'd734, 16'd54814, 16'd40673, 16'd7132, 16'd31718, 16'd57485, 16'd57977, 16'd4219, 16'd12809, 16'd44337, 16'd57715, 16'd53519, 16'd14372, 16'd64895, 16'd33892, 16'd45472, 16'd27573, 16'd35129, 16'd63967, 16'd51323, 16'd125, 16'd23877, 16'd29559, 16'd27857, 16'd45040});
	test_expansion(128'h3aa59ba0f931ed751cebedd5f6c8917f, {16'd31664, 16'd28219, 16'd43247, 16'd55169, 16'd27729, 16'd9763, 16'd53204, 16'd4043, 16'd48516, 16'd55558, 16'd54686, 16'd6815, 16'd52937, 16'd13031, 16'd50293, 16'd35545, 16'd30232, 16'd17179, 16'd62453, 16'd44000, 16'd4869, 16'd21748, 16'd51344, 16'd52564, 16'd57507, 16'd40095});
	test_expansion(128'hc64ad226738d78d4c87e22c0775be81a, {16'd4526, 16'd43546, 16'd52090, 16'd45357, 16'd13896, 16'd53466, 16'd552, 16'd43926, 16'd41709, 16'd30547, 16'd31873, 16'd3151, 16'd65252, 16'd28952, 16'd50109, 16'd15397, 16'd989, 16'd50066, 16'd47149, 16'd8188, 16'd63900, 16'd1766, 16'd2767, 16'd28873, 16'd32703, 16'd52602});
	test_expansion(128'h2907cbae5006721e7467f640942cb7c7, {16'd2990, 16'd50204, 16'd32415, 16'd45999, 16'd57917, 16'd54038, 16'd45627, 16'd36498, 16'd3326, 16'd3018, 16'd33245, 16'd55204, 16'd34824, 16'd49338, 16'd22630, 16'd24803, 16'd58339, 16'd4588, 16'd8535, 16'd31334, 16'd43813, 16'd41819, 16'd62155, 16'd34499, 16'd57773, 16'd10287});
	test_expansion(128'hb2fbae8a59755381e28861034b572971, {16'd17011, 16'd41180, 16'd1711, 16'd49881, 16'd21912, 16'd45386, 16'd1188, 16'd58662, 16'd14075, 16'd22109, 16'd64518, 16'd2487, 16'd48714, 16'd49655, 16'd33097, 16'd46409, 16'd24721, 16'd50731, 16'd25314, 16'd60966, 16'd22369, 16'd29315, 16'd62043, 16'd54830, 16'd6482, 16'd8197});
	test_expansion(128'h1d39d367df8b62202ae55a65f4cb820a, {16'd5641, 16'd55876, 16'd35524, 16'd11175, 16'd38596, 16'd30915, 16'd31919, 16'd57885, 16'd61409, 16'd31398, 16'd46604, 16'd56984, 16'd58909, 16'd46456, 16'd17485, 16'd23998, 16'd22004, 16'd15029, 16'd48421, 16'd15184, 16'd10820, 16'd17933, 16'd59723, 16'd44779, 16'd24671, 16'd50820});
	test_expansion(128'hbf8f5f0675861492790f3015da3bde82, {16'd10102, 16'd57956, 16'd6090, 16'd22427, 16'd37511, 16'd16544, 16'd8539, 16'd57508, 16'd47699, 16'd23884, 16'd42403, 16'd24593, 16'd45118, 16'd57493, 16'd419, 16'd20058, 16'd59809, 16'd3528, 16'd51338, 16'd59422, 16'd7647, 16'd49248, 16'd24057, 16'd42285, 16'd27150, 16'd15128});
	test_expansion(128'hb9db524b9f0faeadd9ffa58aff606bc1, {16'd46046, 16'd16166, 16'd51886, 16'd48825, 16'd64397, 16'd54071, 16'd61953, 16'd25158, 16'd44221, 16'd50959, 16'd59967, 16'd9633, 16'd43982, 16'd46096, 16'd14319, 16'd51342, 16'd20340, 16'd2919, 16'd55010, 16'd21410, 16'd31210, 16'd23645, 16'd36462, 16'd5640, 16'd51273, 16'd35239});
	test_expansion(128'hd01b9ee38951fbc4f0acb89527083402, {16'd23913, 16'd35217, 16'd44877, 16'd50409, 16'd62683, 16'd3396, 16'd60666, 16'd30360, 16'd30023, 16'd36018, 16'd40338, 16'd18526, 16'd11770, 16'd4541, 16'd26828, 16'd57642, 16'd5510, 16'd4689, 16'd21368, 16'd57673, 16'd23128, 16'd23971, 16'd28905, 16'd31207, 16'd50177, 16'd58595});
	test_expansion(128'h62f53f2dbad42ca52a8bfd6faffe4c37, {16'd60892, 16'd40715, 16'd35489, 16'd3745, 16'd55860, 16'd57714, 16'd8686, 16'd63614, 16'd242, 16'd47859, 16'd36372, 16'd22968, 16'd12174, 16'd60731, 16'd49752, 16'd4877, 16'd14144, 16'd31479, 16'd17598, 16'd6558, 16'd54103, 16'd55838, 16'd33888, 16'd22267, 16'd46648, 16'd19430});
	test_expansion(128'h0811e44cb8cdc1bd04920390d007b4bf, {16'd9648, 16'd9965, 16'd57303, 16'd9142, 16'd50478, 16'd22391, 16'd44408, 16'd55401, 16'd64742, 16'd19905, 16'd27975, 16'd1395, 16'd53457, 16'd9335, 16'd62477, 16'd64396, 16'd53363, 16'd24782, 16'd32199, 16'd30786, 16'd59282, 16'd10708, 16'd2459, 16'd17635, 16'd3105, 16'd59836});
	test_expansion(128'h9ae36281f6e80fee7dd9d67c1cc95e71, {16'd33142, 16'd49232, 16'd21078, 16'd63489, 16'd38110, 16'd46490, 16'd7847, 16'd29594, 16'd6583, 16'd25261, 16'd51327, 16'd35876, 16'd55785, 16'd59442, 16'd22881, 16'd51780, 16'd29343, 16'd18535, 16'd8757, 16'd1780, 16'd5737, 16'd17332, 16'd28102, 16'd5714, 16'd59562, 16'd40471});
	test_expansion(128'hfa3fb39c5260097fc5734eed2a205e1e, {16'd15577, 16'd17190, 16'd48253, 16'd20931, 16'd10834, 16'd40415, 16'd16125, 16'd2079, 16'd18392, 16'd48112, 16'd11868, 16'd28290, 16'd34459, 16'd17899, 16'd54002, 16'd29280, 16'd8898, 16'd28768, 16'd40790, 16'd24177, 16'd39239, 16'd58364, 16'd8560, 16'd63371, 16'd62727, 16'd41374});
	test_expansion(128'hcb81f8e7b50ddafc7292b0638f8fddc5, {16'd8354, 16'd53626, 16'd42762, 16'd36718, 16'd28800, 16'd52031, 16'd41969, 16'd61878, 16'd15491, 16'd19460, 16'd54065, 16'd42173, 16'd14901, 16'd415, 16'd53481, 16'd20491, 16'd20218, 16'd54257, 16'd30214, 16'd29645, 16'd15050, 16'd40035, 16'd21599, 16'd54704, 16'd29001, 16'd35300});
	test_expansion(128'h260bdb7c38151f9ed81d8f4c3749a55f, {16'd15979, 16'd39987, 16'd25666, 16'd9974, 16'd39962, 16'd34671, 16'd53488, 16'd14176, 16'd60233, 16'd58749, 16'd16257, 16'd12937, 16'd37839, 16'd42563, 16'd62477, 16'd39324, 16'd22141, 16'd41749, 16'd38080, 16'd50296, 16'd64078, 16'd50167, 16'd30636, 16'd38391, 16'd53040, 16'd45671});
	test_expansion(128'h74b6ce8c97f4213c00e8024a1fa88b65, {16'd48764, 16'd60015, 16'd7808, 16'd63584, 16'd62734, 16'd39695, 16'd17594, 16'd21253, 16'd15453, 16'd12068, 16'd12580, 16'd38572, 16'd23676, 16'd60229, 16'd60724, 16'd31438, 16'd52965, 16'd34875, 16'd36738, 16'd62814, 16'd33959, 16'd61152, 16'd31338, 16'd61899, 16'd21642, 16'd49722});
	test_expansion(128'h99f3d0d0751be66967d8c9d083ae805b, {16'd53557, 16'd63304, 16'd22703, 16'd43583, 16'd22126, 16'd24236, 16'd49874, 16'd26896, 16'd7783, 16'd11027, 16'd8690, 16'd54384, 16'd63090, 16'd1943, 16'd41076, 16'd53422, 16'd45657, 16'd31231, 16'd58296, 16'd54015, 16'd5782, 16'd3462, 16'd11181, 16'd2111, 16'd19875, 16'd18644});
	test_expansion(128'ha57c6c26ede2d98e61c2f2043a3cc00b, {16'd43531, 16'd51987, 16'd21047, 16'd50234, 16'd56777, 16'd29224, 16'd64979, 16'd43963, 16'd56315, 16'd21224, 16'd22288, 16'd9675, 16'd21703, 16'd29924, 16'd44217, 16'd24208, 16'd18748, 16'd19622, 16'd13070, 16'd19152, 16'd30558, 16'd15116, 16'd30610, 16'd43510, 16'd49614, 16'd38773});
	test_expansion(128'h57e583737d8fe3bc147191abc345873d, {16'd33264, 16'd49556, 16'd43203, 16'd27285, 16'd2955, 16'd31576, 16'd8847, 16'd14411, 16'd64332, 16'd25325, 16'd10134, 16'd54744, 16'd32008, 16'd14287, 16'd23865, 16'd7719, 16'd48970, 16'd833, 16'd53689, 16'd48382, 16'd43214, 16'd56171, 16'd51882, 16'd13523, 16'd54293, 16'd46448});
	test_expansion(128'h7b454ffccce860122d2cfbd5577fa31c, {16'd49099, 16'd17694, 16'd61028, 16'd50207, 16'd22437, 16'd26778, 16'd6108, 16'd40905, 16'd22577, 16'd4419, 16'd50816, 16'd53266, 16'd52759, 16'd63748, 16'd18114, 16'd15066, 16'd22456, 16'd13840, 16'd42343, 16'd41878, 16'd53009, 16'd16491, 16'd63936, 16'd60736, 16'd14519, 16'd7298});
	test_expansion(128'hc60e27004fe6f97d37466c4b62c0836e, {16'd52525, 16'd37937, 16'd12576, 16'd34008, 16'd16150, 16'd11555, 16'd14691, 16'd61271, 16'd56198, 16'd62817, 16'd40937, 16'd43120, 16'd42849, 16'd1946, 16'd36949, 16'd18353, 16'd47057, 16'd64240, 16'd11192, 16'd14107, 16'd57245, 16'd19332, 16'd59658, 16'd53575, 16'd56722, 16'd22514});
	test_expansion(128'haee73bd740a549134aaaf36281f4efce, {16'd51205, 16'd2280, 16'd16170, 16'd38219, 16'd51955, 16'd33001, 16'd28952, 16'd15848, 16'd49516, 16'd36919, 16'd21355, 16'd43192, 16'd41520, 16'd50123, 16'd35283, 16'd37464, 16'd12167, 16'd38004, 16'd49393, 16'd55678, 16'd43900, 16'd12449, 16'd11321, 16'd65268, 16'd4558, 16'd8283});
	test_expansion(128'h6bb6d2a46bcb9e1f9742475b052ba95f, {16'd8859, 16'd46614, 16'd37692, 16'd11708, 16'd16947, 16'd28010, 16'd16581, 16'd23628, 16'd64883, 16'd28846, 16'd29646, 16'd20288, 16'd31135, 16'd54674, 16'd41863, 16'd29070, 16'd26656, 16'd32040, 16'd36395, 16'd61219, 16'd52738, 16'd35667, 16'd7126, 16'd38845, 16'd34077, 16'd60405});
	test_expansion(128'h072b4f91dd03f5744e2872dc7fcc7265, {16'd7901, 16'd27341, 16'd62576, 16'd11639, 16'd31540, 16'd1735, 16'd22598, 16'd15717, 16'd51539, 16'd14231, 16'd30490, 16'd59993, 16'd47959, 16'd39317, 16'd45455, 16'd13887, 16'd50906, 16'd15817, 16'd33029, 16'd16869, 16'd17060, 16'd15913, 16'd13171, 16'd7232, 16'd49477, 16'd7604});
	test_expansion(128'h5bbda52a724b4ed9ea5d78e8b45b2290, {16'd30400, 16'd50095, 16'd265, 16'd16839, 16'd29800, 16'd5184, 16'd64243, 16'd44555, 16'd17260, 16'd15562, 16'd2864, 16'd62063, 16'd31885, 16'd34548, 16'd54356, 16'd59504, 16'd51780, 16'd36156, 16'd17207, 16'd42274, 16'd4875, 16'd7208, 16'd37186, 16'd17889, 16'd34455, 16'd48816});
	test_expansion(128'h55cefe93b25f183440012133180953f9, {16'd8101, 16'd60834, 16'd29620, 16'd15605, 16'd14080, 16'd34597, 16'd24476, 16'd9672, 16'd65485, 16'd45390, 16'd3201, 16'd14010, 16'd36194, 16'd31207, 16'd41238, 16'd34794, 16'd33083, 16'd61283, 16'd13113, 16'd12762, 16'd19352, 16'd55511, 16'd42817, 16'd9041, 16'd27515, 16'd42186});
	test_expansion(128'hc9bb87b8076080d817ca3c123e2310b7, {16'd43141, 16'd11481, 16'd57538, 16'd46632, 16'd60893, 16'd23820, 16'd40789, 16'd26268, 16'd21926, 16'd33164, 16'd11726, 16'd18230, 16'd46897, 16'd13419, 16'd49113, 16'd52780, 16'd43751, 16'd47586, 16'd64537, 16'd1275, 16'd8441, 16'd16185, 16'd29463, 16'd24309, 16'd41644, 16'd29161});
	test_expansion(128'h11dd98358b3de330cedc48b27ce8c5e8, {16'd32459, 16'd27091, 16'd49553, 16'd25918, 16'd54596, 16'd40908, 16'd43247, 16'd22893, 16'd14048, 16'd1130, 16'd48236, 16'd59451, 16'd12840, 16'd30071, 16'd50778, 16'd16913, 16'd19994, 16'd28138, 16'd7083, 16'd43547, 16'd14742, 16'd53546, 16'd45842, 16'd55125, 16'd17428, 16'd38106});
	test_expansion(128'h8ef53e1cc04a1e223beefd9549f988da, {16'd38680, 16'd4154, 16'd42047, 16'd31699, 16'd2342, 16'd2485, 16'd22248, 16'd33484, 16'd52860, 16'd58220, 16'd11164, 16'd8045, 16'd8397, 16'd3970, 16'd16516, 16'd29987, 16'd59617, 16'd9576, 16'd44393, 16'd61833, 16'd60264, 16'd17378, 16'd44810, 16'd25401, 16'd29541, 16'd15053});
	test_expansion(128'h07b26e5f4d0b4fa4e60c314c6b252bcf, {16'd24317, 16'd19609, 16'd28065, 16'd40993, 16'd49935, 16'd38316, 16'd37146, 16'd49466, 16'd1642, 16'd38451, 16'd27835, 16'd47212, 16'd48095, 16'd61885, 16'd7820, 16'd42318, 16'd58383, 16'd4949, 16'd52506, 16'd49511, 16'd62684, 16'd17529, 16'd13666, 16'd29873, 16'd38476, 16'd26241});
	test_expansion(128'hc61c055e4c9cc962a4e91effc9250333, {16'd65006, 16'd27825, 16'd30852, 16'd43508, 16'd54676, 16'd32728, 16'd35312, 16'd7109, 16'd36079, 16'd9428, 16'd489, 16'd62205, 16'd2445, 16'd26254, 16'd63689, 16'd22878, 16'd1062, 16'd42847, 16'd27097, 16'd15519, 16'd6032, 16'd58191, 16'd2381, 16'd58666, 16'd35341, 16'd52195});
	test_expansion(128'hcc050c714573d1f3b18f7b63a9da2bba, {16'd41972, 16'd51793, 16'd34684, 16'd37940, 16'd21466, 16'd19463, 16'd30372, 16'd27435, 16'd33265, 16'd4322, 16'd34048, 16'd19121, 16'd63237, 16'd51221, 16'd25920, 16'd26890, 16'd48794, 16'd19642, 16'd7724, 16'd62268, 16'd10374, 16'd51321, 16'd21270, 16'd45626, 16'd49394, 16'd5187});
	test_expansion(128'hbba500ac18d415a3de3cdec04b2b69bf, {16'd22265, 16'd49862, 16'd23619, 16'd65245, 16'd13120, 16'd15664, 16'd10562, 16'd29244, 16'd61165, 16'd8940, 16'd40537, 16'd57202, 16'd34755, 16'd54547, 16'd33473, 16'd37654, 16'd41789, 16'd14960, 16'd8624, 16'd59104, 16'd1162, 16'd26647, 16'd22664, 16'd33644, 16'd46778, 16'd37329});
	test_expansion(128'h9a1404f50edc462992539d43635f0b61, {16'd35692, 16'd11153, 16'd37783, 16'd5199, 16'd4486, 16'd42714, 16'd10211, 16'd2187, 16'd4317, 16'd55284, 16'd53711, 16'd44069, 16'd4624, 16'd10720, 16'd64732, 16'd47528, 16'd10830, 16'd13898, 16'd8138, 16'd3814, 16'd25826, 16'd13281, 16'd30683, 16'd49763, 16'd54140, 16'd41918});
	test_expansion(128'h5fd4df8d06aaf2ffeb60e148fc1cc683, {16'd65110, 16'd6406, 16'd56706, 16'd26286, 16'd57355, 16'd29207, 16'd36253, 16'd28728, 16'd65192, 16'd55872, 16'd32800, 16'd29880, 16'd45923, 16'd6784, 16'd34405, 16'd36132, 16'd55835, 16'd42132, 16'd1505, 16'd31347, 16'd62167, 16'd63997, 16'd41394, 16'd9768, 16'd30248, 16'd1503});
	test_expansion(128'h6069e14143f76cc76b3dd804e0e6725a, {16'd9217, 16'd40566, 16'd20952, 16'd57834, 16'd33353, 16'd57698, 16'd39175, 16'd11892, 16'd12960, 16'd22753, 16'd51056, 16'd4199, 16'd40570, 16'd3612, 16'd57014, 16'd36869, 16'd7591, 16'd51807, 16'd6367, 16'd41032, 16'd55640, 16'd33775, 16'd12573, 16'd31270, 16'd31867, 16'd48523});
	test_expansion(128'h806b1dd29612a8756ee591beb19b3b49, {16'd37038, 16'd41799, 16'd36296, 16'd30318, 16'd64314, 16'd18990, 16'd20491, 16'd60859, 16'd13169, 16'd64869, 16'd3394, 16'd48287, 16'd42360, 16'd61869, 16'd35683, 16'd57992, 16'd4973, 16'd34143, 16'd20994, 16'd56824, 16'd48648, 16'd34467, 16'd3501, 16'd34646, 16'd28847, 16'd59359});
	test_expansion(128'h31eb355e93ef2a5556f509a117e7a29d, {16'd23776, 16'd4733, 16'd36799, 16'd30529, 16'd42887, 16'd8005, 16'd19208, 16'd55934, 16'd62907, 16'd37166, 16'd17636, 16'd23420, 16'd37000, 16'd34805, 16'd30179, 16'd12416, 16'd58244, 16'd34287, 16'd55203, 16'd13770, 16'd58349, 16'd48680, 16'd14648, 16'd57412, 16'd33665, 16'd54613});
	test_expansion(128'h20acdd2c5a9c35e14ecf93a761617b56, {16'd16465, 16'd13234, 16'd14864, 16'd64891, 16'd44693, 16'd63205, 16'd36213, 16'd32041, 16'd39800, 16'd58885, 16'd27866, 16'd13162, 16'd48696, 16'd35025, 16'd40007, 16'd27220, 16'd57906, 16'd63521, 16'd15133, 16'd18151, 16'd39859, 16'd17362, 16'd20642, 16'd47860, 16'd49419, 16'd15721});
	test_expansion(128'h1bf1b345af1c41248df6e79d4b98bb2b, {16'd41023, 16'd12344, 16'd45283, 16'd46162, 16'd29890, 16'd12606, 16'd59430, 16'd40173, 16'd22982, 16'd65369, 16'd28645, 16'd2877, 16'd30856, 16'd34299, 16'd1675, 16'd42730, 16'd45781, 16'd11017, 16'd57171, 16'd43208, 16'd57616, 16'd19245, 16'd13976, 16'd24150, 16'd31562, 16'd21802});
	test_expansion(128'hd6f55e8c0aeb12a6af3ec5e6f16bf73d, {16'd4946, 16'd25360, 16'd20756, 16'd17371, 16'd26960, 16'd64542, 16'd41473, 16'd3815, 16'd54446, 16'd58585, 16'd36280, 16'd40363, 16'd847, 16'd61703, 16'd38763, 16'd29783, 16'd56913, 16'd47134, 16'd59187, 16'd2673, 16'd5156, 16'd7608, 16'd63270, 16'd34775, 16'd28795, 16'd29582});
	test_expansion(128'hbc27e6d7afc8196a17863abd27f9a615, {16'd31190, 16'd37145, 16'd36968, 16'd36292, 16'd2040, 16'd27854, 16'd1258, 16'd10628, 16'd26781, 16'd28783, 16'd22749, 16'd27490, 16'd51388, 16'd58316, 16'd49912, 16'd39492, 16'd6142, 16'd17499, 16'd16665, 16'd16244, 16'd45323, 16'd56829, 16'd44050, 16'd15957, 16'd2509, 16'd45736});
	test_expansion(128'hc02387a976b5c57f73f400cedecc9323, {16'd47417, 16'd2358, 16'd39795, 16'd38885, 16'd3522, 16'd45833, 16'd28350, 16'd51405, 16'd60742, 16'd20031, 16'd52287, 16'd10044, 16'd41183, 16'd54637, 16'd27062, 16'd275, 16'd41802, 16'd13669, 16'd7583, 16'd17262, 16'd50188, 16'd8241, 16'd62121, 16'd23902, 16'd53645, 16'd48774});
	test_expansion(128'h848179be5acfd4392e1a4a2e0f928c1a, {16'd7155, 16'd27674, 16'd52580, 16'd6944, 16'd29390, 16'd25649, 16'd32369, 16'd56502, 16'd44108, 16'd14518, 16'd482, 16'd30978, 16'd34449, 16'd16203, 16'd60579, 16'd25248, 16'd20562, 16'd32869, 16'd18923, 16'd32305, 16'd26623, 16'd45379, 16'd54422, 16'd45179, 16'd35964, 16'd36133});
	test_expansion(128'h2c6b6c18feb6391cd7c4c83c12182516, {16'd41748, 16'd37395, 16'd48653, 16'd22770, 16'd25639, 16'd35232, 16'd30993, 16'd8062, 16'd51946, 16'd34982, 16'd50478, 16'd12424, 16'd4636, 16'd47928, 16'd63846, 16'd58840, 16'd4924, 16'd46599, 16'd29681, 16'd47222, 16'd2092, 16'd6705, 16'd28806, 16'd21406, 16'd30227, 16'd30219});
	test_expansion(128'h332ac3d576dcc6e23cde98762de6cb20, {16'd23846, 16'd28015, 16'd41082, 16'd47333, 16'd29939, 16'd38142, 16'd59522, 16'd21858, 16'd7854, 16'd1302, 16'd38228, 16'd23313, 16'd23108, 16'd41460, 16'd53174, 16'd63662, 16'd29545, 16'd63879, 16'd11978, 16'd62951, 16'd31646, 16'd64865, 16'd33757, 16'd24678, 16'd923, 16'd45520});
	test_expansion(128'h1f9d588f832324436891d236990e5273, {16'd14558, 16'd48864, 16'd63523, 16'd64832, 16'd62144, 16'd18756, 16'd13153, 16'd13383, 16'd42198, 16'd51703, 16'd1067, 16'd52872, 16'd25641, 16'd1970, 16'd42524, 16'd13930, 16'd6222, 16'd41251, 16'd18162, 16'd37525, 16'd1422, 16'd7624, 16'd47694, 16'd57027, 16'd19045, 16'd23149});
	test_expansion(128'h5f55e649477bdbd26023837820803c46, {16'd62995, 16'd26507, 16'd9670, 16'd16176, 16'd34688, 16'd29059, 16'd54000, 16'd55234, 16'd38114, 16'd45229, 16'd51512, 16'd50584, 16'd51064, 16'd7333, 16'd36835, 16'd41707, 16'd193, 16'd57896, 16'd40296, 16'd1670, 16'd51559, 16'd51042, 16'd15130, 16'd61586, 16'd32347, 16'd47814});
	test_expansion(128'h4e26abc26b964290b4a5b8d8cd887f26, {16'd1275, 16'd47645, 16'd37865, 16'd25029, 16'd20385, 16'd42804, 16'd53777, 16'd63214, 16'd46638, 16'd55862, 16'd52067, 16'd44250, 16'd1152, 16'd21061, 16'd57690, 16'd36215, 16'd55449, 16'd29569, 16'd10788, 16'd23876, 16'd29233, 16'd29374, 16'd64311, 16'd52373, 16'd3196, 16'd84});
	test_expansion(128'hf15622941351c24fa1aedf4c508dd59f, {16'd5456, 16'd11763, 16'd32672, 16'd54688, 16'd29945, 16'd54517, 16'd6428, 16'd42990, 16'd54470, 16'd47560, 16'd6821, 16'd12507, 16'd8795, 16'd31805, 16'd38631, 16'd18829, 16'd32254, 16'd55525, 16'd30284, 16'd42674, 16'd18197, 16'd43676, 16'd32009, 16'd60201, 16'd33646, 16'd398});
	test_expansion(128'h0cb49a7c14370039941cca446c7e4e23, {16'd22511, 16'd33894, 16'd53060, 16'd17349, 16'd24856, 16'd64328, 16'd36603, 16'd62295, 16'd13358, 16'd26838, 16'd64225, 16'd5779, 16'd38039, 16'd36187, 16'd16069, 16'd52930, 16'd37572, 16'd56660, 16'd37202, 16'd1055, 16'd51306, 16'd40842, 16'd35590, 16'd40346, 16'd24945, 16'd50034});
	test_expansion(128'hdb0c64589b152a4c5ce6323b4786f56e, {16'd61528, 16'd54905, 16'd58348, 16'd11776, 16'd56365, 16'd36900, 16'd64242, 16'd7352, 16'd55618, 16'd7570, 16'd43895, 16'd37660, 16'd27871, 16'd21101, 16'd53455, 16'd59341, 16'd49038, 16'd54323, 16'd20658, 16'd22103, 16'd6022, 16'd16552, 16'd57507, 16'd58764, 16'd6471, 16'd22607});
	test_expansion(128'h889c5dda1ae038ca6ea6a9b619a59ce5, {16'd9118, 16'd36513, 16'd47499, 16'd1432, 16'd27642, 16'd48407, 16'd20511, 16'd54707, 16'd20652, 16'd28165, 16'd44882, 16'd53898, 16'd46327, 16'd62256, 16'd61502, 16'd27948, 16'd16337, 16'd56354, 16'd45654, 16'd52347, 16'd58032, 16'd39402, 16'd57404, 16'd63855, 16'd18957, 16'd26927});
	test_expansion(128'hc5032b4b88788bef2d52361e74e5c146, {16'd32151, 16'd22821, 16'd5829, 16'd47547, 16'd56501, 16'd50111, 16'd36751, 16'd37527, 16'd55851, 16'd50664, 16'd41632, 16'd33091, 16'd43091, 16'd1745, 16'd14892, 16'd55039, 16'd9639, 16'd30158, 16'd11527, 16'd34686, 16'd20058, 16'd41374, 16'd63506, 16'd63805, 16'd35251, 16'd15065});
	test_expansion(128'h89b9b577efb70f0ae6b3e19f796aed6d, {16'd41695, 16'd55810, 16'd63478, 16'd24144, 16'd26493, 16'd21721, 16'd41574, 16'd34086, 16'd56565, 16'd55025, 16'd56614, 16'd49664, 16'd61267, 16'd10309, 16'd11810, 16'd5228, 16'd19884, 16'd3775, 16'd56422, 16'd22825, 16'd3754, 16'd9118, 16'd10509, 16'd62495, 16'd1152, 16'd24008});
	test_expansion(128'h2ef35cfea7c23f90bb576d8bcb47ddde, {16'd11044, 16'd42498, 16'd29904, 16'd21105, 16'd25699, 16'd26131, 16'd17433, 16'd19261, 16'd49614, 16'd46514, 16'd198, 16'd12264, 16'd48391, 16'd38452, 16'd15504, 16'd59921, 16'd17906, 16'd22159, 16'd24653, 16'd63251, 16'd56576, 16'd45085, 16'd10939, 16'd24761, 16'd21857, 16'd6629});
	test_expansion(128'ha30682253b14294820caf1e43a4d7478, {16'd2276, 16'd9728, 16'd16262, 16'd34451, 16'd20925, 16'd57214, 16'd5163, 16'd56882, 16'd13656, 16'd31636, 16'd59983, 16'd17947, 16'd42131, 16'd8021, 16'd2572, 16'd51524, 16'd62383, 16'd21888, 16'd21904, 16'd31196, 16'd11752, 16'd45464, 16'd60918, 16'd53348, 16'd32251, 16'd56836});
	test_expansion(128'hfdd545b5ef4d2dd989b5ce0c41e9b56f, {16'd39402, 16'd46916, 16'd13997, 16'd33913, 16'd6880, 16'd28725, 16'd14312, 16'd52860, 16'd45939, 16'd30562, 16'd59456, 16'd53870, 16'd30660, 16'd43125, 16'd60002, 16'd23273, 16'd57906, 16'd42086, 16'd20672, 16'd21630, 16'd21871, 16'd22477, 16'd3172, 16'd51695, 16'd19388, 16'd5154});
	test_expansion(128'hd0895427cc924e58fffa2f7a2fe39dfd, {16'd59185, 16'd51510, 16'd33763, 16'd1932, 16'd31568, 16'd65225, 16'd58169, 16'd7556, 16'd63631, 16'd62419, 16'd14267, 16'd57834, 16'd48675, 16'd62485, 16'd18189, 16'd16159, 16'd19928, 16'd55592, 16'd23251, 16'd29946, 16'd38792, 16'd25480, 16'd60727, 16'd39141, 16'd51609, 16'd29162});
	test_expansion(128'h792ff1989e750fcd7ac644b31a6236e1, {16'd24566, 16'd13710, 16'd49712, 16'd25483, 16'd46208, 16'd9069, 16'd14842, 16'd19666, 16'd34348, 16'd605, 16'd41196, 16'd40797, 16'd48819, 16'd5276, 16'd36694, 16'd49224, 16'd47879, 16'd36279, 16'd58680, 16'd58906, 16'd53522, 16'd29672, 16'd3342, 16'd38131, 16'd17914, 16'd8127});
	test_expansion(128'ha31ead212657e3a3f41c1dbacc7c3c53, {16'd62493, 16'd45179, 16'd21175, 16'd6579, 16'd36187, 16'd16642, 16'd28080, 16'd63480, 16'd8563, 16'd37634, 16'd32855, 16'd65400, 16'd65022, 16'd15340, 16'd24205, 16'd51672, 16'd64829, 16'd52345, 16'd13208, 16'd16409, 16'd20523, 16'd22874, 16'd42697, 16'd21759, 16'd58687, 16'd43729});
	test_expansion(128'hf6d5383ec8c7e28d36923b25e252a17b, {16'd48635, 16'd44266, 16'd62489, 16'd34265, 16'd3219, 16'd2111, 16'd38130, 16'd61742, 16'd8765, 16'd4913, 16'd21224, 16'd55114, 16'd3210, 16'd12169, 16'd23306, 16'd4894, 16'd7516, 16'd5799, 16'd5713, 16'd45531, 16'd32764, 16'd24594, 16'd64346, 16'd57539, 16'd64841, 16'd63088});
	test_expansion(128'ha8e17988c13c81ce82f11d4a6120a217, {16'd37578, 16'd22666, 16'd39689, 16'd36879, 16'd49644, 16'd8637, 16'd25427, 16'd29280, 16'd28004, 16'd41746, 16'd18156, 16'd55086, 16'd63402, 16'd46249, 16'd64376, 16'd40344, 16'd5689, 16'd13826, 16'd34958, 16'd46634, 16'd41694, 16'd3486, 16'd60380, 16'd33971, 16'd55364, 16'd25138});
	test_expansion(128'hd06b686bb3ff941fbc74ca6898e3ddb6, {16'd32245, 16'd56659, 16'd59507, 16'd18635, 16'd15137, 16'd18485, 16'd59557, 16'd60412, 16'd19056, 16'd35993, 16'd5173, 16'd60864, 16'd25640, 16'd50555, 16'd17033, 16'd30397, 16'd4211, 16'd18542, 16'd19759, 16'd55786, 16'd5835, 16'd24214, 16'd42272, 16'd50707, 16'd7357, 16'd33637});
	test_expansion(128'h9fe1b55498caa26338e7044c532fc0a8, {16'd45004, 16'd14498, 16'd5924, 16'd55152, 16'd17353, 16'd53482, 16'd49522, 16'd48454, 16'd44015, 16'd63628, 16'd3878, 16'd64965, 16'd61648, 16'd45838, 16'd9747, 16'd18097, 16'd57014, 16'd38163, 16'd35879, 16'd29522, 16'd58897, 16'd27670, 16'd60571, 16'd24062, 16'd65328, 16'd4304});
	test_expansion(128'had628d38a5982cd6fe0b306c09a3478d, {16'd8287, 16'd62485, 16'd47619, 16'd40001, 16'd19418, 16'd65331, 16'd21449, 16'd38438, 16'd65476, 16'd51376, 16'd12699, 16'd61770, 16'd27707, 16'd7201, 16'd13969, 16'd30387, 16'd47944, 16'd2097, 16'd42973, 16'd24600, 16'd43386, 16'd19645, 16'd23616, 16'd16326, 16'd5891, 16'd15526});
	test_expansion(128'h7c5ff23894768752e4d6f61b50a672e3, {16'd29134, 16'd10498, 16'd50625, 16'd2745, 16'd63394, 16'd24188, 16'd36583, 16'd26310, 16'd63344, 16'd39746, 16'd1146, 16'd32916, 16'd17267, 16'd27131, 16'd37285, 16'd725, 16'd41404, 16'd45626, 16'd2798, 16'd41104, 16'd37118, 16'd1277, 16'd27184, 16'd6071, 16'd31819, 16'd24335});
	test_expansion(128'h6926921dfa34167801771f8e4afd6795, {16'd62575, 16'd10346, 16'd41899, 16'd52196, 16'd53500, 16'd14495, 16'd30109, 16'd29806, 16'd39444, 16'd18550, 16'd15009, 16'd63236, 16'd47841, 16'd33058, 16'd46833, 16'd27186, 16'd13756, 16'd23463, 16'd16243, 16'd42508, 16'd7995, 16'd10823, 16'd33500, 16'd64388, 16'd38965, 16'd9328});
	test_expansion(128'hfa6b3b7c8a1126760bc767df49c54b61, {16'd2326, 16'd5722, 16'd2992, 16'd18259, 16'd15483, 16'd9435, 16'd21402, 16'd53341, 16'd59715, 16'd4952, 16'd24717, 16'd41298, 16'd9418, 16'd4049, 16'd20799, 16'd42750, 16'd26772, 16'd54041, 16'd63967, 16'd657, 16'd9274, 16'd24703, 16'd29483, 16'd51851, 16'd53323, 16'd48854});
	test_expansion(128'hc9877acec65964560650ee15f1cc09ba, {16'd5609, 16'd53502, 16'd57412, 16'd8640, 16'd55238, 16'd40196, 16'd59971, 16'd25554, 16'd3428, 16'd38557, 16'd46318, 16'd50372, 16'd16632, 16'd53949, 16'd55888, 16'd4786, 16'd31419, 16'd55219, 16'd47001, 16'd27188, 16'd6368, 16'd23448, 16'd3096, 16'd5297, 16'd15062, 16'd12098});
	test_expansion(128'h4ec50277d0a6451b4aaf0e81f9761b96, {16'd65258, 16'd9805, 16'd36093, 16'd11613, 16'd7561, 16'd1083, 16'd35490, 16'd16110, 16'd723, 16'd19709, 16'd24192, 16'd55131, 16'd14364, 16'd15723, 16'd35986, 16'd11467, 16'd45486, 16'd22738, 16'd61720, 16'd7761, 16'd13271, 16'd9469, 16'd36623, 16'd29487, 16'd17668, 16'd22052});
	test_expansion(128'h402a3f0a55a56c01215b6d08100546b0, {16'd505, 16'd28978, 16'd21938, 16'd59163, 16'd24822, 16'd33527, 16'd17358, 16'd20731, 16'd9611, 16'd7277, 16'd26007, 16'd52080, 16'd25595, 16'd8269, 16'd17437, 16'd63886, 16'd39804, 16'd60103, 16'd13187, 16'd48030, 16'd8378, 16'd5694, 16'd18456, 16'd34561, 16'd37263, 16'd10288});
	test_expansion(128'hd3a461ae211f32b983b708e9fbf9c296, {16'd8975, 16'd11951, 16'd46011, 16'd2796, 16'd2544, 16'd36175, 16'd26862, 16'd15234, 16'd37023, 16'd20863, 16'd56203, 16'd40161, 16'd35862, 16'd24873, 16'd60789, 16'd32795, 16'd58994, 16'd16967, 16'd7809, 16'd33232, 16'd52659, 16'd14582, 16'd47119, 16'd63584, 16'd45808, 16'd34594});
	test_expansion(128'h525faebf1b6105553b35858ce9301cf3, {16'd40259, 16'd1997, 16'd43274, 16'd25503, 16'd16222, 16'd52646, 16'd22144, 16'd57065, 16'd13479, 16'd35307, 16'd27326, 16'd20060, 16'd28561, 16'd12168, 16'd23098, 16'd34839, 16'd39356, 16'd10071, 16'd21013, 16'd23932, 16'd28262, 16'd24117, 16'd17036, 16'd43388, 16'd16967, 16'd26764});
	test_expansion(128'he3d5c90c1cf21a8041ac8f705930d3c6, {16'd29467, 16'd17389, 16'd132, 16'd24702, 16'd14658, 16'd8945, 16'd13192, 16'd41140, 16'd23457, 16'd12891, 16'd33363, 16'd54374, 16'd61642, 16'd51661, 16'd60596, 16'd30274, 16'd50793, 16'd22846, 16'd58876, 16'd15875, 16'd62895, 16'd60927, 16'd3872, 16'd45127, 16'd21422, 16'd60520});
	test_expansion(128'hb2f286188fb9dcaf1917211626957827, {16'd23071, 16'd39247, 16'd29949, 16'd16694, 16'd5830, 16'd59632, 16'd42681, 16'd11986, 16'd53637, 16'd14446, 16'd23375, 16'd10696, 16'd49308, 16'd14928, 16'd38342, 16'd46834, 16'd9461, 16'd23350, 16'd19941, 16'd24485, 16'd62855, 16'd51734, 16'd19168, 16'd45903, 16'd4914, 16'd39457});
	test_expansion(128'hd75d416ee68b48ac87cdaee724061b64, {16'd42300, 16'd41072, 16'd32854, 16'd5070, 16'd51333, 16'd46134, 16'd53272, 16'd53173, 16'd65389, 16'd23587, 16'd34350, 16'd29733, 16'd4440, 16'd42554, 16'd57597, 16'd65195, 16'd53153, 16'd35064, 16'd61922, 16'd36972, 16'd52683, 16'd52724, 16'd60546, 16'd39388, 16'd42293, 16'd42625});
	test_expansion(128'h333b9f4310f62e1af2164f49e6c31095, {16'd54646, 16'd61260, 16'd13935, 16'd56737, 16'd152, 16'd21145, 16'd54686, 16'd38463, 16'd11438, 16'd63061, 16'd63770, 16'd33875, 16'd14902, 16'd51021, 16'd25135, 16'd31801, 16'd20726, 16'd14154, 16'd4303, 16'd19979, 16'd24763, 16'd14136, 16'd29797, 16'd13740, 16'd26001, 16'd54823});
	test_expansion(128'hca7595ac2cc043b4188752851f967694, {16'd28992, 16'd61342, 16'd40573, 16'd29798, 16'd26599, 16'd37900, 16'd759, 16'd16506, 16'd55056, 16'd63898, 16'd17215, 16'd9435, 16'd41538, 16'd16883, 16'd60362, 16'd14038, 16'd35305, 16'd63915, 16'd55989, 16'd4852, 16'd45175, 16'd7957, 16'd63815, 16'd39806, 16'd16472, 16'd36191});
	test_expansion(128'h641bba512bcdbc29cc9bcd53affb9dd0, {16'd20020, 16'd37778, 16'd30853, 16'd6004, 16'd65280, 16'd3760, 16'd6091, 16'd41036, 16'd47588, 16'd42907, 16'd12276, 16'd63862, 16'd3725, 16'd10679, 16'd62841, 16'd9201, 16'd58882, 16'd41396, 16'd3510, 16'd56182, 16'd55053, 16'd61556, 16'd45736, 16'd21639, 16'd19474, 16'd32340});
	test_expansion(128'h3981f604cc46c1314bb4b3abf34b496f, {16'd31552, 16'd49681, 16'd23130, 16'd15632, 16'd37646, 16'd52916, 16'd21341, 16'd49084, 16'd14656, 16'd42660, 16'd33684, 16'd10628, 16'd43283, 16'd56348, 16'd29916, 16'd29619, 16'd45381, 16'd57165, 16'd14600, 16'd39511, 16'd7507, 16'd64862, 16'd40119, 16'd60566, 16'd56682, 16'd6589});
	test_expansion(128'h0cb72325a9192a6a635c980ad221dde5, {16'd94, 16'd18101, 16'd65150, 16'd21230, 16'd12312, 16'd19380, 16'd30218, 16'd56998, 16'd27880, 16'd35920, 16'd4194, 16'd30466, 16'd45960, 16'd12966, 16'd51939, 16'd42884, 16'd53136, 16'd33044, 16'd34360, 16'd10647, 16'd35913, 16'd62591, 16'd27958, 16'd63349, 16'd32798, 16'd28957});
	test_expansion(128'he31d657a0d362ed6e9d4d6e6155b678b, {16'd58240, 16'd32507, 16'd44071, 16'd6, 16'd27213, 16'd53968, 16'd47655, 16'd23096, 16'd16856, 16'd15974, 16'd51123, 16'd33734, 16'd45195, 16'd45769, 16'd23986, 16'd52336, 16'd3205, 16'd59593, 16'd30877, 16'd50294, 16'd26326, 16'd24631, 16'd9448, 16'd5848, 16'd63199, 16'd22490});
	test_expansion(128'h14a4fed250daf08a1dd7af1c14804911, {16'd50665, 16'd24051, 16'd16422, 16'd40279, 16'd53908, 16'd19864, 16'd84, 16'd60537, 16'd21768, 16'd10653, 16'd3604, 16'd58426, 16'd756, 16'd33782, 16'd64258, 16'd54859, 16'd40876, 16'd55761, 16'd52583, 16'd6227, 16'd20181, 16'd30964, 16'd39908, 16'd59873, 16'd20679, 16'd50936});
	test_expansion(128'hb56ae6267d4edc3311c1d37ef777f179, {16'd6483, 16'd21522, 16'd4187, 16'd47880, 16'd51909, 16'd33946, 16'd29529, 16'd63302, 16'd3395, 16'd20747, 16'd53897, 16'd25024, 16'd58112, 16'd42316, 16'd7798, 16'd38425, 16'd44836, 16'd9980, 16'd14205, 16'd22668, 16'd54764, 16'd60396, 16'd16788, 16'd11301, 16'd64694, 16'd56914});
	test_expansion(128'h9036c02b65306e61cf542f2aaf0c22a8, {16'd34773, 16'd12836, 16'd46063, 16'd41608, 16'd60445, 16'd5478, 16'd57471, 16'd4159, 16'd60139, 16'd24156, 16'd17314, 16'd36193, 16'd45297, 16'd55732, 16'd14389, 16'd5768, 16'd27973, 16'd46672, 16'd60322, 16'd48805, 16'd43150, 16'd31721, 16'd53572, 16'd55791, 16'd44863, 16'd10314});
	test_expansion(128'h31e7dd78e4bc694301f594692fa6e491, {16'd59795, 16'd14308, 16'd4033, 16'd816, 16'd58275, 16'd34204, 16'd6257, 16'd37417, 16'd65199, 16'd60934, 16'd8650, 16'd28500, 16'd39445, 16'd33750, 16'd5648, 16'd55958, 16'd27863, 16'd41961, 16'd57389, 16'd21910, 16'd62727, 16'd22493, 16'd31898, 16'd28796, 16'd52701, 16'd46679});
	test_expansion(128'h4a743220103eb2d0d098392388b4bd7b, {16'd40580, 16'd24418, 16'd54108, 16'd48827, 16'd39813, 16'd37983, 16'd25031, 16'd3906, 16'd47218, 16'd6391, 16'd58810, 16'd7594, 16'd31092, 16'd45173, 16'd61941, 16'd48838, 16'd59797, 16'd64536, 16'd41675, 16'd3184, 16'd44493, 16'd13203, 16'd27917, 16'd2601, 16'd37518, 16'd20813});
	test_expansion(128'h4f682681ee6617a89c457efa556154c8, {16'd39890, 16'd54272, 16'd30589, 16'd32255, 16'd28585, 16'd21157, 16'd23982, 16'd29787, 16'd2882, 16'd36892, 16'd56118, 16'd2930, 16'd44736, 16'd28241, 16'd60875, 16'd3635, 16'd28290, 16'd36221, 16'd64115, 16'd16914, 16'd59761, 16'd64214, 16'd6538, 16'd57009, 16'd34405, 16'd49747});
	test_expansion(128'h977b561dfea92c97465cb36a988f9678, {16'd32955, 16'd12976, 16'd9476, 16'd35525, 16'd3908, 16'd22102, 16'd64034, 16'd53095, 16'd12185, 16'd53338, 16'd39548, 16'd4009, 16'd58046, 16'd48190, 16'd54686, 16'd8552, 16'd62015, 16'd18392, 16'd55942, 16'd7973, 16'd48264, 16'd51841, 16'd40192, 16'd13022, 16'd26858, 16'd9113});
	test_expansion(128'h56dc79abcad6be3e65bd02cd282a4f26, {16'd3019, 16'd52220, 16'd51588, 16'd63380, 16'd50968, 16'd16743, 16'd10870, 16'd29556, 16'd34538, 16'd54693, 16'd62996, 16'd54588, 16'd20149, 16'd51505, 16'd14178, 16'd25284, 16'd54911, 16'd7919, 16'd49203, 16'd52689, 16'd38111, 16'd26311, 16'd61336, 16'd33279, 16'd62621, 16'd36001});
	test_expansion(128'h15d29f5e26d42e7095501b92b47aadaf, {16'd19261, 16'd4375, 16'd27567, 16'd7048, 16'd22282, 16'd24232, 16'd26492, 16'd15756, 16'd20829, 16'd30236, 16'd7711, 16'd36528, 16'd4363, 16'd35935, 16'd55539, 16'd34838, 16'd12565, 16'd6701, 16'd18390, 16'd13171, 16'd10563, 16'd21621, 16'd12648, 16'd48021, 16'd38698, 16'd45267});
	test_expansion(128'h23d4bbe9c6d299b80c3e23b791122c6b, {16'd40977, 16'd7036, 16'd52555, 16'd20638, 16'd40404, 16'd10879, 16'd34202, 16'd58056, 16'd26794, 16'd12368, 16'd45398, 16'd30258, 16'd23148, 16'd20946, 16'd59867, 16'd39459, 16'd26204, 16'd8513, 16'd51521, 16'd10139, 16'd11476, 16'd15359, 16'd35979, 16'd18896, 16'd56160, 16'd15520});
	test_expansion(128'h389d48f04e237537be54be74bc7d72e5, {16'd42639, 16'd7321, 16'd20858, 16'd18835, 16'd4184, 16'd11657, 16'd10033, 16'd48957, 16'd59281, 16'd62730, 16'd38358, 16'd51750, 16'd17807, 16'd8034, 16'd1432, 16'd21737, 16'd56264, 16'd59609, 16'd55979, 16'd46969, 16'd30657, 16'd46105, 16'd41986, 16'd35329, 16'd19760, 16'd1296});
	test_expansion(128'h39494b43530048d8ec12aac7a093c49b, {16'd12337, 16'd48755, 16'd44018, 16'd7050, 16'd11399, 16'd20414, 16'd65201, 16'd48561, 16'd17381, 16'd11423, 16'd14104, 16'd58056, 16'd59303, 16'd39279, 16'd34650, 16'd55490, 16'd61049, 16'd21988, 16'd48432, 16'd2978, 16'd30545, 16'd24137, 16'd37202, 16'd43074, 16'd20295, 16'd16460});
	test_expansion(128'h1bd00aecba039cc5ed23c9e243898caa, {16'd4050, 16'd2774, 16'd40768, 16'd33226, 16'd43349, 16'd33780, 16'd23303, 16'd20990, 16'd30221, 16'd54786, 16'd30713, 16'd42185, 16'd38675, 16'd38478, 16'd17404, 16'd8044, 16'd35111, 16'd22454, 16'd10404, 16'd34391, 16'd5104, 16'd18918, 16'd14733, 16'd15153, 16'd33734, 16'd27037});
	test_expansion(128'h973a6763d07e5ce1167309bb855e1028, {16'd8237, 16'd5266, 16'd16480, 16'd30189, 16'd35934, 16'd43589, 16'd28918, 16'd12037, 16'd19914, 16'd53734, 16'd40955, 16'd47029, 16'd63642, 16'd45955, 16'd13278, 16'd19218, 16'd12184, 16'd22767, 16'd32495, 16'd62042, 16'd24341, 16'd27868, 16'd45424, 16'd203, 16'd44142, 16'd54547});
	test_expansion(128'h6349c0ef264c70ff0c589fa3292a486d, {16'd22925, 16'd37803, 16'd28451, 16'd56233, 16'd32222, 16'd43644, 16'd30861, 16'd60321, 16'd63201, 16'd46977, 16'd11672, 16'd44470, 16'd35731, 16'd17102, 16'd20376, 16'd37254, 16'd23629, 16'd23770, 16'd28903, 16'd18917, 16'd7252, 16'd7352, 16'd51477, 16'd56940, 16'd21272, 16'd18399});
	test_expansion(128'hb75e3e41e8f148e5cc03fd8d8817bb50, {16'd10023, 16'd62210, 16'd40944, 16'd50457, 16'd58669, 16'd56114, 16'd50192, 16'd62274, 16'd18487, 16'd30050, 16'd39201, 16'd61268, 16'd61425, 16'd11347, 16'd59961, 16'd44728, 16'd2525, 16'd9851, 16'd4775, 16'd5090, 16'd61382, 16'd7115, 16'd48682, 16'd57810, 16'd36289, 16'd55373});
	test_expansion(128'h192eb1cd42408997d4cd25dcc29f7d81, {16'd21499, 16'd49269, 16'd30433, 16'd58554, 16'd36647, 16'd30894, 16'd12929, 16'd45697, 16'd19815, 16'd47787, 16'd37606, 16'd58683, 16'd8100, 16'd63567, 16'd62217, 16'd14646, 16'd13341, 16'd53842, 16'd64150, 16'd26163, 16'd35334, 16'd43447, 16'd18555, 16'd55716, 16'd7085, 16'd12363});
	test_expansion(128'h15ef3ebfef60019c2b767e6c4e19401d, {16'd49131, 16'd48552, 16'd20017, 16'd44903, 16'd31925, 16'd65515, 16'd59311, 16'd35108, 16'd33902, 16'd15129, 16'd50796, 16'd41894, 16'd29037, 16'd65464, 16'd46692, 16'd59313, 16'd57258, 16'd64975, 16'd37629, 16'd36831, 16'd25930, 16'd17382, 16'd60285, 16'd18832, 16'd8268, 16'd25763});
	test_expansion(128'hce64c5368ca9c9bfc2bf601b90c7653e, {16'd13057, 16'd58445, 16'd19035, 16'd44679, 16'd29439, 16'd25266, 16'd28230, 16'd61923, 16'd17692, 16'd11090, 16'd5630, 16'd20757, 16'd27179, 16'd36619, 16'd9963, 16'd3202, 16'd53418, 16'd59132, 16'd38579, 16'd11533, 16'd4739, 16'd13895, 16'd28201, 16'd22469, 16'd49012, 16'd41588});
	test_expansion(128'hf1a596947479fb774bc70e2d196846d5, {16'd19636, 16'd47875, 16'd27130, 16'd25681, 16'd63047, 16'd62909, 16'd23700, 16'd59823, 16'd46450, 16'd19220, 16'd64192, 16'd5117, 16'd11219, 16'd26117, 16'd15498, 16'd9645, 16'd20783, 16'd60261, 16'd20903, 16'd1256, 16'd52498, 16'd56250, 16'd45195, 16'd17453, 16'd62011, 16'd5493});
	test_expansion(128'h6245a4c0246e44c878752c78c5f84680, {16'd38634, 16'd16164, 16'd23076, 16'd29389, 16'd56326, 16'd49060, 16'd18603, 16'd2326, 16'd43393, 16'd47335, 16'd53152, 16'd54600, 16'd34842, 16'd13017, 16'd35278, 16'd39786, 16'd63758, 16'd15295, 16'd38657, 16'd58504, 16'd16378, 16'd48869, 16'd40886, 16'd33697, 16'd59307, 16'd32375});
	test_expansion(128'h7f4c660fb9635493e23b636d3a9c5f28, {16'd32886, 16'd41309, 16'd2863, 16'd8288, 16'd32865, 16'd59834, 16'd37606, 16'd11224, 16'd38193, 16'd22265, 16'd31709, 16'd27208, 16'd9942, 16'd26407, 16'd11778, 16'd52475, 16'd35742, 16'd63376, 16'd26240, 16'd62707, 16'd24333, 16'd403, 16'd56185, 16'd6283, 16'd30080, 16'd3331});
	test_expansion(128'h0c0a63b6a12987dcc913a38b47a226b5, {16'd23558, 16'd33394, 16'd14994, 16'd12128, 16'd49827, 16'd7051, 16'd24611, 16'd59196, 16'd15006, 16'd36440, 16'd45599, 16'd50126, 16'd9016, 16'd2158, 16'd6694, 16'd16461, 16'd56697, 16'd1285, 16'd22857, 16'd6508, 16'd26551, 16'd20783, 16'd3804, 16'd61061, 16'd42675, 16'd60448});
	test_expansion(128'h8cb45a54f001c0d60c63c2d418d9633f, {16'd57299, 16'd31469, 16'd8901, 16'd50979, 16'd38217, 16'd46230, 16'd14422, 16'd39774, 16'd32673, 16'd3440, 16'd47811, 16'd55327, 16'd7311, 16'd29177, 16'd33681, 16'd19723, 16'd33009, 16'd11580, 16'd13510, 16'd28155, 16'd14399, 16'd45056, 16'd46294, 16'd9920, 16'd3350, 16'd28061});
	test_expansion(128'h32f15877d5f8d1f9a0849049a9c4c0be, {16'd20107, 16'd55725, 16'd27098, 16'd1114, 16'd52612, 16'd52970, 16'd37042, 16'd34081, 16'd48885, 16'd43043, 16'd16607, 16'd24232, 16'd43214, 16'd37789, 16'd50694, 16'd4986, 16'd55881, 16'd58098, 16'd18326, 16'd53244, 16'd10153, 16'd53934, 16'd21601, 16'd14053, 16'd16954, 16'd17901});
	test_expansion(128'h45c39900fd6dc2ae8fe50c634b7cb7fc, {16'd6726, 16'd40416, 16'd56672, 16'd53442, 16'd30606, 16'd22396, 16'd50110, 16'd64823, 16'd43788, 16'd32569, 16'd45320, 16'd29982, 16'd39414, 16'd31957, 16'd43957, 16'd21064, 16'd30723, 16'd6987, 16'd2800, 16'd49857, 16'd12349, 16'd18042, 16'd53137, 16'd50158, 16'd40653, 16'd58139});
	test_expansion(128'h7ecec1532271ed9b81811aaa5cf86796, {16'd22669, 16'd5458, 16'd57404, 16'd52820, 16'd38911, 16'd6917, 16'd35418, 16'd29331, 16'd59345, 16'd26904, 16'd20027, 16'd5837, 16'd27355, 16'd33255, 16'd62248, 16'd3063, 16'd24764, 16'd5766, 16'd54939, 16'd2003, 16'd38698, 16'd24799, 16'd18102, 16'd1039, 16'd38682, 16'd16445});
	test_expansion(128'ha330cff6e30c5a51e9569c1c6ddee314, {16'd18534, 16'd38573, 16'd34401, 16'd37324, 16'd12488, 16'd54003, 16'd40975, 16'd37318, 16'd35225, 16'd62998, 16'd16212, 16'd42434, 16'd18614, 16'd52322, 16'd24481, 16'd35935, 16'd45716, 16'd1185, 16'd47171, 16'd23915, 16'd53590, 16'd47420, 16'd3279, 16'd64015, 16'd1158, 16'd57576});
	test_expansion(128'h204546f002b795b14df84f17962b9c69, {16'd44585, 16'd50533, 16'd44255, 16'd1583, 16'd58471, 16'd42980, 16'd40228, 16'd6081, 16'd48249, 16'd8344, 16'd8672, 16'd60709, 16'd20090, 16'd11653, 16'd14150, 16'd11848, 16'd37682, 16'd34413, 16'd61499, 16'd55815, 16'd21356, 16'd45985, 16'd10939, 16'd31940, 16'd6591, 16'd7486});
	test_expansion(128'h1ef0b76d8b2858ba08adb7734c6814c8, {16'd50600, 16'd46633, 16'd15682, 16'd10821, 16'd54426, 16'd54644, 16'd31581, 16'd57009, 16'd18654, 16'd5253, 16'd61555, 16'd40247, 16'd50455, 16'd40471, 16'd59959, 16'd54576, 16'd26248, 16'd12481, 16'd34781, 16'd64030, 16'd49014, 16'd53538, 16'd26077, 16'd36349, 16'd53971, 16'd48694});
	test_expansion(128'hf8c298c64eda7f87388f0b765076b6e4, {16'd59581, 16'd53720, 16'd3497, 16'd49181, 16'd54536, 16'd18004, 16'd48323, 16'd33017, 16'd36197, 16'd28935, 16'd6691, 16'd39440, 16'd30290, 16'd14780, 16'd47426, 16'd20052, 16'd55430, 16'd41296, 16'd8396, 16'd49710, 16'd11287, 16'd9991, 16'd19954, 16'd52016, 16'd45053, 16'd46640});
	test_expansion(128'hba5ab735cc654769526d41f295644f63, {16'd46635, 16'd19292, 16'd48651, 16'd56607, 16'd64761, 16'd32662, 16'd36697, 16'd2125, 16'd6612, 16'd42902, 16'd36821, 16'd12430, 16'd63628, 16'd55099, 16'd6732, 16'd61217, 16'd34528, 16'd2680, 16'd15834, 16'd57093, 16'd59738, 16'd48454, 16'd5743, 16'd36134, 16'd17010, 16'd10817});
	test_expansion(128'h491c331b136776a6eedb9208d70ac394, {16'd1696, 16'd21864, 16'd4478, 16'd60520, 16'd64625, 16'd24341, 16'd45632, 16'd33503, 16'd44533, 16'd6797, 16'd62816, 16'd52997, 16'd46061, 16'd41103, 16'd57650, 16'd9012, 16'd1496, 16'd20061, 16'd205, 16'd14804, 16'd62848, 16'd41579, 16'd932, 16'd26945, 16'd24085, 16'd27866});
	test_expansion(128'h68ded06d50eef706ff6b320429c1a432, {16'd28448, 16'd56717, 16'd9190, 16'd42050, 16'd19370, 16'd38021, 16'd32451, 16'd19478, 16'd24772, 16'd5855, 16'd33587, 16'd7395, 16'd25351, 16'd50420, 16'd44424, 16'd3520, 16'd44579, 16'd21919, 16'd37568, 16'd5450, 16'd5387, 16'd9158, 16'd65142, 16'd31061, 16'd47155, 16'd47972});
	test_expansion(128'hf0179e9dc2c805cea5a055a2d4d942dc, {16'd54533, 16'd37792, 16'd51542, 16'd14466, 16'd47187, 16'd59307, 16'd4870, 16'd40752, 16'd31583, 16'd54648, 16'd27656, 16'd25557, 16'd49566, 16'd63061, 16'd11904, 16'd21638, 16'd17210, 16'd48420, 16'd54952, 16'd60824, 16'd41910, 16'd35528, 16'd13206, 16'd45623, 16'd10167, 16'd57813});
	test_expansion(128'h0eb38aa35aa8b31f9aaa7a36b651373f, {16'd25169, 16'd1299, 16'd51541, 16'd9510, 16'd54711, 16'd51547, 16'd16732, 16'd46671, 16'd11918, 16'd33994, 16'd26632, 16'd58525, 16'd56807, 16'd7111, 16'd32821, 16'd45163, 16'd16828, 16'd45658, 16'd43021, 16'd39662, 16'd26613, 16'd21751, 16'd50260, 16'd45976, 16'd6249, 16'd46742});
	test_expansion(128'h61c7c9c2f21451cf6af7fa356958a600, {16'd59370, 16'd52021, 16'd42516, 16'd40474, 16'd27395, 16'd54292, 16'd62167, 16'd25999, 16'd32504, 16'd34845, 16'd65227, 16'd53999, 16'd13201, 16'd28244, 16'd46358, 16'd6340, 16'd20963, 16'd18387, 16'd7013, 16'd52338, 16'd1764, 16'd34601, 16'd10844, 16'd30799, 16'd15494, 16'd27381});
	test_expansion(128'hb40a983a2a6439104ec14d49187f41c4, {16'd24039, 16'd14551, 16'd9066, 16'd26061, 16'd62971, 16'd36483, 16'd40786, 16'd52122, 16'd7945, 16'd31213, 16'd46847, 16'd3638, 16'd43060, 16'd783, 16'd64695, 16'd57679, 16'd1100, 16'd54441, 16'd6514, 16'd57846, 16'd62054, 16'd56541, 16'd63158, 16'd2537, 16'd44937, 16'd19238});
	test_expansion(128'he5d49db8cfb796f7040773a3fc18bc10, {16'd27533, 16'd13847, 16'd15514, 16'd46233, 16'd31667, 16'd10400, 16'd23588, 16'd17470, 16'd38131, 16'd26740, 16'd36387, 16'd1344, 16'd35934, 16'd59289, 16'd43896, 16'd40474, 16'd56498, 16'd61282, 16'd15652, 16'd49988, 16'd21678, 16'd36183, 16'd570, 16'd30372, 16'd24617, 16'd15997});
	test_expansion(128'h267a8915fe684af3f3e191840a368536, {16'd61387, 16'd39426, 16'd6139, 16'd47302, 16'd60050, 16'd15462, 16'd1143, 16'd26340, 16'd54585, 16'd37276, 16'd28640, 16'd31698, 16'd55440, 16'd57881, 16'd39665, 16'd41219, 16'd31943, 16'd53250, 16'd23608, 16'd64717, 16'd51200, 16'd9190, 16'd25874, 16'd43406, 16'd43791, 16'd26760});
	test_expansion(128'h970920ad2f0b0428cc96462c60e15f75, {16'd62970, 16'd15030, 16'd45829, 16'd38519, 16'd48971, 16'd12716, 16'd19723, 16'd38269, 16'd47056, 16'd37174, 16'd48843, 16'd12080, 16'd7286, 16'd50333, 16'd64534, 16'd51401, 16'd37178, 16'd12929, 16'd262, 16'd22043, 16'd63052, 16'd11156, 16'd4644, 16'd35629, 16'd9369, 16'd63366});
	test_expansion(128'ha2a5954559c1b35e377aec44ca759256, {16'd26753, 16'd17510, 16'd42470, 16'd38998, 16'd40218, 16'd18950, 16'd35878, 16'd44348, 16'd27504, 16'd4338, 16'd58041, 16'd40468, 16'd8823, 16'd33655, 16'd17042, 16'd1857, 16'd23299, 16'd19474, 16'd25776, 16'd42260, 16'd5405, 16'd56677, 16'd12845, 16'd46505, 16'd35997, 16'd48938});
	test_expansion(128'he9e2dca1bffc309eaa2ecc3d7af7863d, {16'd30224, 16'd13704, 16'd55640, 16'd54931, 16'd42102, 16'd41221, 16'd16369, 16'd3455, 16'd61829, 16'd3316, 16'd42765, 16'd34702, 16'd12992, 16'd20936, 16'd38459, 16'd24942, 16'd8775, 16'd33870, 16'd57932, 16'd25493, 16'd47488, 16'd34773, 16'd65235, 16'd53982, 16'd22760, 16'd33137});
	test_expansion(128'h254ba2431818ac7a5e9a519835f31094, {16'd56684, 16'd58635, 16'd41982, 16'd63382, 16'd4343, 16'd59190, 16'd22360, 16'd42048, 16'd57372, 16'd65519, 16'd56460, 16'd11448, 16'd33325, 16'd41455, 16'd20202, 16'd48519, 16'd41451, 16'd15974, 16'd22158, 16'd53265, 16'd224, 16'd18639, 16'd22946, 16'd57248, 16'd8896, 16'd38054});
	test_expansion(128'h51cee8700132ca49c7d96eb677661e0a, {16'd40369, 16'd53546, 16'd17641, 16'd38094, 16'd52977, 16'd62557, 16'd12868, 16'd22461, 16'd27453, 16'd54967, 16'd61242, 16'd33113, 16'd23244, 16'd18641, 16'd42803, 16'd34970, 16'd10247, 16'd30629, 16'd61475, 16'd4342, 16'd15229, 16'd51168, 16'd12872, 16'd1370, 16'd32912, 16'd27843});
	test_expansion(128'h0ebb2c70d7a732dfa403bac56b6b42b4, {16'd39346, 16'd54981, 16'd6877, 16'd56532, 16'd65280, 16'd46968, 16'd16106, 16'd45317, 16'd5074, 16'd50462, 16'd36454, 16'd17712, 16'd33377, 16'd3208, 16'd55366, 16'd13795, 16'd40382, 16'd27569, 16'd10407, 16'd21491, 16'd24259, 16'd17750, 16'd22029, 16'd11031, 16'd63328, 16'd7179});
	test_expansion(128'heb677fbca44217d1d671b546ae404258, {16'd41278, 16'd11677, 16'd10098, 16'd6452, 16'd57299, 16'd27802, 16'd37489, 16'd25802, 16'd10822, 16'd9590, 16'd34051, 16'd19274, 16'd37018, 16'd60375, 16'd42569, 16'd52997, 16'd52962, 16'd47574, 16'd10268, 16'd26818, 16'd55075, 16'd62179, 16'd22641, 16'd15587, 16'd21166, 16'd62440});
	test_expansion(128'hf54cd91a2f9f1045e347c92681871a5a, {16'd55172, 16'd23471, 16'd797, 16'd57000, 16'd18853, 16'd29576, 16'd5439, 16'd61949, 16'd926, 16'd63993, 16'd29440, 16'd41599, 16'd8995, 16'd10295, 16'd16550, 16'd2748, 16'd33247, 16'd54370, 16'd14717, 16'd63142, 16'd15765, 16'd36640, 16'd12986, 16'd18486, 16'd29145, 16'd27676});
	test_expansion(128'h0dcd67bf7b25b31472f1d6a122bafd39, {16'd52943, 16'd27621, 16'd44614, 16'd27646, 16'd28261, 16'd1325, 16'd36166, 16'd50172, 16'd38441, 16'd32492, 16'd30141, 16'd45479, 16'd11054, 16'd37952, 16'd51410, 16'd4736, 16'd16726, 16'd31679, 16'd24868, 16'd12206, 16'd21287, 16'd49094, 16'd59074, 16'd19673, 16'd13734, 16'd32121});
	test_expansion(128'h1f4c87f38f13fa8862f480f37fd77b64, {16'd2585, 16'd58302, 16'd59066, 16'd65307, 16'd59983, 16'd58020, 16'd4300, 16'd2560, 16'd44504, 16'd36266, 16'd6695, 16'd46982, 16'd27185, 16'd1699, 16'd54383, 16'd36285, 16'd2680, 16'd36300, 16'd49546, 16'd11400, 16'd1976, 16'd9258, 16'd26812, 16'd47244, 16'd26700, 16'd18879});
	test_expansion(128'hf1de1599c088787726512fbff0aebaae, {16'd57718, 16'd63315, 16'd44591, 16'd59230, 16'd29466, 16'd5283, 16'd29236, 16'd56445, 16'd25707, 16'd28186, 16'd49584, 16'd7456, 16'd27546, 16'd51309, 16'd55101, 16'd61344, 16'd38939, 16'd26093, 16'd34752, 16'd34769, 16'd41157, 16'd32625, 16'd11814, 16'd20926, 16'd53514, 16'd16547});
	test_expansion(128'h5630370efc8a94da8c8824babbfbccea, {16'd28986, 16'd4329, 16'd14127, 16'd33718, 16'd19162, 16'd17442, 16'd63247, 16'd30854, 16'd40778, 16'd4249, 16'd37382, 16'd28801, 16'd52321, 16'd58682, 16'd14517, 16'd55966, 16'd14075, 16'd6182, 16'd2564, 16'd26060, 16'd65281, 16'd30557, 16'd29893, 16'd55595, 16'd3125, 16'd24121});
	test_expansion(128'h38960011ae8c72d7429d84a0702e204e, {16'd37827, 16'd35827, 16'd12052, 16'd11389, 16'd18260, 16'd40619, 16'd62679, 16'd13914, 16'd29723, 16'd53531, 16'd18276, 16'd47355, 16'd61843, 16'd27747, 16'd23397, 16'd53900, 16'd44595, 16'd2353, 16'd62825, 16'd59324, 16'd43707, 16'd61334, 16'd10200, 16'd19104, 16'd23563, 16'd7282});
	test_expansion(128'h911bb0915af7311b408bfd53ba0433e8, {16'd32891, 16'd28724, 16'd15543, 16'd30493, 16'd48502, 16'd62043, 16'd64992, 16'd25174, 16'd33398, 16'd24745, 16'd2892, 16'd15152, 16'd13076, 16'd7562, 16'd39842, 16'd49270, 16'd59089, 16'd64813, 16'd51366, 16'd46470, 16'd51705, 16'd40296, 16'd41414, 16'd51536, 16'd28041, 16'd39534});
	test_expansion(128'h8495a471ad86653fb3208ada88390c89, {16'd13497, 16'd27988, 16'd6044, 16'd52667, 16'd19585, 16'd22150, 16'd1560, 16'd15093, 16'd120, 16'd37771, 16'd3464, 16'd35587, 16'd49066, 16'd32598, 16'd37558, 16'd51642, 16'd48133, 16'd18531, 16'd1240, 16'd13500, 16'd7636, 16'd31776, 16'd52526, 16'd36120, 16'd45595, 16'd7238});
	test_expansion(128'hbf6d641db37c7e0aa026414643ed8018, {16'd6927, 16'd14827, 16'd62315, 16'd27393, 16'd39820, 16'd43472, 16'd12208, 16'd43729, 16'd61800, 16'd11350, 16'd25483, 16'd18315, 16'd21366, 16'd3084, 16'd58124, 16'd12005, 16'd25764, 16'd14221, 16'd27497, 16'd14143, 16'd64904, 16'd34199, 16'd36687, 16'd58009, 16'd28543, 16'd4019});
	test_expansion(128'hf60865fc97f1496eaca22cec81e11a0f, {16'd47328, 16'd36700, 16'd40216, 16'd23295, 16'd58949, 16'd24941, 16'd26031, 16'd15190, 16'd41416, 16'd9009, 16'd32816, 16'd51261, 16'd346, 16'd60087, 16'd22911, 16'd13406, 16'd53110, 16'd38994, 16'd15405, 16'd36774, 16'd17187, 16'd27585, 16'd45663, 16'd3748, 16'd23961, 16'd16761});
	test_expansion(128'hc158d2fc5483856b0b908c23ca566b12, {16'd2093, 16'd47037, 16'd27579, 16'd54367, 16'd46605, 16'd59913, 16'd42377, 16'd1596, 16'd58976, 16'd10861, 16'd60553, 16'd12487, 16'd20699, 16'd47535, 16'd30079, 16'd61589, 16'd50876, 16'd11443, 16'd61974, 16'd49736, 16'd12554, 16'd37972, 16'd463, 16'd61369, 16'd17077, 16'd40605});
	test_expansion(128'h1d269f8354af8999a976b7c2f2014db1, {16'd26264, 16'd28749, 16'd38263, 16'd11315, 16'd50972, 16'd39258, 16'd18889, 16'd46548, 16'd58141, 16'd48359, 16'd29116, 16'd36587, 16'd31820, 16'd31648, 16'd17043, 16'd146, 16'd37754, 16'd21949, 16'd10874, 16'd28605, 16'd15912, 16'd45562, 16'd35765, 16'd58375, 16'd53784, 16'd32400});
	test_expansion(128'h9964f869acbbdaae30f42bc481c91edf, {16'd60603, 16'd6177, 16'd12518, 16'd16445, 16'd34949, 16'd17667, 16'd15799, 16'd769, 16'd41334, 16'd3222, 16'd39040, 16'd3847, 16'd1121, 16'd45498, 16'd29424, 16'd23976, 16'd13501, 16'd25173, 16'd43016, 16'd51946, 16'd29745, 16'd28731, 16'd52698, 16'd3849, 16'd54243, 16'd11777});
	test_expansion(128'h127d411ec81f767049d9095929727c93, {16'd14121, 16'd39126, 16'd6060, 16'd48296, 16'd14531, 16'd12543, 16'd36643, 16'd51834, 16'd1331, 16'd26530, 16'd64776, 16'd51403, 16'd22040, 16'd22862, 16'd42954, 16'd225, 16'd5105, 16'd10646, 16'd17927, 16'd17220, 16'd61571, 16'd43974, 16'd13893, 16'd54692, 16'd34068, 16'd16581});
	test_expansion(128'h66eded4142843995f2d6d59752a4cec7, {16'd30417, 16'd18803, 16'd17421, 16'd6469, 16'd40873, 16'd55410, 16'd28514, 16'd64490, 16'd8, 16'd20204, 16'd21772, 16'd28630, 16'd4660, 16'd40101, 16'd2340, 16'd24159, 16'd26186, 16'd9107, 16'd33877, 16'd7851, 16'd30540, 16'd17378, 16'd55795, 16'd3194, 16'd26578, 16'd3896});
	test_expansion(128'h94e05c48fa915814d9fbd6d5bd9407dc, {16'd22528, 16'd36114, 16'd31199, 16'd55315, 16'd55266, 16'd34276, 16'd19919, 16'd40115, 16'd7996, 16'd20244, 16'd11660, 16'd44276, 16'd30534, 16'd32606, 16'd45803, 16'd38270, 16'd40088, 16'd53528, 16'd15940, 16'd1068, 16'd8976, 16'd23644, 16'd1644, 16'd4598, 16'd46855, 16'd57815});
	test_expansion(128'h6616394e485bcbdbed980ccebae64f27, {16'd49860, 16'd61935, 16'd26201, 16'd52378, 16'd30285, 16'd32813, 16'd850, 16'd39477, 16'd17883, 16'd52329, 16'd40971, 16'd17409, 16'd7930, 16'd63997, 16'd10811, 16'd58705, 16'd32060, 16'd58144, 16'd64668, 16'd32227, 16'd12883, 16'd21507, 16'd36927, 16'd19107, 16'd18870, 16'd50521});
	test_expansion(128'h845029cd7fce6f92fd242431f3d0ec78, {16'd24329, 16'd18226, 16'd24679, 16'd20204, 16'd49357, 16'd50774, 16'd39041, 16'd16541, 16'd53759, 16'd26354, 16'd64232, 16'd60321, 16'd63683, 16'd29530, 16'd10975, 16'd54280, 16'd50542, 16'd44123, 16'd62289, 16'd23083, 16'd8825, 16'd62078, 16'd52736, 16'd23467, 16'd47034, 16'd36542});
	test_expansion(128'h1c2a382d195b05f6f92eace47fa202e4, {16'd35011, 16'd59528, 16'd6158, 16'd52722, 16'd34760, 16'd26844, 16'd37782, 16'd32304, 16'd11039, 16'd2473, 16'd47700, 16'd8715, 16'd6664, 16'd348, 16'd60560, 16'd61051, 16'd64442, 16'd6254, 16'd56744, 16'd47352, 16'd41832, 16'd10799, 16'd17496, 16'd49322, 16'd61919, 16'd42338});
	test_expansion(128'h5b3df3433f81ef7be602bd2d3119ba9d, {16'd51493, 16'd36615, 16'd4846, 16'd7208, 16'd8965, 16'd57932, 16'd24565, 16'd63366, 16'd64681, 16'd7457, 16'd54360, 16'd43446, 16'd46032, 16'd42270, 16'd5501, 16'd44172, 16'd19328, 16'd45720, 16'd35219, 16'd49693, 16'd17127, 16'd29241, 16'd30777, 16'd9777, 16'd27640, 16'd56238});
	test_expansion(128'h9d8bdc61876c0d7d856451fcf035ce9c, {16'd18132, 16'd42790, 16'd1500, 16'd4071, 16'd13123, 16'd43059, 16'd42307, 16'd54130, 16'd29064, 16'd53421, 16'd33259, 16'd46567, 16'd40566, 16'd56447, 16'd41705, 16'd55252, 16'd27297, 16'd59972, 16'd52999, 16'd47012, 16'd35557, 16'd6593, 16'd36531, 16'd45581, 16'd44674, 16'd57497});
	test_expansion(128'hb272efc03cadb0de2d475c2692d07186, {16'd63018, 16'd52863, 16'd38654, 16'd59238, 16'd42633, 16'd40110, 16'd24450, 16'd2793, 16'd17267, 16'd26040, 16'd43355, 16'd11097, 16'd65304, 16'd9858, 16'd58386, 16'd50049, 16'd32243, 16'd15180, 16'd7456, 16'd60907, 16'd54469, 16'd13679, 16'd51994, 16'd53436, 16'd34930, 16'd4833});
	test_expansion(128'hd985b9871d1c9b2b7718e13ac9ace3df, {16'd46153, 16'd54326, 16'd18704, 16'd45194, 16'd17649, 16'd2106, 16'd54193, 16'd17084, 16'd22417, 16'd51509, 16'd22360, 16'd25448, 16'd42894, 16'd22984, 16'd12599, 16'd11664, 16'd6025, 16'd7847, 16'd23403, 16'd1599, 16'd36174, 16'd7990, 16'd57237, 16'd13702, 16'd30553, 16'd40934});
	test_expansion(128'hbcc3f7a3107c884c4861b2e5a67b0ed5, {16'd20252, 16'd45300, 16'd29022, 16'd59420, 16'd38552, 16'd55061, 16'd21463, 16'd2940, 16'd32567, 16'd19262, 16'd61148, 16'd29416, 16'd50720, 16'd7179, 16'd49828, 16'd42846, 16'd6683, 16'd9632, 16'd3289, 16'd14788, 16'd16429, 16'd56945, 16'd40747, 16'd27178, 16'd59141, 16'd30949});
	test_expansion(128'h54974da30ef8959bbe4984a06a09d832, {16'd65500, 16'd32615, 16'd49798, 16'd14949, 16'd62012, 16'd58995, 16'd13620, 16'd44580, 16'd50426, 16'd20123, 16'd17888, 16'd55753, 16'd46023, 16'd41708, 16'd62112, 16'd2818, 16'd53908, 16'd31489, 16'd25841, 16'd40404, 16'd19816, 16'd29976, 16'd53657, 16'd48943, 16'd38835, 16'd1456});
	test_expansion(128'h4e9c9d62ea750d0229d9f29b5de35a43, {16'd30891, 16'd34017, 16'd768, 16'd7213, 16'd41758, 16'd45531, 16'd58903, 16'd51497, 16'd4321, 16'd9168, 16'd8471, 16'd54545, 16'd2206, 16'd6062, 16'd41516, 16'd13642, 16'd43482, 16'd48148, 16'd45232, 16'd7455, 16'd63723, 16'd32483, 16'd52785, 16'd13590, 16'd44594, 16'd3874});
	test_expansion(128'h29914037c3259503d476e557201a02d7, {16'd37135, 16'd53422, 16'd49794, 16'd64816, 16'd35800, 16'd1541, 16'd54191, 16'd3837, 16'd12081, 16'd24067, 16'd25546, 16'd59043, 16'd30457, 16'd19966, 16'd1790, 16'd63135, 16'd41425, 16'd57299, 16'd60696, 16'd42756, 16'd35477, 16'd24533, 16'd36731, 16'd59568, 16'd37679, 16'd17122});
	test_expansion(128'h78953974473db24ea5c002f23f120f5d, {16'd15851, 16'd28921, 16'd61100, 16'd22339, 16'd1165, 16'd4854, 16'd41274, 16'd26709, 16'd3046, 16'd44924, 16'd6798, 16'd20044, 16'd10833, 16'd12226, 16'd16544, 16'd41656, 16'd29743, 16'd59343, 16'd33906, 16'd57776, 16'd30088, 16'd39573, 16'd2244, 16'd59725, 16'd31960, 16'd49333});
	test_expansion(128'h23b7464535f3ff877dfd5f68cbe76b22, {16'd36169, 16'd9473, 16'd16473, 16'd50074, 16'd15542, 16'd26453, 16'd4309, 16'd43548, 16'd48094, 16'd15128, 16'd28766, 16'd64464, 16'd29473, 16'd3550, 16'd59206, 16'd44910, 16'd60418, 16'd24716, 16'd21694, 16'd10808, 16'd27583, 16'd61515, 16'd12443, 16'd31156, 16'd42145, 16'd64087});
	test_expansion(128'hb5901ec5ba0cf8c11252a45552bb8b52, {16'd58224, 16'd28090, 16'd53468, 16'd31368, 16'd39883, 16'd53790, 16'd30474, 16'd13695, 16'd63863, 16'd10681, 16'd59534, 16'd63231, 16'd20874, 16'd11572, 16'd61540, 16'd38190, 16'd4557, 16'd18758, 16'd4872, 16'd28446, 16'd15179, 16'd14987, 16'd9762, 16'd36672, 16'd29791, 16'd51662});
	test_expansion(128'h453ffe27692900d73c3792509f383ca3, {16'd64501, 16'd56786, 16'd28956, 16'd53832, 16'd7568, 16'd60568, 16'd54321, 16'd30586, 16'd7802, 16'd32128, 16'd23441, 16'd43158, 16'd24808, 16'd21632, 16'd21576, 16'd32977, 16'd54694, 16'd35055, 16'd19223, 16'd13492, 16'd35262, 16'd11998, 16'd44506, 16'd52979, 16'd45075, 16'd14615});
	test_expansion(128'h0ce932b7784a6dc6b10cedcc4ee8313e, {16'd33073, 16'd6982, 16'd3100, 16'd14582, 16'd6252, 16'd53770, 16'd56413, 16'd48079, 16'd38211, 16'd17996, 16'd26196, 16'd21382, 16'd17608, 16'd58022, 16'd58483, 16'd51558, 16'd49852, 16'd64655, 16'd4165, 16'd45370, 16'd4456, 16'd20688, 16'd64691, 16'd31763, 16'd57577, 16'd54820});
	test_expansion(128'h896765f76198a90ecad414e130b09e31, {16'd38114, 16'd1038, 16'd54778, 16'd8645, 16'd31902, 16'd12545, 16'd12595, 16'd29247, 16'd1180, 16'd65177, 16'd51452, 16'd10226, 16'd19560, 16'd7692, 16'd6025, 16'd50643, 16'd53033, 16'd26159, 16'd65419, 16'd35803, 16'd52076, 16'd54523, 16'd23889, 16'd38401, 16'd52173, 16'd9959});
	test_expansion(128'h78047ac31c6e06f98ab9b09abdecc125, {16'd46471, 16'd23848, 16'd45913, 16'd3324, 16'd40781, 16'd26253, 16'd12536, 16'd33721, 16'd18971, 16'd6685, 16'd12480, 16'd40066, 16'd58932, 16'd32116, 16'd37900, 16'd10139, 16'd60436, 16'd48245, 16'd63328, 16'd62247, 16'd19774, 16'd56730, 16'd38672, 16'd56545, 16'd54940, 16'd52502});
	test_expansion(128'h102168055ec50b7699203f39b9e6c6d1, {16'd50497, 16'd60029, 16'd4784, 16'd5450, 16'd14869, 16'd62314, 16'd28250, 16'd38429, 16'd52709, 16'd56858, 16'd5824, 16'd30233, 16'd16572, 16'd15912, 16'd39086, 16'd42582, 16'd45552, 16'd24339, 16'd23283, 16'd35537, 16'd30420, 16'd35883, 16'd869, 16'd18980, 16'd43872, 16'd16260});
	test_expansion(128'h414c4b77418196fba68efd2f3c0b2bbf, {16'd49076, 16'd10412, 16'd54722, 16'd34440, 16'd24003, 16'd33796, 16'd60474, 16'd25665, 16'd5898, 16'd40328, 16'd63307, 16'd7718, 16'd42193, 16'd26602, 16'd19709, 16'd63730, 16'd26534, 16'd28136, 16'd401, 16'd37077, 16'd42343, 16'd5025, 16'd32525, 16'd57532, 16'd2189, 16'd35498});
	test_expansion(128'h871513e0fbba65ed70d2dc9674478311, {16'd2863, 16'd64939, 16'd31320, 16'd31917, 16'd59569, 16'd38280, 16'd174, 16'd59258, 16'd31507, 16'd55028, 16'd17545, 16'd50207, 16'd23921, 16'd35066, 16'd54660, 16'd50869, 16'd26790, 16'd9774, 16'd17137, 16'd8304, 16'd62891, 16'd25513, 16'd2325, 16'd58970, 16'd9829, 16'd29622});
	test_expansion(128'h4a9fb0579589d378523eb1641cd88252, {16'd21951, 16'd5099, 16'd48, 16'd34220, 16'd55135, 16'd8706, 16'd4621, 16'd3619, 16'd54002, 16'd44042, 16'd23206, 16'd42160, 16'd60241, 16'd44697, 16'd51277, 16'd23455, 16'd2020, 16'd35738, 16'd51249, 16'd55464, 16'd53805, 16'd58601, 16'd2704, 16'd35021, 16'd39616, 16'd46666});
	test_expansion(128'h3b7a80f5dd8a602bd4f667b19df066c8, {16'd49980, 16'd65343, 16'd45065, 16'd41526, 16'd22569, 16'd46497, 16'd28102, 16'd13920, 16'd62052, 16'd29185, 16'd60916, 16'd44686, 16'd5028, 16'd7149, 16'd63756, 16'd22517, 16'd41716, 16'd10022, 16'd3393, 16'd30751, 16'd19050, 16'd26983, 16'd41518, 16'd41817, 16'd46725, 16'd40471});
	test_expansion(128'h5890aa4ffc4746b7c1ba75b4fcd8ce61, {16'd320, 16'd50698, 16'd20384, 16'd11464, 16'd40987, 16'd59221, 16'd17646, 16'd51758, 16'd34127, 16'd20623, 16'd46731, 16'd18874, 16'd36754, 16'd41162, 16'd14317, 16'd61925, 16'd20523, 16'd62843, 16'd61452, 16'd15149, 16'd1053, 16'd62010, 16'd29963, 16'd2193, 16'd19625, 16'd24809});
	test_expansion(128'hddf1c7b4a703876dd8177bd3f5235351, {16'd46521, 16'd31293, 16'd9296, 16'd58130, 16'd63466, 16'd11075, 16'd57246, 16'd47662, 16'd30316, 16'd3224, 16'd64780, 16'd56327, 16'd58050, 16'd41249, 16'd18565, 16'd12476, 16'd34321, 16'd44132, 16'd19619, 16'd35123, 16'd7932, 16'd54135, 16'd24058, 16'd54546, 16'd8661, 16'd30895});
	test_expansion(128'hbe917add6b77cbd1159a056a69f7b39f, {16'd3785, 16'd20333, 16'd65378, 16'd11175, 16'd34010, 16'd42137, 16'd37972, 16'd15543, 16'd37445, 16'd25496, 16'd26658, 16'd53226, 16'd22510, 16'd325, 16'd17332, 16'd52080, 16'd51455, 16'd49796, 16'd18452, 16'd9166, 16'd57591, 16'd47900, 16'd23674, 16'd57133, 16'd48737, 16'd18435});
	test_expansion(128'h6e36a20a4d3cd598a2e4628a83ec478a, {16'd48417, 16'd17652, 16'd60394, 16'd52144, 16'd52975, 16'd30901, 16'd21912, 16'd33033, 16'd56607, 16'd49578, 16'd29876, 16'd34278, 16'd42214, 16'd29319, 16'd13866, 16'd48834, 16'd27204, 16'd32722, 16'd5343, 16'd41296, 16'd13273, 16'd44626, 16'd17071, 16'd36170, 16'd57597, 16'd43892});
	test_expansion(128'hc70e957f74a3aad4d3b4b0d954f25a24, {16'd65029, 16'd58137, 16'd29354, 16'd19055, 16'd54436, 16'd31720, 16'd57166, 16'd41991, 16'd55552, 16'd6985, 16'd46681, 16'd4713, 16'd60435, 16'd15499, 16'd29791, 16'd19890, 16'd18876, 16'd58005, 16'd14679, 16'd19756, 16'd40415, 16'd55348, 16'd48009, 16'd31689, 16'd48654, 16'd15142});
	test_expansion(128'h4957e61fb89597578fae141736d3a085, {16'd27874, 16'd9196, 16'd38360, 16'd16597, 16'd18440, 16'd35061, 16'd16785, 16'd11518, 16'd12086, 16'd41486, 16'd29898, 16'd48643, 16'd38963, 16'd3063, 16'd23250, 16'd58895, 16'd43604, 16'd8556, 16'd50962, 16'd20109, 16'd57754, 16'd55449, 16'd37766, 16'd12336, 16'd42720, 16'd49194});
	test_expansion(128'hf1a171cbc1887da3c9001079ead0c420, {16'd22979, 16'd51585, 16'd4218, 16'd62931, 16'd13690, 16'd25407, 16'd45327, 16'd1323, 16'd28678, 16'd19812, 16'd2170, 16'd33923, 16'd18871, 16'd11920, 16'd2035, 16'd14213, 16'd8543, 16'd56932, 16'd15188, 16'd9549, 16'd60672, 16'd58651, 16'd50981, 16'd27271, 16'd41799, 16'd2851});
	test_expansion(128'he0caca0cd823c0b57ff011d9bfd94129, {16'd22197, 16'd52939, 16'd18189, 16'd29339, 16'd7784, 16'd25182, 16'd57999, 16'd31293, 16'd24668, 16'd7564, 16'd64021, 16'd32384, 16'd12383, 16'd29467, 16'd5153, 16'd57104, 16'd43940, 16'd41681, 16'd35421, 16'd28898, 16'd14924, 16'd22502, 16'd6527, 16'd53616, 16'd51711, 16'd42574});
	test_expansion(128'ha64e66cc7a4f9b6af213f50c5f43ec2b, {16'd64692, 16'd59262, 16'd25069, 16'd36975, 16'd8924, 16'd38600, 16'd52551, 16'd24418, 16'd56342, 16'd43826, 16'd47529, 16'd45243, 16'd39385, 16'd63900, 16'd49854, 16'd53985, 16'd56972, 16'd11382, 16'd55763, 16'd49729, 16'd63478, 16'd14939, 16'd57686, 16'd29873, 16'd15711, 16'd40879});
	test_expansion(128'h009a0ed79b5d4e3c122ee27281026e26, {16'd38759, 16'd48571, 16'd39192, 16'd15914, 16'd52743, 16'd13614, 16'd44049, 16'd17395, 16'd53459, 16'd3701, 16'd32622, 16'd17039, 16'd21112, 16'd19231, 16'd47384, 16'd49080, 16'd52517, 16'd10110, 16'd34854, 16'd37900, 16'd14050, 16'd9220, 16'd18146, 16'd59376, 16'd58714, 16'd37956});
	test_expansion(128'h71e72cd6e7e25f51b6bc944a25252c29, {16'd43668, 16'd62285, 16'd63829, 16'd14949, 16'd4348, 16'd4282, 16'd20075, 16'd27347, 16'd29370, 16'd46190, 16'd2913, 16'd11301, 16'd215, 16'd34253, 16'd20937, 16'd862, 16'd19815, 16'd51280, 16'd6656, 16'd59581, 16'd64664, 16'd64346, 16'd2646, 16'd50664, 16'd33048, 16'd39576});
	test_expansion(128'hf4c56a33248331e41c97d4bf32a59570, {16'd15632, 16'd19372, 16'd38870, 16'd3439, 16'd22870, 16'd34535, 16'd54108, 16'd26609, 16'd60913, 16'd924, 16'd25251, 16'd5009, 16'd25165, 16'd47673, 16'd7897, 16'd52830, 16'd41476, 16'd44640, 16'd3801, 16'd58740, 16'd43979, 16'd25323, 16'd56001, 16'd43424, 16'd28617, 16'd19992});
	test_expansion(128'hcbc4abb5920135289b9096c05bd229e6, {16'd52738, 16'd33959, 16'd14129, 16'd58697, 16'd46271, 16'd39363, 16'd51339, 16'd27075, 16'd59337, 16'd62519, 16'd2040, 16'd60104, 16'd11565, 16'd1743, 16'd4139, 16'd28536, 16'd57131, 16'd29087, 16'd39246, 16'd61543, 16'd5500, 16'd51546, 16'd6943, 16'd80, 16'd41563, 16'd43165});
	test_expansion(128'h198bb3cad9dcd6bdf695853e4f539574, {16'd53602, 16'd65347, 16'd35058, 16'd16204, 16'd13920, 16'd63429, 16'd57052, 16'd21111, 16'd46343, 16'd52816, 16'd33007, 16'd37714, 16'd47457, 16'd39263, 16'd29586, 16'd58654, 16'd43674, 16'd49941, 16'd35092, 16'd24563, 16'd13609, 16'd5858, 16'd49858, 16'd5471, 16'd32621, 16'd26899});
	test_expansion(128'he698b67eed16e1a8c3c1d1cb92d92253, {16'd33103, 16'd18572, 16'd2708, 16'd45203, 16'd6146, 16'd5179, 16'd60913, 16'd37738, 16'd50460, 16'd56642, 16'd64005, 16'd52507, 16'd62871, 16'd59791, 16'd14778, 16'd51374, 16'd20911, 16'd37333, 16'd18496, 16'd53328, 16'd42389, 16'd56037, 16'd35782, 16'd52099, 16'd18232, 16'd42172});
	test_expansion(128'heda4f2e5ba75112ad2b5b9e83398c9e6, {16'd39916, 16'd21343, 16'd61524, 16'd49591, 16'd10618, 16'd29921, 16'd22485, 16'd58875, 16'd47014, 16'd1848, 16'd37000, 16'd62521, 16'd21037, 16'd24215, 16'd51467, 16'd9051, 16'd49823, 16'd20091, 16'd59068, 16'd36576, 16'd51947, 16'd27327, 16'd64110, 16'd61586, 16'd12312, 16'd53418});
	test_expansion(128'h207c82f1c7bab914fe43c21822a3ec9e, {16'd49178, 16'd29032, 16'd43067, 16'd33426, 16'd7938, 16'd2077, 16'd18642, 16'd5217, 16'd23541, 16'd10655, 16'd59381, 16'd40237, 16'd10468, 16'd7581, 16'd19648, 16'd57739, 16'd15880, 16'd30889, 16'd13163, 16'd25624, 16'd20027, 16'd59832, 16'd46104, 16'd2956, 16'd24764, 16'd64103});
	test_expansion(128'h45c28aafaa52da10142dcbdc796ac94b, {16'd62330, 16'd6316, 16'd24504, 16'd34534, 16'd30256, 16'd53758, 16'd1770, 16'd59138, 16'd48663, 16'd62861, 16'd6935, 16'd48137, 16'd1976, 16'd36744, 16'd22434, 16'd8524, 16'd44282, 16'd13936, 16'd1499, 16'd44154, 16'd5768, 16'd7722, 16'd60674, 16'd48129, 16'd25441, 16'd13393});
	test_expansion(128'h134060564672be1d901c7cd1eb9c0873, {16'd52612, 16'd15232, 16'd47187, 16'd14017, 16'd40818, 16'd45206, 16'd8477, 16'd13920, 16'd17826, 16'd61936, 16'd7767, 16'd57252, 16'd30564, 16'd11346, 16'd12715, 16'd39653, 16'd39328, 16'd36498, 16'd32630, 16'd29812, 16'd7118, 16'd47801, 16'd49182, 16'd10212, 16'd4512, 16'd14555});
	test_expansion(128'h9f517e942e6b6a03f64b8735735969f9, {16'd9657, 16'd62208, 16'd16014, 16'd7798, 16'd11140, 16'd4737, 16'd41167, 16'd37900, 16'd63910, 16'd63878, 16'd64140, 16'd4089, 16'd6110, 16'd45807, 16'd55272, 16'd31065, 16'd16912, 16'd18492, 16'd10321, 16'd44771, 16'd34546, 16'd22301, 16'd54307, 16'd48744, 16'd45937, 16'd4383});
	test_expansion(128'h9cbe0b43986689fcfe79c794091c30a7, {16'd43094, 16'd23767, 16'd31757, 16'd32859, 16'd15709, 16'd62821, 16'd21835, 16'd247, 16'd37648, 16'd22354, 16'd17010, 16'd39079, 16'd24105, 16'd24682, 16'd8930, 16'd60795, 16'd16152, 16'd33751, 16'd13307, 16'd16223, 16'd5731, 16'd24595, 16'd8343, 16'd35270, 16'd40854, 16'd2057});
	test_expansion(128'h0a7bd651f623735b1e14e49021c1bd3d, {16'd9649, 16'd49442, 16'd27923, 16'd21651, 16'd26235, 16'd30016, 16'd37854, 16'd28027, 16'd58446, 16'd21580, 16'd3656, 16'd45374, 16'd48749, 16'd5565, 16'd21592, 16'd10117, 16'd62650, 16'd1967, 16'd34370, 16'd29259, 16'd30686, 16'd4248, 16'd19986, 16'd2825, 16'd8676, 16'd24684});
	test_expansion(128'h2a094692cad89c9c0a36c069860a345b, {16'd47180, 16'd51397, 16'd33707, 16'd53917, 16'd61567, 16'd6028, 16'd24882, 16'd52008, 16'd59550, 16'd56352, 16'd4067, 16'd37419, 16'd44633, 16'd45225, 16'd13239, 16'd42840, 16'd34125, 16'd27173, 16'd33755, 16'd36013, 16'd59724, 16'd9353, 16'd12936, 16'd13668, 16'd61457, 16'd14176});
	test_expansion(128'h8f38eb218bc699334e4eaf9030b5a2c4, {16'd12410, 16'd62991, 16'd24320, 16'd16524, 16'd2919, 16'd9560, 16'd24898, 16'd35075, 16'd57822, 16'd33779, 16'd17719, 16'd3418, 16'd4006, 16'd31810, 16'd21386, 16'd30168, 16'd2707, 16'd41140, 16'd393, 16'd9504, 16'd27522, 16'd5556, 16'd6507, 16'd7121, 16'd33766, 16'd47527});
	test_expansion(128'h34e858573b975655454367a17e1212ff, {16'd27402, 16'd11909, 16'd21680, 16'd30494, 16'd20476, 16'd41382, 16'd53975, 16'd30455, 16'd57855, 16'd49573, 16'd42588, 16'd16368, 16'd25355, 16'd42537, 16'd46313, 16'd59051, 16'd1717, 16'd29088, 16'd19579, 16'd28204, 16'd51197, 16'd12191, 16'd52079, 16'd22107, 16'd56720, 16'd2970});
	test_expansion(128'h4cd14d4d17e6c24decb1e9ee5ccb2235, {16'd59862, 16'd38258, 16'd20098, 16'd35129, 16'd24537, 16'd524, 16'd51619, 16'd13620, 16'd53429, 16'd50942, 16'd12803, 16'd58430, 16'd12788, 16'd36871, 16'd24948, 16'd13066, 16'd30751, 16'd14804, 16'd28674, 16'd34203, 16'd16643, 16'd62209, 16'd7774, 16'd16487, 16'd25351, 16'd48668});
	test_expansion(128'hb024f50ff0e2ddfb971b8bfae7343f76, {16'd55038, 16'd61616, 16'd61280, 16'd52272, 16'd12932, 16'd12198, 16'd9078, 16'd54051, 16'd43614, 16'd21278, 16'd65184, 16'd15637, 16'd4473, 16'd7133, 16'd17756, 16'd33095, 16'd14121, 16'd56835, 16'd59593, 16'd24776, 16'd28388, 16'd21869, 16'd58208, 16'd46171, 16'd22575, 16'd24779});
	test_expansion(128'h322ef494bcf664adcd1bf596ea91f5c7, {16'd47415, 16'd27251, 16'd20285, 16'd52322, 16'd32001, 16'd5347, 16'd37408, 16'd49516, 16'd15572, 16'd28048, 16'd36894, 16'd58780, 16'd9714, 16'd1237, 16'd32056, 16'd25017, 16'd23695, 16'd1398, 16'd52776, 16'd2464, 16'd29603, 16'd30490, 16'd15223, 16'd4194, 16'd43789, 16'd41689});
	test_expansion(128'h03d66e189b998c994d9f3b3038ee8ea3, {16'd57775, 16'd6096, 16'd6527, 16'd20530, 16'd8915, 16'd16133, 16'd39001, 16'd41528, 16'd16898, 16'd4547, 16'd51069, 16'd36796, 16'd39861, 16'd26233, 16'd13920, 16'd12177, 16'd25100, 16'd13069, 16'd32147, 16'd30893, 16'd52754, 16'd47920, 16'd33606, 16'd30762, 16'd45683, 16'd35605});
	test_expansion(128'h126f4bcfe0671504086fda9adec930e8, {16'd35623, 16'd34915, 16'd46997, 16'd16480, 16'd44852, 16'd41573, 16'd16079, 16'd49137, 16'd47816, 16'd26423, 16'd26675, 16'd24627, 16'd45289, 16'd45945, 16'd12505, 16'd51574, 16'd64056, 16'd45442, 16'd21318, 16'd62871, 16'd4475, 16'd40835, 16'd45612, 16'd20486, 16'd3589, 16'd41608});
	test_expansion(128'hd0a8cb7d46bff8c641bd28090a340e06, {16'd18869, 16'd1895, 16'd33133, 16'd50420, 16'd4565, 16'd29956, 16'd49039, 16'd43159, 16'd24794, 16'd43292, 16'd32731, 16'd23169, 16'd2874, 16'd26335, 16'd52631, 16'd53247, 16'd27480, 16'd58764, 16'd30526, 16'd37901, 16'd54029, 16'd6434, 16'd9775, 16'd33350, 16'd15683, 16'd14704});
	test_expansion(128'h86eca67fc2ad6336454d35818d140452, {16'd51731, 16'd26482, 16'd40261, 16'd14072, 16'd19808, 16'd4897, 16'd1905, 16'd18028, 16'd47831, 16'd62019, 16'd50106, 16'd52902, 16'd7866, 16'd25680, 16'd12780, 16'd3423, 16'd40264, 16'd44793, 16'd2639, 16'd17595, 16'd10900, 16'd13662, 16'd17492, 16'd41396, 16'd17402, 16'd64409});
	test_expansion(128'h60c638df9d597b77f0dc6b4d1dee43e3, {16'd46950, 16'd59781, 16'd22574, 16'd61408, 16'd62848, 16'd12129, 16'd14952, 16'd57, 16'd13591, 16'd34589, 16'd36253, 16'd13119, 16'd35746, 16'd27005, 16'd9668, 16'd37504, 16'd11806, 16'd5130, 16'd57062, 16'd43959, 16'd32349, 16'd56901, 16'd12895, 16'd62094, 16'd20898, 16'd5006});
	test_expansion(128'h51c7b6d81a14b8858efe33c8b50ce207, {16'd16539, 16'd24077, 16'd7272, 16'd59213, 16'd33247, 16'd14595, 16'd29862, 16'd33793, 16'd8031, 16'd41842, 16'd32104, 16'd8002, 16'd23052, 16'd27434, 16'd35102, 16'd33116, 16'd17015, 16'd62612, 16'd25669, 16'd41704, 16'd60470, 16'd17941, 16'd15905, 16'd25428, 16'd23291, 16'd21662});
	test_expansion(128'h476a93a38dd85b098a812fbf79a12f6b, {16'd54637, 16'd33432, 16'd15941, 16'd1701, 16'd10038, 16'd6380, 16'd61828, 16'd39138, 16'd36636, 16'd45353, 16'd54029, 16'd53602, 16'd28810, 16'd59989, 16'd22960, 16'd53839, 16'd42232, 16'd14194, 16'd24981, 16'd39628, 16'd25965, 16'd55041, 16'd3988, 16'd26055, 16'd4186, 16'd61693});
	test_expansion(128'h9ef75c62db355e1be9f756a91e90d9e1, {16'd59362, 16'd39300, 16'd26484, 16'd7100, 16'd15874, 16'd3726, 16'd22423, 16'd352, 16'd53507, 16'd29977, 16'd54407, 16'd27872, 16'd48947, 16'd7518, 16'd21380, 16'd55024, 16'd63969, 16'd60090, 16'd17694, 16'd19781, 16'd57301, 16'd58631, 16'd28512, 16'd6844, 16'd22913, 16'd45526});
	test_expansion(128'ha635c17e73aca0c0560ba1e2a487d0f3, {16'd56236, 16'd2092, 16'd58840, 16'd34746, 16'd40255, 16'd11912, 16'd40510, 16'd56536, 16'd15229, 16'd65535, 16'd32966, 16'd48238, 16'd38213, 16'd22855, 16'd23943, 16'd36277, 16'd12773, 16'd15608, 16'd3369, 16'd50197, 16'd54445, 16'd55462, 16'd31610, 16'd54538, 16'd17684, 16'd44665});
	test_expansion(128'hc788280f11f9fd6450d8dc8bfcdd1730, {16'd39359, 16'd40023, 16'd19658, 16'd32651, 16'd11936, 16'd11144, 16'd40990, 16'd17169, 16'd57082, 16'd54286, 16'd38775, 16'd55342, 16'd36687, 16'd61485, 16'd2872, 16'd25594, 16'd27269, 16'd5130, 16'd33828, 16'd15042, 16'd560, 16'd57723, 16'd51298, 16'd51560, 16'd7972, 16'd65334});
	test_expansion(128'h18df0c43e693ba6c67231b964be16821, {16'd14049, 16'd13765, 16'd693, 16'd23587, 16'd59272, 16'd61522, 16'd5803, 16'd63968, 16'd38683, 16'd1957, 16'd15686, 16'd18346, 16'd50270, 16'd61470, 16'd27143, 16'd58242, 16'd16577, 16'd57825, 16'd65491, 16'd54479, 16'd47282, 16'd46615, 16'd32084, 16'd48563, 16'd24284, 16'd50540});
	test_expansion(128'h7a7121f346259f2447e1473b6f8b1b43, {16'd38000, 16'd23029, 16'd25262, 16'd36991, 16'd43618, 16'd47293, 16'd26500, 16'd48924, 16'd34749, 16'd44687, 16'd35975, 16'd46086, 16'd38102, 16'd11664, 16'd46852, 16'd45152, 16'd59052, 16'd33289, 16'd33715, 16'd36097, 16'd40735, 16'd17466, 16'd57369, 16'd54347, 16'd61049, 16'd19875});
	test_expansion(128'h28494254e68b4caed6e395e40093fc0d, {16'd3655, 16'd4107, 16'd61687, 16'd38953, 16'd36144, 16'd19242, 16'd46100, 16'd60943, 16'd49772, 16'd51784, 16'd51932, 16'd54745, 16'd4349, 16'd62518, 16'd33967, 16'd21316, 16'd34172, 16'd31818, 16'd390, 16'd34498, 16'd13650, 16'd20506, 16'd15100, 16'd38388, 16'd16531, 16'd5702});
	test_expansion(128'h883f15f9ed259bf091d5c7c6c50be4aa, {16'd51492, 16'd8607, 16'd19920, 16'd52943, 16'd27645, 16'd11751, 16'd55013, 16'd59726, 16'd54375, 16'd23869, 16'd41847, 16'd62524, 16'd26761, 16'd41140, 16'd64933, 16'd44913, 16'd50620, 16'd52192, 16'd22913, 16'd64994, 16'd12934, 16'd14880, 16'd62246, 16'd29938, 16'd19118, 16'd38948});
	test_expansion(128'hb136e5d40f6762b6280248a4aa065b9a, {16'd25836, 16'd8608, 16'd45107, 16'd719, 16'd38070, 16'd6653, 16'd63930, 16'd59203, 16'd17921, 16'd31243, 16'd9354, 16'd16188, 16'd7324, 16'd27467, 16'd45460, 16'd62482, 16'd44324, 16'd32716, 16'd50587, 16'd38524, 16'd55597, 16'd59958, 16'd2395, 16'd32966, 16'd32312, 16'd47056});
	test_expansion(128'h158e4314433b45f9ca587520975a6427, {16'd13870, 16'd30754, 16'd62587, 16'd1231, 16'd50466, 16'd58893, 16'd31918, 16'd54217, 16'd29894, 16'd37419, 16'd27616, 16'd62698, 16'd57130, 16'd1013, 16'd18566, 16'd16407, 16'd48472, 16'd18682, 16'd58354, 16'd32389, 16'd59297, 16'd58981, 16'd48528, 16'd36480, 16'd31677, 16'd40380});
	test_expansion(128'ha954c3d956b50272c771a0ba4e92de45, {16'd47148, 16'd62513, 16'd21224, 16'd729, 16'd38968, 16'd15877, 16'd42936, 16'd21034, 16'd44739, 16'd45482, 16'd8893, 16'd44071, 16'd7447, 16'd53045, 16'd27848, 16'd63927, 16'd52296, 16'd27146, 16'd55100, 16'd21679, 16'd9929, 16'd38409, 16'd55965, 16'd22798, 16'd24341, 16'd60756});
	test_expansion(128'h36cff9a2951d3538b51a945a295f78b1, {16'd57481, 16'd29794, 16'd24998, 16'd31669, 16'd31788, 16'd20120, 16'd818, 16'd64516, 16'd1712, 16'd33439, 16'd56298, 16'd59212, 16'd28016, 16'd17263, 16'd21411, 16'd32892, 16'd24516, 16'd12800, 16'd33296, 16'd2466, 16'd30296, 16'd46789, 16'd7799, 16'd5424, 16'd4115, 16'd8603});
	test_expansion(128'h78b4f3b4f5ca189c28301f12e68bb7e9, {16'd49611, 16'd19184, 16'd1017, 16'd27392, 16'd28636, 16'd55781, 16'd2866, 16'd20086, 16'd11581, 16'd49529, 16'd486, 16'd33179, 16'd52954, 16'd61330, 16'd5761, 16'd40173, 16'd22028, 16'd17501, 16'd24662, 16'd65198, 16'd56828, 16'd56870, 16'd38978, 16'd10671, 16'd16594, 16'd28255});
	test_expansion(128'he370a6bb98f1093187dadd500815e578, {16'd2939, 16'd41506, 16'd64003, 16'd44848, 16'd12900, 16'd21188, 16'd3024, 16'd61070, 16'd46372, 16'd8570, 16'd55367, 16'd7013, 16'd26806, 16'd21552, 16'd62046, 16'd40993, 16'd29023, 16'd13349, 16'd53989, 16'd46956, 16'd21668, 16'd57627, 16'd49894, 16'd38975, 16'd13285, 16'd42387});
	test_expansion(128'h17acadd7072e27444db080844a32bb6c, {16'd58542, 16'd21989, 16'd40647, 16'd32871, 16'd51314, 16'd58833, 16'd38284, 16'd35362, 16'd48317, 16'd39390, 16'd7195, 16'd55975, 16'd6448, 16'd11053, 16'd49510, 16'd1939, 16'd51588, 16'd34387, 16'd24622, 16'd33238, 16'd40845, 16'd55810, 16'd59501, 16'd52548, 16'd47509, 16'd40237});
	test_expansion(128'h82807daaa1a040f74fa23b39f75cbd1d, {16'd19306, 16'd60043, 16'd6309, 16'd55267, 16'd55600, 16'd58614, 16'd31668, 16'd8444, 16'd38291, 16'd17662, 16'd5023, 16'd29739, 16'd4062, 16'd25728, 16'd58065, 16'd23148, 16'd22091, 16'd1502, 16'd43936, 16'd36851, 16'd26086, 16'd49574, 16'd52172, 16'd36023, 16'd24221, 16'd19360});
	test_expansion(128'hc0d34e7e1b2738a82d5f1a9b989fac10, {16'd48318, 16'd53253, 16'd40286, 16'd36985, 16'd43698, 16'd41770, 16'd13745, 16'd33816, 16'd16722, 16'd45066, 16'd52059, 16'd29074, 16'd47842, 16'd18596, 16'd29184, 16'd22125, 16'd34243, 16'd23344, 16'd21737, 16'd4900, 16'd60051, 16'd24270, 16'd318, 16'd56553, 16'd2307, 16'd7229});
	test_expansion(128'hb4b14912d1d8765ccb1aeebed1197c58, {16'd56205, 16'd61482, 16'd24105, 16'd59672, 16'd45347, 16'd26878, 16'd50623, 16'd56088, 16'd13903, 16'd59225, 16'd48545, 16'd36160, 16'd8708, 16'd30947, 16'd59612, 16'd56806, 16'd9675, 16'd50861, 16'd33156, 16'd29340, 16'd19059, 16'd37878, 16'd60153, 16'd53025, 16'd36541, 16'd28906});
	test_expansion(128'h640c90f32964326439baeb4159a29081, {16'd31437, 16'd12657, 16'd61800, 16'd44483, 16'd7430, 16'd34865, 16'd35203, 16'd25530, 16'd34981, 16'd27730, 16'd40562, 16'd63899, 16'd27040, 16'd55403, 16'd10926, 16'd22452, 16'd10991, 16'd54146, 16'd41191, 16'd64406, 16'd26815, 16'd58735, 16'd3476, 16'd49419, 16'd8438, 16'd3531});
	test_expansion(128'h4f8afbb5d9eb4c9f2b64b55e717b1e2f, {16'd47282, 16'd58945, 16'd36505, 16'd13847, 16'd34348, 16'd25190, 16'd41325, 16'd65509, 16'd38957, 16'd39590, 16'd21444, 16'd63721, 16'd25817, 16'd56974, 16'd4989, 16'd10437, 16'd18046, 16'd56546, 16'd59956, 16'd35362, 16'd54778, 16'd61109, 16'd4898, 16'd29920, 16'd54704, 16'd11137});
	test_expansion(128'h7fe0fea96590f6c6897ed88e5243fd0d, {16'd21487, 16'd60485, 16'd33016, 16'd35701, 16'd18491, 16'd855, 16'd60907, 16'd1789, 16'd59449, 16'd52781, 16'd25754, 16'd62161, 16'd26166, 16'd42416, 16'd27646, 16'd27514, 16'd2048, 16'd32846, 16'd47746, 16'd20497, 16'd52816, 16'd22165, 16'd58415, 16'd42701, 16'd43807, 16'd5715});
	test_expansion(128'h9280eec1e4851c19bef46ea8eab15336, {16'd9036, 16'd61643, 16'd63319, 16'd6814, 16'd63336, 16'd32418, 16'd5758, 16'd27173, 16'd8495, 16'd22326, 16'd36873, 16'd18506, 16'd57783, 16'd18467, 16'd44186, 16'd61897, 16'd22965, 16'd29273, 16'd52265, 16'd22493, 16'd43555, 16'd6008, 16'd39592, 16'd11929, 16'd18914, 16'd39010});
	test_expansion(128'he5b15870a3bce80fe37c07454797e8ca, {16'd2499, 16'd40904, 16'd45950, 16'd14112, 16'd16118, 16'd35678, 16'd41130, 16'd6545, 16'd16846, 16'd402, 16'd29797, 16'd31841, 16'd1978, 16'd55059, 16'd21100, 16'd61743, 16'd43987, 16'd2614, 16'd9761, 16'd32180, 16'd52172, 16'd30936, 16'd62340, 16'd45512, 16'd580, 16'd43232});
	test_expansion(128'h7de978635504f9952eff51c894ca8581, {16'd12666, 16'd3947, 16'd21499, 16'd62603, 16'd30432, 16'd31570, 16'd57686, 16'd17560, 16'd27024, 16'd59671, 16'd19592, 16'd5716, 16'd9845, 16'd34545, 16'd28095, 16'd59720, 16'd63683, 16'd5587, 16'd38053, 16'd34631, 16'd22009, 16'd24965, 16'd12580, 16'd39549, 16'd40536, 16'd14447});
	test_expansion(128'hd4dfafa04b7a36ee18ea1a2a892dfa82, {16'd17099, 16'd21001, 16'd45047, 16'd49009, 16'd58929, 16'd20331, 16'd59268, 16'd7134, 16'd46613, 16'd61533, 16'd3930, 16'd60548, 16'd47940, 16'd44942, 16'd26883, 16'd61578, 16'd6755, 16'd65390, 16'd28792, 16'd49184, 16'd35853, 16'd29993, 16'd14476, 16'd23889, 16'd39786, 16'd19527});
	test_expansion(128'h4b487c2915f7bd1f7c03f6883938e605, {16'd1263, 16'd4955, 16'd26014, 16'd50019, 16'd45038, 16'd25058, 16'd3176, 16'd56855, 16'd24712, 16'd46442, 16'd50256, 16'd35596, 16'd4621, 16'd35637, 16'd52962, 16'd37188, 16'd2820, 16'd29728, 16'd18853, 16'd4351, 16'd31078, 16'd19321, 16'd12300, 16'd49473, 16'd61943, 16'd23540});
	test_expansion(128'h7c81df73b73b28882396b3475215bb97, {16'd27952, 16'd46711, 16'd30338, 16'd15680, 16'd51936, 16'd4705, 16'd55767, 16'd20739, 16'd42342, 16'd4439, 16'd50956, 16'd30872, 16'd28183, 16'd39976, 16'd51001, 16'd8605, 16'd62055, 16'd47307, 16'd64486, 16'd36642, 16'd3903, 16'd44181, 16'd9666, 16'd58752, 16'd56707, 16'd35299});
	test_expansion(128'h273014b4dc7d0b7a6c5b61f523e8fe1e, {16'd45095, 16'd35363, 16'd14831, 16'd12090, 16'd43354, 16'd52735, 16'd2937, 16'd13564, 16'd47930, 16'd15048, 16'd12532, 16'd63935, 16'd1622, 16'd48046, 16'd46220, 16'd1195, 16'd42596, 16'd5562, 16'd60301, 16'd58798, 16'd41163, 16'd44141, 16'd23269, 16'd14655, 16'd17585, 16'd37316});
	test_expansion(128'h81ac93e115feb130cf1a28303c466104, {16'd61922, 16'd1123, 16'd36982, 16'd55276, 16'd24772, 16'd7123, 16'd47423, 16'd2879, 16'd21809, 16'd22599, 16'd48855, 16'd39240, 16'd541, 16'd53337, 16'd26118, 16'd13299, 16'd56058, 16'd59276, 16'd31245, 16'd54103, 16'd316, 16'd6638, 16'd44514, 16'd9443, 16'd10667, 16'd22252});
	test_expansion(128'h0606e49c43dcee1c8375d41b63c325bc, {16'd38620, 16'd32213, 16'd36600, 16'd320, 16'd1396, 16'd44548, 16'd38017, 16'd54100, 16'd33647, 16'd12914, 16'd4354, 16'd52002, 16'd45996, 16'd53203, 16'd27551, 16'd19515, 16'd47939, 16'd29416, 16'd22199, 16'd52294, 16'd38840, 16'd20127, 16'd59815, 16'd16678, 16'd32292, 16'd61301});
	test_expansion(128'h121babfb915a775c6a620587298bf567, {16'd61972, 16'd5922, 16'd11408, 16'd39394, 16'd64885, 16'd30231, 16'd21067, 16'd2473, 16'd15951, 16'd21049, 16'd50265, 16'd62611, 16'd58980, 16'd25434, 16'd49216, 16'd8111, 16'd915, 16'd64006, 16'd13233, 16'd38873, 16'd16668, 16'd45582, 16'd6123, 16'd43359, 16'd60491, 16'd41363});
	test_expansion(128'h88f9953335e96f949183d8c501e54c43, {16'd60224, 16'd19660, 16'd22604, 16'd32091, 16'd14786, 16'd46091, 16'd38124, 16'd6160, 16'd3197, 16'd52279, 16'd4533, 16'd29383, 16'd33626, 16'd24675, 16'd24548, 16'd62438, 16'd29125, 16'd636, 16'd2664, 16'd3346, 16'd8948, 16'd65311, 16'd29104, 16'd53332, 16'd65535, 16'd43698});
	test_expansion(128'h8dcc6ba6ae1dbb7412c7160921d8bfbf, {16'd14589, 16'd35740, 16'd33667, 16'd20292, 16'd9586, 16'd12935, 16'd63103, 16'd61019, 16'd37797, 16'd25312, 16'd53871, 16'd33538, 16'd50756, 16'd60959, 16'd63394, 16'd63956, 16'd18814, 16'd29361, 16'd5110, 16'd29359, 16'd48480, 16'd54887, 16'd32682, 16'd50017, 16'd42863, 16'd45644});
	test_expansion(128'he3ca354bae19a4e4c01df43d8fbca499, {16'd27074, 16'd62654, 16'd32658, 16'd14772, 16'd44613, 16'd32590, 16'd64723, 16'd22994, 16'd22046, 16'd27553, 16'd37439, 16'd21476, 16'd65385, 16'd26512, 16'd27593, 16'd27611, 16'd26286, 16'd44561, 16'd36569, 16'd26203, 16'd25146, 16'd22193, 16'd22895, 16'd51613, 16'd50206, 16'd61496});
	test_expansion(128'h209c723792b2899c102e4d64a313d5dc, {16'd35356, 16'd36273, 16'd31442, 16'd31404, 16'd12473, 16'd52383, 16'd47157, 16'd8690, 16'd8730, 16'd52895, 16'd34463, 16'd45265, 16'd42783, 16'd43462, 16'd36530, 16'd35585, 16'd28956, 16'd36943, 16'd35233, 16'd23804, 16'd45019, 16'd16090, 16'd65011, 16'd1731, 16'd19844, 16'd16142});
	test_expansion(128'hb9bd9dd931c460861f6eb79f45a5c6b8, {16'd16349, 16'd52696, 16'd44373, 16'd14455, 16'd29009, 16'd54064, 16'd20123, 16'd1321, 16'd37043, 16'd59939, 16'd58819, 16'd31654, 16'd8557, 16'd12576, 16'd34180, 16'd3867, 16'd37059, 16'd53116, 16'd60314, 16'd24460, 16'd18397, 16'd64260, 16'd39834, 16'd10579, 16'd15177, 16'd44095});
	test_expansion(128'h27cfd3a6b82db4213f3d0934378e1400, {16'd29656, 16'd37459, 16'd56163, 16'd1178, 16'd13140, 16'd13840, 16'd60495, 16'd32463, 16'd62697, 16'd28232, 16'd60030, 16'd47646, 16'd9533, 16'd36582, 16'd22910, 16'd7277, 16'd18974, 16'd723, 16'd28541, 16'd36335, 16'd14645, 16'd62541, 16'd37657, 16'd65445, 16'd55498, 16'd29107});
	test_expansion(128'h804a63a0640f1bca95463d2b14770f1d, {16'd1395, 16'd41824, 16'd59592, 16'd13871, 16'd31380, 16'd8733, 16'd59361, 16'd28712, 16'd2941, 16'd1135, 16'd42697, 16'd59850, 16'd29229, 16'd54742, 16'd62611, 16'd61390, 16'd45495, 16'd4762, 16'd21387, 16'd12895, 16'd56116, 16'd15329, 16'd1300, 16'd63260, 16'd56141, 16'd13917});
	test_expansion(128'hfe33ed637376ed1707a459855b577500, {16'd29561, 16'd56871, 16'd30416, 16'd46458, 16'd568, 16'd1096, 16'd27977, 16'd46265, 16'd45397, 16'd44212, 16'd21274, 16'd47300, 16'd61030, 16'd46791, 16'd6415, 16'd34568, 16'd20260, 16'd41652, 16'd51055, 16'd31257, 16'd54705, 16'd45619, 16'd14013, 16'd24688, 16'd2705, 16'd57975});
	test_expansion(128'h9049875c9bf86df495364efb93dd6185, {16'd41881, 16'd56432, 16'd32384, 16'd51016, 16'd41216, 16'd31777, 16'd1715, 16'd10664, 16'd26170, 16'd27874, 16'd47128, 16'd40165, 16'd47848, 16'd58223, 16'd41003, 16'd47961, 16'd62651, 16'd64752, 16'd52667, 16'd52170, 16'd17250, 16'd3467, 16'd22058, 16'd63462, 16'd24737, 16'd64101});
	test_expansion(128'h1ebc5a94ed962d6e275c87e56bc33166, {16'd58158, 16'd4481, 16'd6081, 16'd19691, 16'd63776, 16'd47915, 16'd4125, 16'd49185, 16'd64238, 16'd23139, 16'd45409, 16'd17279, 16'd26828, 16'd7066, 16'd43343, 16'd53922, 16'd12782, 16'd6917, 16'd4826, 16'd40, 16'd47814, 16'd53308, 16'd33219, 16'd21542, 16'd38767, 16'd9517});
	test_expansion(128'h0fd242e79cf65350f01ce4182cb59967, {16'd41669, 16'd56873, 16'd64825, 16'd12887, 16'd7795, 16'd16485, 16'd39346, 16'd51482, 16'd60814, 16'd51893, 16'd55752, 16'd12273, 16'd23293, 16'd14855, 16'd24085, 16'd23096, 16'd21344, 16'd4337, 16'd37522, 16'd3541, 16'd18876, 16'd17768, 16'd41243, 16'd44056, 16'd11952, 16'd2795});
	test_expansion(128'h44d157747bd8f9297d87808df54a0dba, {16'd21210, 16'd52997, 16'd14552, 16'd24207, 16'd47489, 16'd47459, 16'd42479, 16'd30101, 16'd24054, 16'd44519, 16'd46797, 16'd46923, 16'd16343, 16'd38444, 16'd51330, 16'd33558, 16'd26740, 16'd4446, 16'd30073, 16'd44519, 16'd64194, 16'd29219, 16'd46705, 16'd29004, 16'd20794, 16'd37447});
	test_expansion(128'h9f51ae657edb2be46e496b3460485150, {16'd31695, 16'd36287, 16'd7824, 16'd44163, 16'd59820, 16'd21883, 16'd20656, 16'd47042, 16'd60843, 16'd2804, 16'd49800, 16'd9856, 16'd44603, 16'd48241, 16'd50565, 16'd8155, 16'd23880, 16'd50775, 16'd37269, 16'd47450, 16'd53923, 16'd26748, 16'd16520, 16'd17219, 16'd58313, 16'd25607});
	test_expansion(128'h0ccb9db2edf34b3f90fdd1c3cb9b96df, {16'd55444, 16'd19693, 16'd40170, 16'd46467, 16'd38452, 16'd31330, 16'd52649, 16'd61213, 16'd24643, 16'd62173, 16'd1297, 16'd25372, 16'd733, 16'd54959, 16'd21308, 16'd25655, 16'd56865, 16'd25514, 16'd64504, 16'd14880, 16'd20986, 16'd28176, 16'd37703, 16'd56445, 16'd45295, 16'd24015});
	test_expansion(128'h0c893faa96424f5d72d4081b853eb4c3, {16'd21828, 16'd63324, 16'd23233, 16'd21314, 16'd19731, 16'd38208, 16'd41656, 16'd63698, 16'd38717, 16'd49191, 16'd20834, 16'd56629, 16'd2603, 16'd5604, 16'd24736, 16'd29120, 16'd11044, 16'd22519, 16'd4952, 16'd26846, 16'd45712, 16'd34031, 16'd47110, 16'd29978, 16'd5894, 16'd22063});
	test_expansion(128'hb6e0f73b2499b9d32254213b8fa2b369, {16'd29747, 16'd1272, 16'd56693, 16'd62008, 16'd31958, 16'd39025, 16'd62595, 16'd4363, 16'd45164, 16'd34581, 16'd13601, 16'd20888, 16'd19827, 16'd4555, 16'd11951, 16'd20356, 16'd19193, 16'd52416, 16'd57571, 16'd14264, 16'd48211, 16'd28753, 16'd29524, 16'd33461, 16'd10564, 16'd34385});
	test_expansion(128'h7f771df4570e49ef817a5b3fa6923e51, {16'd46351, 16'd24739, 16'd48716, 16'd49715, 16'd19183, 16'd35004, 16'd21832, 16'd56578, 16'd58712, 16'd25716, 16'd58254, 16'd667, 16'd9408, 16'd20043, 16'd1378, 16'd61032, 16'd63951, 16'd15063, 16'd60767, 16'd61161, 16'd58539, 16'd6302, 16'd29229, 16'd5764, 16'd357, 16'd18366});
	test_expansion(128'h227a1c28bb75063129208bd26674a59b, {16'd30804, 16'd3630, 16'd17297, 16'd23599, 16'd33130, 16'd39931, 16'd22603, 16'd40750, 16'd52167, 16'd9870, 16'd45849, 16'd10489, 16'd54418, 16'd23239, 16'd19963, 16'd7014, 16'd14520, 16'd39236, 16'd39548, 16'd54371, 16'd6601, 16'd8935, 16'd27255, 16'd33009, 16'd59007, 16'd4336});
	test_expansion(128'h6435bb44cb9b15c87331e5b2e8d8d322, {16'd3899, 16'd44074, 16'd51886, 16'd35255, 16'd26062, 16'd34042, 16'd59650, 16'd46354, 16'd43567, 16'd55038, 16'd62125, 16'd8356, 16'd63665, 16'd33800, 16'd4474, 16'd64610, 16'd4626, 16'd19635, 16'd65204, 16'd55182, 16'd26520, 16'd59636, 16'd26206, 16'd56817, 16'd47034, 16'd3602});
	test_expansion(128'h35b644661e924c3bbcf7f0e09f062fe4, {16'd21891, 16'd3323, 16'd13909, 16'd62906, 16'd6391, 16'd35283, 16'd41001, 16'd38371, 16'd34815, 16'd65128, 16'd27562, 16'd35731, 16'd54065, 16'd50447, 16'd21095, 16'd37746, 16'd2133, 16'd45498, 16'd3302, 16'd16184, 16'd24141, 16'd9222, 16'd15807, 16'd63728, 16'd937, 16'd771});
	test_expansion(128'h05d60f0b2c80034954999951e2fc3e6b, {16'd62648, 16'd2291, 16'd11315, 16'd29497, 16'd14363, 16'd23897, 16'd60685, 16'd50933, 16'd29864, 16'd42070, 16'd40243, 16'd9219, 16'd53803, 16'd60444, 16'd44182, 16'd23827, 16'd291, 16'd28001, 16'd463, 16'd62784, 16'd43280, 16'd54066, 16'd59719, 16'd58454, 16'd13611, 16'd29582});
	test_expansion(128'h6c02f35b4b6bba630d0dbbbe171fc7e0, {16'd20650, 16'd219, 16'd49403, 16'd3198, 16'd10878, 16'd15280, 16'd2456, 16'd22549, 16'd20900, 16'd5620, 16'd4439, 16'd51463, 16'd24386, 16'd51605, 16'd38398, 16'd8202, 16'd8821, 16'd61674, 16'd21163, 16'd55284, 16'd22900, 16'd13266, 16'd3143, 16'd11522, 16'd30301, 16'd35578});
	test_expansion(128'h671e3029310b976ec8c3ed734c705450, {16'd40878, 16'd51823, 16'd41532, 16'd58316, 16'd47809, 16'd22276, 16'd21242, 16'd14434, 16'd53909, 16'd30657, 16'd48828, 16'd13273, 16'd30978, 16'd40646, 16'd27305, 16'd23767, 16'd42370, 16'd59027, 16'd26840, 16'd28727, 16'd1602, 16'd30947, 16'd20539, 16'd5959, 16'd30434, 16'd46052});
	test_expansion(128'hd0771b38581a0557a2f01d7333fbfa20, {16'd51828, 16'd32357, 16'd42957, 16'd37765, 16'd18635, 16'd35132, 16'd25082, 16'd57485, 16'd213, 16'd13897, 16'd45559, 16'd4767, 16'd38575, 16'd57631, 16'd30925, 16'd7359, 16'd61776, 16'd48363, 16'd43445, 16'd13081, 16'd43956, 16'd53201, 16'd57317, 16'd43993, 16'd17360, 16'd30648});
	test_expansion(128'h2938b790923bf7b4f09c51ce557c59d9, {16'd25277, 16'd19115, 16'd34422, 16'd11666, 16'd22455, 16'd63276, 16'd12209, 16'd61586, 16'd41471, 16'd25183, 16'd2114, 16'd54569, 16'd3112, 16'd19614, 16'd58359, 16'd5775, 16'd48087, 16'd51095, 16'd45813, 16'd31365, 16'd9505, 16'd47548, 16'd56133, 16'd32703, 16'd57315, 16'd17004});
	test_expansion(128'h5fb3eee933903356648706b74928a65a, {16'd49516, 16'd39427, 16'd15240, 16'd25013, 16'd10371, 16'd49683, 16'd26225, 16'd60168, 16'd59205, 16'd43315, 16'd56187, 16'd42377, 16'd45845, 16'd56795, 16'd59478, 16'd6620, 16'd6077, 16'd35528, 16'd38192, 16'd45123, 16'd30582, 16'd22505, 16'd33294, 16'd7093, 16'd48897, 16'd61711});
	test_expansion(128'h1c4b7a7845176e3264ffe6b13c13928e, {16'd13127, 16'd5981, 16'd41265, 16'd57532, 16'd49795, 16'd35505, 16'd30680, 16'd11556, 16'd11063, 16'd54141, 16'd25208, 16'd52710, 16'd62361, 16'd6980, 16'd41665, 16'd59139, 16'd41194, 16'd36034, 16'd13511, 16'd65364, 16'd8367, 16'd14031, 16'd6282, 16'd6766, 16'd60204, 16'd47411});
	test_expansion(128'h2619cb90f002ffabdd749ec1363f358d, {16'd59252, 16'd8387, 16'd11719, 16'd19836, 16'd55733, 16'd11561, 16'd1116, 16'd44193, 16'd60852, 16'd28029, 16'd64966, 16'd63043, 16'd9080, 16'd63965, 16'd42716, 16'd58664, 16'd37001, 16'd50408, 16'd35446, 16'd1107, 16'd29758, 16'd27987, 16'd5474, 16'd42509, 16'd14878, 16'd12980});
	test_expansion(128'h7279a646e2870e3b4f728ad0c860e8a0, {16'd57876, 16'd45627, 16'd57898, 16'd33073, 16'd32358, 16'd49211, 16'd6397, 16'd30427, 16'd38490, 16'd57168, 16'd54459, 16'd9385, 16'd62455, 16'd20158, 16'd41565, 16'd21488, 16'd30565, 16'd39708, 16'd55660, 16'd14936, 16'd25893, 16'd34266, 16'd28624, 16'd48569, 16'd21829, 16'd32278});
	test_expansion(128'ha42ee324e61ce5c835dcac1363a89c83, {16'd39575, 16'd39639, 16'd37031, 16'd19225, 16'd24323, 16'd60543, 16'd17728, 16'd61544, 16'd44751, 16'd30526, 16'd20511, 16'd7430, 16'd26760, 16'd13903, 16'd65439, 16'd55621, 16'd29963, 16'd51013, 16'd65385, 16'd15460, 16'd8583, 16'd18505, 16'd38267, 16'd15877, 16'd43898, 16'd46828});
	test_expansion(128'h25e047e14cbb57fa914a99659edf1aa7, {16'd46124, 16'd32508, 16'd48916, 16'd58880, 16'd3833, 16'd44906, 16'd26462, 16'd47196, 16'd23936, 16'd1054, 16'd35081, 16'd5890, 16'd2188, 16'd14764, 16'd40843, 16'd13288, 16'd1726, 16'd18378, 16'd54018, 16'd44390, 16'd17716, 16'd44258, 16'd19600, 16'd56114, 16'd24405, 16'd59519});
	test_expansion(128'h8088084bb337fc39b39f88a7d2c56ca9, {16'd15941, 16'd46807, 16'd60375, 16'd37916, 16'd41791, 16'd15706, 16'd62598, 16'd60323, 16'd54252, 16'd38880, 16'd56940, 16'd45664, 16'd54143, 16'd17295, 16'd41898, 16'd30596, 16'd19897, 16'd51529, 16'd50793, 16'd15876, 16'd20220, 16'd19258, 16'd14508, 16'd47597, 16'd37579, 16'd27146});
	test_expansion(128'hff1e4f64fbf1f82b87f6a0abe12bf021, {16'd35033, 16'd56730, 16'd63536, 16'd46407, 16'd36342, 16'd6368, 16'd27782, 16'd59335, 16'd42697, 16'd25872, 16'd50105, 16'd45639, 16'd54203, 16'd61024, 16'd41007, 16'd64445, 16'd29426, 16'd44922, 16'd13681, 16'd43946, 16'd7902, 16'd48364, 16'd14465, 16'd52814, 16'd62103, 16'd41937});
	test_expansion(128'h5ae3079d7431b3a4483fa3b3981f5755, {16'd16726, 16'd59185, 16'd63832, 16'd63810, 16'd17102, 16'd27121, 16'd58131, 16'd40330, 16'd51346, 16'd33865, 16'd29143, 16'd35073, 16'd22374, 16'd59242, 16'd6638, 16'd42200, 16'd33306, 16'd15090, 16'd31508, 16'd7472, 16'd15, 16'd16484, 16'd2560, 16'd48009, 16'd47339, 16'd56249});
	test_expansion(128'hf38220932ccf523f516dafdb70eaa76e, {16'd3377, 16'd14446, 16'd1011, 16'd55636, 16'd34860, 16'd1749, 16'd3782, 16'd60576, 16'd52075, 16'd9343, 16'd47559, 16'd28786, 16'd50206, 16'd60005, 16'd48796, 16'd13124, 16'd35367, 16'd49807, 16'd17667, 16'd60947, 16'd29068, 16'd14260, 16'd58489, 16'd9328, 16'd46007, 16'd24927});
	test_expansion(128'h31794c993d14cdc963660409a6a6a1ad, {16'd50174, 16'd65119, 16'd32076, 16'd1835, 16'd53856, 16'd48812, 16'd61575, 16'd59392, 16'd63073, 16'd47600, 16'd45580, 16'd15819, 16'd19781, 16'd26467, 16'd41301, 16'd1522, 16'd39490, 16'd48036, 16'd28106, 16'd54461, 16'd17715, 16'd15282, 16'd53595, 16'd63615, 16'd4669, 16'd52347});
	test_expansion(128'h9cc453cd19f60d4704ea12b477c13726, {16'd32773, 16'd25931, 16'd36565, 16'd16611, 16'd4857, 16'd21371, 16'd37480, 16'd34141, 16'd59213, 16'd10878, 16'd40318, 16'd37253, 16'd428, 16'd46934, 16'd19405, 16'd47795, 16'd33994, 16'd39945, 16'd9994, 16'd5211, 16'd55474, 16'd11257, 16'd7136, 16'd6024, 16'd56597, 16'd2840});
	test_expansion(128'hb43cd7a433f5f010beb24baf3902c428, {16'd48857, 16'd25127, 16'd26058, 16'd37856, 16'd45027, 16'd34022, 16'd10945, 16'd8336, 16'd34049, 16'd60242, 16'd27405, 16'd27626, 16'd5689, 16'd11728, 16'd61933, 16'd17824, 16'd960, 16'd18420, 16'd17284, 16'd20568, 16'd49459, 16'd55341, 16'd45757, 16'd30008, 16'd438, 16'd44925});
	test_expansion(128'h1543f11e290301ba296fd10d249709a2, {16'd25639, 16'd53370, 16'd34315, 16'd15625, 16'd3196, 16'd49646, 16'd20976, 16'd4369, 16'd4032, 16'd41597, 16'd26914, 16'd38744, 16'd43611, 16'd3723, 16'd62968, 16'd8198, 16'd36900, 16'd55775, 16'd29274, 16'd11939, 16'd18562, 16'd54824, 16'd55109, 16'd38591, 16'd61760, 16'd11464});
	test_expansion(128'he7be2be05c9ad57fb18ac052a6404aa5, {16'd1639, 16'd27873, 16'd25118, 16'd43527, 16'd797, 16'd56121, 16'd65179, 16'd5724, 16'd33376, 16'd10474, 16'd64731, 16'd24555, 16'd37082, 16'd58708, 16'd12207, 16'd44573, 16'd34549, 16'd51351, 16'd53228, 16'd4286, 16'd51386, 16'd37910, 16'd56699, 16'd20607, 16'd54118, 16'd24159});
	test_expansion(128'hcb808422f293035ebe2e1802100c6ad7, {16'd57001, 16'd53753, 16'd25131, 16'd7844, 16'd45245, 16'd19459, 16'd42362, 16'd42070, 16'd38569, 16'd53168, 16'd34595, 16'd16327, 16'd37752, 16'd7062, 16'd48241, 16'd25034, 16'd102, 16'd34134, 16'd59568, 16'd6008, 16'd50146, 16'd3513, 16'd61920, 16'd55855, 16'd40572, 16'd43004});
	test_expansion(128'h0eb777354944264f835d80bef26639aa, {16'd18405, 16'd36493, 16'd43792, 16'd5677, 16'd37219, 16'd10997, 16'd1454, 16'd10610, 16'd38771, 16'd28710, 16'd10949, 16'd63695, 16'd44078, 16'd21582, 16'd12706, 16'd56247, 16'd7361, 16'd64151, 16'd54956, 16'd26478, 16'd53833, 16'd30969, 16'd18205, 16'd15815, 16'd19831, 16'd20536});
	test_expansion(128'h0bbde6c58f9acec2b43cdbf29bed9f92, {16'd64742, 16'd27587, 16'd16369, 16'd14347, 16'd6927, 16'd44704, 16'd14459, 16'd38300, 16'd12375, 16'd52985, 16'd52639, 16'd40605, 16'd6902, 16'd4550, 16'd20546, 16'd37487, 16'd5581, 16'd19543, 16'd46159, 16'd26631, 16'd46177, 16'd31282, 16'd1993, 16'd4856, 16'd2520, 16'd47537});
	test_expansion(128'hb64199b4761458d05c1318d8764d2b23, {16'd18712, 16'd51637, 16'd33520, 16'd50571, 16'd1589, 16'd23393, 16'd65418, 16'd29611, 16'd814, 16'd19313, 16'd43568, 16'd27340, 16'd19361, 16'd35826, 16'd40179, 16'd51656, 16'd35643, 16'd15946, 16'd33590, 16'd63260, 16'd30148, 16'd54751, 16'd22114, 16'd11679, 16'd35333, 16'd9959});
	test_expansion(128'h90e83c571060356d3916df5c676cbb00, {16'd30464, 16'd19340, 16'd30216, 16'd14079, 16'd65061, 16'd61554, 16'd7165, 16'd58371, 16'd51470, 16'd21191, 16'd45034, 16'd10170, 16'd22814, 16'd1568, 16'd47079, 16'd57149, 16'd54329, 16'd55220, 16'd51351, 16'd51771, 16'd50758, 16'd55197, 16'd57960, 16'd18226, 16'd60999, 16'd1306});
	test_expansion(128'hb8ab9ecc0a69da35c850b8deeda99c76, {16'd53637, 16'd13405, 16'd16553, 16'd22209, 16'd6536, 16'd20048, 16'd28031, 16'd56173, 16'd51785, 16'd34756, 16'd28421, 16'd39157, 16'd40102, 16'd60604, 16'd41943, 16'd7706, 16'd20181, 16'd18364, 16'd10725, 16'd54989, 16'd39047, 16'd17596, 16'd42892, 16'd38069, 16'd20369, 16'd8775});
	test_expansion(128'h327df9a3a827c539ecf970bdc7652b16, {16'd41935, 16'd28005, 16'd38999, 16'd33156, 16'd53389, 16'd21711, 16'd16887, 16'd48523, 16'd41100, 16'd57782, 16'd59933, 16'd20567, 16'd19643, 16'd2352, 16'd33428, 16'd60066, 16'd10832, 16'd25222, 16'd63486, 16'd9266, 16'd16891, 16'd11785, 16'd25214, 16'd23266, 16'd23970, 16'd50715});
	test_expansion(128'h5639f113aeafb1e1129356f60eb75dcc, {16'd12476, 16'd48917, 16'd46802, 16'd13956, 16'd14640, 16'd28527, 16'd24486, 16'd15797, 16'd6839, 16'd62810, 16'd43799, 16'd12114, 16'd9406, 16'd63170, 16'd13254, 16'd10762, 16'd61812, 16'd28338, 16'd30816, 16'd47893, 16'd53466, 16'd65293, 16'd56918, 16'd62695, 16'd20828, 16'd25440});
	test_expansion(128'h061f69741628ee693e9845a32a865d0b, {16'd28236, 16'd56634, 16'd13383, 16'd34845, 16'd34420, 16'd25444, 16'd57054, 16'd9798, 16'd14140, 16'd50995, 16'd48440, 16'd33624, 16'd52934, 16'd57378, 16'd24585, 16'd35269, 16'd55946, 16'd19753, 16'd32541, 16'd17489, 16'd12970, 16'd23457, 16'd22907, 16'd10917, 16'd9091, 16'd12482});
	test_expansion(128'hdcdccbf89132a1cb8533b77bdab40ee3, {16'd32394, 16'd27850, 16'd33938, 16'd13622, 16'd47259, 16'd38640, 16'd26191, 16'd14251, 16'd54034, 16'd51788, 16'd33686, 16'd51609, 16'd22033, 16'd22568, 16'd17346, 16'd23, 16'd46799, 16'd46359, 16'd10680, 16'd53879, 16'd27211, 16'd26199, 16'd47404, 16'd42694, 16'd32064, 16'd7539});
	test_expansion(128'hc45fe7c033e60eafa26205375a3cc0d5, {16'd30117, 16'd58905, 16'd7235, 16'd50977, 16'd12962, 16'd55489, 16'd31629, 16'd11821, 16'd50164, 16'd17007, 16'd4779, 16'd790, 16'd32952, 16'd12873, 16'd43232, 16'd58439, 16'd1989, 16'd63636, 16'd50646, 16'd56212, 16'd1417, 16'd56872, 16'd51826, 16'd12283, 16'd10183, 16'd20461});
	test_expansion(128'h80746ddc12c742a3ae8bb1036272c144, {16'd60935, 16'd47740, 16'd21682, 16'd40270, 16'd29395, 16'd41775, 16'd16151, 16'd35966, 16'd38029, 16'd20328, 16'd51811, 16'd39239, 16'd3948, 16'd37727, 16'd38112, 16'd29578, 16'd43866, 16'd33970, 16'd49251, 16'd2596, 16'd24616, 16'd40853, 16'd1351, 16'd47547, 16'd2954, 16'd36073});
	test_expansion(128'hbe59b3bbfb353e3a0b918200f6f5b8a2, {16'd29051, 16'd21960, 16'd15635, 16'd31771, 16'd16872, 16'd5586, 16'd56700, 16'd50007, 16'd27862, 16'd5879, 16'd47933, 16'd64780, 16'd57710, 16'd23999, 16'd14869, 16'd49125, 16'd36464, 16'd30067, 16'd52257, 16'd55151, 16'd21880, 16'd6463, 16'd48755, 16'd18097, 16'd23128, 16'd33678});
	test_expansion(128'h61464096e466f73de91cb8290ea14c3f, {16'd33515, 16'd25464, 16'd64016, 16'd7327, 16'd54830, 16'd62969, 16'd129, 16'd4000, 16'd50984, 16'd21003, 16'd14314, 16'd25327, 16'd27178, 16'd10613, 16'd64726, 16'd31473, 16'd34735, 16'd25076, 16'd63957, 16'd14848, 16'd15499, 16'd16130, 16'd32097, 16'd59397, 16'd2372, 16'd25517});
	test_expansion(128'he462d6d1dba629eb651142b3dd0d241a, {16'd37620, 16'd2933, 16'd31347, 16'd643, 16'd42111, 16'd56561, 16'd5050, 16'd36043, 16'd35098, 16'd903, 16'd29632, 16'd33592, 16'd38165, 16'd61938, 16'd22739, 16'd40745, 16'd54971, 16'd56634, 16'd22058, 16'd35295, 16'd34199, 16'd40042, 16'd4204, 16'd56734, 16'd4886, 16'd35144});
	test_expansion(128'h3e7909057f020b0f88cc215b5118212a, {16'd5280, 16'd8146, 16'd51794, 16'd21227, 16'd15535, 16'd46716, 16'd21491, 16'd28170, 16'd14007, 16'd20337, 16'd9952, 16'd7549, 16'd48832, 16'd46957, 16'd54640, 16'd47021, 16'd37036, 16'd5042, 16'd1822, 16'd62858, 16'd44049, 16'd25222, 16'd40410, 16'd12330, 16'd50909, 16'd2742});
	test_expansion(128'h59877db41a3892fb31a58e5991286d47, {16'd8148, 16'd41233, 16'd45135, 16'd37329, 16'd38445, 16'd13768, 16'd11454, 16'd3258, 16'd64245, 16'd13801, 16'd60367, 16'd26448, 16'd31517, 16'd5280, 16'd16583, 16'd23781, 16'd28846, 16'd50121, 16'd7002, 16'd33538, 16'd53882, 16'd23406, 16'd32655, 16'd31153, 16'd16465, 16'd52270});
	test_expansion(128'h50ed8a3b09d1fae81c5d9fef8d5c417c, {16'd9433, 16'd41474, 16'd23558, 16'd3261, 16'd51913, 16'd12951, 16'd9057, 16'd39282, 16'd9613, 16'd29011, 16'd48582, 16'd21268, 16'd2396, 16'd29341, 16'd19301, 16'd17685, 16'd31549, 16'd21136, 16'd65388, 16'd45430, 16'd3059, 16'd19959, 16'd7242, 16'd15005, 16'd20715, 16'd61831});
	test_expansion(128'hac6e668302a1e0eb0a38e2eea7f848c7, {16'd26875, 16'd53916, 16'd34808, 16'd42523, 16'd18046, 16'd47452, 16'd2428, 16'd51434, 16'd5476, 16'd33316, 16'd576, 16'd61952, 16'd18206, 16'd52577, 16'd62247, 16'd13761, 16'd17841, 16'd15331, 16'd27324, 16'd61925, 16'd31833, 16'd12383, 16'd4179, 16'd40846, 16'd14112, 16'd41295});
	test_expansion(128'hd7fa8c3a5bed4e2c7ac7390c75a5cc14, {16'd45765, 16'd2890, 16'd3625, 16'd64614, 16'd19802, 16'd49795, 16'd41211, 16'd10841, 16'd19289, 16'd28739, 16'd26553, 16'd20301, 16'd36690, 16'd10656, 16'd43331, 16'd48382, 16'd60898, 16'd7224, 16'd23004, 16'd3125, 16'd3744, 16'd23800, 16'd30740, 16'd44343, 16'd53472, 16'd43416});
	test_expansion(128'hfc000a6c7d22e6847878a410d21165bd, {16'd57079, 16'd2748, 16'd54426, 16'd49488, 16'd53342, 16'd34792, 16'd28853, 16'd64505, 16'd30227, 16'd3379, 16'd32352, 16'd7495, 16'd61976, 16'd8119, 16'd46249, 16'd21640, 16'd32467, 16'd44286, 16'd1317, 16'd13561, 16'd35558, 16'd55877, 16'd37870, 16'd43647, 16'd20254, 16'd3171});
	test_expansion(128'h2b4c97b11c7d7e9ba33add8b5b1a6bc3, {16'd18850, 16'd26702, 16'd58695, 16'd8255, 16'd29014, 16'd40713, 16'd32613, 16'd2472, 16'd53542, 16'd65521, 16'd55627, 16'd41018, 16'd9198, 16'd34662, 16'd63977, 16'd35034, 16'd8371, 16'd54183, 16'd35694, 16'd8122, 16'd35691, 16'd61140, 16'd49389, 16'd58450, 16'd61113, 16'd46782});
	test_expansion(128'he58df1360fd68d93b8937333d1f91c67, {16'd32691, 16'd29262, 16'd21133, 16'd1194, 16'd34330, 16'd18319, 16'd11634, 16'd22957, 16'd51797, 16'd17760, 16'd38210, 16'd54245, 16'd35340, 16'd44343, 16'd52006, 16'd25652, 16'd24064, 16'd53949, 16'd7015, 16'd41105, 16'd6993, 16'd51512, 16'd12369, 16'd2470, 16'd63340, 16'd59255});
	test_expansion(128'h0df069d9ec25aeee6ff09a320b2bebd8, {16'd41590, 16'd53541, 16'd22102, 16'd49894, 16'd27636, 16'd26008, 16'd14178, 16'd31424, 16'd37495, 16'd51779, 16'd53506, 16'd44967, 16'd25503, 16'd37210, 16'd33637, 16'd61990, 16'd57328, 16'd34272, 16'd6226, 16'd26964, 16'd19180, 16'd12906, 16'd46465, 16'd21040, 16'd50674, 16'd63512});
	test_expansion(128'h523a9b9a33141c8b1333b5b9cf81dc94, {16'd46175, 16'd2038, 16'd10500, 16'd5133, 16'd50608, 16'd24345, 16'd31053, 16'd12065, 16'd58664, 16'd59724, 16'd2185, 16'd33208, 16'd63130, 16'd32595, 16'd36043, 16'd4348, 16'd49930, 16'd59617, 16'd2161, 16'd36544, 16'd2116, 16'd57212, 16'd59874, 16'd1744, 16'd46938, 16'd49835});
	test_expansion(128'h8ea26ba53c1b2450970a0136fe135387, {16'd12896, 16'd63819, 16'd59130, 16'd61487, 16'd39241, 16'd2477, 16'd16015, 16'd61858, 16'd10798, 16'd49848, 16'd21294, 16'd12675, 16'd29641, 16'd17643, 16'd48068, 16'd25879, 16'd39845, 16'd46680, 16'd19999, 16'd56806, 16'd57017, 16'd12403, 16'd17624, 16'd37561, 16'd12112, 16'd17932});
	test_expansion(128'he7ab89cea25bf6cd5ef63b2e5d80b380, {16'd25259, 16'd32135, 16'd61536, 16'd11266, 16'd1425, 16'd7744, 16'd49213, 16'd6610, 16'd56322, 16'd34700, 16'd47811, 16'd22938, 16'd19325, 16'd15606, 16'd12701, 16'd51814, 16'd16103, 16'd32793, 16'd64905, 16'd209, 16'd24417, 16'd64450, 16'd41341, 16'd22437, 16'd47349, 16'd57422});
	test_expansion(128'h06d5b9c0d337a8af78920353cf1ada13, {16'd36210, 16'd61636, 16'd10839, 16'd42585, 16'd12994, 16'd34521, 16'd43913, 16'd15671, 16'd62032, 16'd4235, 16'd45932, 16'd46557, 16'd58035, 16'd27176, 16'd12437, 16'd59207, 16'd57122, 16'd53051, 16'd33891, 16'd46942, 16'd53532, 16'd51999, 16'd39812, 16'd63454, 16'd17920, 16'd14703});
	test_expansion(128'h1cbd1c68fda63ff29b3e2b28aa2b9e4f, {16'd29955, 16'd64998, 16'd6674, 16'd11926, 16'd41757, 16'd1871, 16'd57000, 16'd55634, 16'd51811, 16'd4499, 16'd10375, 16'd54143, 16'd45675, 16'd23028, 16'd24163, 16'd43917, 16'd3824, 16'd35954, 16'd11494, 16'd10336, 16'd26905, 16'd61958, 16'd2764, 16'd7172, 16'd5771, 16'd64784});
	test_expansion(128'h8d727b86411004009f1caf7b26baee7f, {16'd14602, 16'd43156, 16'd65080, 16'd13386, 16'd7926, 16'd19057, 16'd10092, 16'd62898, 16'd56741, 16'd13439, 16'd54119, 16'd57099, 16'd43916, 16'd15312, 16'd59189, 16'd36918, 16'd9321, 16'd60039, 16'd38382, 16'd38892, 16'd51263, 16'd47888, 16'd41512, 16'd39936, 16'd9898, 16'd50594});
	test_expansion(128'h638f93fa025661b00b7baa7d74ff57e8, {16'd26302, 16'd41178, 16'd9498, 16'd63534, 16'd33207, 16'd2572, 16'd13415, 16'd11424, 16'd28215, 16'd48161, 16'd38531, 16'd35909, 16'd40488, 16'd52905, 16'd60843, 16'd33496, 16'd56949, 16'd34983, 16'd40570, 16'd28272, 16'd23546, 16'd34987, 16'd26620, 16'd56745, 16'd65027, 16'd31954});
	test_expansion(128'h01b6ffd1ca2ec4aee5cc536265497547, {16'd30057, 16'd21516, 16'd54364, 16'd23755, 16'd23918, 16'd55367, 16'd38970, 16'd62174, 16'd61168, 16'd36690, 16'd44326, 16'd54332, 16'd59145, 16'd40402, 16'd62436, 16'd32945, 16'd52483, 16'd63224, 16'd53071, 16'd15654, 16'd40340, 16'd7177, 16'd14441, 16'd9330, 16'd45890, 16'd51686});
	test_expansion(128'h28ead6f101f3d462f569f0265cb1a085, {16'd48043, 16'd30857, 16'd3622, 16'd54035, 16'd37299, 16'd39977, 16'd14598, 16'd50962, 16'd6829, 16'd17287, 16'd53065, 16'd62980, 16'd29895, 16'd35490, 16'd54900, 16'd52356, 16'd42354, 16'd62561, 16'd53908, 16'd27155, 16'd38293, 16'd23351, 16'd11033, 16'd31673, 16'd54364, 16'd24077});
	test_expansion(128'hf5d593fcc57352074eeec6765f8fb759, {16'd2283, 16'd29256, 16'd20345, 16'd16008, 16'd56340, 16'd17362, 16'd44575, 16'd32331, 16'd13041, 16'd44905, 16'd23368, 16'd60928, 16'd63031, 16'd59576, 16'd23229, 16'd7980, 16'd27866, 16'd12744, 16'd51467, 16'd23300, 16'd1427, 16'd59451, 16'd48962, 16'd19769, 16'd24808, 16'd28111});
	test_expansion(128'hdd658d333b5abdb5450dd799fc9439f2, {16'd13992, 16'd36581, 16'd56933, 16'd50648, 16'd47668, 16'd38218, 16'd30623, 16'd20349, 16'd19946, 16'd56406, 16'd6981, 16'd20818, 16'd39611, 16'd20043, 16'd53234, 16'd44553, 16'd4272, 16'd23026, 16'd18771, 16'd32460, 16'd51965, 16'd27217, 16'd59848, 16'd48195, 16'd51180, 16'd26291});
	test_expansion(128'h4e586f944c3dc57b6689e7112942d118, {16'd2779, 16'd63529, 16'd20027, 16'd19141, 16'd6707, 16'd18474, 16'd34848, 16'd29926, 16'd65449, 16'd40761, 16'd11378, 16'd52771, 16'd10129, 16'd9503, 16'd3121, 16'd50029, 16'd5593, 16'd41572, 16'd32993, 16'd14446, 16'd60635, 16'd23267, 16'd64948, 16'd10365, 16'd50803, 16'd39003});
	test_expansion(128'hccb9d7cc4ff28266a60d6a1c331ee227, {16'd23090, 16'd33131, 16'd50388, 16'd65428, 16'd13514, 16'd15538, 16'd11426, 16'd55224, 16'd40511, 16'd23118, 16'd9311, 16'd43714, 16'd13007, 16'd6834, 16'd19387, 16'd59757, 16'd29293, 16'd25147, 16'd24643, 16'd16341, 16'd31172, 16'd60360, 16'd28143, 16'd19447, 16'd20887, 16'd37488});
	test_expansion(128'h2196b83f3df4bba80823a77a267632db, {16'd47571, 16'd50044, 16'd4595, 16'd64818, 16'd60682, 16'd43079, 16'd14953, 16'd51231, 16'd44476, 16'd64928, 16'd28697, 16'd20244, 16'd59705, 16'd62911, 16'd64275, 16'd38241, 16'd33875, 16'd1456, 16'd18533, 16'd29728, 16'd11223, 16'd37178, 16'd62552, 16'd33488, 16'd54650, 16'd13177});
	test_expansion(128'hb59acfbc029f0a1de0701cb228bffe87, {16'd21819, 16'd31493, 16'd27510, 16'd22863, 16'd24411, 16'd45537, 16'd45934, 16'd20252, 16'd36061, 16'd38848, 16'd16868, 16'd6296, 16'd20929, 16'd4409, 16'd28913, 16'd49788, 16'd13997, 16'd6403, 16'd16507, 16'd20371, 16'd11523, 16'd45578, 16'd50307, 16'd43571, 16'd15179, 16'd11967});
	test_expansion(128'h3fc1cfcd7bd05d3a9ff890fed67931d4, {16'd35281, 16'd47743, 16'd37451, 16'd59182, 16'd20613, 16'd18718, 16'd31514, 16'd50485, 16'd52176, 16'd16762, 16'd25685, 16'd13958, 16'd11027, 16'd30808, 16'd22937, 16'd32542, 16'd61572, 16'd19782, 16'd44235, 16'd65108, 16'd9740, 16'd21596, 16'd40686, 16'd11184, 16'd4417, 16'd46494});
	test_expansion(128'h2bdb09a95a2028c547a0699184ff616d, {16'd37397, 16'd2803, 16'd57233, 16'd47960, 16'd31929, 16'd27214, 16'd10393, 16'd57245, 16'd49018, 16'd36810, 16'd39191, 16'd62808, 16'd39617, 16'd53344, 16'd15281, 16'd13532, 16'd29977, 16'd29886, 16'd36924, 16'd50706, 16'd28168, 16'd14462, 16'd31517, 16'd3796, 16'd27423, 16'd41112});
	test_expansion(128'h473df9bc29168422796ada06d4b8b8e0, {16'd48009, 16'd24879, 16'd33802, 16'd48145, 16'd28507, 16'd3795, 16'd52468, 16'd52016, 16'd56453, 16'd8272, 16'd57025, 16'd62926, 16'd29997, 16'd23681, 16'd59973, 16'd52991, 16'd61163, 16'd8285, 16'd47893, 16'd48504, 16'd49813, 16'd57403, 16'd33048, 16'd51421, 16'd6884, 16'd5226});
	test_expansion(128'h6c971b40dd9b36d0725f9d157129d97a, {16'd28959, 16'd36521, 16'd15235, 16'd21109, 16'd51396, 16'd63710, 16'd56631, 16'd62111, 16'd46875, 16'd43729, 16'd18549, 16'd27367, 16'd15227, 16'd59182, 16'd29567, 16'd37060, 16'd49168, 16'd9778, 16'd39226, 16'd3029, 16'd22986, 16'd7793, 16'd58719, 16'd23093, 16'd36729, 16'd25156});
	test_expansion(128'h0bdf3f05a393984d6e7a6790987c73cc, {16'd54852, 16'd38453, 16'd24747, 16'd61699, 16'd20009, 16'd54277, 16'd25392, 16'd53919, 16'd37586, 16'd634, 16'd50177, 16'd16447, 16'd518, 16'd42568, 16'd40990, 16'd11315, 16'd28669, 16'd17170, 16'd3561, 16'd24297, 16'd18738, 16'd48233, 16'd20475, 16'd40188, 16'd32264, 16'd56740});
	test_expansion(128'hdd80942823e0ac7a21c1215bb94d0906, {16'd38868, 16'd16164, 16'd36989, 16'd56162, 16'd14076, 16'd17750, 16'd13599, 16'd23599, 16'd40658, 16'd32873, 16'd19613, 16'd11589, 16'd47382, 16'd12070, 16'd52007, 16'd47208, 16'd3011, 16'd36606, 16'd31979, 16'd3781, 16'd265, 16'd28952, 16'd38750, 16'd41643, 16'd53255, 16'd65303});
	test_expansion(128'h18cc42fd76b0fd3c977eecdaa86b713c, {16'd26160, 16'd26840, 16'd22245, 16'd5489, 16'd346, 16'd21437, 16'd50216, 16'd61541, 16'd47949, 16'd31546, 16'd55565, 16'd46173, 16'd41118, 16'd5149, 16'd22617, 16'd54791, 16'd22784, 16'd55954, 16'd55078, 16'd12435, 16'd16677, 16'd34591, 16'd38077, 16'd38648, 16'd61937, 16'd38571});
	test_expansion(128'hfc254fc6cdaa906ab7c827118737cf89, {16'd59578, 16'd7262, 16'd48931, 16'd29744, 16'd47199, 16'd33973, 16'd64382, 16'd20309, 16'd20817, 16'd34988, 16'd61142, 16'd53767, 16'd40984, 16'd4224, 16'd38856, 16'd65273, 16'd8597, 16'd59983, 16'd37698, 16'd44949, 16'd57787, 16'd59552, 16'd26860, 16'd40056, 16'd29939, 16'd60195});
	test_expansion(128'h651aa97bad98c90b9b2ee41232535369, {16'd13043, 16'd28151, 16'd51617, 16'd62386, 16'd7088, 16'd47608, 16'd36175, 16'd35180, 16'd44788, 16'd1726, 16'd56437, 16'd58363, 16'd5146, 16'd57984, 16'd38073, 16'd25720, 16'd40532, 16'd15943, 16'd22784, 16'd15493, 16'd53019, 16'd11097, 16'd21379, 16'd46369, 16'd59483, 16'd11047});
	test_expansion(128'h48968ac3e4932e6d4983bf767e7763ea, {16'd40695, 16'd63057, 16'd51981, 16'd10918, 16'd43046, 16'd28360, 16'd50062, 16'd9387, 16'd3461, 16'd56304, 16'd46004, 16'd64699, 16'd3315, 16'd28965, 16'd12527, 16'd28726, 16'd58969, 16'd40187, 16'd32268, 16'd60815, 16'd10281, 16'd25, 16'd1780, 16'd58321, 16'd32713, 16'd41669});
	test_expansion(128'h5643e1a12d98ff97b52491f1c3438dee, {16'd1511, 16'd57726, 16'd19094, 16'd967, 16'd15552, 16'd8144, 16'd46563, 16'd59747, 16'd41293, 16'd2295, 16'd9513, 16'd25562, 16'd10541, 16'd22650, 16'd56143, 16'd13136, 16'd20956, 16'd1391, 16'd30847, 16'd18051, 16'd38477, 16'd1402, 16'd31287, 16'd63516, 16'd58073, 16'd13873});
	test_expansion(128'h0649e1c5dba397825e48d72a617a9bd7, {16'd13928, 16'd2746, 16'd11744, 16'd25295, 16'd53531, 16'd60255, 16'd52644, 16'd6576, 16'd12023, 16'd23921, 16'd24832, 16'd25720, 16'd61721, 16'd20588, 16'd12941, 16'd39915, 16'd55060, 16'd7758, 16'd11856, 16'd48816, 16'd17178, 16'd52226, 16'd5756, 16'd27822, 16'd48129, 16'd18087});
	test_expansion(128'h5d8c89604a03018dbbda1c9a0c860c36, {16'd24786, 16'd42579, 16'd47743, 16'd52089, 16'd28808, 16'd61150, 16'd6228, 16'd64296, 16'd7988, 16'd51507, 16'd40920, 16'd58786, 16'd55922, 16'd33098, 16'd25288, 16'd45609, 16'd12699, 16'd27012, 16'd53132, 16'd17736, 16'd60387, 16'd15366, 16'd44796, 16'd40255, 16'd44627, 16'd43631});
	test_expansion(128'h9dd33e6542a7609ab5be12e6658924da, {16'd63484, 16'd45778, 16'd20579, 16'd32694, 16'd61553, 16'd48618, 16'd53497, 16'd17796, 16'd51428, 16'd21400, 16'd32973, 16'd63910, 16'd26758, 16'd11466, 16'd38851, 16'd6791, 16'd23139, 16'd37511, 16'd8780, 16'd15493, 16'd43569, 16'd25719, 16'd53556, 16'd5481, 16'd33156, 16'd55590});
	test_expansion(128'hf9bb1dff2755c281fcdd3d9913e34525, {16'd38604, 16'd36581, 16'd52110, 16'd13665, 16'd41680, 16'd27606, 16'd18030, 16'd63007, 16'd45543, 16'd40936, 16'd13889, 16'd14484, 16'd29297, 16'd60398, 16'd58048, 16'd16784, 16'd57329, 16'd60799, 16'd37035, 16'd61173, 16'd34576, 16'd46143, 16'd51063, 16'd36951, 16'd3050, 16'd50485});
	test_expansion(128'hf6ecec17e7e4f71f769d462f96a2130d, {16'd26005, 16'd22130, 16'd30717, 16'd36424, 16'd39983, 16'd50686, 16'd63064, 16'd18535, 16'd21898, 16'd34578, 16'd55748, 16'd8887, 16'd17063, 16'd43967, 16'd59925, 16'd8697, 16'd30070, 16'd13036, 16'd1590, 16'd15959, 16'd20082, 16'd54997, 16'd43584, 16'd3850, 16'd48349, 16'd14303});
	test_expansion(128'h5f033e5e4b8bbb30805f5a6b9d816774, {16'd3960, 16'd6434, 16'd48855, 16'd15621, 16'd22789, 16'd7544, 16'd28010, 16'd63073, 16'd2419, 16'd55486, 16'd26620, 16'd2231, 16'd7505, 16'd18868, 16'd9074, 16'd57154, 16'd57560, 16'd37472, 16'd42930, 16'd36326, 16'd1061, 16'd46147, 16'd8020, 16'd5275, 16'd26267, 16'd24917});
	test_expansion(128'hbf6bd6d4603bab12dc55eea2a1a983f2, {16'd9620, 16'd36703, 16'd24174, 16'd9601, 16'd45031, 16'd13026, 16'd50202, 16'd3528, 16'd40308, 16'd34805, 16'd8505, 16'd37884, 16'd17239, 16'd6332, 16'd39522, 16'd18298, 16'd15229, 16'd49104, 16'd4533, 16'd29737, 16'd50475, 16'd14952, 16'd26136, 16'd9679, 16'd46286, 16'd53148});
	test_expansion(128'h058e5136d46882cad431937ff3b7f86c, {16'd19818, 16'd61418, 16'd38152, 16'd13304, 16'd20312, 16'd40294, 16'd19301, 16'd29224, 16'd38738, 16'd53880, 16'd38999, 16'd55818, 16'd5378, 16'd12061, 16'd63736, 16'd35919, 16'd62286, 16'd38596, 16'd37100, 16'd20157, 16'd14131, 16'd20450, 16'd56294, 16'd41360, 16'd42589, 16'd40289});
	test_expansion(128'h2a2de0fb08691a46acb051055f6d109e, {16'd44159, 16'd19591, 16'd46259, 16'd40097, 16'd5558, 16'd51349, 16'd2783, 16'd22482, 16'd29364, 16'd1628, 16'd53195, 16'd59209, 16'd46662, 16'd57595, 16'd15666, 16'd4196, 16'd45768, 16'd11972, 16'd62030, 16'd39030, 16'd5982, 16'd3986, 16'd10078, 16'd11506, 16'd38730, 16'd10197});
	test_expansion(128'hacff8a213d040f06f1e72e10fad625cc, {16'd55853, 16'd38367, 16'd33651, 16'd43377, 16'd39913, 16'd40847, 16'd41975, 16'd61113, 16'd39418, 16'd48552, 16'd1796, 16'd25059, 16'd8992, 16'd33897, 16'd11080, 16'd34739, 16'd43793, 16'd34101, 16'd8406, 16'd1998, 16'd60002, 16'd2942, 16'd29776, 16'd55626, 16'd48893, 16'd24102});
	test_expansion(128'he13a01d6b19a9d267cae7be077b05114, {16'd28398, 16'd42493, 16'd24738, 16'd49072, 16'd53095, 16'd5445, 16'd52451, 16'd42336, 16'd38846, 16'd20381, 16'd21846, 16'd22113, 16'd23259, 16'd30826, 16'd45013, 16'd53642, 16'd64614, 16'd7928, 16'd32774, 16'd10141, 16'd46894, 16'd30748, 16'd48644, 16'd2180, 16'd15170, 16'd20036});
	test_expansion(128'h17d1103d779dfef0d3313b2ccbac764e, {16'd19708, 16'd29200, 16'd46756, 16'd45717, 16'd31103, 16'd16649, 16'd38045, 16'd3149, 16'd2210, 16'd30703, 16'd52066, 16'd36139, 16'd45656, 16'd34234, 16'd42036, 16'd27074, 16'd13329, 16'd7952, 16'd65243, 16'd1717, 16'd30387, 16'd55021, 16'd64599, 16'd55219, 16'd24974, 16'd54334});
	test_expansion(128'h657bc180b0ae871ad2b2abe78ba7e6fb, {16'd5972, 16'd53251, 16'd59047, 16'd49018, 16'd48410, 16'd12600, 16'd33770, 16'd15899, 16'd1971, 16'd20520, 16'd43723, 16'd58049, 16'd15316, 16'd55021, 16'd35081, 16'd59719, 16'd37371, 16'd5179, 16'd1250, 16'd52493, 16'd9166, 16'd22109, 16'd17088, 16'd873, 16'd19535, 16'd63859});
	test_expansion(128'hb14d38e400470e19d8e7215266be4281, {16'd12838, 16'd253, 16'd23010, 16'd60077, 16'd27582, 16'd50726, 16'd49174, 16'd44454, 16'd20886, 16'd26761, 16'd44703, 16'd48786, 16'd57994, 16'd524, 16'd4998, 16'd60190, 16'd28222, 16'd18120, 16'd54635, 16'd63700, 16'd2347, 16'd63876, 16'd58350, 16'd7710, 16'd24986, 16'd9055});
	test_expansion(128'hea49569780faf0c5e8b367fc7d0f0a79, {16'd60376, 16'd25816, 16'd59630, 16'd41781, 16'd23543, 16'd21625, 16'd28674, 16'd13992, 16'd35024, 16'd35498, 16'd772, 16'd31923, 16'd50188, 16'd2235, 16'd5563, 16'd31261, 16'd12474, 16'd27725, 16'd35876, 16'd49996, 16'd30472, 16'd41295, 16'd33212, 16'd21716, 16'd13072, 16'd55335});
	test_expansion(128'h79a86e3bbcdf8d3e5baf7f261177279e, {16'd11153, 16'd36348, 16'd49759, 16'd45987, 16'd3650, 16'd50621, 16'd27538, 16'd30354, 16'd45432, 16'd49327, 16'd2022, 16'd10539, 16'd58438, 16'd15026, 16'd21952, 16'd46389, 16'd46717, 16'd9941, 16'd42876, 16'd47632, 16'd42148, 16'd8016, 16'd54133, 16'd46470, 16'd45364, 16'd48567});
	test_expansion(128'h67498f4dcb88db57c4bde6f098f856d6, {16'd11953, 16'd48880, 16'd28754, 16'd14940, 16'd29336, 16'd32288, 16'd5325, 16'd8791, 16'd14989, 16'd43759, 16'd43234, 16'd48842, 16'd26599, 16'd5513, 16'd54213, 16'd7138, 16'd18302, 16'd41232, 16'd51914, 16'd14057, 16'd8898, 16'd29293, 16'd18905, 16'd61312, 16'd18118, 16'd59722});
	test_expansion(128'h7b05d6329b447ffbabe34767027deb26, {16'd45673, 16'd30294, 16'd39222, 16'd9128, 16'd26910, 16'd48350, 16'd55611, 16'd21069, 16'd45754, 16'd57612, 16'd6844, 16'd44694, 16'd12929, 16'd11646, 16'd64576, 16'd16515, 16'd58434, 16'd26727, 16'd54325, 16'd22507, 16'd37246, 16'd26689, 16'd13036, 16'd4541, 16'd42752, 16'd11008});
	test_expansion(128'hbd25194008712492b680316251e8971d, {16'd13522, 16'd64480, 16'd12654, 16'd59561, 16'd35224, 16'd53599, 16'd59038, 16'd16149, 16'd43454, 16'd2203, 16'd24656, 16'd16799, 16'd21117, 16'd34380, 16'd61955, 16'd62403, 16'd8403, 16'd3235, 16'd55461, 16'd55556, 16'd48725, 16'd46808, 16'd48736, 16'd59218, 16'd44267, 16'd13236});
	test_expansion(128'h7d0cbf26eb1c8ab1dcc0e8bdeb2ee9d9, {16'd42221, 16'd6832, 16'd51624, 16'd20915, 16'd21181, 16'd14803, 16'd9329, 16'd10314, 16'd56076, 16'd10135, 16'd47776, 16'd63459, 16'd22170, 16'd272, 16'd31587, 16'd15942, 16'd18438, 16'd11279, 16'd6782, 16'd6402, 16'd47212, 16'd57734, 16'd20902, 16'd55498, 16'd56456, 16'd48547});
	test_expansion(128'h3dcb042c0619cf5103d3bee01d8d2c02, {16'd35407, 16'd3531, 16'd25871, 16'd60969, 16'd23842, 16'd19255, 16'd33546, 16'd4310, 16'd20013, 16'd16990, 16'd63852, 16'd46979, 16'd44135, 16'd13010, 16'd53743, 16'd24923, 16'd61822, 16'd16469, 16'd49004, 16'd37579, 16'd27866, 16'd59607, 16'd29971, 16'd37372, 16'd50401, 16'd39741});
	test_expansion(128'h4b4ee68ae8ba5c0d4819577c19eca99a, {16'd49902, 16'd23558, 16'd39022, 16'd60037, 16'd10270, 16'd52048, 16'd56033, 16'd8003, 16'd13581, 16'd11970, 16'd53750, 16'd36778, 16'd37384, 16'd14686, 16'd39561, 16'd35451, 16'd47170, 16'd47061, 16'd17571, 16'd56347, 16'd47696, 16'd1817, 16'd25620, 16'd25135, 16'd28415, 16'd28921});
	test_expansion(128'h3569f9129e0724319083ed3ec31e8e26, {16'd32805, 16'd61288, 16'd59928, 16'd19799, 16'd47032, 16'd56491, 16'd15653, 16'd33408, 16'd42321, 16'd1078, 16'd6740, 16'd17285, 16'd29202, 16'd536, 16'd46412, 16'd8851, 16'd17190, 16'd6223, 16'd575, 16'd41313, 16'd20442, 16'd33093, 16'd29516, 16'd29828, 16'd42828, 16'd9589});
	test_expansion(128'hee657fab02d095fe1d55de371f59e45d, {16'd49207, 16'd31940, 16'd57068, 16'd53988, 16'd6553, 16'd1073, 16'd53014, 16'd28672, 16'd35007, 16'd33825, 16'd61334, 16'd56886, 16'd59355, 16'd60333, 16'd29453, 16'd64911, 16'd1001, 16'd16876, 16'd43196, 16'd13079, 16'd2936, 16'd65512, 16'd14129, 16'd14286, 16'd35259, 16'd20154});
	test_expansion(128'he2971771681efe993db4bb945dcdef05, {16'd18867, 16'd17598, 16'd20520, 16'd51772, 16'd17846, 16'd22022, 16'd16246, 16'd39765, 16'd5379, 16'd41432, 16'd13364, 16'd11089, 16'd62794, 16'd7363, 16'd46790, 16'd9332, 16'd27266, 16'd8024, 16'd15903, 16'd30154, 16'd46469, 16'd40970, 16'd16478, 16'd9948, 16'd17843, 16'd38316});
	test_expansion(128'h30409cf5fd5dde4a78d042d8c2860cc0, {16'd11593, 16'd47998, 16'd9354, 16'd40107, 16'd43868, 16'd25732, 16'd48613, 16'd49000, 16'd45624, 16'd8519, 16'd33721, 16'd4430, 16'd19000, 16'd27264, 16'd27202, 16'd56708, 16'd52131, 16'd31219, 16'd43125, 16'd37542, 16'd39114, 16'd60781, 16'd64648, 16'd2735, 16'd38241, 16'd45516});
	test_expansion(128'h2c9295d13ec43a3871fbf472b49f4066, {16'd56375, 16'd5604, 16'd38510, 16'd3967, 16'd9216, 16'd18821, 16'd24648, 16'd52216, 16'd65312, 16'd33189, 16'd37265, 16'd7447, 16'd39949, 16'd25391, 16'd63543, 16'd3546, 16'd7404, 16'd44445, 16'd4176, 16'd46599, 16'd49169, 16'd50486, 16'd803, 16'd58120, 16'd49232, 16'd18379});
	test_expansion(128'h0784fca3191c86806e25098f00e9f517, {16'd17039, 16'd35123, 16'd19853, 16'd6673, 16'd63915, 16'd25251, 16'd35913, 16'd63414, 16'd21959, 16'd10559, 16'd41987, 16'd43646, 16'd50539, 16'd32106, 16'd65104, 16'd10134, 16'd20273, 16'd56851, 16'd48023, 16'd23746, 16'd31943, 16'd17066, 16'd8997, 16'd63385, 16'd59268, 16'd59802});
	test_expansion(128'h86406af6b64b63d3c348ce2887119407, {16'd13225, 16'd21305, 16'd29198, 16'd7252, 16'd46921, 16'd12653, 16'd34274, 16'd9728, 16'd46493, 16'd51639, 16'd1109, 16'd10413, 16'd61669, 16'd60800, 16'd47811, 16'd11362, 16'd43217, 16'd5771, 16'd5294, 16'd10443, 16'd31394, 16'd45966, 16'd22763, 16'd19507, 16'd56099, 16'd38678});
	test_expansion(128'h729dc29a602f09ee3f3f5b3d6ff68aa5, {16'd11137, 16'd65078, 16'd44147, 16'd39021, 16'd41689, 16'd24934, 16'd25526, 16'd49883, 16'd29921, 16'd6228, 16'd19097, 16'd56505, 16'd37726, 16'd7022, 16'd50323, 16'd51981, 16'd48329, 16'd32809, 16'd38959, 16'd65044, 16'd18770, 16'd18737, 16'd49878, 16'd64263, 16'd18864, 16'd10157});
	test_expansion(128'h451423a595562d28b62a8557499f909a, {16'd13074, 16'd63720, 16'd58965, 16'd49520, 16'd24330, 16'd6450, 16'd52821, 16'd41094, 16'd46471, 16'd719, 16'd46945, 16'd14076, 16'd37655, 16'd4515, 16'd62092, 16'd59524, 16'd24675, 16'd1488, 16'd60024, 16'd38889, 16'd13809, 16'd55068, 16'd914, 16'd63173, 16'd22665, 16'd58678});
	test_expansion(128'h1b560ed2bd3fa1df96f3fe7aaea8a03c, {16'd11510, 16'd27199, 16'd29337, 16'd11323, 16'd26725, 16'd61969, 16'd62876, 16'd59139, 16'd44573, 16'd18839, 16'd26036, 16'd12944, 16'd56760, 16'd60284, 16'd64542, 16'd42343, 16'd49489, 16'd46943, 16'd30778, 16'd27448, 16'd61546, 16'd878, 16'd47845, 16'd4652, 16'd49608, 16'd39037});
	test_expansion(128'he92c556eec62732ea52c97dc01c90f62, {16'd62269, 16'd29127, 16'd34243, 16'd57795, 16'd61587, 16'd11425, 16'd381, 16'd56195, 16'd55597, 16'd21135, 16'd44301, 16'd40636, 16'd26198, 16'd58684, 16'd60511, 16'd37519, 16'd52280, 16'd13554, 16'd37369, 16'd33467, 16'd34363, 16'd22581, 16'd48797, 16'd404, 16'd5171, 16'd61582});
	test_expansion(128'h8c6b8ecc58fc45949094df05ffeaa378, {16'd48844, 16'd11323, 16'd18144, 16'd63460, 16'd16761, 16'd27457, 16'd30294, 16'd26268, 16'd25247, 16'd51531, 16'd6453, 16'd4502, 16'd11325, 16'd38451, 16'd55674, 16'd36046, 16'd39234, 16'd45112, 16'd16153, 16'd6228, 16'd21099, 16'd56229, 16'd10052, 16'd314, 16'd56830, 16'd6630});
	test_expansion(128'h6c924eef8952714d320062ef4623a4e9, {16'd56225, 16'd46949, 16'd17772, 16'd13538, 16'd22292, 16'd17138, 16'd8016, 16'd38397, 16'd11207, 16'd34883, 16'd54889, 16'd38686, 16'd7311, 16'd5801, 16'd30134, 16'd63432, 16'd61340, 16'd24770, 16'd64617, 16'd3068, 16'd24588, 16'd11232, 16'd36903, 16'd8955, 16'd56324, 16'd62172});
	test_expansion(128'h4c871851e39428a2c35936e742411c06, {16'd20752, 16'd37495, 16'd37869, 16'd38135, 16'd59006, 16'd53998, 16'd22253, 16'd40996, 16'd30639, 16'd7430, 16'd55290, 16'd35210, 16'd9796, 16'd31489, 16'd43019, 16'd35146, 16'd3235, 16'd16503, 16'd24149, 16'd45060, 16'd15884, 16'd64006, 16'd38443, 16'd5943, 16'd27642, 16'd55308});
	test_expansion(128'h1df6ff8bdac6a9c6680afc5693df7406, {16'd36857, 16'd20420, 16'd23630, 16'd18825, 16'd39795, 16'd27358, 16'd33033, 16'd16572, 16'd24672, 16'd12898, 16'd32029, 16'd63068, 16'd1302, 16'd47796, 16'd13553, 16'd33735, 16'd12200, 16'd8093, 16'd20705, 16'd54234, 16'd42529, 16'd60168, 16'd1207, 16'd5693, 16'd32618, 16'd12914});
	test_expansion(128'h6c242e1d7e131a527d1b66d70b820f6e, {16'd30521, 16'd29991, 16'd55215, 16'd57179, 16'd46364, 16'd32572, 16'd19403, 16'd34055, 16'd47487, 16'd2496, 16'd57559, 16'd59228, 16'd13197, 16'd24509, 16'd23773, 16'd16703, 16'd43382, 16'd7229, 16'd42005, 16'd31257, 16'd31314, 16'd4188, 16'd33881, 16'd4504, 16'd3911, 16'd59460});
	test_expansion(128'h354dabd3deed45aa3c7fc66bcde6d75c, {16'd12069, 16'd56150, 16'd31024, 16'd42103, 16'd36022, 16'd41765, 16'd16415, 16'd27112, 16'd9650, 16'd19855, 16'd29724, 16'd236, 16'd27874, 16'd12257, 16'd15935, 16'd54479, 16'd59715, 16'd48113, 16'd5669, 16'd31358, 16'd56651, 16'd50220, 16'd28430, 16'd2205, 16'd12052, 16'd49284});
	test_expansion(128'hb53b180458ffb413cc00192319b2967c, {16'd5438, 16'd9082, 16'd59093, 16'd473, 16'd10692, 16'd35498, 16'd47949, 16'd18325, 16'd19038, 16'd5340, 16'd48108, 16'd16196, 16'd52931, 16'd63536, 16'd24620, 16'd49637, 16'd11204, 16'd38914, 16'd46683, 16'd9642, 16'd40235, 16'd64483, 16'd46439, 16'd2751, 16'd58814, 16'd62743});
	test_expansion(128'h0807a3164c96453e9e9a52258e0688fd, {16'd52251, 16'd28810, 16'd64244, 16'd9503, 16'd9054, 16'd4311, 16'd54450, 16'd38013, 16'd47091, 16'd30774, 16'd52546, 16'd17442, 16'd65089, 16'd1713, 16'd55909, 16'd12534, 16'd43605, 16'd46810, 16'd65521, 16'd13992, 16'd28392, 16'd64316, 16'd53673, 16'd63593, 16'd54233, 16'd5586});
	test_expansion(128'h46f56f34eabb86235b7129ef9729ebcc, {16'd20444, 16'd1300, 16'd37703, 16'd29611, 16'd32083, 16'd30192, 16'd63188, 16'd16248, 16'd27532, 16'd60004, 16'd19881, 16'd20570, 16'd53639, 16'd26357, 16'd45505, 16'd50724, 16'd54616, 16'd786, 16'd62504, 16'd47833, 16'd36258, 16'd54116, 16'd41448, 16'd11997, 16'd28324, 16'd21442});
	test_expansion(128'hd400dd35d8d279cbb99235579d2a5e63, {16'd25557, 16'd33375, 16'd24816, 16'd47060, 16'd21343, 16'd37407, 16'd12474, 16'd17452, 16'd23689, 16'd44692, 16'd44335, 16'd54844, 16'd60453, 16'd62685, 16'd30398, 16'd50146, 16'd46200, 16'd29217, 16'd59754, 16'd4245, 16'd13797, 16'd42996, 16'd49931, 16'd12930, 16'd33405, 16'd37325});
	test_expansion(128'h8971ac6d1dd37e2439666b6ea1deeaf4, {16'd697, 16'd63306, 16'd28260, 16'd52963, 16'd29094, 16'd1267, 16'd25254, 16'd8744, 16'd8220, 16'd11241, 16'd53950, 16'd35599, 16'd60555, 16'd8201, 16'd36949, 16'd10590, 16'd60974, 16'd52330, 16'd10941, 16'd25792, 16'd25715, 16'd53680, 16'd28026, 16'd39091, 16'd32162, 16'd26272});
	test_expansion(128'hc47ede729d550da13390d56c7580e9f2, {16'd61433, 16'd10875, 16'd52816, 16'd22462, 16'd53404, 16'd37148, 16'd38031, 16'd24914, 16'd59437, 16'd3327, 16'd26276, 16'd41370, 16'd24775, 16'd1439, 16'd19596, 16'd38504, 16'd19286, 16'd5714, 16'd16682, 16'd11037, 16'd20605, 16'd26330, 16'd8826, 16'd38342, 16'd13930, 16'd56638});
	test_expansion(128'h3c1b2f95842e5d4ac52d2cb0603bf486, {16'd56705, 16'd7160, 16'd60705, 16'd27908, 16'd10182, 16'd24766, 16'd53046, 16'd61087, 16'd10310, 16'd32351, 16'd42411, 16'd49214, 16'd61339, 16'd16695, 16'd4080, 16'd57824, 16'd59033, 16'd57427, 16'd47985, 16'd46890, 16'd5537, 16'd54533, 16'd42710, 16'd13561, 16'd51234, 16'd27577});
	test_expansion(128'hd7d0f4cd5c1616c203bfa02ffc87768b, {16'd44140, 16'd61330, 16'd2697, 16'd11444, 16'd36464, 16'd35521, 16'd10138, 16'd30272, 16'd26123, 16'd15506, 16'd15911, 16'd28186, 16'd31302, 16'd21635, 16'd20934, 16'd21189, 16'd24384, 16'd30579, 16'd43601, 16'd24151, 16'd57761, 16'd32453, 16'd29966, 16'd55931, 16'd54184, 16'd59592});
	test_expansion(128'hd53cc95deb6bf006df7ce58b691aea60, {16'd18227, 16'd24050, 16'd5763, 16'd48425, 16'd36129, 16'd51769, 16'd14971, 16'd36374, 16'd1079, 16'd47579, 16'd2419, 16'd16070, 16'd31964, 16'd44967, 16'd32022, 16'd32270, 16'd64836, 16'd5504, 16'd51750, 16'd11924, 16'd60224, 16'd52970, 16'd40021, 16'd22288, 16'd45989, 16'd52220});
	test_expansion(128'h7c4cae703209c8b5b4272e150e2a9695, {16'd48527, 16'd51705, 16'd35706, 16'd50444, 16'd65243, 16'd64549, 16'd50052, 16'd30384, 16'd52676, 16'd57245, 16'd51254, 16'd24888, 16'd42776, 16'd26803, 16'd59094, 16'd32280, 16'd1828, 16'd1782, 16'd8803, 16'd37987, 16'd6815, 16'd12264, 16'd32631, 16'd5691, 16'd42651, 16'd25976});
	test_expansion(128'h0b746d0c53f962bbd4c3c97a84a25fd2, {16'd19490, 16'd52356, 16'd30748, 16'd44679, 16'd24380, 16'd20595, 16'd61711, 16'd53009, 16'd6932, 16'd19808, 16'd43055, 16'd31944, 16'd36612, 16'd30094, 16'd37331, 16'd41468, 16'd28838, 16'd46983, 16'd26648, 16'd64583, 16'd37993, 16'd59788, 16'd32927, 16'd50887, 16'd14783, 16'd31180});
	test_expansion(128'hd16eab58ec7f3261adc0cab4d2c4bdba, {16'd1403, 16'd16810, 16'd21540, 16'd49635, 16'd27525, 16'd20067, 16'd33540, 16'd19890, 16'd27042, 16'd21368, 16'd37876, 16'd52593, 16'd31880, 16'd21876, 16'd42888, 16'd17373, 16'd37173, 16'd21666, 16'd41878, 16'd842, 16'd58341, 16'd41878, 16'd50892, 16'd54789, 16'd15797, 16'd62269});
	test_expansion(128'h40709f5dabafd10835b1c7d2fd13e64f, {16'd31169, 16'd45545, 16'd14154, 16'd53129, 16'd62453, 16'd62353, 16'd58630, 16'd25635, 16'd40532, 16'd19119, 16'd30057, 16'd37870, 16'd34063, 16'd49597, 16'd5014, 16'd25855, 16'd53528, 16'd17498, 16'd3134, 16'd25619, 16'd17413, 16'd59778, 16'd15053, 16'd3109, 16'd23059, 16'd6101});
	test_expansion(128'h721bd4e66793380cbe02f61a1a349756, {16'd64081, 16'd59242, 16'd54285, 16'd60775, 16'd51853, 16'd40498, 16'd42511, 16'd48402, 16'd31288, 16'd9684, 16'd54439, 16'd42521, 16'd37479, 16'd63534, 16'd3622, 16'd27247, 16'd63931, 16'd225, 16'd41918, 16'd18194, 16'd10732, 16'd59385, 16'd9437, 16'd18666, 16'd42850, 16'd27883});
	test_expansion(128'hc70d5e8642ed346b56b0b4563b3a7207, {16'd19310, 16'd6578, 16'd23288, 16'd65074, 16'd7405, 16'd47036, 16'd29229, 16'd3646, 16'd1651, 16'd14450, 16'd62445, 16'd27923, 16'd3261, 16'd36348, 16'd49653, 16'd17545, 16'd56007, 16'd16807, 16'd55444, 16'd7228, 16'd56252, 16'd53819, 16'd38793, 16'd56456, 16'd5873, 16'd11547});
	test_expansion(128'h518165d7ad37f0f70508a20d523936a5, {16'd41727, 16'd55573, 16'd25225, 16'd45303, 16'd4835, 16'd27501, 16'd19315, 16'd3987, 16'd25094, 16'd58015, 16'd1240, 16'd13949, 16'd23885, 16'd14136, 16'd27825, 16'd18444, 16'd56653, 16'd37736, 16'd51298, 16'd30184, 16'd57335, 16'd19780, 16'd53851, 16'd16698, 16'd23695, 16'd52601});
	test_expansion(128'ha28ea63e2e841164893ab77fe2aa9a9c, {16'd29314, 16'd48087, 16'd18848, 16'd59122, 16'd60948, 16'd61268, 16'd34495, 16'd36267, 16'd41356, 16'd36195, 16'd29368, 16'd58028, 16'd30899, 16'd44686, 16'd39500, 16'd48700, 16'd13137, 16'd41666, 16'd16871, 16'd3007, 16'd1559, 16'd59842, 16'd11490, 16'd384, 16'd35889, 16'd59798});
	test_expansion(128'h16021bcea725530881a47cc98b13ca04, {16'd58434, 16'd9441, 16'd37595, 16'd60442, 16'd21894, 16'd9779, 16'd45615, 16'd33341, 16'd19409, 16'd28497, 16'd18801, 16'd22803, 16'd9027, 16'd20521, 16'd30235, 16'd65172, 16'd9615, 16'd63282, 16'd15466, 16'd12462, 16'd28317, 16'd22422, 16'd8380, 16'd27049, 16'd31147, 16'd1823});
	test_expansion(128'hb285918ddab8fa9776282e08939b12e2, {16'd54936, 16'd33556, 16'd32986, 16'd61638, 16'd31764, 16'd13913, 16'd50405, 16'd41842, 16'd33067, 16'd6314, 16'd21046, 16'd50776, 16'd35217, 16'd45081, 16'd45506, 16'd31144, 16'd24664, 16'd19615, 16'd20278, 16'd34200, 16'd21114, 16'd2500, 16'd15720, 16'd48664, 16'd61427, 16'd29290});
	test_expansion(128'h1e0b3ea358bbd09921ed8de74b122277, {16'd45607, 16'd21637, 16'd63657, 16'd45851, 16'd21987, 16'd9273, 16'd13737, 16'd1232, 16'd34655, 16'd40057, 16'd52827, 16'd21671, 16'd58933, 16'd57041, 16'd34569, 16'd49114, 16'd19013, 16'd50466, 16'd49776, 16'd51551, 16'd23580, 16'd58815, 16'd43151, 16'd31052, 16'd5235, 16'd21140});
	test_expansion(128'h93bf97e39ba453bd4886a8a94e77de92, {16'd48476, 16'd37138, 16'd16830, 16'd17923, 16'd27136, 16'd62492, 16'd51909, 16'd28863, 16'd13335, 16'd19840, 16'd31589, 16'd10172, 16'd61877, 16'd8849, 16'd56199, 16'd38121, 16'd26814, 16'd62687, 16'd63736, 16'd54574, 16'd2650, 16'd758, 16'd7047, 16'd28324, 16'd26000, 16'd42236});
	test_expansion(128'hce5f41370f783af303c5ac27d872d521, {16'd43555, 16'd50340, 16'd24475, 16'd53300, 16'd39604, 16'd38011, 16'd30391, 16'd49770, 16'd18774, 16'd3895, 16'd8479, 16'd1334, 16'd7036, 16'd27788, 16'd7339, 16'd50801, 16'd25688, 16'd48206, 16'd38251, 16'd19246, 16'd44009, 16'd27860, 16'd36494, 16'd13834, 16'd30515, 16'd6966});
	test_expansion(128'hade7ed8a413537828583ec4da4932907, {16'd60429, 16'd16015, 16'd14755, 16'd63126, 16'd21064, 16'd42712, 16'd795, 16'd9841, 16'd2428, 16'd1293, 16'd17493, 16'd41969, 16'd31719, 16'd49645, 16'd43102, 16'd23062, 16'd13029, 16'd62556, 16'd57656, 16'd13918, 16'd23303, 16'd41702, 16'd10692, 16'd19099, 16'd58109, 16'd23344});
	test_expansion(128'h94b5fd15d17ad02b74826636d3fbe6e9, {16'd58496, 16'd5797, 16'd22458, 16'd2455, 16'd24791, 16'd37498, 16'd40520, 16'd32746, 16'd31120, 16'd63224, 16'd49461, 16'd13890, 16'd17498, 16'd48671, 16'd49085, 16'd6011, 16'd40479, 16'd11450, 16'd19390, 16'd52112, 16'd54452, 16'd8383, 16'd51908, 16'd8287, 16'd60883, 16'd47810});
	test_expansion(128'hcc5645228f9f0d28c34edaee9a14a94f, {16'd45331, 16'd52796, 16'd20955, 16'd65081, 16'd60133, 16'd41067, 16'd36695, 16'd29888, 16'd15611, 16'd46732, 16'd23079, 16'd4715, 16'd25325, 16'd2811, 16'd7286, 16'd21874, 16'd63306, 16'd30473, 16'd36310, 16'd37160, 16'd17099, 16'd28523, 16'd18354, 16'd33644, 16'd48743, 16'd44108});
	test_expansion(128'h1d28bdcbe1f2b5e1acad0930d9789923, {16'd10509, 16'd721, 16'd231, 16'd15868, 16'd49765, 16'd395, 16'd55876, 16'd1869, 16'd51521, 16'd39281, 16'd8052, 16'd20457, 16'd50955, 16'd10088, 16'd14215, 16'd27580, 16'd11503, 16'd58120, 16'd44877, 16'd54939, 16'd364, 16'd34431, 16'd57156, 16'd43913, 16'd12415, 16'd31529});
	test_expansion(128'he3f7832427ffe5ccb498e9fd7b37bcc8, {16'd18827, 16'd54315, 16'd46856, 16'd45673, 16'd46761, 16'd6395, 16'd15042, 16'd53705, 16'd29454, 16'd2134, 16'd246, 16'd23446, 16'd26102, 16'd62532, 16'd38076, 16'd25615, 16'd14774, 16'd64553, 16'd28920, 16'd42629, 16'd30219, 16'd48094, 16'd38569, 16'd58549, 16'd9367, 16'd10082});
	test_expansion(128'h37b6e631cadcd754eb3c828350f4109b, {16'd65117, 16'd26607, 16'd17046, 16'd18508, 16'd26942, 16'd25384, 16'd52689, 16'd58950, 16'd25645, 16'd475, 16'd23124, 16'd45872, 16'd27520, 16'd43603, 16'd34541, 16'd34251, 16'd52996, 16'd18110, 16'd50415, 16'd26145, 16'd21406, 16'd13779, 16'd27086, 16'd55135, 16'd53991, 16'd7916});
	test_expansion(128'h6fbae35937eec4dc048c8306b933ae1d, {16'd6547, 16'd48079, 16'd47138, 16'd21860, 16'd1697, 16'd40767, 16'd27165, 16'd3350, 16'd52175, 16'd8548, 16'd46666, 16'd22793, 16'd3771, 16'd56158, 16'd41021, 16'd11224, 16'd26337, 16'd29235, 16'd32488, 16'd58023, 16'd23725, 16'd51383, 16'd11424, 16'd4480, 16'd32352, 16'd18313});
	test_expansion(128'h35c6cef22bf9e657aeee507e64c80d97, {16'd21787, 16'd23855, 16'd61659, 16'd23420, 16'd1286, 16'd52375, 16'd8659, 16'd9271, 16'd39688, 16'd31466, 16'd1353, 16'd18265, 16'd49125, 16'd26953, 16'd54768, 16'd25897, 16'd52253, 16'd36665, 16'd42358, 16'd4410, 16'd17122, 16'd29127, 16'd16682, 16'd41451, 16'd58527, 16'd9567});
	test_expansion(128'h55581ca57b47c00be935358f5e55a48f, {16'd39709, 16'd16303, 16'd2768, 16'd40450, 16'd36840, 16'd40608, 16'd28616, 16'd51314, 16'd47758, 16'd43863, 16'd16868, 16'd62324, 16'd38802, 16'd60497, 16'd5673, 16'd15255, 16'd27299, 16'd47219, 16'd45512, 16'd38846, 16'd14770, 16'd18415, 16'd29984, 16'd39663, 16'd21239, 16'd38401});
	test_expansion(128'h8453172675bb032fedd085bcb9a42801, {16'd40992, 16'd55843, 16'd22103, 16'd61162, 16'd55819, 16'd33265, 16'd27493, 16'd53945, 16'd37548, 16'd63600, 16'd5650, 16'd10503, 16'd23443, 16'd20042, 16'd249, 16'd11148, 16'd49759, 16'd63983, 16'd32498, 16'd50932, 16'd45172, 16'd47325, 16'd40901, 16'd32658, 16'd57865, 16'd43976});
	test_expansion(128'hc3528e8f27f2c918d1bf1e90fe009a11, {16'd43341, 16'd19062, 16'd27652, 16'd59697, 16'd51543, 16'd45023, 16'd44017, 16'd44289, 16'd10704, 16'd12341, 16'd34499, 16'd56992, 16'd52033, 16'd41056, 16'd57414, 16'd26767, 16'd3414, 16'd9112, 16'd48187, 16'd12805, 16'd65178, 16'd22742, 16'd62210, 16'd22970, 16'd24622, 16'd16201});
	test_expansion(128'hf538b470a40515174afd05c31c4c8444, {16'd55993, 16'd64371, 16'd42916, 16'd2574, 16'd29208, 16'd30566, 16'd55641, 16'd40776, 16'd8024, 16'd37978, 16'd18113, 16'd20402, 16'd1561, 16'd37648, 16'd54647, 16'd11398, 16'd734, 16'd5280, 16'd31910, 16'd58035, 16'd61524, 16'd34878, 16'd59756, 16'd62643, 16'd31730, 16'd1949});
	test_expansion(128'hff6ce805549125c22e55661fe7335db9, {16'd58819, 16'd65290, 16'd29314, 16'd52478, 16'd26099, 16'd27522, 16'd56911, 16'd32042, 16'd63816, 16'd21527, 16'd23650, 16'd31300, 16'd42950, 16'd56261, 16'd56115, 16'd15354, 16'd25138, 16'd8090, 16'd51785, 16'd48390, 16'd44615, 16'd9870, 16'd29570, 16'd62802, 16'd7436, 16'd46459});
	test_expansion(128'he8d9e10e9bce98b57dc2efe7005a6288, {16'd21661, 16'd60977, 16'd46273, 16'd63998, 16'd47095, 16'd54216, 16'd63214, 16'd24591, 16'd20094, 16'd64244, 16'd64649, 16'd380, 16'd50980, 16'd22020, 16'd46036, 16'd61973, 16'd40671, 16'd65528, 16'd50003, 16'd50600, 16'd13711, 16'd379, 16'd42184, 16'd12013, 16'd38214, 16'd45520});
	test_expansion(128'h149e5c2553e036b31fcf7b5431e8d416, {16'd65302, 16'd48502, 16'd52472, 16'd13168, 16'd60769, 16'd39866, 16'd50139, 16'd6465, 16'd6970, 16'd43540, 16'd1153, 16'd24764, 16'd731, 16'd10431, 16'd6641, 16'd54592, 16'd28937, 16'd516, 16'd35225, 16'd45356, 16'd41745, 16'd42826, 16'd48687, 16'd3963, 16'd46969, 16'd15403});
	test_expansion(128'h60e425a8de7f8c4ef868d22ee80aede2, {16'd34138, 16'd34080, 16'd3607, 16'd19385, 16'd8892, 16'd46675, 16'd8989, 16'd65027, 16'd43981, 16'd20948, 16'd3646, 16'd36670, 16'd65123, 16'd8793, 16'd64918, 16'd29755, 16'd626, 16'd45649, 16'd34584, 16'd42720, 16'd43670, 16'd49803, 16'd5830, 16'd23661, 16'd29861, 16'd15768});
	test_expansion(128'he792d14cbbe013166b3f4c06f61ca38e, {16'd62981, 16'd29689, 16'd2389, 16'd53543, 16'd37910, 16'd21390, 16'd37374, 16'd39390, 16'd12871, 16'd48903, 16'd45512, 16'd57054, 16'd51, 16'd9353, 16'd19587, 16'd36512, 16'd4568, 16'd15305, 16'd60281, 16'd32424, 16'd48853, 16'd53724, 16'd27312, 16'd31814, 16'd44047, 16'd6391});
	test_expansion(128'h7f0a955f982f08eaa4a5cb6f34620002, {16'd654, 16'd58430, 16'd54824, 16'd27045, 16'd12914, 16'd60092, 16'd12904, 16'd48820, 16'd30089, 16'd53474, 16'd28384, 16'd8650, 16'd22129, 16'd57134, 16'd51330, 16'd54936, 16'd46151, 16'd20049, 16'd28699, 16'd55359, 16'd37075, 16'd64762, 16'd4846, 16'd31574, 16'd95, 16'd31697});
	test_expansion(128'h73f2e75090839e57fb4f49c724c1e344, {16'd53666, 16'd47214, 16'd8754, 16'd63290, 16'd44658, 16'd29730, 16'd42109, 16'd34002, 16'd41593, 16'd54076, 16'd20469, 16'd28910, 16'd58743, 16'd1247, 16'd29213, 16'd3303, 16'd28702, 16'd30282, 16'd61978, 16'd13111, 16'd32763, 16'd10745, 16'd38318, 16'd16355, 16'd49832, 16'd14749});
	test_expansion(128'hb7b5714285941841145fda9e721dec03, {16'd44333, 16'd59513, 16'd18390, 16'd13598, 16'd54358, 16'd43030, 16'd8834, 16'd8895, 16'd10989, 16'd32030, 16'd41197, 16'd17406, 16'd64006, 16'd25909, 16'd13857, 16'd60656, 16'd34775, 16'd34479, 16'd48880, 16'd10678, 16'd43194, 16'd26655, 16'd44607, 16'd45658, 16'd14906, 16'd39055});
	test_expansion(128'hf873b12c257fe9d38fa650a0dbf5dd89, {16'd39289, 16'd1494, 16'd48038, 16'd25852, 16'd32259, 16'd18182, 16'd6906, 16'd37083, 16'd37902, 16'd19414, 16'd24506, 16'd15905, 16'd27029, 16'd26015, 16'd16883, 16'd20737, 16'd34473, 16'd39818, 16'd32133, 16'd37637, 16'd59663, 16'd14710, 16'd51847, 16'd29654, 16'd22200, 16'd47828});
	test_expansion(128'h314b360d12f056abf39bdf65aebcbae6, {16'd53889, 16'd51984, 16'd45774, 16'd46610, 16'd6513, 16'd23818, 16'd65372, 16'd40477, 16'd27055, 16'd48882, 16'd59308, 16'd40024, 16'd13361, 16'd11933, 16'd60038, 16'd37047, 16'd38433, 16'd33200, 16'd65324, 16'd56339, 16'd63465, 16'd26815, 16'd38914, 16'd8179, 16'd1547, 16'd54288});
	test_expansion(128'h65ceb7a3e294c5f510ac726580677e1c, {16'd9340, 16'd43370, 16'd13067, 16'd43869, 16'd22247, 16'd602, 16'd10734, 16'd18243, 16'd52333, 16'd44396, 16'd30683, 16'd45180, 16'd64090, 16'd29707, 16'd21904, 16'd60938, 16'd46251, 16'd40207, 16'd2256, 16'd28426, 16'd2196, 16'd42506, 16'd28365, 16'd18633, 16'd5491, 16'd55369});
	test_expansion(128'hd9542d247adb4194a83fe828ea899e55, {16'd18153, 16'd44864, 16'd40030, 16'd40901, 16'd17470, 16'd28541, 16'd2964, 16'd54440, 16'd45218, 16'd41445, 16'd16129, 16'd19601, 16'd11442, 16'd23597, 16'd20595, 16'd57955, 16'd17299, 16'd44686, 16'd5164, 16'd18435, 16'd57883, 16'd30377, 16'd12064, 16'd17591, 16'd53922, 16'd9862});
	test_expansion(128'h6600c6c21fc9aade4c31a6422230dd6a, {16'd41538, 16'd50238, 16'd6835, 16'd5502, 16'd52915, 16'd11882, 16'd40902, 16'd62727, 16'd47748, 16'd11396, 16'd35508, 16'd15289, 16'd17066, 16'd736, 16'd10433, 16'd723, 16'd12559, 16'd14515, 16'd51936, 16'd34078, 16'd54948, 16'd63233, 16'd17445, 16'd31561, 16'd54866, 16'd46549});
	test_expansion(128'hb12146e6a8ff1e1fd1e0f94555023db9, {16'd28004, 16'd14632, 16'd33438, 16'd23422, 16'd7905, 16'd48929, 16'd63976, 16'd33148, 16'd52651, 16'd12508, 16'd57431, 16'd22924, 16'd26007, 16'd39535, 16'd38501, 16'd42439, 16'd52956, 16'd53144, 16'd20089, 16'd25701, 16'd37144, 16'd23251, 16'd23094, 16'd9986, 16'd9286, 16'd30046});
	test_expansion(128'he70040e3b3fdba5ea0fe7d0d7a6cc170, {16'd47379, 16'd47027, 16'd22776, 16'd4638, 16'd12350, 16'd10536, 16'd65493, 16'd53008, 16'd19921, 16'd56123, 16'd1147, 16'd3071, 16'd51104, 16'd33482, 16'd9534, 16'd49372, 16'd28405, 16'd30034, 16'd40542, 16'd24607, 16'd26766, 16'd44175, 16'd14935, 16'd50090, 16'd43975, 16'd47956});
	test_expansion(128'hf70b7a71925eab9faf9fc3f73bdd46ea, {16'd62401, 16'd4547, 16'd53609, 16'd909, 16'd54844, 16'd29322, 16'd53677, 16'd63875, 16'd34241, 16'd6050, 16'd50208, 16'd21426, 16'd12265, 16'd60757, 16'd36073, 16'd50666, 16'd6994, 16'd41414, 16'd37073, 16'd51645, 16'd34276, 16'd39030, 16'd531, 16'd55427, 16'd43921, 16'd23317});
	test_expansion(128'h0cdf7b9f951b86d5ec6e11770cee69ff, {16'd13344, 16'd2505, 16'd32783, 16'd21267, 16'd60711, 16'd48955, 16'd43248, 16'd10268, 16'd60657, 16'd30639, 16'd30619, 16'd1273, 16'd27871, 16'd53289, 16'd23971, 16'd11480, 16'd62898, 16'd15095, 16'd10562, 16'd32918, 16'd23573, 16'd27488, 16'd41003, 16'd9641, 16'd8175, 16'd52727});
	test_expansion(128'h04c932f154386974fc49fdd377003cf2, {16'd27170, 16'd10678, 16'd11277, 16'd34639, 16'd63560, 16'd62718, 16'd59013, 16'd44420, 16'd33103, 16'd20197, 16'd47400, 16'd50030, 16'd18450, 16'd12926, 16'd16777, 16'd14910, 16'd43314, 16'd19066, 16'd64236, 16'd583, 16'd61972, 16'd28204, 16'd21217, 16'd40908, 16'd33922, 16'd24079});
	test_expansion(128'h5ba657d9d2bfd8f79be0a5fd461ce471, {16'd29922, 16'd53260, 16'd42518, 16'd37853, 16'd13161, 16'd63990, 16'd18365, 16'd48533, 16'd37760, 16'd9764, 16'd16496, 16'd50803, 16'd54957, 16'd19233, 16'd42388, 16'd20170, 16'd20554, 16'd16368, 16'd29404, 16'd18446, 16'd50452, 16'd16943, 16'd3650, 16'd18670, 16'd50242, 16'd42510});
	test_expansion(128'h8187c5793acab0625df592dff1a40e09, {16'd43063, 16'd62617, 16'd43036, 16'd26553, 16'd61899, 16'd19419, 16'd52639, 16'd4961, 16'd61460, 16'd26775, 16'd10809, 16'd19427, 16'd49941, 16'd11947, 16'd12401, 16'd10124, 16'd820, 16'd42082, 16'd9556, 16'd65173, 16'd3958, 16'd7955, 16'd8620, 16'd11172, 16'd37361, 16'd2024});
	test_expansion(128'h8119aaa4104d7e4feea189b2ca09b218, {16'd37850, 16'd50267, 16'd25330, 16'd9124, 16'd3946, 16'd24498, 16'd7355, 16'd54947, 16'd13560, 16'd26042, 16'd6805, 16'd34084, 16'd60471, 16'd12209, 16'd62318, 16'd61543, 16'd32654, 16'd59161, 16'd47755, 16'd39344, 16'd39991, 16'd52545, 16'd61985, 16'd17349, 16'd53632, 16'd14267});
	test_expansion(128'h689305f192ea8fa35fa0ff89e10b91f5, {16'd19499, 16'd63463, 16'd3083, 16'd54811, 16'd24876, 16'd61532, 16'd42508, 16'd10213, 16'd4070, 16'd56042, 16'd8012, 16'd24229, 16'd26176, 16'd27925, 16'd36074, 16'd40137, 16'd12504, 16'd10426, 16'd56226, 16'd60757, 16'd20609, 16'd38940, 16'd59142, 16'd17253, 16'd64824, 16'd31448});
	test_expansion(128'h2fc76a193445892ab9ac467bcef17162, {16'd63031, 16'd34447, 16'd60560, 16'd36863, 16'd45977, 16'd39965, 16'd50951, 16'd51575, 16'd53326, 16'd33924, 16'd31848, 16'd1555, 16'd63779, 16'd43877, 16'd65369, 16'd36703, 16'd59194, 16'd77, 16'd13330, 16'd35, 16'd47974, 16'd31410, 16'd64616, 16'd49059, 16'd51411, 16'd24051});
	test_expansion(128'hba3d355d4e906fef96d8cb53de6d1c5e, {16'd33479, 16'd10691, 16'd3575, 16'd42615, 16'd25819, 16'd13624, 16'd488, 16'd30740, 16'd33534, 16'd24762, 16'd42105, 16'd61414, 16'd57054, 16'd46860, 16'd1235, 16'd64752, 16'd9408, 16'd28686, 16'd38116, 16'd27902, 16'd20573, 16'd49804, 16'd49842, 16'd3454, 16'd65312, 16'd21839});
	test_expansion(128'h025d21a5184aaba6a5ce291989006770, {16'd21425, 16'd58541, 16'd62463, 16'd11025, 16'd64484, 16'd8921, 16'd28308, 16'd46511, 16'd44392, 16'd27525, 16'd57209, 16'd6599, 16'd48704, 16'd7620, 16'd29784, 16'd27456, 16'd28755, 16'd63407, 16'd3402, 16'd20755, 16'd44040, 16'd17615, 16'd45628, 16'd34913, 16'd42730, 16'd13659});
	test_expansion(128'ha27198efa37b610b94923f0fa6c472c4, {16'd8633, 16'd21948, 16'd59652, 16'd16471, 16'd50596, 16'd24742, 16'd2381, 16'd36625, 16'd51810, 16'd10285, 16'd62927, 16'd53929, 16'd20919, 16'd33835, 16'd40737, 16'd11142, 16'd17897, 16'd62592, 16'd59734, 16'd56336, 16'd6784, 16'd1609, 16'd43908, 16'd63233, 16'd64030, 16'd34265});
	test_expansion(128'h93721144c0c44e064538bbcbed23a7c9, {16'd53507, 16'd37993, 16'd40072, 16'd31241, 16'd17148, 16'd43840, 16'd41940, 16'd37370, 16'd56445, 16'd45049, 16'd25862, 16'd38010, 16'd19034, 16'd45717, 16'd38701, 16'd61580, 16'd45929, 16'd58489, 16'd12911, 16'd40698, 16'd55009, 16'd27616, 16'd44242, 16'd45810, 16'd45901, 16'd27039});
	test_expansion(128'h47f689b39bc969cf3a4553f4481a4ba1, {16'd18806, 16'd226, 16'd8892, 16'd47791, 16'd31475, 16'd61229, 16'd14652, 16'd4540, 16'd55840, 16'd33625, 16'd48663, 16'd30206, 16'd1346, 16'd30992, 16'd31621, 16'd57596, 16'd35079, 16'd25277, 16'd19915, 16'd38765, 16'd620, 16'd35198, 16'd12260, 16'd2330, 16'd17137, 16'd3965});
	test_expansion(128'hdc87b17fa4e9887450469400ffcca971, {16'd41112, 16'd15570, 16'd13182, 16'd11437, 16'd51701, 16'd33902, 16'd39791, 16'd51813, 16'd27604, 16'd61951, 16'd25239, 16'd37494, 16'd44318, 16'd17644, 16'd40047, 16'd4205, 16'd18967, 16'd44815, 16'd57405, 16'd43146, 16'd33868, 16'd2586, 16'd25874, 16'd52640, 16'd43857, 16'd17261});
	test_expansion(128'hf9f5ac4c35f598d89c71d690ad1eb860, {16'd63662, 16'd3058, 16'd37770, 16'd26258, 16'd9131, 16'd41722, 16'd3102, 16'd38953, 16'd9472, 16'd64376, 16'd44810, 16'd18544, 16'd16863, 16'd37130, 16'd29490, 16'd21536, 16'd6136, 16'd4387, 16'd42945, 16'd37825, 16'd24527, 16'd13697, 16'd42191, 16'd27768, 16'd5863, 16'd37500});
	test_expansion(128'hca5b6ddf9b87acea378bc5024853b64f, {16'd58314, 16'd60505, 16'd21778, 16'd62542, 16'd18560, 16'd58432, 16'd63998, 16'd29920, 16'd2409, 16'd24276, 16'd42119, 16'd35052, 16'd22721, 16'd28377, 16'd30697, 16'd4852, 16'd47035, 16'd38867, 16'd26006, 16'd46348, 16'd1870, 16'd53641, 16'd16331, 16'd49016, 16'd47670, 16'd21167});
	test_expansion(128'hb6f64b59be6122ccfff1f6f5dc8e2b9c, {16'd18028, 16'd34468, 16'd61901, 16'd52000, 16'd55111, 16'd46636, 16'd10654, 16'd51761, 16'd9693, 16'd19054, 16'd7623, 16'd34689, 16'd35221, 16'd62573, 16'd34271, 16'd1415, 16'd58961, 16'd25080, 16'd18535, 16'd51482, 16'd20020, 16'd9819, 16'd17362, 16'd25762, 16'd34001, 16'd46845});
	test_expansion(128'hc7c1e80c3faa4fa8dbbc0fe1f11c0f20, {16'd28275, 16'd152, 16'd52852, 16'd37621, 16'd38847, 16'd43393, 16'd63942, 16'd14302, 16'd55350, 16'd45107, 16'd13294, 16'd51198, 16'd56845, 16'd53800, 16'd54495, 16'd7875, 16'd11138, 16'd44418, 16'd18456, 16'd53125, 16'd30311, 16'd8826, 16'd7352, 16'd3100, 16'd45491, 16'd65194});
	test_expansion(128'ha03d2aa577f04aa65efb0200996404c6, {16'd39800, 16'd43695, 16'd28137, 16'd54603, 16'd23655, 16'd52683, 16'd56644, 16'd65208, 16'd18997, 16'd52739, 16'd44778, 16'd54555, 16'd61872, 16'd53825, 16'd52066, 16'd5188, 16'd34678, 16'd25190, 16'd5069, 16'd30486, 16'd8231, 16'd55979, 16'd51923, 16'd57543, 16'd18108, 16'd55642});
	test_expansion(128'h219f71fd96a8f3211edeb1cd4a546223, {16'd59078, 16'd60765, 16'd51016, 16'd42928, 16'd545, 16'd23875, 16'd37627, 16'd23164, 16'd50350, 16'd62342, 16'd2411, 16'd59912, 16'd14210, 16'd36142, 16'd7469, 16'd29608, 16'd54874, 16'd44200, 16'd28117, 16'd40293, 16'd52737, 16'd50801, 16'd42317, 16'd60053, 16'd24123, 16'd33621});
	test_expansion(128'hff10e77e1b40d2ab9db3aca433969f9c, {16'd60617, 16'd61891, 16'd10918, 16'd7754, 16'd18332, 16'd15661, 16'd64636, 16'd57018, 16'd23058, 16'd10003, 16'd51593, 16'd51258, 16'd40497, 16'd63846, 16'd52680, 16'd38399, 16'd50212, 16'd43541, 16'd22524, 16'd3026, 16'd33776, 16'd34661, 16'd15411, 16'd29405, 16'd49026, 16'd18832});
	test_expansion(128'h4035b3d17ffea873586a3151e6da635f, {16'd35811, 16'd60550, 16'd37909, 16'd32889, 16'd62268, 16'd29100, 16'd29912, 16'd46894, 16'd17479, 16'd6597, 16'd58513, 16'd18098, 16'd21533, 16'd42552, 16'd10391, 16'd44083, 16'd14098, 16'd41712, 16'd47890, 16'd6327, 16'd63603, 16'd48759, 16'd32166, 16'd56709, 16'd41939, 16'd14996});
	test_expansion(128'h53929a11e746e48cfe2c3f68cd797029, {16'd12731, 16'd34124, 16'd51946, 16'd27067, 16'd49713, 16'd56605, 16'd4208, 16'd24306, 16'd8629, 16'd40066, 16'd50623, 16'd16639, 16'd14716, 16'd15623, 16'd61213, 16'd41529, 16'd17431, 16'd9821, 16'd3701, 16'd5113, 16'd26508, 16'd38881, 16'd44585, 16'd44252, 16'd587, 16'd38784});
	test_expansion(128'h16b82c8678d985954850b6d3d8015368, {16'd65464, 16'd50956, 16'd1891, 16'd7366, 16'd10255, 16'd4390, 16'd36599, 16'd8810, 16'd31924, 16'd37713, 16'd43188, 16'd4598, 16'd53954, 16'd40655, 16'd55528, 16'd7948, 16'd32344, 16'd56289, 16'd30275, 16'd4571, 16'd15153, 16'd49419, 16'd40445, 16'd58217, 16'd2585, 16'd32121});
	test_expansion(128'hfa003f35672872f8b343ffeb521c9c3a, {16'd58667, 16'd3274, 16'd37061, 16'd53694, 16'd12257, 16'd9326, 16'd60729, 16'd64860, 16'd39185, 16'd37671, 16'd65269, 16'd21322, 16'd32725, 16'd18013, 16'd53158, 16'd2943, 16'd43321, 16'd55695, 16'd36609, 16'd27117, 16'd4278, 16'd17394, 16'd47914, 16'd36709, 16'd51683, 16'd29795});
	test_expansion(128'h6ec1cb4e8f2db3f41e249a2a62c4ade2, {16'd58681, 16'd54376, 16'd18148, 16'd38409, 16'd9218, 16'd59434, 16'd41676, 16'd55842, 16'd47392, 16'd19538, 16'd4036, 16'd56379, 16'd11609, 16'd29197, 16'd7854, 16'd49718, 16'd17892, 16'd34780, 16'd1458, 16'd27192, 16'd60724, 16'd10566, 16'd37554, 16'd18316, 16'd31350, 16'd31340});
	test_expansion(128'h7690cb677925287f103c1d86b40ad3d8, {16'd13464, 16'd64811, 16'd53594, 16'd5040, 16'd19563, 16'd47695, 16'd41777, 16'd62286, 16'd13735, 16'd12798, 16'd28781, 16'd8895, 16'd4442, 16'd14513, 16'd57186, 16'd27162, 16'd52215, 16'd37113, 16'd22393, 16'd39568, 16'd39165, 16'd11095, 16'd12169, 16'd29448, 16'd28127, 16'd22294});
	test_expansion(128'hd04fe0f4c4c95eb24c274b8fe0453d8b, {16'd34204, 16'd32436, 16'd43628, 16'd39141, 16'd31502, 16'd37266, 16'd14721, 16'd51746, 16'd46178, 16'd63042, 16'd52790, 16'd49074, 16'd35895, 16'd5086, 16'd25594, 16'd26948, 16'd29161, 16'd20380, 16'd31145, 16'd53176, 16'd19061, 16'd8959, 16'd21742, 16'd16264, 16'd53907, 16'd9839});
	test_expansion(128'hfe58dc628f6034c615f3fe9c8ffde81c, {16'd23962, 16'd36611, 16'd1947, 16'd64955, 16'd17853, 16'd12146, 16'd41398, 16'd54888, 16'd39763, 16'd16011, 16'd4356, 16'd10238, 16'd25295, 16'd8552, 16'd960, 16'd16496, 16'd22240, 16'd54222, 16'd60731, 16'd26675, 16'd19909, 16'd56467, 16'd63201, 16'd30773, 16'd11475, 16'd22354});
	test_expansion(128'hba6b3e7d4bc2840c96c4583c53668d52, {16'd30702, 16'd61295, 16'd17655, 16'd1284, 16'd57692, 16'd37659, 16'd40882, 16'd20940, 16'd53763, 16'd24551, 16'd50857, 16'd16362, 16'd36478, 16'd9204, 16'd43241, 16'd6643, 16'd56015, 16'd28759, 16'd64331, 16'd46395, 16'd5811, 16'd57226, 16'd41248, 16'd18300, 16'd26351, 16'd7185});
	test_expansion(128'haebe6ace9c79e1cb1c1a09c9b73ea511, {16'd60473, 16'd54099, 16'd13365, 16'd44649, 16'd56642, 16'd44856, 16'd12567, 16'd55225, 16'd39250, 16'd56604, 16'd34472, 16'd63799, 16'd10639, 16'd41170, 16'd53455, 16'd34861, 16'd50583, 16'd6484, 16'd31618, 16'd58757, 16'd5586, 16'd32660, 16'd15840, 16'd47891, 16'd49404, 16'd49051});
	test_expansion(128'h4b4e3bec1948a576e1e5be899d192c72, {16'd32883, 16'd28774, 16'd31192, 16'd49387, 16'd42444, 16'd51468, 16'd59860, 16'd3393, 16'd49475, 16'd30938, 16'd63845, 16'd12373, 16'd13883, 16'd50556, 16'd38631, 16'd53622, 16'd24757, 16'd47576, 16'd51390, 16'd18489, 16'd17438, 16'd25555, 16'd26541, 16'd43492, 16'd50096, 16'd11885});
	test_expansion(128'h050f8f6b9ab599991a2afacd68d30c8a, {16'd42845, 16'd33966, 16'd8208, 16'd41657, 16'd3407, 16'd2153, 16'd52350, 16'd62361, 16'd8305, 16'd64410, 16'd33597, 16'd18926, 16'd60952, 16'd36147, 16'd35583, 16'd1443, 16'd7947, 16'd48363, 16'd6449, 16'd40110, 16'd49009, 16'd61942, 16'd776, 16'd60404, 16'd52245, 16'd64033});
	test_expansion(128'h997fc62d8a0d2846208c75a9e21eca1f, {16'd38512, 16'd33362, 16'd30729, 16'd26627, 16'd64291, 16'd3475, 16'd38937, 16'd11939, 16'd26529, 16'd3532, 16'd40013, 16'd61023, 16'd6895, 16'd30496, 16'd24572, 16'd23697, 16'd62496, 16'd64255, 16'd64432, 16'd29170, 16'd6091, 16'd46059, 16'd19284, 16'd11457, 16'd10166, 16'd59850});
	test_expansion(128'h8b2c0788554529f23e051d1db4b4baf7, {16'd59609, 16'd29732, 16'd6737, 16'd57976, 16'd37042, 16'd64207, 16'd1778, 16'd17307, 16'd1587, 16'd56235, 16'd50384, 16'd15901, 16'd3268, 16'd13920, 16'd17598, 16'd10137, 16'd13553, 16'd60611, 16'd23937, 16'd59223, 16'd20007, 16'd1996, 16'd4370, 16'd60312, 16'd16566, 16'd6725});
	test_expansion(128'h2dbb2ffc95fbf0bc62333060161efb5a, {16'd44928, 16'd11469, 16'd2174, 16'd27178, 16'd43621, 16'd29186, 16'd211, 16'd17697, 16'd18745, 16'd5448, 16'd12446, 16'd1333, 16'd4484, 16'd65313, 16'd9261, 16'd61570, 16'd36371, 16'd18059, 16'd43704, 16'd30657, 16'd54935, 16'd61643, 16'd55761, 16'd29875, 16'd46033, 16'd56050});
	test_expansion(128'h4650f7c425b371cd7ed294932320ddb0, {16'd11491, 16'd4444, 16'd29075, 16'd19776, 16'd1305, 16'd40592, 16'd55261, 16'd6424, 16'd20827, 16'd50381, 16'd57755, 16'd18054, 16'd56999, 16'd13926, 16'd10396, 16'd23816, 16'd54415, 16'd51129, 16'd38191, 16'd32871, 16'd36748, 16'd33842, 16'd55351, 16'd47152, 16'd48836, 16'd25398});
	test_expansion(128'h2f96373b713096e6a757c6e3721575c5, {16'd53849, 16'd5294, 16'd6034, 16'd17337, 16'd20553, 16'd56645, 16'd30054, 16'd50619, 16'd1442, 16'd19797, 16'd15648, 16'd55630, 16'd21768, 16'd46435, 16'd52521, 16'd5350, 16'd8102, 16'd63833, 16'd38192, 16'd58836, 16'd13122, 16'd17179, 16'd3366, 16'd30220, 16'd64514, 16'd57598});
	test_expansion(128'ha738d1cce642951679f8db088f225746, {16'd9888, 16'd39040, 16'd723, 16'd52579, 16'd8832, 16'd17015, 16'd24079, 16'd22043, 16'd40834, 16'd12230, 16'd2125, 16'd28138, 16'd42923, 16'd2397, 16'd9717, 16'd14886, 16'd16000, 16'd2398, 16'd26015, 16'd45246, 16'd34962, 16'd2629, 16'd26100, 16'd4530, 16'd10833, 16'd34402});
	test_expansion(128'h025559d445aa74e6e1715d03027fbc9e, {16'd21044, 16'd22897, 16'd18577, 16'd25204, 16'd37607, 16'd29659, 16'd57151, 16'd61225, 16'd62352, 16'd5605, 16'd20614, 16'd50720, 16'd9416, 16'd25083, 16'd42525, 16'd28573, 16'd56924, 16'd20084, 16'd24067, 16'd46537, 16'd22858, 16'd38486, 16'd1270, 16'd4060, 16'd25210, 16'd38269});
	test_expansion(128'h3e2e5b845f9b92a1645b404c148656c0, {16'd25210, 16'd15002, 16'd54580, 16'd59001, 16'd22769, 16'd47740, 16'd13119, 16'd60312, 16'd29736, 16'd63594, 16'd33268, 16'd59685, 16'd30870, 16'd23470, 16'd64533, 16'd22075, 16'd26301, 16'd10412, 16'd53069, 16'd38223, 16'd13433, 16'd17459, 16'd61104, 16'd6647, 16'd34103, 16'd18524});
	test_expansion(128'h0ad3b49603e67ee42636515e41ee977a, {16'd31206, 16'd4603, 16'd5569, 16'd29183, 16'd36362, 16'd28984, 16'd44592, 16'd53221, 16'd7990, 16'd42724, 16'd35570, 16'd25582, 16'd32371, 16'd23161, 16'd31848, 16'd45901, 16'd40665, 16'd31761, 16'd18611, 16'd24037, 16'd49722, 16'd28844, 16'd18752, 16'd49029, 16'd13002, 16'd51837});
	test_expansion(128'h846ecaf178796a873199c1e58752a71f, {16'd24036, 16'd61227, 16'd56041, 16'd15851, 16'd12844, 16'd57786, 16'd36926, 16'd6085, 16'd20781, 16'd28528, 16'd38898, 16'd29663, 16'd15267, 16'd15552, 16'd41764, 16'd28946, 16'd12500, 16'd25233, 16'd18998, 16'd55044, 16'd50235, 16'd4682, 16'd17029, 16'd48443, 16'd53535, 16'd47207});
	test_expansion(128'h3fd92058291e052327616a0c59276d27, {16'd15748, 16'd60213, 16'd63866, 16'd3709, 16'd53313, 16'd47113, 16'd49583, 16'd16219, 16'd46911, 16'd21510, 16'd54253, 16'd28978, 16'd5422, 16'd20928, 16'd35567, 16'd3062, 16'd23922, 16'd22530, 16'd23521, 16'd23382, 16'd19930, 16'd41692, 16'd49071, 16'd34346, 16'd37001, 16'd37002});
	test_expansion(128'h74e3338bf844ad34e2549b4aec86dfb9, {16'd51924, 16'd27469, 16'd38149, 16'd7991, 16'd62634, 16'd56314, 16'd61306, 16'd13531, 16'd53943, 16'd5648, 16'd49855, 16'd40620, 16'd57411, 16'd56384, 16'd46527, 16'd64204, 16'd47454, 16'd13715, 16'd65351, 16'd46687, 16'd60008, 16'd53723, 16'd46553, 16'd1014, 16'd15259, 16'd53839});
	test_expansion(128'hc5f5cfede7422813e124204051e1656c, {16'd64531, 16'd30652, 16'd13954, 16'd64672, 16'd63203, 16'd41595, 16'd37166, 16'd17390, 16'd18300, 16'd33420, 16'd1371, 16'd13381, 16'd62008, 16'd61755, 16'd50979, 16'd19713, 16'd3746, 16'd64890, 16'd59643, 16'd28254, 16'd12742, 16'd14381, 16'd13437, 16'd46121, 16'd32644, 16'd56724});
	test_expansion(128'hbec0c2997e0f081f9d73a7f3bcb63c35, {16'd36628, 16'd51487, 16'd1930, 16'd3512, 16'd8934, 16'd55551, 16'd17402, 16'd39234, 16'd26647, 16'd47291, 16'd24312, 16'd16725, 16'd4843, 16'd5820, 16'd24955, 16'd4004, 16'd54619, 16'd8329, 16'd2498, 16'd18952, 16'd54428, 16'd59513, 16'd51664, 16'd48541, 16'd26796, 16'd40680});
	test_expansion(128'h1a2a1fb917cd1b56762123965a302a76, {16'd64469, 16'd24111, 16'd43118, 16'd29027, 16'd52723, 16'd58163, 16'd44093, 16'd59767, 16'd26434, 16'd41513, 16'd9021, 16'd65019, 16'd56227, 16'd47784, 16'd58578, 16'd38503, 16'd54721, 16'd2217, 16'd2618, 16'd59295, 16'd45891, 16'd34732, 16'd35350, 16'd2252, 16'd57037, 16'd9751});
	test_expansion(128'h736d9234689c592524db4a97f4b30c8d, {16'd20354, 16'd42485, 16'd47123, 16'd1934, 16'd32035, 16'd13739, 16'd56211, 16'd30192, 16'd1745, 16'd64490, 16'd45405, 16'd46627, 16'd32529, 16'd1836, 16'd57896, 16'd58760, 16'd1208, 16'd16798, 16'd48506, 16'd23900, 16'd13976, 16'd16534, 16'd13313, 16'd35254, 16'd9919, 16'd35849});
	test_expansion(128'h489797a0c2c50aed4202b9ccc935fe47, {16'd32306, 16'd58241, 16'd19191, 16'd64389, 16'd44955, 16'd939, 16'd42253, 16'd49939, 16'd1215, 16'd41734, 16'd7868, 16'd32817, 16'd5418, 16'd48240, 16'd4569, 16'd39067, 16'd27559, 16'd37446, 16'd61604, 16'd6961, 16'd28061, 16'd56109, 16'd38881, 16'd55313, 16'd9510, 16'd15557});
	test_expansion(128'hc5ace2fb2791f9d16cfcc52a54620de8, {16'd49893, 16'd36963, 16'd22593, 16'd34902, 16'd47360, 16'd40577, 16'd17679, 16'd24709, 16'd30237, 16'd56115, 16'd16103, 16'd58235, 16'd28091, 16'd40303, 16'd23015, 16'd9316, 16'd53478, 16'd61188, 16'd50907, 16'd40733, 16'd63426, 16'd38168, 16'd14087, 16'd62976, 16'd27271, 16'd13049});
	test_expansion(128'hb65369b1d0d46ce57fa201e4972779e7, {16'd58316, 16'd34261, 16'd4549, 16'd36610, 16'd56923, 16'd45201, 16'd17664, 16'd35894, 16'd26600, 16'd27143, 16'd21531, 16'd6866, 16'd4825, 16'd35549, 16'd38263, 16'd52897, 16'd59547, 16'd48748, 16'd28451, 16'd23108, 16'd59271, 16'd609, 16'd3712, 16'd15188, 16'd7110, 16'd6007});
	test_expansion(128'he755f163ef61c26f8ba50f6270d50cfb, {16'd9167, 16'd51358, 16'd27989, 16'd52913, 16'd15494, 16'd17058, 16'd5625, 16'd60676, 16'd50222, 16'd56048, 16'd61076, 16'd27164, 16'd12407, 16'd63149, 16'd11878, 16'd39992, 16'd38069, 16'd41025, 16'd20296, 16'd27012, 16'd65465, 16'd52023, 16'd47859, 16'd26132, 16'd18649, 16'd30011});
	test_expansion(128'h6eab3843ad42c56cfd8e7c1e2826b231, {16'd61107, 16'd19773, 16'd2257, 16'd20159, 16'd31488, 16'd5726, 16'd5315, 16'd35501, 16'd48769, 16'd44470, 16'd4765, 16'd39171, 16'd61504, 16'd19635, 16'd18412, 16'd63676, 16'd39912, 16'd47031, 16'd5764, 16'd23675, 16'd1515, 16'd32256, 16'd203, 16'd28790, 16'd12804, 16'd39341});
	test_expansion(128'h10b578970a30b546a06977251d32829e, {16'd15898, 16'd36556, 16'd12814, 16'd10883, 16'd2340, 16'd38843, 16'd56591, 16'd57951, 16'd2733, 16'd47271, 16'd2150, 16'd40958, 16'd49887, 16'd47053, 16'd42421, 16'd51843, 16'd1105, 16'd23000, 16'd6907, 16'd24681, 16'd45987, 16'd54437, 16'd23026, 16'd44573, 16'd17546, 16'd42297});
	test_expansion(128'h6e72df4a7affa9a4cd0bbdc8396cdf67, {16'd38005, 16'd33116, 16'd33597, 16'd51816, 16'd23790, 16'd40188, 16'd52798, 16'd52213, 16'd43342, 16'd57345, 16'd59555, 16'd19148, 16'd45141, 16'd41718, 16'd54623, 16'd17017, 16'd26126, 16'd57333, 16'd17525, 16'd20082, 16'd31086, 16'd13681, 16'd63132, 16'd13242, 16'd48029, 16'd29129});
	test_expansion(128'h05c45d0e64ff239366346895af2eaab4, {16'd10998, 16'd60491, 16'd25646, 16'd23971, 16'd48324, 16'd63838, 16'd9616, 16'd23658, 16'd57995, 16'd60580, 16'd11126, 16'd2821, 16'd44374, 16'd61047, 16'd65256, 16'd9165, 16'd54113, 16'd52083, 16'd28353, 16'd22952, 16'd37526, 16'd29512, 16'd59921, 16'd40528, 16'd65332, 16'd57127});
	test_expansion(128'h8f0f613084cd36b5dc3f5e34e4b23e06, {16'd49612, 16'd27908, 16'd39562, 16'd40035, 16'd1244, 16'd1307, 16'd1115, 16'd16722, 16'd43732, 16'd18784, 16'd12236, 16'd38993, 16'd60733, 16'd16563, 16'd36143, 16'd50580, 16'd41385, 16'd54194, 16'd26214, 16'd26392, 16'd63360, 16'd49343, 16'd5920, 16'd13386, 16'd20135, 16'd32070});
	test_expansion(128'heb2c27881bcaad760321493f9127dbda, {16'd11072, 16'd55347, 16'd39868, 16'd44630, 16'd32881, 16'd24059, 16'd40589, 16'd25491, 16'd24409, 16'd27559, 16'd9381, 16'd33604, 16'd65360, 16'd40267, 16'd24864, 16'd64471, 16'd23471, 16'd47009, 16'd9531, 16'd34000, 16'd49253, 16'd493, 16'd39538, 16'd25399, 16'd16898, 16'd16870});
	test_expansion(128'h8771ca94a8a49c8dd7d17533554da2c7, {16'd64250, 16'd27512, 16'd17565, 16'd47265, 16'd37505, 16'd21163, 16'd46510, 16'd56843, 16'd5536, 16'd44645, 16'd1789, 16'd43402, 16'd59638, 16'd6078, 16'd61029, 16'd60166, 16'd15930, 16'd31582, 16'd35156, 16'd19540, 16'd10895, 16'd50751, 16'd49886, 16'd18918, 16'd42921, 16'd43809});
	test_expansion(128'h692163791c1a5f9c1493e219b54f2047, {16'd34895, 16'd5177, 16'd9622, 16'd5746, 16'd32358, 16'd21243, 16'd46166, 16'd18717, 16'd55242, 16'd33588, 16'd13411, 16'd61889, 16'd22134, 16'd40954, 16'd17033, 16'd23934, 16'd49833, 16'd39810, 16'd6670, 16'd41295, 16'd5525, 16'd20932, 16'd28592, 16'd53670, 16'd42697, 16'd40736});
	test_expansion(128'h1b17b0c0b57343fbe85f6c3f5438a81b, {16'd19127, 16'd14411, 16'd24302, 16'd51899, 16'd50457, 16'd13878, 16'd40676, 16'd43221, 16'd46462, 16'd8002, 16'd40813, 16'd26687, 16'd50524, 16'd49074, 16'd64455, 16'd3419, 16'd16864, 16'd26244, 16'd23804, 16'd45700, 16'd27295, 16'd62285, 16'd43771, 16'd38313, 16'd5926, 16'd16518});
	test_expansion(128'hb3c7ea6fe17c6aab31420012b10bb81f, {16'd34067, 16'd56196, 16'd57273, 16'd40224, 16'd31302, 16'd20018, 16'd47189, 16'd40314, 16'd36691, 16'd31497, 16'd31469, 16'd35242, 16'd2955, 16'd46603, 16'd33615, 16'd9229, 16'd21612, 16'd43374, 16'd27649, 16'd38492, 16'd63351, 16'd21020, 16'd14961, 16'd36539, 16'd9566, 16'd39022});
	test_expansion(128'h17fc565ad6903c04d26228b3a50b7cb6, {16'd5290, 16'd38746, 16'd52803, 16'd61173, 16'd45982, 16'd49331, 16'd46438, 16'd57659, 16'd3063, 16'd58502, 16'd46592, 16'd34968, 16'd32265, 16'd4684, 16'd21586, 16'd31990, 16'd42854, 16'd38205, 16'd51366, 16'd61756, 16'd35813, 16'd17699, 16'd21208, 16'd54097, 16'd41770, 16'd52349});
	test_expansion(128'ha89d2ffaf51681f1b91a90632ec3a694, {16'd37473, 16'd16916, 16'd35640, 16'd49661, 16'd3685, 16'd10302, 16'd16919, 16'd55768, 16'd33649, 16'd35203, 16'd7389, 16'd28860, 16'd31783, 16'd10897, 16'd3100, 16'd62230, 16'd33021, 16'd31699, 16'd47480, 16'd22547, 16'd3798, 16'd2487, 16'd50662, 16'd4239, 16'd12606, 16'd11203});
	test_expansion(128'h17ee59316661195fb99a1ab646308e33, {16'd24500, 16'd25933, 16'd12768, 16'd24096, 16'd31853, 16'd40297, 16'd16142, 16'd53055, 16'd59084, 16'd12765, 16'd31136, 16'd26039, 16'd22461, 16'd58926, 16'd1018, 16'd51052, 16'd11664, 16'd65077, 16'd25528, 16'd15402, 16'd32999, 16'd15951, 16'd21702, 16'd18079, 16'd45436, 16'd28101});
	test_expansion(128'hf71282f108cdb74dd9260648486d3942, {16'd15644, 16'd64520, 16'd41796, 16'd46949, 16'd18713, 16'd43900, 16'd54662, 16'd18481, 16'd50860, 16'd34739, 16'd59606, 16'd51185, 16'd26481, 16'd3664, 16'd27517, 16'd42273, 16'd50792, 16'd30002, 16'd37670, 16'd30333, 16'd50454, 16'd52593, 16'd20003, 16'd13656, 16'd1895, 16'd21244});
	test_expansion(128'hd2d7ee46b88326d55082fca4aa72a1f9, {16'd56487, 16'd46763, 16'd14340, 16'd62955, 16'd58569, 16'd15807, 16'd52160, 16'd48376, 16'd52708, 16'd24959, 16'd37229, 16'd36974, 16'd196, 16'd57848, 16'd5428, 16'd64777, 16'd6528, 16'd32440, 16'd17429, 16'd24263, 16'd3346, 16'd15787, 16'd47239, 16'd35186, 16'd28933, 16'd59721});
	test_expansion(128'hb860176e0b2ded50dfe8c607b24fc94c, {16'd8419, 16'd33730, 16'd23482, 16'd7230, 16'd57436, 16'd16990, 16'd43208, 16'd50522, 16'd16997, 16'd6826, 16'd51921, 16'd23629, 16'd3023, 16'd36587, 16'd17224, 16'd51403, 16'd4708, 16'd33166, 16'd40244, 16'd56951, 16'd56130, 16'd37766, 16'd60336, 16'd35072, 16'd58059, 16'd1989});
	test_expansion(128'hb25b59ce0dcc3dd4b6d034c34c7f855c, {16'd43926, 16'd53989, 16'd23216, 16'd52957, 16'd25792, 16'd21657, 16'd45247, 16'd6839, 16'd6849, 16'd56775, 16'd34763, 16'd27766, 16'd38387, 16'd52245, 16'd17994, 16'd452, 16'd41740, 16'd3856, 16'd64464, 16'd16183, 16'd39220, 16'd41133, 16'd30925, 16'd8489, 16'd15437, 16'd30018});
	test_expansion(128'h04688c24417f2ac99d9d8a6414ecdf45, {16'd36306, 16'd31345, 16'd55716, 16'd10712, 16'd47758, 16'd26972, 16'd16004, 16'd15451, 16'd7846, 16'd57611, 16'd25542, 16'd18981, 16'd6504, 16'd57926, 16'd24255, 16'd42003, 16'd14742, 16'd3577, 16'd48495, 16'd23251, 16'd47822, 16'd1795, 16'd9094, 16'd36755, 16'd10535, 16'd22161});
	test_expansion(128'h7e499396bb91c1adb663483d82b1298a, {16'd52204, 16'd40381, 16'd4573, 16'd21743, 16'd58969, 16'd60429, 16'd51456, 16'd21548, 16'd32242, 16'd28290, 16'd60353, 16'd8995, 16'd62979, 16'd52109, 16'd61473, 16'd47621, 16'd31862, 16'd18348, 16'd32162, 16'd13250, 16'd39664, 16'd45904, 16'd12613, 16'd58551, 16'd27415, 16'd60126});
	test_expansion(128'h9947fe0b1cd87cb11d499f34909fd562, {16'd41774, 16'd1686, 16'd20960, 16'd374, 16'd64163, 16'd39884, 16'd4156, 16'd34735, 16'd39954, 16'd35966, 16'd11620, 16'd42638, 16'd24920, 16'd45002, 16'd2966, 16'd27503, 16'd32433, 16'd44395, 16'd19553, 16'd54294, 16'd10679, 16'd23293, 16'd45837, 16'd37164, 16'd20818, 16'd52522});
	test_expansion(128'h5e46e887ae54945e2d1b7d1869648fd6, {16'd55428, 16'd34032, 16'd20783, 16'd9371, 16'd3138, 16'd15266, 16'd24537, 16'd22018, 16'd33808, 16'd18392, 16'd60482, 16'd5855, 16'd53961, 16'd42394, 16'd4404, 16'd9373, 16'd18949, 16'd61778, 16'd57184, 16'd30531, 16'd45781, 16'd19521, 16'd17842, 16'd6444, 16'd12624, 16'd61192});
	test_expansion(128'h72d8b987bbf60f580649c568fd893868, {16'd5065, 16'd36693, 16'd45508, 16'd64876, 16'd57300, 16'd59383, 16'd18727, 16'd4956, 16'd43092, 16'd14525, 16'd37689, 16'd25185, 16'd37097, 16'd7637, 16'd43343, 16'd42152, 16'd9012, 16'd9158, 16'd46602, 16'd26710, 16'd3772, 16'd21572, 16'd25321, 16'd15837, 16'd45427, 16'd20471});
	test_expansion(128'h488dd0c7d6501f02aa611f46a1f586de, {16'd56545, 16'd4448, 16'd44625, 16'd8297, 16'd26896, 16'd5200, 16'd24044, 16'd30233, 16'd57361, 16'd63499, 16'd29276, 16'd12715, 16'd41419, 16'd36669, 16'd30075, 16'd22696, 16'd6614, 16'd15620, 16'd44985, 16'd51671, 16'd21511, 16'd61252, 16'd37590, 16'd62499, 16'd8271, 16'd7272});
	test_expansion(128'he4e4803743c5bbc063a837579c6cb615, {16'd64951, 16'd28754, 16'd26305, 16'd21785, 16'd25402, 16'd46927, 16'd37356, 16'd34744, 16'd23520, 16'd33743, 16'd4024, 16'd4097, 16'd7185, 16'd25744, 16'd2554, 16'd59381, 16'd3147, 16'd60709, 16'd2068, 16'd12738, 16'd45299, 16'd41089, 16'd16268, 16'd42525, 16'd38194, 16'd50450});
	test_expansion(128'h1a5d0aeb54d35183219e4b6183315699, {16'd4626, 16'd50323, 16'd34335, 16'd15510, 16'd6843, 16'd18495, 16'd60088, 16'd10695, 16'd16238, 16'd12712, 16'd18553, 16'd49276, 16'd23409, 16'd47259, 16'd25273, 16'd56124, 16'd63195, 16'd32025, 16'd54388, 16'd37834, 16'd49112, 16'd48944, 16'd42081, 16'd33587, 16'd14398, 16'd3081});
	test_expansion(128'h866c92337dda370a00698db229bddc85, {16'd25991, 16'd24498, 16'd44897, 16'd62925, 16'd23887, 16'd62144, 16'd39427, 16'd8184, 16'd36674, 16'd45167, 16'd32117, 16'd22485, 16'd9538, 16'd32786, 16'd30485, 16'd948, 16'd42764, 16'd24711, 16'd61582, 16'd42497, 16'd1846, 16'd5319, 16'd39688, 16'd48462, 16'd5753, 16'd44637});
	test_expansion(128'h31a46933eb26f07fa3dade0dcb4fd15d, {16'd2116, 16'd50179, 16'd37144, 16'd53468, 16'd21535, 16'd3936, 16'd874, 16'd51398, 16'd25476, 16'd36034, 16'd59406, 16'd23253, 16'd16746, 16'd8038, 16'd7828, 16'd45451, 16'd39052, 16'd18778, 16'd18784, 16'd57290, 16'd5506, 16'd49578, 16'd25132, 16'd33216, 16'd38769, 16'd10494});
	test_expansion(128'hb32a11df3c6a60698c78ed77727756bf, {16'd51551, 16'd53566, 16'd38369, 16'd44074, 16'd49017, 16'd63515, 16'd42860, 16'd29613, 16'd28397, 16'd35244, 16'd20208, 16'd17121, 16'd51832, 16'd60088, 16'd8711, 16'd50860, 16'd20220, 16'd30328, 16'd7085, 16'd37084, 16'd49593, 16'd52098, 16'd10804, 16'd35383, 16'd9788, 16'd39300});
	test_expansion(128'h639ee793a21eb680569628f061fba6cd, {16'd34681, 16'd12401, 16'd42141, 16'd22912, 16'd24364, 16'd13807, 16'd27776, 16'd61445, 16'd43934, 16'd17374, 16'd2930, 16'd59259, 16'd444, 16'd36335, 16'd44382, 16'd51608, 16'd57094, 16'd61077, 16'd1520, 16'd64177, 16'd44384, 16'd47352, 16'd49298, 16'd2440, 16'd47130, 16'd43929});
	test_expansion(128'hfc1bc35e555bcb7cc49ec635128be259, {16'd2109, 16'd51705, 16'd51656, 16'd44263, 16'd42463, 16'd58229, 16'd3216, 16'd30945, 16'd15712, 16'd11432, 16'd60905, 16'd40461, 16'd21456, 16'd37568, 16'd46613, 16'd9836, 16'd35226, 16'd58807, 16'd30404, 16'd48651, 16'd13853, 16'd29028, 16'd51499, 16'd6319, 16'd21303, 16'd37849});
	test_expansion(128'h7c7d3ebf645d6b3bceffec1588edd353, {16'd50609, 16'd54793, 16'd35050, 16'd55182, 16'd52000, 16'd56190, 16'd37235, 16'd28289, 16'd44521, 16'd22545, 16'd57049, 16'd41088, 16'd39302, 16'd32146, 16'd53161, 16'd62995, 16'd4648, 16'd30282, 16'd9882, 16'd58570, 16'd20443, 16'd7751, 16'd62905, 16'd20364, 16'd18221, 16'd56884});
	test_expansion(128'h23c77abb31e1601242201aacc52c507b, {16'd12293, 16'd13001, 16'd45004, 16'd41871, 16'd47577, 16'd14899, 16'd24711, 16'd40726, 16'd47502, 16'd32483, 16'd20814, 16'd37432, 16'd15510, 16'd45746, 16'd53604, 16'd10633, 16'd2639, 16'd25208, 16'd53574, 16'd52153, 16'd26953, 16'd28307, 16'd59815, 16'd25381, 16'd32255, 16'd8082});
	test_expansion(128'h9824ef0dadfcccc3162de1d5e3868ffe, {16'd65257, 16'd30712, 16'd15748, 16'd42180, 16'd2569, 16'd3538, 16'd24400, 16'd11085, 16'd43874, 16'd23993, 16'd20855, 16'd29218, 16'd48312, 16'd9965, 16'd48456, 16'd43007, 16'd28881, 16'd8475, 16'd10055, 16'd16361, 16'd7154, 16'd37773, 16'd8560, 16'd59156, 16'd28666, 16'd63020});
	test_expansion(128'hc15f072d3fac191a4d14e0db737af71a, {16'd32347, 16'd51794, 16'd20402, 16'd61714, 16'd53686, 16'd62160, 16'd36174, 16'd2412, 16'd44264, 16'd45986, 16'd49956, 16'd56101, 16'd44558, 16'd58714, 16'd63723, 16'd52273, 16'd57871, 16'd8041, 16'd18418, 16'd13583, 16'd45061, 16'd44815, 16'd56332, 16'd39392, 16'd48186, 16'd57646});
	test_expansion(128'h31e45a726f1ff69a3076e812e8556a34, {16'd13675, 16'd57108, 16'd29629, 16'd32901, 16'd32453, 16'd37869, 16'd34526, 16'd17796, 16'd33220, 16'd29183, 16'd7678, 16'd48567, 16'd28446, 16'd22316, 16'd59018, 16'd60911, 16'd42727, 16'd35266, 16'd4319, 16'd4308, 16'd19042, 16'd15734, 16'd43252, 16'd56703, 16'd47655, 16'd33315});
	test_expansion(128'h1dd79d4f57e22b42fff1494a785fdf61, {16'd6539, 16'd24370, 16'd60763, 16'd35859, 16'd11801, 16'd35875, 16'd43729, 16'd26134, 16'd54870, 16'd21520, 16'd34560, 16'd18575, 16'd3251, 16'd26139, 16'd52284, 16'd36861, 16'd63407, 16'd34848, 16'd44144, 16'd41522, 16'd10760, 16'd41983, 16'd51859, 16'd16720, 16'd5668, 16'd29045});
	test_expansion(128'h23d6aa0582580b675b44f24352583d26, {16'd13045, 16'd54376, 16'd40829, 16'd61208, 16'd55706, 16'd62785, 16'd56814, 16'd25271, 16'd48633, 16'd34265, 16'd38619, 16'd64342, 16'd33385, 16'd50871, 16'd6599, 16'd37478, 16'd13911, 16'd2657, 16'd45529, 16'd4522, 16'd59862, 16'd5137, 16'd4798, 16'd48468, 16'd40564, 16'd36228});
	test_expansion(128'hbcdb98183e9022e901fe64a7f0bcc425, {16'd22311, 16'd65489, 16'd44815, 16'd20832, 16'd39483, 16'd11834, 16'd26612, 16'd64118, 16'd48041, 16'd51930, 16'd63050, 16'd34906, 16'd7792, 16'd37813, 16'd6515, 16'd45297, 16'd61607, 16'd16987, 16'd48484, 16'd35882, 16'd13546, 16'd16387, 16'd26391, 16'd16903, 16'd48687, 16'd44601});
	test_expansion(128'h735ae8c5c3ecc54d08d6781ce866459d, {16'd58986, 16'd32460, 16'd11455, 16'd49088, 16'd1748, 16'd29158, 16'd6036, 16'd23389, 16'd19160, 16'd14351, 16'd35957, 16'd39402, 16'd9765, 16'd40386, 16'd64316, 16'd10012, 16'd56950, 16'd42167, 16'd7148, 16'd42960, 16'd13846, 16'd58608, 16'd57807, 16'd59705, 16'd59038, 16'd30284});
	test_expansion(128'h0cccc0b360cc07b0722ccdfd6e5dfb0c, {16'd4081, 16'd32682, 16'd46145, 16'd5598, 16'd45666, 16'd45785, 16'd31339, 16'd17921, 16'd55486, 16'd27546, 16'd30358, 16'd61150, 16'd1349, 16'd30673, 16'd34685, 16'd55476, 16'd2827, 16'd63505, 16'd2928, 16'd42604, 16'd34812, 16'd62886, 16'd32183, 16'd44320, 16'd3663, 16'd25164});
	test_expansion(128'h5c0ee02c7608d3249237631205c6dc0a, {16'd46182, 16'd6214, 16'd47801, 16'd11152, 16'd43977, 16'd3200, 16'd60997, 16'd42442, 16'd7945, 16'd11927, 16'd6424, 16'd48316, 16'd10417, 16'd22758, 16'd53719, 16'd34615, 16'd1490, 16'd14540, 16'd34402, 16'd1206, 16'd27102, 16'd2317, 16'd60714, 16'd33961, 16'd52336, 16'd27966});
	test_expansion(128'habbaef9ee4389a60eea2661afeec5d54, {16'd57597, 16'd5231, 16'd60991, 16'd53964, 16'd56997, 16'd42153, 16'd42374, 16'd46980, 16'd30817, 16'd39969, 16'd4277, 16'd43075, 16'd48098, 16'd4862, 16'd4089, 16'd27305, 16'd54921, 16'd29487, 16'd59769, 16'd60914, 16'd2390, 16'd41119, 16'd14608, 16'd56685, 16'd33267, 16'd28590});
	test_expansion(128'hf640eca9520a2431febd8bbb595850c6, {16'd46142, 16'd1559, 16'd48717, 16'd52990, 16'd53391, 16'd3159, 16'd53767, 16'd18554, 16'd38883, 16'd65399, 16'd30408, 16'd47851, 16'd11430, 16'd27844, 16'd1074, 16'd52639, 16'd648, 16'd57988, 16'd8798, 16'd52941, 16'd37106, 16'd56740, 16'd10383, 16'd57316, 16'd44003, 16'd6915});
	test_expansion(128'h49c54d0bd68c92bdc9f0f71971ac8903, {16'd58381, 16'd29475, 16'd53309, 16'd3324, 16'd12122, 16'd8887, 16'd53622, 16'd13918, 16'd34391, 16'd40130, 16'd39709, 16'd22171, 16'd60212, 16'd26053, 16'd58205, 16'd21697, 16'd40275, 16'd34292, 16'd14266, 16'd32275, 16'd1151, 16'd34961, 16'd21548, 16'd12487, 16'd8845, 16'd50797});
	test_expansion(128'hf59d72bbe7d94ad1d9a25a44887adcde, {16'd63476, 16'd32977, 16'd59414, 16'd42576, 16'd44560, 16'd8748, 16'd27209, 16'd47666, 16'd56128, 16'd47680, 16'd56246, 16'd1434, 16'd31753, 16'd11565, 16'd60038, 16'd39111, 16'd42934, 16'd24794, 16'd10646, 16'd39367, 16'd64431, 16'd52859, 16'd29811, 16'd31705, 16'd46916, 16'd8726});
	test_expansion(128'h847bacc8a0980672c6178ee09d95e0d8, {16'd62762, 16'd35599, 16'd64296, 16'd54618, 16'd38598, 16'd64836, 16'd30170, 16'd32797, 16'd44548, 16'd27731, 16'd60926, 16'd56379, 16'd43106, 16'd5321, 16'd65245, 16'd52922, 16'd61581, 16'd29131, 16'd27072, 16'd25892, 16'd11449, 16'd58679, 16'd19426, 16'd26580, 16'd20278, 16'd8530});
	test_expansion(128'h30285991afb57e00b489af7d2d946f7a, {16'd11159, 16'd52309, 16'd62177, 16'd65261, 16'd22632, 16'd21366, 16'd10224, 16'd22907, 16'd48297, 16'd53144, 16'd46900, 16'd63148, 16'd20156, 16'd49363, 16'd53334, 16'd49709, 16'd39749, 16'd10695, 16'd1155, 16'd60340, 16'd56637, 16'd35211, 16'd23269, 16'd2475, 16'd36494, 16'd21006});
	test_expansion(128'h8bc82add88e4a3009e84df2c01bb4298, {16'd46840, 16'd37717, 16'd12119, 16'd39297, 16'd58055, 16'd48398, 16'd60412, 16'd32300, 16'd32221, 16'd25700, 16'd33867, 16'd63512, 16'd52218, 16'd49748, 16'd41324, 16'd40243, 16'd43434, 16'd50089, 16'd17939, 16'd2355, 16'd45064, 16'd2065, 16'd40216, 16'd18782, 16'd36070, 16'd64430});
	test_expansion(128'he871754de2e90ccf2d4b524c7a93a4ea, {16'd64696, 16'd26036, 16'd29263, 16'd14632, 16'd53119, 16'd18778, 16'd35052, 16'd58980, 16'd43962, 16'd14252, 16'd49511, 16'd22167, 16'd56908, 16'd65002, 16'd20346, 16'd6075, 16'd40399, 16'd22087, 16'd93, 16'd25587, 16'd59025, 16'd39861, 16'd92, 16'd39210, 16'd3444, 16'd25265});
	test_expansion(128'h96fdb3abb3e76db2c9633ba2a456f110, {16'd32491, 16'd43685, 16'd49010, 16'd28324, 16'd17497, 16'd18495, 16'd17900, 16'd54187, 16'd43714, 16'd59756, 16'd41599, 16'd47506, 16'd42587, 16'd56312, 16'd29622, 16'd28316, 16'd39921, 16'd43592, 16'd49366, 16'd39825, 16'd34833, 16'd9073, 16'd60933, 16'd19988, 16'd46152, 16'd43306});
	test_expansion(128'hd737329dd505a82125ee3be2c683a872, {16'd7571, 16'd21872, 16'd62110, 16'd28028, 16'd27343, 16'd58026, 16'd14066, 16'd19951, 16'd7049, 16'd18060, 16'd9835, 16'd45607, 16'd12439, 16'd15219, 16'd56343, 16'd30779, 16'd5095, 16'd50057, 16'd57625, 16'd33631, 16'd18478, 16'd43389, 16'd8094, 16'd38719, 16'd36907, 16'd34128});
	test_expansion(128'hd82e0b68ba3d2607d71a30944335d3f9, {16'd39749, 16'd10021, 16'd20616, 16'd1833, 16'd56903, 16'd55305, 16'd31419, 16'd20383, 16'd958, 16'd12690, 16'd59288, 16'd10989, 16'd42077, 16'd47802, 16'd22454, 16'd16490, 16'd19931, 16'd2266, 16'd3585, 16'd12257, 16'd11238, 16'd2086, 16'd7090, 16'd57048, 16'd24684, 16'd47442});
	test_expansion(128'hc97fc24ab95ebe73de03c0b58c86bbab, {16'd62891, 16'd28932, 16'd55316, 16'd12566, 16'd42940, 16'd28328, 16'd26072, 16'd48921, 16'd3447, 16'd916, 16'd12598, 16'd9873, 16'd16301, 16'd1158, 16'd23906, 16'd5627, 16'd64531, 16'd26862, 16'd53651, 16'd52556, 16'd56174, 16'd46415, 16'd5390, 16'd30324, 16'd11109, 16'd24466});
	test_expansion(128'h21d99167bb156ee4ff0f925cea999629, {16'd10321, 16'd51301, 16'd44508, 16'd28690, 16'd5507, 16'd7796, 16'd54684, 16'd2707, 16'd60337, 16'd60196, 16'd36817, 16'd34183, 16'd3607, 16'd22541, 16'd205, 16'd52325, 16'd64785, 16'd61246, 16'd7990, 16'd47014, 16'd37041, 16'd36266, 16'd32939, 16'd64255, 16'd36214, 16'd17626});
	test_expansion(128'hdede6a4e45ada6fe34e17b279cf5d175, {16'd25844, 16'd2998, 16'd35395, 16'd38685, 16'd5294, 16'd38077, 16'd35919, 16'd24959, 16'd26859, 16'd46473, 16'd1467, 16'd39294, 16'd57608, 16'd20231, 16'd2269, 16'd33684, 16'd63364, 16'd46306, 16'd2823, 16'd58188, 16'd23552, 16'd16369, 16'd17066, 16'd58055, 16'd64567, 16'd16634});
	test_expansion(128'h57be9410bc18b2a3755b3ff97be056c4, {16'd36148, 16'd27982, 16'd32176, 16'd40233, 16'd57233, 16'd13521, 16'd48695, 16'd60704, 16'd20279, 16'd35006, 16'd62527, 16'd6197, 16'd9859, 16'd53801, 16'd12872, 16'd36892, 16'd573, 16'd54540, 16'd56757, 16'd55542, 16'd23877, 16'd34905, 16'd20405, 16'd61476, 16'd63991, 16'd7267});
	test_expansion(128'he9e9e653045b58b2349d60d9fcf2325d, {16'd58381, 16'd4108, 16'd30324, 16'd35408, 16'd51917, 16'd42133, 16'd51966, 16'd23221, 16'd38400, 16'd9356, 16'd64801, 16'd38537, 16'd50176, 16'd45232, 16'd11037, 16'd25117, 16'd45119, 16'd56682, 16'd14802, 16'd33271, 16'd21308, 16'd47521, 16'd54808, 16'd35443, 16'd37283, 16'd12452});
	test_expansion(128'h018492678845fe38da9d9043bd3c801a, {16'd54704, 16'd540, 16'd50738, 16'd21487, 16'd26945, 16'd18760, 16'd20508, 16'd49645, 16'd22470, 16'd16559, 16'd41721, 16'd41290, 16'd1759, 16'd41098, 16'd27595, 16'd6888, 16'd30150, 16'd29617, 16'd58507, 16'd65132, 16'd48783, 16'd43745, 16'd46421, 16'd32424, 16'd32933, 16'd7540});
	test_expansion(128'h02e683a46e6b3397aec3e325bff170c5, {16'd47084, 16'd63667, 16'd31996, 16'd28105, 16'd12232, 16'd6408, 16'd9420, 16'd29159, 16'd7218, 16'd29735, 16'd22206, 16'd60105, 16'd39309, 16'd57468, 16'd26015, 16'd86, 16'd33447, 16'd22518, 16'd37840, 16'd41600, 16'd13180, 16'd55438, 16'd57990, 16'd33289, 16'd38515, 16'd31004});
	test_expansion(128'hfe0c694039f756ffe6290b5aa25ec89d, {16'd35462, 16'd59499, 16'd30204, 16'd55481, 16'd14637, 16'd3739, 16'd11686, 16'd29771, 16'd53405, 16'd9931, 16'd44000, 16'd22680, 16'd47522, 16'd62884, 16'd5503, 16'd496, 16'd7536, 16'd44320, 16'd46679, 16'd57396, 16'd21070, 16'd63760, 16'd39674, 16'd42955, 16'd6314, 16'd63393});
	test_expansion(128'h15f3ff70944bb13829bd4f92151da323, {16'd63790, 16'd14401, 16'd3993, 16'd44915, 16'd55440, 16'd5959, 16'd11355, 16'd24507, 16'd3356, 16'd55485, 16'd41366, 16'd3620, 16'd19473, 16'd38430, 16'd30955, 16'd28122, 16'd64345, 16'd47918, 16'd31053, 16'd49087, 16'd51784, 16'd59404, 16'd3265, 16'd4894, 16'd12796, 16'd65496});
	test_expansion(128'h87b8b5c867753f8942fbc355b7251c24, {16'd22321, 16'd28717, 16'd16206, 16'd53238, 16'd13626, 16'd41667, 16'd36358, 16'd58228, 16'd27133, 16'd28877, 16'd27085, 16'd27552, 16'd59594, 16'd26326, 16'd44961, 16'd31432, 16'd12505, 16'd47860, 16'd21523, 16'd48268, 16'd36150, 16'd16384, 16'd15729, 16'd17982, 16'd38670, 16'd28033});
	test_expansion(128'h054b27f7d744234ee9a27d06658ed778, {16'd54495, 16'd9560, 16'd23972, 16'd7159, 16'd61071, 16'd63995, 16'd36564, 16'd50208, 16'd3867, 16'd21002, 16'd20675, 16'd12536, 16'd57446, 16'd5266, 16'd17726, 16'd46422, 16'd18275, 16'd60318, 16'd53599, 16'd14821, 16'd3980, 16'd61892, 16'd64693, 16'd31652, 16'd35100, 16'd65245});
	test_expansion(128'he11269c73179cb1b7b34a57a25e3f0eb, {16'd37856, 16'd25567, 16'd22681, 16'd10663, 16'd30783, 16'd19157, 16'd24909, 16'd57975, 16'd10684, 16'd58396, 16'd12631, 16'd37447, 16'd52891, 16'd59695, 16'd2041, 16'd5731, 16'd25633, 16'd46613, 16'd39203, 16'd52795, 16'd48546, 16'd28856, 16'd38759, 16'd61444, 16'd27855, 16'd32655});
	test_expansion(128'hd3da7384b50ad9bc02d36611e248e2ea, {16'd5362, 16'd3035, 16'd38824, 16'd54341, 16'd60848, 16'd56685, 16'd58244, 16'd4966, 16'd27319, 16'd13537, 16'd63706, 16'd42727, 16'd61294, 16'd46780, 16'd5386, 16'd27949, 16'd48387, 16'd7218, 16'd5196, 16'd45636, 16'd56899, 16'd38041, 16'd1220, 16'd15642, 16'd6584, 16'd64066});
	test_expansion(128'h3fd7a4477ef692c31c9f7118b884eb07, {16'd62858, 16'd23794, 16'd37399, 16'd27341, 16'd50197, 16'd65507, 16'd8178, 16'd63411, 16'd14506, 16'd56923, 16'd39147, 16'd4675, 16'd63823, 16'd3300, 16'd27033, 16'd29432, 16'd36234, 16'd43452, 16'd23993, 16'd59112, 16'd10917, 16'd52282, 16'd13892, 16'd43206, 16'd57471, 16'd64490});
	test_expansion(128'ha3dfc2cbb525743cdc3dd7d4d56ef030, {16'd141, 16'd50811, 16'd24140, 16'd60773, 16'd253, 16'd1746, 16'd45210, 16'd45053, 16'd26534, 16'd52806, 16'd13359, 16'd35896, 16'd14185, 16'd37757, 16'd3274, 16'd10276, 16'd5135, 16'd48431, 16'd9420, 16'd37767, 16'd49654, 16'd65265, 16'd38199, 16'd25201, 16'd21699, 16'd1924});
	test_expansion(128'h8e9c64cf681ef96ee3a2e693487412dd, {16'd39931, 16'd13259, 16'd45771, 16'd1656, 16'd32304, 16'd45685, 16'd51275, 16'd14913, 16'd55938, 16'd50068, 16'd26440, 16'd31500, 16'd15469, 16'd13321, 16'd61716, 16'd30376, 16'd57328, 16'd56210, 16'd48821, 16'd36359, 16'd18506, 16'd61434, 16'd29402, 16'd49181, 16'd21118, 16'd26007});
	test_expansion(128'hae54e389927d8040f190fc1ec6e225fb, {16'd22500, 16'd10312, 16'd34010, 16'd55370, 16'd7235, 16'd19641, 16'd33147, 16'd14407, 16'd15614, 16'd48282, 16'd61865, 16'd40643, 16'd1493, 16'd7512, 16'd1932, 16'd29219, 16'd63275, 16'd58016, 16'd623, 16'd51775, 16'd25048, 16'd55315, 16'd29853, 16'd59191, 16'd63956, 16'd55862});
	test_expansion(128'h35067d6f9043ff609ecbfa0534dc05dd, {16'd19466, 16'd17406, 16'd17583, 16'd34135, 16'd21679, 16'd22514, 16'd43175, 16'd5612, 16'd27236, 16'd33752, 16'd52698, 16'd51827, 16'd23368, 16'd35878, 16'd49642, 16'd19378, 16'd20670, 16'd5937, 16'd30137, 16'd38173, 16'd61514, 16'd63635, 16'd56748, 16'd2086, 16'd42739, 16'd35343});
	test_expansion(128'h1a9df4f31f9d557d333a7c28f7bbbe63, {16'd33220, 16'd36838, 16'd37996, 16'd39673, 16'd14969, 16'd2786, 16'd64478, 16'd47590, 16'd49329, 16'd6493, 16'd9004, 16'd28295, 16'd59489, 16'd17134, 16'd32782, 16'd6100, 16'd7442, 16'd46314, 16'd46335, 16'd7772, 16'd50237, 16'd29266, 16'd32796, 16'd19069, 16'd7841, 16'd53726});
	test_expansion(128'h887de5841cad4fb15ef1ced026005e05, {16'd58369, 16'd9015, 16'd13439, 16'd59313, 16'd54577, 16'd53697, 16'd42651, 16'd40331, 16'd24657, 16'd10307, 16'd53463, 16'd48130, 16'd65357, 16'd60597, 16'd22624, 16'd5370, 16'd19358, 16'd24005, 16'd56171, 16'd26384, 16'd21423, 16'd29228, 16'd29054, 16'd31879, 16'd13807, 16'd38074});
	test_expansion(128'h5b73929da3f1908ab16e1fff56dd9c5e, {16'd38364, 16'd35055, 16'd4954, 16'd50609, 16'd25989, 16'd27229, 16'd18564, 16'd58794, 16'd60713, 16'd50852, 16'd21126, 16'd60572, 16'd29095, 16'd53620, 16'd25821, 16'd45821, 16'd58272, 16'd24422, 16'd41525, 16'd50768, 16'd20097, 16'd45368, 16'd62654, 16'd56717, 16'd35997, 16'd49238});
	test_expansion(128'hbe136acd691e81daf15a1a80d2a35622, {16'd20009, 16'd19701, 16'd34325, 16'd31316, 16'd33211, 16'd33900, 16'd63868, 16'd32295, 16'd12959, 16'd21273, 16'd3237, 16'd17172, 16'd23287, 16'd20009, 16'd8802, 16'd64236, 16'd32794, 16'd47470, 16'd57034, 16'd6406, 16'd27937, 16'd37188, 16'd19018, 16'd46573, 16'd35356, 16'd27102});
	test_expansion(128'he7ff9ee8b2af0b3e0e54a660c5e0e421, {16'd2046, 16'd58219, 16'd8689, 16'd12279, 16'd22441, 16'd15650, 16'd29151, 16'd33839, 16'd13266, 16'd33117, 16'd29347, 16'd46600, 16'd48061, 16'd17068, 16'd27021, 16'd880, 16'd1159, 16'd19288, 16'd59201, 16'd56908, 16'd9987, 16'd49888, 16'd16386, 16'd49258, 16'd38589, 16'd48931});
	test_expansion(128'hd2135b1f20a4cb23c7bb69cf19df5e8b, {16'd37621, 16'd22905, 16'd40980, 16'd29527, 16'd64665, 16'd16577, 16'd32180, 16'd50343, 16'd31909, 16'd14390, 16'd31356, 16'd35612, 16'd34445, 16'd20495, 16'd3352, 16'd8300, 16'd31993, 16'd2125, 16'd40211, 16'd38398, 16'd18880, 16'd32574, 16'd32914, 16'd52214, 16'd579, 16'd3589});
	test_expansion(128'haf94fe07c068e91743e25d85c7031aca, {16'd12183, 16'd40188, 16'd38764, 16'd24280, 16'd29902, 16'd42326, 16'd31586, 16'd14173, 16'd42689, 16'd1342, 16'd47342, 16'd19991, 16'd37546, 16'd14129, 16'd59454, 16'd58484, 16'd26151, 16'd32680, 16'd47092, 16'd44563, 16'd34815, 16'd34311, 16'd38399, 16'd333, 16'd45685, 16'd27473});
	test_expansion(128'h6396fd839a3c16d849b144bfecc8d24f, {16'd33411, 16'd38801, 16'd65431, 16'd43051, 16'd48985, 16'd64311, 16'd3384, 16'd51197, 16'd43445, 16'd25576, 16'd19375, 16'd49680, 16'd47691, 16'd47056, 16'd35114, 16'd17763, 16'd45920, 16'd39164, 16'd26535, 16'd42406, 16'd60520, 16'd35785, 16'd58092, 16'd59830, 16'd7910, 16'd44690});
	test_expansion(128'h8f23934dc9d1bd424b3f74b5f7ab506c, {16'd3861, 16'd62679, 16'd9342, 16'd15564, 16'd65517, 16'd27111, 16'd28939, 16'd48764, 16'd58237, 16'd914, 16'd11300, 16'd26495, 16'd29309, 16'd29365, 16'd4184, 16'd63362, 16'd5471, 16'd36383, 16'd28860, 16'd34686, 16'd17427, 16'd50980, 16'd50763, 16'd47319, 16'd22418, 16'd13278});
	test_expansion(128'he0c2e5174d0d71087f219a5560b09747, {16'd46333, 16'd41305, 16'd26938, 16'd16010, 16'd53145, 16'd52532, 16'd62456, 16'd35608, 16'd22371, 16'd38949, 16'd14030, 16'd40394, 16'd56134, 16'd1411, 16'd44455, 16'd8476, 16'd39902, 16'd7803, 16'd51294, 16'd31826, 16'd51069, 16'd36748, 16'd8455, 16'd5391, 16'd62303, 16'd1383});
	test_expansion(128'h8b64b4985b8072d965c93bc031c937bb, {16'd59284, 16'd16945, 16'd10880, 16'd380, 16'd48146, 16'd10459, 16'd22555, 16'd13426, 16'd64060, 16'd54277, 16'd9403, 16'd595, 16'd10068, 16'd43697, 16'd61154, 16'd59382, 16'd4720, 16'd51247, 16'd56963, 16'd22979, 16'd48275, 16'd58449, 16'd16877, 16'd9018, 16'd9346, 16'd61446});
	test_expansion(128'hfdd47c924a376a62960bf4006650afaf, {16'd24704, 16'd62064, 16'd15627, 16'd26678, 16'd23570, 16'd5973, 16'd65047, 16'd59665, 16'd37945, 16'd7440, 16'd53897, 16'd11243, 16'd55115, 16'd62962, 16'd35267, 16'd56198, 16'd44862, 16'd4570, 16'd57740, 16'd24701, 16'd34276, 16'd63359, 16'd18267, 16'd30852, 16'd61175, 16'd22656});
	test_expansion(128'h80ab031248f2516351148c33afd5108d, {16'd26741, 16'd42577, 16'd47388, 16'd44837, 16'd48187, 16'd27400, 16'd37082, 16'd32282, 16'd64021, 16'd1129, 16'd12205, 16'd58596, 16'd35284, 16'd27488, 16'd43652, 16'd55142, 16'd59712, 16'd15048, 16'd37808, 16'd18601, 16'd19235, 16'd33474, 16'd18588, 16'd36006, 16'd52903, 16'd14216});
	test_expansion(128'hb610646f1b0b18dae6d5127fc54ecbd7, {16'd42461, 16'd34350, 16'd50234, 16'd13440, 16'd8303, 16'd22804, 16'd31331, 16'd19062, 16'd34781, 16'd59839, 16'd42073, 16'd5498, 16'd37237, 16'd62150, 16'd24830, 16'd21463, 16'd54568, 16'd20323, 16'd34855, 16'd55248, 16'd48476, 16'd60610, 16'd14442, 16'd8224, 16'd31199, 16'd42564});
	test_expansion(128'hce6ec733cd22581672df1ac2689b35d2, {16'd6657, 16'd10396, 16'd46675, 16'd15623, 16'd11440, 16'd24917, 16'd10455, 16'd61780, 16'd58146, 16'd58870, 16'd11259, 16'd60372, 16'd656, 16'd64158, 16'd63080, 16'd17243, 16'd19127, 16'd16131, 16'd57150, 16'd50352, 16'd4711, 16'd60328, 16'd51290, 16'd56661, 16'd57953, 16'd20668});
	test_expansion(128'hc4c8fd0b86ecd52f2112b83dc7436d0b, {16'd19425, 16'd56722, 16'd7246, 16'd29911, 16'd2880, 16'd422, 16'd50221, 16'd64976, 16'd60679, 16'd45796, 16'd10710, 16'd56107, 16'd24281, 16'd6613, 16'd35858, 16'd19605, 16'd12083, 16'd7819, 16'd52701, 16'd27088, 16'd35131, 16'd45511, 16'd25680, 16'd16651, 16'd58792, 16'd64000});
	test_expansion(128'h0823a7db6e58c828d2c3456139af9917, {16'd29783, 16'd48387, 16'd33972, 16'd57896, 16'd44083, 16'd38879, 16'd41672, 16'd49334, 16'd25739, 16'd47550, 16'd3026, 16'd49074, 16'd18419, 16'd47429, 16'd8101, 16'd525, 16'd16403, 16'd54626, 16'd47532, 16'd63404, 16'd47529, 16'd16545, 16'd2287, 16'd15679, 16'd62866, 16'd3246});
	test_expansion(128'h83afbff49ae75b22b6fe72376803dc06, {16'd60169, 16'd34258, 16'd58179, 16'd20675, 16'd47058, 16'd29969, 16'd4645, 16'd12230, 16'd5821, 16'd65110, 16'd29279, 16'd19506, 16'd56736, 16'd6704, 16'd22257, 16'd54722, 16'd38266, 16'd3980, 16'd55995, 16'd48660, 16'd14941, 16'd2161, 16'd34435, 16'd16173, 16'd18940, 16'd51288});
	test_expansion(128'he0fe3a0a273a5a87d281b79cf74f25fd, {16'd11362, 16'd65467, 16'd57681, 16'd61425, 16'd59498, 16'd5753, 16'd44499, 16'd15649, 16'd122, 16'd50711, 16'd28553, 16'd59399, 16'd11376, 16'd15860, 16'd24209, 16'd56909, 16'd51664, 16'd48400, 16'd16124, 16'd35005, 16'd40361, 16'd3440, 16'd60497, 16'd37932, 16'd24145, 16'd25002});
	test_expansion(128'h9121e9f6596d5bec957be939e4ea7383, {16'd9146, 16'd51102, 16'd33129, 16'd6886, 16'd34958, 16'd13674, 16'd64693, 16'd21210, 16'd52592, 16'd49749, 16'd24970, 16'd44647, 16'd31256, 16'd48901, 16'd34132, 16'd64395, 16'd46878, 16'd51382, 16'd19834, 16'd3815, 16'd5644, 16'd10122, 16'd20983, 16'd53495, 16'd33940, 16'd25080});
	test_expansion(128'ha965872b953fa9ad1ad99aee664631d8, {16'd51607, 16'd2605, 16'd26079, 16'd25221, 16'd49190, 16'd13277, 16'd55335, 16'd7407, 16'd35950, 16'd56130, 16'd50812, 16'd55925, 16'd64707, 16'd33039, 16'd56598, 16'd17242, 16'd6060, 16'd44201, 16'd8727, 16'd32775, 16'd20313, 16'd64700, 16'd5322, 16'd16531, 16'd17918, 16'd42106});
	test_expansion(128'h31bea79a313c77e04e5803e5a8d37810, {16'd65066, 16'd18573, 16'd210, 16'd50687, 16'd63943, 16'd49278, 16'd51357, 16'd16860, 16'd29793, 16'd11359, 16'd22111, 16'd43297, 16'd50230, 16'd55943, 16'd46392, 16'd16621, 16'd12382, 16'd34453, 16'd37535, 16'd37968, 16'd58689, 16'd3939, 16'd32115, 16'd21161, 16'd12924, 16'd64285});
	test_expansion(128'hb93e0c3d7e83b3df159fbb8cfe3ccd07, {16'd42084, 16'd25589, 16'd59108, 16'd38279, 16'd41613, 16'd54514, 16'd5825, 16'd41967, 16'd54382, 16'd50030, 16'd64395, 16'd37814, 16'd23459, 16'd39167, 16'd43300, 16'd28961, 16'd44920, 16'd37328, 16'd37966, 16'd43162, 16'd8713, 16'd8929, 16'd47484, 16'd20967, 16'd57908, 16'd32922});
	test_expansion(128'h9862f76073f37d09e06ea04e45b674c8, {16'd49825, 16'd14589, 16'd18367, 16'd42967, 16'd57328, 16'd36967, 16'd25068, 16'd7172, 16'd1905, 16'd16301, 16'd5373, 16'd25626, 16'd20616, 16'd3104, 16'd14338, 16'd14091, 16'd44668, 16'd23270, 16'd35505, 16'd3537, 16'd41736, 16'd32588, 16'd39657, 16'd41496, 16'd31872, 16'd25203});
	test_expansion(128'h4e89b1f3fd9574069a7a315740040f1f, {16'd1693, 16'd16525, 16'd14577, 16'd56829, 16'd29141, 16'd48394, 16'd34688, 16'd24699, 16'd12052, 16'd55828, 16'd34980, 16'd57931, 16'd55428, 16'd8259, 16'd32771, 16'd18213, 16'd51544, 16'd44661, 16'd56270, 16'd16152, 16'd10802, 16'd62005, 16'd45901, 16'd62433, 16'd26188, 16'd6994});
	test_expansion(128'h93fd363747553a1f5cbf8a3336619d5e, {16'd21604, 16'd5662, 16'd35816, 16'd3847, 16'd11013, 16'd57108, 16'd29518, 16'd18241, 16'd22269, 16'd40098, 16'd45413, 16'd33587, 16'd40303, 16'd49314, 16'd40070, 16'd62393, 16'd37201, 16'd1111, 16'd3553, 16'd65216, 16'd22180, 16'd16970, 16'd14452, 16'd33427, 16'd33314, 16'd9751});
	test_expansion(128'hb6e1fc62ab014b31c1f9e46a0d220982, {16'd18769, 16'd53709, 16'd5045, 16'd37640, 16'd27344, 16'd4847, 16'd46305, 16'd40347, 16'd37733, 16'd31630, 16'd22719, 16'd48469, 16'd25604, 16'd11587, 16'd28996, 16'd9320, 16'd29320, 16'd58767, 16'd57891, 16'd22592, 16'd3196, 16'd35819, 16'd37608, 16'd46581, 16'd3116, 16'd15447});
	test_expansion(128'ha7f677677748bcfaae02cd2d4487e959, {16'd2994, 16'd7957, 16'd29103, 16'd52256, 16'd47596, 16'd58833, 16'd29354, 16'd4825, 16'd49248, 16'd4107, 16'd47701, 16'd29374, 16'd26866, 16'd17422, 16'd34073, 16'd52416, 16'd40591, 16'd9020, 16'd38591, 16'd7043, 16'd29659, 16'd54850, 16'd40590, 16'd1662, 16'd32620, 16'd50440});
	test_expansion(128'hfda775f8ec3c8c10122a5888c782ebaf, {16'd38530, 16'd16621, 16'd45032, 16'd46143, 16'd41471, 16'd22162, 16'd34370, 16'd27696, 16'd48489, 16'd9677, 16'd37065, 16'd24880, 16'd34765, 16'd46245, 16'd23939, 16'd1226, 16'd4504, 16'd29235, 16'd60897, 16'd23879, 16'd60836, 16'd15980, 16'd19470, 16'd64270, 16'd17966, 16'd15129});
	test_expansion(128'hd9bc3495490e084a17298c5b74a24bb4, {16'd20369, 16'd32779, 16'd40318, 16'd34732, 16'd60795, 16'd48588, 16'd23702, 16'd56984, 16'd33304, 16'd50579, 16'd13860, 16'd23748, 16'd50727, 16'd55662, 16'd49141, 16'd17692, 16'd47513, 16'd9454, 16'd16147, 16'd3116, 16'd58914, 16'd25581, 16'd57442, 16'd60200, 16'd20356, 16'd21390});
	test_expansion(128'h91043c661a479ee85ce0f5700f1c88b0, {16'd22550, 16'd34590, 16'd21689, 16'd48506, 16'd18239, 16'd5215, 16'd29904, 16'd37318, 16'd46535, 16'd36550, 16'd51969, 16'd25422, 16'd61206, 16'd42681, 16'd2229, 16'd57534, 16'd42331, 16'd20456, 16'd13905, 16'd11830, 16'd63593, 16'd18998, 16'd35964, 16'd44923, 16'd14295, 16'd61036});
	test_expansion(128'hd59bc38dd83049ef340d7f081fca8f82, {16'd8886, 16'd28971, 16'd39551, 16'd54973, 16'd17742, 16'd25295, 16'd49752, 16'd41786, 16'd35316, 16'd35122, 16'd64710, 16'd4243, 16'd26275, 16'd58393, 16'd31500, 16'd61143, 16'd47189, 16'd39895, 16'd24837, 16'd45872, 16'd58945, 16'd17623, 16'd1251, 16'd17391, 16'd61421, 16'd35305});
	test_expansion(128'he8b90a22c21d865f394f89d9fc4a5512, {16'd25953, 16'd19631, 16'd64863, 16'd29455, 16'd53187, 16'd35360, 16'd25935, 16'd62378, 16'd50619, 16'd49908, 16'd32050, 16'd28181, 16'd2357, 16'd2515, 16'd12775, 16'd43715, 16'd18401, 16'd51470, 16'd43645, 16'd44109, 16'd53328, 16'd43799, 16'd54823, 16'd26173, 16'd51715, 16'd5702});
	test_expansion(128'h5de053e8066dbf99b63cfd12c278dac8, {16'd25786, 16'd19486, 16'd19323, 16'd21131, 16'd351, 16'd23807, 16'd2153, 16'd9745, 16'd44855, 16'd40769, 16'd16135, 16'd27608, 16'd33203, 16'd41239, 16'd24819, 16'd64851, 16'd37311, 16'd25791, 16'd58762, 16'd37244, 16'd19241, 16'd33871, 16'd32736, 16'd28333, 16'd7544, 16'd61003});
	test_expansion(128'haa8ea0f8b97acb40a134515fbcf21de3, {16'd13963, 16'd37797, 16'd58077, 16'd30500, 16'd48670, 16'd37232, 16'd47351, 16'd49990, 16'd41851, 16'd52602, 16'd27736, 16'd45775, 16'd32210, 16'd32122, 16'd29208, 16'd62003, 16'd52743, 16'd11077, 16'd26286, 16'd47312, 16'd65059, 16'd65409, 16'd14574, 16'd18595, 16'd58583, 16'd41801});
	test_expansion(128'h9da7e87b633a5febef721e30641be559, {16'd51734, 16'd1646, 16'd7814, 16'd48839, 16'd11042, 16'd7254, 16'd27332, 16'd6771, 16'd24393, 16'd58437, 16'd59654, 16'd38143, 16'd55211, 16'd2261, 16'd34453, 16'd59136, 16'd53801, 16'd43142, 16'd24448, 16'd21629, 16'd4296, 16'd27815, 16'd40037, 16'd48387, 16'd2561, 16'd19842});
	test_expansion(128'hbfe1aa5e1929ee8fd70b81009abbb786, {16'd9674, 16'd36545, 16'd42406, 16'd34069, 16'd16273, 16'd64992, 16'd50561, 16'd63521, 16'd43529, 16'd4111, 16'd13268, 16'd43253, 16'd2422, 16'd35698, 16'd19404, 16'd6826, 16'd33263, 16'd54887, 16'd22570, 16'd1611, 16'd55615, 16'd17096, 16'd23728, 16'd58504, 16'd28032, 16'd60318});
	test_expansion(128'h3121c22be393662244cbf7f197c067f7, {16'd27164, 16'd26344, 16'd51359, 16'd35493, 16'd28914, 16'd36060, 16'd14153, 16'd40619, 16'd55255, 16'd31938, 16'd8530, 16'd40309, 16'd14868, 16'd10320, 16'd2388, 16'd18689, 16'd39142, 16'd9647, 16'd49014, 16'd16899, 16'd14429, 16'd21413, 16'd18300, 16'd21222, 16'd43078, 16'd12605});
	test_expansion(128'hc7aacedebba0ea1d3502217b587f1793, {16'd41486, 16'd9187, 16'd20381, 16'd55035, 16'd60044, 16'd13018, 16'd7678, 16'd12078, 16'd55361, 16'd15437, 16'd43938, 16'd61193, 16'd26645, 16'd53616, 16'd58067, 16'd65077, 16'd34473, 16'd50352, 16'd27380, 16'd16228, 16'd23902, 16'd63330, 16'd38350, 16'd55131, 16'd2271, 16'd19296});
	test_expansion(128'h9eeac8481045b9375c65f774df7dfd95, {16'd55937, 16'd38060, 16'd56545, 16'd1947, 16'd20753, 16'd14666, 16'd8135, 16'd36173, 16'd23899, 16'd12288, 16'd20242, 16'd16704, 16'd58847, 16'd31786, 16'd52254, 16'd42598, 16'd31530, 16'd45885, 16'd7244, 16'd47234, 16'd22530, 16'd42118, 16'd33846, 16'd56869, 16'd24952, 16'd55881});
	test_expansion(128'ha63401be1f51b3d18e3ff948a9d7abd4, {16'd18809, 16'd33816, 16'd4447, 16'd60242, 16'd34442, 16'd15250, 16'd47065, 16'd59106, 16'd11401, 16'd40251, 16'd32838, 16'd62543, 16'd4985, 16'd4129, 16'd5373, 16'd6954, 16'd11508, 16'd48757, 16'd18849, 16'd49742, 16'd10821, 16'd10629, 16'd23484, 16'd29637, 16'd15475, 16'd1216});
	test_expansion(128'hda4daa5d49b92630da756dad14e09cd0, {16'd41019, 16'd33507, 16'd51053, 16'd59282, 16'd62672, 16'd41901, 16'd8832, 16'd17807, 16'd3075, 16'd18387, 16'd6887, 16'd47803, 16'd8141, 16'd9449, 16'd44996, 16'd64829, 16'd60824, 16'd6335, 16'd22615, 16'd3845, 16'd41390, 16'd188, 16'd22393, 16'd19396, 16'd44550, 16'd62922});
	test_expansion(128'hfea1d01bb1979288b5e957a58ef52c49, {16'd17048, 16'd13859, 16'd29370, 16'd27490, 16'd36871, 16'd53210, 16'd58973, 16'd26627, 16'd57801, 16'd56611, 16'd19764, 16'd3842, 16'd43823, 16'd35383, 16'd24459, 16'd58086, 16'd24709, 16'd2618, 16'd62039, 16'd6789, 16'd26423, 16'd17441, 16'd17509, 16'd38631, 16'd1920, 16'd56985});
	test_expansion(128'h4860988517405632454ff6e66cd83047, {16'd46944, 16'd15742, 16'd55836, 16'd7662, 16'd55525, 16'd18992, 16'd6440, 16'd50828, 16'd5716, 16'd21680, 16'd36685, 16'd21953, 16'd33683, 16'd10626, 16'd1040, 16'd22267, 16'd18426, 16'd22732, 16'd63228, 16'd49665, 16'd25176, 16'd64309, 16'd4357, 16'd10781, 16'd41846, 16'd61874});
	test_expansion(128'hc8657d3395d29f0e820ef41fd01beab2, {16'd21401, 16'd54986, 16'd32699, 16'd21946, 16'd44, 16'd37612, 16'd22578, 16'd17486, 16'd63646, 16'd31177, 16'd37592, 16'd10234, 16'd55488, 16'd6001, 16'd59556, 16'd31606, 16'd39107, 16'd51572, 16'd44396, 16'd34020, 16'd60549, 16'd33701, 16'd18060, 16'd54033, 16'd57930, 16'd6098});
	test_expansion(128'hc7796293ef94b2e8e44d295ee0acf6ed, {16'd39672, 16'd18245, 16'd43998, 16'd15321, 16'd29067, 16'd1460, 16'd50427, 16'd55321, 16'd40280, 16'd35772, 16'd50849, 16'd51407, 16'd4772, 16'd60860, 16'd42382, 16'd29309, 16'd39973, 16'd56556, 16'd31056, 16'd41343, 16'd36003, 16'd27440, 16'd46367, 16'd25178, 16'd30383, 16'd21291});
	test_expansion(128'h01b1efc6b47bb2a349883bfe3a055be5, {16'd34326, 16'd60841, 16'd3668, 16'd12413, 16'd13740, 16'd1219, 16'd51970, 16'd37848, 16'd41731, 16'd45302, 16'd20981, 16'd52894, 16'd62803, 16'd17157, 16'd43640, 16'd5088, 16'd14272, 16'd36157, 16'd3763, 16'd53287, 16'd57666, 16'd44646, 16'd30035, 16'd30287, 16'd41476, 16'd13289});
	test_expansion(128'hdfc5d8e605081b67956ae6b6f7cc96fe, {16'd27592, 16'd46329, 16'd23636, 16'd51374, 16'd16936, 16'd54766, 16'd55144, 16'd29077, 16'd48954, 16'd5329, 16'd58487, 16'd29871, 16'd23580, 16'd22568, 16'd56480, 16'd43219, 16'd15944, 16'd42056, 16'd57678, 16'd51022, 16'd24151, 16'd21027, 16'd5855, 16'd55964, 16'd261, 16'd55153});
	test_expansion(128'haf88f46a7f844adfa66ddfa34da4287e, {16'd53614, 16'd45394, 16'd25556, 16'd14621, 16'd57001, 16'd28815, 16'd44973, 16'd38102, 16'd22401, 16'd55660, 16'd10757, 16'd59649, 16'd41391, 16'd21686, 16'd12844, 16'd46167, 16'd55463, 16'd37041, 16'd34512, 16'd57576, 16'd51901, 16'd36530, 16'd30973, 16'd1518, 16'd64463, 16'd50511});
	test_expansion(128'h5f0f1475af5588d0320b4162993e656a, {16'd62166, 16'd30792, 16'd59811, 16'd52752, 16'd10499, 16'd37264, 16'd58692, 16'd53902, 16'd47408, 16'd2129, 16'd55217, 16'd29981, 16'd12367, 16'd19486, 16'd28239, 16'd62095, 16'd29467, 16'd51376, 16'd54831, 16'd33418, 16'd17948, 16'd13602, 16'd2716, 16'd33651, 16'd39516, 16'd60087});
	test_expansion(128'h4f39c387b94d2efc4cd91fc4c912644e, {16'd10148, 16'd5176, 16'd60426, 16'd10209, 16'd8416, 16'd3618, 16'd60167, 16'd24472, 16'd30961, 16'd24968, 16'd34462, 16'd54558, 16'd64879, 16'd50921, 16'd30483, 16'd8244, 16'd45296, 16'd41536, 16'd55789, 16'd36686, 16'd53485, 16'd17716, 16'd11408, 16'd52267, 16'd59163, 16'd62616});
	test_expansion(128'hc9e1853af28ffbc6009e348d50f8bab7, {16'd42826, 16'd14507, 16'd21851, 16'd36920, 16'd24251, 16'd21093, 16'd30661, 16'd53231, 16'd24075, 16'd22318, 16'd49272, 16'd11378, 16'd51175, 16'd9172, 16'd38946, 16'd27283, 16'd45091, 16'd21118, 16'd51194, 16'd20280, 16'd48436, 16'd49682, 16'd36704, 16'd11622, 16'd8753, 16'd682});
	test_expansion(128'h3efb189c78b11b74d87f9f38a0e43242, {16'd42134, 16'd64405, 16'd26678, 16'd34934, 16'd21749, 16'd28669, 16'd59987, 16'd29886, 16'd28066, 16'd46489, 16'd23431, 16'd12687, 16'd9287, 16'd20410, 16'd13085, 16'd6090, 16'd33582, 16'd31068, 16'd24034, 16'd38610, 16'd48041, 16'd33637, 16'd63953, 16'd45547, 16'd43365, 16'd34212});
	test_expansion(128'h583eea7e5d04bddefd8baf6bde05eb3e, {16'd41700, 16'd60183, 16'd57806, 16'd64864, 16'd59022, 16'd15164, 16'd45508, 16'd60568, 16'd18218, 16'd62454, 16'd33697, 16'd60065, 16'd48510, 16'd12517, 16'd30355, 16'd20442, 16'd10800, 16'd1951, 16'd26635, 16'd46813, 16'd3327, 16'd25180, 16'd42427, 16'd43718, 16'd51008, 16'd3700});
	test_expansion(128'hb4dfff21ef9e059c8656bdc84b95ed16, {16'd26617, 16'd4018, 16'd10344, 16'd20742, 16'd22381, 16'd22484, 16'd26761, 16'd11781, 16'd64349, 16'd35201, 16'd14079, 16'd64045, 16'd57550, 16'd4033, 16'd60733, 16'd7934, 16'd24393, 16'd39704, 16'd19387, 16'd12533, 16'd32220, 16'd63859, 16'd38591, 16'd2402, 16'd30927, 16'd16008});
	test_expansion(128'hb3c95eb016b899061107b8750f2afd5b, {16'd61816, 16'd25754, 16'd54375, 16'd3468, 16'd11826, 16'd21168, 16'd10021, 16'd42785, 16'd9956, 16'd796, 16'd28861, 16'd34458, 16'd59916, 16'd49253, 16'd32555, 16'd21600, 16'd1523, 16'd6473, 16'd64581, 16'd3565, 16'd14295, 16'd22272, 16'd31791, 16'd52583, 16'd56325, 16'd4949});
	test_expansion(128'h1541fdd1404c95f4039abbe52f45ad79, {16'd58958, 16'd36970, 16'd8282, 16'd48276, 16'd50181, 16'd17978, 16'd25409, 16'd38197, 16'd36262, 16'd53418, 16'd1961, 16'd54168, 16'd44206, 16'd48129, 16'd4743, 16'd27034, 16'd16459, 16'd2955, 16'd15422, 16'd16108, 16'd61886, 16'd15697, 16'd36584, 16'd64280, 16'd12317, 16'd26584});
	test_expansion(128'h779956f656d22cd5bb7b0fdd8dc2266b, {16'd57802, 16'd48981, 16'd26156, 16'd6349, 16'd8817, 16'd36694, 16'd52830, 16'd12551, 16'd23848, 16'd37536, 16'd20594, 16'd34784, 16'd42141, 16'd33935, 16'd3520, 16'd25478, 16'd49508, 16'd13876, 16'd1995, 16'd24798, 16'd46477, 16'd47009, 16'd42911, 16'd34939, 16'd39086, 16'd48843});
	test_expansion(128'h54a1786ac08003b3e8602cf278727747, {16'd9115, 16'd18419, 16'd63657, 16'd55666, 16'd1432, 16'd33096, 16'd27571, 16'd25373, 16'd14439, 16'd1729, 16'd15066, 16'd34005, 16'd29650, 16'd3173, 16'd14204, 16'd58867, 16'd34648, 16'd56813, 16'd6718, 16'd9039, 16'd51865, 16'd24238, 16'd44704, 16'd62847, 16'd12703, 16'd40792});
	test_expansion(128'h88cc514e94ebb9daf30e28c8dc6f9e3f, {16'd6955, 16'd48335, 16'd52598, 16'd56553, 16'd64631, 16'd24444, 16'd18171, 16'd58243, 16'd35479, 16'd63775, 16'd41579, 16'd10055, 16'd53263, 16'd12290, 16'd54231, 16'd60272, 16'd16252, 16'd39836, 16'd13826, 16'd41378, 16'd48540, 16'd12910, 16'd18089, 16'd11074, 16'd47174, 16'd42874});
	test_expansion(128'hf9cc6504e1c9fd3b3f42f9ab92f78bf5, {16'd24262, 16'd39806, 16'd51270, 16'd56166, 16'd54031, 16'd65103, 16'd44315, 16'd4222, 16'd38124, 16'd11897, 16'd64203, 16'd10864, 16'd47293, 16'd57538, 16'd60623, 16'd41171, 16'd33163, 16'd42758, 16'd14208, 16'd30736, 16'd10082, 16'd14480, 16'd25465, 16'd60159, 16'd12443, 16'd8266});
	test_expansion(128'h912e4cd9816191681a69020ffdd90a0e, {16'd38143, 16'd10193, 16'd59667, 16'd24655, 16'd26080, 16'd40306, 16'd9402, 16'd1632, 16'd49029, 16'd31344, 16'd18813, 16'd6098, 16'd15026, 16'd7823, 16'd2675, 16'd39681, 16'd38059, 16'd30755, 16'd135, 16'd14195, 16'd56426, 16'd24912, 16'd15218, 16'd53837, 16'd8076, 16'd9993});
	test_expansion(128'h187a58fb080231c9166f19055f8aa9c0, {16'd40172, 16'd28576, 16'd42887, 16'd48416, 16'd64899, 16'd611, 16'd44954, 16'd55047, 16'd14824, 16'd40560, 16'd191, 16'd14797, 16'd11925, 16'd47691, 16'd6502, 16'd8542, 16'd64348, 16'd42611, 16'd40389, 16'd4201, 16'd37850, 16'd59695, 16'd12302, 16'd20218, 16'd32357, 16'd8651});
	test_expansion(128'hb4587a619c16a8e995db859732931f37, {16'd35440, 16'd26824, 16'd13310, 16'd38402, 16'd18168, 16'd53851, 16'd62309, 16'd34007, 16'd380, 16'd20673, 16'd1781, 16'd59471, 16'd36410, 16'd5031, 16'd22721, 16'd48469, 16'd1434, 16'd60435, 16'd13868, 16'd2087, 16'd3231, 16'd3196, 16'd44830, 16'd2251, 16'd42114, 16'd13157});
	test_expansion(128'hb4ba0b019492489c6808d3b23487c3bf, {16'd44244, 16'd7291, 16'd58494, 16'd25472, 16'd59441, 16'd16176, 16'd27809, 16'd47439, 16'd15602, 16'd1476, 16'd3487, 16'd55847, 16'd48555, 16'd26383, 16'd26262, 16'd42326, 16'd32194, 16'd60789, 16'd7127, 16'd32339, 16'd21741, 16'd1450, 16'd26303, 16'd25906, 16'd22388, 16'd6455});
	test_expansion(128'hc67c56e68e0c9bef7b9eeafdb63dab5d, {16'd7454, 16'd44990, 16'd20813, 16'd4730, 16'd46913, 16'd36086, 16'd7787, 16'd48847, 16'd62235, 16'd8365, 16'd45800, 16'd39152, 16'd42066, 16'd7112, 16'd59858, 16'd22658, 16'd16019, 16'd44328, 16'd54016, 16'd22916, 16'd37023, 16'd22793, 16'd25049, 16'd64128, 16'd6166, 16'd22902});
	test_expansion(128'h6dd55ad96413bee133af86260d6d5e51, {16'd40011, 16'd31604, 16'd33144, 16'd19324, 16'd16616, 16'd32109, 16'd24833, 16'd47233, 16'd52809, 16'd63745, 16'd2765, 16'd5478, 16'd58955, 16'd13233, 16'd50133, 16'd51130, 16'd40805, 16'd44308, 16'd43421, 16'd43067, 16'd42233, 16'd45536, 16'd44977, 16'd10230, 16'd7795, 16'd12363});
	test_expansion(128'h07ac7343a0d0cb8ee10bbb1647db5364, {16'd26176, 16'd58511, 16'd10673, 16'd42002, 16'd59493, 16'd47723, 16'd47265, 16'd44486, 16'd34779, 16'd31886, 16'd38113, 16'd25445, 16'd59493, 16'd57395, 16'd3164, 16'd5166, 16'd5947, 16'd8570, 16'd10196, 16'd44872, 16'd49943, 16'd65434, 16'd6516, 16'd16629, 16'd47991, 16'd12913});
	test_expansion(128'h14f04fa2d235edc6e125efcd99ced078, {16'd43666, 16'd8133, 16'd46922, 16'd36528, 16'd3818, 16'd1136, 16'd48530, 16'd4711, 16'd59406, 16'd54920, 16'd61380, 16'd31687, 16'd8840, 16'd42605, 16'd44941, 16'd13619, 16'd48101, 16'd46088, 16'd59475, 16'd61591, 16'd63855, 16'd34871, 16'd35656, 16'd21455, 16'd42723, 16'd61491});
	test_expansion(128'h394456b7af5305b5b7f497a4a5d99845, {16'd21306, 16'd52246, 16'd48500, 16'd35264, 16'd64528, 16'd28088, 16'd37037, 16'd7415, 16'd42052, 16'd64845, 16'd11962, 16'd12721, 16'd14957, 16'd63460, 16'd1463, 16'd33948, 16'd52853, 16'd52780, 16'd22440, 16'd7858, 16'd27322, 16'd62119, 16'd20424, 16'd38147, 16'd54893, 16'd24604});
	test_expansion(128'h26df01c686b06f86564e26695b3a747a, {16'd58017, 16'd48167, 16'd53400, 16'd49991, 16'd57057, 16'd37308, 16'd10071, 16'd36719, 16'd33748, 16'd48032, 16'd64701, 16'd26207, 16'd10195, 16'd64649, 16'd46759, 16'd15761, 16'd38100, 16'd19131, 16'd60742, 16'd51146, 16'd46307, 16'd63633, 16'd62013, 16'd54088, 16'd47937, 16'd41424});
	test_expansion(128'h008691ca359d90801c1d1e8e17f4e948, {16'd6262, 16'd24998, 16'd19150, 16'd53912, 16'd31895, 16'd10519, 16'd24099, 16'd36814, 16'd40708, 16'd1263, 16'd62989, 16'd36152, 16'd64415, 16'd29264, 16'd19609, 16'd33522, 16'd16205, 16'd12991, 16'd863, 16'd49039, 16'd30639, 16'd56733, 16'd45287, 16'd44479, 16'd59227, 16'd26246});
	test_expansion(128'h81db845a6476e62f5ac99fae4f2bc1e4, {16'd54789, 16'd21872, 16'd36746, 16'd7561, 16'd22814, 16'd48755, 16'd15142, 16'd55509, 16'd13809, 16'd62663, 16'd1598, 16'd36415, 16'd34019, 16'd20202, 16'd33773, 16'd47557, 16'd55610, 16'd2581, 16'd17628, 16'd63040, 16'd5290, 16'd33771, 16'd57218, 16'd11974, 16'd9182, 16'd14632});
	test_expansion(128'he586f884bc21b82a5dc99fc4701bbfdb, {16'd48652, 16'd46713, 16'd37468, 16'd29675, 16'd31595, 16'd27, 16'd26442, 16'd10883, 16'd33364, 16'd40222, 16'd6854, 16'd34792, 16'd42037, 16'd22638, 16'd12650, 16'd37873, 16'd44813, 16'd38, 16'd6950, 16'd12868, 16'd21966, 16'd4882, 16'd16570, 16'd53727, 16'd6557, 16'd19196});
	test_expansion(128'h65bb3d02777653f86acf0ea57c16a709, {16'd56718, 16'd62235, 16'd5888, 16'd11415, 16'd34095, 16'd38080, 16'd30191, 16'd21187, 16'd24718, 16'd22138, 16'd56184, 16'd26072, 16'd22144, 16'd35162, 16'd58933, 16'd226, 16'd43867, 16'd52647, 16'd19319, 16'd12187, 16'd48170, 16'd53935, 16'd26618, 16'd22536, 16'd6195, 16'd9918});
	test_expansion(128'h1f502283582fb1036ac788aee60ff215, {16'd64181, 16'd63124, 16'd48654, 16'd59630, 16'd16846, 16'd30110, 16'd56913, 16'd53598, 16'd65331, 16'd55778, 16'd62501, 16'd42272, 16'd63688, 16'd48479, 16'd5135, 16'd3574, 16'd58523, 16'd14262, 16'd64548, 16'd37724, 16'd53062, 16'd21246, 16'd64622, 16'd64559, 16'd30420, 16'd3679});
	test_expansion(128'h9ee696832eba1ab32f71a25d5ef0eb60, {16'd33170, 16'd57270, 16'd7615, 16'd12399, 16'd20787, 16'd14133, 16'd42365, 16'd20370, 16'd37229, 16'd58066, 16'd27063, 16'd16877, 16'd9410, 16'd45298, 16'd15550, 16'd24842, 16'd18084, 16'd62508, 16'd42198, 16'd50231, 16'd62964, 16'd44881, 16'd53558, 16'd21571, 16'd14628, 16'd41922});
	test_expansion(128'h5a5391f7a313f2b4bca3eed64a5aa565, {16'd2496, 16'd54812, 16'd32817, 16'd32524, 16'd3147, 16'd55873, 16'd26607, 16'd45163, 16'd44718, 16'd22729, 16'd9299, 16'd3236, 16'd53467, 16'd14951, 16'd1893, 16'd47266, 16'd11201, 16'd22562, 16'd49021, 16'd56312, 16'd7973, 16'd40905, 16'd45493, 16'd27513, 16'd59054, 16'd10136});
	test_expansion(128'ha3079313fa4252a92ef1360698575e92, {16'd30968, 16'd2606, 16'd10614, 16'd35654, 16'd50782, 16'd41119, 16'd56486, 16'd53249, 16'd42506, 16'd62605, 16'd54300, 16'd48304, 16'd20931, 16'd47483, 16'd54534, 16'd43243, 16'd21484, 16'd33712, 16'd43039, 16'd29987, 16'd27433, 16'd8118, 16'd23147, 16'd29147, 16'd19928, 16'd64777});
	test_expansion(128'h1f13e080b7ee01641170bb4e9fcfaeb2, {16'd62423, 16'd3901, 16'd40126, 16'd46504, 16'd14822, 16'd16930, 16'd21144, 16'd53995, 16'd30001, 16'd38344, 16'd58180, 16'd59723, 16'd44080, 16'd19572, 16'd23570, 16'd33774, 16'd17233, 16'd30967, 16'd15407, 16'd17587, 16'd612, 16'd47542, 16'd11417, 16'd56460, 16'd50316, 16'd14652});
	test_expansion(128'h56211ebf39d5099e76dfdb2371216f05, {16'd54553, 16'd9297, 16'd33606, 16'd40203, 16'd5985, 16'd12800, 16'd5447, 16'd60174, 16'd22152, 16'd22702, 16'd60764, 16'd62481, 16'd29105, 16'd50686, 16'd49826, 16'd10380, 16'd48859, 16'd19061, 16'd54496, 16'd7175, 16'd45180, 16'd18938, 16'd54529, 16'd51765, 16'd17139, 16'd54570});
	test_expansion(128'h516490d450c227a755e1293b581f9ecd, {16'd30979, 16'd33836, 16'd26721, 16'd56749, 16'd658, 16'd52871, 16'd7757, 16'd61349, 16'd36610, 16'd28261, 16'd29929, 16'd19313, 16'd27275, 16'd63190, 16'd47392, 16'd8586, 16'd44888, 16'd26913, 16'd52551, 16'd11960, 16'd51325, 16'd60182, 16'd6810, 16'd64999, 16'd36736, 16'd56359});
	test_expansion(128'h2913d04a93ecabd882a9d768f26008e6, {16'd37670, 16'd45564, 16'd17071, 16'd62287, 16'd52623, 16'd19489, 16'd51443, 16'd16455, 16'd12175, 16'd51404, 16'd24977, 16'd53468, 16'd20285, 16'd26806, 16'd10576, 16'd5725, 16'd37868, 16'd14204, 16'd44987, 16'd31198, 16'd58471, 16'd7481, 16'd31628, 16'd36924, 16'd26861, 16'd5469});
	test_expansion(128'he70790a4d1a5cbb6fbead728e21d456f, {16'd36066, 16'd32650, 16'd8436, 16'd51630, 16'd27878, 16'd52376, 16'd15427, 16'd54178, 16'd57238, 16'd34809, 16'd10251, 16'd9095, 16'd38924, 16'd7041, 16'd10796, 16'd51579, 16'd4334, 16'd46877, 16'd36517, 16'd33503, 16'd20511, 16'd45984, 16'd13729, 16'd48043, 16'd29842, 16'd34548});
	test_expansion(128'hd9df588473b0918fc1bf9680d331c6fb, {16'd23482, 16'd57207, 16'd13523, 16'd17625, 16'd33735, 16'd6765, 16'd60769, 16'd59682, 16'd14236, 16'd27640, 16'd45790, 16'd50639, 16'd61036, 16'd24342, 16'd49551, 16'd9704, 16'd28013, 16'd63384, 16'd48494, 16'd4098, 16'd26644, 16'd18863, 16'd45255, 16'd48353, 16'd36584, 16'd30169});
	test_expansion(128'h540b81c6e284999de9845dbd22df9304, {16'd30090, 16'd9005, 16'd28049, 16'd10712, 16'd48770, 16'd47847, 16'd47657, 16'd13540, 16'd40479, 16'd37885, 16'd40077, 16'd65188, 16'd54367, 16'd631, 16'd39733, 16'd13876, 16'd6360, 16'd7607, 16'd55299, 16'd35532, 16'd63605, 16'd30040, 16'd954, 16'd27924, 16'd52243, 16'd52030});
	test_expansion(128'h6598380aa55e6c5fa411e7b9e0f2f497, {16'd54239, 16'd50554, 16'd7321, 16'd15375, 16'd25451, 16'd8660, 16'd62785, 16'd37266, 16'd9172, 16'd47954, 16'd54346, 16'd22845, 16'd2211, 16'd22351, 16'd24275, 16'd2461, 16'd15307, 16'd49997, 16'd22065, 16'd44770, 16'd11877, 16'd55401, 16'd48139, 16'd54695, 16'd24349, 16'd7128});
	test_expansion(128'h0ec305b6f6c0395160f20d14fff094b0, {16'd268, 16'd29124, 16'd20612, 16'd9469, 16'd34732, 16'd34086, 16'd24082, 16'd13757, 16'd19548, 16'd58850, 16'd32640, 16'd36255, 16'd39879, 16'd19212, 16'd32647, 16'd52704, 16'd5352, 16'd58431, 16'd55094, 16'd52567, 16'd45090, 16'd42951, 16'd15847, 16'd32168, 16'd9429, 16'd48890});
	test_expansion(128'hce1b9313558129f18d9279615eacccaa, {16'd52778, 16'd38483, 16'd61223, 16'd7644, 16'd27521, 16'd22417, 16'd5431, 16'd59293, 16'd30233, 16'd18167, 16'd8908, 16'd42041, 16'd32460, 16'd40905, 16'd47234, 16'd52933, 16'd33824, 16'd45044, 16'd23357, 16'd59869, 16'd45951, 16'd46410, 16'd40578, 16'd8107, 16'd26898, 16'd13737});
	test_expansion(128'h72d8f3960f6f5761987ec9020fa4383a, {16'd60741, 16'd41914, 16'd46594, 16'd27260, 16'd45615, 16'd8216, 16'd11487, 16'd65481, 16'd39733, 16'd56344, 16'd13417, 16'd23233, 16'd58609, 16'd45077, 16'd56237, 16'd3919, 16'd32956, 16'd1027, 16'd26542, 16'd48343, 16'd23320, 16'd22933, 16'd11774, 16'd44156, 16'd52809, 16'd62011});
	test_expansion(128'h2d2a2445dd7ec87b07d5ed532fe2777f, {16'd50268, 16'd8160, 16'd59009, 16'd43425, 16'd25441, 16'd36536, 16'd63600, 16'd37238, 16'd25347, 16'd30513, 16'd45223, 16'd54794, 16'd52154, 16'd39200, 16'd48158, 16'd54272, 16'd57920, 16'd58216, 16'd44478, 16'd42984, 16'd9754, 16'd43886, 16'd183, 16'd49514, 16'd10610, 16'd65415});
	test_expansion(128'h40bf22c3484b9654ac1d7568d08d7355, {16'd43781, 16'd63921, 16'd2502, 16'd49675, 16'd19765, 16'd42949, 16'd53624, 16'd4396, 16'd59458, 16'd2590, 16'd64362, 16'd3325, 16'd59253, 16'd10999, 16'd21939, 16'd58071, 16'd25432, 16'd51771, 16'd31071, 16'd6444, 16'd51241, 16'd40598, 16'd43790, 16'd41535, 16'd18906, 16'd5522});
	test_expansion(128'ha1ec45aa5100268503b01561cc222fc0, {16'd24928, 16'd15472, 16'd19893, 16'd40715, 16'd6421, 16'd16008, 16'd42962, 16'd41639, 16'd47911, 16'd15878, 16'd59681, 16'd56522, 16'd33615, 16'd31339, 16'd37159, 16'd49468, 16'd6622, 16'd49431, 16'd22958, 16'd58397, 16'd8615, 16'd48139, 16'd35907, 16'd50849, 16'd51123, 16'd13442});
	test_expansion(128'h691bc9f61eaafa2f8d2c697f9b859543, {16'd6124, 16'd26906, 16'd40747, 16'd59330, 16'd2294, 16'd48849, 16'd19430, 16'd33868, 16'd42185, 16'd32286, 16'd14711, 16'd13017, 16'd30061, 16'd7395, 16'd36215, 16'd52018, 16'd6040, 16'd13667, 16'd624, 16'd25972, 16'd36729, 16'd57061, 16'd24056, 16'd31576, 16'd3779, 16'd732});
	test_expansion(128'h39e9e88c2a796f93f30e2ff259f85bc6, {16'd30602, 16'd44441, 16'd59575, 16'd63363, 16'd14203, 16'd58757, 16'd60189, 16'd8841, 16'd10810, 16'd7838, 16'd13265, 16'd17821, 16'd38937, 16'd3087, 16'd20029, 16'd31115, 16'd36257, 16'd2720, 16'd52688, 16'd42991, 16'd32549, 16'd58078, 16'd33955, 16'd29185, 16'd4890, 16'd12738});
	test_expansion(128'h7b0d9683893799f5710e17dea15dc9ab, {16'd47947, 16'd9117, 16'd42851, 16'd48558, 16'd3359, 16'd47926, 16'd5995, 16'd15103, 16'd53417, 16'd5679, 16'd55462, 16'd45711, 16'd22673, 16'd61672, 16'd54228, 16'd43262, 16'd32133, 16'd8879, 16'd53500, 16'd8069, 16'd62058, 16'd22253, 16'd63434, 16'd59834, 16'd52060, 16'd34005});
	test_expansion(128'h37a7fe32efaf8aafb04fc29fa5a3e9fc, {16'd58278, 16'd22789, 16'd23468, 16'd46983, 16'd46341, 16'd30392, 16'd24488, 16'd18620, 16'd57011, 16'd63738, 16'd32260, 16'd19401, 16'd17572, 16'd16436, 16'd3510, 16'd54498, 16'd30850, 16'd16671, 16'd56036, 16'd52178, 16'd55519, 16'd3478, 16'd18495, 16'd16157, 16'd37351, 16'd19141});
	test_expansion(128'h27a400e32932790c41d0f93a3eaed9fa, {16'd19410, 16'd24582, 16'd33032, 16'd6986, 16'd9214, 16'd22217, 16'd62509, 16'd29997, 16'd40006, 16'd3910, 16'd5010, 16'd51835, 16'd63259, 16'd53419, 16'd63699, 16'd24625, 16'd17725, 16'd442, 16'd187, 16'd7489, 16'd51724, 16'd39340, 16'd42903, 16'd14908, 16'd64807, 16'd22061});
	test_expansion(128'h2f0c558d79d6f24d88fd00f6bb03ed55, {16'd16575, 16'd60717, 16'd13065, 16'd53937, 16'd28744, 16'd53922, 16'd15862, 16'd43598, 16'd23689, 16'd41765, 16'd32546, 16'd50436, 16'd21751, 16'd13934, 16'd19853, 16'd39703, 16'd8511, 16'd33872, 16'd43054, 16'd52829, 16'd64102, 16'd54957, 16'd63216, 16'd19317, 16'd50588, 16'd22036});
	test_expansion(128'hfca1ef7349aa6870cd833264ada1db4a, {16'd55284, 16'd42620, 16'd44748, 16'd27865, 16'd57845, 16'd60400, 16'd10772, 16'd30026, 16'd44079, 16'd13469, 16'd28059, 16'd9595, 16'd49335, 16'd37569, 16'd41859, 16'd15536, 16'd60155, 16'd58918, 16'd57701, 16'd31950, 16'd41906, 16'd45126, 16'd38950, 16'd38337, 16'd13945, 16'd37968});
	test_expansion(128'h1f47075da2c0957e1a96123103c5f41b, {16'd22047, 16'd36185, 16'd47070, 16'd18959, 16'd11957, 16'd2205, 16'd43831, 16'd52305, 16'd41215, 16'd16910, 16'd8183, 16'd54820, 16'd40229, 16'd18350, 16'd46071, 16'd17584, 16'd55324, 16'd39182, 16'd51016, 16'd24324, 16'd55544, 16'd56134, 16'd9235, 16'd57169, 16'd15538, 16'd6233});
	test_expansion(128'h6f733ea13de48bb4de9ab93c773b9f8b, {16'd54497, 16'd42621, 16'd41078, 16'd40147, 16'd19919, 16'd33817, 16'd17462, 16'd36452, 16'd16416, 16'd6932, 16'd48083, 16'd8133, 16'd45237, 16'd139, 16'd45253, 16'd15333, 16'd1661, 16'd51428, 16'd22164, 16'd47498, 16'd374, 16'd58859, 16'd28632, 16'd35279, 16'd51245, 16'd18024});
	test_expansion(128'h86f28770f7d1e0216ab4f831a05702fd, {16'd26180, 16'd22549, 16'd29929, 16'd40359, 16'd54084, 16'd6947, 16'd53476, 16'd21991, 16'd63106, 16'd1080, 16'd46522, 16'd57737, 16'd11842, 16'd51523, 16'd8562, 16'd7922, 16'd10788, 16'd14528, 16'd63482, 16'd35150, 16'd47326, 16'd62491, 16'd51912, 16'd6014, 16'd55541, 16'd12103});
	test_expansion(128'hb132170c1791f4fe0a2272f9ecfee41a, {16'd26551, 16'd60943, 16'd56917, 16'd65111, 16'd5078, 16'd32900, 16'd64324, 16'd15364, 16'd2293, 16'd29130, 16'd49079, 16'd5659, 16'd20037, 16'd55675, 16'd27361, 16'd55969, 16'd57669, 16'd51043, 16'd18835, 16'd30894, 16'd5620, 16'd46361, 16'd39465, 16'd11237, 16'd6639, 16'd3319});
	test_expansion(128'h05fed590a89e119cd06f71456937da45, {16'd40916, 16'd42755, 16'd14141, 16'd57183, 16'd32644, 16'd64603, 16'd4145, 16'd42714, 16'd1405, 16'd56262, 16'd9373, 16'd7114, 16'd61320, 16'd10204, 16'd9341, 16'd4702, 16'd6226, 16'd24032, 16'd39751, 16'd51002, 16'd25720, 16'd14708, 16'd62855, 16'd19558, 16'd39248, 16'd6343});
	test_expansion(128'h0a79c6bb45cff65c73132330c5263ce6, {16'd7200, 16'd46242, 16'd8961, 16'd57571, 16'd39224, 16'd55965, 16'd45293, 16'd43785, 16'd10021, 16'd26500, 16'd21128, 16'd44823, 16'd24702, 16'd41623, 16'd40513, 16'd34403, 16'd5920, 16'd12475, 16'd48851, 16'd11934, 16'd36201, 16'd27492, 16'd31239, 16'd12990, 16'd12218, 16'd33914});
	test_expansion(128'h3ddbade4ef00918f3e5cc19af20b7679, {16'd16426, 16'd59767, 16'd32685, 16'd4945, 16'd9989, 16'd17266, 16'd65319, 16'd3878, 16'd63105, 16'd2016, 16'd44901, 16'd62514, 16'd55025, 16'd3571, 16'd12128, 16'd9601, 16'd43820, 16'd18029, 16'd43938, 16'd25637, 16'd54985, 16'd4337, 16'd15898, 16'd54056, 16'd64404, 16'd34237});
	test_expansion(128'hb0c31dee1befe20c84f72eb014cb067e, {16'd46402, 16'd38906, 16'd60233, 16'd42171, 16'd37230, 16'd21991, 16'd38540, 16'd48499, 16'd11747, 16'd48824, 16'd17238, 16'd15292, 16'd55166, 16'd41942, 16'd37186, 16'd40315, 16'd49316, 16'd35317, 16'd59597, 16'd18117, 16'd40248, 16'd19076, 16'd54849, 16'd5721, 16'd52851, 16'd904});
	test_expansion(128'h7da0140f5045b32dd643075045ab4938, {16'd24458, 16'd2495, 16'd36799, 16'd39261, 16'd47895, 16'd29952, 16'd4012, 16'd46189, 16'd52901, 16'd31179, 16'd55423, 16'd40180, 16'd41057, 16'd7899, 16'd48967, 16'd56051, 16'd24629, 16'd618, 16'd49150, 16'd27569, 16'd56050, 16'd44923, 16'd8516, 16'd59371, 16'd60706, 16'd11185});
	test_expansion(128'hb3739bc476d01d31918caa064f44d184, {16'd16911, 16'd48688, 16'd347, 16'd17009, 16'd62356, 16'd39718, 16'd4771, 16'd58354, 16'd17759, 16'd4748, 16'd14154, 16'd47845, 16'd56618, 16'd35192, 16'd17696, 16'd57823, 16'd8156, 16'd45374, 16'd65081, 16'd51031, 16'd30023, 16'd30418, 16'd13487, 16'd30673, 16'd5044, 16'd33264});
	test_expansion(128'h882ed8309565e3dd4b35e3d1b4f0bd75, {16'd48133, 16'd44579, 16'd17189, 16'd12347, 16'd37900, 16'd39968, 16'd17978, 16'd18822, 16'd13933, 16'd16684, 16'd23486, 16'd44339, 16'd17951, 16'd32113, 16'd39149, 16'd4502, 16'd3440, 16'd59096, 16'd38453, 16'd8335, 16'd43895, 16'd24739, 16'd8143, 16'd23325, 16'd20303, 16'd5463});
	test_expansion(128'h49635e9d9eccb8a403bc92879b8405c8, {16'd61044, 16'd46506, 16'd12431, 16'd22564, 16'd10458, 16'd13376, 16'd340, 16'd710, 16'd63051, 16'd54066, 16'd21041, 16'd23347, 16'd57800, 16'd52543, 16'd13916, 16'd7074, 16'd36551, 16'd54013, 16'd13830, 16'd57747, 16'd10022, 16'd5170, 16'd13483, 16'd18535, 16'd32776, 16'd59778});
	test_expansion(128'hbafd0c91dbded3cafdc0e8196d0f3e49, {16'd33218, 16'd5287, 16'd17636, 16'd43480, 16'd36699, 16'd48916, 16'd52862, 16'd44619, 16'd34945, 16'd29539, 16'd6526, 16'd12179, 16'd52051, 16'd59347, 16'd14459, 16'd39638, 16'd33593, 16'd40909, 16'd49844, 16'd20002, 16'd56227, 16'd54469, 16'd29708, 16'd24654, 16'd62403, 16'd54848});
	test_expansion(128'hc4c2e45ec9ad2a0735a100c0130c83dd, {16'd2954, 16'd88, 16'd9213, 16'd1124, 16'd29076, 16'd1590, 16'd33031, 16'd44695, 16'd57735, 16'd35599, 16'd40756, 16'd39878, 16'd22998, 16'd2636, 16'd23208, 16'd6326, 16'd12377, 16'd1509, 16'd50152, 16'd58275, 16'd32662, 16'd23394, 16'd2432, 16'd65054, 16'd51543, 16'd32694});
	test_expansion(128'ha6214d829fb81e692730b4fcac8c2c72, {16'd64732, 16'd5888, 16'd51963, 16'd47376, 16'd48400, 16'd38414, 16'd45062, 16'd28658, 16'd44970, 16'd46191, 16'd32880, 16'd34046, 16'd4931, 16'd41741, 16'd764, 16'd21747, 16'd11421, 16'd12539, 16'd39529, 16'd30289, 16'd59799, 16'd48037, 16'd10492, 16'd25718, 16'd50533, 16'd13292});
	test_expansion(128'h6a10c37605bed5c7c734452b287999c5, {16'd27787, 16'd58271, 16'd6906, 16'd23642, 16'd62842, 16'd18848, 16'd28740, 16'd16820, 16'd14591, 16'd59364, 16'd7215, 16'd7244, 16'd13138, 16'd5433, 16'd25423, 16'd10261, 16'd49869, 16'd28282, 16'd25261, 16'd28356, 16'd19663, 16'd10337, 16'd37190, 16'd32783, 16'd26214, 16'd35334});
	test_expansion(128'h8063d9636a3562467be2c23d6d992a02, {16'd55657, 16'd6887, 16'd54333, 16'd41457, 16'd24431, 16'd29884, 16'd59940, 16'd49789, 16'd7281, 16'd11149, 16'd42691, 16'd59760, 16'd22102, 16'd32942, 16'd65391, 16'd49775, 16'd12447, 16'd46204, 16'd27563, 16'd4670, 16'd60550, 16'd34561, 16'd56504, 16'd33517, 16'd29651, 16'd48148});
	test_expansion(128'hdb38d89f6198e2544115ff73d77821b4, {16'd30140, 16'd21072, 16'd28213, 16'd5797, 16'd28385, 16'd17898, 16'd13432, 16'd55822, 16'd59339, 16'd24799, 16'd32484, 16'd12560, 16'd52844, 16'd9636, 16'd46170, 16'd7023, 16'd45221, 16'd63605, 16'd26716, 16'd56040, 16'd36089, 16'd8681, 16'd44924, 16'd19916, 16'd7247, 16'd65163});
	test_expansion(128'h5dca562a9ca3829cfd99d097970072d4, {16'd44871, 16'd22439, 16'd17673, 16'd22006, 16'd65081, 16'd50505, 16'd47033, 16'd22405, 16'd49687, 16'd55314, 16'd59108, 16'd63174, 16'd38415, 16'd16545, 16'd41465, 16'd13419, 16'd35486, 16'd46414, 16'd38363, 16'd43528, 16'd7173, 16'd38784, 16'd10954, 16'd20990, 16'd27439, 16'd59931});
	test_expansion(128'he8def6bbefd5b87495aaac76a5aa0f0f, {16'd8452, 16'd17118, 16'd27871, 16'd56533, 16'd34535, 16'd64601, 16'd508, 16'd24156, 16'd55116, 16'd49019, 16'd63884, 16'd25543, 16'd9485, 16'd24877, 16'd64992, 16'd5638, 16'd16279, 16'd6352, 16'd9209, 16'd911, 16'd53482, 16'd29753, 16'd4667, 16'd61308, 16'd19013, 16'd24234});
	test_expansion(128'had73e813b0ca159d884b07f95498224f, {16'd11739, 16'd5444, 16'd55035, 16'd12772, 16'd22779, 16'd31539, 16'd63792, 16'd25433, 16'd21661, 16'd52532, 16'd46743, 16'd52220, 16'd57525, 16'd32389, 16'd30016, 16'd28638, 16'd65063, 16'd10988, 16'd14056, 16'd14482, 16'd28374, 16'd56550, 16'd44726, 16'd24474, 16'd56175, 16'd24092});
	test_expansion(128'hef749ad8dec0155d322fb21f77618d46, {16'd24183, 16'd59395, 16'd25240, 16'd1968, 16'd18547, 16'd35176, 16'd40872, 16'd43450, 16'd58332, 16'd62422, 16'd63871, 16'd30418, 16'd37729, 16'd17184, 16'd38523, 16'd33381, 16'd22385, 16'd61284, 16'd16590, 16'd19827, 16'd51955, 16'd1726, 16'd64568, 16'd63404, 16'd38370, 16'd30759});
	test_expansion(128'h2e07fe436020fbf18d32581b988f5265, {16'd59065, 16'd54160, 16'd21958, 16'd3016, 16'd17585, 16'd47842, 16'd33533, 16'd46723, 16'd372, 16'd6945, 16'd6743, 16'd20134, 16'd41440, 16'd23934, 16'd10870, 16'd32925, 16'd53086, 16'd14845, 16'd12979, 16'd12954, 16'd2210, 16'd25768, 16'd24077, 16'd5152, 16'd60712, 16'd25709});
	test_expansion(128'h69f9c3ef36d10f7399c00f48723c1453, {16'd18263, 16'd50249, 16'd8761, 16'd37171, 16'd11250, 16'd27600, 16'd34111, 16'd29598, 16'd64555, 16'd20609, 16'd42558, 16'd269, 16'd53007, 16'd34036, 16'd20248, 16'd51863, 16'd35495, 16'd24179, 16'd62973, 16'd6790, 16'd54640, 16'd49270, 16'd61858, 16'd56685, 16'd57313, 16'd56998});
	test_expansion(128'hb41da7dcaf08042d085def4f6c796c03, {16'd34920, 16'd39830, 16'd41899, 16'd24421, 16'd14207, 16'd48652, 16'd63508, 16'd51438, 16'd51766, 16'd13673, 16'd33586, 16'd23540, 16'd478, 16'd54404, 16'd11536, 16'd16449, 16'd28741, 16'd16316, 16'd33000, 16'd11102, 16'd31079, 16'd38420, 16'd23908, 16'd45899, 16'd26181, 16'd38304});
	test_expansion(128'h90634919ea416b64cd58f4eb293222c1, {16'd9970, 16'd38519, 16'd5462, 16'd6429, 16'd28935, 16'd38651, 16'd45197, 16'd26178, 16'd7875, 16'd54450, 16'd835, 16'd39027, 16'd56802, 16'd47560, 16'd22244, 16'd12811, 16'd10957, 16'd18430, 16'd32317, 16'd54870, 16'd7028, 16'd35453, 16'd52585, 16'd31085, 16'd31887, 16'd57920});
	test_expansion(128'h04c7548df7c9f2a9229444c1a494b18a, {16'd28777, 16'd60097, 16'd11758, 16'd9269, 16'd1435, 16'd56922, 16'd64740, 16'd8880, 16'd49506, 16'd64376, 16'd17219, 16'd15831, 16'd14011, 16'd18501, 16'd15104, 16'd50565, 16'd45895, 16'd18088, 16'd3290, 16'd50639, 16'd55762, 16'd45535, 16'd40893, 16'd47271, 16'd26204, 16'd6437});
	test_expansion(128'h305314718e8ec3b47bc8e8866a4ae7e3, {16'd56372, 16'd47201, 16'd32571, 16'd36747, 16'd9393, 16'd18707, 16'd20839, 16'd49628, 16'd29529, 16'd65029, 16'd58172, 16'd63893, 16'd54921, 16'd6245, 16'd61993, 16'd35335, 16'd37992, 16'd29283, 16'd17047, 16'd36001, 16'd62316, 16'd37520, 16'd41217, 16'd27552, 16'd28599, 16'd50591});
	test_expansion(128'h916b0d1bc8ec465f537680538b1f8209, {16'd1727, 16'd2438, 16'd32891, 16'd33043, 16'd37732, 16'd29954, 16'd7789, 16'd16451, 16'd4596, 16'd48463, 16'd62959, 16'd46875, 16'd61987, 16'd57681, 16'd5428, 16'd18609, 16'd42863, 16'd43012, 16'd19348, 16'd57881, 16'd47385, 16'd15969, 16'd16353, 16'd11762, 16'd62862, 16'd8497});
	test_expansion(128'hed301b48049e250f105c8fe989f7a206, {16'd6079, 16'd37303, 16'd37739, 16'd49292, 16'd39739, 16'd56119, 16'd43008, 16'd56805, 16'd33896, 16'd43426, 16'd3689, 16'd64560, 16'd43891, 16'd19425, 16'd37117, 16'd27752, 16'd35594, 16'd49238, 16'd15450, 16'd24073, 16'd38870, 16'd37682, 16'd21394, 16'd65184, 16'd55838, 16'd49750});
	test_expansion(128'h6c218667187c64f62af1ce5de115c6cb, {16'd42931, 16'd50044, 16'd10431, 16'd37688, 16'd31147, 16'd51195, 16'd10510, 16'd29035, 16'd37507, 16'd45579, 16'd4919, 16'd3416, 16'd58192, 16'd759, 16'd18404, 16'd3345, 16'd21828, 16'd49344, 16'd11833, 16'd3958, 16'd61687, 16'd64024, 16'd29612, 16'd42682, 16'd10484, 16'd53134});
	test_expansion(128'h3d248675a3315251a10c21d73a64735d, {16'd55270, 16'd47046, 16'd65223, 16'd63607, 16'd47240, 16'd65280, 16'd6768, 16'd58491, 16'd7040, 16'd52909, 16'd39065, 16'd63214, 16'd25236, 16'd26708, 16'd13303, 16'd59975, 16'd45980, 16'd20344, 16'd45477, 16'd39153, 16'd21903, 16'd31320, 16'd41442, 16'd32899, 16'd32548, 16'd41635});
	test_expansion(128'hd32dddab8a86ca475289957f0495114f, {16'd19777, 16'd24462, 16'd14683, 16'd54027, 16'd26757, 16'd20628, 16'd43850, 16'd29581, 16'd50154, 16'd49789, 16'd9510, 16'd7776, 16'd62880, 16'd29703, 16'd57673, 16'd41182, 16'd28181, 16'd17936, 16'd35476, 16'd40759, 16'd16306, 16'd21653, 16'd57002, 16'd47672, 16'd29074, 16'd45554});
	test_expansion(128'h7007586292580fba1280b39fbc1af5f9, {16'd45010, 16'd54749, 16'd28240, 16'd64887, 16'd12587, 16'd63, 16'd29359, 16'd39181, 16'd65284, 16'd61605, 16'd63129, 16'd8032, 16'd28784, 16'd20928, 16'd14715, 16'd39898, 16'd16775, 16'd36119, 16'd52680, 16'd55849, 16'd51963, 16'd10348, 16'd18915, 16'd15290, 16'd5035, 16'd23831});
	test_expansion(128'h8891693c54103dc3ac1534418c45ec25, {16'd5682, 16'd49226, 16'd10601, 16'd12922, 16'd48755, 16'd10178, 16'd57396, 16'd45016, 16'd34546, 16'd23903, 16'd50263, 16'd34370, 16'd44571, 16'd62584, 16'd30230, 16'd32772, 16'd50368, 16'd27555, 16'd65207, 16'd58297, 16'd28110, 16'd43731, 16'd21421, 16'd5180, 16'd41693, 16'd32045});
	test_expansion(128'h3c8d8e7a80d35e7f74779654c2f30fb2, {16'd59497, 16'd16348, 16'd13238, 16'd6316, 16'd24295, 16'd12641, 16'd45896, 16'd9059, 16'd55456, 16'd12786, 16'd42708, 16'd56020, 16'd926, 16'd61698, 16'd1024, 16'd52668, 16'd744, 16'd49817, 16'd62733, 16'd7941, 16'd10925, 16'd33009, 16'd4861, 16'd5587, 16'd30933, 16'd55505});
	test_expansion(128'h8c2181d3ab9d4a4640db690ffa5a5960, {16'd44453, 16'd39006, 16'd58301, 16'd31158, 16'd59326, 16'd40001, 16'd3392, 16'd57816, 16'd59312, 16'd55319, 16'd20359, 16'd10074, 16'd37019, 16'd14689, 16'd9942, 16'd17375, 16'd8213, 16'd13659, 16'd35372, 16'd41485, 16'd37562, 16'd34489, 16'd7935, 16'd40946, 16'd38716, 16'd3916});
	test_expansion(128'h180be1af0f37f45d4d820b5c20082e32, {16'd24112, 16'd8881, 16'd25623, 16'd301, 16'd32729, 16'd36694, 16'd18465, 16'd24702, 16'd13374, 16'd64872, 16'd63114, 16'd7874, 16'd54932, 16'd438, 16'd11261, 16'd36716, 16'd15324, 16'd21710, 16'd45556, 16'd61409, 16'd26604, 16'd8204, 16'd17192, 16'd3513, 16'd11260, 16'd64041});
	test_expansion(128'ha350cba7e547084d3cd8d9e9544de88a, {16'd28017, 16'd44048, 16'd64783, 16'd15552, 16'd9222, 16'd56481, 16'd20094, 16'd41385, 16'd60938, 16'd65313, 16'd6571, 16'd35174, 16'd34634, 16'd60243, 16'd51079, 16'd997, 16'd30288, 16'd22391, 16'd42970, 16'd63957, 16'd26810, 16'd26120, 16'd31929, 16'd18450, 16'd26062, 16'd12});
	test_expansion(128'h33fc37df1a376a8ab83d9172546773a5, {16'd41828, 16'd6359, 16'd60315, 16'd426, 16'd9594, 16'd34170, 16'd40921, 16'd57051, 16'd48455, 16'd39824, 16'd43020, 16'd32192, 16'd28734, 16'd10474, 16'd35775, 16'd17408, 16'd58147, 16'd10989, 16'd34660, 16'd33342, 16'd49435, 16'd59437, 16'd1248, 16'd10309, 16'd57794, 16'd17552});
	test_expansion(128'h82440ade1e9e3e995c12e4529f6d491d, {16'd36735, 16'd30942, 16'd2206, 16'd50835, 16'd64544, 16'd33784, 16'd48720, 16'd34831, 16'd34117, 16'd954, 16'd24498, 16'd32106, 16'd12803, 16'd24990, 16'd44753, 16'd52279, 16'd42503, 16'd3231, 16'd37632, 16'd33489, 16'd44722, 16'd3706, 16'd44269, 16'd11633, 16'd56882, 16'd57310});
	test_expansion(128'hfa56c73c31dd74797aa2b5894315e438, {16'd48714, 16'd16684, 16'd59034, 16'd14590, 16'd51542, 16'd19586, 16'd9896, 16'd9576, 16'd55973, 16'd36139, 16'd62591, 16'd1385, 16'd52618, 16'd46139, 16'd12296, 16'd43553, 16'd46508, 16'd29452, 16'd5341, 16'd51509, 16'd57387, 16'd37448, 16'd18307, 16'd3052, 16'd43965, 16'd260});
	test_expansion(128'he4f2db26dc6133071dfd050713e1e3b1, {16'd3576, 16'd6009, 16'd61096, 16'd61489, 16'd22545, 16'd37127, 16'd19339, 16'd5612, 16'd5213, 16'd28854, 16'd1354, 16'd39432, 16'd20655, 16'd14804, 16'd38754, 16'd49353, 16'd403, 16'd13013, 16'd6217, 16'd42160, 16'd50540, 16'd33566, 16'd12438, 16'd8377, 16'd11564, 16'd16132});
	test_expansion(128'h799372ef2ff1c905909f395427fe89ca, {16'd62018, 16'd60320, 16'd40599, 16'd15085, 16'd56051, 16'd54354, 16'd54252, 16'd5239, 16'd53268, 16'd29451, 16'd29855, 16'd18859, 16'd22246, 16'd5088, 16'd47852, 16'd61159, 16'd21984, 16'd23215, 16'd58881, 16'd28038, 16'd20991, 16'd62809, 16'd1771, 16'd55329, 16'd7906, 16'd64858});
	test_expansion(128'h2b2362009c74dc4be1e5c56830640748, {16'd16194, 16'd57935, 16'd42019, 16'd9175, 16'd42110, 16'd16361, 16'd10048, 16'd8540, 16'd6247, 16'd25260, 16'd42545, 16'd38219, 16'd34501, 16'd27633, 16'd59611, 16'd43033, 16'd44190, 16'd7462, 16'd41217, 16'd63938, 16'd24960, 16'd16314, 16'd20501, 16'd56465, 16'd39899, 16'd34736});
	test_expansion(128'hcf2533ce36744252acb6cc25d91f5b3d, {16'd3181, 16'd60605, 16'd4068, 16'd58704, 16'd51643, 16'd12745, 16'd28648, 16'd32084, 16'd2583, 16'd45529, 16'd19416, 16'd5092, 16'd57308, 16'd35449, 16'd8754, 16'd55880, 16'd43316, 16'd6537, 16'd57254, 16'd61355, 16'd39239, 16'd60621, 16'd719, 16'd16099, 16'd46312, 16'd9961});
	test_expansion(128'h4f9eb0d9948bec5f45ef9a59e060e59c, {16'd4334, 16'd8064, 16'd32120, 16'd30509, 16'd30242, 16'd54806, 16'd46544, 16'd56428, 16'd12583, 16'd50280, 16'd2442, 16'd41490, 16'd51197, 16'd16429, 16'd50860, 16'd11849, 16'd31165, 16'd29115, 16'd51574, 16'd43650, 16'd20068, 16'd51981, 16'd5707, 16'd28754, 16'd7974, 16'd58799});
	test_expansion(128'h07436bddb877b9b31ee596593b889f73, {16'd17828, 16'd2192, 16'd45138, 16'd6685, 16'd25226, 16'd29398, 16'd63695, 16'd34914, 16'd48791, 16'd19059, 16'd26398, 16'd57233, 16'd44619, 16'd30750, 16'd35875, 16'd41538, 16'd33619, 16'd52778, 16'd679, 16'd9853, 16'd31452, 16'd36152, 16'd53515, 16'd53047, 16'd55047, 16'd25998});
	test_expansion(128'hcf70303e83cc5bf355fdacf57b2b62da, {16'd16011, 16'd45726, 16'd22222, 16'd54060, 16'd3932, 16'd42669, 16'd51205, 16'd9632, 16'd53933, 16'd55848, 16'd2941, 16'd5751, 16'd48210, 16'd37153, 16'd1100, 16'd12657, 16'd20572, 16'd50949, 16'd56745, 16'd45904, 16'd32476, 16'd64197, 16'd48606, 16'd8914, 16'd56482, 16'd31714});
	test_expansion(128'hab0a07737af96052a9964fafee6add5a, {16'd22285, 16'd27197, 16'd41695, 16'd7389, 16'd9016, 16'd2251, 16'd50780, 16'd63008, 16'd38385, 16'd38393, 16'd23032, 16'd26261, 16'd12764, 16'd45189, 16'd14815, 16'd21575, 16'd8922, 16'd25199, 16'd63800, 16'd64386, 16'd8899, 16'd9229, 16'd33446, 16'd2400, 16'd14109, 16'd46612});
	test_expansion(128'h1db55423b741c5f4040f54bb79e513f7, {16'd15186, 16'd48396, 16'd54379, 16'd47341, 16'd41761, 16'd32838, 16'd39909, 16'd50623, 16'd59761, 16'd28776, 16'd15070, 16'd92, 16'd33845, 16'd30062, 16'd9450, 16'd12607, 16'd40649, 16'd54567, 16'd6866, 16'd22831, 16'd28444, 16'd11124, 16'd30207, 16'd38161, 16'd62266, 16'd22568});
	test_expansion(128'h728f3662bc80cbd0ad6f733e511cf971, {16'd48806, 16'd4896, 16'd10179, 16'd59694, 16'd27261, 16'd48980, 16'd53880, 16'd42114, 16'd2745, 16'd63216, 16'd28800, 16'd20998, 16'd10021, 16'd31436, 16'd6046, 16'd36741, 16'd25949, 16'd51563, 16'd48315, 16'd11015, 16'd3337, 16'd16553, 16'd45846, 16'd34509, 16'd40019, 16'd20718});
	test_expansion(128'h7e31a990233febe0e5c64e3f50400afb, {16'd21171, 16'd64010, 16'd22463, 16'd8192, 16'd19548, 16'd43549, 16'd43865, 16'd6748, 16'd35691, 16'd42387, 16'd64164, 16'd27596, 16'd3237, 16'd44828, 16'd22544, 16'd40741, 16'd60867, 16'd26401, 16'd55117, 16'd28003, 16'd30585, 16'd19023, 16'd25600, 16'd14917, 16'd17347, 16'd47979});
	test_expansion(128'h57d2e5fff32a90e0d9709b02fcdf3446, {16'd42481, 16'd45155, 16'd42613, 16'd47534, 16'd24319, 16'd55457, 16'd15447, 16'd8434, 16'd31062, 16'd8610, 16'd63829, 16'd5963, 16'd39871, 16'd2286, 16'd59725, 16'd55401, 16'd57974, 16'd35030, 16'd43129, 16'd36133, 16'd44903, 16'd37976, 16'd39648, 16'd42610, 16'd15897, 16'd7231});
	test_expansion(128'h7b3d722c89e38d8bf3dd4d4a8155a6c7, {16'd53318, 16'd53987, 16'd8190, 16'd3652, 16'd61244, 16'd14268, 16'd53856, 16'd57296, 16'd59237, 16'd7331, 16'd17923, 16'd3528, 16'd29236, 16'd320, 16'd29474, 16'd3413, 16'd18270, 16'd4705, 16'd26581, 16'd40013, 16'd265, 16'd46222, 16'd21023, 16'd11651, 16'd34475, 16'd51521});
	test_expansion(128'h4bc7740d10c71cf198c38e8e807c1c05, {16'd24017, 16'd58691, 16'd8929, 16'd25476, 16'd37102, 16'd56564, 16'd51006, 16'd5960, 16'd33320, 16'd914, 16'd20814, 16'd64427, 16'd29003, 16'd60620, 16'd51064, 16'd14670, 16'd50520, 16'd19060, 16'd28893, 16'd59671, 16'd52405, 16'd40351, 16'd43386, 16'd29554, 16'd24337, 16'd2857});
	test_expansion(128'h8488ebe58880d62918c7de14e3109b2c, {16'd35420, 16'd42019, 16'd28256, 16'd48054, 16'd24042, 16'd63163, 16'd27838, 16'd23566, 16'd27485, 16'd24325, 16'd8416, 16'd37312, 16'd32839, 16'd35960, 16'd55053, 16'd43784, 16'd12137, 16'd27090, 16'd54422, 16'd52270, 16'd18695, 16'd927, 16'd55098, 16'd59504, 16'd25601, 16'd1533});
	test_expansion(128'h290404a883e6dc78226d363cf189e510, {16'd42248, 16'd60825, 16'd6741, 16'd58596, 16'd42393, 16'd19636, 16'd47782, 16'd55456, 16'd31239, 16'd41742, 16'd2721, 16'd26228, 16'd35715, 16'd24266, 16'd28841, 16'd38146, 16'd45634, 16'd27692, 16'd58143, 16'd2611, 16'd19396, 16'd12102, 16'd54571, 16'd8123, 16'd60646, 16'd10730});
	test_expansion(128'hb06428d2c0c1c94a1975fc7023da5445, {16'd10339, 16'd36746, 16'd10898, 16'd60323, 16'd65199, 16'd10836, 16'd49898, 16'd4378, 16'd28281, 16'd11142, 16'd45962, 16'd51811, 16'd37998, 16'd52638, 16'd32276, 16'd22325, 16'd29995, 16'd27343, 16'd56202, 16'd45151, 16'd57577, 16'd23586, 16'd5003, 16'd56187, 16'd6805, 16'd28742});
	test_expansion(128'hc3c6d1b25d16bafd1d89b34faf617cd0, {16'd1607, 16'd64215, 16'd14992, 16'd58153, 16'd43942, 16'd37533, 16'd27305, 16'd39314, 16'd39169, 16'd64244, 16'd34742, 16'd45309, 16'd38087, 16'd53873, 16'd8820, 16'd26517, 16'd37802, 16'd63818, 16'd56886, 16'd56579, 16'd43836, 16'd47283, 16'd33324, 16'd61257, 16'd1424, 16'd42800});
	test_expansion(128'hab60d8a7336f534075bcad4d1cbd742a, {16'd27307, 16'd250, 16'd13674, 16'd58116, 16'd23002, 16'd19493, 16'd29413, 16'd59498, 16'd35117, 16'd25179, 16'd22875, 16'd47993, 16'd61612, 16'd4212, 16'd383, 16'd37362, 16'd9328, 16'd29075, 16'd18298, 16'd28341, 16'd41245, 16'd36066, 16'd16297, 16'd48459, 16'd37425, 16'd54098});
	test_expansion(128'h4e756fe9ac40ee4045f641131f971b4d, {16'd42969, 16'd24774, 16'd12398, 16'd1168, 16'd64687, 16'd1106, 16'd53310, 16'd62529, 16'd19684, 16'd14188, 16'd17031, 16'd7674, 16'd9806, 16'd18084, 16'd55989, 16'd6990, 16'd2090, 16'd1761, 16'd59787, 16'd7, 16'd29263, 16'd59033, 16'd53962, 16'd28509, 16'd55197, 16'd52679});
	test_expansion(128'hada6434d746bddb6cfa5c7a205c75470, {16'd55235, 16'd27027, 16'd55804, 16'd11835, 16'd49153, 16'd40390, 16'd12403, 16'd37279, 16'd35578, 16'd5202, 16'd26535, 16'd62212, 16'd51763, 16'd51793, 16'd11756, 16'd26550, 16'd22776, 16'd58087, 16'd42602, 16'd48733, 16'd9177, 16'd55397, 16'd3920, 16'd38864, 16'd20012, 16'd8136});
	test_expansion(128'hff2ac9048024c53485d3bba8ac9b9071, {16'd47275, 16'd23877, 16'd12540, 16'd4235, 16'd11430, 16'd23660, 16'd9395, 16'd11268, 16'd27697, 16'd20786, 16'd21953, 16'd43726, 16'd29859, 16'd50673, 16'd26803, 16'd54810, 16'd30813, 16'd32297, 16'd12354, 16'd57861, 16'd39269, 16'd24308, 16'd30581, 16'd15895, 16'd1111, 16'd30191});
	test_expansion(128'h04d38030bb9e31c7dc928cd18ae2fa07, {16'd21393, 16'd22694, 16'd42862, 16'd10403, 16'd63244, 16'd53298, 16'd53027, 16'd54376, 16'd41321, 16'd64068, 16'd9437, 16'd6491, 16'd2233, 16'd43941, 16'd23127, 16'd28797, 16'd57038, 16'd20171, 16'd63403, 16'd48944, 16'd1434, 16'd41160, 16'd1165, 16'd35231, 16'd36814, 16'd31096});
	test_expansion(128'h4976795da10953d6b83c76682d500925, {16'd46964, 16'd53675, 16'd44028, 16'd32839, 16'd25652, 16'd62309, 16'd62368, 16'd57197, 16'd15165, 16'd40355, 16'd30840, 16'd58632, 16'd31187, 16'd28896, 16'd51112, 16'd48177, 16'd61694, 16'd22700, 16'd8769, 16'd48335, 16'd36491, 16'd37760, 16'd61161, 16'd15763, 16'd1401, 16'd56190});
	test_expansion(128'ha281c1a9c984bb274e6bf306add128f4, {16'd14490, 16'd5702, 16'd44805, 16'd21553, 16'd45522, 16'd41911, 16'd15940, 16'd33695, 16'd39314, 16'd31925, 16'd36104, 16'd48381, 16'd55840, 16'd57829, 16'd32696, 16'd59361, 16'd61038, 16'd34927, 16'd64607, 16'd487, 16'd38492, 16'd57663, 16'd30162, 16'd64349, 16'd51893, 16'd15327});
	test_expansion(128'h6a7f96b8c8547565f37cc1868c921b2a, {16'd31158, 16'd42891, 16'd34526, 16'd59814, 16'd42785, 16'd18880, 16'd63364, 16'd34189, 16'd51167, 16'd31536, 16'd1726, 16'd60430, 16'd64845, 16'd33886, 16'd57542, 16'd61614, 16'd27907, 16'd58734, 16'd7253, 16'd22579, 16'd57475, 16'd43551, 16'd59207, 16'd11353, 16'd37832, 16'd16440});
	test_expansion(128'h3823db99dc0268110633910d75ae5dc4, {16'd856, 16'd17309, 16'd49458, 16'd47982, 16'd30450, 16'd45446, 16'd29885, 16'd49586, 16'd6477, 16'd8267, 16'd58018, 16'd22118, 16'd34483, 16'd13532, 16'd51924, 16'd42946, 16'd33447, 16'd57320, 16'd55300, 16'd36238, 16'd7252, 16'd51489, 16'd23344, 16'd6993, 16'd2933, 16'd14352});
	test_expansion(128'hb56c1d4945da97e32a7dc6090b69a25a, {16'd54223, 16'd46406, 16'd4825, 16'd28063, 16'd16709, 16'd56123, 16'd47514, 16'd42294, 16'd43711, 16'd110, 16'd40942, 16'd58210, 16'd4403, 16'd33209, 16'd22922, 16'd59008, 16'd28098, 16'd40637, 16'd23957, 16'd20840, 16'd2438, 16'd37845, 16'd14879, 16'd34804, 16'd46221, 16'd2495});
	test_expansion(128'h9f6534fb73891aa0851e45fe8f8107c5, {16'd13606, 16'd22582, 16'd64840, 16'd48462, 16'd60343, 16'd51966, 16'd55543, 16'd43304, 16'd13741, 16'd43570, 16'd53126, 16'd4010, 16'd5683, 16'd31210, 16'd26682, 16'd9391, 16'd4484, 16'd44499, 16'd18825, 16'd10177, 16'd34419, 16'd7968, 16'd19628, 16'd41863, 16'd53155, 16'd19538});
	test_expansion(128'h065d71247fde936378bd36f2f02b5082, {16'd9540, 16'd14083, 16'd34843, 16'd4017, 16'd52280, 16'd50942, 16'd56210, 16'd13836, 16'd28892, 16'd16410, 16'd37361, 16'd28533, 16'd34720, 16'd32150, 16'd23401, 16'd18639, 16'd10167, 16'd10749, 16'd63796, 16'd31825, 16'd41819, 16'd19986, 16'd11760, 16'd61744, 16'd42454, 16'd10731});
	test_expansion(128'h063888383c7780f2ce3057783a2c7122, {16'd3478, 16'd23201, 16'd8142, 16'd9059, 16'd19097, 16'd12146, 16'd60590, 16'd23230, 16'd35124, 16'd13964, 16'd48517, 16'd44556, 16'd9040, 16'd15377, 16'd4663, 16'd37243, 16'd23781, 16'd47674, 16'd12267, 16'd39082, 16'd5395, 16'd64067, 16'd31440, 16'd41598, 16'd41555, 16'd31219});
	test_expansion(128'h17307fc2c0baf242b4696b6095b0e7cc, {16'd50476, 16'd23426, 16'd45028, 16'd6210, 16'd29212, 16'd52812, 16'd34627, 16'd9019, 16'd24349, 16'd39907, 16'd54912, 16'd6343, 16'd28089, 16'd35379, 16'd47458, 16'd63335, 16'd24408, 16'd55379, 16'd38544, 16'd40030, 16'd31657, 16'd60458, 16'd30197, 16'd41441, 16'd29107, 16'd41549});
	test_expansion(128'h6dc0cfab46877fe3a63118b89b9a8476, {16'd16570, 16'd30000, 16'd36802, 16'd64277, 16'd64475, 16'd22787, 16'd59975, 16'd5436, 16'd48909, 16'd8587, 16'd24049, 16'd63744, 16'd22775, 16'd44323, 16'd1148, 16'd53707, 16'd52951, 16'd12872, 16'd7022, 16'd46360, 16'd30796, 16'd1378, 16'd23201, 16'd23125, 16'd52802, 16'd14001});
	test_expansion(128'h0e1424069b44e148fc02d922b2771438, {16'd54925, 16'd57612, 16'd17223, 16'd44186, 16'd46010, 16'd56099, 16'd44593, 16'd17704, 16'd15485, 16'd25448, 16'd42001, 16'd28758, 16'd62870, 16'd61969, 16'd45789, 16'd15726, 16'd13350, 16'd41414, 16'd10877, 16'd39369, 16'd44866, 16'd8889, 16'd4520, 16'd42151, 16'd20870, 16'd48762});
	test_expansion(128'h0f19c78bc60267c54e7af7a8e4f258b4, {16'd22476, 16'd8408, 16'd39225, 16'd20486, 16'd51890, 16'd56195, 16'd57374, 16'd24609, 16'd9977, 16'd6528, 16'd6137, 16'd47655, 16'd1452, 16'd4382, 16'd33574, 16'd43200, 16'd48896, 16'd51704, 16'd14138, 16'd20094, 16'd28874, 16'd10047, 16'd41675, 16'd8369, 16'd24332, 16'd51366});
	test_expansion(128'hb029e145e2ce3d853f1bb490ef1e98b5, {16'd50851, 16'd2271, 16'd50318, 16'd44262, 16'd10135, 16'd22041, 16'd27050, 16'd27495, 16'd32204, 16'd44339, 16'd22497, 16'd36942, 16'd8205, 16'd35283, 16'd40583, 16'd28384, 16'd43398, 16'd42415, 16'd49012, 16'd4981, 16'd31954, 16'd45982, 16'd7226, 16'd12543, 16'd17314, 16'd46241});
	test_expansion(128'hc02ab97466ad8712f60fec9079c39342, {16'd2204, 16'd53120, 16'd57308, 16'd44134, 16'd42267, 16'd29976, 16'd20642, 16'd47560, 16'd17703, 16'd59585, 16'd11256, 16'd30040, 16'd57658, 16'd30306, 16'd20378, 16'd49119, 16'd23269, 16'd48196, 16'd12553, 16'd54878, 16'd5979, 16'd50420, 16'd62194, 16'd19531, 16'd42942, 16'd11673});
	test_expansion(128'hff32f84dfbc401c442c89eb3f66546ba, {16'd15231, 16'd28997, 16'd9710, 16'd17270, 16'd4153, 16'd13237, 16'd22330, 16'd6439, 16'd63156, 16'd18957, 16'd7614, 16'd63252, 16'd15288, 16'd30786, 16'd25641, 16'd17643, 16'd18657, 16'd547, 16'd31622, 16'd39421, 16'd41724, 16'd15472, 16'd54481, 16'd53234, 16'd3319, 16'd15770});
	test_expansion(128'ha8bbc69f48157984d5b21ef6fdadad92, {16'd3615, 16'd37464, 16'd53024, 16'd48853, 16'd21578, 16'd9396, 16'd40089, 16'd27202, 16'd29839, 16'd6179, 16'd32341, 16'd2586, 16'd21771, 16'd39102, 16'd48577, 16'd8378, 16'd37088, 16'd63861, 16'd36974, 16'd42100, 16'd50714, 16'd17550, 16'd21350, 16'd33427, 16'd51754, 16'd46624});
	test_expansion(128'hb4d374368d00e4e300d70c7bd62874dc, {16'd36133, 16'd42257, 16'd44920, 16'd9399, 16'd24713, 16'd56316, 16'd11910, 16'd11583, 16'd41684, 16'd975, 16'd2213, 16'd64292, 16'd17253, 16'd59009, 16'd50651, 16'd51930, 16'd19575, 16'd25394, 16'd61997, 16'd37728, 16'd35945, 16'd5528, 16'd25330, 16'd28698, 16'd60012, 16'd44026});
	test_expansion(128'ha8ca8bd785089bcff6282719180ae583, {16'd52241, 16'd46077, 16'd44552, 16'd208, 16'd8603, 16'd15800, 16'd6838, 16'd14020, 16'd21016, 16'd27614, 16'd52487, 16'd29666, 16'd2067, 16'd13121, 16'd32511, 16'd47344, 16'd21902, 16'd21397, 16'd55994, 16'd64123, 16'd62890, 16'd29807, 16'd62896, 16'd29266, 16'd22306, 16'd36867});
	test_expansion(128'h8e47674caff01881bd7b89f96d4f7fa2, {16'd32409, 16'd65013, 16'd58539, 16'd59950, 16'd61308, 16'd20416, 16'd146, 16'd48080, 16'd58716, 16'd54561, 16'd40281, 16'd34176, 16'd48140, 16'd31535, 16'd43505, 16'd22151, 16'd15241, 16'd40697, 16'd7110, 16'd19284, 16'd44291, 16'd40919, 16'd46452, 16'd23822, 16'd55587, 16'd51464});
	test_expansion(128'h83165b81c811ec840b11044372c58236, {16'd22655, 16'd34483, 16'd14434, 16'd12779, 16'd42268, 16'd37038, 16'd37732, 16'd14570, 16'd37315, 16'd58639, 16'd48902, 16'd38, 16'd37834, 16'd9398, 16'd13714, 16'd56592, 16'd27392, 16'd12105, 16'd39781, 16'd50385, 16'd8788, 16'd9254, 16'd43701, 16'd36410, 16'd53573, 16'd20349});
	test_expansion(128'h07aa4a1bf8789a1acdbf7beb743fc03d, {16'd61582, 16'd41688, 16'd37232, 16'd51939, 16'd21646, 16'd58183, 16'd15911, 16'd17475, 16'd45369, 16'd42043, 16'd9251, 16'd9244, 16'd5974, 16'd12536, 16'd37396, 16'd40178, 16'd19745, 16'd2531, 16'd661, 16'd22719, 16'd18100, 16'd47868, 16'd36730, 16'd65406, 16'd32459, 16'd28902});
	test_expansion(128'h69c35b03b44a4ee2c1040cd67ee68709, {16'd20324, 16'd52223, 16'd45313, 16'd14053, 16'd31013, 16'd24586, 16'd25624, 16'd27959, 16'd61223, 16'd43288, 16'd37869, 16'd47879, 16'd30949, 16'd47360, 16'd53781, 16'd15630, 16'd60667, 16'd59934, 16'd33074, 16'd38413, 16'd50345, 16'd1599, 16'd1108, 16'd23074, 16'd31899, 16'd23715});
	test_expansion(128'he0e9f55a95135dd43c8f9184469de5be, {16'd23081, 16'd37773, 16'd6990, 16'd4279, 16'd3252, 16'd10213, 16'd27410, 16'd15117, 16'd22061, 16'd44125, 16'd64677, 16'd17220, 16'd42643, 16'd59739, 16'd34681, 16'd41871, 16'd39372, 16'd28964, 16'd58655, 16'd36710, 16'd34229, 16'd64231, 16'd38627, 16'd42660, 16'd41967, 16'd2242});
	test_expansion(128'h8788f5165e837aaf6c8b8c937f38d156, {16'd8420, 16'd20853, 16'd51489, 16'd51270, 16'd60957, 16'd14368, 16'd62642, 16'd37110, 16'd14152, 16'd28862, 16'd23958, 16'd61185, 16'd27723, 16'd4765, 16'd60029, 16'd48298, 16'd43853, 16'd42661, 16'd9021, 16'd38222, 16'd9855, 16'd33083, 16'd9851, 16'd29440, 16'd25616, 16'd47565});
	test_expansion(128'hcc488b3820327996d2a47054580909c5, {16'd37086, 16'd41621, 16'd52029, 16'd23364, 16'd4086, 16'd13965, 16'd21901, 16'd45481, 16'd58004, 16'd18835, 16'd378, 16'd32791, 16'd25109, 16'd60345, 16'd19452, 16'd8830, 16'd62506, 16'd25538, 16'd55889, 16'd16245, 16'd212, 16'd61551, 16'd6207, 16'd20528, 16'd58389, 16'd6450});
	test_expansion(128'h135d7ccb9cd3811aa59c3d26817f6e00, {16'd28749, 16'd34808, 16'd7021, 16'd10958, 16'd62389, 16'd37757, 16'd22602, 16'd42868, 16'd9841, 16'd47166, 16'd48679, 16'd49049, 16'd15617, 16'd7133, 16'd28662, 16'd29760, 16'd40200, 16'd21112, 16'd64949, 16'd29138, 16'd5236, 16'd30075, 16'd31176, 16'd10504, 16'd49049, 16'd3086});
	test_expansion(128'h22534edc8be2e758680213301748ceb3, {16'd65484, 16'd44210, 16'd63561, 16'd53967, 16'd36784, 16'd36447, 16'd61725, 16'd53261, 16'd58255, 16'd22196, 16'd50679, 16'd33568, 16'd10933, 16'd33162, 16'd55932, 16'd26995, 16'd4517, 16'd58228, 16'd1541, 16'd53070, 16'd9921, 16'd8404, 16'd6006, 16'd24996, 16'd64021, 16'd2952});
	test_expansion(128'h740fb489566e56b08a8d6de65f424a4f, {16'd48395, 16'd15559, 16'd5261, 16'd55188, 16'd62209, 16'd50332, 16'd50180, 16'd38999, 16'd405, 16'd56122, 16'd27390, 16'd48734, 16'd18331, 16'd14714, 16'd14374, 16'd16787, 16'd30566, 16'd24554, 16'd42743, 16'd47687, 16'd36461, 16'd34617, 16'd764, 16'd20229, 16'd1794, 16'd62112});
	test_expansion(128'h32898372cd76ad51f58044a2eeaf08a3, {16'd39306, 16'd61832, 16'd12871, 16'd10710, 16'd50457, 16'd2098, 16'd35199, 16'd29057, 16'd1880, 16'd23031, 16'd642, 16'd33719, 16'd22513, 16'd8198, 16'd11471, 16'd14509, 16'd16378, 16'd29258, 16'd6977, 16'd65263, 16'd57826, 16'd6239, 16'd51596, 16'd48023, 16'd57255, 16'd34755});
	test_expansion(128'h4cadb220e177a468c7b9493de7e61e71, {16'd37675, 16'd28782, 16'd46657, 16'd56511, 16'd53215, 16'd25383, 16'd20806, 16'd12849, 16'd32562, 16'd10891, 16'd41136, 16'd39539, 16'd37352, 16'd35645, 16'd1221, 16'd18169, 16'd8912, 16'd14826, 16'd63619, 16'd58105, 16'd14027, 16'd40533, 16'd24677, 16'd55848, 16'd20617, 16'd50422});
	test_expansion(128'h560873a4be38f87e7b8f313a887fe47b, {16'd55200, 16'd23723, 16'd46506, 16'd17560, 16'd62988, 16'd5660, 16'd56519, 16'd53662, 16'd37937, 16'd34949, 16'd765, 16'd57846, 16'd13479, 16'd35550, 16'd9289, 16'd45379, 16'd35077, 16'd10332, 16'd23004, 16'd7833, 16'd32349, 16'd32194, 16'd50949, 16'd5611, 16'd64795, 16'd22867});
	test_expansion(128'hee46f07bc9e4a8a8b30f261112d6f243, {16'd55657, 16'd43982, 16'd18907, 16'd54769, 16'd60920, 16'd48128, 16'd7800, 16'd64302, 16'd15610, 16'd38278, 16'd42263, 16'd54299, 16'd3632, 16'd42250, 16'd27025, 16'd65252, 16'd37202, 16'd15307, 16'd12523, 16'd13619, 16'd9305, 16'd60155, 16'd8568, 16'd56564, 16'd36783, 16'd21719});
	test_expansion(128'h59464de2436bc99ea075c461b5d5c2c1, {16'd21498, 16'd37426, 16'd21164, 16'd52752, 16'd39749, 16'd30285, 16'd60390, 16'd12162, 16'd32063, 16'd33541, 16'd33539, 16'd57965, 16'd6700, 16'd38050, 16'd7672, 16'd2415, 16'd14160, 16'd24324, 16'd27655, 16'd19156, 16'd19373, 16'd35363, 16'd3887, 16'd52656, 16'd13010, 16'd12064});
	test_expansion(128'h0710d473f4388a1aa91c7d6dbed848d9, {16'd59892, 16'd18017, 16'd52423, 16'd17330, 16'd5235, 16'd18686, 16'd3339, 16'd13357, 16'd57664, 16'd61883, 16'd3029, 16'd47656, 16'd43888, 16'd65079, 16'd44730, 16'd30312, 16'd18326, 16'd22299, 16'd48047, 16'd37371, 16'd51188, 16'd42363, 16'd64041, 16'd14258, 16'd62637, 16'd20330});
	test_expansion(128'hd1ef960a02db069e2326e5c2e176ea7b, {16'd41791, 16'd3920, 16'd26396, 16'd11730, 16'd731, 16'd21635, 16'd29538, 16'd11669, 16'd64795, 16'd17624, 16'd58569, 16'd47520, 16'd8772, 16'd1235, 16'd24644, 16'd57314, 16'd46685, 16'd55248, 16'd58678, 16'd54068, 16'd12359, 16'd32037, 16'd23019, 16'd21513, 16'd13178, 16'd45130});
	test_expansion(128'h300dc2b4f41ce869f20ba63fa99de1c8, {16'd46250, 16'd55974, 16'd38442, 16'd4690, 16'd45979, 16'd40274, 16'd33432, 16'd27487, 16'd15820, 16'd21710, 16'd27224, 16'd25640, 16'd52118, 16'd31568, 16'd22697, 16'd54295, 16'd18797, 16'd3222, 16'd18865, 16'd35606, 16'd29460, 16'd52982, 16'd19795, 16'd48335, 16'd51057, 16'd29740});
	test_expansion(128'hc2071bc14d8e2a449fa86bda81c87e90, {16'd8072, 16'd6642, 16'd29428, 16'd36781, 16'd36014, 16'd50836, 16'd36092, 16'd35424, 16'd46635, 16'd46732, 16'd27840, 16'd27106, 16'd45751, 16'd27762, 16'd51605, 16'd39510, 16'd28509, 16'd45956, 16'd14711, 16'd14873, 16'd45748, 16'd61848, 16'd62408, 16'd27150, 16'd3290, 16'd21767});
	test_expansion(128'h5633496c6722121f6de4202d1832ddf7, {16'd35365, 16'd873, 16'd40956, 16'd55026, 16'd14380, 16'd9612, 16'd54933, 16'd4536, 16'd215, 16'd44753, 16'd26313, 16'd18369, 16'd36105, 16'd5814, 16'd64423, 16'd8255, 16'd61491, 16'd5628, 16'd54374, 16'd31913, 16'd6150, 16'd25841, 16'd16213, 16'd29294, 16'd52133, 16'd17547});
	test_expansion(128'h6d177cb16b72c4d56ab6d4b04fe6d840, {16'd50007, 16'd15655, 16'd58305, 16'd37240, 16'd21389, 16'd57607, 16'd64431, 16'd34363, 16'd23781, 16'd11710, 16'd21082, 16'd2481, 16'd44304, 16'd29345, 16'd24551, 16'd15583, 16'd62710, 16'd4567, 16'd34114, 16'd36096, 16'd65194, 16'd13335, 16'd44930, 16'd47464, 16'd3086, 16'd1712});
	test_expansion(128'h7889f94daa1c7dd26df3a3d238949b93, {16'd43953, 16'd51307, 16'd43140, 16'd9398, 16'd2062, 16'd46851, 16'd62651, 16'd57932, 16'd2744, 16'd2879, 16'd53512, 16'd43514, 16'd54753, 16'd40793, 16'd61920, 16'd48603, 16'd9522, 16'd1544, 16'd41585, 16'd19661, 16'd10814, 16'd25203, 16'd13764, 16'd32386, 16'd34204, 16'd7288});
	test_expansion(128'h1e8d42ebfee3b8ba53d088a4e082ad0b, {16'd56945, 16'd3787, 16'd39723, 16'd52358, 16'd25196, 16'd4467, 16'd12009, 16'd8275, 16'd42305, 16'd21068, 16'd51457, 16'd38689, 16'd6644, 16'd65368, 16'd43718, 16'd10615, 16'd42971, 16'd28092, 16'd58534, 16'd464, 16'd55997, 16'd19212, 16'd31286, 16'd41993, 16'd6040, 16'd47675});
	test_expansion(128'h6b39b624a40d28becfea54794fe8fffb, {16'd41272, 16'd12088, 16'd36479, 16'd17282, 16'd14264, 16'd38887, 16'd63587, 16'd50728, 16'd1783, 16'd63080, 16'd27864, 16'd40921, 16'd65291, 16'd35029, 16'd38135, 16'd16949, 16'd53322, 16'd13917, 16'd49591, 16'd7507, 16'd30359, 16'd18743, 16'd8740, 16'd57545, 16'd45793, 16'd6670});
	test_expansion(128'h8387c26850dc7733a3fb89a3c63494f9, {16'd23763, 16'd63791, 16'd1063, 16'd15579, 16'd38586, 16'd47442, 16'd42222, 16'd32189, 16'd550, 16'd19813, 16'd32900, 16'd22943, 16'd62739, 16'd65019, 16'd22324, 16'd26136, 16'd30513, 16'd23838, 16'd9411, 16'd3324, 16'd16425, 16'd48206, 16'd24790, 16'd58006, 16'd12336, 16'd12512});
	test_expansion(128'hd0c5d0b9ebdeb3c373c3ebc944e6c13a, {16'd60365, 16'd50159, 16'd35480, 16'd7495, 16'd29351, 16'd30485, 16'd20073, 16'd12853, 16'd44030, 16'd2236, 16'd6343, 16'd58900, 16'd25399, 16'd30154, 16'd23860, 16'd49795, 16'd4556, 16'd54805, 16'd39446, 16'd32872, 16'd14747, 16'd6893, 16'd27788, 16'd64475, 16'd8033, 16'd51241});
	test_expansion(128'h4fdedaee82982e130fab8213532ae0ee, {16'd14956, 16'd45457, 16'd27825, 16'd41901, 16'd15936, 16'd59226, 16'd63948, 16'd24563, 16'd25932, 16'd8360, 16'd49168, 16'd33986, 16'd32374, 16'd51263, 16'd39171, 16'd4428, 16'd43786, 16'd14141, 16'd61739, 16'd16518, 16'd56908, 16'd10952, 16'd54946, 16'd32622, 16'd57879, 16'd23621});
	test_expansion(128'hfc65898d137be654d74a346dfbab90c4, {16'd42475, 16'd23918, 16'd42584, 16'd55260, 16'd7143, 16'd54862, 16'd22697, 16'd9051, 16'd13016, 16'd34723, 16'd60220, 16'd43563, 16'd41435, 16'd39967, 16'd53485, 16'd51872, 16'd49234, 16'd6169, 16'd55061, 16'd3490, 16'd6235, 16'd24951, 16'd41133, 16'd38280, 16'd36095, 16'd60489});
	test_expansion(128'hd5d4213efd7ab26f2e9d0466384d58de, {16'd15412, 16'd39758, 16'd19818, 16'd36599, 16'd11117, 16'd22979, 16'd8328, 16'd37093, 16'd42311, 16'd13938, 16'd27534, 16'd27213, 16'd39123, 16'd198, 16'd38093, 16'd5263, 16'd50471, 16'd45868, 16'd9748, 16'd50122, 16'd29684, 16'd9991, 16'd32601, 16'd56218, 16'd13362, 16'd34299});
	test_expansion(128'hd13aa5378a190bfdb14c7562d936fdf9, {16'd21933, 16'd27107, 16'd51576, 16'd39540, 16'd61610, 16'd14609, 16'd3575, 16'd40616, 16'd22640, 16'd56063, 16'd21831, 16'd118, 16'd36170, 16'd17668, 16'd20651, 16'd58742, 16'd59168, 16'd1585, 16'd436, 16'd13945, 16'd24558, 16'd39396, 16'd46666, 16'd56679, 16'd21545, 16'd21903});
	test_expansion(128'h99589603779b0872bf1b0154a621bc4c, {16'd53909, 16'd61179, 16'd30046, 16'd8167, 16'd38002, 16'd36145, 16'd52520, 16'd33259, 16'd9442, 16'd32745, 16'd6927, 16'd54056, 16'd11495, 16'd59610, 16'd60599, 16'd18783, 16'd64170, 16'd50313, 16'd40150, 16'd32704, 16'd23091, 16'd38856, 16'd19357, 16'd4802, 16'd64156, 16'd6959});
	test_expansion(128'h006cc7abbbb3cdc5612ad94d9e1ad26a, {16'd24395, 16'd24002, 16'd44816, 16'd38139, 16'd7330, 16'd35551, 16'd53275, 16'd58955, 16'd18124, 16'd43410, 16'd41142, 16'd55578, 16'd16809, 16'd49242, 16'd37177, 16'd20340, 16'd24279, 16'd56689, 16'd29790, 16'd17958, 16'd2362, 16'd47454, 16'd14153, 16'd18620, 16'd17346, 16'd10972});
	test_expansion(128'h12eeab244b4fa5a6b765d25bc7da8559, {16'd17109, 16'd29703, 16'd15656, 16'd12685, 16'd31005, 16'd11833, 16'd18621, 16'd28051, 16'd37680, 16'd56994, 16'd31801, 16'd24637, 16'd32264, 16'd14948, 16'd61740, 16'd30047, 16'd14596, 16'd46095, 16'd32796, 16'd46656, 16'd289, 16'd63554, 16'd31172, 16'd11872, 16'd31012, 16'd51493});
	test_expansion(128'hf7444d718f0f4ada8aa9b32a3569ae2b, {16'd41124, 16'd59945, 16'd48152, 16'd3670, 16'd31525, 16'd10637, 16'd244, 16'd59010, 16'd30746, 16'd21215, 16'd58549, 16'd5542, 16'd26882, 16'd2097, 16'd18256, 16'd1204, 16'd51569, 16'd6351, 16'd54990, 16'd17454, 16'd26068, 16'd18393, 16'd29047, 16'd40104, 16'd59734, 16'd47144});
	test_expansion(128'h769e0fbc97e1d93dec122c0cb422a3ac, {16'd5185, 16'd51443, 16'd65251, 16'd31977, 16'd39370, 16'd54725, 16'd60602, 16'd52108, 16'd13574, 16'd3396, 16'd32148, 16'd42817, 16'd1742, 16'd10439, 16'd62542, 16'd47425, 16'd37602, 16'd11468, 16'd64486, 16'd7082, 16'd62336, 16'd65246, 16'd13266, 16'd58058, 16'd3787, 16'd8213});
	test_expansion(128'hc29f976a5b197dba25d5ac770309cf5f, {16'd61057, 16'd31655, 16'd3658, 16'd61667, 16'd42791, 16'd19353, 16'd37663, 16'd40300, 16'd15855, 16'd51164, 16'd27823, 16'd29197, 16'd31019, 16'd25935, 16'd57364, 16'd53311, 16'd33535, 16'd10361, 16'd44572, 16'd4323, 16'd43045, 16'd36327, 16'd27010, 16'd21684, 16'd54347, 16'd58851});
	test_expansion(128'h490db2c179dbe0773a26ac45e752709e, {16'd30895, 16'd46518, 16'd3456, 16'd8391, 16'd38894, 16'd4729, 16'd41527, 16'd65243, 16'd47692, 16'd13150, 16'd45909, 16'd28364, 16'd56970, 16'd52962, 16'd51816, 16'd54004, 16'd7715, 16'd59927, 16'd61772, 16'd39800, 16'd60350, 16'd60212, 16'd45624, 16'd5825, 16'd27546, 16'd63236});
	test_expansion(128'h704004d6f82a585949cadcb58561befc, {16'd17227, 16'd63142, 16'd30032, 16'd49668, 16'd44179, 16'd24843, 16'd36784, 16'd27161, 16'd55730, 16'd17599, 16'd374, 16'd14674, 16'd32372, 16'd41966, 16'd18257, 16'd33048, 16'd53533, 16'd61455, 16'd30677, 16'd20890, 16'd26136, 16'd38821, 16'd43, 16'd5962, 16'd11767, 16'd8929});
	test_expansion(128'h8dae326d05e5fbfda75e308754704f88, {16'd16015, 16'd4533, 16'd33810, 16'd15150, 16'd8950, 16'd42595, 16'd10537, 16'd63054, 16'd17500, 16'd55516, 16'd55259, 16'd25985, 16'd10650, 16'd11601, 16'd49663, 16'd5879, 16'd6897, 16'd5782, 16'd21153, 16'd58187, 16'd14883, 16'd21600, 16'd55257, 16'd15331, 16'd52133, 16'd57627});
	test_expansion(128'ha5caaad58534fbb3eee11d5963e08f10, {16'd54834, 16'd58605, 16'd60237, 16'd53261, 16'd2078, 16'd25612, 16'd9899, 16'd29513, 16'd31903, 16'd18818, 16'd31441, 16'd38487, 16'd46070, 16'd51808, 16'd1673, 16'd42170, 16'd54288, 16'd22539, 16'd59224, 16'd35891, 16'd5676, 16'd44627, 16'd63018, 16'd46517, 16'd163, 16'd25040});
	test_expansion(128'h5c46146f6056dbd3b58cc45b0a5f6e1a, {16'd8778, 16'd48918, 16'd33664, 16'd44219, 16'd26169, 16'd58138, 16'd6748, 16'd62434, 16'd19825, 16'd61668, 16'd48375, 16'd55008, 16'd61499, 16'd50165, 16'd40862, 16'd1745, 16'd56540, 16'd30825, 16'd17797, 16'd17273, 16'd25133, 16'd40633, 16'd39829, 16'd33563, 16'd17429, 16'd6467});
	test_expansion(128'hebf48b08cb3a250084324f3c34be7df5, {16'd21554, 16'd51432, 16'd41591, 16'd63349, 16'd42143, 16'd43375, 16'd60669, 16'd28293, 16'd938, 16'd21177, 16'd27377, 16'd863, 16'd4025, 16'd34181, 16'd43349, 16'd7163, 16'd46473, 16'd50699, 16'd11429, 16'd26913, 16'd37836, 16'd4512, 16'd7026, 16'd36038, 16'd44500, 16'd64289});
	test_expansion(128'hcb151c03e86c5cf95ff0a434a0d1803f, {16'd40896, 16'd42118, 16'd54468, 16'd39799, 16'd12756, 16'd47856, 16'd37030, 16'd20376, 16'd45153, 16'd26535, 16'd52370, 16'd12457, 16'd38108, 16'd13762, 16'd51564, 16'd29994, 16'd21016, 16'd52326, 16'd26023, 16'd65218, 16'd21867, 16'd10494, 16'd1363, 16'd45954, 16'd661, 16'd64733});
	test_expansion(128'h2f21b58a033c3ad8ad7304c73ef47dc2, {16'd27895, 16'd2492, 16'd22756, 16'd44832, 16'd20638, 16'd51962, 16'd24642, 16'd49026, 16'd22853, 16'd64746, 16'd30117, 16'd54231, 16'd24298, 16'd56764, 16'd14053, 16'd51979, 16'd8569, 16'd40663, 16'd30578, 16'd57505, 16'd106, 16'd491, 16'd37248, 16'd7167, 16'd58268, 16'd13938});
	test_expansion(128'h9dfafca86e32d9a0dcd12c4f70397054, {16'd4379, 16'd37666, 16'd35963, 16'd4510, 16'd57808, 16'd4553, 16'd47671, 16'd12578, 16'd50192, 16'd7247, 16'd485, 16'd24479, 16'd7575, 16'd48398, 16'd24693, 16'd30207, 16'd47563, 16'd14122, 16'd28227, 16'd4634, 16'd40849, 16'd31282, 16'd3533, 16'd43679, 16'd47398, 16'd48669});
	test_expansion(128'h245b9782d1fba55c70632c49dbc2183f, {16'd60666, 16'd1046, 16'd16505, 16'd384, 16'd10339, 16'd2651, 16'd22611, 16'd12691, 16'd720, 16'd20801, 16'd10321, 16'd64914, 16'd9288, 16'd31860, 16'd784, 16'd45514, 16'd61773, 16'd2748, 16'd44455, 16'd42128, 16'd48975, 16'd15286, 16'd28517, 16'd23894, 16'd63519, 16'd15851});
	test_expansion(128'ha269401ea95b61105345730dc1c685de, {16'd11516, 16'd50598, 16'd28415, 16'd64960, 16'd61973, 16'd46110, 16'd55994, 16'd12331, 16'd1742, 16'd99, 16'd63658, 16'd63534, 16'd32548, 16'd18525, 16'd43192, 16'd63127, 16'd58254, 16'd55393, 16'd17682, 16'd57076, 16'd9810, 16'd21043, 16'd4062, 16'd59525, 16'd32855, 16'd3616});
	test_expansion(128'h961f004458f8cbb68c84a20a9e6ac66d, {16'd34644, 16'd6249, 16'd32463, 16'd28309, 16'd49158, 16'd21147, 16'd23566, 16'd20032, 16'd57760, 16'd57841, 16'd18686, 16'd55778, 16'd61328, 16'd11937, 16'd36761, 16'd6876, 16'd63936, 16'd5633, 16'd2346, 16'd10125, 16'd60234, 16'd15333, 16'd17283, 16'd22015, 16'd56079, 16'd26807});
	test_expansion(128'h80a873fd4af8515fcbc2895ec839da39, {16'd29969, 16'd57157, 16'd31719, 16'd49873, 16'd32899, 16'd8264, 16'd18807, 16'd50123, 16'd31771, 16'd23578, 16'd61379, 16'd1188, 16'd99, 16'd59486, 16'd19109, 16'd63661, 16'd18014, 16'd44627, 16'd2643, 16'd44541, 16'd64717, 16'd17752, 16'd34239, 16'd10783, 16'd7513, 16'd21880});
	test_expansion(128'hb2b3c65e3aa96c90c60bbdfcb4467696, {16'd54774, 16'd10560, 16'd49919, 16'd36133, 16'd11952, 16'd20486, 16'd13812, 16'd62240, 16'd35129, 16'd44650, 16'd51139, 16'd52068, 16'd33671, 16'd42111, 16'd44006, 16'd18661, 16'd33863, 16'd27992, 16'd35072, 16'd6483, 16'd49045, 16'd16860, 16'd62993, 16'd8582, 16'd64444, 16'd11667});
	test_expansion(128'h02f48d020cb9ea394b86ba5ca1ce1e31, {16'd61958, 16'd56894, 16'd45917, 16'd33012, 16'd53569, 16'd51507, 16'd3286, 16'd31264, 16'd22185, 16'd16119, 16'd53477, 16'd52985, 16'd19245, 16'd30473, 16'd2553, 16'd1053, 16'd12689, 16'd11869, 16'd20989, 16'd61778, 16'd54596, 16'd22486, 16'd64882, 16'd54075, 16'd30588, 16'd461});
	test_expansion(128'h56fd69546a377ec99505a7265dc0c887, {16'd33473, 16'd34877, 16'd58863, 16'd57605, 16'd46418, 16'd8501, 16'd49579, 16'd7622, 16'd27442, 16'd14903, 16'd20001, 16'd15154, 16'd42841, 16'd17474, 16'd48630, 16'd22186, 16'd62138, 16'd15096, 16'd60432, 16'd9255, 16'd21230, 16'd43438, 16'd3464, 16'd54447, 16'd2922, 16'd63379});
	test_expansion(128'h206569080a125d63eba7dd50dfa5e1ee, {16'd42535, 16'd30109, 16'd13097, 16'd50463, 16'd24385, 16'd41931, 16'd44242, 16'd34694, 16'd61133, 16'd50352, 16'd62486, 16'd46689, 16'd54916, 16'd5011, 16'd12627, 16'd4025, 16'd42686, 16'd8748, 16'd40045, 16'd36831, 16'd39973, 16'd12686, 16'd2484, 16'd58250, 16'd1542, 16'd56205});
	test_expansion(128'hd87ac283e9e37a53914a558887e61e19, {16'd7826, 16'd19863, 16'd22305, 16'd13460, 16'd26010, 16'd29796, 16'd50664, 16'd45709, 16'd10146, 16'd30993, 16'd51450, 16'd20537, 16'd13810, 16'd46598, 16'd15539, 16'd39395, 16'd13224, 16'd24080, 16'd28206, 16'd48174, 16'd64382, 16'd51589, 16'd17211, 16'd2251, 16'd28821, 16'd63443});
	test_expansion(128'h6c44916cb82d42c25dcc94971968a54a, {16'd56669, 16'd4211, 16'd54789, 16'd6336, 16'd41637, 16'd62390, 16'd6054, 16'd32802, 16'd44928, 16'd26651, 16'd38809, 16'd24359, 16'd54922, 16'd47644, 16'd60304, 16'd12321, 16'd5374, 16'd5434, 16'd30812, 16'd31328, 16'd39955, 16'd9213, 16'd27636, 16'd63618, 16'd37314, 16'd9888});
	test_expansion(128'h791d2e415be10db21f5f0f0f7d1545e0, {16'd13187, 16'd13358, 16'd70, 16'd21597, 16'd40804, 16'd45099, 16'd4309, 16'd40303, 16'd42436, 16'd15817, 16'd37448, 16'd26274, 16'd46489, 16'd18816, 16'd58488, 16'd22975, 16'd35620, 16'd59472, 16'd4668, 16'd12009, 16'd19795, 16'd23018, 16'd35176, 16'd9686, 16'd20344, 16'd46982});
	test_expansion(128'h391d89e3ac39feb27ce7c6876ef31f8b, {16'd32482, 16'd7143, 16'd50271, 16'd12684, 16'd59602, 16'd58169, 16'd35598, 16'd47867, 16'd10519, 16'd58625, 16'd59841, 16'd40335, 16'd39033, 16'd20108, 16'd43298, 16'd8701, 16'd33023, 16'd18152, 16'd12509, 16'd20289, 16'd33169, 16'd3955, 16'd60748, 16'd7387, 16'd60701, 16'd43008});
	test_expansion(128'h9771baec6a877a670c1448b0cd500a08, {16'd62647, 16'd7685, 16'd61600, 16'd7295, 16'd38531, 16'd6475, 16'd61490, 16'd62106, 16'd55408, 16'd13963, 16'd17318, 16'd59365, 16'd23504, 16'd50916, 16'd35328, 16'd39472, 16'd40290, 16'd30582, 16'd25719, 16'd62626, 16'd62164, 16'd7431, 16'd22862, 16'd17539, 16'd26689, 16'd47785});
	test_expansion(128'hf6921ce43c748ca8ace4f79dd33058e6, {16'd28050, 16'd24473, 16'd15928, 16'd50796, 16'd8706, 16'd45754, 16'd24983, 16'd63255, 16'd61781, 16'd63842, 16'd23733, 16'd64753, 16'd23370, 16'd19632, 16'd48823, 16'd54531, 16'd63888, 16'd7397, 16'd19803, 16'd60499, 16'd30368, 16'd23894, 16'd36636, 16'd30321, 16'd24900, 16'd18863});
	test_expansion(128'hb108c958a190cc7b620661c3fb0383da, {16'd36095, 16'd55448, 16'd64071, 16'd42093, 16'd23214, 16'd28266, 16'd17661, 16'd1144, 16'd52788, 16'd17444, 16'd55356, 16'd50198, 16'd59927, 16'd1861, 16'd17416, 16'd5486, 16'd10198, 16'd24931, 16'd24534, 16'd65319, 16'd64676, 16'd53353, 16'd24180, 16'd43672, 16'd26309, 16'd23574});
	test_expansion(128'h39a65a034bf565f028c48086008d0716, {16'd53032, 16'd56301, 16'd44070, 16'd56217, 16'd20096, 16'd59420, 16'd58848, 16'd13327, 16'd2892, 16'd34067, 16'd8842, 16'd5686, 16'd34031, 16'd3817, 16'd57119, 16'd14334, 16'd22895, 16'd38785, 16'd39346, 16'd20832, 16'd65113, 16'd34751, 16'd42263, 16'd40964, 16'd34135, 16'd14006});
	test_expansion(128'had9e8b8292f8935a4f3c0a694e38fb7d, {16'd43901, 16'd52421, 16'd29164, 16'd55846, 16'd34961, 16'd62656, 16'd63401, 16'd53393, 16'd14578, 16'd30514, 16'd38259, 16'd6003, 16'd48582, 16'd12482, 16'd35065, 16'd22008, 16'd46708, 16'd39892, 16'd5477, 16'd11376, 16'd6552, 16'd50885, 16'd12320, 16'd21176, 16'd15382, 16'd4290});
	test_expansion(128'heb50a8de680fb157f5d3e819149bf8c3, {16'd37417, 16'd747, 16'd53423, 16'd63839, 16'd52439, 16'd26908, 16'd20644, 16'd5447, 16'd36772, 16'd23328, 16'd54589, 16'd5044, 16'd32819, 16'd18388, 16'd56546, 16'd10821, 16'd20032, 16'd17459, 16'd58861, 16'd45385, 16'd51616, 16'd4442, 16'd42451, 16'd55250, 16'd25159, 16'd7753});
	test_expansion(128'hdc05f0556936a6c4ab6d91dd341cbeb3, {16'd39060, 16'd26763, 16'd34058, 16'd30961, 16'd19689, 16'd52334, 16'd37334, 16'd36669, 16'd52434, 16'd51727, 16'd39963, 16'd42226, 16'd20255, 16'd51439, 16'd57824, 16'd57683, 16'd29725, 16'd31403, 16'd27026, 16'd49881, 16'd61466, 16'd36409, 16'd20208, 16'd53163, 16'd21434, 16'd64574});
	test_expansion(128'h43fc10d0fc6fe024fe213fb23ca36954, {16'd10746, 16'd6206, 16'd61855, 16'd6960, 16'd40319, 16'd14620, 16'd10621, 16'd55489, 16'd33312, 16'd11390, 16'd18053, 16'd56543, 16'd10223, 16'd9494, 16'd52852, 16'd20623, 16'd55613, 16'd52836, 16'd40451, 16'd6378, 16'd28948, 16'd27914, 16'd55094, 16'd7683, 16'd52511, 16'd22872});
	test_expansion(128'h3d42edf3830d785fe34b7794ab700ea0, {16'd11416, 16'd60109, 16'd53873, 16'd45447, 16'd54619, 16'd42802, 16'd49497, 16'd39907, 16'd18301, 16'd5099, 16'd20009, 16'd55011, 16'd17456, 16'd30671, 16'd57040, 16'd17748, 16'd31825, 16'd15041, 16'd54400, 16'd10522, 16'd18707, 16'd12497, 16'd30102, 16'd43301, 16'd59529, 16'd5180});
	test_expansion(128'h636a76f45f29d5cff0e314ca47982de0, {16'd27065, 16'd32702, 16'd44534, 16'd59072, 16'd12341, 16'd5482, 16'd50011, 16'd18582, 16'd4340, 16'd58599, 16'd30569, 16'd17367, 16'd61678, 16'd27389, 16'd21824, 16'd22152, 16'd33974, 16'd29, 16'd40099, 16'd34258, 16'd3723, 16'd2569, 16'd2215, 16'd63730, 16'd485, 16'd7623});
	test_expansion(128'he7fbb55c4c994e26b9d80ae662b5e736, {16'd55066, 16'd63914, 16'd61757, 16'd60272, 16'd56850, 16'd37330, 16'd16932, 16'd64039, 16'd61614, 16'd51196, 16'd26599, 16'd7405, 16'd44438, 16'd7553, 16'd41534, 16'd35760, 16'd12313, 16'd59984, 16'd15057, 16'd6852, 16'd55187, 16'd55354, 16'd23477, 16'd33174, 16'd44054, 16'd60462});
	test_expansion(128'hb15803d90382a334005e60560a6264f8, {16'd34567, 16'd12556, 16'd44209, 16'd3996, 16'd16930, 16'd11718, 16'd60295, 16'd31413, 16'd9815, 16'd40779, 16'd22946, 16'd36179, 16'd24550, 16'd22156, 16'd20204, 16'd29885, 16'd8187, 16'd28495, 16'd34801, 16'd65110, 16'd43032, 16'd42032, 16'd5792, 16'd31608, 16'd4, 16'd9134});
	test_expansion(128'h3b9b2ca179fc9e21b228cce31b6fd244, {16'd5658, 16'd35634, 16'd16083, 16'd53468, 16'd32559, 16'd30447, 16'd17315, 16'd27922, 16'd37494, 16'd3579, 16'd45546, 16'd40245, 16'd39189, 16'd47833, 16'd22077, 16'd41416, 16'd28432, 16'd2730, 16'd35238, 16'd14873, 16'd12261, 16'd24627, 16'd65434, 16'd46087, 16'd47139, 16'd23912});
	test_expansion(128'h2b5b2692581f26cb7b4ff05eb04d2902, {16'd61592, 16'd53930, 16'd22532, 16'd21356, 16'd12456, 16'd5015, 16'd50955, 16'd48435, 16'd57510, 16'd28864, 16'd2756, 16'd186, 16'd15076, 16'd62592, 16'd50619, 16'd16797, 16'd15374, 16'd15487, 16'd3206, 16'd23410, 16'd28631, 16'd57700, 16'd10243, 16'd38612, 16'd36309, 16'd8769});
	test_expansion(128'hcfe2b5873a7a29f665fefd3d486c6883, {16'd37780, 16'd38896, 16'd822, 16'd61366, 16'd2712, 16'd11279, 16'd5308, 16'd60886, 16'd30596, 16'd35932, 16'd29646, 16'd40356, 16'd41754, 16'd64246, 16'd52786, 16'd39371, 16'd55719, 16'd65332, 16'd64132, 16'd62361, 16'd1368, 16'd62245, 16'd52262, 16'd56401, 16'd29806, 16'd2151});
	test_expansion(128'hb6610145ff5d2ce2da3d48453c26b9a9, {16'd14578, 16'd1417, 16'd30752, 16'd21828, 16'd33873, 16'd43216, 16'd64720, 16'd26600, 16'd54598, 16'd13777, 16'd53179, 16'd10968, 16'd604, 16'd64219, 16'd9605, 16'd28822, 16'd3726, 16'd12356, 16'd51772, 16'd45134, 16'd62779, 16'd41277, 16'd62113, 16'd48797, 16'd51471, 16'd46877});
	test_expansion(128'h4994240562f12eff443c787b0e5a0668, {16'd59988, 16'd23420, 16'd42279, 16'd22570, 16'd19732, 16'd22495, 16'd1576, 16'd58669, 16'd23920, 16'd59749, 16'd23327, 16'd52473, 16'd20898, 16'd47089, 16'd12294, 16'd61849, 16'd33169, 16'd21284, 16'd59471, 16'd42963, 16'd59626, 16'd16019, 16'd41529, 16'd45420, 16'd54117, 16'd39223});
	test_expansion(128'h57912732ae34839ce7e194220ea08e60, {16'd41653, 16'd46480, 16'd46817, 16'd25479, 16'd5792, 16'd51779, 16'd4486, 16'd1259, 16'd6826, 16'd55900, 16'd9086, 16'd48589, 16'd209, 16'd39302, 16'd45006, 16'd21429, 16'd35610, 16'd35628, 16'd56087, 16'd4051, 16'd62772, 16'd25749, 16'd16468, 16'd50284, 16'd30602, 16'd61024});
	test_expansion(128'hca887ea2fe6953891b034a4aa76c2ef8, {16'd64724, 16'd24018, 16'd872, 16'd27772, 16'd60082, 16'd34884, 16'd55064, 16'd31805, 16'd57968, 16'd38520, 16'd52540, 16'd61239, 16'd33321, 16'd11352, 16'd32976, 16'd24455, 16'd46997, 16'd32128, 16'd36244, 16'd8413, 16'd50583, 16'd6836, 16'd49236, 16'd36187, 16'd549, 16'd32005});
	test_expansion(128'h205d1eb8c5c2f4e8900ab7c57b1469dc, {16'd56080, 16'd51915, 16'd3922, 16'd59454, 16'd14510, 16'd60690, 16'd15357, 16'd14571, 16'd62539, 16'd35142, 16'd31845, 16'd14741, 16'd38717, 16'd26809, 16'd8660, 16'd53157, 16'd11957, 16'd11471, 16'd43524, 16'd19936, 16'd53349, 16'd14398, 16'd10359, 16'd45939, 16'd47966, 16'd3690});
	test_expansion(128'haec6be47eac56620b40e21b94fe8a6a6, {16'd22613, 16'd53737, 16'd15636, 16'd54538, 16'd22861, 16'd24186, 16'd10102, 16'd43209, 16'd29471, 16'd2395, 16'd5624, 16'd5209, 16'd47479, 16'd18527, 16'd27732, 16'd45346, 16'd20230, 16'd24159, 16'd23599, 16'd59609, 16'd47094, 16'd52207, 16'd50574, 16'd24957, 16'd14639, 16'd14041});
	test_expansion(128'h357983fdbcd3cad9400c4115b210ab1f, {16'd30199, 16'd24802, 16'd4729, 16'd11384, 16'd28628, 16'd39163, 16'd10808, 16'd17084, 16'd39629, 16'd56824, 16'd40590, 16'd9581, 16'd14538, 16'd59655, 16'd1604, 16'd48683, 16'd59684, 16'd63100, 16'd16746, 16'd1076, 16'd14109, 16'd15371, 16'd11536, 16'd22368, 16'd52360, 16'd11863});
	test_expansion(128'h2d8c19d007770e0dcfdef40fc666cb16, {16'd52274, 16'd30489, 16'd21284, 16'd15886, 16'd1353, 16'd45023, 16'd53979, 16'd3010, 16'd36278, 16'd11112, 16'd28691, 16'd42445, 16'd11059, 16'd55318, 16'd6913, 16'd63699, 16'd7298, 16'd12594, 16'd57227, 16'd60351, 16'd25332, 16'd60702, 16'd56205, 16'd55305, 16'd7644, 16'd30688});
	test_expansion(128'h27486c88f114cf2ebdc776fcd2c7bc43, {16'd65247, 16'd34152, 16'd2313, 16'd6523, 16'd24526, 16'd46929, 16'd19747, 16'd14156, 16'd9396, 16'd55741, 16'd61214, 16'd40569, 16'd23116, 16'd51135, 16'd5771, 16'd42497, 16'd15318, 16'd26092, 16'd32616, 16'd3815, 16'd3779, 16'd53271, 16'd44246, 16'd13300, 16'd42128, 16'd60391});
	test_expansion(128'h0dbe30864a277f77c2319e03b1f1547d, {16'd6044, 16'd45577, 16'd796, 16'd57814, 16'd4877, 16'd49196, 16'd8271, 16'd29391, 16'd28213, 16'd39890, 16'd21789, 16'd3572, 16'd55328, 16'd22777, 16'd20378, 16'd1009, 16'd14219, 16'd32075, 16'd8797, 16'd52117, 16'd18260, 16'd54059, 16'd51295, 16'd3906, 16'd41459, 16'd47146});
	test_expansion(128'h3bd9d5edaff0f9e09762774460c52f10, {16'd49254, 16'd4330, 16'd42874, 16'd24997, 16'd47728, 16'd16832, 16'd47887, 16'd53294, 16'd38769, 16'd49846, 16'd14957, 16'd44328, 16'd29603, 16'd56969, 16'd59943, 16'd24578, 16'd36968, 16'd20191, 16'd62494, 16'd22090, 16'd42113, 16'd53898, 16'd19708, 16'd17320, 16'd12639, 16'd43002});
	test_expansion(128'h30dfe08f87a592971a969d37e678a6fb, {16'd54844, 16'd6284, 16'd21535, 16'd50475, 16'd9548, 16'd54266, 16'd5121, 16'd20817, 16'd17052, 16'd12711, 16'd27887, 16'd53675, 16'd43820, 16'd15743, 16'd15848, 16'd49516, 16'd49375, 16'd44438, 16'd34374, 16'd50408, 16'd60777, 16'd47341, 16'd20602, 16'd23447, 16'd23419, 16'd58068});
	test_expansion(128'h171b58733f337194b9cae0751fec16d8, {16'd28765, 16'd59862, 16'd58021, 16'd45197, 16'd62215, 16'd29485, 16'd37910, 16'd55393, 16'd28590, 16'd24618, 16'd18703, 16'd29938, 16'd20618, 16'd46441, 16'd243, 16'd8422, 16'd37857, 16'd55750, 16'd60193, 16'd53299, 16'd60707, 16'd7348, 16'd42942, 16'd58572, 16'd57624, 16'd20638});
	test_expansion(128'hc349e0a0132cc98ea28b7612cc06f561, {16'd13304, 16'd14994, 16'd50431, 16'd11512, 16'd16928, 16'd35228, 16'd48, 16'd33526, 16'd63673, 16'd39689, 16'd28684, 16'd33065, 16'd1470, 16'd43020, 16'd27165, 16'd14876, 16'd20442, 16'd61591, 16'd10854, 16'd9906, 16'd37098, 16'd54764, 16'd37949, 16'd21343, 16'd45462, 16'd11483});
	test_expansion(128'h4a95decc4b000016068d497b9d8021b0, {16'd6931, 16'd62843, 16'd18803, 16'd20800, 16'd10122, 16'd57139, 16'd22562, 16'd49361, 16'd39249, 16'd3470, 16'd45852, 16'd62713, 16'd39262, 16'd12377, 16'd30524, 16'd17890, 16'd34185, 16'd36249, 16'd60604, 16'd33092, 16'd4327, 16'd11881, 16'd19363, 16'd3441, 16'd1800, 16'd51524});
	test_expansion(128'hbcf179be055dbb4497d07f5741a4cfa9, {16'd7591, 16'd12809, 16'd26471, 16'd53037, 16'd3175, 16'd45729, 16'd50599, 16'd55583, 16'd56474, 16'd28474, 16'd33508, 16'd47898, 16'd30470, 16'd7106, 16'd57718, 16'd61567, 16'd42156, 16'd28334, 16'd51454, 16'd3306, 16'd31537, 16'd45441, 16'd422, 16'd29012, 16'd41836, 16'd12016});
	test_expansion(128'hdd37b0d47bd49728e30c7e10c43d825c, {16'd49159, 16'd12605, 16'd38957, 16'd10907, 16'd56216, 16'd48685, 16'd36018, 16'd61979, 16'd27755, 16'd65267, 16'd38765, 16'd35928, 16'd7232, 16'd50723, 16'd40391, 16'd52724, 16'd30280, 16'd9365, 16'd27974, 16'd10923, 16'd59577, 16'd48850, 16'd62795, 16'd28342, 16'd59118, 16'd44717});
	test_expansion(128'h84336c8fb09dbfc4b98bab746963a548, {16'd64115, 16'd56269, 16'd38374, 16'd11298, 16'd40755, 16'd28898, 16'd36658, 16'd10786, 16'd19237, 16'd5557, 16'd55225, 16'd33060, 16'd35554, 16'd4116, 16'd45288, 16'd55934, 16'd37836, 16'd2866, 16'd22217, 16'd26561, 16'd32852, 16'd56990, 16'd60752, 16'd42033, 16'd41442, 16'd47274});
	test_expansion(128'hdca63c68bdc40d5971adfc58df662856, {16'd62999, 16'd20014, 16'd26127, 16'd24846, 16'd8921, 16'd39556, 16'd12107, 16'd42012, 16'd30168, 16'd25508, 16'd15224, 16'd9508, 16'd38434, 16'd33860, 16'd26756, 16'd41690, 16'd40828, 16'd17239, 16'd28816, 16'd8595, 16'd1393, 16'd7383, 16'd2439, 16'd36163, 16'd38347, 16'd17940});
	test_expansion(128'h631c8419a902a8dcf6698e8963a27763, {16'd30390, 16'd54623, 16'd48101, 16'd53894, 16'd16620, 16'd38323, 16'd37453, 16'd30312, 16'd56828, 16'd17236, 16'd38671, 16'd38298, 16'd8088, 16'd51470, 16'd26542, 16'd43647, 16'd12984, 16'd12156, 16'd39275, 16'd32970, 16'd2631, 16'd50698, 16'd49516, 16'd48655, 16'd49556, 16'd48302});
	test_expansion(128'hdf0e9cc1c49bfc83a0e6538d26193e9f, {16'd44028, 16'd58230, 16'd33966, 16'd18553, 16'd50338, 16'd34446, 16'd52704, 16'd8701, 16'd32098, 16'd14644, 16'd63784, 16'd40174, 16'd31997, 16'd22867, 16'd45274, 16'd4964, 16'd5418, 16'd42034, 16'd34075, 16'd48197, 16'd41324, 16'd35098, 16'd53800, 16'd57790, 16'd25016, 16'd45182});
	test_expansion(128'hab8f0017ba18989f2a822f68bf97ca2a, {16'd21044, 16'd60262, 16'd15829, 16'd58532, 16'd54649, 16'd37493, 16'd62096, 16'd49586, 16'd61168, 16'd20844, 16'd34663, 16'd18520, 16'd57610, 16'd54609, 16'd20374, 16'd31206, 16'd47160, 16'd16444, 16'd46381, 16'd41936, 16'd52124, 16'd17851, 16'd16051, 16'd46249, 16'd19561, 16'd18461});
	test_expansion(128'h0d935b8677107cdb1d4ac0aa28157bd9, {16'd60969, 16'd56026, 16'd53097, 16'd20563, 16'd59614, 16'd23669, 16'd53220, 16'd48617, 16'd22441, 16'd45017, 16'd32003, 16'd52585, 16'd33788, 16'd56982, 16'd5996, 16'd17224, 16'd63200, 16'd5491, 16'd14790, 16'd28305, 16'd9724, 16'd19573, 16'd11883, 16'd50426, 16'd51462, 16'd25244});
	test_expansion(128'ha8c4205f459c2020fd140b8773c74c5e, {16'd33502, 16'd3413, 16'd32938, 16'd53549, 16'd56970, 16'd20410, 16'd37098, 16'd40468, 16'd33407, 16'd60684, 16'd39243, 16'd38485, 16'd18217, 16'd41726, 16'd2285, 16'd28931, 16'd41188, 16'd21596, 16'd39111, 16'd1421, 16'd17897, 16'd55175, 16'd26336, 16'd19750, 16'd35168, 16'd7360});
	test_expansion(128'hf81108d8aa5e2794d2f8260741aaa0ba, {16'd48705, 16'd6290, 16'd19357, 16'd21967, 16'd25995, 16'd1295, 16'd15466, 16'd15045, 16'd46003, 16'd28673, 16'd56052, 16'd35732, 16'd41030, 16'd4399, 16'd17398, 16'd8637, 16'd11592, 16'd52100, 16'd59497, 16'd56835, 16'd49447, 16'd43005, 16'd44318, 16'd10582, 16'd3343, 16'd59908});
	test_expansion(128'h7f26732382d9b7031e5a19dddaecf7f1, {16'd17413, 16'd62228, 16'd28338, 16'd58974, 16'd30699, 16'd41454, 16'd1036, 16'd21509, 16'd54360, 16'd59029, 16'd47589, 16'd59688, 16'd23484, 16'd40230, 16'd50051, 16'd61330, 16'd28674, 16'd31595, 16'd26534, 16'd21155, 16'd47358, 16'd26797, 16'd34314, 16'd8516, 16'd54186, 16'd54930});
	test_expansion(128'hfc798871d0fdb68e301c445df6bf0724, {16'd14268, 16'd17426, 16'd21358, 16'd22236, 16'd233, 16'd28815, 16'd64902, 16'd27281, 16'd52967, 16'd9645, 16'd29380, 16'd29085, 16'd44392, 16'd62831, 16'd44976, 16'd9852, 16'd43518, 16'd13640, 16'd4546, 16'd42160, 16'd62645, 16'd39154, 16'd42183, 16'd15245, 16'd525, 16'd61048});
	test_expansion(128'he0c45c74f8018d868351f177f0fb642e, {16'd22580, 16'd6189, 16'd19105, 16'd41335, 16'd34265, 16'd56993, 16'd59796, 16'd60974, 16'd54228, 16'd31498, 16'd4904, 16'd38491, 16'd29075, 16'd59959, 16'd49547, 16'd65315, 16'd46817, 16'd6523, 16'd10653, 16'd38079, 16'd55081, 16'd24609, 16'd5784, 16'd63349, 16'd33805, 16'd3513});
	test_expansion(128'h9c07028152ab17b0fdd9744c4eb7679e, {16'd56616, 16'd15763, 16'd53157, 16'd17634, 16'd9128, 16'd35382, 16'd58712, 16'd13622, 16'd61811, 16'd50828, 16'd34218, 16'd14855, 16'd44328, 16'd54574, 16'd55360, 16'd38657, 16'd26408, 16'd10200, 16'd25046, 16'd6117, 16'd27460, 16'd30557, 16'd64271, 16'd10246, 16'd40548, 16'd31332});
	test_expansion(128'h9aa0f7c0d9ee45376e53fc8c2f2e5418, {16'd1165, 16'd63950, 16'd52327, 16'd39592, 16'd37467, 16'd13442, 16'd1458, 16'd22178, 16'd20187, 16'd33691, 16'd19287, 16'd48101, 16'd2426, 16'd34475, 16'd63663, 16'd51608, 16'd32424, 16'd46772, 16'd28998, 16'd35163, 16'd52162, 16'd26125, 16'd47313, 16'd22165, 16'd16720, 16'd29558});
	test_expansion(128'hc3269372df564f3b6319e09542d56cce, {16'd17027, 16'd50939, 16'd4104, 16'd14821, 16'd7956, 16'd21383, 16'd61317, 16'd49948, 16'd39537, 16'd33727, 16'd59093, 16'd59795, 16'd34204, 16'd54128, 16'd35683, 16'd59452, 16'd41326, 16'd45536, 16'd38452, 16'd39692, 16'd12120, 16'd42849, 16'd41490, 16'd26404, 16'd19515, 16'd4249});
	test_expansion(128'h0855723df2b6583ef49f33baf7926c1f, {16'd50845, 16'd29942, 16'd52407, 16'd63368, 16'd42223, 16'd47407, 16'd47536, 16'd2267, 16'd15827, 16'd23902, 16'd20669, 16'd61347, 16'd48764, 16'd10530, 16'd54591, 16'd89, 16'd36726, 16'd42774, 16'd21717, 16'd41291, 16'd47490, 16'd8934, 16'd18663, 16'd30480, 16'd1386, 16'd4282});
	test_expansion(128'hf1d47837ef15b4ef86656a6e1b8f9044, {16'd22681, 16'd35983, 16'd38220, 16'd29464, 16'd50262, 16'd46930, 16'd34409, 16'd49197, 16'd29888, 16'd54671, 16'd56387, 16'd51566, 16'd35325, 16'd2617, 16'd14178, 16'd24034, 16'd49448, 16'd64171, 16'd17177, 16'd28876, 16'd4655, 16'd52402, 16'd16621, 16'd7392, 16'd8471, 16'd62535});
	test_expansion(128'h82dd92cce8f8f984b09779a9ed065898, {16'd54145, 16'd37019, 16'd9195, 16'd18451, 16'd2699, 16'd63815, 16'd52202, 16'd22133, 16'd42303, 16'd20122, 16'd50944, 16'd7937, 16'd64706, 16'd25370, 16'd24336, 16'd58528, 16'd56735, 16'd19378, 16'd4300, 16'd25165, 16'd37192, 16'd16457, 16'd30601, 16'd50754, 16'd3925, 16'd6680});
	test_expansion(128'h1973f8e74d78ae7afe4aa3f04f40c4e1, {16'd51198, 16'd10510, 16'd2581, 16'd61403, 16'd34386, 16'd34514, 16'd16665, 16'd64103, 16'd13389, 16'd43385, 16'd26876, 16'd11790, 16'd49634, 16'd3316, 16'd57933, 16'd13612, 16'd27352, 16'd24438, 16'd18124, 16'd15128, 16'd21552, 16'd33363, 16'd2609, 16'd3807, 16'd10302, 16'd2089});
	test_expansion(128'h36413c72fccc9072502de6eed9407b3e, {16'd42671, 16'd31264, 16'd58434, 16'd43836, 16'd20867, 16'd59694, 16'd18048, 16'd22126, 16'd58149, 16'd30473, 16'd60512, 16'd21469, 16'd34714, 16'd59616, 16'd65294, 16'd27327, 16'd55252, 16'd32286, 16'd30113, 16'd15725, 16'd63319, 16'd34859, 16'd49215, 16'd1901, 16'd30013, 16'd8237});
	test_expansion(128'h6aa0348d7220fa726471741f8253dd69, {16'd1189, 16'd7847, 16'd33006, 16'd282, 16'd13141, 16'd41340, 16'd7933, 16'd54416, 16'd29161, 16'd36766, 16'd26316, 16'd29231, 16'd56590, 16'd58975, 16'd2724, 16'd56756, 16'd27230, 16'd50747, 16'd28269, 16'd599, 16'd605, 16'd6473, 16'd11574, 16'd48235, 16'd35471, 16'd7151});
	test_expansion(128'h5a87b5478b664f426a087a32f36c93a6, {16'd3396, 16'd49116, 16'd20844, 16'd61067, 16'd37962, 16'd15057, 16'd7806, 16'd41584, 16'd39837, 16'd54728, 16'd41233, 16'd40622, 16'd4513, 16'd29105, 16'd1223, 16'd45070, 16'd16745, 16'd59739, 16'd2533, 16'd29516, 16'd39098, 16'd60240, 16'd41874, 16'd13675, 16'd8247, 16'd16983});
	test_expansion(128'h7af148ffb810b17305385376370e9020, {16'd29459, 16'd39050, 16'd26793, 16'd9317, 16'd11599, 16'd5438, 16'd19654, 16'd25717, 16'd54838, 16'd8920, 16'd13760, 16'd18180, 16'd55521, 16'd55881, 16'd10199, 16'd45767, 16'd41036, 16'd50960, 16'd15362, 16'd7016, 16'd32785, 16'd62687, 16'd11965, 16'd38988, 16'd25427, 16'd45068});
	test_expansion(128'hbcedaa562a8fe713a653efe6ec0b2093, {16'd53660, 16'd13334, 16'd64031, 16'd47905, 16'd12402, 16'd9147, 16'd23042, 16'd48641, 16'd62355, 16'd61153, 16'd42667, 16'd16376, 16'd3876, 16'd19374, 16'd4850, 16'd38908, 16'd24911, 16'd29135, 16'd41745, 16'd21129, 16'd55142, 16'd62445, 16'd33266, 16'd14559, 16'd60579, 16'd62659});
	test_expansion(128'heb8d6f9f464ea97b77513649220fd6f6, {16'd23193, 16'd24867, 16'd31943, 16'd20875, 16'd43209, 16'd43605, 16'd11009, 16'd62309, 16'd58978, 16'd29019, 16'd32699, 16'd35868, 16'd45236, 16'd25108, 16'd43590, 16'd33677, 16'd54260, 16'd61027, 16'd45425, 16'd25645, 16'd18278, 16'd52521, 16'd35772, 16'd23260, 16'd10201, 16'd64484});
	test_expansion(128'h5f4613cdc2c03068a009dae0fc9fc930, {16'd40023, 16'd9602, 16'd44173, 16'd30045, 16'd55684, 16'd51860, 16'd28567, 16'd41305, 16'd4712, 16'd661, 16'd21089, 16'd20717, 16'd14307, 16'd30918, 16'd32392, 16'd58436, 16'd23431, 16'd36904, 16'd8419, 16'd19888, 16'd1972, 16'd63947, 16'd54203, 16'd3907, 16'd16165, 16'd7262});
	test_expansion(128'h79f6eb42a4ef8dcc983bdea063c8f433, {16'd54585, 16'd33043, 16'd26246, 16'd437, 16'd50668, 16'd61313, 16'd26243, 16'd64558, 16'd46846, 16'd35423, 16'd8357, 16'd82, 16'd27950, 16'd20207, 16'd30782, 16'd4511, 16'd8625, 16'd19236, 16'd59288, 16'd17086, 16'd40211, 16'd49884, 16'd24180, 16'd49828, 16'd9152, 16'd48315});
	test_expansion(128'h4ac8d0bc3081b1173ad978fdd011906a, {16'd48718, 16'd7756, 16'd5152, 16'd64652, 16'd12839, 16'd40623, 16'd43996, 16'd30606, 16'd44086, 16'd19036, 16'd28079, 16'd44321, 16'd45553, 16'd55225, 16'd29267, 16'd8274, 16'd25639, 16'd28965, 16'd63047, 16'd52266, 16'd58792, 16'd42616, 16'd39962, 16'd14065, 16'd18926, 16'd39398});
	test_expansion(128'h6790ecbaa63a58bf4909bfb372276851, {16'd30560, 16'd31028, 16'd12466, 16'd14940, 16'd343, 16'd32635, 16'd3298, 16'd22390, 16'd3981, 16'd17842, 16'd49320, 16'd27890, 16'd60379, 16'd31631, 16'd62325, 16'd17519, 16'd42424, 16'd18077, 16'd48549, 16'd19016, 16'd18502, 16'd16201, 16'd36315, 16'd32751, 16'd5135, 16'd24884});
	test_expansion(128'h49d22cc34c3f0d9631e55304520aa16a, {16'd46809, 16'd18803, 16'd37043, 16'd33051, 16'd15000, 16'd58064, 16'd51493, 16'd34257, 16'd63008, 16'd8659, 16'd9985, 16'd16684, 16'd15981, 16'd13003, 16'd62863, 16'd62009, 16'd31498, 16'd2620, 16'd39463, 16'd45679, 16'd34622, 16'd16375, 16'd6481, 16'd11883, 16'd25077, 16'd36956});
	test_expansion(128'h39c324c0e44f923d88b1c7c4eae39249, {16'd5819, 16'd47723, 16'd13213, 16'd28974, 16'd47720, 16'd4353, 16'd27623, 16'd45895, 16'd6499, 16'd49489, 16'd11082, 16'd56828, 16'd14330, 16'd20457, 16'd29268, 16'd60699, 16'd6261, 16'd12617, 16'd40509, 16'd49983, 16'd58376, 16'd57335, 16'd45273, 16'd13946, 16'd36763, 16'd22600});
	test_expansion(128'h853d78c6cc8465767ac62bcde37d86a6, {16'd16111, 16'd57023, 16'd50101, 16'd3568, 16'd23448, 16'd27223, 16'd20228, 16'd50378, 16'd11334, 16'd59631, 16'd28505, 16'd45691, 16'd3475, 16'd3842, 16'd60398, 16'd22534, 16'd57453, 16'd46780, 16'd48102, 16'd2519, 16'd28334, 16'd10971, 16'd11300, 16'd33446, 16'd19761, 16'd29580});
	test_expansion(128'h5fc8c8d5e0ffa8274f9baaa58ba20e52, {16'd41171, 16'd25711, 16'd652, 16'd35495, 16'd44363, 16'd42830, 16'd44441, 16'd43035, 16'd60291, 16'd11539, 16'd41764, 16'd7379, 16'd52946, 16'd1914, 16'd15161, 16'd52126, 16'd62705, 16'd47851, 16'd29611, 16'd31632, 16'd2988, 16'd19373, 16'd36083, 16'd52066, 16'd34261, 16'd17848});
	test_expansion(128'h205a485fec2c768e176873c49924c6b7, {16'd55452, 16'd43641, 16'd57033, 16'd27002, 16'd53266, 16'd40065, 16'd37947, 16'd47884, 16'd28681, 16'd15950, 16'd9343, 16'd17525, 16'd10566, 16'd50144, 16'd37888, 16'd8292, 16'd57578, 16'd38447, 16'd5507, 16'd488, 16'd22005, 16'd4789, 16'd2259, 16'd42194, 16'd1325, 16'd23965});
	test_expansion(128'ha2f075056827aefe890709463f240fd8, {16'd24951, 16'd33323, 16'd11176, 16'd39467, 16'd27762, 16'd20414, 16'd42010, 16'd15688, 16'd18796, 16'd56543, 16'd13567, 16'd9157, 16'd42765, 16'd42945, 16'd55603, 16'd55796, 16'd46102, 16'd40821, 16'd38420, 16'd4027, 16'd13642, 16'd3620, 16'd53805, 16'd61239, 16'd13045, 16'd8107});
	test_expansion(128'he458e89460850fbe5cd3ab2abf4cdb7e, {16'd54257, 16'd6818, 16'd63720, 16'd10606, 16'd23555, 16'd50702, 16'd62825, 16'd24081, 16'd40691, 16'd42261, 16'd12029, 16'd48900, 16'd12443, 16'd17943, 16'd47340, 16'd39002, 16'd29587, 16'd50966, 16'd17313, 16'd27396, 16'd17810, 16'd5720, 16'd35147, 16'd22387, 16'd27624, 16'd37247});
	test_expansion(128'h873ba7313e90db3dd87385eedc4fd2fb, {16'd34431, 16'd48282, 16'd3203, 16'd6758, 16'd34060, 16'd12362, 16'd8648, 16'd50353, 16'd47429, 16'd40405, 16'd15918, 16'd39283, 16'd51664, 16'd46250, 16'd1294, 16'd58080, 16'd16621, 16'd8896, 16'd8124, 16'd55698, 16'd22887, 16'd12963, 16'd24670, 16'd49962, 16'd7242, 16'd4873});
	test_expansion(128'hee8700d057d7778e220c2575a7152631, {16'd55953, 16'd49972, 16'd23936, 16'd46938, 16'd62538, 16'd4812, 16'd18010, 16'd12176, 16'd12147, 16'd42502, 16'd22588, 16'd41698, 16'd39760, 16'd10904, 16'd27086, 16'd19549, 16'd1021, 16'd1193, 16'd57700, 16'd24419, 16'd33474, 16'd34197, 16'd47290, 16'd17866, 16'd23997, 16'd9439});
	test_expansion(128'hb4a5c4ec3cde2d9f52f29b5e45fdc57e, {16'd50558, 16'd60639, 16'd64350, 16'd32810, 16'd42168, 16'd54669, 16'd30729, 16'd44691, 16'd9910, 16'd39640, 16'd52794, 16'd52475, 16'd58897, 16'd32391, 16'd39357, 16'd3814, 16'd45247, 16'd19887, 16'd38541, 16'd40232, 16'd58290, 16'd33314, 16'd25393, 16'd57260, 16'd16482, 16'd20881});
	test_expansion(128'h845c913f3aa5801cded14389aab1e496, {16'd50422, 16'd56201, 16'd28684, 16'd12762, 16'd3172, 16'd44758, 16'd33501, 16'd35564, 16'd12428, 16'd40416, 16'd62686, 16'd46475, 16'd1131, 16'd13765, 16'd13726, 16'd53896, 16'd19211, 16'd17598, 16'd34668, 16'd27350, 16'd20958, 16'd62986, 16'd9536, 16'd9824, 16'd51829, 16'd33976});
	test_expansion(128'he51ea4cc5b5d1d0bf1aafdb9df5fe15d, {16'd59645, 16'd9707, 16'd60293, 16'd60840, 16'd53242, 16'd35920, 16'd25447, 16'd14721, 16'd44494, 16'd60853, 16'd65148, 16'd32083, 16'd22733, 16'd34973, 16'd29561, 16'd26695, 16'd9066, 16'd7285, 16'd52454, 16'd63156, 16'd60012, 16'd30155, 16'd61579, 16'd58689, 16'd6958, 16'd51952});
	test_expansion(128'h15c3d812affb1c2ecdf6d1ec74d1c00b, {16'd5959, 16'd299, 16'd36125, 16'd40190, 16'd8228, 16'd13863, 16'd21866, 16'd55428, 16'd3010, 16'd1879, 16'd50415, 16'd37757, 16'd18715, 16'd51225, 16'd29697, 16'd1676, 16'd54346, 16'd30712, 16'd22617, 16'd17728, 16'd43648, 16'd23285, 16'd5321, 16'd23302, 16'd63770, 16'd50994});
	test_expansion(128'hd83cb9b6b5861897f982265af632524c, {16'd14939, 16'd3464, 16'd10001, 16'd13425, 16'd8843, 16'd53894, 16'd57562, 16'd52737, 16'd31324, 16'd33561, 16'd44134, 16'd4952, 16'd41092, 16'd53092, 16'd18978, 16'd7376, 16'd18635, 16'd24974, 16'd14285, 16'd4147, 16'd10386, 16'd50767, 16'd1684, 16'd36014, 16'd23903, 16'd34144});
	test_expansion(128'h585aa97e3fb3e64084c820e446f0f4d7, {16'd28556, 16'd35254, 16'd38042, 16'd18530, 16'd50058, 16'd12509, 16'd21128, 16'd17731, 16'd49441, 16'd26684, 16'd22088, 16'd63354, 16'd23251, 16'd27500, 16'd15490, 16'd33782, 16'd45223, 16'd7762, 16'd64367, 16'd19531, 16'd56809, 16'd29004, 16'd53898, 16'd37832, 16'd32499, 16'd33661});
	test_expansion(128'h6d68e2758d914831ae8b0c68a9d1a37c, {16'd39921, 16'd4943, 16'd2321, 16'd12301, 16'd26067, 16'd686, 16'd10711, 16'd10615, 16'd34304, 16'd12450, 16'd52975, 16'd1525, 16'd46520, 16'd45787, 16'd24895, 16'd40124, 16'd53287, 16'd3972, 16'd1900, 16'd24196, 16'd54129, 16'd62024, 16'd17145, 16'd18448, 16'd46077, 16'd35070});
	test_expansion(128'hf7f8b8950a5ba11374604c1c8a6b470f, {16'd64250, 16'd21910, 16'd28188, 16'd29890, 16'd22781, 16'd58087, 16'd56170, 16'd44760, 16'd63422, 16'd34032, 16'd32420, 16'd32433, 16'd24641, 16'd6094, 16'd50863, 16'd9139, 16'd34862, 16'd1453, 16'd13760, 16'd52734, 16'd56416, 16'd31884, 16'd22336, 16'd40306, 16'd62935, 16'd35570});
	test_expansion(128'h547dfa985003f650f0daa9304f5e5846, {16'd561, 16'd42381, 16'd3866, 16'd18173, 16'd57700, 16'd25151, 16'd61712, 16'd30288, 16'd60988, 16'd38602, 16'd37343, 16'd45165, 16'd58020, 16'd54204, 16'd21688, 16'd50458, 16'd60801, 16'd63051, 16'd3923, 16'd64371, 16'd17159, 16'd57766, 16'd36387, 16'd5551, 16'd54589, 16'd2373});
	test_expansion(128'h9c8c1caa71f6f860a55c7ad24de8433b, {16'd43320, 16'd64772, 16'd33424, 16'd57372, 16'd29990, 16'd19993, 16'd47306, 16'd49840, 16'd13275, 16'd10018, 16'd49983, 16'd2800, 16'd6171, 16'd42085, 16'd47131, 16'd22892, 16'd34960, 16'd1775, 16'd63792, 16'd25430, 16'd47063, 16'd57250, 16'd1681, 16'd8404, 16'd23267, 16'd14249});
	test_expansion(128'h9481def3d5aad0d51e7e045e3ca6ba14, {16'd61204, 16'd52322, 16'd40527, 16'd42756, 16'd53037, 16'd51920, 16'd45622, 16'd3103, 16'd19266, 16'd10657, 16'd36251, 16'd52433, 16'd55531, 16'd57015, 16'd25608, 16'd64624, 16'd53020, 16'd57111, 16'd27403, 16'd14714, 16'd20962, 16'd61317, 16'd16607, 16'd60759, 16'd13796, 16'd15211});
	test_expansion(128'h9d1cc29a072acccf830f75f681106fc0, {16'd22747, 16'd45934, 16'd5426, 16'd37054, 16'd28507, 16'd33788, 16'd30064, 16'd23147, 16'd13829, 16'd23188, 16'd44620, 16'd33588, 16'd58627, 16'd51966, 16'd45239, 16'd29581, 16'd41843, 16'd55100, 16'd28882, 16'd32832, 16'd59465, 16'd43509, 16'd43095, 16'd5137, 16'd46565, 16'd60960});
	test_expansion(128'h94a46ebb49ad3024fe31e4c932657a78, {16'd12979, 16'd48907, 16'd44795, 16'd18473, 16'd11749, 16'd19296, 16'd11007, 16'd19193, 16'd61545, 16'd63330, 16'd65288, 16'd65444, 16'd12723, 16'd8874, 16'd32786, 16'd36783, 16'd40329, 16'd5160, 16'd6548, 16'd58699, 16'd62486, 16'd24325, 16'd22703, 16'd20524, 16'd32265, 16'd53552});
	test_expansion(128'h896e805b8232e5e1a5c27221a89cfc75, {16'd4630, 16'd62852, 16'd14872, 16'd21886, 16'd10140, 16'd43851, 16'd21580, 16'd11983, 16'd15611, 16'd23278, 16'd18834, 16'd34647, 16'd56702, 16'd57869, 16'd57951, 16'd15451, 16'd39679, 16'd38076, 16'd44607, 16'd38854, 16'd7114, 16'd22420, 16'd46836, 16'd3062, 16'd17877, 16'd4322});
	test_expansion(128'h89a672332066fa683a7ad7ec8c9b509e, {16'd59857, 16'd25807, 16'd33254, 16'd39430, 16'd22642, 16'd17094, 16'd4620, 16'd16579, 16'd16224, 16'd32066, 16'd47675, 16'd17850, 16'd24416, 16'd64437, 16'd57117, 16'd30087, 16'd17127, 16'd64982, 16'd6550, 16'd28143, 16'd672, 16'd42641, 16'd6713, 16'd12625, 16'd20414, 16'd54981});
	test_expansion(128'hffd6cb3a6a6f9fb3b686655a0856d11e, {16'd55241, 16'd6056, 16'd54890, 16'd3826, 16'd40143, 16'd44467, 16'd41342, 16'd1256, 16'd33584, 16'd30024, 16'd60803, 16'd7153, 16'd58429, 16'd12095, 16'd42264, 16'd65511, 16'd23695, 16'd4252, 16'd49991, 16'd26579, 16'd38776, 16'd10151, 16'd24766, 16'd23734, 16'd64159, 16'd11753});
	test_expansion(128'hda2f7ac9c6e19f696dabbcf928df4b3e, {16'd63436, 16'd55935, 16'd57914, 16'd16213, 16'd34593, 16'd27901, 16'd4004, 16'd32630, 16'd26459, 16'd18599, 16'd25874, 16'd42209, 16'd65115, 16'd22320, 16'd31665, 16'd16874, 16'd2322, 16'd27693, 16'd51745, 16'd10950, 16'd15727, 16'd48981, 16'd41477, 16'd26649, 16'd16314, 16'd22647});
	test_expansion(128'h8ece6e811c7b7fd6404f25735d2a680b, {16'd60625, 16'd33711, 16'd61864, 16'd35806, 16'd51237, 16'd50229, 16'd26171, 16'd65506, 16'd18255, 16'd37523, 16'd48158, 16'd47050, 16'd7808, 16'd48425, 16'd61571, 16'd26339, 16'd10554, 16'd61137, 16'd56559, 16'd24728, 16'd64114, 16'd33882, 16'd23818, 16'd29775, 16'd143, 16'd33095});
	test_expansion(128'h4ed06aa41b7fcb6fc7d497496e78f8d2, {16'd49450, 16'd36052, 16'd11458, 16'd61000, 16'd5286, 16'd58820, 16'd20911, 16'd20924, 16'd61896, 16'd40757, 16'd8370, 16'd53416, 16'd43944, 16'd33150, 16'd41263, 16'd39777, 16'd4387, 16'd14061, 16'd25753, 16'd5373, 16'd64119, 16'd61980, 16'd26204, 16'd797, 16'd58430, 16'd27202});
	test_expansion(128'hbce643f3d9da599fcce28eabc12dcabc, {16'd63498, 16'd61737, 16'd7834, 16'd38977, 16'd40397, 16'd17654, 16'd33488, 16'd32120, 16'd17094, 16'd62334, 16'd62302, 16'd50054, 16'd19703, 16'd13304, 16'd32260, 16'd7777, 16'd62966, 16'd30914, 16'd18071, 16'd25184, 16'd35059, 16'd6294, 16'd56927, 16'd39489, 16'd17774, 16'd20484});
	test_expansion(128'h9b76f0e4da873f6a6a468fae74eafdc7, {16'd9188, 16'd10220, 16'd57544, 16'd38855, 16'd25342, 16'd57025, 16'd26745, 16'd44906, 16'd46939, 16'd20462, 16'd34648, 16'd28390, 16'd58727, 16'd25451, 16'd21559, 16'd7203, 16'd16780, 16'd5149, 16'd19384, 16'd48607, 16'd6731, 16'd14032, 16'd15105, 16'd35317, 16'd47206, 16'd47642});
	test_expansion(128'hf5f7076f1f26e44b2cb5c8bcaff4df16, {16'd49138, 16'd30022, 16'd13702, 16'd60249, 16'd24472, 16'd304, 16'd41919, 16'd34004, 16'd52121, 16'd795, 16'd12903, 16'd1126, 16'd9091, 16'd42688, 16'd8621, 16'd58802, 16'd14816, 16'd2953, 16'd6890, 16'd6999, 16'd44724, 16'd17090, 16'd57237, 16'd26371, 16'd1382, 16'd58011});
	test_expansion(128'h2793f61cb83a206da1d939477dff953e, {16'd9767, 16'd29770, 16'd22119, 16'd34588, 16'd8044, 16'd21449, 16'd59004, 16'd5754, 16'd16410, 16'd10893, 16'd8729, 16'd39148, 16'd61018, 16'd41864, 16'd60587, 16'd8587, 16'd55191, 16'd30249, 16'd30256, 16'd42948, 16'd37640, 16'd2128, 16'd38429, 16'd60359, 16'd64914, 16'd40393});
	test_expansion(128'h1a6777eb323927e98a419f4b82a0bd70, {16'd59171, 16'd16745, 16'd35568, 16'd50659, 16'd62393, 16'd42364, 16'd4511, 16'd54943, 16'd19086, 16'd34585, 16'd41021, 16'd42592, 16'd18660, 16'd34071, 16'd15954, 16'd37973, 16'd57612, 16'd39696, 16'd39771, 16'd7880, 16'd21674, 16'd26016, 16'd52953, 16'd584, 16'd16712, 16'd48731});
	test_expansion(128'h0a0d89b06c79c95b34cc7e84d2fa00ae, {16'd39401, 16'd19272, 16'd2873, 16'd44256, 16'd8024, 16'd7485, 16'd6562, 16'd22364, 16'd43736, 16'd16738, 16'd58880, 16'd48321, 16'd13958, 16'd25294, 16'd32606, 16'd21156, 16'd54259, 16'd12488, 16'd4836, 16'd28270, 16'd47565, 16'd46848, 16'd34864, 16'd36656, 16'd52597, 16'd51895});
	test_expansion(128'hc2b4dd0a007496ef42958a021fb10977, {16'd36570, 16'd31229, 16'd19054, 16'd8678, 16'd40559, 16'd16700, 16'd56816, 16'd59153, 16'd52650, 16'd26994, 16'd34433, 16'd56020, 16'd46594, 16'd60809, 16'd59575, 16'd1574, 16'd31376, 16'd32337, 16'd5469, 16'd18598, 16'd30715, 16'd22108, 16'd60766, 16'd24800, 16'd37982, 16'd62870});
	test_expansion(128'h90a8268485ed47fa4a755201bfc02232, {16'd15775, 16'd55937, 16'd37806, 16'd28131, 16'd28633, 16'd33665, 16'd41515, 16'd60165, 16'd25770, 16'd59450, 16'd17512, 16'd8760, 16'd1176, 16'd9893, 16'd53709, 16'd22749, 16'd16685, 16'd35479, 16'd1720, 16'd61149, 16'd26054, 16'd7561, 16'd65167, 16'd26754, 16'd3150, 16'd41355});
	test_expansion(128'h881d9c4eddff29dad14b52ef647dc30c, {16'd47883, 16'd38035, 16'd63673, 16'd20401, 16'd60598, 16'd12368, 16'd52461, 16'd3366, 16'd22793, 16'd38057, 16'd256, 16'd26925, 16'd60606, 16'd17603, 16'd1770, 16'd39616, 16'd50192, 16'd16818, 16'd58020, 16'd40858, 16'd20826, 16'd14760, 16'd45622, 16'd45939, 16'd64123, 16'd6866});
	test_expansion(128'h4d3997f5788b5cc0d78e8b60d517f048, {16'd63538, 16'd4263, 16'd24022, 16'd931, 16'd47429, 16'd24671, 16'd28477, 16'd38029, 16'd52694, 16'd43944, 16'd10063, 16'd61564, 16'd45995, 16'd45702, 16'd57766, 16'd57445, 16'd41561, 16'd49279, 16'd14088, 16'd11492, 16'd30469, 16'd252, 16'd20415, 16'd56631, 16'd18331, 16'd51813});
	test_expansion(128'hd3a116f9b383a85373ccbc253adae2e0, {16'd2066, 16'd24981, 16'd36650, 16'd35848, 16'd57358, 16'd44821, 16'd60049, 16'd53520, 16'd41102, 16'd18525, 16'd37491, 16'd9219, 16'd6533, 16'd26753, 16'd18356, 16'd56384, 16'd2293, 16'd63370, 16'd846, 16'd2985, 16'd3820, 16'd19614, 16'd31833, 16'd20453, 16'd21363, 16'd14232});
	test_expansion(128'h7ff18e671d3c4b409babcf750410e92a, {16'd22564, 16'd38787, 16'd45550, 16'd44544, 16'd45435, 16'd28265, 16'd43135, 16'd32045, 16'd11089, 16'd36, 16'd29640, 16'd31690, 16'd65314, 16'd65513, 16'd58250, 16'd3575, 16'd20151, 16'd44721, 16'd31106, 16'd23902, 16'd28659, 16'd2230, 16'd58591, 16'd3195, 16'd61597, 16'd50821});
	test_expansion(128'hc04a0ce70ff13f0ce9676976c89ba66d, {16'd23374, 16'd9636, 16'd23653, 16'd57987, 16'd49761, 16'd50956, 16'd61179, 16'd45493, 16'd25269, 16'd16928, 16'd42530, 16'd52651, 16'd63489, 16'd3279, 16'd24021, 16'd61835, 16'd62426, 16'd29389, 16'd24122, 16'd10844, 16'd51958, 16'd54922, 16'd28165, 16'd58905, 16'd52807, 16'd45238});
	test_expansion(128'h21715ca376c794242bf3f41f1fbf9c9c, {16'd52631, 16'd41315, 16'd50566, 16'd37040, 16'd52444, 16'd30526, 16'd57585, 16'd20137, 16'd48203, 16'd62392, 16'd39104, 16'd9122, 16'd60976, 16'd52172, 16'd34448, 16'd26205, 16'd64044, 16'd36710, 16'd49878, 16'd7902, 16'd13027, 16'd13767, 16'd62634, 16'd26627, 16'd64879, 16'd53558});
	test_expansion(128'h9be17f4b82fd449a5f2110792ace36f3, {16'd39646, 16'd29226, 16'd9238, 16'd51577, 16'd63510, 16'd566, 16'd56961, 16'd31036, 16'd22134, 16'd7689, 16'd16264, 16'd18914, 16'd20757, 16'd7439, 16'd4041, 16'd63636, 16'd63001, 16'd5829, 16'd46340, 16'd16138, 16'd35819, 16'd18491, 16'd46697, 16'd6976, 16'd61398, 16'd4548});
	test_expansion(128'h80b473ac5a6438046b6147ee140cc5a3, {16'd13243, 16'd2537, 16'd42155, 16'd56762, 16'd29959, 16'd33771, 16'd5296, 16'd27158, 16'd53085, 16'd35240, 16'd6644, 16'd30925, 16'd41824, 16'd47373, 16'd55891, 16'd64524, 16'd27909, 16'd58675, 16'd51704, 16'd54177, 16'd57368, 16'd59674, 16'd41712, 16'd20449, 16'd45807, 16'd58816});
	test_expansion(128'hf174cd54f37d9c32b90697c0d72d8fe2, {16'd45094, 16'd55749, 16'd35323, 16'd23257, 16'd45459, 16'd36613, 16'd30078, 16'd55850, 16'd4487, 16'd47722, 16'd17906, 16'd62128, 16'd17787, 16'd15673, 16'd46920, 16'd9984, 16'd32530, 16'd33887, 16'd1319, 16'd17819, 16'd9421, 16'd50768, 16'd2053, 16'd8245, 16'd32994, 16'd63872});
	test_expansion(128'h242b3d84e22fae2341f368600bec5399, {16'd419, 16'd64363, 16'd45888, 16'd55102, 16'd64990, 16'd53881, 16'd14328, 16'd51766, 16'd65404, 16'd45765, 16'd62101, 16'd30781, 16'd39285, 16'd59986, 16'd48621, 16'd43517, 16'd58620, 16'd8945, 16'd10236, 16'd28646, 16'd28921, 16'd58093, 16'd27432, 16'd61584, 16'd47436, 16'd4910});
	test_expansion(128'h36656a480b82fb72968c6610cdd84067, {16'd6558, 16'd63006, 16'd5190, 16'd26730, 16'd57644, 16'd64726, 16'd692, 16'd33718, 16'd21048, 16'd57751, 16'd28982, 16'd61929, 16'd58875, 16'd61873, 16'd27661, 16'd12030, 16'd474, 16'd8045, 16'd15726, 16'd48487, 16'd24871, 16'd62954, 16'd47116, 16'd27365, 16'd17325, 16'd18697});
	test_expansion(128'hca4fe755fb3f1f13c6a6113c70128f15, {16'd48805, 16'd16309, 16'd57772, 16'd53638, 16'd2935, 16'd46861, 16'd13573, 16'd64014, 16'd57942, 16'd31665, 16'd7572, 16'd41480, 16'd10179, 16'd4563, 16'd29811, 16'd6575, 16'd42973, 16'd8391, 16'd64725, 16'd50105, 16'd44189, 16'd19629, 16'd38362, 16'd47334, 16'd6872, 16'd38127});
	test_expansion(128'h017fd306d618eb0a9114f8ce39832deb, {16'd37778, 16'd29291, 16'd25768, 16'd47892, 16'd40967, 16'd8160, 16'd8848, 16'd38785, 16'd29467, 16'd1947, 16'd46674, 16'd12542, 16'd63115, 16'd26121, 16'd24892, 16'd15257, 16'd26456, 16'd13991, 16'd11602, 16'd27376, 16'd10372, 16'd19451, 16'd58605, 16'd62598, 16'd26538, 16'd6669});
	test_expansion(128'hf7ea02b2e93945ebe5f4e52bc0dfac2a, {16'd36301, 16'd44664, 16'd54644, 16'd6101, 16'd12250, 16'd25118, 16'd51027, 16'd34400, 16'd23793, 16'd55522, 16'd30854, 16'd387, 16'd59152, 16'd44913, 16'd12777, 16'd28521, 16'd20599, 16'd51197, 16'd25102, 16'd807, 16'd35470, 16'd29116, 16'd26801, 16'd43966, 16'd45443, 16'd65044});
	test_expansion(128'hf3edf92ee0930d15d6d01b37c84e7a8b, {16'd56201, 16'd35176, 16'd22858, 16'd59798, 16'd10358, 16'd27766, 16'd33151, 16'd24766, 16'd949, 16'd35263, 16'd20239, 16'd53235, 16'd8534, 16'd17043, 16'd61288, 16'd34229, 16'd50748, 16'd33312, 16'd33258, 16'd7326, 16'd1494, 16'd49789, 16'd28942, 16'd50991, 16'd19974, 16'd6974});
	test_expansion(128'h3027d13fb04ed03b9228f65975411063, {16'd54615, 16'd37044, 16'd5943, 16'd988, 16'd55377, 16'd46845, 16'd64601, 16'd62404, 16'd594, 16'd39279, 16'd7977, 16'd32732, 16'd13074, 16'd48187, 16'd60074, 16'd49164, 16'd58358, 16'd29375, 16'd50312, 16'd44738, 16'd33837, 16'd3685, 16'd44430, 16'd9015, 16'd13142, 16'd23317});
	test_expansion(128'h56182b0789f781574c1080fc48bf3e5b, {16'd64977, 16'd38594, 16'd52309, 16'd49646, 16'd37104, 16'd47242, 16'd37383, 16'd2267, 16'd61929, 16'd45332, 16'd28656, 16'd11390, 16'd29851, 16'd49092, 16'd5548, 16'd44661, 16'd50643, 16'd37700, 16'd41779, 16'd60669, 16'd32971, 16'd20849, 16'd12090, 16'd18811, 16'd61723, 16'd17458});
	test_expansion(128'h22fa9620df9481ac44d4e5f8bdb2a5ee, {16'd41457, 16'd1266, 16'd31277, 16'd34311, 16'd49664, 16'd57992, 16'd21544, 16'd19444, 16'd58953, 16'd48354, 16'd14915, 16'd34164, 16'd13925, 16'd748, 16'd10148, 16'd51084, 16'd42992, 16'd19726, 16'd61599, 16'd64640, 16'd47476, 16'd52805, 16'd6100, 16'd34187, 16'd6466, 16'd32045});
	test_expansion(128'h5b89557cb77d22f5d71ac68c4fca464d, {16'd56731, 16'd51740, 16'd28547, 16'd20631, 16'd24534, 16'd10457, 16'd10558, 16'd58046, 16'd19013, 16'd29818, 16'd63904, 16'd11673, 16'd19541, 16'd43106, 16'd13586, 16'd52039, 16'd51343, 16'd35704, 16'd42282, 16'd9502, 16'd49874, 16'd62270, 16'd23897, 16'd8654, 16'd37153, 16'd46497});
	test_expansion(128'h48fc4d572ae2b4aa73c4d105653bd3a2, {16'd44073, 16'd9294, 16'd61000, 16'd51240, 16'd11314, 16'd24999, 16'd39064, 16'd11069, 16'd24953, 16'd57257, 16'd15215, 16'd11491, 16'd42639, 16'd1508, 16'd19537, 16'd1278, 16'd8766, 16'd8379, 16'd57, 16'd676, 16'd55682, 16'd26871, 16'd64647, 16'd61831, 16'd57209, 16'd26760});
	test_expansion(128'h7bbd6f8b0b15aceb308be29a2128cbad, {16'd42759, 16'd31491, 16'd63439, 16'd54885, 16'd22583, 16'd61417, 16'd32525, 16'd52603, 16'd34929, 16'd34749, 16'd30753, 16'd26026, 16'd24889, 16'd33282, 16'd28327, 16'd26843, 16'd15058, 16'd8639, 16'd38063, 16'd45927, 16'd28053, 16'd9312, 16'd40231, 16'd19156, 16'd40910, 16'd61046});
	test_expansion(128'hfa76ca69fc96825767e5ec3d8c88c2c6, {16'd31072, 16'd28996, 16'd9576, 16'd63917, 16'd64229, 16'd47327, 16'd36560, 16'd23298, 16'd39784, 16'd36369, 16'd65162, 16'd6339, 16'd4132, 16'd21197, 16'd11244, 16'd31045, 16'd33260, 16'd52121, 16'd57831, 16'd25629, 16'd50873, 16'd26265, 16'd29339, 16'd12636, 16'd36907, 16'd29647});
	test_expansion(128'h64393fa499eccdc16b94a8efe82f82f5, {16'd47549, 16'd37351, 16'd63741, 16'd54287, 16'd62713, 16'd24054, 16'd55923, 16'd43503, 16'd57006, 16'd3585, 16'd12182, 16'd36425, 16'd55169, 16'd59436, 16'd41848, 16'd44949, 16'd3995, 16'd2315, 16'd42976, 16'd62953, 16'd28341, 16'd24489, 16'd47091, 16'd11346, 16'd10888, 16'd27871});
	test_expansion(128'h5eb082f693ef172e9106e435bfb53dd4, {16'd10647, 16'd2459, 16'd40097, 16'd7162, 16'd25246, 16'd8501, 16'd17029, 16'd35207, 16'd35132, 16'd19933, 16'd25667, 16'd31440, 16'd29241, 16'd17466, 16'd28780, 16'd44084, 16'd10210, 16'd45108, 16'd36290, 16'd53284, 16'd47256, 16'd48012, 16'd24502, 16'd60820, 16'd30241, 16'd35260});
	test_expansion(128'hbc8ad0e37c848e97f2dd75ea0da0cd72, {16'd10244, 16'd32974, 16'd33248, 16'd54655, 16'd53711, 16'd38676, 16'd59354, 16'd19748, 16'd9549, 16'd19777, 16'd38749, 16'd28709, 16'd18906, 16'd41970, 16'd17778, 16'd61226, 16'd11375, 16'd52551, 16'd59373, 16'd16674, 16'd24017, 16'd27229, 16'd64258, 16'd1835, 16'd21618, 16'd49445});
	test_expansion(128'h05f6bc2ff6fe677374ec2264543b209c, {16'd36988, 16'd46709, 16'd4752, 16'd49609, 16'd17661, 16'd64953, 16'd25024, 16'd31920, 16'd42675, 16'd51853, 16'd57033, 16'd51668, 16'd1404, 16'd5187, 16'd53864, 16'd65187, 16'd41132, 16'd42844, 16'd23960, 16'd37531, 16'd7734, 16'd40252, 16'd46973, 16'd24209, 16'd56692, 16'd35246});
	test_expansion(128'heeea1b180e314029b79972c47980d22c, {16'd29742, 16'd52706, 16'd508, 16'd56002, 16'd15043, 16'd13173, 16'd4513, 16'd37318, 16'd45908, 16'd28469, 16'd52269, 16'd26028, 16'd1052, 16'd47191, 16'd43093, 16'd52489, 16'd6720, 16'd30682, 16'd23690, 16'd50406, 16'd62951, 16'd28801, 16'd31285, 16'd54596, 16'd18767, 16'd34380});
	test_expansion(128'h57482e773785e7a65919cc49eaca792c, {16'd62101, 16'd36909, 16'd38056, 16'd59011, 16'd55252, 16'd64942, 16'd32411, 16'd36372, 16'd57309, 16'd4340, 16'd23054, 16'd32189, 16'd41939, 16'd43940, 16'd8255, 16'd53362, 16'd1346, 16'd55757, 16'd16684, 16'd59941, 16'd20865, 16'd3928, 16'd39256, 16'd63067, 16'd64209, 16'd41032});
	test_expansion(128'h4f5aeea9d358ed22326d5813519fc579, {16'd40601, 16'd31790, 16'd28856, 16'd64706, 16'd45407, 16'd24218, 16'd13510, 16'd33765, 16'd35545, 16'd31745, 16'd60659, 16'd43994, 16'd33016, 16'd40476, 16'd36684, 16'd43309, 16'd41865, 16'd23450, 16'd32079, 16'd17746, 16'd12746, 16'd27993, 16'd6859, 16'd29962, 16'd35045, 16'd59092});
	test_expansion(128'h4aab45710c3ad33f99f9d287c92c4b81, {16'd39834, 16'd13414, 16'd32592, 16'd3224, 16'd50518, 16'd33697, 16'd40560, 16'd51354, 16'd54153, 16'd37558, 16'd17029, 16'd35485, 16'd47655, 16'd1070, 16'd61746, 16'd35717, 16'd3470, 16'd29812, 16'd48449, 16'd47958, 16'd53003, 16'd8106, 16'd15834, 16'd13284, 16'd19840, 16'd27941});
	test_expansion(128'h6a29d715e1b43e7a1aadc5768e994220, {16'd34679, 16'd30304, 16'd13373, 16'd19106, 16'd56813, 16'd45690, 16'd30743, 16'd43856, 16'd64670, 16'd13543, 16'd25203, 16'd20564, 16'd12270, 16'd32440, 16'd46693, 16'd32071, 16'd15431, 16'd44226, 16'd1034, 16'd39484, 16'd43065, 16'd11603, 16'd21566, 16'd39239, 16'd17435, 16'd46949});
	test_expansion(128'h6408bba72c06aeff92ba5946313d223a, {16'd32257, 16'd17612, 16'd28863, 16'd48399, 16'd60226, 16'd36319, 16'd28084, 16'd44017, 16'd37066, 16'd22593, 16'd32031, 16'd58320, 16'd32946, 16'd58548, 16'd41055, 16'd29842, 16'd17590, 16'd18835, 16'd20484, 16'd17303, 16'd42364, 16'd5386, 16'd55305, 16'd8113, 16'd34319, 16'd60060});
	test_expansion(128'heb493e0ac9bc2c30d77d0c9dfd6dd3f2, {16'd15504, 16'd40519, 16'd44519, 16'd53969, 16'd9259, 16'd20312, 16'd45923, 16'd7438, 16'd45916, 16'd48644, 16'd48637, 16'd3651, 16'd26408, 16'd16201, 16'd55179, 16'd61708, 16'd33015, 16'd63380, 16'd13085, 16'd29152, 16'd35358, 16'd12140, 16'd63379, 16'd51498, 16'd56371, 16'd52315});
	test_expansion(128'h1ffa20284f71ba34bf73636d9ef217fa, {16'd3816, 16'd16423, 16'd20859, 16'd17250, 16'd64488, 16'd16059, 16'd58110, 16'd22576, 16'd51871, 16'd11225, 16'd19887, 16'd2793, 16'd14005, 16'd39393, 16'd22515, 16'd56078, 16'd38363, 16'd55684, 16'd64123, 16'd21585, 16'd5043, 16'd45650, 16'd43641, 16'd6824, 16'd7900, 16'd65128});
	test_expansion(128'h4881e60bebcb27a8c62fbcd6fb57039e, {16'd52770, 16'd8949, 16'd6478, 16'd6079, 16'd20415, 16'd40668, 16'd41665, 16'd17249, 16'd6323, 16'd849, 16'd3811, 16'd33999, 16'd14664, 16'd34082, 16'd22979, 16'd59597, 16'd53089, 16'd43453, 16'd62488, 16'd3885, 16'd28411, 16'd61667, 16'd30938, 16'd33448, 16'd60324, 16'd57412});
	test_expansion(128'h54097860252622f37a3bbb1fb23425ad, {16'd33979, 16'd18055, 16'd19030, 16'd15954, 16'd5639, 16'd51040, 16'd52720, 16'd9963, 16'd16620, 16'd44352, 16'd60027, 16'd39494, 16'd47235, 16'd13413, 16'd11626, 16'd48364, 16'd43891, 16'd54538, 16'd10296, 16'd63210, 16'd23748, 16'd18518, 16'd10333, 16'd3, 16'd16489, 16'd35243});
	test_expansion(128'hfe3f62da45b2391452a1b97b5dcb3555, {16'd8206, 16'd50666, 16'd2383, 16'd20381, 16'd45221, 16'd4167, 16'd44843, 16'd8531, 16'd57716, 16'd8858, 16'd4894, 16'd57251, 16'd31529, 16'd10513, 16'd40835, 16'd4677, 16'd44576, 16'd25714, 16'd62787, 16'd48845, 16'd55735, 16'd22967, 16'd56188, 16'd64539, 16'd5798, 16'd2027});
	test_expansion(128'hb2d3a3010923468e19948ff98b8bddd2, {16'd50207, 16'd47031, 16'd943, 16'd14253, 16'd27416, 16'd42749, 16'd15433, 16'd13002, 16'd18048, 16'd61622, 16'd5958, 16'd48846, 16'd44468, 16'd45576, 16'd19060, 16'd61600, 16'd51468, 16'd28386, 16'd50683, 16'd6812, 16'd14798, 16'd32417, 16'd25641, 16'd48770, 16'd11172, 16'd3555});
	test_expansion(128'hc535b9cbc064b88d09c7b9b70d06d31e, {16'd51887, 16'd23272, 16'd261, 16'd15216, 16'd5593, 16'd61989, 16'd3391, 16'd64488, 16'd54641, 16'd36988, 16'd23571, 16'd41369, 16'd49577, 16'd52558, 16'd45781, 16'd7535, 16'd54899, 16'd55606, 16'd55221, 16'd27048, 16'd54176, 16'd6830, 16'd41301, 16'd54243, 16'd27967, 16'd56802});
	test_expansion(128'h5ad820a7ed6f605ac4069502b20431f6, {16'd6046, 16'd26768, 16'd54656, 16'd26632, 16'd31061, 16'd49641, 16'd45136, 16'd43005, 16'd1471, 16'd11713, 16'd48557, 16'd34647, 16'd24427, 16'd62602, 16'd58332, 16'd43597, 16'd13392, 16'd20608, 16'd24175, 16'd42334, 16'd23300, 16'd33071, 16'd60563, 16'd41366, 16'd57568, 16'd21016});
	test_expansion(128'hc0e308dd4887e565acab216657770ccd, {16'd40620, 16'd25766, 16'd8116, 16'd39236, 16'd33255, 16'd19919, 16'd62223, 16'd48797, 16'd61247, 16'd63471, 16'd16895, 16'd34129, 16'd14905, 16'd63278, 16'd10257, 16'd1813, 16'd32852, 16'd53666, 16'd29428, 16'd38314, 16'd37417, 16'd33727, 16'd54864, 16'd23444, 16'd17476, 16'd47899});
	test_expansion(128'h189660f454a45ef9ed87d8210dfa1154, {16'd14388, 16'd58121, 16'd49665, 16'd20675, 16'd27795, 16'd29885, 16'd54737, 16'd13374, 16'd50660, 16'd44816, 16'd8939, 16'd16261, 16'd49398, 16'd6194, 16'd63819, 16'd13239, 16'd24498, 16'd55215, 16'd49981, 16'd14869, 16'd51762, 16'd62033, 16'd37172, 16'd1251, 16'd44462, 16'd55315});
	test_expansion(128'hc27181eaadf901601f64b35ae1661a59, {16'd43549, 16'd13340, 16'd22851, 16'd54049, 16'd26383, 16'd30890, 16'd25049, 16'd41391, 16'd42424, 16'd4340, 16'd64693, 16'd45251, 16'd30937, 16'd40032, 16'd1368, 16'd24091, 16'd59665, 16'd57972, 16'd11650, 16'd38741, 16'd12504, 16'd21403, 16'd35371, 16'd49867, 16'd35999, 16'd2831});
	test_expansion(128'h4ba62146fc329ec02a94440a8ca39631, {16'd47385, 16'd10181, 16'd60799, 16'd53670, 16'd46140, 16'd16211, 16'd8556, 16'd27990, 16'd21432, 16'd11572, 16'd48271, 16'd11730, 16'd40116, 16'd50688, 16'd54462, 16'd51916, 16'd62913, 16'd1031, 16'd3740, 16'd53569, 16'd45049, 16'd54529, 16'd15517, 16'd35950, 16'd43292, 16'd3045});
	test_expansion(128'he5b7a2283a56b6a3cdb77c155875d909, {16'd62879, 16'd54667, 16'd29346, 16'd30304, 16'd32500, 16'd26622, 16'd25628, 16'd11081, 16'd9168, 16'd47591, 16'd5943, 16'd47607, 16'd7916, 16'd61182, 16'd62588, 16'd54559, 16'd15463, 16'd32167, 16'd56380, 16'd15589, 16'd58010, 16'd30980, 16'd31237, 16'd47534, 16'd61890, 16'd46533});
	test_expansion(128'h8e921fdcf246f377d8348a05e92a3e57, {16'd45860, 16'd7567, 16'd46783, 16'd3443, 16'd19122, 16'd23571, 16'd2899, 16'd31396, 16'd16219, 16'd21871, 16'd58529, 16'd5132, 16'd28628, 16'd19154, 16'd58008, 16'd16753, 16'd673, 16'd61163, 16'd38363, 16'd28297, 16'd40149, 16'd35636, 16'd52636, 16'd34685, 16'd23842, 16'd14138});
	test_expansion(128'h12e7ca858c8cab45c846bce3b3e5f48f, {16'd33554, 16'd56055, 16'd62872, 16'd59116, 16'd25661, 16'd27640, 16'd64224, 16'd52037, 16'd30861, 16'd37913, 16'd53970, 16'd49756, 16'd28443, 16'd194, 16'd29995, 16'd37737, 16'd59264, 16'd8599, 16'd11882, 16'd59089, 16'd17685, 16'd3094, 16'd54852, 16'd4649, 16'd15503, 16'd60754});
	test_expansion(128'h48b7e2ff98d29285bb31edf26fc51da9, {16'd16251, 16'd56044, 16'd23738, 16'd4187, 16'd9532, 16'd26375, 16'd33291, 16'd31734, 16'd40115, 16'd62232, 16'd5248, 16'd26237, 16'd28392, 16'd62649, 16'd40244, 16'd46647, 16'd4268, 16'd21424, 16'd7227, 16'd63236, 16'd58821, 16'd40528, 16'd48063, 16'd56655, 16'd52328, 16'd9627});
	test_expansion(128'h6287a4b1801214977c2deed0b81bbe88, {16'd56002, 16'd19648, 16'd21849, 16'd60183, 16'd48399, 16'd49746, 16'd65504, 16'd8714, 16'd17534, 16'd55346, 16'd44887, 16'd46675, 16'd10504, 16'd44679, 16'd21242, 16'd49463, 16'd3745, 16'd56924, 16'd58027, 16'd38946, 16'd53910, 16'd8506, 16'd42166, 16'd59702, 16'd63849, 16'd35809});
	test_expansion(128'hb29e3cdd4bc467f9f895f57b111223c1, {16'd56772, 16'd50350, 16'd14838, 16'd24975, 16'd64105, 16'd63772, 16'd37440, 16'd58471, 16'd20248, 16'd11036, 16'd53206, 16'd60504, 16'd16106, 16'd29698, 16'd11306, 16'd9540, 16'd56638, 16'd44412, 16'd26918, 16'd62888, 16'd48046, 16'd19539, 16'd50344, 16'd40360, 16'd9281, 16'd2223});
	test_expansion(128'he41e2a6623cf09ed7d4f61b1ff9700c7, {16'd56038, 16'd25767, 16'd61908, 16'd60589, 16'd29705, 16'd1659, 16'd59917, 16'd58326, 16'd45779, 16'd27166, 16'd60435, 16'd28724, 16'd12209, 16'd41025, 16'd35983, 16'd35076, 16'd11778, 16'd36363, 16'd19626, 16'd1560, 16'd4790, 16'd22973, 16'd1528, 16'd42850, 16'd48848, 16'd25292});
	test_expansion(128'hd2d8cdc5ebc4901e854e8c2477129ecf, {16'd49295, 16'd5002, 16'd10529, 16'd59051, 16'd64401, 16'd62208, 16'd62302, 16'd55575, 16'd36381, 16'd24212, 16'd9091, 16'd3905, 16'd44261, 16'd59791, 16'd3437, 16'd25265, 16'd7692, 16'd19139, 16'd31675, 16'd15264, 16'd40226, 16'd19890, 16'd33606, 16'd23110, 16'd6702, 16'd60397});
	test_expansion(128'h729b283ee7ac6a943a0f3c3bf3360aa9, {16'd29263, 16'd60539, 16'd19156, 16'd38941, 16'd58631, 16'd62785, 16'd21634, 16'd24900, 16'd55120, 16'd61568, 16'd9038, 16'd302, 16'd57283, 16'd4048, 16'd1842, 16'd34991, 16'd39380, 16'd41571, 16'd29692, 16'd43087, 16'd48328, 16'd15786, 16'd29893, 16'd7098, 16'd44846, 16'd48060});
	test_expansion(128'hc4de5bebf15f230f0c6735615aa4cb7e, {16'd11291, 16'd49260, 16'd53085, 16'd58083, 16'd4952, 16'd3783, 16'd14533, 16'd58000, 16'd42982, 16'd24610, 16'd2120, 16'd55509, 16'd53087, 16'd20947, 16'd31344, 16'd41853, 16'd57693, 16'd21762, 16'd38653, 16'd46963, 16'd36238, 16'd53515, 16'd59918, 16'd6170, 16'd60429, 16'd6016});
	test_expansion(128'h03185c6d243119e983808aa4a1eca77f, {16'd23023, 16'd42296, 16'd50132, 16'd874, 16'd61080, 16'd32056, 16'd5587, 16'd11917, 16'd59275, 16'd37901, 16'd61333, 16'd6513, 16'd29525, 16'd57111, 16'd40319, 16'd48688, 16'd51248, 16'd8838, 16'd42819, 16'd28048, 16'd2992, 16'd35747, 16'd5361, 16'd34768, 16'd50568, 16'd60740});
	test_expansion(128'h540b7bd47e4a2a5fa3f543c50eb7dc05, {16'd3880, 16'd29869, 16'd55015, 16'd53427, 16'd52023, 16'd31956, 16'd20397, 16'd7061, 16'd43714, 16'd18706, 16'd17015, 16'd46070, 16'd34377, 16'd20063, 16'd50669, 16'd16134, 16'd52904, 16'd57938, 16'd7601, 16'd26174, 16'd31886, 16'd8963, 16'd4254, 16'd41545, 16'd7751, 16'd36767});
	test_expansion(128'hcb92f489ad3f4602b5b70a3fa60b7bb5, {16'd46569, 16'd7274, 16'd51181, 16'd20262, 16'd28777, 16'd18602, 16'd62302, 16'd37239, 16'd16019, 16'd14336, 16'd52841, 16'd43718, 16'd47070, 16'd8910, 16'd44483, 16'd1051, 16'd20758, 16'd57310, 16'd38436, 16'd9127, 16'd55731, 16'd36816, 16'd58302, 16'd10338, 16'd4536, 16'd10540});
	test_expansion(128'h1e79c79a18304c68e45a43b1acd0c3b5, {16'd49548, 16'd49176, 16'd25178, 16'd62961, 16'd46127, 16'd20624, 16'd20728, 16'd42935, 16'd15438, 16'd20966, 16'd62862, 16'd38910, 16'd33183, 16'd24963, 16'd19195, 16'd43053, 16'd34076, 16'd58520, 16'd25734, 16'd62399, 16'd13169, 16'd3273, 16'd24370, 16'd31410, 16'd26897, 16'd42656});
	test_expansion(128'h0e815fe39fd624fbfc0ce9b514a4faa6, {16'd28077, 16'd50638, 16'd21488, 16'd52394, 16'd48385, 16'd30611, 16'd28377, 16'd39894, 16'd898, 16'd61326, 16'd26781, 16'd9873, 16'd4661, 16'd38648, 16'd145, 16'd36410, 16'd31625, 16'd161, 16'd4932, 16'd6634, 16'd9844, 16'd41448, 16'd32347, 16'd35250, 16'd10140, 16'd41405});
	test_expansion(128'hb4fe1e8286959c08cd73f6ae65d2ad0b, {16'd40237, 16'd6684, 16'd14844, 16'd61191, 16'd35613, 16'd44145, 16'd34993, 16'd45804, 16'd170, 16'd43585, 16'd24744, 16'd26766, 16'd47896, 16'd57260, 16'd24265, 16'd60588, 16'd26563, 16'd7829, 16'd19065, 16'd16347, 16'd63740, 16'd54111, 16'd19977, 16'd19417, 16'd21269, 16'd5360});
	test_expansion(128'h683a3a636357feb93f3b76f40aa17a6b, {16'd40196, 16'd23010, 16'd44190, 16'd3698, 16'd27387, 16'd50409, 16'd3902, 16'd50728, 16'd42793, 16'd52608, 16'd31117, 16'd12295, 16'd58283, 16'd38329, 16'd47028, 16'd31401, 16'd31643, 16'd60927, 16'd37237, 16'd55868, 16'd49531, 16'd19847, 16'd48022, 16'd7445, 16'd28278, 16'd13652});
	test_expansion(128'h401106deb4829c3601c059f0ac22b560, {16'd45383, 16'd13599, 16'd64543, 16'd43475, 16'd58161, 16'd18878, 16'd8457, 16'd40741, 16'd35843, 16'd22508, 16'd33378, 16'd48674, 16'd8138, 16'd31385, 16'd3420, 16'd53956, 16'd14191, 16'd63071, 16'd22189, 16'd814, 16'd20884, 16'd47867, 16'd63726, 16'd44048, 16'd39943, 16'd27001});
	test_expansion(128'hdd8cc45f44974bd5df28109b79391271, {16'd60000, 16'd513, 16'd35463, 16'd41040, 16'd6926, 16'd6150, 16'd41614, 16'd25391, 16'd64350, 16'd46208, 16'd19104, 16'd54800, 16'd51247, 16'd26987, 16'd54190, 16'd42920, 16'd26775, 16'd41356, 16'd5907, 16'd40721, 16'd21270, 16'd30645, 16'd10092, 16'd27317, 16'd46913, 16'd51753});
	test_expansion(128'hf1f45d59597ced905de03379d55ee698, {16'd53237, 16'd17088, 16'd14996, 16'd55405, 16'd17393, 16'd30929, 16'd30226, 16'd9335, 16'd30821, 16'd33455, 16'd38254, 16'd43365, 16'd14167, 16'd60014, 16'd22150, 16'd40849, 16'd60232, 16'd3560, 16'd39871, 16'd32964, 16'd19166, 16'd56976, 16'd8777, 16'd14815, 16'd49213, 16'd18186});
	test_expansion(128'hf1be798ae89fe578849c5bcb014bb31b, {16'd60038, 16'd40740, 16'd33347, 16'd57254, 16'd12640, 16'd10577, 16'd63566, 16'd9595, 16'd61027, 16'd38344, 16'd38790, 16'd64302, 16'd37014, 16'd58816, 16'd30911, 16'd25547, 16'd35271, 16'd36417, 16'd25569, 16'd28536, 16'd372, 16'd2215, 16'd56330, 16'd31474, 16'd31474, 16'd64217});
	test_expansion(128'hd280b4eb0417d73036f31f67a46cb3a5, {16'd22666, 16'd1960, 16'd5862, 16'd57145, 16'd53661, 16'd262, 16'd29803, 16'd1189, 16'd31531, 16'd57756, 16'd40491, 16'd28479, 16'd41474, 16'd51098, 16'd3773, 16'd7843, 16'd30281, 16'd23735, 16'd47581, 16'd14344, 16'd11517, 16'd60026, 16'd10596, 16'd15654, 16'd34613, 16'd63511});
	test_expansion(128'hd6445fcd0fe8cbc5e22198176792a44a, {16'd46672, 16'd20332, 16'd50954, 16'd64786, 16'd1462, 16'd32988, 16'd20558, 16'd46359, 16'd60518, 16'd15898, 16'd1663, 16'd64950, 16'd48715, 16'd17190, 16'd33256, 16'd30732, 16'd28208, 16'd56899, 16'd16879, 16'd52579, 16'd1194, 16'd58990, 16'd24411, 16'd55499, 16'd17067, 16'd10783});
	test_expansion(128'haa186537a7c7b3180f6bf209585facbc, {16'd57757, 16'd21532, 16'd30221, 16'd63685, 16'd56367, 16'd8140, 16'd24170, 16'd18372, 16'd52866, 16'd18293, 16'd40556, 16'd63674, 16'd18588, 16'd45947, 16'd46915, 16'd10164, 16'd13506, 16'd57192, 16'd1168, 16'd34682, 16'd55463, 16'd57288, 16'd34769, 16'd25724, 16'd57723, 16'd58858});
	test_expansion(128'h2a1d2c9fca6f9da5ffa73252b7dcf490, {16'd7956, 16'd43406, 16'd31441, 16'd47628, 16'd31516, 16'd49212, 16'd44486, 16'd23536, 16'd65201, 16'd54698, 16'd26301, 16'd7920, 16'd49203, 16'd58520, 16'd21653, 16'd33005, 16'd6129, 16'd43235, 16'd17833, 16'd61434, 16'd25462, 16'd33887, 16'd53045, 16'd21209, 16'd34906, 16'd34124});
	test_expansion(128'h7cd9e576f63cb47b4df9c93743ca3f73, {16'd47772, 16'd17402, 16'd39086, 16'd25909, 16'd21066, 16'd34202, 16'd49335, 16'd18073, 16'd18093, 16'd55465, 16'd10596, 16'd29035, 16'd34326, 16'd64125, 16'd26078, 16'd23422, 16'd5780, 16'd54679, 16'd41004, 16'd10763, 16'd27472, 16'd52924, 16'd37026, 16'd4800, 16'd10902, 16'd29356});
	test_expansion(128'hbef5002fd51af39aae89e2ecff8c6714, {16'd32710, 16'd30363, 16'd30132, 16'd65346, 16'd52255, 16'd3281, 16'd61204, 16'd37440, 16'd55267, 16'd40278, 16'd8385, 16'd41441, 16'd26456, 16'd8809, 16'd59094, 16'd38075, 16'd59795, 16'd9620, 16'd60204, 16'd46920, 16'd2742, 16'd31365, 16'd36460, 16'd56088, 16'd9967, 16'd29920});
	test_expansion(128'hcfc0e34f41d2af115111454b1addc051, {16'd54260, 16'd29551, 16'd16997, 16'd34823, 16'd9202, 16'd18799, 16'd31358, 16'd58013, 16'd31505, 16'd8837, 16'd12714, 16'd54989, 16'd59985, 16'd55361, 16'd62109, 16'd39948, 16'd35879, 16'd63424, 16'd41960, 16'd7934, 16'd58442, 16'd24022, 16'd49744, 16'd11363, 16'd39033, 16'd19774});
	test_expansion(128'h0ea396af4ff50f00d36a6304f73b4899, {16'd42139, 16'd42733, 16'd27201, 16'd1625, 16'd52252, 16'd35804, 16'd134, 16'd27515, 16'd52124, 16'd42534, 16'd11462, 16'd2970, 16'd35684, 16'd18982, 16'd37193, 16'd55496, 16'd17023, 16'd41611, 16'd31460, 16'd49397, 16'd49776, 16'd55467, 16'd16511, 16'd42946, 16'd17074, 16'd10574});
	test_expansion(128'h83e18b915160335eab224c3403e14748, {16'd20484, 16'd59168, 16'd39542, 16'd15731, 16'd25300, 16'd12118, 16'd43846, 16'd60494, 16'd11795, 16'd6798, 16'd65352, 16'd63185, 16'd53243, 16'd21276, 16'd52003, 16'd843, 16'd42181, 16'd61107, 16'd36650, 16'd14922, 16'd45814, 16'd49044, 16'd43239, 16'd64724, 16'd38622, 16'd63437});
	test_expansion(128'hb2a721c760e0956041ca17cac5cff735, {16'd52141, 16'd30656, 16'd45616, 16'd40675, 16'd5682, 16'd62579, 16'd11305, 16'd5371, 16'd45403, 16'd23023, 16'd57919, 16'd54357, 16'd25866, 16'd563, 16'd56977, 16'd3142, 16'd42669, 16'd64907, 16'd48429, 16'd64504, 16'd65478, 16'd62254, 16'd16866, 16'd281, 16'd42417, 16'd15558});
	test_expansion(128'hc53948129009b06d31adaa10807145a8, {16'd50309, 16'd37860, 16'd28612, 16'd11018, 16'd3944, 16'd8123, 16'd61107, 16'd46182, 16'd18333, 16'd9520, 16'd31502, 16'd23309, 16'd5149, 16'd61101, 16'd38628, 16'd13214, 16'd11175, 16'd14729, 16'd26983, 16'd57490, 16'd49670, 16'd4426, 16'd47570, 16'd43148, 16'd3962, 16'd29225});
	test_expansion(128'h5b17b92d595c9c1402c132c5e89ef494, {16'd58069, 16'd7432, 16'd59685, 16'd37198, 16'd57392, 16'd4076, 16'd61055, 16'd63276, 16'd34058, 16'd56992, 16'd16657, 16'd54053, 16'd35631, 16'd42569, 16'd44809, 16'd47514, 16'd52565, 16'd8830, 16'd12426, 16'd14965, 16'd17279, 16'd62075, 16'd36961, 16'd64015, 16'd51166, 16'd39378});
	test_expansion(128'h610758c3287302a0676bb0a62bb6f4c2, {16'd27749, 16'd47608, 16'd59597, 16'd31240, 16'd17004, 16'd29168, 16'd63924, 16'd15980, 16'd2861, 16'd35783, 16'd43110, 16'd49663, 16'd5893, 16'd11151, 16'd23816, 16'd26259, 16'd40237, 16'd51252, 16'd39334, 16'd5594, 16'd8855, 16'd38271, 16'd10871, 16'd14773, 16'd43930, 16'd28171});
	test_expansion(128'h4919f930f43c60345eb8e735e915187b, {16'd11551, 16'd63222, 16'd39262, 16'd18119, 16'd48550, 16'd49177, 16'd46291, 16'd7225, 16'd45811, 16'd18581, 16'd60153, 16'd30170, 16'd37668, 16'd3820, 16'd30381, 16'd30258, 16'd42825, 16'd63414, 16'd15612, 16'd38840, 16'd30079, 16'd13817, 16'd26342, 16'd42083, 16'd8093, 16'd5159});
	test_expansion(128'h5e5cef1eed74810c622f76c64e01045e, {16'd20198, 16'd47412, 16'd49483, 16'd64002, 16'd16576, 16'd6797, 16'd61448, 16'd60250, 16'd20740, 16'd39412, 16'd1516, 16'd35180, 16'd7234, 16'd7348, 16'd45070, 16'd21104, 16'd10955, 16'd12321, 16'd1703, 16'd3086, 16'd41764, 16'd11752, 16'd12816, 16'd51624, 16'd19956, 16'd19268});
	test_expansion(128'h9988e8e687ec21531e4202645fe6dade, {16'd39444, 16'd47322, 16'd11035, 16'd22105, 16'd22340, 16'd50905, 16'd494, 16'd34404, 16'd23095, 16'd22623, 16'd42359, 16'd64151, 16'd34686, 16'd20755, 16'd23632, 16'd4242, 16'd41590, 16'd9930, 16'd59392, 16'd17163, 16'd25140, 16'd34734, 16'd10672, 16'd46645, 16'd17905, 16'd34050});
	test_expansion(128'h0a4b9ed832035fe8068c7456aaa0a147, {16'd38532, 16'd20922, 16'd24452, 16'd32327, 16'd55330, 16'd8811, 16'd9345, 16'd13221, 16'd341, 16'd11963, 16'd64896, 16'd30552, 16'd42128, 16'd43824, 16'd11323, 16'd41509, 16'd26454, 16'd31798, 16'd5496, 16'd51851, 16'd53911, 16'd41432, 16'd4976, 16'd53203, 16'd6794, 16'd21712});
	test_expansion(128'h2727e62d08f13981984812ba3eb8ac34, {16'd8246, 16'd43917, 16'd28830, 16'd14279, 16'd55280, 16'd55279, 16'd45797, 16'd16889, 16'd60175, 16'd48826, 16'd26677, 16'd62658, 16'd32863, 16'd58308, 16'd6423, 16'd1507, 16'd34646, 16'd12323, 16'd26850, 16'd9593, 16'd51152, 16'd19943, 16'd36018, 16'd12617, 16'd11842, 16'd51020});
	test_expansion(128'hd469b80a3bc6d34fe1155d6f0266161d, {16'd43463, 16'd51014, 16'd8794, 16'd39917, 16'd10208, 16'd8879, 16'd37677, 16'd8185, 16'd48038, 16'd29694, 16'd41957, 16'd11879, 16'd47066, 16'd58757, 16'd5739, 16'd27236, 16'd4431, 16'd15381, 16'd50685, 16'd59081, 16'd55852, 16'd51583, 16'd32990, 16'd32140, 16'd3029, 16'd4932});
	test_expansion(128'h594526bf69de9dc068205d9a69e18107, {16'd37261, 16'd4388, 16'd12217, 16'd41987, 16'd33287, 16'd55210, 16'd41175, 16'd11291, 16'd49102, 16'd41613, 16'd29517, 16'd31867, 16'd49498, 16'd19026, 16'd63675, 16'd34143, 16'd24277, 16'd51638, 16'd13800, 16'd6188, 16'd32983, 16'd48463, 16'd30807, 16'd58798, 16'd58146, 16'd41200});
	test_expansion(128'h8d5d717b2b73cf2fe25d60c46107bf73, {16'd51154, 16'd24333, 16'd16633, 16'd45690, 16'd65000, 16'd17599, 16'd8513, 16'd52474, 16'd1689, 16'd28355, 16'd6833, 16'd28825, 16'd59223, 16'd29518, 16'd53939, 16'd2081, 16'd64644, 16'd2070, 16'd20170, 16'd23027, 16'd25286, 16'd57712, 16'd26166, 16'd6233, 16'd33838, 16'd25599});
	test_expansion(128'hf501a8981003015acba29cd41afac112, {16'd20182, 16'd29915, 16'd61685, 16'd55210, 16'd14753, 16'd9272, 16'd11338, 16'd31630, 16'd55227, 16'd52049, 16'd30263, 16'd42096, 16'd8728, 16'd9053, 16'd56675, 16'd49297, 16'd23207, 16'd8753, 16'd3785, 16'd12349, 16'd47383, 16'd24871, 16'd51158, 16'd29852, 16'd7437, 16'd17173});
	test_expansion(128'hd22ed6aa947f2d4571905f9d638519d6, {16'd59488, 16'd21845, 16'd63312, 16'd25749, 16'd47605, 16'd38279, 16'd22593, 16'd28521, 16'd48335, 16'd18760, 16'd24956, 16'd27930, 16'd61078, 16'd65335, 16'd34926, 16'd12140, 16'd39829, 16'd60751, 16'd4826, 16'd61516, 16'd4690, 16'd5315, 16'd50654, 16'd24408, 16'd37047, 16'd4093});
	test_expansion(128'hcbdf7bf7612960cde34b7f18ebf78361, {16'd34058, 16'd18074, 16'd44848, 16'd32367, 16'd21123, 16'd37780, 16'd35563, 16'd53934, 16'd64291, 16'd64359, 16'd56818, 16'd52329, 16'd20890, 16'd36301, 16'd53893, 16'd53914, 16'd28992, 16'd19027, 16'd34219, 16'd52407, 16'd52126, 16'd65210, 16'd60947, 16'd8010, 16'd41773, 16'd64637});
	test_expansion(128'h3c8f258cbdad288df34e0f16172b4082, {16'd39921, 16'd28654, 16'd4297, 16'd41004, 16'd62683, 16'd46582, 16'd49141, 16'd41624, 16'd63483, 16'd63039, 16'd38168, 16'd52008, 16'd22554, 16'd11716, 16'd34419, 16'd528, 16'd30807, 16'd37192, 16'd31747, 16'd59009, 16'd59719, 16'd24963, 16'd7927, 16'd51411, 16'd31149, 16'd17512});
	test_expansion(128'h8bc69155014d7729769434186bbad820, {16'd31804, 16'd7698, 16'd60028, 16'd47477, 16'd35801, 16'd14838, 16'd34468, 16'd28353, 16'd24980, 16'd60133, 16'd33227, 16'd56815, 16'd57440, 16'd59740, 16'd10548, 16'd28512, 16'd47306, 16'd30362, 16'd55973, 16'd34120, 16'd36043, 16'd43870, 16'd8306, 16'd5741, 16'd23932, 16'd19513});
	test_expansion(128'ha6f457e2d7a7b609a4fab742a52b45ba, {16'd54010, 16'd287, 16'd5785, 16'd60365, 16'd48198, 16'd33373, 16'd49828, 16'd28708, 16'd24023, 16'd42826, 16'd26054, 16'd46609, 16'd63483, 16'd6944, 16'd26072, 16'd52274, 16'd18757, 16'd25540, 16'd4800, 16'd19382, 16'd36975, 16'd4481, 16'd43815, 16'd30957, 16'd43, 16'd21110});
	test_expansion(128'hbeded5a67ec763a059309bbe398b344e, {16'd12569, 16'd5197, 16'd21710, 16'd58646, 16'd3990, 16'd24997, 16'd32913, 16'd34148, 16'd38791, 16'd60577, 16'd33283, 16'd62867, 16'd60676, 16'd12576, 16'd10694, 16'd51221, 16'd13096, 16'd35503, 16'd58035, 16'd51323, 16'd11110, 16'd5337, 16'd30720, 16'd11877, 16'd8635, 16'd27999});
	test_expansion(128'h4e7664d14574e485db5a67e72278b332, {16'd20390, 16'd31041, 16'd8933, 16'd49381, 16'd22525, 16'd62309, 16'd50846, 16'd33179, 16'd6291, 16'd14697, 16'd12889, 16'd24487, 16'd24890, 16'd59214, 16'd18382, 16'd50427, 16'd61459, 16'd45988, 16'd15663, 16'd62710, 16'd41579, 16'd15348, 16'd26407, 16'd17287, 16'd17271, 16'd48154});
	test_expansion(128'haa577feb14b3c3569c325f92012d25b3, {16'd46325, 16'd9644, 16'd22399, 16'd677, 16'd32352, 16'd12527, 16'd22218, 16'd62356, 16'd17611, 16'd35396, 16'd48313, 16'd46584, 16'd38924, 16'd56166, 16'd56887, 16'd43542, 16'd30674, 16'd814, 16'd36929, 16'd39871, 16'd63535, 16'd64915, 16'd59325, 16'd2511, 16'd43515, 16'd23061});
	test_expansion(128'h790df2c7a3b429a960944633a4f8b0fa, {16'd21195, 16'd16454, 16'd49556, 16'd70, 16'd19175, 16'd19378, 16'd29318, 16'd50052, 16'd55424, 16'd41709, 16'd52041, 16'd59152, 16'd55921, 16'd29733, 16'd21502, 16'd37522, 16'd49780, 16'd15375, 16'd34400, 16'd7228, 16'd5838, 16'd34652, 16'd42946, 16'd16181, 16'd28073, 16'd40574});
	test_expansion(128'h6755efc10e1c2bea33e4c5f95716a92a, {16'd55611, 16'd65352, 16'd63620, 16'd4930, 16'd20288, 16'd21560, 16'd60442, 16'd31896, 16'd32336, 16'd58126, 16'd53959, 16'd10799, 16'd57860, 16'd51301, 16'd42065, 16'd57249, 16'd249, 16'd32698, 16'd19234, 16'd59650, 16'd17961, 16'd45763, 16'd10894, 16'd13349, 16'd31737, 16'd20765});
	test_expansion(128'hd6265a0704758005e15a0637787bafc7, {16'd41542, 16'd27281, 16'd4376, 16'd44017, 16'd44670, 16'd54284, 16'd40997, 16'd60416, 16'd10103, 16'd4352, 16'd41244, 16'd65386, 16'd60726, 16'd10634, 16'd64923, 16'd46879, 16'd20212, 16'd7081, 16'd44807, 16'd2759, 16'd20334, 16'd33307, 16'd61028, 16'd55943, 16'd56763, 16'd27382});
	test_expansion(128'h4348e3631bb87d4a5ec2637e88a0757d, {16'd37728, 16'd30220, 16'd26994, 16'd63443, 16'd37636, 16'd17703, 16'd52487, 16'd7483, 16'd54702, 16'd48569, 16'd22494, 16'd53176, 16'd6659, 16'd62797, 16'd29799, 16'd47470, 16'd58767, 16'd27014, 16'd44321, 16'd14691, 16'd9289, 16'd41693, 16'd17028, 16'd1012, 16'd53892, 16'd14066});
	test_expansion(128'hf62905a7b61cb787cc7e06085fc5b5f9, {16'd38500, 16'd48909, 16'd42232, 16'd29628, 16'd18288, 16'd12170, 16'd28379, 16'd55843, 16'd54918, 16'd1545, 16'd13623, 16'd51890, 16'd23042, 16'd34141, 16'd39684, 16'd36285, 16'd29073, 16'd2781, 16'd21176, 16'd55172, 16'd58658, 16'd8090, 16'd39697, 16'd50388, 16'd19680, 16'd24279});
	test_expansion(128'h2b184a5891d16b4b7086c34eb1f9dfd6, {16'd40857, 16'd42641, 16'd6588, 16'd41172, 16'd6951, 16'd33563, 16'd31271, 16'd19111, 16'd45664, 16'd31872, 16'd37450, 16'd47471, 16'd8129, 16'd28084, 16'd6497, 16'd51119, 16'd33957, 16'd8073, 16'd34093, 16'd54038, 16'd41864, 16'd52726, 16'd63925, 16'd32028, 16'd10677, 16'd4519});
	test_expansion(128'h79cba87dd03959c45949a1b600ce165e, {16'd10700, 16'd4796, 16'd7637, 16'd24583, 16'd15761, 16'd61243, 16'd7908, 16'd48101, 16'd49008, 16'd34730, 16'd33715, 16'd25214, 16'd52598, 16'd31549, 16'd2594, 16'd39986, 16'd43837, 16'd29924, 16'd11726, 16'd32684, 16'd7194, 16'd25715, 16'd21568, 16'd41917, 16'd46745, 16'd40120});
	test_expansion(128'h022c1cc86c581c915379f494aed1add2, {16'd6647, 16'd10637, 16'd14469, 16'd27374, 16'd60732, 16'd54982, 16'd58638, 16'd34623, 16'd4972, 16'd24138, 16'd31232, 16'd28999, 16'd19832, 16'd45268, 16'd59989, 16'd32234, 16'd55972, 16'd34146, 16'd45831, 16'd41310, 16'd50665, 16'd1382, 16'd16171, 16'd3897, 16'd34706, 16'd55981});
	test_expansion(128'h9a6dc08735bc5183ef7082e986f248ac, {16'd25162, 16'd14249, 16'd51463, 16'd11198, 16'd16253, 16'd17236, 16'd4965, 16'd3428, 16'd28556, 16'd54193, 16'd13545, 16'd61981, 16'd39309, 16'd63529, 16'd43343, 16'd45192, 16'd56343, 16'd64422, 16'd61654, 16'd25521, 16'd42700, 16'd53689, 16'd52372, 16'd51926, 16'd26560, 16'd57940});
	test_expansion(128'he79c95be69f2ab10f3291d8256dbd781, {16'd16113, 16'd23058, 16'd38802, 16'd18920, 16'd44487, 16'd46860, 16'd1190, 16'd26188, 16'd1878, 16'd35699, 16'd30660, 16'd29119, 16'd63089, 16'd45816, 16'd19004, 16'd19406, 16'd45204, 16'd48012, 16'd14871, 16'd32717, 16'd17380, 16'd6219, 16'd9930, 16'd38808, 16'd14110, 16'd7286});
	test_expansion(128'h6b30e21f11eabb5dcdbe9b1a011372df, {16'd53002, 16'd56587, 16'd42931, 16'd22984, 16'd65387, 16'd44366, 16'd8410, 16'd59198, 16'd55519, 16'd59976, 16'd33421, 16'd51387, 16'd726, 16'd7030, 16'd990, 16'd60171, 16'd57656, 16'd41518, 16'd9662, 16'd6765, 16'd14844, 16'd65452, 16'd18033, 16'd6268, 16'd19669, 16'd15645});
	test_expansion(128'h7304b3b209faaa130497513b33037d24, {16'd63067, 16'd56320, 16'd8578, 16'd26725, 16'd12923, 16'd53602, 16'd3984, 16'd59935, 16'd25143, 16'd14922, 16'd26316, 16'd33417, 16'd40183, 16'd64089, 16'd31734, 16'd8374, 16'd35647, 16'd57390, 16'd23365, 16'd46605, 16'd3927, 16'd62164, 16'd51534, 16'd5748, 16'd54868, 16'd37945});
	test_expansion(128'h93c7a92a3b4664a73e5e0e2775c291af, {16'd50325, 16'd18864, 16'd45939, 16'd53164, 16'd23029, 16'd14053, 16'd64491, 16'd57730, 16'd52236, 16'd25586, 16'd61725, 16'd64796, 16'd2857, 16'd48200, 16'd15137, 16'd62086, 16'd48815, 16'd47248, 16'd27254, 16'd50990, 16'd50441, 16'd2630, 16'd56642, 16'd13042, 16'd38030, 16'd54792});
	test_expansion(128'hedd1fc34e7e87c41dc88c2ea9a833bd4, {16'd63822, 16'd27114, 16'd46141, 16'd41323, 16'd45164, 16'd63376, 16'd6340, 16'd51439, 16'd26814, 16'd3653, 16'd8343, 16'd26861, 16'd44920, 16'd37783, 16'd34449, 16'd63784, 16'd1024, 16'd16319, 16'd48097, 16'd60019, 16'd54214, 16'd8616, 16'd46325, 16'd27216, 16'd20051, 16'd48001});
	test_expansion(128'h2a59fd099326283b1a9122829b60f117, {16'd52116, 16'd29270, 16'd55040, 16'd37576, 16'd29621, 16'd847, 16'd54709, 16'd43609, 16'd56686, 16'd46433, 16'd46567, 16'd46859, 16'd31162, 16'd13851, 16'd42430, 16'd26004, 16'd65058, 16'd20348, 16'd40152, 16'd49648, 16'd41191, 16'd26929, 16'd47339, 16'd34611, 16'd58971, 16'd34190});
	test_expansion(128'h08b9ec8828cc527ac2a1d1188e85bcec, {16'd34460, 16'd63815, 16'd20095, 16'd13940, 16'd63247, 16'd30448, 16'd60172, 16'd52494, 16'd12644, 16'd39640, 16'd46217, 16'd37546, 16'd37594, 16'd16808, 16'd10184, 16'd43898, 16'd3752, 16'd49111, 16'd30306, 16'd24164, 16'd52271, 16'd59733, 16'd48619, 16'd50520, 16'd43185, 16'd33762});
	test_expansion(128'h91da556d1db475c2e72ed6e739c51989, {16'd1479, 16'd51066, 16'd11928, 16'd45678, 16'd22819, 16'd14440, 16'd38613, 16'd56533, 16'd17785, 16'd64544, 16'd16122, 16'd33368, 16'd51590, 16'd12539, 16'd65275, 16'd27455, 16'd44148, 16'd44449, 16'd50105, 16'd39717, 16'd21080, 16'd57200, 16'd7476, 16'd41433, 16'd11122, 16'd13990});
	test_expansion(128'hb14b96f29273578a808f54ce09f2d0e3, {16'd46386, 16'd21978, 16'd57118, 16'd41702, 16'd59559, 16'd52958, 16'd48479, 16'd36570, 16'd34122, 16'd15315, 16'd51210, 16'd53816, 16'd13909, 16'd13383, 16'd64336, 16'd24983, 16'd3877, 16'd38957, 16'd39012, 16'd48814, 16'd30980, 16'd12632, 16'd9976, 16'd32964, 16'd63740, 16'd30591});
	test_expansion(128'hb8302167478df35b11c773a12ca18ba7, {16'd59052, 16'd9895, 16'd58885, 16'd47632, 16'd1117, 16'd17347, 16'd49747, 16'd39219, 16'd38477, 16'd1263, 16'd22369, 16'd56571, 16'd58437, 16'd23686, 16'd33476, 16'd14389, 16'd63341, 16'd38867, 16'd35077, 16'd6950, 16'd41517, 16'd24396, 16'd40125, 16'd62788, 16'd61066, 16'd29152});
	test_expansion(128'h1234491e87ccf3fb1abb7f288a336749, {16'd16435, 16'd11948, 16'd1090, 16'd3904, 16'd42161, 16'd52519, 16'd54186, 16'd14182, 16'd16294, 16'd1205, 16'd53931, 16'd639, 16'd22332, 16'd54443, 16'd41039, 16'd761, 16'd46141, 16'd30776, 16'd38164, 16'd9610, 16'd23532, 16'd18655, 16'd56525, 16'd7630, 16'd9506, 16'd11742});
	test_expansion(128'hcc5d45da778eaf242350062bf99e0bb6, {16'd16137, 16'd36549, 16'd22491, 16'd59847, 16'd54596, 16'd23802, 16'd58859, 16'd59762, 16'd13653, 16'd17579, 16'd60436, 16'd11581, 16'd51930, 16'd38617, 16'd22393, 16'd40120, 16'd28065, 16'd62959, 16'd59203, 16'd64193, 16'd8430, 16'd61189, 16'd32859, 16'd58854, 16'd36969, 16'd56878});
	test_expansion(128'h373fe803ff27c60ae77b4b9f631eaf8a, {16'd894, 16'd57876, 16'd46545, 16'd17821, 16'd4490, 16'd60984, 16'd2522, 16'd58938, 16'd3153, 16'd8689, 16'd17984, 16'd13748, 16'd17049, 16'd3383, 16'd6384, 16'd14515, 16'd56701, 16'd3773, 16'd5663, 16'd20248, 16'd4637, 16'd49969, 16'd35524, 16'd49384, 16'd47305, 16'd18870});
	test_expansion(128'haea71feccdbc2ffcf5b10be0eda0f2c4, {16'd42423, 16'd2980, 16'd49700, 16'd27589, 16'd17252, 16'd48877, 16'd2802, 16'd60040, 16'd15956, 16'd40753, 16'd52473, 16'd11803, 16'd45415, 16'd59838, 16'd58344, 16'd6188, 16'd47484, 16'd32677, 16'd9491, 16'd28836, 16'd10720, 16'd5410, 16'd46063, 16'd6758, 16'd52075, 16'd5292});
	test_expansion(128'hf343cdf23bf83ab1868762986e1aebb1, {16'd2828, 16'd4974, 16'd59133, 16'd64779, 16'd52193, 16'd5369, 16'd30328, 16'd57049, 16'd29236, 16'd28222, 16'd27033, 16'd28126, 16'd48083, 16'd25418, 16'd57646, 16'd29684, 16'd33937, 16'd41488, 16'd49610, 16'd3859, 16'd33328, 16'd23615, 16'd38970, 16'd43673, 16'd38872, 16'd40663});
	test_expansion(128'h6a618c16fc90911cb2889942fb84c8f6, {16'd41382, 16'd21183, 16'd35276, 16'd43084, 16'd52385, 16'd5977, 16'd17353, 16'd26996, 16'd57711, 16'd9071, 16'd8683, 16'd17212, 16'd4203, 16'd32215, 16'd55363, 16'd61488, 16'd56663, 16'd18291, 16'd13512, 16'd13011, 16'd63387, 16'd27073, 16'd18342, 16'd49606, 16'd11869, 16'd34019});
	test_expansion(128'h8f47d080d267a9da00ec47f9abf4e4a9, {16'd46486, 16'd41218, 16'd32121, 16'd32026, 16'd63677, 16'd5402, 16'd57820, 16'd16994, 16'd44835, 16'd49864, 16'd1026, 16'd15986, 16'd44712, 16'd20853, 16'd28663, 16'd2396, 16'd24237, 16'd23411, 16'd30731, 16'd49817, 16'd20428, 16'd33874, 16'd45299, 16'd54141, 16'd21741, 16'd53285});
	test_expansion(128'h32ebc2799591c7655c62994b6a7dd7a9, {16'd7955, 16'd49272, 16'd61930, 16'd7260, 16'd41071, 16'd16192, 16'd57290, 16'd42301, 16'd17649, 16'd6584, 16'd37310, 16'd65288, 16'd58491, 16'd53395, 16'd20672, 16'd13943, 16'd15625, 16'd51393, 16'd23358, 16'd59644, 16'd3348, 16'd8831, 16'd29537, 16'd32802, 16'd35461, 16'd54871});
	test_expansion(128'h662df4568793e8130c23845495148e2f, {16'd22881, 16'd7438, 16'd33826, 16'd49783, 16'd37085, 16'd35304, 16'd40287, 16'd49449, 16'd19997, 16'd64354, 16'd47098, 16'd63077, 16'd22978, 16'd40894, 16'd16532, 16'd45897, 16'd10369, 16'd22064, 16'd3014, 16'd51759, 16'd9530, 16'd25369, 16'd49984, 16'd16716, 16'd32406, 16'd59225});
	test_expansion(128'he720a25406b14543d72c3f102870e38d, {16'd27103, 16'd5023, 16'd43915, 16'd8495, 16'd6172, 16'd2612, 16'd31177, 16'd62687, 16'd37334, 16'd52116, 16'd3401, 16'd37627, 16'd1074, 16'd55406, 16'd29129, 16'd5028, 16'd37560, 16'd8367, 16'd56716, 16'd48213, 16'd52994, 16'd54817, 16'd54052, 16'd33624, 16'd57555, 16'd3976});
	test_expansion(128'h713a5efa941dd3edc2f66b5762f3bcef, {16'd28562, 16'd45534, 16'd54081, 16'd8085, 16'd64062, 16'd17527, 16'd56128, 16'd46545, 16'd47798, 16'd22024, 16'd32202, 16'd52860, 16'd48990, 16'd61197, 16'd55019, 16'd62477, 16'd62729, 16'd31999, 16'd53464, 16'd64100, 16'd38965, 16'd64728, 16'd39525, 16'd43806, 16'd16302, 16'd4379});
	test_expansion(128'h6742308a84db07c27d3d1444fed15244, {16'd21507, 16'd9421, 16'd2370, 16'd58235, 16'd65306, 16'd26770, 16'd28742, 16'd24284, 16'd25202, 16'd58942, 16'd38433, 16'd2354, 16'd3227, 16'd60700, 16'd33100, 16'd1832, 16'd57970, 16'd20327, 16'd64926, 16'd31560, 16'd2168, 16'd48495, 16'd36302, 16'd18801, 16'd57099, 16'd6501});
	test_expansion(128'h28c4cfd0f54b112a54363fd63a330a53, {16'd39513, 16'd8889, 16'd27361, 16'd42568, 16'd48939, 16'd26312, 16'd59748, 16'd39871, 16'd42947, 16'd56193, 16'd52984, 16'd8169, 16'd15301, 16'd50768, 16'd27541, 16'd25291, 16'd37998, 16'd59227, 16'd57894, 16'd56608, 16'd32450, 16'd58961, 16'd39176, 16'd10521, 16'd46092, 16'd35755});
	test_expansion(128'hf0b68a83b415a824088f2aacb0c1df7e, {16'd28011, 16'd15659, 16'd59630, 16'd42045, 16'd44957, 16'd18990, 16'd56789, 16'd41942, 16'd58736, 16'd30290, 16'd53789, 16'd14619, 16'd43607, 16'd12460, 16'd48682, 16'd55665, 16'd4888, 16'd58037, 16'd44640, 16'd40241, 16'd21176, 16'd5013, 16'd16813, 16'd29875, 16'd55524, 16'd47988});
	test_expansion(128'h2b7cc67f4cc7521ac4d4043be9078663, {16'd60016, 16'd63134, 16'd30790, 16'd38831, 16'd10011, 16'd56067, 16'd42110, 16'd65019, 16'd46326, 16'd43205, 16'd49875, 16'd48190, 16'd40822, 16'd50660, 16'd27847, 16'd59132, 16'd64111, 16'd10647, 16'd26977, 16'd12495, 16'd33728, 16'd8171, 16'd8087, 16'd3912, 16'd4557, 16'd43129});
	test_expansion(128'hf4de4891a750e50fcf6f2cd165fe7a15, {16'd63542, 16'd6460, 16'd24530, 16'd50626, 16'd16300, 16'd43433, 16'd13050, 16'd26400, 16'd12432, 16'd18768, 16'd61716, 16'd19108, 16'd28457, 16'd2172, 16'd42112, 16'd26132, 16'd10640, 16'd38097, 16'd5191, 16'd53694, 16'd2010, 16'd18596, 16'd36092, 16'd2936, 16'd24861, 16'd53069});
	test_expansion(128'h0e75de7d111537b5ef33e20902dfbc50, {16'd52383, 16'd54671, 16'd9077, 16'd5863, 16'd62635, 16'd44515, 16'd26687, 16'd3716, 16'd55216, 16'd60508, 16'd58930, 16'd23298, 16'd53556, 16'd11913, 16'd18529, 16'd51783, 16'd55310, 16'd22943, 16'd8716, 16'd47785, 16'd2424, 16'd48543, 16'd776, 16'd62011, 16'd45764, 16'd54690});
	test_expansion(128'hddc81187e23157e5163bb697c98864b9, {16'd25616, 16'd35552, 16'd38986, 16'd54628, 16'd42431, 16'd33573, 16'd4825, 16'd9913, 16'd44536, 16'd55315, 16'd39051, 16'd5666, 16'd2835, 16'd44467, 16'd12077, 16'd12720, 16'd50942, 16'd55251, 16'd12734, 16'd36673, 16'd45633, 16'd42145, 16'd49373, 16'd20232, 16'd58103, 16'd16050});
	test_expansion(128'he8008eef6227f30f9eb07ad2f9bdc24c, {16'd10832, 16'd16795, 16'd53364, 16'd62447, 16'd20865, 16'd18606, 16'd63766, 16'd27138, 16'd22036, 16'd24928, 16'd32259, 16'd46027, 16'd13937, 16'd56678, 16'd16049, 16'd10693, 16'd19180, 16'd46133, 16'd10654, 16'd39542, 16'd47409, 16'd62705, 16'd63560, 16'd1154, 16'd11554, 16'd4283});
	test_expansion(128'h95ae88fc1c25edfb570d7ca32a681145, {16'd57777, 16'd11100, 16'd10486, 16'd45610, 16'd29266, 16'd21273, 16'd32595, 16'd65036, 16'd48760, 16'd41822, 16'd12592, 16'd52004, 16'd4014, 16'd32059, 16'd40797, 16'd42808, 16'd62721, 16'd18653, 16'd53334, 16'd51941, 16'd8848, 16'd25388, 16'd53266, 16'd32855, 16'd56593, 16'd64923});
	test_expansion(128'h5db83e91e83857efd86f14d97eb819e7, {16'd55971, 16'd26514, 16'd38357, 16'd27356, 16'd35936, 16'd6844, 16'd15562, 16'd31204, 16'd58030, 16'd12511, 16'd52367, 16'd48542, 16'd24626, 16'd39545, 16'd35359, 16'd36692, 16'd47586, 16'd14630, 16'd3150, 16'd41480, 16'd8837, 16'd21554, 16'd47120, 16'd53050, 16'd35163, 16'd7575});
	test_expansion(128'h2e0d0c5fa976c261524fd9f55197eb0b, {16'd31966, 16'd60624, 16'd61764, 16'd12961, 16'd20385, 16'd46814, 16'd32986, 16'd36147, 16'd57303, 16'd26216, 16'd33613, 16'd53402, 16'd46145, 16'd26432, 16'd58340, 16'd42558, 16'd1849, 16'd63451, 16'd53714, 16'd29411, 16'd9152, 16'd16282, 16'd7000, 16'd25379, 16'd61677, 16'd3091});
	test_expansion(128'h95bc6cb29b52e3d2045409f7684f736e, {16'd5352, 16'd50326, 16'd54395, 16'd28063, 16'd52933, 16'd27791, 16'd31400, 16'd37753, 16'd60902, 16'd6767, 16'd2029, 16'd5336, 16'd19132, 16'd21259, 16'd10249, 16'd63591, 16'd50094, 16'd19863, 16'd52205, 16'd58913, 16'd27760, 16'd47908, 16'd38832, 16'd34574, 16'd26466, 16'd4869});
	test_expansion(128'h138898736595547fefca0a9b8f5f5451, {16'd59888, 16'd13925, 16'd16746, 16'd37169, 16'd31176, 16'd13165, 16'd45776, 16'd18665, 16'd46619, 16'd24743, 16'd58621, 16'd59292, 16'd37428, 16'd41753, 16'd52195, 16'd14855, 16'd61330, 16'd51068, 16'd13253, 16'd25351, 16'd65467, 16'd20740, 16'd26079, 16'd31220, 16'd57044, 16'd8438});
	test_expansion(128'hd3cc3f2fd68cd50f3728b50fd8588ba8, {16'd51096, 16'd34706, 16'd34837, 16'd60505, 16'd45960, 16'd36373, 16'd17435, 16'd40598, 16'd15445, 16'd45885, 16'd9619, 16'd14201, 16'd54267, 16'd27851, 16'd58819, 16'd35860, 16'd49778, 16'd62352, 16'd20885, 16'd50442, 16'd29642, 16'd63433, 16'd31770, 16'd17575, 16'd45099, 16'd11693});
	test_expansion(128'heeec4c9464c18c53d6675b018614c1c3, {16'd23753, 16'd62887, 16'd46376, 16'd63889, 16'd23083, 16'd49730, 16'd51177, 16'd41172, 16'd47747, 16'd46729, 16'd55721, 16'd29986, 16'd47701, 16'd16568, 16'd6478, 16'd35697, 16'd10988, 16'd65382, 16'd11521, 16'd46989, 16'd10532, 16'd52963, 16'd57092, 16'd55098, 16'd42593, 16'd44079});
	test_expansion(128'h41afb48f5383d230de8ac9d12087ad50, {16'd37393, 16'd7456, 16'd36631, 16'd40106, 16'd13177, 16'd11642, 16'd50364, 16'd24547, 16'd40922, 16'd41380, 16'd10913, 16'd8562, 16'd27473, 16'd33481, 16'd2231, 16'd31800, 16'd13447, 16'd19954, 16'd39683, 16'd36582, 16'd31183, 16'd40807, 16'd4632, 16'd16103, 16'd29414, 16'd39451});
	test_expansion(128'h2ce6354bc364e2e70f6a50a898c1616a, {16'd65125, 16'd59137, 16'd18333, 16'd40014, 16'd15347, 16'd42654, 16'd49561, 16'd60997, 16'd21000, 16'd42356, 16'd56124, 16'd22306, 16'd17006, 16'd43799, 16'd15960, 16'd52533, 16'd6941, 16'd51752, 16'd4397, 16'd15921, 16'd37373, 16'd37133, 16'd58667, 16'd2751, 16'd39928, 16'd56359});
	test_expansion(128'hc4a5e841dac2b02b622c03c14d4d9c07, {16'd18274, 16'd14975, 16'd16470, 16'd59035, 16'd38459, 16'd63607, 16'd38627, 16'd17346, 16'd8352, 16'd38216, 16'd48155, 16'd25953, 16'd26371, 16'd9605, 16'd5724, 16'd41702, 16'd5508, 16'd43047, 16'd20267, 16'd60714, 16'd22071, 16'd54599, 16'd55595, 16'd46110, 16'd12907, 16'd7819});
	test_expansion(128'hf222c0b9ba9326b55a7a0d836cdce84b, {16'd57826, 16'd56255, 16'd23724, 16'd47065, 16'd24721, 16'd31295, 16'd60863, 16'd8350, 16'd46546, 16'd25397, 16'd29983, 16'd36581, 16'd34024, 16'd21591, 16'd17251, 16'd15415, 16'd63351, 16'd46628, 16'd65228, 16'd7312, 16'd2933, 16'd42, 16'd42515, 16'd42788, 16'd3162, 16'd24993});
	test_expansion(128'he3018cce9fefd37db8da141c2babaf3f, {16'd33318, 16'd65084, 16'd3736, 16'd62479, 16'd42493, 16'd63164, 16'd40265, 16'd4767, 16'd48657, 16'd22240, 16'd28015, 16'd56685, 16'd4110, 16'd8747, 16'd3794, 16'd13514, 16'd15742, 16'd9820, 16'd39591, 16'd13798, 16'd49533, 16'd48008, 16'd49039, 16'd62030, 16'd48391, 16'd59704});
	test_expansion(128'hdd62d18921953f061e6a73cb4a8f3130, {16'd22070, 16'd60164, 16'd43928, 16'd3493, 16'd32215, 16'd57829, 16'd9608, 16'd56634, 16'd41139, 16'd44170, 16'd28850, 16'd7260, 16'd32887, 16'd18778, 16'd56755, 16'd1384, 16'd16455, 16'd8310, 16'd63564, 16'd34975, 16'd58447, 16'd120, 16'd40518, 16'd8450, 16'd25714, 16'd38258});
	test_expansion(128'hcab1782a07a2e34d3f112b8bc6b7e2d5, {16'd61899, 16'd32594, 16'd59196, 16'd12886, 16'd30652, 16'd36387, 16'd20638, 16'd51634, 16'd33394, 16'd55158, 16'd21801, 16'd35379, 16'd61534, 16'd13495, 16'd28238, 16'd39083, 16'd47505, 16'd51078, 16'd37620, 16'd37692, 16'd31866, 16'd29818, 16'd25536, 16'd11962, 16'd62199, 16'd9571});
	test_expansion(128'hd91e81c16010516ab9bbc7f6cd148394, {16'd61131, 16'd7260, 16'd1942, 16'd27754, 16'd16627, 16'd45374, 16'd65472, 16'd44190, 16'd55706, 16'd27601, 16'd25560, 16'd41019, 16'd27138, 16'd48512, 16'd59189, 16'd25457, 16'd3969, 16'd13855, 16'd51414, 16'd9679, 16'd26900, 16'd8175, 16'd2377, 16'd44744, 16'd638, 16'd55004});
	test_expansion(128'h74d874a7ad2d09a7e8411fdbc0aeef7c, {16'd18271, 16'd41005, 16'd46366, 16'd32063, 16'd59833, 16'd55741, 16'd32369, 16'd49183, 16'd9596, 16'd19752, 16'd6873, 16'd2266, 16'd63734, 16'd58276, 16'd54870, 16'd13860, 16'd27967, 16'd38464, 16'd26372, 16'd13820, 16'd46560, 16'd10804, 16'd16264, 16'd40195, 16'd44387, 16'd8850});
	test_expansion(128'h70f6a97d590f0caafbb83f49db365bfe, {16'd16521, 16'd6584, 16'd34352, 16'd47248, 16'd1016, 16'd44222, 16'd31268, 16'd58698, 16'd16588, 16'd32922, 16'd27021, 16'd18963, 16'd54054, 16'd38821, 16'd16722, 16'd30791, 16'd41335, 16'd2404, 16'd8746, 16'd25909, 16'd14686, 16'd19704, 16'd62063, 16'd34385, 16'd22720, 16'd45900});
	test_expansion(128'h6d5bfe1235da1f0690cc5113f555760a, {16'd6884, 16'd6298, 16'd37323, 16'd4517, 16'd37935, 16'd57136, 16'd18610, 16'd6910, 16'd37280, 16'd42188, 16'd38036, 16'd48614, 16'd18966, 16'd4864, 16'd36434, 16'd2782, 16'd43388, 16'd64232, 16'd65408, 16'd38935, 16'd49242, 16'd57665, 16'd56206, 16'd46002, 16'd1255, 16'd30189});
	test_expansion(128'hbb581d2a005ae0fb430dd309e7ecafa2, {16'd59618, 16'd65139, 16'd49903, 16'd2781, 16'd59064, 16'd59980, 16'd7336, 16'd5031, 16'd52510, 16'd62173, 16'd63438, 16'd64941, 16'd55313, 16'd56650, 16'd39563, 16'd50442, 16'd6933, 16'd62273, 16'd62942, 16'd52924, 16'd58047, 16'd37123, 16'd15237, 16'd30476, 16'd1274, 16'd5580});
	test_expansion(128'h357cbff4c30b59436bf1233de68bbca4, {16'd36143, 16'd41269, 16'd7015, 16'd27165, 16'd5533, 16'd39602, 16'd24229, 16'd14881, 16'd59054, 16'd4386, 16'd56605, 16'd8150, 16'd57942, 16'd23471, 16'd8992, 16'd41606, 16'd1525, 16'd15870, 16'd6145, 16'd35107, 16'd4748, 16'd35236, 16'd26333, 16'd32536, 16'd40626, 16'd24463});
	test_expansion(128'hb9fba7f2f6e57930fc079130e5a3802f, {16'd9536, 16'd52250, 16'd60754, 16'd37326, 16'd37911, 16'd22039, 16'd51643, 16'd12615, 16'd38142, 16'd39915, 16'd49292, 16'd7292, 16'd53998, 16'd50477, 16'd57746, 16'd50649, 16'd51388, 16'd5037, 16'd9338, 16'd44481, 16'd57552, 16'd56709, 16'd10009, 16'd43675, 16'd31118, 16'd18287});
	test_expansion(128'h0f2b4bd5a053f1aa42e8b41b6c751a08, {16'd32626, 16'd53581, 16'd15726, 16'd38323, 16'd15597, 16'd40466, 16'd3074, 16'd46401, 16'd28319, 16'd33184, 16'd16653, 16'd34656, 16'd1934, 16'd50013, 16'd62396, 16'd64875, 16'd51549, 16'd61903, 16'd13206, 16'd6598, 16'd59054, 16'd13365, 16'd2988, 16'd11931, 16'd5942, 16'd16488});
	test_expansion(128'h55dfbed3956c2f147731557de03598f0, {16'd24158, 16'd35621, 16'd5100, 16'd19457, 16'd42992, 16'd48417, 16'd45810, 16'd64965, 16'd12867, 16'd53062, 16'd59343, 16'd64333, 16'd51965, 16'd27352, 16'd17439, 16'd52235, 16'd35573, 16'd51088, 16'd11756, 16'd51117, 16'd30351, 16'd54894, 16'd15441, 16'd12947, 16'd32361, 16'd36175});
	test_expansion(128'hab5c6a42085d2b4a409051011a4a4f4a, {16'd51995, 16'd58494, 16'd56795, 16'd61047, 16'd30728, 16'd37195, 16'd62448, 16'd27901, 16'd40915, 16'd59556, 16'd21332, 16'd50566, 16'd4588, 16'd2718, 16'd12914, 16'd41100, 16'd42309, 16'd30549, 16'd62293, 16'd23604, 16'd32915, 16'd29164, 16'd9586, 16'd23995, 16'd48668, 16'd61247});
	test_expansion(128'h878e3cc9ca8ccebae822d043de0563d6, {16'd27406, 16'd10831, 16'd61968, 16'd6721, 16'd21623, 16'd53838, 16'd31289, 16'd59280, 16'd16853, 16'd28003, 16'd18206, 16'd10134, 16'd37592, 16'd9249, 16'd56624, 16'd47291, 16'd41713, 16'd29901, 16'd52291, 16'd18043, 16'd50722, 16'd441, 16'd3789, 16'd34789, 16'd65052, 16'd24562});
	test_expansion(128'haf62bc0fda8582c07a1ecd17afdac3bc, {16'd17469, 16'd59744, 16'd6287, 16'd48767, 16'd32381, 16'd9820, 16'd29431, 16'd49264, 16'd35613, 16'd21211, 16'd31368, 16'd58770, 16'd36575, 16'd31712, 16'd11945, 16'd23645, 16'd64972, 16'd53537, 16'd24309, 16'd29797, 16'd56302, 16'd39399, 16'd57738, 16'd32922, 16'd44927, 16'd3129});
	test_expansion(128'h5201a2625b24103260f6720ee0fca598, {16'd6704, 16'd2714, 16'd61318, 16'd11486, 16'd61340, 16'd43980, 16'd20698, 16'd4113, 16'd43563, 16'd54010, 16'd54432, 16'd48193, 16'd21795, 16'd30526, 16'd52666, 16'd49050, 16'd54180, 16'd53202, 16'd1721, 16'd18209, 16'd22904, 16'd56889, 16'd31845, 16'd10021, 16'd51525, 16'd10629});
	test_expansion(128'h826d91b17cecb455681f12fdda0015a1, {16'd36040, 16'd22692, 16'd3281, 16'd58554, 16'd48842, 16'd34858, 16'd11855, 16'd46052, 16'd44482, 16'd45205, 16'd12347, 16'd18184, 16'd50518, 16'd27495, 16'd32908, 16'd41566, 16'd40823, 16'd21905, 16'd12281, 16'd15356, 16'd54009, 16'd27130, 16'd35988, 16'd19220, 16'd5688, 16'd30993});
	test_expansion(128'hcec144b1f48b684dd5666faec935fca3, {16'd28190, 16'd37993, 16'd9092, 16'd40322, 16'd49399, 16'd3371, 16'd22183, 16'd7281, 16'd2362, 16'd45927, 16'd17271, 16'd8865, 16'd30662, 16'd25678, 16'd48748, 16'd6901, 16'd14156, 16'd55075, 16'd3771, 16'd28939, 16'd18065, 16'd48532, 16'd15655, 16'd62556, 16'd47918, 16'd10893});
	test_expansion(128'heb9981abca844fcc6f626fec4e7fb7c8, {16'd29600, 16'd48803, 16'd14865, 16'd34706, 16'd6565, 16'd59387, 16'd4600, 16'd15621, 16'd51437, 16'd35933, 16'd10859, 16'd5745, 16'd16643, 16'd22716, 16'd17833, 16'd34810, 16'd61887, 16'd8444, 16'd51855, 16'd15702, 16'd52383, 16'd7246, 16'd55461, 16'd15996, 16'd26901, 16'd290});
	test_expansion(128'h433d4a4ca585bc798d1ea2fa616f2154, {16'd47487, 16'd3267, 16'd17623, 16'd10935, 16'd60419, 16'd35899, 16'd59111, 16'd36601, 16'd8295, 16'd49411, 16'd18810, 16'd20991, 16'd45598, 16'd46456, 16'd24063, 16'd3809, 16'd16328, 16'd27876, 16'd15750, 16'd24075, 16'd1634, 16'd53566, 16'd47871, 16'd12961, 16'd17708, 16'd13045});
	test_expansion(128'h3a02e4b7e79c040d86240ef8dacd2f16, {16'd17508, 16'd57348, 16'd11750, 16'd21952, 16'd63093, 16'd32218, 16'd19322, 16'd20742, 16'd39483, 16'd20250, 16'd61697, 16'd53803, 16'd9313, 16'd14001, 16'd9621, 16'd43541, 16'd11275, 16'd12271, 16'd51274, 16'd36380, 16'd7431, 16'd22166, 16'd58959, 16'd10662, 16'd64713, 16'd62214});
	test_expansion(128'h780d9c37ffaa75d4c38cd9dd2ec724de, {16'd24395, 16'd36992, 16'd31538, 16'd3878, 16'd20053, 16'd54984, 16'd19858, 16'd10246, 16'd33250, 16'd21558, 16'd4683, 16'd18250, 16'd60961, 16'd21583, 16'd20657, 16'd19887, 16'd30296, 16'd62829, 16'd41640, 16'd54294, 16'd11227, 16'd21140, 16'd48992, 16'd4184, 16'd424, 16'd56424});
	test_expansion(128'h3dad4431da19539df4d3d8bde9fc0405, {16'd21070, 16'd58453, 16'd13564, 16'd10696, 16'd22562, 16'd5116, 16'd37211, 16'd21104, 16'd31785, 16'd35611, 16'd32341, 16'd63278, 16'd64852, 16'd25223, 16'd59715, 16'd59128, 16'd36494, 16'd15381, 16'd57644, 16'd2419, 16'd6414, 16'd8166, 16'd39074, 16'd48659, 16'd29936, 16'd10967});
	test_expansion(128'h96b584293a2f79ab522045f0f5a41200, {16'd31385, 16'd55197, 16'd34294, 16'd4917, 16'd10332, 16'd16306, 16'd27274, 16'd17755, 16'd26747, 16'd54562, 16'd64945, 16'd24316, 16'd34910, 16'd17375, 16'd42644, 16'd13975, 16'd38878, 16'd54939, 16'd9679, 16'd43569, 16'd15856, 16'd4032, 16'd3793, 16'd20124, 16'd6341, 16'd13147});
	test_expansion(128'h152147f9142af30bbd3eefe13feef993, {16'd53425, 16'd5117, 16'd50066, 16'd61545, 16'd51315, 16'd24315, 16'd45545, 16'd9348, 16'd32893, 16'd62216, 16'd22883, 16'd8763, 16'd50509, 16'd53280, 16'd51138, 16'd29588, 16'd62178, 16'd7533, 16'd37835, 16'd3826, 16'd59076, 16'd14899, 16'd42311, 16'd27848, 16'd22938, 16'd58659});
	test_expansion(128'h424898ff859ac86c536cea8c2b769734, {16'd43834, 16'd8088, 16'd39919, 16'd34222, 16'd1881, 16'd822, 16'd36891, 16'd25098, 16'd41174, 16'd11369, 16'd52132, 16'd1245, 16'd23167, 16'd48179, 16'd59723, 16'd49338, 16'd34147, 16'd8415, 16'd45171, 16'd33963, 16'd5663, 16'd63264, 16'd20963, 16'd8651, 16'd6751, 16'd26517});
	test_expansion(128'h73770d4f2e5b51f1b94bd5bfe94ef633, {16'd5701, 16'd13398, 16'd23055, 16'd14555, 16'd16308, 16'd19961, 16'd57307, 16'd9989, 16'd24111, 16'd56433, 16'd23541, 16'd5926, 16'd24127, 16'd55821, 16'd21460, 16'd21155, 16'd3451, 16'd12940, 16'd56217, 16'd5848, 16'd11699, 16'd56509, 16'd23217, 16'd19677, 16'd32748, 16'd37798});
	test_expansion(128'h1ead9227661f047d85bf4154faef499b, {16'd38049, 16'd42774, 16'd62663, 16'd41952, 16'd27585, 16'd64843, 16'd39659, 16'd48538, 16'd54451, 16'd1291, 16'd8340, 16'd6694, 16'd56163, 16'd9669, 16'd59789, 16'd36096, 16'd23176, 16'd25235, 16'd23084, 16'd36767, 16'd31063, 16'd23001, 16'd7349, 16'd2874, 16'd3127, 16'd543});
	test_expansion(128'h2d697a395fdd6a909de34c77a8c43a19, {16'd60084, 16'd2442, 16'd33017, 16'd32699, 16'd158, 16'd55264, 16'd20701, 16'd52545, 16'd12085, 16'd8307, 16'd8273, 16'd52309, 16'd15941, 16'd25537, 16'd37079, 16'd45551, 16'd2679, 16'd23566, 16'd21402, 16'd7719, 16'd30698, 16'd33899, 16'd990, 16'd32557, 16'd233, 16'd19608});
	test_expansion(128'hd4e9710420b5312d36ed18cd8b842090, {16'd21094, 16'd29557, 16'd6512, 16'd60649, 16'd52033, 16'd38476, 16'd32348, 16'd60900, 16'd32134, 16'd63301, 16'd27823, 16'd1644, 16'd10381, 16'd10097, 16'd37408, 16'd3605, 16'd33842, 16'd56240, 16'd4954, 16'd32121, 16'd45743, 16'd61788, 16'd43509, 16'd22482, 16'd30683, 16'd48850});
	test_expansion(128'ha9ba9af815727fe7c1379a808d049051, {16'd42174, 16'd43133, 16'd64826, 16'd23411, 16'd22706, 16'd28155, 16'd28645, 16'd40886, 16'd52130, 16'd53910, 16'd14615, 16'd57073, 16'd48266, 16'd59321, 16'd57894, 16'd49223, 16'd45800, 16'd42428, 16'd18775, 16'd55307, 16'd6663, 16'd61439, 16'd51284, 16'd29172, 16'd42685, 16'd51985});
	test_expansion(128'h5176b0103f7e947ee26fbbd2c49ebe95, {16'd59048, 16'd61411, 16'd64139, 16'd32845, 16'd45670, 16'd26060, 16'd63984, 16'd20670, 16'd44369, 16'd21546, 16'd22800, 16'd51392, 16'd29398, 16'd56778, 16'd35694, 16'd21074, 16'd43289, 16'd34246, 16'd42373, 16'd53267, 16'd20220, 16'd57914, 16'd45714, 16'd33268, 16'd4802, 16'd6957});
	test_expansion(128'hbcc64036e22b420289697328f5a094c6, {16'd47077, 16'd46037, 16'd46178, 16'd57262, 16'd5979, 16'd14138, 16'd8629, 16'd64780, 16'd28177, 16'd56895, 16'd64945, 16'd14105, 16'd57653, 16'd377, 16'd6267, 16'd19120, 16'd56963, 16'd63027, 16'd23490, 16'd55513, 16'd15265, 16'd52332, 16'd41363, 16'd44969, 16'd39565, 16'd37271});
	test_expansion(128'hcf36fc45b60a0b94fcb97d49b8c9556d, {16'd20341, 16'd51770, 16'd32269, 16'd29903, 16'd43758, 16'd29484, 16'd7743, 16'd64843, 16'd13549, 16'd13314, 16'd6846, 16'd29702, 16'd36381, 16'd29284, 16'd49794, 16'd55636, 16'd38507, 16'd10672, 16'd56968, 16'd60004, 16'd26411, 16'd17519, 16'd30178, 16'd57205, 16'd44579, 16'd10140});
	test_expansion(128'h748cc48775b59daecc8abbe97acc0358, {16'd27144, 16'd3556, 16'd15505, 16'd29755, 16'd50605, 16'd55338, 16'd15143, 16'd4863, 16'd1323, 16'd2365, 16'd52375, 16'd27840, 16'd22958, 16'd42355, 16'd20345, 16'd27602, 16'd20817, 16'd38055, 16'd362, 16'd52017, 16'd24790, 16'd40589, 16'd55363, 16'd16566, 16'd11409, 16'd44635});
	test_expansion(128'ha5fe725232d849b69b7529ea6d42237c, {16'd16983, 16'd9446, 16'd50588, 16'd36155, 16'd8772, 16'd49969, 16'd14491, 16'd16078, 16'd59862, 16'd36497, 16'd4868, 16'd13998, 16'd63648, 16'd59393, 16'd12825, 16'd14754, 16'd41201, 16'd24648, 16'd43534, 16'd12315, 16'd2981, 16'd45289, 16'd51854, 16'd11769, 16'd21275, 16'd46228});
	test_expansion(128'h2a35c6de153388d293d48a31aded4341, {16'd24065, 16'd62531, 16'd62299, 16'd47695, 16'd3699, 16'd33633, 16'd64956, 16'd19027, 16'd52594, 16'd47974, 16'd4273, 16'd45907, 16'd4498, 16'd38560, 16'd3250, 16'd9319, 16'd34014, 16'd20921, 16'd31870, 16'd40366, 16'd35818, 16'd19585, 16'd57431, 16'd51589, 16'd48924, 16'd31791});
	test_expansion(128'hb12a43d295565cab373218c4f5c9fb62, {16'd5913, 16'd33228, 16'd55406, 16'd27388, 16'd64455, 16'd36568, 16'd6391, 16'd56647, 16'd40146, 16'd48409, 16'd59799, 16'd10337, 16'd32660, 16'd31395, 16'd18001, 16'd42617, 16'd62687, 16'd31765, 16'd58624, 16'd61159, 16'd52431, 16'd11559, 16'd18449, 16'd52184, 16'd45319, 16'd34829});
	test_expansion(128'h208c7e12313a5cbad35f14af1fa32d86, {16'd41918, 16'd22100, 16'd29329, 16'd11920, 16'd40763, 16'd43539, 16'd65064, 16'd47274, 16'd63215, 16'd51330, 16'd41958, 16'd29781, 16'd25368, 16'd61983, 16'd33771, 16'd38012, 16'd27188, 16'd16288, 16'd11478, 16'd15970, 16'd45919, 16'd9771, 16'd28546, 16'd56185, 16'd17918, 16'd62815});
	test_expansion(128'h6ef9a2c3f1a2abf8a301573bb003c48a, {16'd46248, 16'd12806, 16'd59544, 16'd29336, 16'd8732, 16'd40704, 16'd11043, 16'd22898, 16'd59148, 16'd49384, 16'd26813, 16'd11554, 16'd60358, 16'd56522, 16'd57134, 16'd994, 16'd49250, 16'd49578, 16'd46148, 16'd62899, 16'd9584, 16'd7167, 16'd25989, 16'd12134, 16'd3192, 16'd22331});
	test_expansion(128'h5648df8e3ce0f58683de1c0428679996, {16'd14965, 16'd57406, 16'd24888, 16'd33806, 16'd32928, 16'd9900, 16'd23009, 16'd11143, 16'd49495, 16'd8465, 16'd214, 16'd49906, 16'd33923, 16'd3287, 16'd24106, 16'd7490, 16'd10655, 16'd19559, 16'd11809, 16'd2326, 16'd11747, 16'd51933, 16'd6567, 16'd44328, 16'd44452, 16'd57741});
	test_expansion(128'h24f0a86454e40a8cd98021f0d0d33c34, {16'd9222, 16'd7803, 16'd43434, 16'd45581, 16'd38592, 16'd27958, 16'd20106, 16'd7775, 16'd43673, 16'd37943, 16'd5695, 16'd476, 16'd57844, 16'd23872, 16'd3865, 16'd17384, 16'd17637, 16'd33509, 16'd55615, 16'd3353, 16'd13066, 16'd50871, 16'd45677, 16'd36344, 16'd7690, 16'd15339});
	test_expansion(128'h6de3fb2e825cf596e2fddba5f6e2811a, {16'd1369, 16'd12543, 16'd48631, 16'd31967, 16'd12157, 16'd2723, 16'd13502, 16'd14997, 16'd46152, 16'd8943, 16'd13950, 16'd50, 16'd63503, 16'd38398, 16'd24221, 16'd3157, 16'd57879, 16'd51072, 16'd34357, 16'd14036, 16'd4506, 16'd8925, 16'd14278, 16'd26088, 16'd18849, 16'd19595});
	test_expansion(128'hedfac50abbf747d14b89d45c84585382, {16'd9809, 16'd42553, 16'd44672, 16'd62595, 16'd9322, 16'd61299, 16'd40311, 16'd49731, 16'd5261, 16'd41123, 16'd30292, 16'd27455, 16'd28750, 16'd27429, 16'd20417, 16'd17336, 16'd21667, 16'd20929, 16'd48092, 16'd14408, 16'd32256, 16'd33796, 16'd9097, 16'd54574, 16'd49385, 16'd25128});
	test_expansion(128'h668edfbab160c248b956eecfbb40f260, {16'd17651, 16'd28025, 16'd1149, 16'd7848, 16'd4238, 16'd15946, 16'd2882, 16'd12831, 16'd5353, 16'd62419, 16'd38787, 16'd62888, 16'd21231, 16'd19724, 16'd16252, 16'd27704, 16'd9851, 16'd29485, 16'd64166, 16'd25132, 16'd28547, 16'd1852, 16'd4489, 16'd43090, 16'd23643, 16'd19823});
	test_expansion(128'h43bcbb6a8a0536e21af6c407b90e518b, {16'd34317, 16'd6548, 16'd48050, 16'd19933, 16'd35720, 16'd30649, 16'd51965, 16'd8216, 16'd7295, 16'd14195, 16'd34498, 16'd951, 16'd42937, 16'd33665, 16'd3397, 16'd33223, 16'd15705, 16'd9183, 16'd54190, 16'd29246, 16'd14678, 16'd6378, 16'd30336, 16'd32471, 16'd13852, 16'd49126});
	test_expansion(128'hec9c83c48c0a5e3c8ba242c76812950d, {16'd2506, 16'd37161, 16'd11165, 16'd20361, 16'd33547, 16'd52182, 16'd56647, 16'd2290, 16'd45681, 16'd42892, 16'd13100, 16'd59655, 16'd5644, 16'd6380, 16'd6530, 16'd63101, 16'd51849, 16'd45761, 16'd51569, 16'd60397, 16'd46668, 16'd9033, 16'd61595, 16'd8205, 16'd64110, 16'd61650});
	test_expansion(128'h74dc945f18e716767d989d5a03c7b8c6, {16'd54, 16'd64003, 16'd38940, 16'd46074, 16'd47790, 16'd41439, 16'd25484, 16'd33739, 16'd9839, 16'd6509, 16'd25839, 16'd10324, 16'd4827, 16'd25606, 16'd29309, 16'd52873, 16'd22808, 16'd65400, 16'd59644, 16'd48384, 16'd28000, 16'd44074, 16'd38981, 16'd23612, 16'd36910, 16'd34679});
	test_expansion(128'hd8b7fe4b263c82080260f99a6b4021d9, {16'd43097, 16'd14518, 16'd6999, 16'd12226, 16'd17478, 16'd60380, 16'd6855, 16'd6898, 16'd45370, 16'd53101, 16'd18934, 16'd14870, 16'd32525, 16'd34951, 16'd7609, 16'd481, 16'd17426, 16'd51835, 16'd13536, 16'd12340, 16'd3655, 16'd1235, 16'd39929, 16'd34335, 16'd55165, 16'd61402});
	test_expansion(128'hd8cc18783655cdf82434f143256570aa, {16'd41962, 16'd2429, 16'd3638, 16'd48951, 16'd48521, 16'd36868, 16'd47241, 16'd65289, 16'd27273, 16'd12890, 16'd49892, 16'd1625, 16'd26564, 16'd37316, 16'd55610, 16'd17870, 16'd49306, 16'd56446, 16'd11476, 16'd17486, 16'd19693, 16'd40499, 16'd30585, 16'd57899, 16'd35850, 16'd5729});
	test_expansion(128'h60274f43d19e2fdfdd65e36542f43a32, {16'd55129, 16'd23832, 16'd40672, 16'd26794, 16'd41351, 16'd64147, 16'd9370, 16'd17502, 16'd26613, 16'd46343, 16'd56666, 16'd48883, 16'd26321, 16'd29428, 16'd20441, 16'd39861, 16'd39447, 16'd38134, 16'd9854, 16'd53206, 16'd32158, 16'd61726, 16'd5061, 16'd63469, 16'd46701, 16'd29689});
	test_expansion(128'h2b50c6eb122c2b2f3fc3a8904e9df624, {16'd1285, 16'd24487, 16'd46326, 16'd7673, 16'd587, 16'd39564, 16'd17547, 16'd55468, 16'd4523, 16'd10493, 16'd41643, 16'd11821, 16'd36398, 16'd26370, 16'd65476, 16'd64616, 16'd30428, 16'd37415, 16'd38238, 16'd6042, 16'd41351, 16'd61314, 16'd14550, 16'd39128, 16'd43346, 16'd1928});
	test_expansion(128'h2b34451153af7690d057888d328068b6, {16'd40473, 16'd14162, 16'd24628, 16'd26798, 16'd22676, 16'd38690, 16'd64958, 16'd13011, 16'd9061, 16'd11012, 16'd26725, 16'd21219, 16'd61115, 16'd49124, 16'd16945, 16'd29747, 16'd11355, 16'd5698, 16'd16314, 16'd24911, 16'd45318, 16'd54946, 16'd30253, 16'd16506, 16'd455, 16'd24897});
	test_expansion(128'hffabb44ce4cefa74246bf0cb932f809f, {16'd38588, 16'd37518, 16'd19202, 16'd3908, 16'd12918, 16'd53562, 16'd37257, 16'd3810, 16'd26261, 16'd61445, 16'd63355, 16'd21555, 16'd39490, 16'd45057, 16'd10880, 16'd11243, 16'd17982, 16'd7614, 16'd12762, 16'd62575, 16'd61379, 16'd36683, 16'd36574, 16'd45968, 16'd9002, 16'd33341});
	test_expansion(128'h05a4c8507c51c8bb39d9628ef351e05a, {16'd50724, 16'd51717, 16'd23495, 16'd35767, 16'd39505, 16'd44167, 16'd16972, 16'd1542, 16'd49696, 16'd34944, 16'd28112, 16'd57870, 16'd63712, 16'd35675, 16'd59092, 16'd1782, 16'd1806, 16'd27631, 16'd22176, 16'd4913, 16'd40472, 16'd47003, 16'd40498, 16'd14578, 16'd40100, 16'd34046});
	test_expansion(128'hd0aa914dbd547d39a3a155453f40987c, {16'd7786, 16'd45248, 16'd3888, 16'd30721, 16'd15685, 16'd50744, 16'd55804, 16'd41663, 16'd44221, 16'd45369, 16'd49997, 16'd25814, 16'd3344, 16'd47814, 16'd44735, 16'd48671, 16'd22133, 16'd32365, 16'd16840, 16'd35223, 16'd59910, 16'd28467, 16'd3269, 16'd3052, 16'd32621, 16'd46905});
	test_expansion(128'h22e8e565a81ea45f58ee3fec5ba047d8, {16'd31391, 16'd11884, 16'd39012, 16'd46313, 16'd63467, 16'd61208, 16'd48626, 16'd59470, 16'd43299, 16'd59641, 16'd53873, 16'd29781, 16'd34516, 16'd6369, 16'd44447, 16'd40102, 16'd41393, 16'd29767, 16'd39171, 16'd58460, 16'd1031, 16'd3163, 16'd16644, 16'd44358, 16'd34649, 16'd7000});
	test_expansion(128'h57fc752a488e8d80fb93251829183753, {16'd31906, 16'd4776, 16'd45683, 16'd21866, 16'd22014, 16'd65039, 16'd26191, 16'd7276, 16'd2875, 16'd45864, 16'd13424, 16'd57123, 16'd11491, 16'd30873, 16'd59728, 16'd48376, 16'd13375, 16'd10300, 16'd49981, 16'd35518, 16'd23108, 16'd42497, 16'd36595, 16'd64338, 16'd16572, 16'd46744});
	test_expansion(128'h8444dc31e212f762b9df44b73e0ce047, {16'd63501, 16'd61800, 16'd57893, 16'd17666, 16'd19301, 16'd7275, 16'd45233, 16'd29206, 16'd19872, 16'd6737, 16'd38959, 16'd57612, 16'd12575, 16'd6583, 16'd22545, 16'd3055, 16'd39392, 16'd324, 16'd49844, 16'd28309, 16'd13179, 16'd6282, 16'd36732, 16'd41607, 16'd54175, 16'd35303});
	test_expansion(128'hc54f6f7492371cddd0d416e93ce520db, {16'd56083, 16'd23793, 16'd56539, 16'd29857, 16'd65193, 16'd35696, 16'd53969, 16'd47777, 16'd20134, 16'd7033, 16'd27880, 16'd7675, 16'd23712, 16'd17436, 16'd6256, 16'd33896, 16'd24340, 16'd15016, 16'd64859, 16'd59919, 16'd62636, 16'd28555, 16'd24825, 16'd23951, 16'd45988, 16'd21719});
	test_expansion(128'hf2630523c068d869fda1e0024735947c, {16'd14877, 16'd13139, 16'd23619, 16'd54189, 16'd36531, 16'd45620, 16'd11398, 16'd57240, 16'd16691, 16'd42084, 16'd21821, 16'd31867, 16'd42367, 16'd4769, 16'd63368, 16'd26566, 16'd11585, 16'd46918, 16'd49255, 16'd61885, 16'd6171, 16'd15339, 16'd21938, 16'd16122, 16'd50219, 16'd11748});
	test_expansion(128'hba7310884fbf111d54ac9bdc78df6eab, {16'd61402, 16'd5823, 16'd41820, 16'd41229, 16'd37866, 16'd1682, 16'd36698, 16'd65196, 16'd12120, 16'd12546, 16'd31769, 16'd35247, 16'd10716, 16'd36743, 16'd10925, 16'd46187, 16'd60296, 16'd5127, 16'd60288, 16'd18967, 16'd59161, 16'd21351, 16'd3198, 16'd29716, 16'd37395, 16'd62307});
	test_expansion(128'h796126e884cab63d3ad1d3d45864fe28, {16'd23215, 16'd28214, 16'd32375, 16'd54852, 16'd52040, 16'd63025, 16'd6830, 16'd6540, 16'd45822, 16'd13192, 16'd49299, 16'd61280, 16'd64152, 16'd13644, 16'd3083, 16'd50088, 16'd22692, 16'd14811, 16'd13586, 16'd12330, 16'd28587, 16'd9305, 16'd36185, 16'd47082, 16'd36497, 16'd40908});
	test_expansion(128'hf1e48c3d5168a81ee8d0935969ef5cc2, {16'd25273, 16'd54346, 16'd18586, 16'd37526, 16'd36807, 16'd2817, 16'd35694, 16'd55932, 16'd4360, 16'd63684, 16'd22603, 16'd23748, 16'd4315, 16'd52823, 16'd13876, 16'd4901, 16'd63262, 16'd51740, 16'd7004, 16'd7063, 16'd27372, 16'd54387, 16'd36009, 16'd48464, 16'd30031, 16'd12233});
	test_expansion(128'h86f1c026158eb46d6fa0fb79a3dc733c, {16'd43509, 16'd27942, 16'd51639, 16'd23735, 16'd53526, 16'd7879, 16'd24593, 16'd3391, 16'd35583, 16'd44255, 16'd14444, 16'd292, 16'd5995, 16'd9919, 16'd56454, 16'd21012, 16'd19915, 16'd8474, 16'd33081, 16'd65157, 16'd1075, 16'd44251, 16'd14034, 16'd24934, 16'd1382, 16'd54027});
	test_expansion(128'h720aae6453e316b842132d357dd8a1d4, {16'd23883, 16'd45449, 16'd18289, 16'd37218, 16'd16425, 16'd37680, 16'd16545, 16'd47813, 16'd47603, 16'd62405, 16'd56764, 16'd37052, 16'd14950, 16'd8570, 16'd41703, 16'd48889, 16'd7927, 16'd63326, 16'd34084, 16'd19203, 16'd8552, 16'd57253, 16'd39456, 16'd11463, 16'd58935, 16'd18774});
	test_expansion(128'h11375acd93d7863965b0d930097829f9, {16'd23531, 16'd40169, 16'd20150, 16'd47521, 16'd4395, 16'd12870, 16'd9059, 16'd40924, 16'd25881, 16'd63291, 16'd42023, 16'd4377, 16'd29560, 16'd57822, 16'd55960, 16'd12640, 16'd31764, 16'd33640, 16'd59183, 16'd44577, 16'd11751, 16'd17776, 16'd18091, 16'd43836, 16'd10765, 16'd15267});
	test_expansion(128'h18e5f08a73a972ba9f533ea22993f831, {16'd28840, 16'd48995, 16'd57155, 16'd58846, 16'd4214, 16'd59567, 16'd10243, 16'd14557, 16'd50569, 16'd19816, 16'd36237, 16'd13734, 16'd29257, 16'd52375, 16'd60012, 16'd11904, 16'd5295, 16'd47651, 16'd16224, 16'd37090, 16'd3435, 16'd50859, 16'd44004, 16'd64741, 16'd32412, 16'd23462});
	test_expansion(128'h14282eaed0563c62ea731232945cf009, {16'd32967, 16'd32987, 16'd46207, 16'd31616, 16'd33919, 16'd19320, 16'd18814, 16'd53871, 16'd28411, 16'd3290, 16'd5756, 16'd43789, 16'd15553, 16'd38732, 16'd38305, 16'd26365, 16'd37992, 16'd62345, 16'd48774, 16'd6086, 16'd26913, 16'd6025, 16'd1274, 16'd2607, 16'd59282, 16'd4198});
	test_expansion(128'hbffa81b7e29ef08ad508d018cdc90cf6, {16'd38340, 16'd49147, 16'd5881, 16'd7685, 16'd51036, 16'd32531, 16'd45483, 16'd40480, 16'd56646, 16'd65111, 16'd43138, 16'd22802, 16'd32148, 16'd27294, 16'd1010, 16'd13093, 16'd37937, 16'd5907, 16'd56260, 16'd22597, 16'd34296, 16'd40445, 16'd2397, 16'd23006, 16'd55557, 16'd54112});
	test_expansion(128'hb4173c1b83baa6851229c59c43b49369, {16'd60261, 16'd3781, 16'd53651, 16'd58310, 16'd5550, 16'd14151, 16'd7091, 16'd17706, 16'd32380, 16'd7484, 16'd58823, 16'd34815, 16'd12461, 16'd28965, 16'd18708, 16'd54973, 16'd16428, 16'd32351, 16'd52554, 16'd38196, 16'd15017, 16'd36802, 16'd29511, 16'd42387, 16'd62536, 16'd63706});
	test_expansion(128'hea8c90daa1de24af50ad636b4a29106a, {16'd56787, 16'd43319, 16'd57702, 16'd39428, 16'd44877, 16'd9759, 16'd50857, 16'd29585, 16'd38244, 16'd22619, 16'd30018, 16'd59258, 16'd40150, 16'd20595, 16'd44650, 16'd55002, 16'd20109, 16'd31361, 16'd53919, 16'd59497, 16'd65471, 16'd48619, 16'd51284, 16'd7906, 16'd39784, 16'd24249});
	test_expansion(128'h631bb24d2d64be3b1b2115170c0a1aaa, {16'd58877, 16'd50333, 16'd59114, 16'd59549, 16'd24264, 16'd53769, 16'd200, 16'd24834, 16'd58811, 16'd57204, 16'd31547, 16'd41159, 16'd62793, 16'd30990, 16'd43521, 16'd3523, 16'd15139, 16'd43542, 16'd24094, 16'd31527, 16'd15090, 16'd20480, 16'd63681, 16'd20179, 16'd26772, 16'd2676});
	test_expansion(128'hc5ce49f609004a0976f6439ebce899eb, {16'd10209, 16'd12566, 16'd6205, 16'd49660, 16'd47711, 16'd16545, 16'd24819, 16'd56051, 16'd64612, 16'd36667, 16'd9928, 16'd16112, 16'd2144, 16'd10895, 16'd48182, 16'd45798, 16'd60371, 16'd6317, 16'd51570, 16'd30717, 16'd64712, 16'd57129, 16'd38551, 16'd337, 16'd10295, 16'd27382});
	test_expansion(128'hef916bb548a77a473bdafb101f3cbd07, {16'd6508, 16'd51712, 16'd12701, 16'd11857, 16'd6831, 16'd50650, 16'd47548, 16'd55427, 16'd46978, 16'd9927, 16'd14416, 16'd62546, 16'd21495, 16'd18146, 16'd7743, 16'd25997, 16'd57067, 16'd59920, 16'd30466, 16'd11576, 16'd17076, 16'd3069, 16'd28151, 16'd46356, 16'd49681, 16'd51582});
	test_expansion(128'h8fdc557d093797f55635a1776780ad1a, {16'd35620, 16'd61093, 16'd63272, 16'd3921, 16'd5983, 16'd54690, 16'd53185, 16'd19910, 16'd64877, 16'd40209, 16'd34267, 16'd15622, 16'd42002, 16'd56483, 16'd711, 16'd21863, 16'd1860, 16'd33081, 16'd59882, 16'd54120, 16'd34910, 16'd8606, 16'd57616, 16'd7390, 16'd6156, 16'd55934});
	test_expansion(128'h70cb62f24cf6eb354b522a1d356f6908, {16'd62603, 16'd50729, 16'd42638, 16'd57660, 16'd13874, 16'd4405, 16'd45624, 16'd36628, 16'd39217, 16'd10106, 16'd23962, 16'd40326, 16'd24116, 16'd44197, 16'd57382, 16'd31272, 16'd6347, 16'd4962, 16'd49142, 16'd29150, 16'd2093, 16'd28613, 16'd5350, 16'd7989, 16'd28113, 16'd38697});
	test_expansion(128'hb8d8e92b6b1640b5b894d577fdd6bb8d, {16'd58218, 16'd48139, 16'd57967, 16'd34287, 16'd16821, 16'd2802, 16'd27404, 16'd11624, 16'd46299, 16'd24638, 16'd56341, 16'd56802, 16'd63811, 16'd51222, 16'd19028, 16'd58357, 16'd59227, 16'd16924, 16'd12227, 16'd4022, 16'd10501, 16'd43736, 16'd38299, 16'd45848, 16'd20847, 16'd15608});
	test_expansion(128'hf8244d25c3e6f7b3f1083d3905d8a834, {16'd17139, 16'd14911, 16'd19751, 16'd20318, 16'd51873, 16'd62668, 16'd59495, 16'd28536, 16'd35077, 16'd42738, 16'd39146, 16'd50583, 16'd11007, 16'd62332, 16'd6418, 16'd13978, 16'd64965, 16'd48024, 16'd56162, 16'd9173, 16'd6827, 16'd35328, 16'd53457, 16'd3144, 16'd54476, 16'd29474});
	test_expansion(128'h2dcbafd0ec4545b5f7deede8b2d09cd0, {16'd53696, 16'd58369, 16'd17805, 16'd43234, 16'd37177, 16'd54794, 16'd24485, 16'd19164, 16'd6921, 16'd59181, 16'd62572, 16'd25120, 16'd2911, 16'd60109, 16'd17455, 16'd18528, 16'd26994, 16'd46166, 16'd51139, 16'd56786, 16'd1283, 16'd50487, 16'd6744, 16'd57795, 16'd57289, 16'd35351});
	test_expansion(128'ha42bc3013e9149b97c4ffc2d45238a3b, {16'd35289, 16'd45087, 16'd16904, 16'd38591, 16'd25949, 16'd2395, 16'd55814, 16'd16596, 16'd60861, 16'd20531, 16'd10426, 16'd41564, 16'd48487, 16'd13434, 16'd52381, 16'd65147, 16'd17027, 16'd17001, 16'd8016, 16'd2817, 16'd7831, 16'd325, 16'd47744, 16'd2335, 16'd45108, 16'd22187});
	test_expansion(128'h8550aadc4073b5075a7abdb6e4ea3480, {16'd49332, 16'd36803, 16'd25179, 16'd12538, 16'd33296, 16'd45621, 16'd42563, 16'd50841, 16'd19145, 16'd3155, 16'd44439, 16'd11988, 16'd3122, 16'd50507, 16'd31742, 16'd63679, 16'd44684, 16'd19351, 16'd54874, 16'd4841, 16'd20969, 16'd45102, 16'd1904, 16'd14919, 16'd5379, 16'd3103});
	test_expansion(128'hc06a01b55072fe46aad913354c8223a0, {16'd54220, 16'd22095, 16'd11147, 16'd55266, 16'd18561, 16'd65253, 16'd39018, 16'd63806, 16'd22319, 16'd22694, 16'd63362, 16'd22287, 16'd37656, 16'd15195, 16'd6528, 16'd36770, 16'd6333, 16'd50201, 16'd64076, 16'd27571, 16'd57817, 16'd61923, 16'd58792, 16'd4740, 16'd17107, 16'd17109});
	test_expansion(128'he8a071221e27894642efdf53ff10eca4, {16'd48436, 16'd65456, 16'd45145, 16'd64348, 16'd38005, 16'd3954, 16'd33239, 16'd36515, 16'd24850, 16'd37191, 16'd30499, 16'd43753, 16'd25240, 16'd542, 16'd53502, 16'd53007, 16'd52420, 16'd4505, 16'd48242, 16'd54127, 16'd8473, 16'd18342, 16'd11278, 16'd20927, 16'd3748, 16'd25705});
	test_expansion(128'hd022b909e4a156672a11e40a25716aab, {16'd39163, 16'd16096, 16'd24013, 16'd62598, 16'd26055, 16'd13319, 16'd5736, 16'd19406, 16'd23238, 16'd31872, 16'd27141, 16'd32006, 16'd19578, 16'd9284, 16'd34674, 16'd11000, 16'd56163, 16'd29410, 16'd25656, 16'd40353, 16'd48606, 16'd59452, 16'd47691, 16'd51288, 16'd44568, 16'd40168});
	test_expansion(128'h474f7c1d850c7e270e264c4cb42fa86d, {16'd1055, 16'd59073, 16'd21883, 16'd60174, 16'd39455, 16'd28306, 16'd39726, 16'd17475, 16'd63378, 16'd57941, 16'd29251, 16'd4827, 16'd46047, 16'd41368, 16'd61637, 16'd1520, 16'd43350, 16'd5148, 16'd40743, 16'd605, 16'd52754, 16'd15535, 16'd606, 16'd51920, 16'd14738, 16'd21238});
	test_expansion(128'hc1206b890bed85f6b8bd83bb198a7f9d, {16'd11250, 16'd20379, 16'd17299, 16'd32801, 16'd36672, 16'd58304, 16'd55722, 16'd50040, 16'd28538, 16'd10575, 16'd18010, 16'd48461, 16'd14415, 16'd32492, 16'd60507, 16'd34472, 16'd7637, 16'd49915, 16'd56111, 16'd52519, 16'd57976, 16'd20507, 16'd8185, 16'd28785, 16'd58733, 16'd15829});
	test_expansion(128'hbafe87e2d6dba9ae006ac278e63ef755, {16'd6301, 16'd22171, 16'd28287, 16'd38729, 16'd10583, 16'd26675, 16'd45358, 16'd32422, 16'd52616, 16'd36569, 16'd26247, 16'd44635, 16'd32259, 16'd53812, 16'd54510, 16'd13499, 16'd13132, 16'd40916, 16'd16150, 16'd64179, 16'd20747, 16'd51895, 16'd9306, 16'd40443, 16'd9060, 16'd9867});
	test_expansion(128'h3a54cd8454e13ee36b94541c22d751c6, {16'd52588, 16'd26075, 16'd18461, 16'd13433, 16'd8332, 16'd3871, 16'd7875, 16'd33386, 16'd25782, 16'd27259, 16'd17999, 16'd50980, 16'd52292, 16'd56174, 16'd53693, 16'd6206, 16'd46894, 16'd46816, 16'd13344, 16'd29349, 16'd18212, 16'd23004, 16'd59026, 16'd57589, 16'd38026, 16'd61011});
	test_expansion(128'h358bbb4750ae59130bf09b78c12e7664, {16'd60340, 16'd22801, 16'd8600, 16'd35311, 16'd43599, 16'd16711, 16'd10679, 16'd23167, 16'd51357, 16'd42932, 16'd54521, 16'd12357, 16'd1432, 16'd24512, 16'd4370, 16'd25448, 16'd45988, 16'd26527, 16'd13247, 16'd54776, 16'd26539, 16'd42363, 16'd27740, 16'd4242, 16'd17134, 16'd14234});
	test_expansion(128'h3f7d917405571bb09956e9f01e25a42a, {16'd25953, 16'd14921, 16'd63597, 16'd34485, 16'd37493, 16'd22262, 16'd13170, 16'd16388, 16'd41758, 16'd21355, 16'd15504, 16'd49580, 16'd28588, 16'd9508, 16'd58227, 16'd44356, 16'd62378, 16'd983, 16'd17071, 16'd45079, 16'd42509, 16'd42409, 16'd28169, 16'd9537, 16'd42677, 16'd43337});
	test_expansion(128'h42d67b83f8948c1de947efe547d1244b, {16'd34688, 16'd62305, 16'd13787, 16'd5093, 16'd50948, 16'd19, 16'd58843, 16'd23072, 16'd62736, 16'd5973, 16'd1393, 16'd10585, 16'd64996, 16'd6615, 16'd49121, 16'd19379, 16'd34133, 16'd18242, 16'd16923, 16'd18416, 16'd16675, 16'd3168, 16'd24218, 16'd3860, 16'd27949, 16'd17164});
	test_expansion(128'h971eac067ed5755036d17b423db80ed6, {16'd43550, 16'd46535, 16'd18808, 16'd15747, 16'd2346, 16'd32, 16'd21516, 16'd63490, 16'd29394, 16'd54266, 16'd13879, 16'd176, 16'd52530, 16'd9301, 16'd58558, 16'd2222, 16'd29560, 16'd57262, 16'd24846, 16'd13850, 16'd31390, 16'd62716, 16'd54167, 16'd7351, 16'd30758, 16'd51458});
	test_expansion(128'h51b55fccdb7a5341e0f98cbcad0ac8e7, {16'd32578, 16'd20538, 16'd1490, 16'd2451, 16'd43492, 16'd29937, 16'd31403, 16'd53990, 16'd12359, 16'd8564, 16'd24310, 16'd20514, 16'd41933, 16'd4627, 16'd58055, 16'd429, 16'd3912, 16'd32723, 16'd10966, 16'd5275, 16'd57353, 16'd36588, 16'd59059, 16'd27384, 16'd55972, 16'd45482});
	test_expansion(128'h74d11ece883dd05e35fc3ff0f4e46f5c, {16'd2624, 16'd64017, 16'd53345, 16'd13560, 16'd7777, 16'd46214, 16'd30770, 16'd27050, 16'd25311, 16'd6647, 16'd49807, 16'd56950, 16'd61088, 16'd4761, 16'd55180, 16'd6501, 16'd26495, 16'd19796, 16'd28675, 16'd55330, 16'd2966, 16'd64628, 16'd13929, 16'd1537, 16'd64889, 16'd20065});
	test_expansion(128'ha9a0a6a3b529a392499baad272208774, {16'd20767, 16'd29808, 16'd36607, 16'd13112, 16'd59134, 16'd29357, 16'd10503, 16'd50370, 16'd44637, 16'd63371, 16'd20346, 16'd17017, 16'd54456, 16'd56791, 16'd33625, 16'd38067, 16'd48959, 16'd24212, 16'd31856, 16'd29078, 16'd55780, 16'd40050, 16'd197, 16'd51868, 16'd11653, 16'd61393});
	test_expansion(128'h6ce1378b809f8d0d021fd7b650d1ec7a, {16'd55891, 16'd20835, 16'd54830, 16'd55797, 16'd9022, 16'd44566, 16'd30932, 16'd53495, 16'd18648, 16'd59091, 16'd16611, 16'd53552, 16'd24008, 16'd7521, 16'd33659, 16'd38315, 16'd59496, 16'd60546, 16'd39985, 16'd7980, 16'd16285, 16'd26712, 16'd155, 16'd15748, 16'd12488, 16'd1110});
	test_expansion(128'h6266455ecf3abdbad88cf561aa586344, {16'd37906, 16'd13550, 16'd28916, 16'd1008, 16'd41760, 16'd30967, 16'd61287, 16'd4709, 16'd27831, 16'd50722, 16'd53161, 16'd10005, 16'd33991, 16'd403, 16'd22018, 16'd12608, 16'd61276, 16'd56056, 16'd26968, 16'd9041, 16'd61369, 16'd10208, 16'd60448, 16'd5092, 16'd56542, 16'd53842});
	test_expansion(128'h1c221f54de2f191c68a486450c134cba, {16'd57426, 16'd61197, 16'd25691, 16'd32478, 16'd59533, 16'd28495, 16'd28075, 16'd50136, 16'd60224, 16'd35400, 16'd17793, 16'd28728, 16'd25309, 16'd36175, 16'd22017, 16'd33007, 16'd42886, 16'd37647, 16'd23897, 16'd18704, 16'd5175, 16'd42646, 16'd47774, 16'd57287, 16'd50617, 16'd17780});
	test_expansion(128'hc460f64b405f732ce6656baa9282c3c0, {16'd46042, 16'd28268, 16'd11786, 16'd40412, 16'd53390, 16'd62081, 16'd51208, 16'd14487, 16'd50959, 16'd22060, 16'd62202, 16'd17977, 16'd37275, 16'd55749, 16'd38410, 16'd63712, 16'd20994, 16'd37860, 16'd22371, 16'd13651, 16'd39712, 16'd12795, 16'd41696, 16'd22146, 16'd29450, 16'd37213});
	test_expansion(128'hfc439dbe113d336177f1f04114924543, {16'd21654, 16'd34742, 16'd40386, 16'd48859, 16'd9352, 16'd49073, 16'd7635, 16'd55011, 16'd43879, 16'd1820, 16'd24569, 16'd1635, 16'd18811, 16'd58436, 16'd34895, 16'd14847, 16'd27052, 16'd58835, 16'd15273, 16'd9380, 16'd58344, 16'd63862, 16'd47792, 16'd13904, 16'd53950, 16'd5328});
	test_expansion(128'hc0df168f10a878e0bb56ec1774157936, {16'd54417, 16'd29974, 16'd54226, 16'd54045, 16'd12566, 16'd53589, 16'd63216, 16'd10430, 16'd59973, 16'd63951, 16'd10762, 16'd62535, 16'd50342, 16'd10565, 16'd22134, 16'd46313, 16'd10234, 16'd59432, 16'd35623, 16'd35578, 16'd55093, 16'd46571, 16'd18980, 16'd50114, 16'd55041, 16'd57330});
	test_expansion(128'h3a6739f951d7859a1bea0db468b3f4c4, {16'd52762, 16'd43583, 16'd26913, 16'd60832, 16'd45361, 16'd52186, 16'd57773, 16'd53902, 16'd21570, 16'd29827, 16'd19312, 16'd16077, 16'd5898, 16'd32437, 16'd30340, 16'd62452, 16'd39621, 16'd30364, 16'd12212, 16'd36195, 16'd38946, 16'd49764, 16'd13948, 16'd21253, 16'd19924, 16'd6146});
	test_expansion(128'h4efb1653bd7a1ec3eddb7151696fb3fa, {16'd21734, 16'd55490, 16'd38807, 16'd43728, 16'd50139, 16'd56423, 16'd20919, 16'd45391, 16'd1736, 16'd64032, 16'd26837, 16'd17513, 16'd23320, 16'd34437, 16'd32122, 16'd5285, 16'd35489, 16'd57941, 16'd59680, 16'd48227, 16'd35158, 16'd54757, 16'd46710, 16'd24389, 16'd33553, 16'd48738});
	test_expansion(128'h1909d3b9bbba876a6b7884efa70e031a, {16'd28698, 16'd36535, 16'd23779, 16'd12701, 16'd18362, 16'd52502, 16'd45771, 16'd58638, 16'd51533, 16'd31047, 16'd39381, 16'd29654, 16'd20505, 16'd13712, 16'd6389, 16'd56939, 16'd56444, 16'd19681, 16'd65334, 16'd662, 16'd12030, 16'd16085, 16'd39785, 16'd34469, 16'd54679, 16'd50163});
	test_expansion(128'h0d634ed4b8995576b3cc6e1a92e21670, {16'd57537, 16'd30165, 16'd15921, 16'd53607, 16'd24832, 16'd49383, 16'd30702, 16'd33956, 16'd25854, 16'd43137, 16'd50215, 16'd43207, 16'd35688, 16'd25919, 16'd75, 16'd52428, 16'd34657, 16'd17474, 16'd38052, 16'd26953, 16'd34579, 16'd33105, 16'd7930, 16'd13724, 16'd8240, 16'd46382});
	test_expansion(128'h9525bff5c01dd6d58671fbe50f37a9f6, {16'd9362, 16'd61222, 16'd41885, 16'd9782, 16'd10036, 16'd61250, 16'd43665, 16'd20088, 16'd54857, 16'd34698, 16'd53060, 16'd13030, 16'd24007, 16'd64126, 16'd37180, 16'd60300, 16'd52852, 16'd27077, 16'd19752, 16'd17649, 16'd13489, 16'd4296, 16'd4855, 16'd34290, 16'd63349, 16'd11402});
	test_expansion(128'h2da5db2ee0f2d671c8018b9acd5198d6, {16'd6029, 16'd41819, 16'd52160, 16'd58666, 16'd37838, 16'd55629, 16'd10369, 16'd58894, 16'd12983, 16'd45910, 16'd39011, 16'd29321, 16'd41112, 16'd13129, 16'd54219, 16'd31640, 16'd7512, 16'd50268, 16'd20, 16'd13398, 16'd12145, 16'd50783, 16'd25373, 16'd60049, 16'd31335, 16'd51594});
	test_expansion(128'h33388b1ffa83a3ecbd306a71c784ff03, {16'd45566, 16'd14491, 16'd6594, 16'd34170, 16'd39616, 16'd37798, 16'd45753, 16'd51903, 16'd34551, 16'd54277, 16'd20504, 16'd34423, 16'd27910, 16'd4741, 16'd53958, 16'd38654, 16'd31817, 16'd60271, 16'd5171, 16'd47687, 16'd5470, 16'd8412, 16'd48264, 16'd63946, 16'd44645, 16'd31399});
	test_expansion(128'hcb8c6f2389b6b341498d8e29937d2a9b, {16'd5804, 16'd10339, 16'd20019, 16'd24539, 16'd21197, 16'd34297, 16'd4393, 16'd54324, 16'd44618, 16'd4064, 16'd47327, 16'd11803, 16'd47722, 16'd51670, 16'd34238, 16'd13191, 16'd9665, 16'd48525, 16'd21180, 16'd51163, 16'd36965, 16'd52971, 16'd49556, 16'd31686, 16'd12909, 16'd2471});
	test_expansion(128'hb4e70c03474be72c198ea97af408121b, {16'd19859, 16'd62479, 16'd7865, 16'd55831, 16'd8233, 16'd48278, 16'd7512, 16'd42924, 16'd39328, 16'd6862, 16'd45403, 16'd53116, 16'd38620, 16'd35534, 16'd1944, 16'd55813, 16'd63919, 16'd16548, 16'd18628, 16'd17749, 16'd29110, 16'd13440, 16'd44760, 16'd39323, 16'd62882, 16'd64313});
	test_expansion(128'h79d1cb028e830e0287fcf261ac10a687, {16'd25064, 16'd7040, 16'd32007, 16'd14, 16'd3244, 16'd19947, 16'd1686, 16'd64610, 16'd63389, 16'd17081, 16'd46251, 16'd31889, 16'd10384, 16'd1163, 16'd15035, 16'd20659, 16'd56780, 16'd40272, 16'd255, 16'd746, 16'd54966, 16'd44370, 16'd51947, 16'd56635, 16'd50816, 16'd59162});
	test_expansion(128'ha423f537aa5cb4f8ced3c08f1c1b77ef, {16'd51346, 16'd11242, 16'd64120, 16'd28482, 16'd53857, 16'd43440, 16'd13514, 16'd21732, 16'd57688, 16'd29233, 16'd24572, 16'd35314, 16'd34945, 16'd64396, 16'd6965, 16'd15898, 16'd29965, 16'd49947, 16'd49073, 16'd49511, 16'd63182, 16'd65533, 16'd48265, 16'd38846, 16'd53131, 16'd54084});
	test_expansion(128'hefe1735f2c5fe7ed76d3261107ea65ec, {16'd20313, 16'd51953, 16'd6115, 16'd4272, 16'd17384, 16'd60851, 16'd13809, 16'd40227, 16'd61474, 16'd28023, 16'd34527, 16'd50168, 16'd47241, 16'd25594, 16'd4483, 16'd59389, 16'd51387, 16'd1658, 16'd6682, 16'd8520, 16'd53758, 16'd15833, 16'd24351, 16'd6172, 16'd7605, 16'd32413});
	test_expansion(128'he23d253425aee19e080c0ec0388e65a4, {16'd22708, 16'd13574, 16'd7846, 16'd22611, 16'd6549, 16'd26778, 16'd17385, 16'd27893, 16'd65006, 16'd42394, 16'd38621, 16'd13256, 16'd55693, 16'd45022, 16'd14688, 16'd13228, 16'd48985, 16'd49734, 16'd42433, 16'd57036, 16'd16605, 16'd57535, 16'd35829, 16'd3008, 16'd16132, 16'd28237});
	test_expansion(128'hbbc85b0038c291acddf65bacd0f27fde, {16'd39152, 16'd15369, 16'd43629, 16'd31604, 16'd24578, 16'd21247, 16'd45371, 16'd36738, 16'd62514, 16'd47937, 16'd9040, 16'd59591, 16'd32844, 16'd20933, 16'd36000, 16'd9536, 16'd18596, 16'd43497, 16'd60329, 16'd5516, 16'd47020, 16'd57695, 16'd63568, 16'd53383, 16'd9065, 16'd9860});
	test_expansion(128'hd390540a8ebbf1332251324be59db4ae, {16'd11789, 16'd39851, 16'd27881, 16'd41951, 16'd28587, 16'd15697, 16'd34183, 16'd31924, 16'd13780, 16'd22415, 16'd28879, 16'd48944, 16'd13190, 16'd27691, 16'd20471, 16'd2748, 16'd19300, 16'd1783, 16'd12534, 16'd12193, 16'd17441, 16'd59180, 16'd56534, 16'd26461, 16'd54574, 16'd28982});
	test_expansion(128'hdce4413262f9fb9d7cefa0dc976e5ad8, {16'd491, 16'd21774, 16'd54902, 16'd9746, 16'd8283, 16'd63190, 16'd20092, 16'd7704, 16'd10022, 16'd25546, 16'd39952, 16'd61245, 16'd6124, 16'd32657, 16'd36403, 16'd38526, 16'd25730, 16'd30781, 16'd49451, 16'd52765, 16'd14132, 16'd47953, 16'd43603, 16'd5351, 16'd64698, 16'd59194});
	test_expansion(128'hc8f420735caafd2701c5cb63628dac63, {16'd65424, 16'd8744, 16'd42398, 16'd43919, 16'd8515, 16'd11980, 16'd59635, 16'd25916, 16'd23460, 16'd36620, 16'd42588, 16'd52960, 16'd7373, 16'd22378, 16'd2009, 16'd43473, 16'd17382, 16'd12529, 16'd1934, 16'd21202, 16'd7049, 16'd58840, 16'd45617, 16'd46138, 16'd43028, 16'd20567});
	test_expansion(128'h37a465072c495911221050cf20e75c69, {16'd20501, 16'd12924, 16'd889, 16'd7713, 16'd31397, 16'd54169, 16'd8343, 16'd55907, 16'd61460, 16'd47457, 16'd3034, 16'd20921, 16'd14999, 16'd43777, 16'd64915, 16'd50001, 16'd48812, 16'd46612, 16'd41039, 16'd6410, 16'd25420, 16'd46575, 16'd26714, 16'd17509, 16'd30653, 16'd54090});
	test_expansion(128'hea7b72038f50cb95ed69ff237abd6c7c, {16'd60211, 16'd58255, 16'd52484, 16'd6042, 16'd19067, 16'd60370, 16'd64746, 16'd58066, 16'd1718, 16'd45088, 16'd37153, 16'd26631, 16'd61567, 16'd33954, 16'd33648, 16'd11163, 16'd48821, 16'd39814, 16'd3783, 16'd12603, 16'd51018, 16'd54022, 16'd16011, 16'd62979, 16'd36620, 16'd2647});
	test_expansion(128'h3afc126bd5b2155ca62fce66f51ef6aa, {16'd29906, 16'd49747, 16'd56849, 16'd9534, 16'd48918, 16'd25417, 16'd38331, 16'd23280, 16'd37219, 16'd37406, 16'd34990, 16'd26781, 16'd39564, 16'd25428, 16'd27367, 16'd36830, 16'd6866, 16'd16285, 16'd38369, 16'd61359, 16'd5343, 16'd6328, 16'd26595, 16'd45851, 16'd15857, 16'd18051});
	test_expansion(128'h53e872ee742e06661c3a77672ed94aa2, {16'd45439, 16'd40981, 16'd58762, 16'd47374, 16'd158, 16'd61802, 16'd50882, 16'd54943, 16'd31788, 16'd61398, 16'd27990, 16'd6251, 16'd65073, 16'd59876, 16'd12557, 16'd17500, 16'd2332, 16'd52684, 16'd13891, 16'd53868, 16'd21315, 16'd1383, 16'd62607, 16'd26344, 16'd53660, 16'd6253});
	test_expansion(128'ha5e587f35af1d7c39c8edc32301df576, {16'd15264, 16'd22229, 16'd8660, 16'd25749, 16'd55016, 16'd30038, 16'd11011, 16'd25406, 16'd56965, 16'd683, 16'd61210, 16'd50886, 16'd39090, 16'd11104, 16'd5973, 16'd7593, 16'd16429, 16'd63393, 16'd61886, 16'd17334, 16'd60645, 16'd840, 16'd26784, 16'd10344, 16'd9204, 16'd10995});
	test_expansion(128'he03bce6fbd5aa0786f90f5e990b96e12, {16'd29088, 16'd11371, 16'd2523, 16'd5262, 16'd44462, 16'd4606, 16'd36676, 16'd8727, 16'd49863, 16'd24801, 16'd64254, 16'd32572, 16'd41097, 16'd59594, 16'd26152, 16'd5470, 16'd35032, 16'd16939, 16'd26973, 16'd12677, 16'd5105, 16'd61231, 16'd6919, 16'd7531, 16'd44864, 16'd58600});
	test_expansion(128'h3e33d91c4bc01f4546212dbf5c05a27f, {16'd32612, 16'd60426, 16'd10858, 16'd47316, 16'd39933, 16'd19738, 16'd60515, 16'd44478, 16'd45550, 16'd19943, 16'd46344, 16'd176, 16'd14290, 16'd23337, 16'd32309, 16'd30417, 16'd26368, 16'd57194, 16'd5817, 16'd28156, 16'd19960, 16'd56077, 16'd45596, 16'd47284, 16'd36295, 16'd38349});
	test_expansion(128'h525b098a8457f3276b2d31f02e8db0e7, {16'd49657, 16'd36143, 16'd56977, 16'd16179, 16'd47324, 16'd12327, 16'd44907, 16'd46868, 16'd17518, 16'd43134, 16'd25694, 16'd10356, 16'd8940, 16'd56843, 16'd51624, 16'd65235, 16'd24792, 16'd29074, 16'd31364, 16'd55073, 16'd4239, 16'd6635, 16'd31298, 16'd62894, 16'd2231, 16'd54700});
	test_expansion(128'hf745cdb2d95702023efaf50117cdd800, {16'd21064, 16'd28100, 16'd51342, 16'd27375, 16'd27745, 16'd45383, 16'd17164, 16'd19743, 16'd62725, 16'd62096, 16'd15995, 16'd5913, 16'd35051, 16'd4532, 16'd5416, 16'd59845, 16'd46320, 16'd54295, 16'd8277, 16'd49734, 16'd40468, 16'd29128, 16'd14633, 16'd36444, 16'd26783, 16'd48794});
	test_expansion(128'h68fddc8d697838ab413f86b5da778ab6, {16'd12047, 16'd31397, 16'd15891, 16'd61810, 16'd49509, 16'd35557, 16'd11702, 16'd7732, 16'd28204, 16'd44092, 16'd597, 16'd44297, 16'd28995, 16'd928, 16'd50021, 16'd15294, 16'd3229, 16'd814, 16'd19714, 16'd51975, 16'd58020, 16'd54127, 16'd26772, 16'd11347, 16'd40664, 16'd16889});
	test_expansion(128'he22ebbfd69d7eb07631d5f21bb567414, {16'd41964, 16'd42684, 16'd57585, 16'd12398, 16'd62234, 16'd59491, 16'd8008, 16'd18544, 16'd36844, 16'd65205, 16'd2020, 16'd16817, 16'd63464, 16'd7967, 16'd14287, 16'd42776, 16'd39031, 16'd8663, 16'd29263, 16'd5829, 16'd33431, 16'd6123, 16'd7800, 16'd51555, 16'd36286, 16'd42736});
	test_expansion(128'hbbeb9fe50c534f1cdb5385a188329056, {16'd53271, 16'd23971, 16'd55830, 16'd65283, 16'd26379, 16'd7226, 16'd43303, 16'd31654, 16'd58575, 16'd27649, 16'd3029, 16'd1406, 16'd53557, 16'd41015, 16'd36604, 16'd24365, 16'd35106, 16'd33105, 16'd55803, 16'd31376, 16'd21656, 16'd39039, 16'd10149, 16'd27897, 16'd55189, 16'd38636});
	test_expansion(128'he4154a80e1daebe1886cc711c36c5550, {16'd1584, 16'd7738, 16'd46233, 16'd34889, 16'd13581, 16'd24561, 16'd13467, 16'd57345, 16'd34532, 16'd34508, 16'd7244, 16'd45839, 16'd2068, 16'd55660, 16'd22451, 16'd59955, 16'd10486, 16'd31740, 16'd59998, 16'd27148, 16'd42622, 16'd58653, 16'd58640, 16'd27952, 16'd6596, 16'd62194});
	test_expansion(128'h9cf2969082e09922c15bc1c71a418106, {16'd47722, 16'd32335, 16'd5021, 16'd8858, 16'd14632, 16'd58569, 16'd4103, 16'd17666, 16'd16566, 16'd40198, 16'd551, 16'd60655, 16'd8445, 16'd7415, 16'd1448, 16'd37321, 16'd38488, 16'd7942, 16'd54166, 16'd34359, 16'd2353, 16'd54136, 16'd65131, 16'd26234, 16'd45692, 16'd10832});
	test_expansion(128'h58196a66fda795a09d2ab95c5f6cf32f, {16'd65220, 16'd1114, 16'd358, 16'd28062, 16'd6335, 16'd41645, 16'd32388, 16'd61418, 16'd22702, 16'd41360, 16'd55888, 16'd45057, 16'd55349, 16'd22632, 16'd10786, 16'd15663, 16'd52297, 16'd55364, 16'd55090, 16'd35147, 16'd15689, 16'd42229, 16'd15547, 16'd15354, 16'd42829, 16'd21270});
	test_expansion(128'h961e175808be13c01f9f17c5f915c8c1, {16'd44854, 16'd62372, 16'd42918, 16'd28217, 16'd773, 16'd51261, 16'd3964, 16'd58840, 16'd56092, 16'd6782, 16'd29233, 16'd48321, 16'd12031, 16'd50335, 16'd25544, 16'd51964, 16'd25855, 16'd41319, 16'd46864, 16'd14498, 16'd19468, 16'd59687, 16'd23082, 16'd4992, 16'd33965, 16'd44072});
	test_expansion(128'h484376a4b9df116fec347816bb3fdf84, {16'd4733, 16'd28097, 16'd21113, 16'd13600, 16'd6753, 16'd54089, 16'd40096, 16'd30936, 16'd3026, 16'd57993, 16'd31151, 16'd1648, 16'd38867, 16'd17334, 16'd33031, 16'd12723, 16'd65311, 16'd56463, 16'd1054, 16'd8568, 16'd58018, 16'd29448, 16'd566, 16'd33374, 16'd61976, 16'd51629});
	test_expansion(128'h2006470ff13fca34b6917985cb0e6096, {16'd30601, 16'd31063, 16'd25292, 16'd13672, 16'd25949, 16'd46296, 16'd24304, 16'd8604, 16'd39438, 16'd20695, 16'd50433, 16'd37534, 16'd58841, 16'd51028, 16'd52345, 16'd27883, 16'd45214, 16'd55643, 16'd15115, 16'd23842, 16'd24840, 16'd57731, 16'd18516, 16'd2782, 16'd57585, 16'd43883});
	test_expansion(128'hbaa7177b272fc47682a1197b60176fd0, {16'd55453, 16'd45803, 16'd48045, 16'd40824, 16'd33737, 16'd53937, 16'd50997, 16'd42824, 16'd1548, 16'd57176, 16'd18527, 16'd52640, 16'd61383, 16'd56869, 16'd61727, 16'd33475, 16'd45053, 16'd64427, 16'd25740, 16'd61601, 16'd15374, 16'd13458, 16'd40280, 16'd41779, 16'd56051, 16'd26232});
	test_expansion(128'h5d13230eb628b6527b42ddf2163f9cc5, {16'd39324, 16'd40874, 16'd20615, 16'd25260, 16'd19122, 16'd13789, 16'd60563, 16'd30507, 16'd4286, 16'd18142, 16'd45432, 16'd45246, 16'd40938, 16'd3709, 16'd32212, 16'd22632, 16'd17559, 16'd50180, 16'd15164, 16'd1569, 16'd34917, 16'd64334, 16'd5151, 16'd54603, 16'd37841, 16'd12115});
	test_expansion(128'h638f4e70feb37c52b23cef5800a4f91f, {16'd32516, 16'd3379, 16'd7813, 16'd20614, 16'd10282, 16'd64820, 16'd16074, 16'd55680, 16'd51930, 16'd39004, 16'd37219, 16'd32799, 16'd43605, 16'd62656, 16'd47566, 16'd40395, 16'd28391, 16'd8767, 16'd45214, 16'd53674, 16'd21894, 16'd52421, 16'd38774, 16'd15628, 16'd4154, 16'd29448});
	test_expansion(128'h77e0e24916688a8e80c319f6ff654ff2, {16'd28741, 16'd25399, 16'd24955, 16'd13283, 16'd5026, 16'd31031, 16'd63137, 16'd44983, 16'd28967, 16'd13731, 16'd18358, 16'd14629, 16'd23935, 16'd38070, 16'd64999, 16'd61511, 16'd47954, 16'd45373, 16'd60173, 16'd29635, 16'd52073, 16'd38239, 16'd62918, 16'd58209, 16'd33444, 16'd19995});
	test_expansion(128'h065c7e42859a9e738d456505e1219541, {16'd64056, 16'd47141, 16'd9031, 16'd45771, 16'd7307, 16'd45683, 16'd14767, 16'd62650, 16'd22554, 16'd35239, 16'd35582, 16'd59852, 16'd62375, 16'd26933, 16'd29887, 16'd57842, 16'd31812, 16'd22981, 16'd62896, 16'd52812, 16'd61656, 16'd55220, 16'd14697, 16'd17933, 16'd54625, 16'd55258});
	test_expansion(128'h9de88b5e73456226b7d9b1bc2ad75c52, {16'd17632, 16'd46745, 16'd29401, 16'd31355, 16'd64271, 16'd60798, 16'd9123, 16'd7021, 16'd39755, 16'd50421, 16'd8050, 16'd11376, 16'd46292, 16'd787, 16'd5112, 16'd30289, 16'd5050, 16'd42019, 16'd27304, 16'd31362, 16'd25757, 16'd51671, 16'd29471, 16'd31414, 16'd47842, 16'd37138});
	test_expansion(128'he3148460816bf910b8706c8bd74266e6, {16'd53660, 16'd59001, 16'd59411, 16'd40242, 16'd15532, 16'd59615, 16'd19941, 16'd57935, 16'd39717, 16'd53021, 16'd58908, 16'd13543, 16'd41580, 16'd13391, 16'd1519, 16'd50060, 16'd55095, 16'd52570, 16'd51394, 16'd58542, 16'd27299, 16'd62261, 16'd42449, 16'd23978, 16'd16394, 16'd27664});
	test_expansion(128'he633561952b3e3807e01ea534c9ccaf5, {16'd61430, 16'd28986, 16'd18231, 16'd15707, 16'd24131, 16'd37058, 16'd28409, 16'd21112, 16'd41564, 16'd12771, 16'd10143, 16'd7528, 16'd59558, 16'd31952, 16'd52970, 16'd17703, 16'd36653, 16'd31089, 16'd23732, 16'd34728, 16'd46060, 16'd42719, 16'd63537, 16'd21701, 16'd59050, 16'd60160});
	test_expansion(128'h0d29ff49ff94e159b37ed0061a333e22, {16'd21904, 16'd32080, 16'd17021, 16'd62375, 16'd33206, 16'd20097, 16'd1600, 16'd27200, 16'd34541, 16'd56265, 16'd15497, 16'd35925, 16'd8429, 16'd32192, 16'd28646, 16'd56217, 16'd25881, 16'd42238, 16'd10564, 16'd50203, 16'd29003, 16'd13569, 16'd3944, 16'd8857, 16'd149, 16'd56220});
	test_expansion(128'hf06c98733c04193b7d145124a90c5cb0, {16'd50885, 16'd9940, 16'd42090, 16'd26632, 16'd24866, 16'd63433, 16'd39583, 16'd34447, 16'd58234, 16'd5763, 16'd56843, 16'd56240, 16'd1760, 16'd5735, 16'd25584, 16'd42644, 16'd22213, 16'd25012, 16'd21764, 16'd32355, 16'd7153, 16'd16756, 16'd6386, 16'd4004, 16'd47328, 16'd47809});
	test_expansion(128'h06357d2912fb0f8610d5213131b8e3ea, {16'd49853, 16'd15036, 16'd45109, 16'd4710, 16'd30016, 16'd50246, 16'd7379, 16'd49958, 16'd20549, 16'd29138, 16'd22999, 16'd34860, 16'd61547, 16'd50317, 16'd20030, 16'd34135, 16'd41962, 16'd22126, 16'd38135, 16'd30577, 16'd21505, 16'd25046, 16'd17789, 16'd45042, 16'd32545, 16'd59319});
	test_expansion(128'h23347e8d59855edc595c7498b7754cb7, {16'd33402, 16'd3399, 16'd38839, 16'd59678, 16'd1681, 16'd59183, 16'd8448, 16'd61761, 16'd36120, 16'd38363, 16'd54657, 16'd37, 16'd63684, 16'd41, 16'd13662, 16'd51713, 16'd51345, 16'd59409, 16'd24862, 16'd13965, 16'd64080, 16'd36510, 16'd11349, 16'd36830, 16'd49231, 16'd17511});
	test_expansion(128'hf4fff660fb6eb1f2f1b6446365fd3e2c, {16'd62384, 16'd20510, 16'd63954, 16'd46807, 16'd59362, 16'd26922, 16'd20231, 16'd27020, 16'd48977, 16'd5522, 16'd16400, 16'd31596, 16'd6496, 16'd6015, 16'd12040, 16'd56101, 16'd28712, 16'd4432, 16'd36895, 16'd49963, 16'd20364, 16'd2909, 16'd57005, 16'd60955, 16'd64819, 16'd40881});
	test_expansion(128'h7d90c6cbd73007e4bacd31cafbd22c70, {16'd13664, 16'd1197, 16'd30922, 16'd42325, 16'd11610, 16'd10841, 16'd16170, 16'd5494, 16'd6308, 16'd62557, 16'd57912, 16'd56644, 16'd30737, 16'd46740, 16'd40435, 16'd28698, 16'd60008, 16'd40286, 16'd49559, 16'd16687, 16'd36412, 16'd48070, 16'd35697, 16'd64539, 16'd29247, 16'd9188});
	test_expansion(128'hac1db536db314214358edf947f0a9293, {16'd30836, 16'd44104, 16'd26963, 16'd11769, 16'd54006, 16'd27952, 16'd27820, 16'd53565, 16'd28819, 16'd55153, 16'd31650, 16'd32290, 16'd30768, 16'd56110, 16'd31022, 16'd9218, 16'd45548, 16'd2447, 16'd61176, 16'd17331, 16'd2362, 16'd65514, 16'd13407, 16'd41569, 16'd53975, 16'd20564});
	test_expansion(128'he4a593b141c8484f59f9c09995f452cb, {16'd20257, 16'd11288, 16'd52807, 16'd11224, 16'd32257, 16'd43640, 16'd64402, 16'd20881, 16'd29423, 16'd30862, 16'd60069, 16'd48339, 16'd18541, 16'd11259, 16'd46961, 16'd57909, 16'd8161, 16'd32237, 16'd32841, 16'd14915, 16'd43293, 16'd48455, 16'd27335, 16'd40756, 16'd9481, 16'd59510});
	test_expansion(128'ha01b14fe041910c41638973d94b1a8a8, {16'd5719, 16'd10084, 16'd33810, 16'd22729, 16'd56671, 16'd41935, 16'd31098, 16'd2995, 16'd35224, 16'd36140, 16'd64977, 16'd44948, 16'd5941, 16'd47315, 16'd61803, 16'd5718, 16'd60634, 16'd10191, 16'd16395, 16'd64560, 16'd27469, 16'd293, 16'd57612, 16'd54447, 16'd55770, 16'd37229});
	test_expansion(128'he0f7b3cb92f94b884ff7469aa1ef7d45, {16'd14603, 16'd32648, 16'd37845, 16'd61637, 16'd11600, 16'd52677, 16'd52527, 16'd42601, 16'd32492, 16'd17290, 16'd26934, 16'd14881, 16'd42611, 16'd49864, 16'd39862, 16'd23756, 16'd47598, 16'd36554, 16'd8921, 16'd49221, 16'd32546, 16'd50603, 16'd42293, 16'd9010, 16'd44289, 16'd38928});
	test_expansion(128'h81bfe5dc4bec482898bb51c24a0e9e8d, {16'd23401, 16'd27141, 16'd39153, 16'd20993, 16'd27127, 16'd52316, 16'd33822, 16'd24867, 16'd9930, 16'd33908, 16'd38030, 16'd1318, 16'd2275, 16'd55770, 16'd609, 16'd43162, 16'd999, 16'd62574, 16'd7971, 16'd27323, 16'd52151, 16'd38292, 16'd14658, 16'd41551, 16'd4351, 16'd49090});
	test_expansion(128'ha7448004d32d5855e30bc51b92cb3e78, {16'd19281, 16'd53218, 16'd54622, 16'd45067, 16'd43691, 16'd3487, 16'd8794, 16'd40646, 16'd34320, 16'd62959, 16'd45973, 16'd46149, 16'd12643, 16'd14374, 16'd14393, 16'd22227, 16'd10863, 16'd8858, 16'd23407, 16'd13280, 16'd47195, 16'd51155, 16'd41556, 16'd11947, 16'd14027, 16'd61951});
	test_expansion(128'h2248ee0ac3b747db3f8b303a8f5bc569, {16'd3632, 16'd36517, 16'd53015, 16'd35938, 16'd15366, 16'd16792, 16'd78, 16'd53554, 16'd63884, 16'd26036, 16'd38775, 16'd39854, 16'd1157, 16'd40475, 16'd31854, 16'd20044, 16'd5256, 16'd30029, 16'd36010, 16'd43510, 16'd28240, 16'd41200, 16'd429, 16'd46894, 16'd57825, 16'd31387});
	test_expansion(128'h8aefa5631b13f5a0196c64c9a6be8428, {16'd55914, 16'd61822, 16'd53309, 16'd10422, 16'd42827, 16'd11135, 16'd22355, 16'd3830, 16'd39508, 16'd57464, 16'd13363, 16'd34440, 16'd50208, 16'd55540, 16'd31775, 16'd52663, 16'd44530, 16'd53059, 16'd14701, 16'd50665, 16'd42631, 16'd5196, 16'd16720, 16'd9995, 16'd32759, 16'd28761});
	test_expansion(128'h68d6bb920bf28c386de7a74b8bf96129, {16'd1944, 16'd8029, 16'd27480, 16'd58355, 16'd19431, 16'd35315, 16'd30878, 16'd62285, 16'd13774, 16'd7209, 16'd40768, 16'd20746, 16'd4955, 16'd13967, 16'd38426, 16'd50159, 16'd11089, 16'd22614, 16'd59240, 16'd53004, 16'd14941, 16'd28185, 16'd34479, 16'd17776, 16'd27475, 16'd54265});
	test_expansion(128'he37fa414df68fb236979a3c3f095678d, {16'd20905, 16'd25785, 16'd27119, 16'd39548, 16'd33575, 16'd51968, 16'd49403, 16'd59752, 16'd64338, 16'd52206, 16'd15298, 16'd13615, 16'd31085, 16'd52880, 16'd22308, 16'd35199, 16'd10050, 16'd43785, 16'd37352, 16'd38459, 16'd43879, 16'd38600, 16'd7810, 16'd50758, 16'd47680, 16'd5488});
	test_expansion(128'h21409a1d868ea44c17a5b7592ebaef87, {16'd20589, 16'd6644, 16'd44120, 16'd49952, 16'd21575, 16'd3090, 16'd34810, 16'd45600, 16'd11381, 16'd41356, 16'd65490, 16'd27535, 16'd59385, 16'd39206, 16'd33679, 16'd25964, 16'd24163, 16'd62938, 16'd43561, 16'd12509, 16'd33562, 16'd16891, 16'd42769, 16'd65285, 16'd30871, 16'd9073});
	test_expansion(128'h204f688fe0d086d93ed486b459f58cb6, {16'd39927, 16'd41593, 16'd22213, 16'd41778, 16'd63970, 16'd65101, 16'd55356, 16'd34927, 16'd36409, 16'd5386, 16'd49788, 16'd2223, 16'd47393, 16'd30840, 16'd51235, 16'd56457, 16'd41760, 16'd38609, 16'd4254, 16'd51979, 16'd57333, 16'd5136, 16'd18899, 16'd58426, 16'd37774, 16'd60814});
	test_expansion(128'h6b3acad965c4bb8131aeee7c446c6a6d, {16'd20882, 16'd14164, 16'd21293, 16'd44199, 16'd64138, 16'd57862, 16'd18742, 16'd55394, 16'd48456, 16'd48119, 16'd1390, 16'd55323, 16'd13343, 16'd43052, 16'd57097, 16'd43929, 16'd62142, 16'd53019, 16'd36703, 16'd10035, 16'd17963, 16'd48053, 16'd41338, 16'd49481, 16'd7759, 16'd53985});
	test_expansion(128'hf73571a9056c730aebd45f55b692f09d, {16'd52251, 16'd43315, 16'd19315, 16'd46340, 16'd26790, 16'd41594, 16'd51898, 16'd46224, 16'd14570, 16'd39288, 16'd55140, 16'd7913, 16'd27839, 16'd54607, 16'd14294, 16'd59724, 16'd54541, 16'd14550, 16'd14632, 16'd51398, 16'd56322, 16'd12640, 16'd12892, 16'd54725, 16'd49187, 16'd52781});
	test_expansion(128'h67cbf8469d08d96ba58b24111814ab28, {16'd34499, 16'd23672, 16'd64134, 16'd7085, 16'd44576, 16'd25221, 16'd54708, 16'd33821, 16'd2746, 16'd7080, 16'd21986, 16'd18363, 16'd54917, 16'd40522, 16'd59889, 16'd29311, 16'd53212, 16'd42486, 16'd61348, 16'd19723, 16'd19367, 16'd3009, 16'd46086, 16'd57960, 16'd14125, 16'd8444});
	test_expansion(128'he7e9cd1fa6a27c4b5718dc84ee20c318, {16'd57384, 16'd25767, 16'd39703, 16'd10779, 16'd14521, 16'd2382, 16'd37041, 16'd386, 16'd29952, 16'd47887, 16'd62838, 16'd52103, 16'd2045, 16'd53616, 16'd46090, 16'd53242, 16'd61637, 16'd57712, 16'd22339, 16'd6211, 16'd31563, 16'd52484, 16'd13740, 16'd35431, 16'd19583, 16'd55497});
	test_expansion(128'h5bc421395b5a3ea28f434eeecff6bf2b, {16'd13343, 16'd38442, 16'd31352, 16'd57191, 16'd61014, 16'd29304, 16'd61736, 16'd64351, 16'd37781, 16'd41142, 16'd50143, 16'd11867, 16'd61133, 16'd35436, 16'd34055, 16'd53696, 16'd16450, 16'd51490, 16'd22689, 16'd31296, 16'd48421, 16'd15402, 16'd39697, 16'd55830, 16'd37612, 16'd58800});
	test_expansion(128'hbf88de598438588e394c36256402a261, {16'd41374, 16'd33701, 16'd35825, 16'd28823, 16'd18052, 16'd3355, 16'd61237, 16'd29971, 16'd41769, 16'd45859, 16'd55561, 16'd48164, 16'd44812, 16'd3277, 16'd4199, 16'd27575, 16'd33356, 16'd44583, 16'd1552, 16'd18855, 16'd15567, 16'd36345, 16'd49037, 16'd188, 16'd22824, 16'd31777});
	test_expansion(128'h896dcd83b6286feb6c7710a61f8e0afe, {16'd21515, 16'd21843, 16'd23847, 16'd48427, 16'd64561, 16'd21559, 16'd25770, 16'd3668, 16'd1704, 16'd5451, 16'd29819, 16'd24452, 16'd53704, 16'd54338, 16'd46030, 16'd13923, 16'd43860, 16'd31640, 16'd26609, 16'd20560, 16'd12435, 16'd2605, 16'd34564, 16'd649, 16'd46209, 16'd40901});
	test_expansion(128'h097b0e086d63e44325f90120d657350e, {16'd15121, 16'd45383, 16'd40714, 16'd34752, 16'd8855, 16'd1832, 16'd49656, 16'd40818, 16'd31656, 16'd60794, 16'd23767, 16'd56853, 16'd54998, 16'd19783, 16'd4214, 16'd21396, 16'd12243, 16'd54483, 16'd41902, 16'd7784, 16'd23024, 16'd49529, 16'd48949, 16'd30485, 16'd22078, 16'd20847});
	test_expansion(128'h37f3c4e165b4396cae3a028d6bd45520, {16'd64736, 16'd57654, 16'd19170, 16'd59835, 16'd28646, 16'd20253, 16'd18260, 16'd40514, 16'd42887, 16'd11673, 16'd54838, 16'd10727, 16'd46979, 16'd62892, 16'd15429, 16'd44435, 16'd50639, 16'd25855, 16'd23348, 16'd50935, 16'd40455, 16'd47616, 16'd22809, 16'd21004, 16'd7445, 16'd30466});
	test_expansion(128'ha2afb22f018e8c32fd3944a64361e426, {16'd52768, 16'd45652, 16'd53102, 16'd47844, 16'd59505, 16'd65383, 16'd22184, 16'd24985, 16'd29477, 16'd4372, 16'd46013, 16'd50952, 16'd29749, 16'd54729, 16'd47249, 16'd35039, 16'd48828, 16'd58132, 16'd52677, 16'd52642, 16'd52127, 16'd44023, 16'd50634, 16'd52520, 16'd10281, 16'd3088});
	test_expansion(128'h809eb95ea239fb68103c71d1a3f2a2ff, {16'd50452, 16'd11700, 16'd7933, 16'd47473, 16'd37443, 16'd47407, 16'd20441, 16'd31338, 16'd1438, 16'd8787, 16'd58982, 16'd65295, 16'd17865, 16'd48715, 16'd8014, 16'd2841, 16'd28124, 16'd15182, 16'd312, 16'd15712, 16'd1496, 16'd558, 16'd7213, 16'd57984, 16'd55975, 16'd45895});
	test_expansion(128'hb6f96a5f7f1b610ae290c5c9028217c3, {16'd58801, 16'd15400, 16'd35391, 16'd14566, 16'd10816, 16'd49808, 16'd25074, 16'd33979, 16'd4876, 16'd13100, 16'd18274, 16'd13681, 16'd59754, 16'd35622, 16'd16366, 16'd48447, 16'd53562, 16'd26405, 16'd28776, 16'd14164, 16'd15618, 16'd43608, 16'd52031, 16'd58419, 16'd19440, 16'd43714});
	test_expansion(128'hadf552c4a35e0e7f6cbfecf485b1e8c8, {16'd26484, 16'd16178, 16'd45591, 16'd11190, 16'd26101, 16'd14259, 16'd26274, 16'd56788, 16'd78, 16'd52429, 16'd30453, 16'd15274, 16'd13217, 16'd29391, 16'd23794, 16'd16131, 16'd14080, 16'd47477, 16'd16430, 16'd62216, 16'd48547, 16'd32141, 16'd26644, 16'd56618, 16'd42587, 16'd61222});
	test_expansion(128'hbf8abc1abfeb67fd00dc15715d3d6ad9, {16'd6042, 16'd45542, 16'd19292, 16'd13905, 16'd62917, 16'd4204, 16'd30400, 16'd55435, 16'd34914, 16'd63442, 16'd15907, 16'd50602, 16'd26137, 16'd28927, 16'd10956, 16'd45829, 16'd61359, 16'd43694, 16'd6533, 16'd56070, 16'd49543, 16'd30077, 16'd338, 16'd46316, 16'd59528, 16'd31689});
	test_expansion(128'hbbe17cef7bc90fed9d6c78460e0d3a14, {16'd25010, 16'd59970, 16'd55898, 16'd54901, 16'd63437, 16'd31167, 16'd27770, 16'd49511, 16'd61303, 16'd41543, 16'd63736, 16'd9027, 16'd53114, 16'd40494, 16'd48250, 16'd9198, 16'd20885, 16'd59402, 16'd20502, 16'd4537, 16'd11243, 16'd1279, 16'd24077, 16'd24148, 16'd57832, 16'd62031});
	test_expansion(128'h5bac9baba6d4c85d07cc26a41798299b, {16'd36307, 16'd25925, 16'd32482, 16'd39673, 16'd30984, 16'd53070, 16'd62298, 16'd21294, 16'd56346, 16'd42024, 16'd35213, 16'd18518, 16'd43243, 16'd3510, 16'd20313, 16'd9944, 16'd54177, 16'd56077, 16'd43665, 16'd28460, 16'd27229, 16'd63063, 16'd9490, 16'd22646, 16'd56371, 16'd41639});
	test_expansion(128'h5d4e64ec2d351823e7b5636f4583363d, {16'd8326, 16'd7300, 16'd27097, 16'd50171, 16'd22911, 16'd65443, 16'd11103, 16'd28221, 16'd57983, 16'd448, 16'd21369, 16'd57843, 16'd8882, 16'd14031, 16'd22128, 16'd53722, 16'd34871, 16'd12555, 16'd30312, 16'd1224, 16'd50514, 16'd61228, 16'd13566, 16'd11048, 16'd65077, 16'd1228});
	test_expansion(128'hc286b7e932e84780973f195a6d11f116, {16'd63772, 16'd56755, 16'd61498, 16'd48780, 16'd9546, 16'd7716, 16'd50181, 16'd12452, 16'd10366, 16'd2398, 16'd50455, 16'd28256, 16'd34501, 16'd5848, 16'd6626, 16'd14617, 16'd3805, 16'd63450, 16'd48643, 16'd28739, 16'd43900, 16'd3232, 16'd63235, 16'd51884, 16'd14002, 16'd54444});
	test_expansion(128'h77db6616fa448c5f7893812562a24f6d, {16'd44206, 16'd18326, 16'd32405, 16'd57904, 16'd59237, 16'd5059, 16'd49107, 16'd8485, 16'd14467, 16'd44619, 16'd13271, 16'd61707, 16'd38358, 16'd34753, 16'd60140, 16'd11049, 16'd45370, 16'd47836, 16'd4642, 16'd16748, 16'd52713, 16'd50284, 16'd49672, 16'd58502, 16'd63352, 16'd59113});
	test_expansion(128'h1f223a1a4bee910cb9845334dce6c518, {16'd17269, 16'd30935, 16'd27996, 16'd47611, 16'd27317, 16'd38122, 16'd61887, 16'd60867, 16'd18047, 16'd9519, 16'd5391, 16'd3598, 16'd58740, 16'd5120, 16'd1679, 16'd33484, 16'd13603, 16'd51513, 16'd44077, 16'd24359, 16'd39122, 16'd10634, 16'd38193, 16'd24527, 16'd38019, 16'd5898});
	test_expansion(128'h1a073949ba658d9cded8b211722fee57, {16'd46278, 16'd39658, 16'd19879, 16'd55902, 16'd41035, 16'd43691, 16'd47315, 16'd31156, 16'd43468, 16'd61966, 16'd58043, 16'd61982, 16'd25148, 16'd47148, 16'd62597, 16'd48766, 16'd61061, 16'd51320, 16'd48019, 16'd55916, 16'd37556, 16'd14061, 16'd49771, 16'd62432, 16'd24723, 16'd54207});
	test_expansion(128'hdefabaeec04f8f80cb1996e8db2e97bc, {16'd5563, 16'd44199, 16'd6219, 16'd23269, 16'd32853, 16'd32095, 16'd61447, 16'd18922, 16'd55271, 16'd64737, 16'd51792, 16'd37536, 16'd13757, 16'd55790, 16'd47519, 16'd2748, 16'd63780, 16'd2847, 16'd35890, 16'd8557, 16'd19525, 16'd58827, 16'd51246, 16'd16644, 16'd581, 16'd55128});
	test_expansion(128'h9a4a43912c5753bc4778dec5480361fe, {16'd19875, 16'd37958, 16'd42458, 16'd27667, 16'd11919, 16'd8730, 16'd27901, 16'd14339, 16'd24033, 16'd57726, 16'd6528, 16'd39163, 16'd55465, 16'd31228, 16'd35986, 16'd26608, 16'd46763, 16'd34142, 16'd51902, 16'd22994, 16'd53190, 16'd29382, 16'd35858, 16'd29363, 16'd53423, 16'd37809});
	test_expansion(128'h7ffce19e67ac24e4629ae6213896c08d, {16'd33448, 16'd8170, 16'd27768, 16'd11190, 16'd56546, 16'd782, 16'd25858, 16'd25521, 16'd20820, 16'd64151, 16'd56944, 16'd59031, 16'd5444, 16'd45286, 16'd25940, 16'd17262, 16'd29278, 16'd8872, 16'd6832, 16'd56081, 16'd63613, 16'd23643, 16'd15148, 16'd46571, 16'd3305, 16'd28756});
	test_expansion(128'h63e1a478be4242e811a97b052abd8d56, {16'd49028, 16'd13842, 16'd30345, 16'd34259, 16'd19165, 16'd49944, 16'd51270, 16'd12894, 16'd34287, 16'd44557, 16'd25699, 16'd11541, 16'd19218, 16'd59455, 16'd37254, 16'd40530, 16'd4265, 16'd37158, 16'd46569, 16'd7047, 16'd14387, 16'd17360, 16'd40683, 16'd2875, 16'd51688, 16'd17397});
	test_expansion(128'h6f8866214331065c43910ea5d7ae4aab, {16'd57411, 16'd7383, 16'd38000, 16'd5583, 16'd54210, 16'd26636, 16'd51041, 16'd29178, 16'd33929, 16'd1794, 16'd34461, 16'd57377, 16'd34693, 16'd28688, 16'd22458, 16'd1684, 16'd1907, 16'd17129, 16'd41444, 16'd43718, 16'd62645, 16'd5808, 16'd32832, 16'd10149, 16'd31062, 16'd12713});
	test_expansion(128'h3da715e06540331a58ccea90a692ede9, {16'd38315, 16'd43118, 16'd10916, 16'd26451, 16'd60340, 16'd47371, 16'd14613, 16'd54228, 16'd60431, 16'd9446, 16'd34808, 16'd52310, 16'd48852, 16'd14431, 16'd25803, 16'd27820, 16'd18379, 16'd4160, 16'd53289, 16'd64872, 16'd5554, 16'd52808, 16'd40548, 16'd48427, 16'd51295, 16'd27540});
	test_expansion(128'hcda34510202f2afba0b53b8de5b8aec1, {16'd62723, 16'd546, 16'd55634, 16'd7303, 16'd7801, 16'd1039, 16'd59636, 16'd27379, 16'd8524, 16'd26621, 16'd35809, 16'd12227, 16'd48352, 16'd24244, 16'd35504, 16'd63224, 16'd17329, 16'd12946, 16'd30474, 16'd57004, 16'd34488, 16'd65456, 16'd26946, 16'd58546, 16'd44866, 16'd33334});
	test_expansion(128'h8b7e210f249cf351414b871552f11ba8, {16'd4317, 16'd12858, 16'd5899, 16'd17470, 16'd47298, 16'd12568, 16'd32291, 16'd23721, 16'd12309, 16'd51942, 16'd13961, 16'd41699, 16'd37246, 16'd9289, 16'd19975, 16'd27054, 16'd63007, 16'd62629, 16'd45999, 16'd21664, 16'd6404, 16'd42855, 16'd47033, 16'd47090, 16'd65432, 16'd63959});
	test_expansion(128'hd289f2415e0aed53ac7d60f1f0e06340, {16'd56175, 16'd18967, 16'd34124, 16'd10279, 16'd23610, 16'd39029, 16'd41357, 16'd12981, 16'd64472, 16'd34085, 16'd12161, 16'd29157, 16'd48822, 16'd29039, 16'd47978, 16'd55552, 16'd57484, 16'd7120, 16'd53231, 16'd12507, 16'd10592, 16'd47268, 16'd3109, 16'd38221, 16'd25448, 16'd17519});
	test_expansion(128'hde91358a3868562502a170d25006d1dc, {16'd22452, 16'd7775, 16'd61046, 16'd60976, 16'd14912, 16'd5247, 16'd53376, 16'd24514, 16'd37824, 16'd48730, 16'd36688, 16'd16551, 16'd51191, 16'd7633, 16'd54292, 16'd19982, 16'd11749, 16'd45518, 16'd34223, 16'd65326, 16'd9410, 16'd14757, 16'd44570, 16'd27801, 16'd58425, 16'd60601});
	test_expansion(128'h53d77657ccbc89085763a9b66d8f1329, {16'd34255, 16'd44744, 16'd15884, 16'd5183, 16'd48147, 16'd40318, 16'd36373, 16'd18489, 16'd58969, 16'd47422, 16'd58552, 16'd63366, 16'd16893, 16'd34504, 16'd37975, 16'd8535, 16'd1971, 16'd21897, 16'd7112, 16'd38912, 16'd38942, 16'd25566, 16'd50847, 16'd23950, 16'd60029, 16'd25761});
	test_expansion(128'h82b00f5f340e00c4af46d544506d55c7, {16'd55177, 16'd54700, 16'd28597, 16'd51713, 16'd50588, 16'd44411, 16'd41906, 16'd48267, 16'd27921, 16'd63105, 16'd24553, 16'd5233, 16'd27172, 16'd20421, 16'd58517, 16'd60274, 16'd19492, 16'd2155, 16'd14309, 16'd3275, 16'd61111, 16'd12684, 16'd54250, 16'd24544, 16'd26625, 16'd43795});
	test_expansion(128'h0aa03b7c7c6bd9ed93014e370745d5ee, {16'd48376, 16'd36777, 16'd57583, 16'd60804, 16'd34547, 16'd20245, 16'd15559, 16'd35577, 16'd15276, 16'd39978, 16'd4345, 16'd58682, 16'd48873, 16'd16440, 16'd38889, 16'd29336, 16'd32451, 16'd32705, 16'd22529, 16'd48304, 16'd52422, 16'd12432, 16'd61911, 16'd25250, 16'd25201, 16'd11419});
	test_expansion(128'h964e3dc7c9c41fd3ed66b113325f6810, {16'd753, 16'd57794, 16'd33577, 16'd4388, 16'd3029, 16'd2063, 16'd51523, 16'd34759, 16'd40019, 16'd25616, 16'd43146, 16'd37258, 16'd58964, 16'd47667, 16'd43479, 16'd2081, 16'd38401, 16'd5642, 16'd15314, 16'd62102, 16'd25694, 16'd56564, 16'd43138, 16'd64579, 16'd52777, 16'd21184});
	test_expansion(128'hbc185ce025856188824288c82882896f, {16'd23009, 16'd52760, 16'd20336, 16'd8703, 16'd50289, 16'd13821, 16'd19658, 16'd8391, 16'd43471, 16'd479, 16'd19540, 16'd27148, 16'd56997, 16'd51235, 16'd54689, 16'd28011, 16'd16322, 16'd7090, 16'd42075, 16'd26145, 16'd36455, 16'd63934, 16'd40866, 16'd59883, 16'd36076, 16'd54479});
	test_expansion(128'hdae8deed8808cb6ad8a407b993c1c710, {16'd15521, 16'd32691, 16'd16249, 16'd14235, 16'd45397, 16'd21473, 16'd8861, 16'd61657, 16'd42901, 16'd47963, 16'd51565, 16'd3266, 16'd16978, 16'd61183, 16'd29880, 16'd2772, 16'd22116, 16'd31137, 16'd21069, 16'd36208, 16'd46703, 16'd17840, 16'd40612, 16'd34960, 16'd2403, 16'd15843});
	test_expansion(128'h707271b32842fd98229f8db40c12aa44, {16'd3778, 16'd11446, 16'd14070, 16'd64349, 16'd23837, 16'd12103, 16'd36380, 16'd11561, 16'd59044, 16'd11394, 16'd34337, 16'd12611, 16'd43057, 16'd6421, 16'd20396, 16'd45334, 16'd52760, 16'd60498, 16'd41918, 16'd22494, 16'd23513, 16'd51272, 16'd4809, 16'd29624, 16'd49918, 16'd41449});
	test_expansion(128'h8d7c81324a92be5a0080f5a265a8aa12, {16'd6859, 16'd63652, 16'd12089, 16'd30279, 16'd21866, 16'd1867, 16'd7571, 16'd24111, 16'd55119, 16'd53128, 16'd4100, 16'd18042, 16'd52318, 16'd65012, 16'd9270, 16'd17826, 16'd55713, 16'd16701, 16'd38070, 16'd11399, 16'd39520, 16'd32942, 16'd21445, 16'd44478, 16'd15854, 16'd37250});
	test_expansion(128'hf85148b959206a10d28f09f04e5b1745, {16'd1173, 16'd8909, 16'd56487, 16'd48163, 16'd40727, 16'd35283, 16'd14143, 16'd32641, 16'd12994, 16'd19715, 16'd15615, 16'd40768, 16'd25352, 16'd40557, 16'd20464, 16'd34055, 16'd47830, 16'd6961, 16'd9876, 16'd26854, 16'd49579, 16'd6906, 16'd49960, 16'd4549, 16'd18657, 16'd1725});
	test_expansion(128'h729f14b40e489f27d36ddbdfe041fe1d, {16'd30244, 16'd64649, 16'd23322, 16'd54354, 16'd22640, 16'd42127, 16'd37131, 16'd58155, 16'd25411, 16'd13638, 16'd10094, 16'd16771, 16'd60889, 16'd12961, 16'd7246, 16'd63033, 16'd58182, 16'd17931, 16'd39783, 16'd39899, 16'd37819, 16'd168, 16'd40011, 16'd18335, 16'd61594, 16'd26280});
	test_expansion(128'ha44b923257a9b9dddf139b6ac9967701, {16'd21229, 16'd53788, 16'd43455, 16'd44423, 16'd52496, 16'd44443, 16'd15729, 16'd38497, 16'd43460, 16'd1073, 16'd1565, 16'd6224, 16'd54964, 16'd16878, 16'd50876, 16'd2206, 16'd7658, 16'd31937, 16'd27653, 16'd17413, 16'd54950, 16'd33664, 16'd22044, 16'd11105, 16'd32634, 16'd57157});
	test_expansion(128'hc703da11db9a289ed861ab0493813e9d, {16'd17386, 16'd22670, 16'd11148, 16'd65345, 16'd41164, 16'd64281, 16'd51145, 16'd28359, 16'd26792, 16'd24255, 16'd60596, 16'd58560, 16'd6631, 16'd50729, 16'd12827, 16'd62372, 16'd30700, 16'd41954, 16'd35161, 16'd9520, 16'd62397, 16'd63004, 16'd22946, 16'd50600, 16'd19104, 16'd20681});
	test_expansion(128'h10aedaf9e575d437206d61c5460f5345, {16'd12130, 16'd38574, 16'd19390, 16'd3855, 16'd54624, 16'd47745, 16'd4857, 16'd24482, 16'd15406, 16'd38124, 16'd55961, 16'd59709, 16'd34308, 16'd21103, 16'd15364, 16'd50716, 16'd25798, 16'd39517, 16'd11166, 16'd59730, 16'd45022, 16'd38554, 16'd29650, 16'd41656, 16'd36532, 16'd25848});
	test_expansion(128'h616c0eb36a1ac1c86ad3ef4d276df401, {16'd49434, 16'd63587, 16'd50151, 16'd12729, 16'd53210, 16'd21234, 16'd49687, 16'd53655, 16'd59009, 16'd59013, 16'd39992, 16'd14580, 16'd24030, 16'd50194, 16'd19028, 16'd35209, 16'd3124, 16'd39276, 16'd29749, 16'd29860, 16'd15192, 16'd29839, 16'd1351, 16'd4217, 16'd4159, 16'd2020});
	test_expansion(128'h6502c2def783567bdb577002608a593b, {16'd20588, 16'd55786, 16'd33704, 16'd39891, 16'd13239, 16'd13779, 16'd35038, 16'd50357, 16'd5108, 16'd6111, 16'd13440, 16'd21011, 16'd55597, 16'd19930, 16'd53995, 16'd47039, 16'd25036, 16'd24953, 16'd45670, 16'd46936, 16'd51257, 16'd63428, 16'd45807, 16'd22244, 16'd14858, 16'd62420});
	test_expansion(128'he8a24b0951998f32668a62177ee42b24, {16'd17693, 16'd8035, 16'd16612, 16'd18258, 16'd55317, 16'd11602, 16'd48362, 16'd47064, 16'd37468, 16'd52589, 16'd28767, 16'd15951, 16'd17578, 16'd24825, 16'd56056, 16'd16706, 16'd64882, 16'd35417, 16'd36573, 16'd33455, 16'd40951, 16'd27777, 16'd57370, 16'd51844, 16'd55438, 16'd34877});
	test_expansion(128'h1e19ad0ba5ea12a36d8c1fa43218b269, {16'd54012, 16'd2067, 16'd58959, 16'd9430, 16'd3638, 16'd45348, 16'd2922, 16'd47421, 16'd27392, 16'd8643, 16'd58181, 16'd27770, 16'd64046, 16'd35747, 16'd3526, 16'd22721, 16'd11000, 16'd26712, 16'd4436, 16'd6632, 16'd45050, 16'd214, 16'd28372, 16'd56981, 16'd25827, 16'd51932});
	test_expansion(128'he4cbed06612d7e3b51932f29e957a434, {16'd59078, 16'd62935, 16'd60525, 16'd4690, 16'd14231, 16'd8984, 16'd45249, 16'd15608, 16'd14752, 16'd60341, 16'd38082, 16'd30856, 16'd43385, 16'd64000, 16'd27504, 16'd13209, 16'd57356, 16'd4276, 16'd58074, 16'd45536, 16'd62396, 16'd18717, 16'd13109, 16'd43361, 16'd9698, 16'd27410});
	test_expansion(128'h9b8c98ad987a4e7240ff02ff95c1cf6e, {16'd51953, 16'd44532, 16'd11012, 16'd60485, 16'd34437, 16'd55148, 16'd25476, 16'd56699, 16'd1251, 16'd16961, 16'd28185, 16'd10838, 16'd58442, 16'd7744, 16'd10334, 16'd29465, 16'd32429, 16'd46295, 16'd32463, 16'd13088, 16'd60261, 16'd54635, 16'd20560, 16'd36845, 16'd25445, 16'd54160});
	test_expansion(128'hecdb822c8c9e5131352edfd67f1c77c7, {16'd42327, 16'd5564, 16'd41213, 16'd9525, 16'd29402, 16'd60448, 16'd27951, 16'd58303, 16'd16848, 16'd9165, 16'd61153, 16'd26723, 16'd21659, 16'd41016, 16'd33673, 16'd58795, 16'd39309, 16'd58464, 16'd55999, 16'd13796, 16'd61847, 16'd44694, 16'd6455, 16'd58726, 16'd41426, 16'd46160});
	test_expansion(128'h5242f5d279f1711dd38656cb88d60690, {16'd30748, 16'd55273, 16'd64174, 16'd3354, 16'd6096, 16'd11036, 16'd55170, 16'd19900, 16'd31004, 16'd23028, 16'd31100, 16'd16724, 16'd42285, 16'd57832, 16'd61714, 16'd23962, 16'd55893, 16'd45512, 16'd43784, 16'd18207, 16'd17966, 16'd21663, 16'd43442, 16'd3759, 16'd28341, 16'd38856});
	test_expansion(128'hf778ab9d3e55e6eb4bccd8f381d8a20d, {16'd18185, 16'd22591, 16'd55348, 16'd35107, 16'd42592, 16'd55350, 16'd46659, 16'd60816, 16'd46384, 16'd5994, 16'd8457, 16'd64145, 16'd25974, 16'd55897, 16'd28027, 16'd61801, 16'd35716, 16'd33874, 16'd55927, 16'd17992, 16'd53209, 16'd54669, 16'd14027, 16'd21931, 16'd43098, 16'd28651});
	test_expansion(128'h1d9e166da4733986eec8b91bbc38a594, {16'd49882, 16'd13718, 16'd8631, 16'd57222, 16'd22178, 16'd5140, 16'd52999, 16'd20714, 16'd30753, 16'd35369, 16'd1626, 16'd15320, 16'd18885, 16'd40583, 16'd65396, 16'd17802, 16'd23732, 16'd52806, 16'd21207, 16'd3005, 16'd15670, 16'd14681, 16'd56735, 16'd41662, 16'd61102, 16'd970});
	test_expansion(128'hc610058f0b26ed4cda9ee43ba682ed8c, {16'd20599, 16'd21286, 16'd15773, 16'd62930, 16'd38652, 16'd31840, 16'd37928, 16'd16799, 16'd15754, 16'd44043, 16'd7572, 16'd31296, 16'd39024, 16'd59011, 16'd12137, 16'd46773, 16'd16500, 16'd29054, 16'd41156, 16'd58288, 16'd31451, 16'd57006, 16'd50318, 16'd28225, 16'd933, 16'd20157});
	test_expansion(128'h7597b8777dcd86ea0c6b1d6deef91193, {16'd23791, 16'd3351, 16'd40339, 16'd41379, 16'd53759, 16'd63716, 16'd51094, 16'd27983, 16'd40477, 16'd62676, 16'd44798, 16'd63952, 16'd63374, 16'd15762, 16'd8502, 16'd44424, 16'd54922, 16'd60318, 16'd11063, 16'd47736, 16'd42908, 16'd22114, 16'd28661, 16'd29776, 16'd35167, 16'd4287});
	test_expansion(128'h6713028870c7c25aa4e2ab7525e83639, {16'd45163, 16'd39012, 16'd11828, 16'd53054, 16'd2741, 16'd3429, 16'd11957, 16'd53024, 16'd3029, 16'd9727, 16'd32666, 16'd56435, 16'd63867, 16'd24088, 16'd43138, 16'd49667, 16'd46166, 16'd44085, 16'd56104, 16'd24553, 16'd50718, 16'd21441, 16'd15985, 16'd62501, 16'd35144, 16'd42138});
	test_expansion(128'hfac5c63b4ac817afdf7f76482d1fc4f9, {16'd60865, 16'd54933, 16'd10419, 16'd43267, 16'd44342, 16'd49372, 16'd26472, 16'd62734, 16'd35082, 16'd35534, 16'd28982, 16'd2981, 16'd3484, 16'd3716, 16'd16669, 16'd43746, 16'd3916, 16'd40945, 16'd31729, 16'd14357, 16'd6083, 16'd26560, 16'd33228, 16'd42918, 16'd16878, 16'd54531});
	test_expansion(128'h5a02333e1a70af0c73a99fe4ab4c9334, {16'd5226, 16'd25361, 16'd9468, 16'd37812, 16'd30008, 16'd64543, 16'd55917, 16'd2330, 16'd35998, 16'd63362, 16'd19069, 16'd57707, 16'd1725, 16'd3699, 16'd9408, 16'd26865, 16'd56200, 16'd40970, 16'd54043, 16'd24910, 16'd55793, 16'd39867, 16'd11547, 16'd43316, 16'd50449, 16'd28236});
	test_expansion(128'h92c1138ca4cca0b876e54556ee2e282c, {16'd60427, 16'd57780, 16'd29384, 16'd5726, 16'd28430, 16'd25478, 16'd62488, 16'd11030, 16'd54672, 16'd35041, 16'd54954, 16'd40491, 16'd21559, 16'd29883, 16'd64359, 16'd41948, 16'd50054, 16'd3147, 16'd5247, 16'd8325, 16'd53404, 16'd24961, 16'd65519, 16'd33845, 16'd41345, 16'd29042});
	test_expansion(128'h2b3174226f3589315690171b23794594, {16'd11069, 16'd47449, 16'd48501, 16'd969, 16'd28081, 16'd44586, 16'd39203, 16'd5313, 16'd13914, 16'd20126, 16'd35337, 16'd5158, 16'd11623, 16'd22830, 16'd6668, 16'd5937, 16'd30055, 16'd51250, 16'd8240, 16'd62010, 16'd24790, 16'd51843, 16'd27862, 16'd40581, 16'd42296, 16'd6879});
	test_expansion(128'he40c4a8a4bd183fcd5eb7f74a6c09e94, {16'd47115, 16'd37576, 16'd60680, 16'd53213, 16'd16253, 16'd633, 16'd40225, 16'd61507, 16'd35854, 16'd62865, 16'd48137, 16'd62448, 16'd3766, 16'd20535, 16'd37670, 16'd44709, 16'd38764, 16'd57502, 16'd41140, 16'd21542, 16'd19947, 16'd41116, 16'd64952, 16'd63092, 16'd58531, 16'd46293});
	test_expansion(128'h1084f8b0e52bab8dfb7fdaa823f34d0d, {16'd28136, 16'd15141, 16'd22718, 16'd4111, 16'd42444, 16'd14264, 16'd19954, 16'd32536, 16'd54836, 16'd34116, 16'd61921, 16'd6498, 16'd62135, 16'd7704, 16'd39936, 16'd19153, 16'd6635, 16'd63415, 16'd2868, 16'd41854, 16'd26478, 16'd21486, 16'd12948, 16'd49475, 16'd47089, 16'd19370});
	test_expansion(128'hff0cffeb7b6fdb005374a3e7c03bc06b, {16'd2314, 16'd4528, 16'd4746, 16'd56739, 16'd37630, 16'd23618, 16'd43736, 16'd1801, 16'd25771, 16'd60480, 16'd64776, 16'd38571, 16'd22561, 16'd7267, 16'd46174, 16'd832, 16'd9581, 16'd22401, 16'd1150, 16'd62115, 16'd19737, 16'd64363, 16'd36570, 16'd59548, 16'd56463, 16'd962});
	test_expansion(128'h2af08b7d3594567f813e3b134cffcd14, {16'd47191, 16'd32411, 16'd62026, 16'd33105, 16'd40869, 16'd28505, 16'd28647, 16'd6004, 16'd11583, 16'd10494, 16'd9607, 16'd10957, 16'd36095, 16'd32943, 16'd39964, 16'd39631, 16'd33509, 16'd56896, 16'd3864, 16'd6703, 16'd56585, 16'd61186, 16'd50130, 16'd22791, 16'd28445, 16'd7043});
	test_expansion(128'hdefc2743d7e841c3fbd0d265fa1f7fbe, {16'd31611, 16'd18485, 16'd53589, 16'd49919, 16'd36544, 16'd8494, 16'd45350, 16'd5446, 16'd61979, 16'd47448, 16'd154, 16'd61670, 16'd3465, 16'd6970, 16'd22151, 16'd21133, 16'd29948, 16'd3597, 16'd53301, 16'd21286, 16'd30746, 16'd3453, 16'd3107, 16'd30459, 16'd24978, 16'd15405});
	test_expansion(128'h9eb0230a894f7e88c5b9b2ef94a3ab1b, {16'd10171, 16'd38366, 16'd35153, 16'd28716, 16'd10960, 16'd34619, 16'd61220, 16'd36272, 16'd7170, 16'd3716, 16'd45420, 16'd25696, 16'd58437, 16'd52376, 16'd46030, 16'd50462, 16'd10752, 16'd9523, 16'd65133, 16'd30981, 16'd49366, 16'd18336, 16'd62618, 16'd43229, 16'd45077, 16'd4781});
	test_expansion(128'h85d6d62c581fcb351660e88d4ce01dd0, {16'd58545, 16'd22216, 16'd8460, 16'd56681, 16'd53448, 16'd40822, 16'd3871, 16'd26318, 16'd28527, 16'd33372, 16'd26748, 16'd42403, 16'd25850, 16'd63511, 16'd53660, 16'd45239, 16'd47338, 16'd38020, 16'd46656, 16'd35197, 16'd59661, 16'd2921, 16'd25329, 16'd58228, 16'd7467, 16'd36160});
	test_expansion(128'hb94fc77db58ab6445c5be5cdfa3de061, {16'd6862, 16'd32, 16'd43713, 16'd27018, 16'd12770, 16'd7813, 16'd10584, 16'd35935, 16'd20401, 16'd13760, 16'd42092, 16'd43655, 16'd17803, 16'd21734, 16'd58087, 16'd59308, 16'd29178, 16'd36386, 16'd6894, 16'd23720, 16'd15257, 16'd49241, 16'd16358, 16'd12247, 16'd22659, 16'd11256});
	test_expansion(128'h56352d546bc7d2e19e16abfd9377e503, {16'd35585, 16'd19226, 16'd37504, 16'd26977, 16'd22718, 16'd42865, 16'd31203, 16'd57108, 16'd27571, 16'd27363, 16'd40169, 16'd41053, 16'd58237, 16'd52929, 16'd29506, 16'd35866, 16'd22465, 16'd35816, 16'd57023, 16'd49387, 16'd21161, 16'd32375, 16'd4235, 16'd60574, 16'd1356, 16'd39894});
	test_expansion(128'h34d05d9ef4f1c7765f32abf746926504, {16'd19486, 16'd64958, 16'd3426, 16'd25064, 16'd6977, 16'd11835, 16'd40648, 16'd52963, 16'd14173, 16'd27059, 16'd38756, 16'd59603, 16'd47682, 16'd60025, 16'd32146, 16'd20795, 16'd12002, 16'd7126, 16'd31939, 16'd14438, 16'd51248, 16'd22130, 16'd7262, 16'd48817, 16'd59910, 16'd56513});
	test_expansion(128'h84eb095d9a7280b01406e6ab3c6717fa, {16'd62871, 16'd37787, 16'd62841, 16'd48061, 16'd57273, 16'd12560, 16'd34472, 16'd65, 16'd23958, 16'd24337, 16'd4772, 16'd24288, 16'd25217, 16'd57278, 16'd12206, 16'd4546, 16'd52714, 16'd917, 16'd58247, 16'd31326, 16'd22223, 16'd48678, 16'd14703, 16'd15075, 16'd27780, 16'd26399});
	test_expansion(128'hb348040e75e15feb6700dd2d60b65f3f, {16'd57275, 16'd33801, 16'd21079, 16'd1368, 16'd55238, 16'd65285, 16'd31553, 16'd19410, 16'd4991, 16'd38072, 16'd38060, 16'd45662, 16'd48403, 16'd45565, 16'd28653, 16'd21311, 16'd46737, 16'd25679, 16'd58537, 16'd22140, 16'd38440, 16'd31587, 16'd65402, 16'd47697, 16'd19635, 16'd10231});
	test_expansion(128'h5e5bf380f8e57c74268a56a125681b36, {16'd1981, 16'd24719, 16'd30602, 16'd26306, 16'd37297, 16'd52533, 16'd47680, 16'd5303, 16'd14598, 16'd12331, 16'd50833, 16'd8283, 16'd14492, 16'd36541, 16'd26357, 16'd58568, 16'd39473, 16'd27094, 16'd17032, 16'd54541, 16'd9446, 16'd29095, 16'd13199, 16'd51261, 16'd48414, 16'd50814});
	test_expansion(128'hba293cb8b28cab55b794532d67a20fdf, {16'd39425, 16'd54172, 16'd21500, 16'd33318, 16'd28431, 16'd1989, 16'd8977, 16'd775, 16'd49947, 16'd49026, 16'd16346, 16'd16262, 16'd8481, 16'd65309, 16'd5544, 16'd33839, 16'd8096, 16'd32282, 16'd10136, 16'd9820, 16'd24963, 16'd42763, 16'd9425, 16'd57886, 16'd32520, 16'd29514});
	test_expansion(128'hc25463184f962fec6f286644ec40ecc7, {16'd14679, 16'd31563, 16'd7979, 16'd61678, 16'd51290, 16'd61083, 16'd19825, 16'd51477, 16'd65430, 16'd16601, 16'd36884, 16'd13713, 16'd54780, 16'd52923, 16'd25605, 16'd35519, 16'd18996, 16'd25161, 16'd6512, 16'd50791, 16'd54600, 16'd11349, 16'd53730, 16'd36504, 16'd48056, 16'd13613});
	test_expansion(128'h6c950044e1e8baef9cd9efcca0d83186, {16'd64214, 16'd56724, 16'd60439, 16'd9266, 16'd46029, 16'd10606, 16'd32612, 16'd43021, 16'd5165, 16'd28927, 16'd45501, 16'd7753, 16'd29936, 16'd40101, 16'd56857, 16'd5248, 16'd30820, 16'd48119, 16'd42678, 16'd16927, 16'd38279, 16'd60276, 16'd19592, 16'd64046, 16'd37279, 16'd28888});
	test_expansion(128'h9857ab94078f2549788b1e25e1b04295, {16'd47779, 16'd55978, 16'd16603, 16'd29335, 16'd59059, 16'd5904, 16'd24796, 16'd14438, 16'd4487, 16'd41510, 16'd40667, 16'd37572, 16'd44879, 16'd58758, 16'd21100, 16'd58952, 16'd65437, 16'd3954, 16'd60466, 16'd44253, 16'd21749, 16'd12252, 16'd24483, 16'd59013, 16'd163, 16'd2163});
	test_expansion(128'ha013c784d8115fd54412283c23c6a1f0, {16'd54804, 16'd64881, 16'd35242, 16'd30182, 16'd7294, 16'd62970, 16'd42575, 16'd17654, 16'd742, 16'd25592, 16'd55968, 16'd37620, 16'd61409, 16'd142, 16'd9112, 16'd44251, 16'd45083, 16'd35218, 16'd52557, 16'd46695, 16'd30958, 16'd46133, 16'd11088, 16'd35180, 16'd19845, 16'd54253});
	test_expansion(128'hc891d38ed692a88daddb576e167998d9, {16'd31597, 16'd2715, 16'd50755, 16'd60508, 16'd26297, 16'd26526, 16'd49883, 16'd52087, 16'd20625, 16'd62534, 16'd31320, 16'd49382, 16'd45124, 16'd42711, 16'd27078, 16'd15893, 16'd22821, 16'd58789, 16'd8391, 16'd9074, 16'd56091, 16'd12831, 16'd29927, 16'd6520, 16'd21540, 16'd25997});
	test_expansion(128'h33fa576da7c3ad30360ac5012e20b409, {16'd53165, 16'd50594, 16'd39137, 16'd50015, 16'd51233, 16'd20435, 16'd5173, 16'd36446, 16'd15858, 16'd31847, 16'd52659, 16'd2631, 16'd42618, 16'd4986, 16'd42592, 16'd30186, 16'd43009, 16'd27086, 16'd20107, 16'd61266, 16'd61183, 16'd46057, 16'd64138, 16'd17119, 16'd40773, 16'd25677});
	test_expansion(128'hf071df65f5a2fe6fa7635c609ddfca4e, {16'd50813, 16'd53873, 16'd30300, 16'd52873, 16'd41071, 16'd1101, 16'd45716, 16'd58252, 16'd38292, 16'd30149, 16'd48057, 16'd63974, 16'd64127, 16'd41956, 16'd52078, 16'd28786, 16'd45944, 16'd5195, 16'd27359, 16'd18514, 16'd44600, 16'd4569, 16'd40689, 16'd37805, 16'd23979, 16'd2987});
	test_expansion(128'h0e78b0924da11dcb23d454002698f18e, {16'd4796, 16'd56254, 16'd50632, 16'd24108, 16'd13292, 16'd55281, 16'd40385, 16'd21620, 16'd53457, 16'd19357, 16'd17522, 16'd22480, 16'd25514, 16'd19935, 16'd11524, 16'd24181, 16'd20061, 16'd34465, 16'd35221, 16'd38175, 16'd10521, 16'd31418, 16'd59280, 16'd27451, 16'd60659, 16'd49916});
	test_expansion(128'hc83c8b536793cd87d2478b61a85096f3, {16'd12542, 16'd15604, 16'd17958, 16'd44274, 16'd33470, 16'd34926, 16'd46959, 16'd18624, 16'd63783, 16'd60589, 16'd48662, 16'd29793, 16'd23820, 16'd30632, 16'd24155, 16'd31237, 16'd19076, 16'd59586, 16'd4177, 16'd51406, 16'd41483, 16'd24140, 16'd18030, 16'd6145, 16'd40484, 16'd12814});
	test_expansion(128'hd1c1dc6c88d1a90f6a20ec98d163f7b7, {16'd9935, 16'd52108, 16'd39607, 16'd56140, 16'd20537, 16'd19855, 16'd5262, 16'd65030, 16'd22662, 16'd11849, 16'd21928, 16'd35879, 16'd31625, 16'd4272, 16'd5102, 16'd19248, 16'd2795, 16'd37423, 16'd34326, 16'd50164, 16'd2445, 16'd21981, 16'd5398, 16'd31532, 16'd31997, 16'd10510});
	test_expansion(128'h864f509811285106c4b2177c14c87620, {16'd30940, 16'd26645, 16'd35482, 16'd56377, 16'd45202, 16'd22847, 16'd51263, 16'd49983, 16'd56782, 16'd25829, 16'd18368, 16'd51620, 16'd9955, 16'd54985, 16'd57185, 16'd42192, 16'd49813, 16'd12486, 16'd57617, 16'd50379, 16'd22308, 16'd59065, 16'd34765, 16'd8802, 16'd3465, 16'd39490});
	test_expansion(128'h65886bb59678d239977e2a442d3af7a4, {16'd64400, 16'd52642, 16'd45657, 16'd36070, 16'd17865, 16'd10671, 16'd32424, 16'd2154, 16'd9027, 16'd14564, 16'd28065, 16'd51625, 16'd61539, 16'd18297, 16'd15999, 16'd34674, 16'd17573, 16'd63823, 16'd41083, 16'd7245, 16'd54799, 16'd33280, 16'd12678, 16'd4388, 16'd41391, 16'd7821});
	test_expansion(128'h3e06ad7065e886124077b97d9d925ede, {16'd64234, 16'd59641, 16'd64711, 16'd61548, 16'd45753, 16'd15316, 16'd23303, 16'd34986, 16'd31898, 16'd48566, 16'd4114, 16'd5879, 16'd23708, 16'd11237, 16'd64724, 16'd49729, 16'd38124, 16'd41614, 16'd39606, 16'd51421, 16'd10185, 16'd57155, 16'd23409, 16'd33168, 16'd27205, 16'd15737});
	test_expansion(128'h55420e5012938d5f8716fa419826a5af, {16'd11298, 16'd22363, 16'd47284, 16'd17427, 16'd60457, 16'd57875, 16'd19029, 16'd6133, 16'd19213, 16'd8225, 16'd20901, 16'd39812, 16'd4000, 16'd64015, 16'd33370, 16'd29482, 16'd24441, 16'd35274, 16'd12382, 16'd35830, 16'd33614, 16'd60373, 16'd25781, 16'd3574, 16'd43835, 16'd54256});
	test_expansion(128'hf6252fc07cedf849d8d5b83c8931f14a, {16'd2225, 16'd31094, 16'd3177, 16'd22951, 16'd20341, 16'd14956, 16'd21830, 16'd39710, 16'd28383, 16'd3932, 16'd3083, 16'd48759, 16'd53335, 16'd14863, 16'd59327, 16'd24241, 16'd20939, 16'd42856, 16'd33900, 16'd39919, 16'd19329, 16'd338, 16'd43382, 16'd5583, 16'd42665, 16'd5958});
	test_expansion(128'hc1a73e165c847f83e8964330976ad3b5, {16'd37981, 16'd47252, 16'd61933, 16'd27489, 16'd36349, 16'd58768, 16'd11598, 16'd26655, 16'd37883, 16'd39030, 16'd10358, 16'd50339, 16'd20206, 16'd29131, 16'd14346, 16'd43396, 16'd9454, 16'd52487, 16'd50159, 16'd33983, 16'd44035, 16'd32383, 16'd39241, 16'd17, 16'd40851, 16'd58138});
	test_expansion(128'h373f9b76c021012411e7723b0926477b, {16'd65236, 16'd42672, 16'd52378, 16'd46500, 16'd38029, 16'd17374, 16'd30092, 16'd5779, 16'd63865, 16'd24461, 16'd18940, 16'd30819, 16'd10335, 16'd34754, 16'd46017, 16'd8538, 16'd33952, 16'd27325, 16'd46042, 16'd63573, 16'd43983, 16'd39660, 16'd53655, 16'd62100, 16'd55235, 16'd37559});
	test_expansion(128'h0c40ce7dc8c0c3f22781fd9b2745e6c2, {16'd26569, 16'd11079, 16'd45792, 16'd31694, 16'd20949, 16'd3749, 16'd13715, 16'd45337, 16'd44308, 16'd40082, 16'd32697, 16'd43599, 16'd35550, 16'd19474, 16'd55306, 16'd8093, 16'd36304, 16'd37411, 16'd58552, 16'd3159, 16'd11374, 16'd2153, 16'd19382, 16'd54968, 16'd42159, 16'd60922});
	test_expansion(128'h1c3b9d91dc9c008ed507d14234eb2ad5, {16'd39062, 16'd22629, 16'd28610, 16'd47929, 16'd732, 16'd22990, 16'd54008, 16'd56705, 16'd33137, 16'd12505, 16'd30681, 16'd20543, 16'd58798, 16'd40710, 16'd33671, 16'd23573, 16'd28295, 16'd46044, 16'd24499, 16'd8870, 16'd10943, 16'd45707, 16'd33536, 16'd1951, 16'd44838, 16'd52310});
	test_expansion(128'hfd8de115e2cdddff30a343d12bab0c8b, {16'd65209, 16'd11402, 16'd35013, 16'd52578, 16'd13892, 16'd44225, 16'd21964, 16'd25040, 16'd56050, 16'd23410, 16'd60201, 16'd61046, 16'd58529, 16'd17, 16'd9163, 16'd19487, 16'd50254, 16'd61762, 16'd10475, 16'd47724, 16'd33275, 16'd51377, 16'd38068, 16'd6680, 16'd52757, 16'd48249});
	test_expansion(128'h93e8f7c74ddd19fd6610c5e93ac7d43a, {16'd20270, 16'd50762, 16'd52033, 16'd2292, 16'd1541, 16'd33754, 16'd57948, 16'd37947, 16'd14503, 16'd23803, 16'd52457, 16'd17370, 16'd36015, 16'd63959, 16'd45297, 16'd44255, 16'd1829, 16'd44504, 16'd54941, 16'd28227, 16'd61489, 16'd24862, 16'd89, 16'd33036, 16'd62220, 16'd25983});
	test_expansion(128'h78b1ab446c764c6943eaf017700077df, {16'd56411, 16'd13399, 16'd5928, 16'd63806, 16'd52870, 16'd35991, 16'd25764, 16'd61628, 16'd2123, 16'd24358, 16'd32288, 16'd9548, 16'd7573, 16'd61243, 16'd5254, 16'd4994, 16'd54590, 16'd56954, 16'd59516, 16'd20776, 16'd60888, 16'd19749, 16'd27143, 16'd35925, 16'd64242, 16'd62970});
	test_expansion(128'h1bcd3123f56b75da665e8bbb2657beb4, {16'd8415, 16'd24153, 16'd16176, 16'd8076, 16'd30170, 16'd12652, 16'd46235, 16'd27528, 16'd54060, 16'd43503, 16'd61342, 16'd43427, 16'd24778, 16'd28973, 16'd58048, 16'd6560, 16'd41878, 16'd60675, 16'd19613, 16'd61439, 16'd24338, 16'd5563, 16'd41601, 16'd8500, 16'd33475, 16'd41416});
	test_expansion(128'h849664f507151d097302c899e86d5ed2, {16'd32603, 16'd50818, 16'd3912, 16'd58075, 16'd32759, 16'd2061, 16'd12092, 16'd53430, 16'd37800, 16'd10449, 16'd27630, 16'd63296, 16'd59181, 16'd30968, 16'd8016, 16'd4548, 16'd31008, 16'd59841, 16'd63773, 16'd45639, 16'd12391, 16'd57955, 16'd61426, 16'd1901, 16'd30805, 16'd35929});
	test_expansion(128'h4ea80f0e335aa558762b4ee4143d9e9a, {16'd47452, 16'd32309, 16'd52246, 16'd62099, 16'd39244, 16'd23020, 16'd2048, 16'd50156, 16'd65345, 16'd39208, 16'd56872, 16'd9021, 16'd24784, 16'd58351, 16'd5862, 16'd50818, 16'd6246, 16'd48525, 16'd33924, 16'd45051, 16'd26588, 16'd56837, 16'd53062, 16'd35995, 16'd43773, 16'd27921});
	test_expansion(128'hc70bfacc31c6398cdce0510b9c9ade00, {16'd12095, 16'd55078, 16'd53146, 16'd58308, 16'd6523, 16'd2741, 16'd20967, 16'd46157, 16'd3126, 16'd24484, 16'd1168, 16'd42299, 16'd9718, 16'd6653, 16'd7508, 16'd59586, 16'd38655, 16'd62909, 16'd34676, 16'd17837, 16'd37740, 16'd47914, 16'd25558, 16'd29911, 16'd46400, 16'd53932});
	test_expansion(128'hddfb67fd010271d2e3b090d3e935fc54, {16'd35257, 16'd17502, 16'd62468, 16'd30644, 16'd7139, 16'd17144, 16'd55228, 16'd2748, 16'd17112, 16'd60543, 16'd60115, 16'd29343, 16'd38275, 16'd36656, 16'd33850, 16'd50465, 16'd2383, 16'd7132, 16'd42276, 16'd15791, 16'd12359, 16'd40326, 16'd54790, 16'd49985, 16'd26523, 16'd22474});
	test_expansion(128'h0f51cca47b7f98abc713d953f3d66b87, {16'd31052, 16'd5371, 16'd37789, 16'd49774, 16'd36466, 16'd37657, 16'd27441, 16'd35131, 16'd44921, 16'd63992, 16'd36457, 16'd4134, 16'd36961, 16'd58308, 16'd42012, 16'd9195, 16'd11790, 16'd22039, 16'd52538, 16'd6968, 16'd51005, 16'd1355, 16'd39091, 16'd7673, 16'd31072, 16'd49481});
	test_expansion(128'h8900d3959d7cc52b2d9d4165e498d95a, {16'd15883, 16'd11042, 16'd53457, 16'd64679, 16'd38914, 16'd30560, 16'd58733, 16'd1962, 16'd51825, 16'd47910, 16'd18659, 16'd1795, 16'd13900, 16'd58098, 16'd40062, 16'd55528, 16'd5276, 16'd24142, 16'd27669, 16'd24067, 16'd48443, 16'd58539, 16'd30689, 16'd52384, 16'd34528, 16'd40618});
	test_expansion(128'he81a564ca532239ae3a84f4ef637be71, {16'd48472, 16'd22906, 16'd31400, 16'd15659, 16'd48162, 16'd547, 16'd20047, 16'd60705, 16'd47958, 16'd21262, 16'd47678, 16'd25563, 16'd24183, 16'd2207, 16'd20522, 16'd17133, 16'd60846, 16'd11460, 16'd31101, 16'd13798, 16'd1643, 16'd33124, 16'd21817, 16'd6273, 16'd7635, 16'd24677});
	test_expansion(128'h791509b54f37c25998b77916644b279b, {16'd33292, 16'd8240, 16'd18753, 16'd48990, 16'd11297, 16'd46783, 16'd7609, 16'd52272, 16'd19933, 16'd32607, 16'd29362, 16'd40411, 16'd58117, 16'd3417, 16'd24858, 16'd2451, 16'd33979, 16'd8746, 16'd1286, 16'd13767, 16'd59200, 16'd56265, 16'd38895, 16'd20538, 16'd37462, 16'd47273});
	test_expansion(128'h755cd8330836d541b565e73807936c8e, {16'd43105, 16'd40178, 16'd51874, 16'd9265, 16'd12886, 16'd51110, 16'd43255, 16'd6848, 16'd12282, 16'd22526, 16'd27228, 16'd46870, 16'd60615, 16'd59661, 16'd36445, 16'd20839, 16'd4090, 16'd15054, 16'd25845, 16'd37557, 16'd25816, 16'd18484, 16'd33149, 16'd48990, 16'd15257, 16'd23423});
	test_expansion(128'hbd9fa17555c4fce39a3679bb2f56ec1e, {16'd47062, 16'd6358, 16'd667, 16'd51550, 16'd20821, 16'd27392, 16'd61685, 16'd30618, 16'd50674, 16'd21194, 16'd60540, 16'd36184, 16'd34281, 16'd19633, 16'd8467, 16'd53042, 16'd43976, 16'd60748, 16'd37730, 16'd12436, 16'd6633, 16'd35343, 16'd47305, 16'd48412, 16'd47915, 16'd14761});
	test_expansion(128'h981ecd169f234f208a4cadee0931a796, {16'd51496, 16'd33486, 16'd23870, 16'd7751, 16'd30589, 16'd6957, 16'd11594, 16'd25082, 16'd33700, 16'd4902, 16'd22176, 16'd33659, 16'd14152, 16'd31199, 16'd62102, 16'd49434, 16'd52890, 16'd30233, 16'd20762, 16'd28377, 16'd1875, 16'd41558, 16'd27922, 16'd26035, 16'd34681, 16'd52038});
	test_expansion(128'hcc94ce95fac513e47dd8129f9bd43c8b, {16'd9490, 16'd51437, 16'd18966, 16'd688, 16'd39785, 16'd25583, 16'd18751, 16'd344, 16'd11458, 16'd25551, 16'd12196, 16'd13852, 16'd52226, 16'd38322, 16'd7151, 16'd35306, 16'd11916, 16'd10628, 16'd20472, 16'd4372, 16'd15555, 16'd38782, 16'd49869, 16'd57346, 16'd39647, 16'd1592});
	test_expansion(128'h4ff7f2bf08650fdbeb803badf5cb419b, {16'd28835, 16'd32202, 16'd4256, 16'd4140, 16'd14894, 16'd13494, 16'd3245, 16'd11946, 16'd62915, 16'd633, 16'd10581, 16'd4736, 16'd31268, 16'd44451, 16'd58433, 16'd33173, 16'd58870, 16'd49966, 16'd5996, 16'd1636, 16'd50027, 16'd49772, 16'd1151, 16'd4243, 16'd33118, 16'd50877});
	test_expansion(128'hb2845054412819f818432cbba2425c66, {16'd54626, 16'd30428, 16'd28463, 16'd46387, 16'd9115, 16'd11096, 16'd3621, 16'd62350, 16'd49517, 16'd55894, 16'd26621, 16'd58933, 16'd31810, 16'd40172, 16'd12869, 16'd40479, 16'd63940, 16'd45377, 16'd2822, 16'd33823, 16'd49925, 16'd31395, 16'd3947, 16'd20601, 16'd18890, 16'd32526});
	test_expansion(128'hfcc38ea097a47f55a033938d6bc8e672, {16'd6963, 16'd28702, 16'd55299, 16'd42465, 16'd33055, 16'd46477, 16'd29693, 16'd28419, 16'd50566, 16'd8948, 16'd51843, 16'd5968, 16'd21710, 16'd37126, 16'd32266, 16'd17994, 16'd46012, 16'd40605, 16'd38877, 16'd50087, 16'd13215, 16'd21113, 16'd42183, 16'd30874, 16'd1761, 16'd27167});
	test_expansion(128'h90aac02c499d0a7d90f0f09c6778e96e, {16'd17637, 16'd54882, 16'd37809, 16'd62755, 16'd24690, 16'd55126, 16'd43747, 16'd44407, 16'd24057, 16'd61486, 16'd4650, 16'd13974, 16'd57887, 16'd36458, 16'd57383, 16'd13333, 16'd52943, 16'd44260, 16'd9669, 16'd31774, 16'd37268, 16'd53282, 16'd48128, 16'd46524, 16'd39588, 16'd23965});
	test_expansion(128'h8c231dcd813777f290d75da6acbeb65b, {16'd44733, 16'd41328, 16'd12191, 16'd28609, 16'd51105, 16'd33747, 16'd34010, 16'd43734, 16'd37244, 16'd6819, 16'd59888, 16'd62239, 16'd50979, 16'd12448, 16'd35252, 16'd50993, 16'd9919, 16'd24212, 16'd45403, 16'd24277, 16'd47533, 16'd4981, 16'd31331, 16'd52156, 16'd43917, 16'd38766});
	test_expansion(128'h7af41c8640b35cf547971fb73ed1f540, {16'd39162, 16'd32851, 16'd54072, 16'd25810, 16'd31094, 16'd14804, 16'd50992, 16'd27357, 16'd46674, 16'd23053, 16'd55871, 16'd2063, 16'd45796, 16'd43472, 16'd49747, 16'd58287, 16'd11525, 16'd29818, 16'd52686, 16'd39335, 16'd21374, 16'd41708, 16'd61962, 16'd60886, 16'd34806, 16'd41762});
	test_expansion(128'hfeffa6db54fbbd0694552bbbe17f9987, {16'd9017, 16'd57444, 16'd50294, 16'd53866, 16'd12735, 16'd23402, 16'd62955, 16'd38407, 16'd33812, 16'd55347, 16'd25188, 16'd29331, 16'd53065, 16'd63642, 16'd35105, 16'd24398, 16'd39482, 16'd41856, 16'd18189, 16'd10512, 16'd18395, 16'd13754, 16'd7439, 16'd64643, 16'd54549, 16'd19821});
	test_expansion(128'h0fc9c40458f44f3184c24ce83c93a95e, {16'd56234, 16'd49757, 16'd56009, 16'd39181, 16'd56800, 16'd30816, 16'd56370, 16'd53332, 16'd48188, 16'd10828, 16'd2119, 16'd18435, 16'd20506, 16'd42985, 16'd10919, 16'd22390, 16'd20370, 16'd63349, 16'd25261, 16'd9713, 16'd29820, 16'd51909, 16'd47202, 16'd27345, 16'd31391, 16'd59618});
	test_expansion(128'h7cd1988a8bc25e0d22920c9de0b9df98, {16'd17475, 16'd28765, 16'd9404, 16'd13578, 16'd62146, 16'd12434, 16'd32485, 16'd50747, 16'd35344, 16'd41955, 16'd51342, 16'd37373, 16'd13234, 16'd35234, 16'd60392, 16'd30985, 16'd48275, 16'd38183, 16'd58988, 16'd16735, 16'd7857, 16'd55444, 16'd7094, 16'd25404, 16'd49363, 16'd7762});
	test_expansion(128'h85ed88f18cbbc6a84d1ebc858109d11c, {16'd38737, 16'd54845, 16'd12895, 16'd19437, 16'd29693, 16'd13378, 16'd15393, 16'd62378, 16'd37718, 16'd29504, 16'd2801, 16'd4923, 16'd4644, 16'd30325, 16'd46036, 16'd6173, 16'd20316, 16'd33780, 16'd25921, 16'd49599, 16'd15791, 16'd49339, 16'd2107, 16'd12327, 16'd65084, 16'd10364});
	test_expansion(128'haba5a4b72850bea9177a75b20ad6ed6a, {16'd28364, 16'd31359, 16'd9496, 16'd31260, 16'd27588, 16'd41732, 16'd60913, 16'd52623, 16'd22142, 16'd49132, 16'd44764, 16'd3952, 16'd19336, 16'd8330, 16'd40760, 16'd59483, 16'd32459, 16'd11820, 16'd23782, 16'd62389, 16'd39346, 16'd6308, 16'd60743, 16'd49709, 16'd52994, 16'd23220});
	test_expansion(128'h6417ca900f75b6564db01704ed260205, {16'd16516, 16'd43531, 16'd51010, 16'd52396, 16'd41983, 16'd4070, 16'd18526, 16'd65415, 16'd35108, 16'd30409, 16'd59345, 16'd38490, 16'd5052, 16'd22878, 16'd10890, 16'd9650, 16'd25789, 16'd56267, 16'd47203, 16'd16190, 16'd23835, 16'd63384, 16'd13867, 16'd29237, 16'd11397, 16'd33420});
	test_expansion(128'h9daab857dde8ac4950a7bf0e204ca778, {16'd16110, 16'd14629, 16'd1210, 16'd39289, 16'd33245, 16'd6537, 16'd24555, 16'd145, 16'd47895, 16'd31944, 16'd19981, 16'd32409, 16'd58700, 16'd39918, 16'd32452, 16'd4290, 16'd20409, 16'd15422, 16'd40928, 16'd58167, 16'd8772, 16'd27113, 16'd45280, 16'd59053, 16'd39976, 16'd41311});
	test_expansion(128'hceebedcbcb8a63162ae68998dab3a12b, {16'd50105, 16'd5848, 16'd54757, 16'd21999, 16'd41746, 16'd1142, 16'd2396, 16'd56640, 16'd49417, 16'd16659, 16'd38566, 16'd37319, 16'd20073, 16'd5136, 16'd6749, 16'd24224, 16'd65300, 16'd14668, 16'd10372, 16'd13587, 16'd46674, 16'd3819, 16'd43255, 16'd20100, 16'd50856, 16'd25371});
	test_expansion(128'hab918446cd6f57df32ef93deee7c6f8a, {16'd13570, 16'd12838, 16'd64826, 16'd4285, 16'd52609, 16'd13316, 16'd58736, 16'd6439, 16'd61268, 16'd21802, 16'd25675, 16'd50320, 16'd50788, 16'd14121, 16'd13305, 16'd50740, 16'd32807, 16'd10736, 16'd1421, 16'd44757, 16'd25776, 16'd58697, 16'd33803, 16'd17123, 16'd41146, 16'd23873});
	test_expansion(128'h558f3f74a18e0432cb5e916d17dd35d0, {16'd22850, 16'd51052, 16'd37356, 16'd27199, 16'd64596, 16'd50017, 16'd25885, 16'd27454, 16'd11322, 16'd49641, 16'd59552, 16'd20956, 16'd54048, 16'd23366, 16'd47993, 16'd44214, 16'd39690, 16'd54434, 16'd55013, 16'd33007, 16'd9099, 16'd36466, 16'd55096, 16'd12488, 16'd26088, 16'd13555});
	test_expansion(128'h6807c60763c7c7b2c0c0407a80de00e6, {16'd18245, 16'd12817, 16'd31007, 16'd46225, 16'd23358, 16'd11313, 16'd38827, 16'd45936, 16'd49276, 16'd6533, 16'd21710, 16'd42939, 16'd11018, 16'd11419, 16'd62666, 16'd63654, 16'd30282, 16'd2483, 16'd24861, 16'd6589, 16'd7590, 16'd2741, 16'd11145, 16'd55798, 16'd3736, 16'd20859});
	test_expansion(128'hb66791329693da8d2ab0a909c8861429, {16'd31964, 16'd35742, 16'd62280, 16'd15646, 16'd56154, 16'd18588, 16'd40023, 16'd64668, 16'd47458, 16'd50877, 16'd10393, 16'd26769, 16'd55738, 16'd36370, 16'd61557, 16'd18731, 16'd37847, 16'd20996, 16'd6058, 16'd52478, 16'd64688, 16'd31585, 16'd39928, 16'd753, 16'd46669, 16'd35313});
	test_expansion(128'h56dea350d25f38e2f98520afa357d951, {16'd19487, 16'd28531, 16'd23531, 16'd59959, 16'd27266, 16'd26426, 16'd46544, 16'd17302, 16'd10668, 16'd34903, 16'd59633, 16'd60277, 16'd37433, 16'd58876, 16'd5388, 16'd22104, 16'd34834, 16'd18717, 16'd48884, 16'd41184, 16'd23866, 16'd51141, 16'd10567, 16'd39981, 16'd36624, 16'd26089});
	test_expansion(128'he86a65f12c0a04de69024ba8b702efff, {16'd24912, 16'd59880, 16'd51314, 16'd8853, 16'd36514, 16'd44443, 16'd51986, 16'd49085, 16'd17179, 16'd36224, 16'd1493, 16'd50343, 16'd41932, 16'd54051, 16'd9112, 16'd7932, 16'd16457, 16'd11616, 16'd46562, 16'd7728, 16'd38711, 16'd64024, 16'd59433, 16'd63001, 16'd6985, 16'd40144});
	test_expansion(128'h24810706aab0968792a3adb8b94c3980, {16'd25150, 16'd42090, 16'd65267, 16'd9439, 16'd54047, 16'd25689, 16'd8345, 16'd58955, 16'd38229, 16'd18928, 16'd27452, 16'd62237, 16'd40132, 16'd10733, 16'd50727, 16'd46213, 16'd15898, 16'd58535, 16'd27734, 16'd49314, 16'd22122, 16'd31969, 16'd4859, 16'd2296, 16'd5649, 16'd41128});
	test_expansion(128'h212bcba42b7758ca807b68c3a313cdeb, {16'd14995, 16'd43274, 16'd32877, 16'd24846, 16'd63041, 16'd5612, 16'd56252, 16'd42876, 16'd15757, 16'd23412, 16'd62308, 16'd7724, 16'd22649, 16'd22800, 16'd25594, 16'd33389, 16'd62542, 16'd32942, 16'd9434, 16'd35854, 16'd38759, 16'd22674, 16'd329, 16'd59147, 16'd42087, 16'd11580});
	test_expansion(128'hf2a89975ffb143145b1918c477e13c4a, {16'd62393, 16'd28623, 16'd43125, 16'd15873, 16'd19629, 16'd13900, 16'd22615, 16'd56378, 16'd57863, 16'd36366, 16'd16353, 16'd12139, 16'd54950, 16'd54689, 16'd61634, 16'd18542, 16'd49323, 16'd55324, 16'd45535, 16'd3700, 16'd32259, 16'd38535, 16'd62518, 16'd3385, 16'd26366, 16'd15475});
	test_expansion(128'h567b95bfb98dfd60a07bd09a6bbc4b9f, {16'd45259, 16'd63428, 16'd24925, 16'd12827, 16'd45715, 16'd18678, 16'd15183, 16'd31872, 16'd11717, 16'd35942, 16'd7195, 16'd12321, 16'd49298, 16'd44674, 16'd4, 16'd56631, 16'd21647, 16'd22511, 16'd32331, 16'd45416, 16'd44741, 16'd18503, 16'd44522, 16'd24630, 16'd45474, 16'd49127});
	test_expansion(128'he39dd95ce69b1fe9a03d3240f7ac9521, {16'd26662, 16'd34700, 16'd52568, 16'd47371, 16'd1321, 16'd42037, 16'd14526, 16'd91, 16'd29361, 16'd1132, 16'd27927, 16'd15664, 16'd2872, 16'd52708, 16'd43415, 16'd5110, 16'd34654, 16'd29688, 16'd36041, 16'd23689, 16'd12641, 16'd63903, 16'd2496, 16'd61175, 16'd40363, 16'd40612});
	test_expansion(128'h2d6a7c34839b415d7fce359113858e5c, {16'd21224, 16'd25207, 16'd28394, 16'd12784, 16'd1928, 16'd15270, 16'd64741, 16'd63589, 16'd36015, 16'd53357, 16'd39660, 16'd22171, 16'd35047, 16'd50595, 16'd47279, 16'd26546, 16'd10921, 16'd44179, 16'd4199, 16'd58108, 16'd14128, 16'd49272, 16'd28071, 16'd38048, 16'd9837, 16'd19883});
	test_expansion(128'ha43cf8dce3f74084b7d9f249e6087f5e, {16'd48205, 16'd39522, 16'd1705, 16'd11357, 16'd29750, 16'd34801, 16'd41451, 16'd42685, 16'd21510, 16'd33664, 16'd59143, 16'd7696, 16'd13276, 16'd62589, 16'd65158, 16'd4256, 16'd48546, 16'd60768, 16'd23279, 16'd33497, 16'd44890, 16'd22261, 16'd20341, 16'd17151, 16'd39189, 16'd45547});
	test_expansion(128'hf4a6707445f708c5d2a762280895f3ae, {16'd30832, 16'd60332, 16'd9727, 16'd31013, 16'd52996, 16'd13526, 16'd44009, 16'd21067, 16'd23269, 16'd63182, 16'd21301, 16'd51798, 16'd19402, 16'd57990, 16'd44913, 16'd17749, 16'd7679, 16'd51227, 16'd35534, 16'd1390, 16'd34728, 16'd33731, 16'd48467, 16'd26427, 16'd23487, 16'd42985});
	test_expansion(128'h050289ee06f8e2c6a44af231e94ab0fe, {16'd21118, 16'd58270, 16'd61295, 16'd26724, 16'd43359, 16'd40623, 16'd371, 16'd1427, 16'd41219, 16'd30059, 16'd58007, 16'd5274, 16'd27222, 16'd62151, 16'd63843, 16'd45676, 16'd58968, 16'd32754, 16'd45264, 16'd5548, 16'd11744, 16'd550, 16'd13526, 16'd36270, 16'd45510, 16'd3350});
	test_expansion(128'h5750961863b1c5d1a806ba834021496d, {16'd42979, 16'd28956, 16'd31039, 16'd65401, 16'd13250, 16'd12399, 16'd38958, 16'd29407, 16'd59178, 16'd2730, 16'd17488, 16'd57683, 16'd58675, 16'd3056, 16'd36968, 16'd26324, 16'd18933, 16'd52524, 16'd35710, 16'd12499, 16'd23116, 16'd60534, 16'd27245, 16'd58843, 16'd47122, 16'd54604});
	test_expansion(128'hd45229bd6880acec77fb1ad0409bbeb7, {16'd1602, 16'd52235, 16'd7738, 16'd11894, 16'd42652, 16'd37174, 16'd49097, 16'd52822, 16'd42468, 16'd15447, 16'd43478, 16'd60364, 16'd59716, 16'd33284, 16'd2807, 16'd63167, 16'd4490, 16'd7770, 16'd38470, 16'd47718, 16'd26259, 16'd48598, 16'd26110, 16'd56112, 16'd2754, 16'd65442});
	test_expansion(128'hd3368a05315f4e4627afcfd51509aba1, {16'd50789, 16'd57169, 16'd38704, 16'd55303, 16'd16175, 16'd57481, 16'd22284, 16'd13252, 16'd7167, 16'd29567, 16'd38246, 16'd3217, 16'd461, 16'd27015, 16'd39622, 16'd24809, 16'd61427, 16'd22359, 16'd62841, 16'd55811, 16'd6113, 16'd59664, 16'd27273, 16'd65371, 16'd62155, 16'd50618});
	test_expansion(128'h92b047eefa99ea11241eb4a370a77aa3, {16'd42567, 16'd50536, 16'd59824, 16'd29070, 16'd504, 16'd49223, 16'd16620, 16'd7556, 16'd684, 16'd13320, 16'd26453, 16'd20580, 16'd2098, 16'd59048, 16'd4509, 16'd40475, 16'd18196, 16'd51587, 16'd64002, 16'd48778, 16'd28125, 16'd39156, 16'd27738, 16'd63708, 16'd40655, 16'd37008});
	test_expansion(128'hcd9bb6b22d7c58f33ac5bac1e515c2b5, {16'd35696, 16'd29427, 16'd55306, 16'd52000, 16'd30073, 16'd57892, 16'd55952, 16'd29242, 16'd29885, 16'd10394, 16'd58588, 16'd52918, 16'd41249, 16'd12600, 16'd50157, 16'd33975, 16'd26080, 16'd8957, 16'd44537, 16'd152, 16'd62065, 16'd26149, 16'd55000, 16'd65189, 16'd41768, 16'd48251});
	test_expansion(128'h6c6342bd4efb74722922cc4bb7112387, {16'd30401, 16'd19584, 16'd51181, 16'd16920, 16'd63553, 16'd2883, 16'd28013, 16'd4554, 16'd16896, 16'd58858, 16'd54531, 16'd42721, 16'd11191, 16'd16305, 16'd29552, 16'd54237, 16'd7774, 16'd19422, 16'd39509, 16'd49004, 16'd48347, 16'd43471, 16'd60521, 16'd54727, 16'd37836, 16'd35804});
	test_expansion(128'hd59f0119a5d3779128b42a7b2b618f1e, {16'd33186, 16'd39987, 16'd55510, 16'd31584, 16'd25252, 16'd19866, 16'd17962, 16'd63295, 16'd43823, 16'd34259, 16'd56553, 16'd18972, 16'd8809, 16'd65406, 16'd41895, 16'd23995, 16'd49346, 16'd50622, 16'd58918, 16'd18471, 16'd42716, 16'd56440, 16'd60479, 16'd28843, 16'd29133, 16'd59605});
	test_expansion(128'h93bcd72c69dd32c44620d81b20c11170, {16'd45917, 16'd50796, 16'd19815, 16'd45614, 16'd33142, 16'd37081, 16'd9381, 16'd30822, 16'd44192, 16'd2830, 16'd59319, 16'd64405, 16'd64450, 16'd45235, 16'd31142, 16'd36266, 16'd42082, 16'd50264, 16'd2792, 16'd25470, 16'd36402, 16'd32647, 16'd24046, 16'd10828, 16'd3098, 16'd57187});
	test_expansion(128'he95b5eb445bc68bae22f70e2f576bc47, {16'd53951, 16'd37623, 16'd21015, 16'd47302, 16'd63896, 16'd9670, 16'd16103, 16'd20897, 16'd30741, 16'd21263, 16'd53395, 16'd4678, 16'd31598, 16'd34058, 16'd55225, 16'd10952, 16'd51574, 16'd25146, 16'd21151, 16'd12195, 16'd46479, 16'd37727, 16'd2482, 16'd46860, 16'd50876, 16'd16802});
	test_expansion(128'h89e22ffae434618d1095d977c8458b14, {16'd31183, 16'd36632, 16'd57310, 16'd6664, 16'd54937, 16'd33737, 16'd842, 16'd44372, 16'd62780, 16'd1729, 16'd64243, 16'd59571, 16'd33978, 16'd16712, 16'd50771, 16'd33246, 16'd3527, 16'd1146, 16'd58056, 16'd17178, 16'd17729, 16'd2049, 16'd16883, 16'd9489, 16'd15710, 16'd20832});
	test_expansion(128'h85ce6e7d95b88aa0dbff455ba0dfa4b5, {16'd62143, 16'd44533, 16'd43814, 16'd53414, 16'd62971, 16'd5131, 16'd5211, 16'd20991, 16'd19331, 16'd6141, 16'd15949, 16'd59726, 16'd65200, 16'd33188, 16'd46195, 16'd31207, 16'd49595, 16'd31255, 16'd18802, 16'd49227, 16'd61043, 16'd57338, 16'd60592, 16'd44215, 16'd31190, 16'd15592});
	test_expansion(128'ha4bd827a81be824a80e7d0b8c2bc4865, {16'd5282, 16'd5532, 16'd56933, 16'd11053, 16'd63019, 16'd7082, 16'd9053, 16'd20426, 16'd34595, 16'd31931, 16'd59311, 16'd45234, 16'd56033, 16'd54753, 16'd57895, 16'd25189, 16'd60221, 16'd24087, 16'd29782, 16'd29765, 16'd12990, 16'd53070, 16'd9160, 16'd18274, 16'd46685, 16'd38116});
	test_expansion(128'h17120579c0103871b44d9138bed4f8c6, {16'd45654, 16'd37754, 16'd38979, 16'd22859, 16'd23930, 16'd16015, 16'd1650, 16'd9479, 16'd35701, 16'd14507, 16'd19818, 16'd63808, 16'd26900, 16'd13124, 16'd27325, 16'd17991, 16'd3498, 16'd12817, 16'd24694, 16'd41966, 16'd17194, 16'd1930, 16'd11694, 16'd5572, 16'd58429, 16'd25140});
	test_expansion(128'hbb55c118b07d159e0373bb531a27bcd9, {16'd24335, 16'd33512, 16'd37370, 16'd48759, 16'd20421, 16'd29976, 16'd62734, 16'd10080, 16'd36573, 16'd54848, 16'd34531, 16'd50544, 16'd60531, 16'd46055, 16'd43614, 16'd6623, 16'd35941, 16'd15594, 16'd30464, 16'd52309, 16'd1144, 16'd22495, 16'd56332, 16'd8473, 16'd46386, 16'd12660});
	test_expansion(128'h27b4afbb759f41fb0ebff152195d8c36, {16'd9235, 16'd28769, 16'd12061, 16'd17034, 16'd6867, 16'd5949, 16'd10149, 16'd37897, 16'd33806, 16'd13526, 16'd40465, 16'd31631, 16'd64295, 16'd34337, 16'd34748, 16'd34142, 16'd18311, 16'd44620, 16'd40168, 16'd39951, 16'd54948, 16'd2886, 16'd36638, 16'd46966, 16'd25352, 16'd11515});
	test_expansion(128'h0d3b18e8c97ca61cc55a7962c53eba6f, {16'd843, 16'd14040, 16'd28708, 16'd18633, 16'd31538, 16'd10788, 16'd61358, 16'd57601, 16'd46812, 16'd61493, 16'd44463, 16'd65471, 16'd61401, 16'd59291, 16'd42321, 16'd23743, 16'd52477, 16'd37459, 16'd62740, 16'd27808, 16'd18183, 16'd4348, 16'd64778, 16'd43172, 16'd24779, 16'd15079});
	test_expansion(128'hc98ab947d70324711281a661c9b03070, {16'd52935, 16'd19249, 16'd11316, 16'd14373, 16'd65125, 16'd15147, 16'd27130, 16'd49569, 16'd56656, 16'd50536, 16'd20638, 16'd29938, 16'd61761, 16'd15926, 16'd62705, 16'd56476, 16'd22175, 16'd46092, 16'd59932, 16'd59214, 16'd55893, 16'd32215, 16'd23433, 16'd26637, 16'd53175, 16'd60971});
	test_expansion(128'h9cc13dbb82a5c9e741a18b2a56708013, {16'd48327, 16'd497, 16'd34094, 16'd35089, 16'd47475, 16'd56078, 16'd58327, 16'd58406, 16'd651, 16'd17253, 16'd28668, 16'd33795, 16'd21286, 16'd42483, 16'd20706, 16'd48872, 16'd887, 16'd30078, 16'd44569, 16'd16532, 16'd18736, 16'd11271, 16'd55710, 16'd28624, 16'd37685, 16'd59743});
	test_expansion(128'hd055fb854160dccf889a536eee9dbe9f, {16'd5057, 16'd43650, 16'd10390, 16'd54287, 16'd31431, 16'd60369, 16'd47297, 16'd56063, 16'd3616, 16'd6876, 16'd57946, 16'd8771, 16'd57552, 16'd1736, 16'd25503, 16'd37324, 16'd34773, 16'd43626, 16'd44838, 16'd2943, 16'd35103, 16'd75, 16'd57358, 16'd53372, 16'd34975, 16'd13407});
	test_expansion(128'h17e0ff478a2688879df7e2e9ac990354, {16'd41486, 16'd49643, 16'd54457, 16'd34276, 16'd18749, 16'd43959, 16'd55893, 16'd18443, 16'd43106, 16'd59226, 16'd10170, 16'd32334, 16'd33647, 16'd57391, 16'd20521, 16'd31782, 16'd57661, 16'd56615, 16'd61777, 16'd8239, 16'd21727, 16'd34781, 16'd2516, 16'd16076, 16'd6658, 16'd5215});
	test_expansion(128'h978ed886d5913300e3d248538c563337, {16'd53103, 16'd1397, 16'd31591, 16'd12234, 16'd30370, 16'd36237, 16'd65479, 16'd58374, 16'd27404, 16'd44547, 16'd12581, 16'd18124, 16'd43249, 16'd39475, 16'd11927, 16'd50620, 16'd1298, 16'd31337, 16'd2889, 16'd27480, 16'd35103, 16'd48968, 16'd20226, 16'd7533, 16'd63257, 16'd60627});
	test_expansion(128'hcfb4c45115f8593cb2378c449f12e41d, {16'd42302, 16'd5331, 16'd8983, 16'd26466, 16'd58685, 16'd10365, 16'd56086, 16'd40730, 16'd12291, 16'd8064, 16'd7362, 16'd23931, 16'd64696, 16'd64511, 16'd57032, 16'd62855, 16'd38639, 16'd3999, 16'd27790, 16'd36065, 16'd17413, 16'd359, 16'd38630, 16'd50053, 16'd60970, 16'd61174});
	test_expansion(128'hf2a8c676c9b5b476f68c9fcb2b395f8d, {16'd41863, 16'd9272, 16'd6497, 16'd7799, 16'd47895, 16'd37644, 16'd45590, 16'd19590, 16'd64196, 16'd42610, 16'd51902, 16'd25274, 16'd47087, 16'd272, 16'd58516, 16'd48058, 16'd55119, 16'd63595, 16'd53817, 16'd55900, 16'd9520, 16'd54859, 16'd27873, 16'd12907, 16'd12596, 16'd28875});
	test_expansion(128'hc457d0c5ecc9207433df90e2b80b1f98, {16'd4352, 16'd15583, 16'd42383, 16'd22800, 16'd7640, 16'd27875, 16'd60625, 16'd13716, 16'd54002, 16'd50704, 16'd13365, 16'd57033, 16'd43344, 16'd65273, 16'd1931, 16'd62679, 16'd40724, 16'd41531, 16'd64533, 16'd5784, 16'd59104, 16'd12037, 16'd45398, 16'd7268, 16'd22633, 16'd30051});
	test_expansion(128'h2d76fa927525de46f554903693cd9a8d, {16'd25843, 16'd50751, 16'd51508, 16'd58700, 16'd33556, 16'd55418, 16'd11939, 16'd54937, 16'd59855, 16'd22829, 16'd45077, 16'd41106, 16'd63363, 16'd258, 16'd59729, 16'd42943, 16'd22811, 16'd5737, 16'd17333, 16'd15232, 16'd6847, 16'd25316, 16'd42985, 16'd63384, 16'd14100, 16'd49506});
	test_expansion(128'h01d766994d1f561130415965acc7520a, {16'd22240, 16'd38381, 16'd30055, 16'd20617, 16'd42588, 16'd62656, 16'd37406, 16'd34612, 16'd57870, 16'd43112, 16'd48121, 16'd61349, 16'd50272, 16'd9545, 16'd35026, 16'd25595, 16'd38408, 16'd49385, 16'd64397, 16'd32017, 16'd31256, 16'd12674, 16'd16414, 16'd48808, 16'd29723, 16'd10480});
	test_expansion(128'he9e658d72a004c54d1324feac635fcfe, {16'd48058, 16'd65168, 16'd37990, 16'd44674, 16'd53052, 16'd41528, 16'd29302, 16'd13975, 16'd51185, 16'd30494, 16'd46722, 16'd38296, 16'd19285, 16'd9822, 16'd26427, 16'd25086, 16'd41399, 16'd29267, 16'd55945, 16'd51097, 16'd38315, 16'd42428, 16'd46299, 16'd13656, 16'd61252, 16'd11906});
	test_expansion(128'h82f29c99ce0b6c59ebfb3725a85471c2, {16'd8874, 16'd34590, 16'd18445, 16'd29046, 16'd32837, 16'd19001, 16'd35910, 16'd52989, 16'd23578, 16'd25999, 16'd18395, 16'd42884, 16'd25761, 16'd55574, 16'd53598, 16'd35587, 16'd29341, 16'd61, 16'd12495, 16'd34905, 16'd34597, 16'd54026, 16'd6154, 16'd36991, 16'd61088, 16'd24601});
	test_expansion(128'h3031e23a7db153c73a0ffbdbaf795545, {16'd37983, 16'd60781, 16'd18484, 16'd65378, 16'd13749, 16'd25313, 16'd6018, 16'd31549, 16'd45331, 16'd15070, 16'd55778, 16'd50601, 16'd3799, 16'd28213, 16'd6268, 16'd28477, 16'd27192, 16'd4828, 16'd22150, 16'd50899, 16'd44750, 16'd43000, 16'd63435, 16'd13960, 16'd32490, 16'd39348});
	test_expansion(128'h751d391c8f2e7caff5147627630a8789, {16'd1485, 16'd22115, 16'd52617, 16'd32790, 16'd20341, 16'd33402, 16'd7084, 16'd65022, 16'd47206, 16'd43123, 16'd54366, 16'd18724, 16'd63789, 16'd37770, 16'd27005, 16'd25830, 16'd40032, 16'd6846, 16'd14726, 16'd12593, 16'd19521, 16'd3954, 16'd59588, 16'd30292, 16'd32681, 16'd17143});
	test_expansion(128'h3d0685c946582dbc4b729595ccf92b42, {16'd5249, 16'd12925, 16'd13745, 16'd18079, 16'd29888, 16'd15153, 16'd19007, 16'd19165, 16'd30403, 16'd56697, 16'd13021, 16'd7096, 16'd2665, 16'd13760, 16'd51007, 16'd38596, 16'd4431, 16'd27510, 16'd45834, 16'd41144, 16'd49315, 16'd15619, 16'd42428, 16'd5890, 16'd19992, 16'd28276});
	test_expansion(128'h495c00048d9bdb8070e161c2c18a1a99, {16'd51469, 16'd43605, 16'd40294, 16'd29617, 16'd12209, 16'd2479, 16'd32652, 16'd18508, 16'd42169, 16'd61995, 16'd17651, 16'd25138, 16'd6699, 16'd9535, 16'd41407, 16'd59029, 16'd12021, 16'd19472, 16'd58272, 16'd16986, 16'd553, 16'd60546, 16'd27338, 16'd46217, 16'd63280, 16'd60624});
	test_expansion(128'h36c94eb395ec5cd9cc2ee9589ff6acb9, {16'd556, 16'd51635, 16'd35589, 16'd54996, 16'd52047, 16'd34531, 16'd18280, 16'd836, 16'd45080, 16'd13196, 16'd963, 16'd61619, 16'd41359, 16'd262, 16'd49697, 16'd49451, 16'd9936, 16'd32282, 16'd58431, 16'd23915, 16'd18903, 16'd26779, 16'd60741, 16'd22973, 16'd42869, 16'd42188});
	test_expansion(128'hbf2310e486c544053e291780766a1a68, {16'd23700, 16'd1208, 16'd15228, 16'd19333, 16'd16042, 16'd5234, 16'd49399, 16'd25028, 16'd1970, 16'd39107, 16'd58413, 16'd63555, 16'd11128, 16'd59505, 16'd2263, 16'd12085, 16'd47614, 16'd26380, 16'd50889, 16'd3665, 16'd37870, 16'd9874, 16'd34646, 16'd54747, 16'd17045, 16'd8323});
	test_expansion(128'h649f3298440048745eb7886b34135ccd, {16'd34544, 16'd43189, 16'd31528, 16'd29957, 16'd48682, 16'd26267, 16'd2304, 16'd1294, 16'd21148, 16'd47351, 16'd50310, 16'd56445, 16'd12052, 16'd50911, 16'd58029, 16'd37971, 16'd38668, 16'd52163, 16'd10990, 16'd28330, 16'd49067, 16'd4500, 16'd1280, 16'd56196, 16'd55232, 16'd60145});
	test_expansion(128'h5a8dce3a8957d8c10f05114abaee3d41, {16'd29442, 16'd44337, 16'd17463, 16'd29451, 16'd34664, 16'd25362, 16'd59372, 16'd4362, 16'd5975, 16'd26463, 16'd22706, 16'd19642, 16'd29557, 16'd38294, 16'd47838, 16'd57494, 16'd11205, 16'd21992, 16'd40060, 16'd41831, 16'd6338, 16'd61248, 16'd53173, 16'd34718, 16'd1795, 16'd47938});
	test_expansion(128'hc9f16c3c48bbbcd6cc9e76a895037718, {16'd26981, 16'd25593, 16'd2182, 16'd63388, 16'd53843, 16'd14580, 16'd18830, 16'd50076, 16'd18439, 16'd22820, 16'd61075, 16'd43195, 16'd17425, 16'd59131, 16'd7420, 16'd63023, 16'd42395, 16'd39225, 16'd37913, 16'd59763, 16'd13087, 16'd20270, 16'd42725, 16'd40407, 16'd25547, 16'd1843});
	test_expansion(128'hb197c936004fef187153d4e140bb5ebe, {16'd43910, 16'd11918, 16'd37983, 16'd61622, 16'd28474, 16'd9028, 16'd60598, 16'd31865, 16'd41253, 16'd40188, 16'd60248, 16'd64258, 16'd38630, 16'd57087, 16'd52366, 16'd58128, 16'd51234, 16'd26336, 16'd35350, 16'd9706, 16'd29799, 16'd16214, 16'd4432, 16'd54269, 16'd1333, 16'd1830});
	test_expansion(128'h65c2e5be50c2b8dfc8e402a19916ab0b, {16'd53923, 16'd46613, 16'd5405, 16'd46398, 16'd32989, 16'd14420, 16'd11745, 16'd29379, 16'd37802, 16'd18289, 16'd46166, 16'd25168, 16'd45549, 16'd24513, 16'd42478, 16'd42845, 16'd46084, 16'd54156, 16'd3717, 16'd60917, 16'd1460, 16'd11063, 16'd29839, 16'd19639, 16'd9268, 16'd38055});
	test_expansion(128'h7f3b20754b74cd64524f8d9607f80a3c, {16'd10904, 16'd39246, 16'd54663, 16'd4798, 16'd49633, 16'd35890, 16'd17727, 16'd57831, 16'd62781, 16'd32833, 16'd49883, 16'd10673, 16'd28095, 16'd12235, 16'd3325, 16'd47472, 16'd25299, 16'd53319, 16'd54674, 16'd241, 16'd42926, 16'd30987, 16'd14535, 16'd19610, 16'd61905, 16'd59440});
	test_expansion(128'h144716cfde6b99fa675b006b95e1e75b, {16'd7541, 16'd54337, 16'd2302, 16'd28194, 16'd37498, 16'd19496, 16'd37651, 16'd46499, 16'd22851, 16'd1113, 16'd62505, 16'd65250, 16'd34671, 16'd3968, 16'd8955, 16'd14222, 16'd60006, 16'd6730, 16'd61523, 16'd61584, 16'd31161, 16'd59889, 16'd18433, 16'd53533, 16'd25953, 16'd46446});
	test_expansion(128'h77b2a3751568f07deefa08a0dac29c76, {16'd15157, 16'd42558, 16'd29651, 16'd52464, 16'd36566, 16'd1675, 16'd62257, 16'd61321, 16'd13477, 16'd60120, 16'd57058, 16'd34216, 16'd58132, 16'd21158, 16'd6859, 16'd23662, 16'd60646, 16'd39002, 16'd40753, 16'd6239, 16'd26720, 16'd42377, 16'd10487, 16'd35390, 16'd17561, 16'd21021});
	test_expansion(128'ha502c546fbba63230ae0f1b36d9f1785, {16'd38275, 16'd28601, 16'd32612, 16'd62157, 16'd60168, 16'd47239, 16'd19681, 16'd18661, 16'd22767, 16'd61069, 16'd30726, 16'd27163, 16'd21685, 16'd62446, 16'd22696, 16'd1200, 16'd24339, 16'd56014, 16'd2468, 16'd22297, 16'd11247, 16'd40225, 16'd29423, 16'd63847, 16'd5551, 16'd15059});
	test_expansion(128'h0cf337dde3e23cec1cc78d0b4a3f07b3, {16'd38825, 16'd62042, 16'd3564, 16'd65219, 16'd61468, 16'd34864, 16'd62000, 16'd48532, 16'd36605, 16'd5558, 16'd23454, 16'd25127, 16'd716, 16'd18651, 16'd60245, 16'd60153, 16'd40990, 16'd3163, 16'd47173, 16'd30730, 16'd21695, 16'd10117, 16'd8502, 16'd36221, 16'd15665, 16'd56192});
	test_expansion(128'h5f4c48d012f27b116f7d8edc7f584628, {16'd18998, 16'd65271, 16'd30167, 16'd34252, 16'd42491, 16'd11374, 16'd33010, 16'd59924, 16'd58176, 16'd315, 16'd40849, 16'd39696, 16'd33139, 16'd33728, 16'd13344, 16'd10196, 16'd19913, 16'd20342, 16'd30018, 16'd61767, 16'd40969, 16'd7760, 16'd30170, 16'd58802, 16'd52755, 16'd32341});
	test_expansion(128'h472c007d9784fe7487fab70aa05eeb81, {16'd24401, 16'd34259, 16'd3332, 16'd63184, 16'd47024, 16'd30978, 16'd15385, 16'd10297, 16'd43754, 16'd13250, 16'd46580, 16'd51423, 16'd46078, 16'd54017, 16'd41580, 16'd44284, 16'd37636, 16'd22743, 16'd20281, 16'd37564, 16'd44090, 16'd46445, 16'd48296, 16'd5648, 16'd5224, 16'd43156});
	test_expansion(128'hc2db17d1e37574c0fd3611a94675ae6d, {16'd40339, 16'd40063, 16'd22235, 16'd44799, 16'd10252, 16'd56313, 16'd23386, 16'd37528, 16'd15658, 16'd7163, 16'd1034, 16'd9566, 16'd63252, 16'd12613, 16'd57734, 16'd9913, 16'd42481, 16'd10143, 16'd5898, 16'd43253, 16'd34712, 16'd57679, 16'd18394, 16'd12344, 16'd845, 16'd7417});
	test_expansion(128'h6e510487c90b5d95a51cd0803402a2a3, {16'd48094, 16'd57289, 16'd32129, 16'd21897, 16'd33763, 16'd61488, 16'd61480, 16'd31808, 16'd43524, 16'd65062, 16'd45888, 16'd38890, 16'd11883, 16'd61789, 16'd22202, 16'd13204, 16'd22005, 16'd26243, 16'd20791, 16'd17786, 16'd18068, 16'd32949, 16'd31938, 16'd38159, 16'd29250, 16'd45207});
	test_expansion(128'h4e29542caf0fd6bc1164e2a12bb839b2, {16'd53766, 16'd11120, 16'd34850, 16'd22416, 16'd43365, 16'd63264, 16'd63979, 16'd61432, 16'd34875, 16'd58629, 16'd58770, 16'd55746, 16'd19869, 16'd51795, 16'd61128, 16'd16468, 16'd22093, 16'd5772, 16'd37577, 16'd56547, 16'd23462, 16'd60300, 16'd53730, 16'd65245, 16'd18345, 16'd48597});
	test_expansion(128'h207c803c5ecfb7f840b48c83253a032d, {16'd27713, 16'd65124, 16'd48285, 16'd52246, 16'd14387, 16'd8671, 16'd35414, 16'd57880, 16'd24170, 16'd53919, 16'd38541, 16'd58787, 16'd63866, 16'd12878, 16'd9947, 16'd50376, 16'd39866, 16'd23593, 16'd62543, 16'd53835, 16'd16625, 16'd52049, 16'd16546, 16'd25537, 16'd51507, 16'd10334});
	test_expansion(128'h7bc00dc8f3338bdae8ca82a7b933ab08, {16'd64342, 16'd35619, 16'd56271, 16'd63496, 16'd45484, 16'd3247, 16'd46552, 16'd30205, 16'd60357, 16'd46218, 16'd61659, 16'd60526, 16'd4547, 16'd42702, 16'd55755, 16'd10549, 16'd63270, 16'd57325, 16'd54708, 16'd10751, 16'd35583, 16'd2670, 16'd35581, 16'd41499, 16'd43541, 16'd47804});
	test_expansion(128'ha2f8b80ec11c1c33ece6174addd6b578, {16'd21447, 16'd5567, 16'd58692, 16'd41852, 16'd30502, 16'd50286, 16'd37528, 16'd52724, 16'd50172, 16'd1648, 16'd45322, 16'd61092, 16'd47414, 16'd6835, 16'd4438, 16'd63597, 16'd44519, 16'd27378, 16'd53634, 16'd8084, 16'd47336, 16'd13920, 16'd13404, 16'd59902, 16'd14419, 16'd56642});
	test_expansion(128'hd25debaa2e030619008c7984408a031f, {16'd48102, 16'd23908, 16'd15341, 16'd17060, 16'd52550, 16'd43036, 16'd52357, 16'd40560, 16'd9909, 16'd48465, 16'd2441, 16'd717, 16'd7406, 16'd27447, 16'd12339, 16'd46421, 16'd22617, 16'd49444, 16'd28395, 16'd65143, 16'd43653, 16'd9801, 16'd65218, 16'd48166, 16'd36486, 16'd39124});
	test_expansion(128'had96435ae7d395d7d472d8574c35775a, {16'd6870, 16'd13482, 16'd10126, 16'd42844, 16'd64502, 16'd30587, 16'd40717, 16'd17650, 16'd8827, 16'd61621, 16'd25084, 16'd4394, 16'd7165, 16'd43360, 16'd48233, 16'd51873, 16'd45565, 16'd2036, 16'd12961, 16'd46969, 16'd27191, 16'd21565, 16'd46873, 16'd29675, 16'd49831, 16'd44336});
	test_expansion(128'ha0e2143867eaf02fc264cd45c883e9aa, {16'd63462, 16'd52970, 16'd2527, 16'd59839, 16'd43721, 16'd13754, 16'd31858, 16'd29311, 16'd17505, 16'd51866, 16'd51107, 16'd4698, 16'd31672, 16'd5016, 16'd9408, 16'd37431, 16'd26222, 16'd8448, 16'd62516, 16'd48720, 16'd42249, 16'd37554, 16'd19355, 16'd10458, 16'd63545, 16'd27554});
	test_expansion(128'hf4520258e9a419158fe0a0d8f05d504b, {16'd233, 16'd51994, 16'd44645, 16'd62295, 16'd6245, 16'd15764, 16'd20172, 16'd52242, 16'd60686, 16'd33890, 16'd10975, 16'd8835, 16'd52211, 16'd43176, 16'd10725, 16'd61566, 16'd7059, 16'd59597, 16'd25, 16'd25312, 16'd31503, 16'd58799, 16'd16273, 16'd15313, 16'd17647, 16'd32088});
	test_expansion(128'h1ac4b4199154a31cad50962e0811225c, {16'd2877, 16'd3078, 16'd56135, 16'd27175, 16'd14597, 16'd10127, 16'd59143, 16'd61139, 16'd34180, 16'd33582, 16'd25013, 16'd56886, 16'd46396, 16'd40358, 16'd51395, 16'd49834, 16'd24293, 16'd63055, 16'd19730, 16'd51474, 16'd47769, 16'd50920, 16'd42927, 16'd28473, 16'd61853, 16'd34887});
	test_expansion(128'h3281f0a70681e9c1887f42d09e31e0a6, {16'd28545, 16'd29013, 16'd9431, 16'd39533, 16'd22391, 16'd19119, 16'd30378, 16'd36006, 16'd30821, 16'd26326, 16'd46514, 16'd47757, 16'd5534, 16'd57941, 16'd14982, 16'd56326, 16'd1900, 16'd52653, 16'd52769, 16'd17160, 16'd51495, 16'd35256, 16'd26569, 16'd15376, 16'd54997, 16'd49719});
	test_expansion(128'hf061ea5206b1d05cf6809ebb6f1f68c1, {16'd15018, 16'd42612, 16'd52183, 16'd37783, 16'd21640, 16'd6381, 16'd64670, 16'd9927, 16'd54144, 16'd37842, 16'd36955, 16'd41681, 16'd35957, 16'd7358, 16'd60626, 16'd21003, 16'd32379, 16'd19337, 16'd33904, 16'd43620, 16'd59802, 16'd57428, 16'd10622, 16'd60945, 16'd50535, 16'd37290});
	test_expansion(128'h83b8909b87c5c68ceb57152320edc21f, {16'd28791, 16'd32019, 16'd26778, 16'd46745, 16'd52080, 16'd16020, 16'd34997, 16'd59824, 16'd13204, 16'd52198, 16'd20940, 16'd54601, 16'd32579, 16'd6605, 16'd18502, 16'd62520, 16'd63350, 16'd23623, 16'd36233, 16'd55559, 16'd28946, 16'd50972, 16'd16595, 16'd58813, 16'd31067, 16'd45878});
	test_expansion(128'h410a9cf2f7711e78b6e58598ca6f4124, {16'd53243, 16'd64386, 16'd3932, 16'd16372, 16'd36785, 16'd42428, 16'd64753, 16'd48174, 16'd42471, 16'd41985, 16'd14491, 16'd28120, 16'd35541, 16'd16250, 16'd54385, 16'd32009, 16'd32258, 16'd39249, 16'd14681, 16'd5937, 16'd48202, 16'd41333, 16'd15052, 16'd49558, 16'd63197, 16'd2650});
	test_expansion(128'hab5618947d537cbbd65cc0739e459a55, {16'd31380, 16'd1254, 16'd40711, 16'd46107, 16'd19891, 16'd40096, 16'd13345, 16'd10179, 16'd25535, 16'd188, 16'd42028, 16'd6416, 16'd52292, 16'd9095, 16'd50841, 16'd50095, 16'd24007, 16'd1227, 16'd24428, 16'd62121, 16'd35505, 16'd18176, 16'd20372, 16'd23626, 16'd54089, 16'd2990});
	test_expansion(128'hc0fe4ac33fc4310edc4dfc4a3f3f60f4, {16'd33002, 16'd32647, 16'd63561, 16'd44064, 16'd54497, 16'd30851, 16'd19086, 16'd29825, 16'd3076, 16'd11950, 16'd18377, 16'd35334, 16'd59914, 16'd62603, 16'd35669, 16'd22507, 16'd32280, 16'd43874, 16'd11903, 16'd35744, 16'd59470, 16'd14642, 16'd62762, 16'd39447, 16'd63412, 16'd7106});
	test_expansion(128'hb7dc25cedb90ec10555662817e1279ec, {16'd36697, 16'd29292, 16'd10210, 16'd61859, 16'd49886, 16'd47202, 16'd42815, 16'd39668, 16'd18822, 16'd21227, 16'd44505, 16'd55444, 16'd21917, 16'd15332, 16'd9868, 16'd38205, 16'd21765, 16'd50991, 16'd3913, 16'd46608, 16'd7130, 16'd18144, 16'd62204, 16'd47798, 16'd52757, 16'd1834});
	test_expansion(128'hdc73cd2d0e4fecfef6f953bb5d9966e6, {16'd50952, 16'd58591, 16'd18544, 16'd34524, 16'd29118, 16'd14253, 16'd5295, 16'd56759, 16'd14085, 16'd30117, 16'd1471, 16'd64570, 16'd24617, 16'd37265, 16'd8520, 16'd21556, 16'd52472, 16'd33354, 16'd7012, 16'd22968, 16'd54396, 16'd6640, 16'd18087, 16'd57721, 16'd46622, 16'd47209});
	test_expansion(128'ha0cdcca6fbf063a4b772e3055017934d, {16'd65111, 16'd14172, 16'd41225, 16'd36167, 16'd27665, 16'd10809, 16'd33925, 16'd13696, 16'd13669, 16'd1041, 16'd65127, 16'd64627, 16'd48287, 16'd19545, 16'd51693, 16'd16607, 16'd47654, 16'd18862, 16'd36689, 16'd36238, 16'd13249, 16'd39391, 16'd54097, 16'd18566, 16'd26767, 16'd26188});
	test_expansion(128'hee5e1073a9dae493ac1a75a3437897d7, {16'd24684, 16'd52569, 16'd36353, 16'd11314, 16'd22265, 16'd57016, 16'd38811, 16'd1021, 16'd58672, 16'd15507, 16'd24967, 16'd33347, 16'd23987, 16'd33636, 16'd13144, 16'd21517, 16'd24969, 16'd52589, 16'd12355, 16'd52889, 16'd55627, 16'd56671, 16'd40115, 16'd54868, 16'd24498, 16'd25044});
	test_expansion(128'h91484bd6843605f58232524cb55f9d63, {16'd15836, 16'd46671, 16'd43601, 16'd25781, 16'd8921, 16'd56372, 16'd53905, 16'd40590, 16'd41948, 16'd20607, 16'd16216, 16'd2852, 16'd42293, 16'd60433, 16'd18500, 16'd55491, 16'd42758, 16'd57543, 16'd10707, 16'd36902, 16'd42550, 16'd12196, 16'd38105, 16'd26109, 16'd30346, 16'd61632});
	test_expansion(128'h0c0c975faa665c7533f807191329e488, {16'd55737, 16'd18473, 16'd55456, 16'd11255, 16'd53956, 16'd1871, 16'd14893, 16'd51537, 16'd12800, 16'd30161, 16'd25203, 16'd51139, 16'd33330, 16'd11776, 16'd50414, 16'd50332, 16'd57766, 16'd31498, 16'd20781, 16'd53183, 16'd50397, 16'd45338, 16'd13653, 16'd24976, 16'd32878, 16'd41997});
	test_expansion(128'h8bb2f9ee306d8b039c1ed56b81109caa, {16'd48300, 16'd16036, 16'd63344, 16'd26664, 16'd40246, 16'd55318, 16'd45141, 16'd33718, 16'd62499, 16'd8381, 16'd8024, 16'd36888, 16'd63843, 16'd12613, 16'd39995, 16'd14453, 16'd37316, 16'd39922, 16'd38716, 16'd62531, 16'd46138, 16'd33667, 16'd50079, 16'd54070, 16'd36171, 16'd40108});
	test_expansion(128'h436ebf9b0cdc04b7ecc735c893b62ef7, {16'd29406, 16'd30439, 16'd3652, 16'd7658, 16'd39693, 16'd23989, 16'd51393, 16'd51950, 16'd40349, 16'd63534, 16'd44939, 16'd52626, 16'd4566, 16'd30175, 16'd21041, 16'd62130, 16'd54361, 16'd3555, 16'd5985, 16'd37322, 16'd22798, 16'd22605, 16'd43342, 16'd16874, 16'd3643, 16'd40729});
	test_expansion(128'hf7f75e824883c262e3a0749b15b403b5, {16'd21807, 16'd10832, 16'd39681, 16'd63752, 16'd35052, 16'd12616, 16'd3396, 16'd58313, 16'd54886, 16'd65348, 16'd12457, 16'd62015, 16'd14030, 16'd19142, 16'd17244, 16'd13284, 16'd5474, 16'd51400, 16'd65456, 16'd54493, 16'd2446, 16'd40596, 16'd24009, 16'd53734, 16'd38085, 16'd41957});
	test_expansion(128'he4c306066ff299b327f3cca73a1697aa, {16'd34729, 16'd62612, 16'd53201, 16'd50724, 16'd42352, 16'd17305, 16'd56929, 16'd58515, 16'd19906, 16'd27840, 16'd37210, 16'd14438, 16'd53326, 16'd17965, 16'd42538, 16'd23288, 16'd49240, 16'd30662, 16'd32913, 16'd2423, 16'd46692, 16'd37837, 16'd17996, 16'd11735, 16'd13238, 16'd56299});
	test_expansion(128'h54d9db84ba3f1dfe54ffec1d62ee20b1, {16'd37985, 16'd12026, 16'd52978, 16'd11677, 16'd24561, 16'd21037, 16'd38824, 16'd28329, 16'd4795, 16'd60263, 16'd41048, 16'd27973, 16'd64800, 16'd61117, 16'd27151, 16'd22706, 16'd48018, 16'd5414, 16'd42824, 16'd19471, 16'd22487, 16'd18160, 16'd60230, 16'd1204, 16'd41581, 16'd14984});
	test_expansion(128'he98d9c05b5565a16103ecd87b6b1912d, {16'd14152, 16'd3172, 16'd2067, 16'd38765, 16'd64457, 16'd18951, 16'd10036, 16'd44659, 16'd52952, 16'd20078, 16'd35669, 16'd7979, 16'd57575, 16'd28134, 16'd2941, 16'd59922, 16'd61177, 16'd30554, 16'd33135, 16'd52993, 16'd61467, 16'd15167, 16'd45384, 16'd23296, 16'd45406, 16'd54954});
	test_expansion(128'h224cf43aead75d1fff0b3b09eb376c3e, {16'd12007, 16'd23561, 16'd30247, 16'd57602, 16'd20198, 16'd25026, 16'd49770, 16'd46951, 16'd25228, 16'd42283, 16'd40050, 16'd19281, 16'd20130, 16'd4916, 16'd39466, 16'd51653, 16'd8286, 16'd27710, 16'd29328, 16'd47052, 16'd38325, 16'd59116, 16'd48098, 16'd49857, 16'd52738, 16'd5590});
	test_expansion(128'h648412a2a07cea68f6e52786950df822, {16'd58301, 16'd48860, 16'd24513, 16'd36638, 16'd1849, 16'd17257, 16'd41838, 16'd4003, 16'd39769, 16'd56274, 16'd47399, 16'd8285, 16'd43147, 16'd52557, 16'd19841, 16'd43158, 16'd19254, 16'd21896, 16'd9572, 16'd17803, 16'd7882, 16'd37339, 16'd57910, 16'd22459, 16'd11403, 16'd31354});
	test_expansion(128'hffe6f0af2a355e1c40057758d758b973, {16'd39326, 16'd31299, 16'd9354, 16'd60848, 16'd8872, 16'd41357, 16'd38632, 16'd8024, 16'd39293, 16'd25643, 16'd17228, 16'd17931, 16'd33284, 16'd1516, 16'd55986, 16'd47536, 16'd45850, 16'd34183, 16'd847, 16'd64322, 16'd51310, 16'd49343, 16'd38471, 16'd26701, 16'd55534, 16'd17185});
	test_expansion(128'hb0f25699d78a1937ed61abb42bf21544, {16'd45931, 16'd62798, 16'd19892, 16'd19487, 16'd15322, 16'd41270, 16'd42619, 16'd5910, 16'd35131, 16'd40220, 16'd13173, 16'd38337, 16'd21488, 16'd37859, 16'd35699, 16'd49890, 16'd54976, 16'd23748, 16'd12502, 16'd2608, 16'd28257, 16'd14031, 16'd14659, 16'd22185, 16'd16309, 16'd15540});
	test_expansion(128'h52dc8b03f4db8d1a3c2592e9a85052a4, {16'd13794, 16'd50085, 16'd21015, 16'd57046, 16'd32842, 16'd17360, 16'd2191, 16'd2321, 16'd4456, 16'd4203, 16'd55931, 16'd6140, 16'd12599, 16'd37089, 16'd21809, 16'd33694, 16'd51909, 16'd646, 16'd18217, 16'd63126, 16'd31644, 16'd26562, 16'd37728, 16'd53199, 16'd3564, 16'd64602});
	test_expansion(128'h7c477169fc5115f6f2806834f10e77cd, {16'd27176, 16'd52177, 16'd27368, 16'd32105, 16'd37750, 16'd22931, 16'd44312, 16'd45708, 16'd57742, 16'd49273, 16'd63581, 16'd45788, 16'd3136, 16'd43302, 16'd3461, 16'd51372, 16'd63977, 16'd1386, 16'd8084, 16'd57248, 16'd27684, 16'd14003, 16'd46850, 16'd47955, 16'd22430, 16'd62304});
	test_expansion(128'h866aeb4094b3ed2349ec406c4d2da593, {16'd55356, 16'd5006, 16'd24250, 16'd36236, 16'd61420, 16'd10702, 16'd51855, 16'd8587, 16'd22809, 16'd59555, 16'd20474, 16'd52427, 16'd16446, 16'd47027, 16'd39589, 16'd30971, 16'd65200, 16'd19178, 16'd4853, 16'd2619, 16'd62323, 16'd30434, 16'd21973, 16'd53167, 16'd56283, 16'd32468});
	test_expansion(128'h3ac5009ee3717f35323d0670f801953b, {16'd38966, 16'd12579, 16'd53965, 16'd65308, 16'd2877, 16'd58796, 16'd20680, 16'd17354, 16'd52731, 16'd40623, 16'd54533, 16'd45763, 16'd62386, 16'd54932, 16'd45921, 16'd23256, 16'd7995, 16'd48287, 16'd9795, 16'd28632, 16'd19917, 16'd54710, 16'd51691, 16'd3962, 16'd39511, 16'd43147});
	test_expansion(128'h44c2392ab7bd812e176b6ba9449b8c8c, {16'd59959, 16'd55224, 16'd7399, 16'd41353, 16'd48142, 16'd62814, 16'd15520, 16'd43193, 16'd53403, 16'd2789, 16'd6845, 16'd51654, 16'd44452, 16'd17026, 16'd20842, 16'd22838, 16'd19737, 16'd7769, 16'd12398, 16'd24369, 16'd3645, 16'd5742, 16'd25848, 16'd39736, 16'd29527, 16'd33454});
	test_expansion(128'hb7cbfe76b7af4acc3a8e7329d06c1066, {16'd24271, 16'd22443, 16'd54718, 16'd8227, 16'd30182, 16'd49516, 16'd45233, 16'd26770, 16'd30485, 16'd29171, 16'd12473, 16'd38698, 16'd20385, 16'd30195, 16'd49526, 16'd23317, 16'd61268, 16'd23944, 16'd57499, 16'd8698, 16'd50316, 16'd35496, 16'd35526, 16'd43819, 16'd21784, 16'd14229});
	test_expansion(128'hb89ed3ee881c1bc9dbd4233da915125e, {16'd52532, 16'd9043, 16'd49427, 16'd40109, 16'd43649, 16'd7307, 16'd12262, 16'd40325, 16'd35823, 16'd22753, 16'd58784, 16'd27305, 16'd39657, 16'd51876, 16'd42813, 16'd58122, 16'd52756, 16'd22775, 16'd20352, 16'd63392, 16'd13213, 16'd18585, 16'd21536, 16'd49615, 16'd14342, 16'd48103});
	test_expansion(128'h54c34f64efa653a3ad1d96eaf2e5e38f, {16'd35944, 16'd11948, 16'd49574, 16'd26310, 16'd59320, 16'd34727, 16'd58772, 16'd38724, 16'd34053, 16'd9490, 16'd14985, 16'd43312, 16'd44408, 16'd21443, 16'd4974, 16'd6441, 16'd32113, 16'd10776, 16'd13155, 16'd31650, 16'd13988, 16'd43527, 16'd65226, 16'd46145, 16'd5271, 16'd46914});
	test_expansion(128'ha14bd9571b0ad758305ec14823ae3aeb, {16'd56975, 16'd25246, 16'd30379, 16'd56277, 16'd23914, 16'd1789, 16'd29398, 16'd56795, 16'd40669, 16'd46536, 16'd41488, 16'd64765, 16'd20431, 16'd25311, 16'd44585, 16'd1494, 16'd1664, 16'd2690, 16'd7863, 16'd3011, 16'd59714, 16'd45769, 16'd53844, 16'd15597, 16'd53241, 16'd39420});
	test_expansion(128'h1f22e2e9e5a591c0e794a951413e21e1, {16'd34359, 16'd35339, 16'd5068, 16'd55812, 16'd27801, 16'd53830, 16'd11406, 16'd15424, 16'd54942, 16'd3838, 16'd35123, 16'd11396, 16'd39979, 16'd51572, 16'd38045, 16'd26850, 16'd54877, 16'd25252, 16'd34602, 16'd34638, 16'd46688, 16'd57425, 16'd55736, 16'd4263, 16'd58575, 16'd35836});
	test_expansion(128'h20ea84901e6eedc3e8a5e79a2cd073f9, {16'd56309, 16'd47791, 16'd6452, 16'd60181, 16'd14407, 16'd15385, 16'd45809, 16'd53007, 16'd37719, 16'd28281, 16'd46178, 16'd36356, 16'd26570, 16'd3886, 16'd49649, 16'd16992, 16'd19188, 16'd14786, 16'd44230, 16'd18085, 16'd62586, 16'd12163, 16'd9629, 16'd40943, 16'd52990, 16'd54196});
	test_expansion(128'h85c09c6c40fe491c660cf8627972759e, {16'd6914, 16'd21856, 16'd7980, 16'd20882, 16'd32695, 16'd62258, 16'd3388, 16'd959, 16'd58934, 16'd23479, 16'd55942, 16'd27319, 16'd13714, 16'd741, 16'd6980, 16'd62313, 16'd8340, 16'd26712, 16'd25812, 16'd35205, 16'd32957, 16'd26181, 16'd12857, 16'd7327, 16'd32890, 16'd55695});
	test_expansion(128'hfc939a9d13e0f0e726963e6a305bbcd6, {16'd55219, 16'd8151, 16'd37310, 16'd1725, 16'd29228, 16'd23099, 16'd56283, 16'd22137, 16'd45334, 16'd23270, 16'd65413, 16'd46376, 16'd45985, 16'd64263, 16'd16315, 16'd15700, 16'd6029, 16'd57509, 16'd19146, 16'd22363, 16'd16084, 16'd35997, 16'd47955, 16'd16501, 16'd27066, 16'd56446});
	test_expansion(128'h5c62bbb418681c463e0203b31c66ce4e, {16'd13199, 16'd64786, 16'd35676, 16'd10909, 16'd12491, 16'd42290, 16'd42151, 16'd57032, 16'd36768, 16'd3501, 16'd62930, 16'd49939, 16'd26602, 16'd2571, 16'd35759, 16'd37089, 16'd41608, 16'd40820, 16'd51938, 16'd1176, 16'd27093, 16'd60147, 16'd53046, 16'd40728, 16'd10952, 16'd5391});
	test_expansion(128'h2c2b0d0030c455f4ed0fa1806464f6b5, {16'd27370, 16'd30708, 16'd18177, 16'd19884, 16'd55932, 16'd61058, 16'd4480, 16'd27096, 16'd49643, 16'd21208, 16'd21383, 16'd5163, 16'd64536, 16'd27189, 16'd16661, 16'd56380, 16'd53070, 16'd42464, 16'd16193, 16'd6820, 16'd9629, 16'd28293, 16'd44399, 16'd25986, 16'd61221, 16'd19671});
	test_expansion(128'hc77d9f8dcb7b3fc4959be818f92e783d, {16'd1217, 16'd50793, 16'd58595, 16'd26300, 16'd37723, 16'd26465, 16'd8574, 16'd31044, 16'd64423, 16'd48491, 16'd20118, 16'd33729, 16'd43025, 16'd45928, 16'd53778, 16'd41059, 16'd34419, 16'd17726, 16'd57638, 16'd47206, 16'd18061, 16'd61269, 16'd45503, 16'd55883, 16'd16140, 16'd10665});
	test_expansion(128'h33bf1408896749054e8c9406c2d85ae7, {16'd20976, 16'd44440, 16'd41696, 16'd32919, 16'd32745, 16'd53309, 16'd20238, 16'd18298, 16'd41859, 16'd13833, 16'd57224, 16'd8882, 16'd6526, 16'd48441, 16'd18609, 16'd23921, 16'd49826, 16'd15450, 16'd9782, 16'd13574, 16'd36566, 16'd38666, 16'd48562, 16'd16461, 16'd31153, 16'd7705});
	test_expansion(128'h5e6fe6c306e5218b47f4bb6d02468762, {16'd7371, 16'd42399, 16'd53868, 16'd34074, 16'd27041, 16'd32171, 16'd40767, 16'd21297, 16'd4398, 16'd10561, 16'd8345, 16'd42654, 16'd52636, 16'd45973, 16'd65142, 16'd11068, 16'd45853, 16'd15719, 16'd16201, 16'd64774, 16'd5901, 16'd47316, 16'd56927, 16'd29667, 16'd533, 16'd19827});
	test_expansion(128'h9ca9f859a663e4abfbe88a352323a7f1, {16'd15922, 16'd5376, 16'd155, 16'd31262, 16'd50895, 16'd24748, 16'd7897, 16'd61917, 16'd20448, 16'd16992, 16'd901, 16'd55552, 16'd24, 16'd58085, 16'd35220, 16'd27565, 16'd22998, 16'd57912, 16'd9090, 16'd56552, 16'd3073, 16'd4135, 16'd2205, 16'd63712, 16'd47039, 16'd35111});
	test_expansion(128'h464664d2daad939c50c30fd867197832, {16'd16750, 16'd52888, 16'd9046, 16'd49917, 16'd52077, 16'd32800, 16'd3254, 16'd41841, 16'd31731, 16'd56020, 16'd13172, 16'd1787, 16'd16085, 16'd50948, 16'd43306, 16'd65356, 16'd61326, 16'd37675, 16'd40797, 16'd9487, 16'd41537, 16'd18334, 16'd46183, 16'd10628, 16'd4795, 16'd24214});
	test_expansion(128'h13e6f76978e7efefb0b3e6c84b5279e3, {16'd13787, 16'd43252, 16'd64885, 16'd65451, 16'd62436, 16'd11020, 16'd35901, 16'd27212, 16'd34780, 16'd25217, 16'd18574, 16'd33451, 16'd41379, 16'd26619, 16'd6134, 16'd65085, 16'd58418, 16'd46603, 16'd64580, 16'd10482, 16'd54980, 16'd14772, 16'd18329, 16'd25573, 16'd63767, 16'd48119});
	test_expansion(128'hb2f44a941e0a8cb7a9da3b1a50965fae, {16'd47479, 16'd34519, 16'd5583, 16'd25781, 16'd22979, 16'd57638, 16'd47229, 16'd51115, 16'd53929, 16'd8670, 16'd52244, 16'd3805, 16'd60340, 16'd57657, 16'd3382, 16'd34842, 16'd56465, 16'd30691, 16'd16270, 16'd14806, 16'd27878, 16'd59284, 16'd20998, 16'd34161, 16'd34588, 16'd19455});
	test_expansion(128'h80cf5ffc0d9dfa8e2cb6eb59df3d4ff4, {16'd4219, 16'd16398, 16'd41409, 16'd43758, 16'd7476, 16'd33700, 16'd29809, 16'd52343, 16'd6527, 16'd45057, 16'd61928, 16'd45428, 16'd58901, 16'd26935, 16'd60839, 16'd5230, 16'd61759, 16'd27798, 16'd60846, 16'd38998, 16'd47852, 16'd25368, 16'd53108, 16'd45964, 16'd11915, 16'd32666});
	test_expansion(128'h697e57da518c98e3fe4607dfe7122a6d, {16'd4192, 16'd3407, 16'd51875, 16'd4060, 16'd58879, 16'd14782, 16'd33636, 16'd20863, 16'd6403, 16'd34409, 16'd11134, 16'd52651, 16'd50007, 16'd18850, 16'd21099, 16'd24355, 16'd23687, 16'd23751, 16'd22095, 16'd18071, 16'd12392, 16'd52347, 16'd40986, 16'd19709, 16'd56254, 16'd30891});
	test_expansion(128'h4f438b7300c9d76188a7994bcc3b683f, {16'd4343, 16'd21466, 16'd9373, 16'd57118, 16'd6576, 16'd55343, 16'd62391, 16'd47057, 16'd27730, 16'd37322, 16'd41609, 16'd58228, 16'd16115, 16'd2579, 16'd42043, 16'd64747, 16'd25170, 16'd60216, 16'd59869, 16'd27915, 16'd28688, 16'd16792, 16'd1208, 16'd27409, 16'd43447, 16'd1232});
	test_expansion(128'hfe8e135e46c45334ebd08d532ee80e0c, {16'd6333, 16'd49949, 16'd23598, 16'd12793, 16'd31952, 16'd629, 16'd42165, 16'd45058, 16'd24290, 16'd51507, 16'd1052, 16'd18621, 16'd16763, 16'd49063, 16'd8727, 16'd62617, 16'd58090, 16'd12511, 16'd57668, 16'd33809, 16'd61617, 16'd6617, 16'd23852, 16'd4677, 16'd59843, 16'd33348});
	test_expansion(128'he26ff863b40c213f21056340edc53ebd, {16'd1045, 16'd60631, 16'd8739, 16'd55708, 16'd65058, 16'd27407, 16'd47484, 16'd15884, 16'd35640, 16'd62640, 16'd47951, 16'd19201, 16'd11803, 16'd54012, 16'd17654, 16'd54333, 16'd13362, 16'd35537, 16'd35103, 16'd9372, 16'd5375, 16'd1382, 16'd21137, 16'd21864, 16'd18629, 16'd23088});
	test_expansion(128'h891ae79871e9bee0833201227745a21c, {16'd20906, 16'd43339, 16'd48591, 16'd50874, 16'd48657, 16'd16991, 16'd32464, 16'd4470, 16'd50327, 16'd24220, 16'd38621, 16'd26170, 16'd33816, 16'd20294, 16'd11593, 16'd47767, 16'd6934, 16'd41480, 16'd17134, 16'd9367, 16'd54320, 16'd62951, 16'd16382, 16'd6191, 16'd9460, 16'd50232});
	test_expansion(128'h2ab711f3d0bc60eb04d54c3daddb7e18, {16'd20084, 16'd39671, 16'd45669, 16'd62116, 16'd32248, 16'd65329, 16'd16716, 16'd9735, 16'd49064, 16'd5180, 16'd28025, 16'd1530, 16'd2179, 16'd9392, 16'd23362, 16'd311, 16'd7563, 16'd7049, 16'd44114, 16'd5908, 16'd29703, 16'd38171, 16'd51559, 16'd46464, 16'd58431, 16'd11398});
	test_expansion(128'h98a8b209e3310dab025c197d14c3a921, {16'd12368, 16'd33801, 16'd44076, 16'd47202, 16'd59223, 16'd13306, 16'd5775, 16'd20982, 16'd62668, 16'd11352, 16'd54808, 16'd35570, 16'd32387, 16'd11046, 16'd63196, 16'd10416, 16'd62806, 16'd30395, 16'd62128, 16'd36581, 16'd31984, 16'd14620, 16'd43135, 16'd28677, 16'd56309, 16'd51815});
	test_expansion(128'hbfbf4e8a3b7531cd4900c19437d8c7a3, {16'd46318, 16'd15749, 16'd43584, 16'd44929, 16'd62635, 16'd10034, 16'd604, 16'd1628, 16'd37295, 16'd29442, 16'd54883, 16'd13698, 16'd45032, 16'd53703, 16'd6125, 16'd64175, 16'd57345, 16'd48411, 16'd26490, 16'd4788, 16'd62623, 16'd19307, 16'd27480, 16'd5528, 16'd46993, 16'd51891});
	test_expansion(128'h18c243d1ef2bbc7e6ef6e2f4b36626fe, {16'd55100, 16'd1492, 16'd38405, 16'd63274, 16'd44877, 16'd31570, 16'd27902, 16'd47753, 16'd60884, 16'd53862, 16'd60993, 16'd4912, 16'd60028, 16'd26004, 16'd52107, 16'd32072, 16'd51928, 16'd38374, 16'd29483, 16'd60011, 16'd25070, 16'd12554, 16'd45635, 16'd36691, 16'd41853, 16'd5474});
	test_expansion(128'hd12ef909148d7e227062ab3a15e55ef2, {16'd17097, 16'd59347, 16'd10728, 16'd35976, 16'd46372, 16'd23339, 16'd11669, 16'd47998, 16'd19472, 16'd55260, 16'd61284, 16'd8185, 16'd38298, 16'd43903, 16'd63789, 16'd36306, 16'd20553, 16'd56827, 16'd8155, 16'd43123, 16'd17313, 16'd1744, 16'd36453, 16'd58854, 16'd23316, 16'd63071});
	test_expansion(128'h87e1cd664cfac2cd45b0583974ed0393, {16'd8814, 16'd6080, 16'd35668, 16'd1673, 16'd26894, 16'd36517, 16'd3137, 16'd11293, 16'd18732, 16'd20614, 16'd8353, 16'd4069, 16'd58297, 16'd40165, 16'd82, 16'd45509, 16'd13277, 16'd29859, 16'd37379, 16'd13104, 16'd52793, 16'd24752, 16'd2163, 16'd14951, 16'd63889, 16'd13964});
	test_expansion(128'hfe2b80b0ba16cecdd0cd3fb8f18598c9, {16'd31282, 16'd33946, 16'd17063, 16'd16000, 16'd2144, 16'd61146, 16'd65526, 16'd57409, 16'd56053, 16'd56333, 16'd35877, 16'd27952, 16'd27767, 16'd55874, 16'd17754, 16'd302, 16'd11024, 16'd31757, 16'd19780, 16'd33104, 16'd9771, 16'd32251, 16'd33688, 16'd1257, 16'd4935, 16'd22822});
	test_expansion(128'h23c262421b4555d2f84383f894b2f01c, {16'd39874, 16'd28498, 16'd35663, 16'd23168, 16'd22039, 16'd45626, 16'd22831, 16'd64507, 16'd1424, 16'd24891, 16'd1253, 16'd53088, 16'd16100, 16'd24444, 16'd36694, 16'd13102, 16'd53980, 16'd32475, 16'd46604, 16'd8615, 16'd18094, 16'd27170, 16'd59930, 16'd49721, 16'd55768, 16'd52627});
	test_expansion(128'h177870203a09212d5ef7808b67e91964, {16'd34162, 16'd50559, 16'd54151, 16'd59689, 16'd43698, 16'd12047, 16'd22094, 16'd27452, 16'd45424, 16'd44484, 16'd19465, 16'd47047, 16'd25284, 16'd51755, 16'd59832, 16'd25475, 16'd63909, 16'd43133, 16'd19059, 16'd19226, 16'd31055, 16'd38560, 16'd46257, 16'd51843, 16'd28521, 16'd14825});
	test_expansion(128'hb3922465b5fd5bee4a5a71dfc8fcf4ec, {16'd37595, 16'd14031, 16'd60018, 16'd18990, 16'd41928, 16'd13113, 16'd56595, 16'd47075, 16'd36845, 16'd17603, 16'd61204, 16'd16359, 16'd32847, 16'd51761, 16'd52498, 16'd25197, 16'd45957, 16'd5864, 16'd64756, 16'd8302, 16'd43376, 16'd44603, 16'd10768, 16'd56814, 16'd61545, 16'd13298});
	test_expansion(128'h883a4f8f59829afee542d08ba57c7272, {16'd54995, 16'd22758, 16'd63460, 16'd7177, 16'd36167, 16'd11940, 16'd49569, 16'd38640, 16'd19484, 16'd5644, 16'd13142, 16'd40901, 16'd7153, 16'd38812, 16'd2838, 16'd46413, 16'd34182, 16'd34612, 16'd19602, 16'd61567, 16'd27674, 16'd25959, 16'd47979, 16'd47837, 16'd29633, 16'd44948});
	test_expansion(128'h396616d9d54a2139e55e156c45b2303e, {16'd4102, 16'd52767, 16'd4566, 16'd18746, 16'd39747, 16'd500, 16'd2367, 16'd42042, 16'd62796, 16'd56736, 16'd58896, 16'd62792, 16'd55838, 16'd20099, 16'd27455, 16'd48736, 16'd24234, 16'd14571, 16'd48189, 16'd60242, 16'd11276, 16'd15434, 16'd37032, 16'd41417, 16'd58597, 16'd9816});
	test_expansion(128'haf5b2128729322f1dd05d4c5fd6fb731, {16'd52125, 16'd60202, 16'd22049, 16'd9798, 16'd1035, 16'd34544, 16'd15987, 16'd44817, 16'd59754, 16'd20145, 16'd37710, 16'd40022, 16'd42879, 16'd59763, 16'd55771, 16'd11997, 16'd53403, 16'd41732, 16'd3237, 16'd30903, 16'd33437, 16'd4091, 16'd42305, 16'd35528, 16'd27508, 16'd64952});
	test_expansion(128'he1adc5ea02e55cebc5e2e08edde9e00f, {16'd41474, 16'd785, 16'd28781, 16'd35704, 16'd37554, 16'd7175, 16'd48295, 16'd65244, 16'd6065, 16'd13175, 16'd23532, 16'd15431, 16'd11861, 16'd26378, 16'd22693, 16'd64895, 16'd51003, 16'd40728, 16'd62590, 16'd1915, 16'd61708, 16'd51840, 16'd19896, 16'd56361, 16'd38631, 16'd24903});
	test_expansion(128'h334c953e0ad1f996df419b419092af8e, {16'd20994, 16'd14391, 16'd43679, 16'd23541, 16'd14379, 16'd46069, 16'd43144, 16'd60685, 16'd34563, 16'd59193, 16'd18092, 16'd60968, 16'd62487, 16'd10067, 16'd32241, 16'd16227, 16'd64159, 16'd36993, 16'd22041, 16'd51462, 16'd57315, 16'd20122, 16'd45756, 16'd53225, 16'd50114, 16'd55482});
	test_expansion(128'h5753fdbb6743e0f92d95218eb6991c90, {16'd61751, 16'd60162, 16'd22948, 16'd55507, 16'd63109, 16'd52983, 16'd43916, 16'd52304, 16'd30964, 16'd11814, 16'd58151, 16'd33018, 16'd54850, 16'd43885, 16'd48783, 16'd18546, 16'd30969, 16'd23541, 16'd19291, 16'd4478, 16'd43719, 16'd47651, 16'd2488, 16'd29286, 16'd46172, 16'd56596});
	test_expansion(128'h6a893544aa0ae304be4be68259015ae5, {16'd51678, 16'd59020, 16'd5087, 16'd11620, 16'd52397, 16'd30184, 16'd48568, 16'd14852, 16'd20266, 16'd30933, 16'd32578, 16'd14074, 16'd39941, 16'd51194, 16'd45992, 16'd61445, 16'd13235, 16'd51071, 16'd41325, 16'd13900, 16'd61943, 16'd48643, 16'd36795, 16'd65450, 16'd37557, 16'd36063});
	test_expansion(128'h62fcfc3bff5fe1e85885bed209ff0f17, {16'd47458, 16'd21633, 16'd12143, 16'd32572, 16'd50952, 16'd46842, 16'd3201, 16'd18976, 16'd49381, 16'd11172, 16'd32407, 16'd62803, 16'd43609, 16'd6068, 16'd52014, 16'd11864, 16'd30146, 16'd44663, 16'd6155, 16'd21301, 16'd64695, 16'd23375, 16'd62102, 16'd5357, 16'd54971, 16'd2294});
	test_expansion(128'h9b6a4c6858ced78c86a430b0f341409d, {16'd316, 16'd60540, 16'd30640, 16'd26160, 16'd23094, 16'd11312, 16'd28903, 16'd13343, 16'd61002, 16'd55069, 16'd31634, 16'd14558, 16'd35350, 16'd59424, 16'd62513, 16'd11576, 16'd18959, 16'd37232, 16'd38603, 16'd6680, 16'd38820, 16'd40479, 16'd29742, 16'd42718, 16'd10342, 16'd26416});
	test_expansion(128'hd30b9728ecaa3a2cd06cccc6fefcd454, {16'd34513, 16'd64880, 16'd18623, 16'd60090, 16'd19740, 16'd55029, 16'd45226, 16'd57433, 16'd39334, 16'd47499, 16'd43061, 16'd50932, 16'd38940, 16'd545, 16'd26337, 16'd55886, 16'd10058, 16'd16062, 16'd45064, 16'd866, 16'd3081, 16'd38972, 16'd57172, 16'd22380, 16'd8839, 16'd11951});
	test_expansion(128'h458c84855cd78bcf62748a7db13db7e0, {16'd63524, 16'd33423, 16'd38746, 16'd55836, 16'd63020, 16'd25100, 16'd40286, 16'd42811, 16'd21461, 16'd41061, 16'd62114, 16'd57464, 16'd32201, 16'd9150, 16'd58920, 16'd9654, 16'd31909, 16'd58328, 16'd1553, 16'd18137, 16'd25226, 16'd48262, 16'd62154, 16'd16755, 16'd46954, 16'd34240});
	test_expansion(128'h35d3212d9bc36e930adb941734ef331c, {16'd36587, 16'd49208, 16'd31565, 16'd54021, 16'd62567, 16'd11477, 16'd59747, 16'd11160, 16'd15389, 16'd21410, 16'd38669, 16'd53684, 16'd48372, 16'd40130, 16'd63411, 16'd32034, 16'd20883, 16'd23221, 16'd23904, 16'd7652, 16'd6141, 16'd33155, 16'd29413, 16'd22437, 16'd10622, 16'd56465});
	test_expansion(128'he0a8e2042f587388cd670ce59944798d, {16'd8411, 16'd46972, 16'd32925, 16'd27013, 16'd62162, 16'd36951, 16'd35895, 16'd25492, 16'd44923, 16'd40030, 16'd30744, 16'd25140, 16'd58428, 16'd57772, 16'd49341, 16'd8368, 16'd6934, 16'd48543, 16'd13984, 16'd48724, 16'd58966, 16'd20586, 16'd41931, 16'd15051, 16'd23616, 16'd18994});
	test_expansion(128'h282cbe314c0af306fcba8e676a327e51, {16'd19532, 16'd37989, 16'd36196, 16'd31257, 16'd47509, 16'd22762, 16'd2557, 16'd56808, 16'd29000, 16'd64653, 16'd37057, 16'd33060, 16'd49682, 16'd25853, 16'd43826, 16'd33039, 16'd29864, 16'd57311, 16'd14347, 16'd34738, 16'd45000, 16'd47835, 16'd25760, 16'd5752, 16'd18860, 16'd59291});
	test_expansion(128'h8b0482681bbd111b4911986e3a9ec138, {16'd54471, 16'd25757, 16'd6418, 16'd10425, 16'd56846, 16'd27567, 16'd36815, 16'd39187, 16'd59122, 16'd15116, 16'd52568, 16'd37011, 16'd40832, 16'd56603, 16'd55879, 16'd46999, 16'd35916, 16'd50645, 16'd2965, 16'd16580, 16'd213, 16'd43256, 16'd30705, 16'd42116, 16'd13889, 16'd16357});
	test_expansion(128'hb6bf4941414554be6bb737b6ab997ad6, {16'd12688, 16'd7115, 16'd48888, 16'd61307, 16'd42786, 16'd64070, 16'd12759, 16'd52021, 16'd10835, 16'd32666, 16'd24957, 16'd57234, 16'd26768, 16'd55265, 16'd30862, 16'd41132, 16'd57953, 16'd4020, 16'd36830, 16'd20535, 16'd52322, 16'd36636, 16'd47007, 16'd63108, 16'd53133, 16'd32392});
	test_expansion(128'h63d592497786cdde6c7da3608a20156a, {16'd23367, 16'd62825, 16'd12243, 16'd64856, 16'd22556, 16'd57194, 16'd2389, 16'd2350, 16'd47716, 16'd29187, 16'd6290, 16'd62036, 16'd56194, 16'd17610, 16'd58025, 16'd15135, 16'd8848, 16'd2390, 16'd35377, 16'd53891, 16'd57550, 16'd34356, 16'd40084, 16'd55376, 16'd5800, 16'd33609});
	test_expansion(128'h6471316cd7985ad7a1e5e564094a6f7f, {16'd4535, 16'd21902, 16'd28312, 16'd10714, 16'd34136, 16'd42377, 16'd16125, 16'd30788, 16'd64961, 16'd37820, 16'd22934, 16'd61330, 16'd36464, 16'd10092, 16'd51893, 16'd10309, 16'd11929, 16'd29852, 16'd44373, 16'd34360, 16'd36659, 16'd26491, 16'd162, 16'd12835, 16'd54272, 16'd25889});
	test_expansion(128'h66ca558c8b7d0ecbc23145603d2c83c0, {16'd31803, 16'd40615, 16'd15474, 16'd8631, 16'd28394, 16'd33599, 16'd52539, 16'd48332, 16'd32831, 16'd22167, 16'd52820, 16'd46864, 16'd50649, 16'd26662, 16'd16220, 16'd6456, 16'd6298, 16'd15301, 16'd61447, 16'd52495, 16'd28149, 16'd49320, 16'd61365, 16'd8374, 16'd1582, 16'd12805});
	test_expansion(128'hde1e4017edf9f722e066dddd3d543ece, {16'd11582, 16'd55018, 16'd23928, 16'd22722, 16'd44161, 16'd17367, 16'd57079, 16'd38106, 16'd18954, 16'd16826, 16'd1986, 16'd48331, 16'd45488, 16'd33685, 16'd10872, 16'd35342, 16'd25351, 16'd29885, 16'd64685, 16'd46039, 16'd58564, 16'd47458, 16'd51138, 16'd54290, 16'd20961, 16'd412});
	test_expansion(128'hcfe530862c9f130bf8959e6e8733f0a4, {16'd59898, 16'd38928, 16'd6938, 16'd12515, 16'd64496, 16'd7608, 16'd10535, 16'd39484, 16'd43787, 16'd44853, 16'd34206, 16'd41254, 16'd43863, 16'd49650, 16'd37022, 16'd5482, 16'd44367, 16'd61530, 16'd2210, 16'd7782, 16'd46622, 16'd21947, 16'd20836, 16'd61358, 16'd64791, 16'd59972});
	test_expansion(128'hbc6cae85c23a216bb4d2aab242115e65, {16'd14802, 16'd11346, 16'd22581, 16'd38772, 16'd5515, 16'd4792, 16'd37944, 16'd45133, 16'd13179, 16'd27748, 16'd4297, 16'd36245, 16'd7540, 16'd59500, 16'd34039, 16'd42399, 16'd40326, 16'd49015, 16'd47646, 16'd27171, 16'd41440, 16'd19136, 16'd10210, 16'd10385, 16'd20955, 16'd26872});
	test_expansion(128'hda66623c259dccde1ef94f327737d8a0, {16'd31615, 16'd14933, 16'd5272, 16'd21132, 16'd27883, 16'd52966, 16'd15520, 16'd49317, 16'd871, 16'd38325, 16'd13730, 16'd57871, 16'd8261, 16'd1406, 16'd15754, 16'd20193, 16'd10876, 16'd39183, 16'd61919, 16'd65408, 16'd7354, 16'd8326, 16'd39112, 16'd32204, 16'd45470, 16'd32908});
	test_expansion(128'h0819e055baf03d4253197ecc99f17965, {16'd17913, 16'd54425, 16'd18491, 16'd6029, 16'd13055, 16'd60617, 16'd37951, 16'd14451, 16'd7609, 16'd12585, 16'd6194, 16'd41042, 16'd16949, 16'd59511, 16'd27816, 16'd3395, 16'd43825, 16'd22553, 16'd40786, 16'd46558, 16'd19400, 16'd29738, 16'd41998, 16'd26530, 16'd59948, 16'd37657});
	test_expansion(128'ha8363c2fd4d9b2985957671991d591f0, {16'd62078, 16'd47511, 16'd44037, 16'd41558, 16'd39269, 16'd44131, 16'd18572, 16'd33031, 16'd6805, 16'd24752, 16'd24127, 16'd62385, 16'd27415, 16'd28121, 16'd11641, 16'd48374, 16'd55150, 16'd7205, 16'd18640, 16'd54723, 16'd41117, 16'd44103, 16'd23220, 16'd33195, 16'd29163, 16'd18951});
	test_expansion(128'h633551551ba978f47a9c9d6198817dcf, {16'd21480, 16'd61479, 16'd56665, 16'd39379, 16'd32279, 16'd34018, 16'd11299, 16'd24056, 16'd48433, 16'd59426, 16'd4784, 16'd44513, 16'd14063, 16'd31829, 16'd28786, 16'd14067, 16'd25913, 16'd65234, 16'd4726, 16'd37078, 16'd15740, 16'd7765, 16'd42115, 16'd62265, 16'd52129, 16'd36663});
	test_expansion(128'hcd8ce53623127338dea58d52336076fa, {16'd55486, 16'd17399, 16'd14975, 16'd19469, 16'd40499, 16'd55025, 16'd48628, 16'd39661, 16'd49802, 16'd16773, 16'd50318, 16'd14928, 16'd55295, 16'd55332, 16'd11109, 16'd48985, 16'd37085, 16'd51011, 16'd9881, 16'd16364, 16'd53970, 16'd445, 16'd27475, 16'd25665, 16'd77, 16'd2223});
	test_expansion(128'hb5cf9cf804f3a73a204df9c622ca1977, {16'd33191, 16'd846, 16'd25464, 16'd28979, 16'd3882, 16'd55011, 16'd12601, 16'd28099, 16'd31665, 16'd444, 16'd32017, 16'd39655, 16'd44266, 16'd5253, 16'd19662, 16'd17436, 16'd44355, 16'd40280, 16'd19620, 16'd60760, 16'd31806, 16'd64185, 16'd64820, 16'd22072, 16'd8824, 16'd54109});
	test_expansion(128'hc56ade46094a666ea09efbcc43d5f07e, {16'd58596, 16'd38386, 16'd57168, 16'd25372, 16'd422, 16'd38109, 16'd5606, 16'd50133, 16'd765, 16'd8484, 16'd27971, 16'd30976, 16'd34434, 16'd20403, 16'd34357, 16'd46298, 16'd64672, 16'd29627, 16'd20015, 16'd37462, 16'd18223, 16'd13965, 16'd29978, 16'd42369, 16'd40432, 16'd51746});
	test_expansion(128'hca1949abdb56a8f54327c2847c4287d0, {16'd27081, 16'd13581, 16'd34389, 16'd57264, 16'd37222, 16'd45650, 16'd28481, 16'd47081, 16'd31372, 16'd8923, 16'd20331, 16'd26510, 16'd12912, 16'd24490, 16'd21168, 16'd65301, 16'd24518, 16'd62810, 16'd62278, 16'd32185, 16'd41525, 16'd24775, 16'd62018, 16'd23251, 16'd5697, 16'd56778});
	test_expansion(128'h524a93e6f7c8e456b37b7d4a091f8024, {16'd48861, 16'd29827, 16'd32359, 16'd60032, 16'd46677, 16'd56754, 16'd61439, 16'd42402, 16'd9365, 16'd16819, 16'd19679, 16'd40852, 16'd65338, 16'd17629, 16'd12295, 16'd34803, 16'd30659, 16'd14053, 16'd30504, 16'd41485, 16'd3526, 16'd2448, 16'd31212, 16'd40705, 16'd51665, 16'd12732});
	test_expansion(128'hac8dec057d78c4168df80736fc2c86a5, {16'd26723, 16'd37774, 16'd31242, 16'd56952, 16'd16272, 16'd19824, 16'd12856, 16'd53067, 16'd52055, 16'd47255, 16'd52018, 16'd20468, 16'd42537, 16'd9563, 16'd44440, 16'd57833, 16'd31231, 16'd35083, 16'd24818, 16'd61672, 16'd14276, 16'd13227, 16'd54302, 16'd20782, 16'd21872, 16'd3463});
	test_expansion(128'hdf9c735b9bc433d3dc56b466d2ebb96e, {16'd22383, 16'd61480, 16'd63625, 16'd33712, 16'd29485, 16'd53896, 16'd61326, 16'd57775, 16'd59963, 16'd49989, 16'd865, 16'd5146, 16'd43623, 16'd52111, 16'd52236, 16'd1130, 16'd55147, 16'd62193, 16'd59706, 16'd38417, 16'd3129, 16'd34424, 16'd42251, 16'd58012, 16'd50728, 16'd4129});
	test_expansion(128'ha851cd851bd49f0f28da7a9e683acd4e, {16'd12233, 16'd11161, 16'd4054, 16'd1763, 16'd4887, 16'd29331, 16'd21587, 16'd5440, 16'd26615, 16'd64706, 16'd54870, 16'd8758, 16'd9066, 16'd43585, 16'd3076, 16'd24319, 16'd55829, 16'd61615, 16'd28848, 16'd62073, 16'd26692, 16'd53546, 16'd18145, 16'd36086, 16'd50256, 16'd40196});
	test_expansion(128'ha0d37338a9d2308bf0f3f628d0c1ff98, {16'd33113, 16'd24582, 16'd36486, 16'd339, 16'd64046, 16'd38066, 16'd52673, 16'd52155, 16'd36592, 16'd3849, 16'd64772, 16'd23782, 16'd47088, 16'd59568, 16'd49102, 16'd42665, 16'd61840, 16'd20852, 16'd28799, 16'd53541, 16'd19318, 16'd48217, 16'd41819, 16'd4208, 16'd7713, 16'd13648});
	test_expansion(128'hb55fd199485d78e7d219ff8ed0df76a3, {16'd50617, 16'd56418, 16'd23294, 16'd19222, 16'd42716, 16'd53567, 16'd9380, 16'd29506, 16'd35361, 16'd40754, 16'd45287, 16'd45751, 16'd39565, 16'd59136, 16'd50601, 16'd37399, 16'd60672, 16'd10952, 16'd9467, 16'd62452, 16'd20771, 16'd42470, 16'd42122, 16'd54374, 16'd58229, 16'd44884});
	test_expansion(128'h81d230126c28a83573522191211af19a, {16'd52927, 16'd18047, 16'd36419, 16'd56765, 16'd13355, 16'd14490, 16'd34829, 16'd2573, 16'd20395, 16'd19660, 16'd39362, 16'd10615, 16'd12104, 16'd20043, 16'd37876, 16'd56148, 16'd40767, 16'd53571, 16'd16295, 16'd22136, 16'd48445, 16'd56942, 16'd41110, 16'd27552, 16'd51711, 16'd47});
	test_expansion(128'h7390b43510ccd3c63457531a2c0a6482, {16'd2110, 16'd43018, 16'd54589, 16'd62374, 16'd13214, 16'd65530, 16'd48627, 16'd50588, 16'd48635, 16'd10950, 16'd7913, 16'd51252, 16'd49970, 16'd51197, 16'd5897, 16'd3727, 16'd7873, 16'd54812, 16'd58018, 16'd364, 16'd14102, 16'd14988, 16'd17916, 16'd342, 16'd48689, 16'd52875});
	test_expansion(128'h1abc1242299d25ac43df6cf790ae6b0f, {16'd4269, 16'd15459, 16'd27243, 16'd2383, 16'd51781, 16'd31999, 16'd3525, 16'd1368, 16'd4957, 16'd53750, 16'd33508, 16'd2524, 16'd36588, 16'd9537, 16'd13204, 16'd41785, 16'd10537, 16'd3495, 16'd4218, 16'd47572, 16'd3398, 16'd32839, 16'd49333, 16'd52036, 16'd45907, 16'd44355});
	test_expansion(128'hcbdc154e99f1f3cc45a55eb0e03e3490, {16'd29175, 16'd32573, 16'd4379, 16'd15263, 16'd14275, 16'd17154, 16'd50790, 16'd29390, 16'd59327, 16'd33282, 16'd30167, 16'd20367, 16'd52981, 16'd53873, 16'd58371, 16'd51110, 16'd26518, 16'd16365, 16'd26273, 16'd16204, 16'd13281, 16'd33257, 16'd44665, 16'd17670, 16'd38659, 16'd10189});
	test_expansion(128'h85fa3b058b2f5a838bfd4361ee5c4d8a, {16'd6640, 16'd23412, 16'd52356, 16'd20778, 16'd49975, 16'd62351, 16'd57275, 16'd23192, 16'd16574, 16'd62046, 16'd17347, 16'd16116, 16'd54442, 16'd47493, 16'd29730, 16'd36044, 16'd2211, 16'd38162, 16'd34073, 16'd21051, 16'd63186, 16'd37263, 16'd49493, 16'd241, 16'd64058, 16'd22470});
	test_expansion(128'h10de35cef621df03c5e2e278e47c3b35, {16'd25903, 16'd49690, 16'd12301, 16'd29363, 16'd3745, 16'd47986, 16'd23772, 16'd12978, 16'd7960, 16'd35016, 16'd4773, 16'd26989, 16'd18192, 16'd59934, 16'd24226, 16'd62537, 16'd34347, 16'd21398, 16'd48789, 16'd27169, 16'd60094, 16'd45767, 16'd45088, 16'd8947, 16'd60518, 16'd37635});
	test_expansion(128'h06f327a87def25582f23e5d1ccc58d6f, {16'd62155, 16'd63141, 16'd29286, 16'd51451, 16'd45922, 16'd26882, 16'd6914, 16'd49059, 16'd65360, 16'd37014, 16'd42960, 16'd41710, 16'd3086, 16'd32347, 16'd14566, 16'd24951, 16'd279, 16'd25464, 16'd52660, 16'd10842, 16'd21144, 16'd52809, 16'd44026, 16'd47425, 16'd37640, 16'd12807});
	test_expansion(128'hafb13edf53a61133f7f6bf16a1d1fc36, {16'd63186, 16'd10503, 16'd48108, 16'd56251, 16'd50194, 16'd57137, 16'd5838, 16'd4223, 16'd25442, 16'd4682, 16'd47136, 16'd22735, 16'd51579, 16'd52364, 16'd9533, 16'd19683, 16'd61713, 16'd2113, 16'd8438, 16'd40255, 16'd16472, 16'd28309, 16'd2688, 16'd13959, 16'd43366, 16'd10567});
	test_expansion(128'h688d8dd52f153546cfc2aa5f1f851ad4, {16'd41192, 16'd29840, 16'd60783, 16'd2147, 16'd11139, 16'd41546, 16'd36851, 16'd15635, 16'd58683, 16'd38900, 16'd49002, 16'd26135, 16'd20561, 16'd26938, 16'd15414, 16'd5473, 16'd19205, 16'd55863, 16'd51676, 16'd34053, 16'd31453, 16'd63582, 16'd10667, 16'd989, 16'd52500, 16'd27950});
	test_expansion(128'h98c571babc618829d572ba990b0355d7, {16'd2089, 16'd39923, 16'd29298, 16'd58729, 16'd31310, 16'd46917, 16'd33203, 16'd5893, 16'd33089, 16'd761, 16'd29080, 16'd1241, 16'd4229, 16'd36679, 16'd7318, 16'd33987, 16'd30141, 16'd1331, 16'd37591, 16'd53957, 16'd53238, 16'd19665, 16'd21133, 16'd64614, 16'd32325, 16'd54339});
	test_expansion(128'h7dc66ab1b234c9cd00fc06c3a457c651, {16'd44355, 16'd30434, 16'd20645, 16'd26987, 16'd52918, 16'd53206, 16'd18794, 16'd32629, 16'd45448, 16'd11738, 16'd8079, 16'd64637, 16'd60910, 16'd53254, 16'd17031, 16'd31400, 16'd31055, 16'd51795, 16'd13544, 16'd41710, 16'd56613, 16'd24478, 16'd31149, 16'd6957, 16'd16491, 16'd6109});
	test_expansion(128'ha1cb41ba577c1aafbf5161e0a4f8cda9, {16'd20861, 16'd14442, 16'd26826, 16'd34879, 16'd56830, 16'd65481, 16'd61562, 16'd1978, 16'd22904, 16'd23829, 16'd57051, 16'd218, 16'd65274, 16'd16217, 16'd16615, 16'd46310, 16'd5026, 16'd45833, 16'd27451, 16'd30761, 16'd55379, 16'd26730, 16'd47333, 16'd53992, 16'd177, 16'd30411});
	test_expansion(128'hf9c7b5dd7479877e197b8349022b87e2, {16'd14185, 16'd61023, 16'd47533, 16'd48740, 16'd45036, 16'd36222, 16'd62199, 16'd42062, 16'd7525, 16'd45387, 16'd43522, 16'd13613, 16'd9559, 16'd62844, 16'd58713, 16'd49562, 16'd7934, 16'd54930, 16'd21460, 16'd56548, 16'd64485, 16'd47626, 16'd30880, 16'd25903, 16'd57560, 16'd64826});
	test_expansion(128'h58634d30a9a392e7dc8b7793d9630e5f, {16'd58417, 16'd31070, 16'd13939, 16'd50720, 16'd56828, 16'd60803, 16'd60517, 16'd9173, 16'd33767, 16'd12662, 16'd48833, 16'd22832, 16'd51795, 16'd19517, 16'd28457, 16'd34749, 16'd25563, 16'd34354, 16'd54350, 16'd4725, 16'd28458, 16'd1214, 16'd65235, 16'd2255, 16'd17529, 16'd39683});
	test_expansion(128'ha75cd70bdf4e017bcb514a981826d5fa, {16'd5091, 16'd29425, 16'd7883, 16'd65153, 16'd16430, 16'd2990, 16'd9306, 16'd13081, 16'd29868, 16'd39779, 16'd58511, 16'd23495, 16'd20250, 16'd39358, 16'd58548, 16'd30920, 16'd13016, 16'd26572, 16'd20432, 16'd48058, 16'd22812, 16'd31252, 16'd36625, 16'd25260, 16'd10018, 16'd50112});
	test_expansion(128'ha0be2282c093d1c252c9af21d0cffd31, {16'd13052, 16'd38158, 16'd40678, 16'd23841, 16'd55313, 16'd6752, 16'd8124, 16'd38585, 16'd8338, 16'd30096, 16'd62138, 16'd123, 16'd44415, 16'd42132, 16'd49354, 16'd21767, 16'd31479, 16'd6021, 16'd46785, 16'd24742, 16'd62096, 16'd34867, 16'd40157, 16'd17694, 16'd22386, 16'd8004});
	test_expansion(128'hd51a1a1ba1659acb3ea762001033955e, {16'd49526, 16'd23494, 16'd39933, 16'd50175, 16'd10829, 16'd52513, 16'd10504, 16'd39531, 16'd41778, 16'd61751, 16'd35137, 16'd33603, 16'd2481, 16'd11121, 16'd35171, 16'd22467, 16'd54720, 16'd23664, 16'd59360, 16'd2869, 16'd1825, 16'd19310, 16'd56277, 16'd21397, 16'd865, 16'd56543});
	test_expansion(128'h2edfc7f00fda70663b71bc5a50f72a1a, {16'd33929, 16'd19132, 16'd19243, 16'd48540, 16'd23417, 16'd44456, 16'd27059, 16'd8862, 16'd7108, 16'd31565, 16'd9313, 16'd54285, 16'd17429, 16'd42650, 16'd19404, 16'd18373, 16'd51878, 16'd51718, 16'd56490, 16'd10691, 16'd49329, 16'd33280, 16'd40151, 16'd19570, 16'd40857, 16'd18150});
	test_expansion(128'h0095123e79b60249abd5a04625b11d15, {16'd57487, 16'd6994, 16'd63354, 16'd53007, 16'd5230, 16'd3646, 16'd1854, 16'd8892, 16'd6056, 16'd13682, 16'd55233, 16'd22235, 16'd18643, 16'd51027, 16'd37723, 16'd38409, 16'd4916, 16'd21656, 16'd47425, 16'd16898, 16'd27501, 16'd35753, 16'd15105, 16'd20680, 16'd37404, 16'd56935});
	test_expansion(128'he51b10068b0a4c1f28701031e2491f05, {16'd52681, 16'd51911, 16'd28740, 16'd45960, 16'd16523, 16'd42728, 16'd40404, 16'd4587, 16'd59718, 16'd5715, 16'd53452, 16'd46972, 16'd4782, 16'd46474, 16'd34985, 16'd15148, 16'd33855, 16'd43022, 16'd9493, 16'd18917, 16'd52077, 16'd10501, 16'd57559, 16'd5564, 16'd13751, 16'd55454});
	test_expansion(128'hd35df1fd078911c09f787e6ba4b951f5, {16'd42082, 16'd56548, 16'd41997, 16'd54421, 16'd5027, 16'd49469, 16'd59784, 16'd10677, 16'd65202, 16'd45801, 16'd11687, 16'd53880, 16'd46245, 16'd51048, 16'd23000, 16'd41886, 16'd21298, 16'd19558, 16'd18721, 16'd59759, 16'd62444, 16'd61251, 16'd48944, 16'd28216, 16'd21476, 16'd6084});
	test_expansion(128'ha04e123c8e49cf283a662c391f149a58, {16'd47444, 16'd55046, 16'd23963, 16'd55808, 16'd11485, 16'd4255, 16'd55992, 16'd2545, 16'd33466, 16'd26409, 16'd5990, 16'd16084, 16'd37088, 16'd7343, 16'd9096, 16'd54390, 16'd13344, 16'd51445, 16'd58935, 16'd54687, 16'd51344, 16'd59829, 16'd5159, 16'd58070, 16'd39736, 16'd32549});
	test_expansion(128'h62c31dcda2f7c89934aaff3954f00de3, {16'd2612, 16'd37001, 16'd9343, 16'd40977, 16'd46874, 16'd42779, 16'd35593, 16'd28244, 16'd11462, 16'd36851, 16'd39184, 16'd19783, 16'd404, 16'd31899, 16'd13166, 16'd28606, 16'd12540, 16'd18804, 16'd21450, 16'd59083, 16'd27083, 16'd18553, 16'd30700, 16'd62820, 16'd36501, 16'd41522});
	test_expansion(128'h7bed080c8603e30a9df6eb22a4512cfa, {16'd54044, 16'd4715, 16'd1427, 16'd43012, 16'd7094, 16'd19494, 16'd51681, 16'd56111, 16'd17275, 16'd57848, 16'd33252, 16'd17433, 16'd38281, 16'd44287, 16'd13414, 16'd10984, 16'd5791, 16'd30273, 16'd47194, 16'd24777, 16'd20440, 16'd62706, 16'd17638, 16'd997, 16'd61372, 16'd55888});
	test_expansion(128'he17fe7a1af80fc7cd9406cbde89e980f, {16'd368, 16'd56446, 16'd22343, 16'd49932, 16'd60215, 16'd47542, 16'd58568, 16'd37302, 16'd55138, 16'd3854, 16'd48838, 16'd53334, 16'd49519, 16'd35693, 16'd27748, 16'd788, 16'd17590, 16'd65334, 16'd28283, 16'd64432, 16'd64550, 16'd19760, 16'd42735, 16'd41075, 16'd4067, 16'd57088});
	test_expansion(128'hf1644236148ca89c25feb1086bb943dc, {16'd48654, 16'd14448, 16'd17585, 16'd41195, 16'd43260, 16'd22694, 16'd6373, 16'd20350, 16'd19895, 16'd20199, 16'd37791, 16'd6417, 16'd8717, 16'd5848, 16'd41829, 16'd7578, 16'd13363, 16'd16625, 16'd33953, 16'd2773, 16'd22048, 16'd58466, 16'd56622, 16'd54738, 16'd3934, 16'd12980});
	test_expansion(128'hb32ea857df5c388c704211a78b0bf1d9, {16'd13215, 16'd47936, 16'd12231, 16'd44233, 16'd50586, 16'd34352, 16'd31969, 16'd62975, 16'd32858, 16'd52136, 16'd3311, 16'd3126, 16'd56806, 16'd55165, 16'd18896, 16'd51257, 16'd12404, 16'd27320, 16'd2746, 16'd39880, 16'd30673, 16'd35875, 16'd11141, 16'd40779, 16'd27681, 16'd56779});
	test_expansion(128'h75a191a8bbade7433d6860c33eddff3d, {16'd14741, 16'd40802, 16'd26114, 16'd36765, 16'd49958, 16'd8344, 16'd16632, 16'd44555, 16'd49077, 16'd126, 16'd585, 16'd11225, 16'd21114, 16'd27110, 16'd41191, 16'd64989, 16'd7687, 16'd18478, 16'd43461, 16'd29399, 16'd62012, 16'd36841, 16'd56240, 16'd54780, 16'd32253, 16'd17276});
	test_expansion(128'h42265f2b432edef646322e9db7ed75fa, {16'd57876, 16'd34392, 16'd19390, 16'd17259, 16'd35472, 16'd24598, 16'd25107, 16'd5052, 16'd36868, 16'd5214, 16'd20340, 16'd46876, 16'd5410, 16'd2951, 16'd19592, 16'd46724, 16'd59985, 16'd57713, 16'd22841, 16'd11057, 16'd8377, 16'd20728, 16'd50184, 16'd38642, 16'd63904, 16'd15547});
	test_expansion(128'h4abe2fba6888e5ce2fa24b95973cdab2, {16'd55543, 16'd56516, 16'd39428, 16'd8244, 16'd3660, 16'd35610, 16'd17471, 16'd39296, 16'd55852, 16'd13874, 16'd30443, 16'd58385, 16'd2870, 16'd7748, 16'd20549, 16'd9674, 16'd60162, 16'd54688, 16'd4739, 16'd2022, 16'd29109, 16'd54358, 16'd27215, 16'd35422, 16'd59911, 16'd64420});
	test_expansion(128'he4591b4c88bb0d0e86ebcde71e00e1f2, {16'd32498, 16'd40755, 16'd5545, 16'd12000, 16'd43052, 16'd27460, 16'd6982, 16'd31375, 16'd8106, 16'd54349, 16'd1157, 16'd23244, 16'd41210, 16'd34000, 16'd34528, 16'd34740, 16'd40531, 16'd53299, 16'd6475, 16'd43387, 16'd23036, 16'd15420, 16'd19501, 16'd8455, 16'd21827, 16'd2365});
	test_expansion(128'ha8ba9d8561c1ca2f9c74f75d7e62eff3, {16'd57328, 16'd1263, 16'd22335, 16'd57534, 16'd3901, 16'd61012, 16'd43524, 16'd61476, 16'd60817, 16'd58499, 16'd35163, 16'd58433, 16'd42685, 16'd25939, 16'd38765, 16'd31826, 16'd13385, 16'd55420, 16'd37666, 16'd42419, 16'd38637, 16'd34667, 16'd39683, 16'd58071, 16'd5440, 16'd24695});
	test_expansion(128'h2c9a17c8ad41827ae3f2d9f273265ce4, {16'd15773, 16'd46361, 16'd27707, 16'd29126, 16'd27597, 16'd49454, 16'd30448, 16'd12390, 16'd65369, 16'd54007, 16'd39508, 16'd43789, 16'd48231, 16'd58131, 16'd61837, 16'd63486, 16'd51934, 16'd15171, 16'd29170, 16'd48440, 16'd44158, 16'd16490, 16'd30330, 16'd63283, 16'd8736, 16'd35443});
	test_expansion(128'hb61f839c9f57eb186d1673d2d5a04bf4, {16'd5307, 16'd60964, 16'd62365, 16'd10002, 16'd16116, 16'd1051, 16'd46077, 16'd40276, 16'd1942, 16'd11022, 16'd26052, 16'd32073, 16'd43489, 16'd17652, 16'd16311, 16'd41666, 16'd6387, 16'd33740, 16'd44105, 16'd18981, 16'd15777, 16'd1569, 16'd26071, 16'd6648, 16'd7434, 16'd46926});
	test_expansion(128'hea7716c93a4e639cb468d0cbdafb278e, {16'd57904, 16'd11261, 16'd48907, 16'd35141, 16'd42120, 16'd19321, 16'd62558, 16'd63654, 16'd17502, 16'd56802, 16'd21983, 16'd43460, 16'd41308, 16'd64742, 16'd40856, 16'd24079, 16'd17043, 16'd28719, 16'd50365, 16'd2887, 16'd16238, 16'd33863, 16'd52009, 16'd807, 16'd29984, 16'd17177});
	test_expansion(128'hc19bb32cfdb31ec8634e5961158660f3, {16'd9691, 16'd48122, 16'd7402, 16'd13675, 16'd17607, 16'd8533, 16'd53319, 16'd14148, 16'd29199, 16'd7147, 16'd57436, 16'd28333, 16'd11564, 16'd42666, 16'd31196, 16'd6887, 16'd6015, 16'd55809, 16'd62943, 16'd24299, 16'd17424, 16'd49358, 16'd30023, 16'd50143, 16'd452, 16'd31972});
	test_expansion(128'h4eb1b8f30cedf49e9da1de0b7512118b, {16'd39873, 16'd34284, 16'd54484, 16'd51307, 16'd27571, 16'd34775, 16'd25350, 16'd18624, 16'd52495, 16'd11486, 16'd36324, 16'd3552, 16'd26450, 16'd58011, 16'd4540, 16'd42477, 16'd38326, 16'd54080, 16'd27604, 16'd13516, 16'd40216, 16'd17917, 16'd18820, 16'd44152, 16'd64702, 16'd15018});
	test_expansion(128'h2aebee18f03effea3c9c5f7fcd6d1e34, {16'd42168, 16'd61085, 16'd7678, 16'd20480, 16'd57855, 16'd14152, 16'd4106, 16'd34137, 16'd54299, 16'd35702, 16'd24839, 16'd22910, 16'd46117, 16'd5440, 16'd32277, 16'd56191, 16'd58838, 16'd17286, 16'd59104, 16'd35919, 16'd44929, 16'd57573, 16'd64881, 16'd11086, 16'd47731, 16'd30966});
	test_expansion(128'h52f77f7ff3e113e3e14ebe1f79108525, {16'd32002, 16'd34562, 16'd23321, 16'd35084, 16'd37291, 16'd7, 16'd11670, 16'd37485, 16'd20493, 16'd30590, 16'd44364, 16'd40650, 16'd30076, 16'd33097, 16'd32958, 16'd26158, 16'd57557, 16'd49600, 16'd20842, 16'd22213, 16'd7152, 16'd6541, 16'd42126, 16'd29116, 16'd4434, 16'd24698});
	test_expansion(128'hbd7e68454059736fa9234b19dde0af54, {16'd55553, 16'd2055, 16'd64793, 16'd2469, 16'd59917, 16'd20551, 16'd64527, 16'd8301, 16'd16631, 16'd155, 16'd29031, 16'd1942, 16'd45568, 16'd31898, 16'd44538, 16'd47558, 16'd3634, 16'd32402, 16'd40984, 16'd26169, 16'd17601, 16'd59936, 16'd23474, 16'd41194, 16'd50955, 16'd25338});
	test_expansion(128'h90a20cef92c828456d55b7f491f14ab5, {16'd4082, 16'd32774, 16'd35082, 16'd25945, 16'd9175, 16'd34424, 16'd1670, 16'd1932, 16'd44925, 16'd14303, 16'd51318, 16'd19574, 16'd32794, 16'd28147, 16'd23982, 16'd39109, 16'd56706, 16'd8301, 16'd35805, 16'd60080, 16'd16798, 16'd39791, 16'd57623, 16'd31154, 16'd23415, 16'd59017});
	test_expansion(128'he25afe0455c0c0599f3aaa58c9c34ee8, {16'd7050, 16'd60484, 16'd33859, 16'd13356, 16'd18593, 16'd29363, 16'd11576, 16'd56852, 16'd1608, 16'd32256, 16'd7426, 16'd33813, 16'd45981, 16'd31236, 16'd28811, 16'd27518, 16'd36606, 16'd32313, 16'd52819, 16'd50376, 16'd42038, 16'd25691, 16'd22649, 16'd2786, 16'd1573, 16'd61563});
	test_expansion(128'hba6955410f096add0d7e5a800f521d5d, {16'd41709, 16'd15842, 16'd41664, 16'd18722, 16'd2777, 16'd57894, 16'd56178, 16'd24973, 16'd22468, 16'd5222, 16'd38887, 16'd40821, 16'd45802, 16'd58012, 16'd8095, 16'd23546, 16'd65408, 16'd59088, 16'd10929, 16'd30941, 16'd7380, 16'd34790, 16'd31230, 16'd35756, 16'd16222, 16'd9895});
	test_expansion(128'h6fc705d75b9528f292f87a88600893bc, {16'd36414, 16'd55784, 16'd43433, 16'd60234, 16'd37263, 16'd24034, 16'd17760, 16'd31324, 16'd50455, 16'd36629, 16'd37042, 16'd61043, 16'd5637, 16'd21676, 16'd57951, 16'd57971, 16'd9424, 16'd15295, 16'd2292, 16'd29260, 16'd13231, 16'd46031, 16'd48651, 16'd47706, 16'd1001, 16'd13147});
	test_expansion(128'heb40e7552233942ea801c568c8eae052, {16'd39589, 16'd8595, 16'd15409, 16'd24515, 16'd45636, 16'd38526, 16'd34460, 16'd64919, 16'd15962, 16'd6931, 16'd16927, 16'd914, 16'd17510, 16'd45497, 16'd56104, 16'd34010, 16'd10602, 16'd12680, 16'd9557, 16'd61238, 16'd9490, 16'd8964, 16'd37618, 16'd64552, 16'd52118, 16'd27156});
	test_expansion(128'ha431687cd6218dded92770437ee55f62, {16'd26958, 16'd55408, 16'd12320, 16'd36460, 16'd42299, 16'd48368, 16'd48736, 16'd1113, 16'd9631, 16'd17116, 16'd59076, 16'd60134, 16'd25084, 16'd25649, 16'd37603, 16'd20505, 16'd28547, 16'd11192, 16'd44007, 16'd19537, 16'd20761, 16'd24495, 16'd58709, 16'd65168, 16'd16560, 16'd29764});
	test_expansion(128'h5a65515e18fab72822a6b595de7862c1, {16'd62853, 16'd46511, 16'd49440, 16'd61193, 16'd3342, 16'd13044, 16'd39107, 16'd65289, 16'd1331, 16'd49316, 16'd59325, 16'd12179, 16'd65309, 16'd48508, 16'd18913, 16'd29668, 16'd21708, 16'd58433, 16'd21820, 16'd14477, 16'd28622, 16'd62339, 16'd64559, 16'd7506, 16'd62200, 16'd64514});
	test_expansion(128'h5ddefac0d50bb7a94e52736224e1554b, {16'd20229, 16'd35705, 16'd24023, 16'd46858, 16'd22104, 16'd36202, 16'd1262, 16'd21781, 16'd15388, 16'd40575, 16'd6530, 16'd60244, 16'd29437, 16'd63778, 16'd15186, 16'd45409, 16'd19024, 16'd710, 16'd19310, 16'd212, 16'd58488, 16'd64265, 16'd47776, 16'd42090, 16'd48352, 16'd63712});
	test_expansion(128'h9c6caad58e9ffe822212d2ba73ef55cc, {16'd17716, 16'd33472, 16'd30160, 16'd8659, 16'd12511, 16'd36446, 16'd31085, 16'd34489, 16'd748, 16'd64668, 16'd1985, 16'd38873, 16'd36628, 16'd32621, 16'd26564, 16'd5850, 16'd28892, 16'd49359, 16'd30472, 16'd32044, 16'd53504, 16'd13566, 16'd615, 16'd24739, 16'd19280, 16'd11315});
	test_expansion(128'he64449208dda0c8e4e0c5e01bd6eca49, {16'd43060, 16'd41046, 16'd30651, 16'd31150, 16'd33109, 16'd44988, 16'd30394, 16'd19706, 16'd9615, 16'd10845, 16'd53903, 16'd7629, 16'd57787, 16'd25139, 16'd57082, 16'd16914, 16'd24508, 16'd62899, 16'd49910, 16'd35559, 16'd8452, 16'd24699, 16'd62244, 16'd7748, 16'd2127, 16'd1870});
	test_expansion(128'hc4e0f287f2eb392ce01efd746b793ba0, {16'd38617, 16'd35671, 16'd35436, 16'd42646, 16'd64281, 16'd11083, 16'd54074, 16'd49734, 16'd60212, 16'd43407, 16'd37001, 16'd50885, 16'd48315, 16'd17657, 16'd38117, 16'd11222, 16'd43760, 16'd25620, 16'd46852, 16'd24846, 16'd38799, 16'd1563, 16'd14266, 16'd62215, 16'd46712, 16'd56530});
	test_expansion(128'h42f075bbee7b3e9fc31faeec2b6e8abc, {16'd38218, 16'd41693, 16'd10345, 16'd48764, 16'd32246, 16'd17940, 16'd46340, 16'd23201, 16'd3488, 16'd41882, 16'd31087, 16'd41027, 16'd40954, 16'd22554, 16'd6417, 16'd17514, 16'd24748, 16'd14474, 16'd24396, 16'd39499, 16'd25967, 16'd23706, 16'd60265, 16'd33202, 16'd12114, 16'd31599});
	test_expansion(128'h73d36152309a51da60ba45755faf13ca, {16'd5454, 16'd14033, 16'd29064, 16'd1241, 16'd812, 16'd39949, 16'd56544, 16'd15078, 16'd24149, 16'd55232, 16'd46874, 16'd38999, 16'd61958, 16'd59333, 16'd30744, 16'd59360, 16'd12028, 16'd47036, 16'd61228, 16'd62442, 16'd2145, 16'd46376, 16'd34921, 16'd52996, 16'd62155, 16'd63513});
	test_expansion(128'ha62e32d9997dc81b7463a269131998a2, {16'd39747, 16'd12301, 16'd48736, 16'd52591, 16'd7545, 16'd53916, 16'd2017, 16'd63589, 16'd37374, 16'd22910, 16'd61835, 16'd33475, 16'd59107, 16'd61809, 16'd61273, 16'd36476, 16'd46334, 16'd15229, 16'd15197, 16'd22931, 16'd5150, 16'd57563, 16'd27909, 16'd23433, 16'd61998, 16'd32662});
	test_expansion(128'h7d2f9fd8c590ff7c2f806703cfefae66, {16'd48221, 16'd21095, 16'd17239, 16'd62807, 16'd51915, 16'd10625, 16'd52755, 16'd11319, 16'd35172, 16'd5175, 16'd23948, 16'd37464, 16'd28146, 16'd58556, 16'd46791, 16'd19847, 16'd45504, 16'd21204, 16'd48363, 16'd48995, 16'd743, 16'd57598, 16'd61207, 16'd8922, 16'd37819, 16'd49873});
	test_expansion(128'h557a4e1e13222ddbb2451dbe04137850, {16'd51963, 16'd11155, 16'd31832, 16'd61241, 16'd42621, 16'd44738, 16'd15869, 16'd55190, 16'd43254, 16'd55569, 16'd14113, 16'd40421, 16'd55546, 16'd35240, 16'd33019, 16'd2459, 16'd20816, 16'd27837, 16'd61619, 16'd20714, 16'd1604, 16'd56971, 16'd12132, 16'd53536, 16'd11273, 16'd27787});
	test_expansion(128'h80ed7ed48dcbdc5d3e92de6661339ea4, {16'd6289, 16'd48061, 16'd41996, 16'd9752, 16'd27034, 16'd56635, 16'd22521, 16'd64902, 16'd25850, 16'd3711, 16'd34420, 16'd50554, 16'd25472, 16'd52135, 16'd34652, 16'd33428, 16'd13669, 16'd20337, 16'd36602, 16'd7839, 16'd15586, 16'd45756, 16'd15349, 16'd53652, 16'd31327, 16'd24695});
	test_expansion(128'h94e0ffc362404a8c43a865b040543748, {16'd13276, 16'd374, 16'd47275, 16'd42240, 16'd43048, 16'd61283, 16'd11958, 16'd22275, 16'd19931, 16'd40073, 16'd39198, 16'd59923, 16'd5287, 16'd31110, 16'd27316, 16'd45296, 16'd6051, 16'd40552, 16'd43899, 16'd52841, 16'd19771, 16'd13210, 16'd60199, 16'd29364, 16'd11384, 16'd9550});
	test_expansion(128'h9e72a9f57940f76d8b7ddda27c78dd7d, {16'd56990, 16'd19266, 16'd15265, 16'd65453, 16'd26191, 16'd43343, 16'd40510, 16'd48588, 16'd34469, 16'd34435, 16'd59537, 16'd64749, 16'd1179, 16'd58447, 16'd15558, 16'd62267, 16'd24214, 16'd44344, 16'd21211, 16'd51412, 16'd7235, 16'd14131, 16'd23340, 16'd12987, 16'd39267, 16'd44070});
	test_expansion(128'h1525a70db31f8dde9611f388e715cd60, {16'd24038, 16'd17684, 16'd14217, 16'd41266, 16'd36163, 16'd37108, 16'd21911, 16'd8686, 16'd58369, 16'd55841, 16'd223, 16'd49760, 16'd31656, 16'd58218, 16'd41016, 16'd63714, 16'd15483, 16'd36283, 16'd52831, 16'd58006, 16'd1337, 16'd27150, 16'd47706, 16'd35222, 16'd54480, 16'd7945});
	test_expansion(128'h55c54b43802ae8141f4b09f2445df7f8, {16'd53938, 16'd51978, 16'd48378, 16'd30865, 16'd52977, 16'd47908, 16'd60831, 16'd65289, 16'd9020, 16'd50976, 16'd36800, 16'd3169, 16'd40813, 16'd18367, 16'd7338, 16'd35146, 16'd15188, 16'd51317, 16'd27677, 16'd48455, 16'd34438, 16'd2029, 16'd23814, 16'd9707, 16'd20256, 16'd28494});
	test_expansion(128'h352e6197854c5243186ba26ad0245802, {16'd41661, 16'd17054, 16'd59885, 16'd55487, 16'd40978, 16'd43299, 16'd24558, 16'd28197, 16'd55423, 16'd13220, 16'd35345, 16'd6661, 16'd57162, 16'd41263, 16'd41671, 16'd29051, 16'd7829, 16'd40445, 16'd61198, 16'd60341, 16'd27116, 16'd45395, 16'd21767, 16'd31347, 16'd31511, 16'd2230});
	test_expansion(128'h25f5176c170f37b2562afb85976aee1a, {16'd60285, 16'd3179, 16'd52283, 16'd26934, 16'd54691, 16'd18731, 16'd25618, 16'd60009, 16'd4319, 16'd44653, 16'd4456, 16'd15860, 16'd26103, 16'd48127, 16'd44285, 16'd33972, 16'd11273, 16'd47928, 16'd48629, 16'd13963, 16'd53789, 16'd62695, 16'd7141, 16'd49379, 16'd40356, 16'd7773});
	test_expansion(128'he9261eefb7d3c3e0dc9405343f66e83a, {16'd62585, 16'd61552, 16'd52353, 16'd54662, 16'd12945, 16'd6950, 16'd33801, 16'd64441, 16'd20937, 16'd40374, 16'd37686, 16'd35134, 16'd42554, 16'd13273, 16'd40457, 16'd47915, 16'd7800, 16'd46402, 16'd55055, 16'd48606, 16'd52578, 16'd62796, 16'd30498, 16'd1352, 16'd36078, 16'd40699});
	test_expansion(128'habfa684d39f5ebf721a55ae62e6bd7d5, {16'd53815, 16'd26102, 16'd58142, 16'd21556, 16'd33372, 16'd26755, 16'd59574, 16'd44281, 16'd21825, 16'd62412, 16'd23510, 16'd52029, 16'd25284, 16'd50318, 16'd21430, 16'd33573, 16'd37456, 16'd15416, 16'd32998, 16'd17233, 16'd61794, 16'd58966, 16'd15628, 16'd21758, 16'd45742, 16'd32601});
	test_expansion(128'h4e1ecc17e192983e130c00e65ae81896, {16'd37112, 16'd8887, 16'd4128, 16'd22153, 16'd53892, 16'd24877, 16'd13957, 16'd2889, 16'd7765, 16'd63175, 16'd36858, 16'd11534, 16'd63742, 16'd57158, 16'd22932, 16'd53646, 16'd33807, 16'd15131, 16'd11380, 16'd37391, 16'd2648, 16'd22663, 16'd26728, 16'd28039, 16'd44927, 16'd54343});
	test_expansion(128'h01ab8747504f42178250749abb3b08c9, {16'd57990, 16'd65333, 16'd40533, 16'd1383, 16'd24461, 16'd43708, 16'd63644, 16'd26212, 16'd8487, 16'd47374, 16'd20053, 16'd60703, 16'd57215, 16'd57082, 16'd27424, 16'd39532, 16'd57801, 16'd36583, 16'd49791, 16'd1176, 16'd49346, 16'd39241, 16'd38114, 16'd158, 16'd43139, 16'd43964});
	test_expansion(128'h26039f1c84501de28c828272bdbb46a7, {16'd52196, 16'd5183, 16'd292, 16'd30193, 16'd57926, 16'd41321, 16'd10474, 16'd57288, 16'd55286, 16'd41711, 16'd38109, 16'd42695, 16'd4383, 16'd20691, 16'd26284, 16'd35230, 16'd62833, 16'd45950, 16'd3088, 16'd5952, 16'd50631, 16'd29672, 16'd29037, 16'd12631, 16'd27662, 16'd54840});
	test_expansion(128'h83ce7459ae407aba9d25f8e84bf71d3c, {16'd20122, 16'd15463, 16'd44839, 16'd42317, 16'd28056, 16'd51250, 16'd5043, 16'd34222, 16'd5260, 16'd15098, 16'd20367, 16'd52370, 16'd7848, 16'd57312, 16'd28189, 16'd16326, 16'd17491, 16'd13575, 16'd49139, 16'd54261, 16'd24492, 16'd31062, 16'd21865, 16'd12380, 16'd9446, 16'd1141});
	test_expansion(128'h354a2e63b58c63570cc62d5f9f3a09dc, {16'd3766, 16'd34320, 16'd50151, 16'd8499, 16'd50887, 16'd28065, 16'd64770, 16'd55410, 16'd61873, 16'd59676, 16'd34934, 16'd24140, 16'd48634, 16'd19413, 16'd31047, 16'd8468, 16'd26542, 16'd14155, 16'd37133, 16'd51740, 16'd62202, 16'd26188, 16'd5426, 16'd13835, 16'd47731, 16'd60496});
	test_expansion(128'h14099c1990dd5d12f9820ed7df983a2d, {16'd37642, 16'd26739, 16'd47891, 16'd47049, 16'd23840, 16'd36517, 16'd43193, 16'd1713, 16'd52911, 16'd35165, 16'd41343, 16'd6840, 16'd60525, 16'd4386, 16'd20394, 16'd65005, 16'd28207, 16'd62732, 16'd5473, 16'd48718, 16'd43086, 16'd56745, 16'd52715, 16'd11710, 16'd8699, 16'd53082});
	test_expansion(128'h0e71c47a93f6cd6fca848d13bb574bb7, {16'd35611, 16'd20554, 16'd4893, 16'd63354, 16'd32379, 16'd45594, 16'd58158, 16'd23691, 16'd32586, 16'd56822, 16'd62384, 16'd24730, 16'd273, 16'd39070, 16'd63937, 16'd11085, 16'd43240, 16'd55434, 16'd21840, 16'd182, 16'd7305, 16'd45610, 16'd18956, 16'd24967, 16'd20256, 16'd49288});
	test_expansion(128'he434afb9f88e0f54df01874dbdd152e6, {16'd667, 16'd34179, 16'd20058, 16'd38604, 16'd3602, 16'd56072, 16'd16980, 16'd22350, 16'd50385, 16'd10672, 16'd42802, 16'd58377, 16'd61027, 16'd55898, 16'd50358, 16'd9800, 16'd44475, 16'd25985, 16'd36982, 16'd1641, 16'd63223, 16'd41904, 16'd12349, 16'd28060, 16'd9532, 16'd62455});
	test_expansion(128'h1eec005b44ecf0c5218c1c1259d34aca, {16'd44586, 16'd16040, 16'd25224, 16'd49161, 16'd55968, 16'd12608, 16'd30190, 16'd9330, 16'd23721, 16'd9830, 16'd22759, 16'd25998, 16'd56581, 16'd23210, 16'd42530, 16'd36356, 16'd62688, 16'd41521, 16'd4640, 16'd11167, 16'd46028, 16'd37390, 16'd60276, 16'd28509, 16'd43805, 16'd27214});
	test_expansion(128'h206fb46347e1ed6211072d4a505a8044, {16'd8665, 16'd5534, 16'd46351, 16'd34529, 16'd42723, 16'd22258, 16'd44287, 16'd16253, 16'd24708, 16'd35775, 16'd60243, 16'd58240, 16'd55881, 16'd52533, 16'd4103, 16'd64918, 16'd19874, 16'd5593, 16'd27332, 16'd65364, 16'd57932, 16'd3157, 16'd994, 16'd55933, 16'd64548, 16'd15642});
	test_expansion(128'hf0e31ca3f1eb1c87df009393a83f7d04, {16'd52517, 16'd2437, 16'd29005, 16'd55034, 16'd59452, 16'd39441, 16'd36739, 16'd15538, 16'd36966, 16'd16184, 16'd17830, 16'd1345, 16'd2300, 16'd36168, 16'd26625, 16'd61655, 16'd18389, 16'd61853, 16'd48230, 16'd43403, 16'd16335, 16'd28074, 16'd6508, 16'd28266, 16'd6771, 16'd18319});
	test_expansion(128'ha9f6a12de11065d99c1cf51b35bcfcbe, {16'd28091, 16'd36604, 16'd50238, 16'd14679, 16'd28425, 16'd58272, 16'd23084, 16'd31562, 16'd41197, 16'd41754, 16'd59924, 16'd25807, 16'd52646, 16'd54794, 16'd58941, 16'd31766, 16'd63635, 16'd3941, 16'd26549, 16'd30243, 16'd47106, 16'd39345, 16'd3430, 16'd50023, 16'd48390, 16'd47320});
	test_expansion(128'h67deca990354978a160972ce2aa49479, {16'd18793, 16'd21629, 16'd45528, 16'd29516, 16'd51074, 16'd57582, 16'd31851, 16'd8764, 16'd28674, 16'd36355, 16'd251, 16'd50462, 16'd30330, 16'd19632, 16'd28097, 16'd53369, 16'd33804, 16'd53343, 16'd1847, 16'd36904, 16'd54059, 16'd5561, 16'd36952, 16'd43644, 16'd7134, 16'd23252});
	test_expansion(128'heb3d756505ea39055cbfacd44127ec5f, {16'd64631, 16'd17116, 16'd62715, 16'd14697, 16'd35570, 16'd54587, 16'd41734, 16'd32083, 16'd27917, 16'd36977, 16'd11911, 16'd52525, 16'd39303, 16'd64800, 16'd17568, 16'd24034, 16'd50754, 16'd12086, 16'd59733, 16'd41250, 16'd33672, 16'd30824, 16'd58281, 16'd50558, 16'd54194, 16'd34881});
	test_expansion(128'h1fbf8438cc4c02c8fcb4342bf9f2b4b0, {16'd15196, 16'd43589, 16'd10211, 16'd20836, 16'd44440, 16'd17791, 16'd13648, 16'd2009, 16'd48777, 16'd3558, 16'd55193, 16'd7889, 16'd1100, 16'd9860, 16'd3133, 16'd58338, 16'd41018, 16'd62583, 16'd54180, 16'd36646, 16'd22783, 16'd21177, 16'd31454, 16'd50822, 16'd12539, 16'd35582});
	test_expansion(128'h72043083a700ece8c9485d19c44577a2, {16'd18774, 16'd53016, 16'd24430, 16'd35598, 16'd14810, 16'd51333, 16'd3988, 16'd27, 16'd6025, 16'd50810, 16'd57456, 16'd16316, 16'd31745, 16'd58129, 16'd57802, 16'd16004, 16'd20722, 16'd472, 16'd2440, 16'd20595, 16'd54155, 16'd9797, 16'd60765, 16'd54444, 16'd22134, 16'd48932});
	test_expansion(128'hadf7819ab2faba56359553266f3b0a0d, {16'd36525, 16'd58604, 16'd64935, 16'd4283, 16'd42266, 16'd35829, 16'd32650, 16'd41725, 16'd9308, 16'd54440, 16'd63453, 16'd3681, 16'd33912, 16'd7007, 16'd26598, 16'd27432, 16'd54665, 16'd32206, 16'd10542, 16'd12997, 16'd43173, 16'd57803, 16'd55148, 16'd14283, 16'd59299, 16'd2702});
	test_expansion(128'ha266d856aa4533c653142379bd2ff3e0, {16'd23262, 16'd33104, 16'd40686, 16'd42617, 16'd25560, 16'd20475, 16'd30490, 16'd60322, 16'd1713, 16'd34031, 16'd40641, 16'd59749, 16'd60646, 16'd59825, 16'd59577, 16'd4098, 16'd64373, 16'd41471, 16'd62353, 16'd20913, 16'd46816, 16'd2709, 16'd26072, 16'd39210, 16'd43116, 16'd27983});
	test_expansion(128'h45d6cff2f338ae5d8fd931b83273d133, {16'd62545, 16'd61179, 16'd6265, 16'd44975, 16'd65380, 16'd36427, 16'd2555, 16'd5907, 16'd24577, 16'd15770, 16'd51350, 16'd34850, 16'd26640, 16'd6248, 16'd47686, 16'd14084, 16'd49499, 16'd12803, 16'd57032, 16'd31819, 16'd28040, 16'd7298, 16'd40961, 16'd56021, 16'd4319, 16'd27498});
	test_expansion(128'ha4bdbac3dde147be07b84577928299f1, {16'd41704, 16'd22609, 16'd43264, 16'd54422, 16'd27949, 16'd58404, 16'd32612, 16'd60606, 16'd57264, 16'd48583, 16'd1341, 16'd46489, 16'd53897, 16'd19581, 16'd51208, 16'd63775, 16'd6847, 16'd60024, 16'd42965, 16'd3212, 16'd37999, 16'd17234, 16'd30163, 16'd42137, 16'd63690, 16'd21630});
	test_expansion(128'he61805622f0852278b6f1b00346b0f90, {16'd20209, 16'd40180, 16'd9738, 16'd36849, 16'd61487, 16'd13600, 16'd50443, 16'd15826, 16'd26911, 16'd8277, 16'd8504, 16'd26221, 16'd28537, 16'd9732, 16'd36751, 16'd35424, 16'd43478, 16'd53777, 16'd33100, 16'd32746, 16'd30753, 16'd33490, 16'd25815, 16'd2135, 16'd57248, 16'd5545});
	test_expansion(128'hb961eacd2d57f5dc72fbf6d503a5dd3a, {16'd25490, 16'd57214, 16'd40735, 16'd48883, 16'd45768, 16'd61155, 16'd45338, 16'd39071, 16'd16550, 16'd20778, 16'd60183, 16'd20622, 16'd50149, 16'd18288, 16'd46472, 16'd27796, 16'd30180, 16'd29598, 16'd21196, 16'd64746, 16'd743, 16'd41548, 16'd813, 16'd17711, 16'd1844, 16'd42429});
	test_expansion(128'hb5283071d72c961b4fcd138003345eaf, {16'd35094, 16'd39487, 16'd65011, 16'd29551, 16'd48006, 16'd21240, 16'd919, 16'd64301, 16'd30547, 16'd39972, 16'd62218, 16'd26842, 16'd13628, 16'd39655, 16'd29315, 16'd29922, 16'd2478, 16'd38717, 16'd42504, 16'd25985, 16'd35683, 16'd31134, 16'd2034, 16'd46282, 16'd19908, 16'd1385});
	test_expansion(128'hfcfa35d3b64117fdc626cca9beb4b1d2, {16'd44242, 16'd24684, 16'd60032, 16'd1663, 16'd39663, 16'd12816, 16'd5016, 16'd27099, 16'd18278, 16'd3489, 16'd1212, 16'd42965, 16'd62731, 16'd40433, 16'd27677, 16'd26486, 16'd7039, 16'd47482, 16'd65267, 16'd4430, 16'd15835, 16'd45220, 16'd62603, 16'd11167, 16'd28051, 16'd14668});
	test_expansion(128'hb5f5f6ff85dc6e0c4fdd002e152206c7, {16'd28095, 16'd42406, 16'd23504, 16'd56165, 16'd8520, 16'd5685, 16'd7955, 16'd2858, 16'd51292, 16'd38287, 16'd24189, 16'd55928, 16'd5002, 16'd30463, 16'd42123, 16'd17974, 16'd17959, 16'd10205, 16'd14506, 16'd15122, 16'd49009, 16'd25359, 16'd17706, 16'd42045, 16'd28664, 16'd12461});
	test_expansion(128'h534e50d84ffec295b8067cbeb4ca8b37, {16'd11243, 16'd46307, 16'd60286, 16'd64240, 16'd29595, 16'd27804, 16'd4445, 16'd56255, 16'd42766, 16'd59229, 16'd58865, 16'd51449, 16'd30936, 16'd63729, 16'd53276, 16'd12354, 16'd60087, 16'd14710, 16'd17299, 16'd14462, 16'd17608, 16'd54228, 16'd46966, 16'd2871, 16'd46991, 16'd6672});
	test_expansion(128'hb1c0ff93ef576f13e7f13ce79377d7b5, {16'd10632, 16'd53382, 16'd25118, 16'd45135, 16'd25327, 16'd63170, 16'd41067, 16'd63950, 16'd60482, 16'd46589, 16'd21277, 16'd58779, 16'd30659, 16'd27585, 16'd61527, 16'd60743, 16'd44593, 16'd56260, 16'd9163, 16'd60201, 16'd52618, 16'd42560, 16'd21467, 16'd30865, 16'd19249, 16'd45472});
	test_expansion(128'h54cb7f0c2a53516cb65a0b9e34cdb832, {16'd20869, 16'd24577, 16'd55516, 16'd59796, 16'd43434, 16'd2198, 16'd23215, 16'd18440, 16'd35131, 16'd4181, 16'd10840, 16'd7628, 16'd2890, 16'd39872, 16'd9704, 16'd46465, 16'd54504, 16'd25359, 16'd23164, 16'd59081, 16'd50163, 16'd37305, 16'd57575, 16'd40918, 16'd49163, 16'd40294});
	test_expansion(128'h2a0a5becf485ddff3cdbaa805347e067, {16'd5682, 16'd6883, 16'd26467, 16'd15882, 16'd29346, 16'd23382, 16'd24, 16'd50449, 16'd39182, 16'd52645, 16'd2197, 16'd23433, 16'd9754, 16'd28240, 16'd32787, 16'd13027, 16'd44112, 16'd25356, 16'd3120, 16'd52006, 16'd55352, 16'd37592, 16'd33680, 16'd10248, 16'd3822, 16'd32622});
	test_expansion(128'h7e1ae636e2fd0ecbb58a0c8145cafa4e, {16'd7889, 16'd42446, 16'd54996, 16'd36799, 16'd9141, 16'd45844, 16'd232, 16'd43268, 16'd23518, 16'd24879, 16'd35699, 16'd28113, 16'd48892, 16'd58364, 16'd11259, 16'd10359, 16'd62396, 16'd28799, 16'd19760, 16'd34325, 16'd64944, 16'd28780, 16'd46097, 16'd14579, 16'd17143, 16'd14831});
	test_expansion(128'h943d92f453756b922181cfacf03c5825, {16'd57528, 16'd20181, 16'd36877, 16'd49706, 16'd9358, 16'd41933, 16'd17111, 16'd28384, 16'd23552, 16'd63087, 16'd32276, 16'd40365, 16'd44716, 16'd21474, 16'd13301, 16'd22620, 16'd1032, 16'd43661, 16'd33456, 16'd15434, 16'd1679, 16'd20248, 16'd4102, 16'd43055, 16'd33862, 16'd22608});
	test_expansion(128'h38ad8480cb1c489dd372178c58695183, {16'd4833, 16'd42188, 16'd19022, 16'd39889, 16'd23198, 16'd23916, 16'd51013, 16'd42885, 16'd244, 16'd30895, 16'd57646, 16'd34457, 16'd13370, 16'd51258, 16'd41601, 16'd32626, 16'd53951, 16'd38546, 16'd52927, 16'd49256, 16'd24837, 16'd25480, 16'd60654, 16'd3882, 16'd52043, 16'd32818});
	test_expansion(128'hcda889485ad8a33216388fbc5f72fb11, {16'd24754, 16'd45047, 16'd21210, 16'd23879, 16'd16459, 16'd48037, 16'd40358, 16'd11140, 16'd59899, 16'd29030, 16'd31756, 16'd51769, 16'd34539, 16'd47947, 16'd39723, 16'd3830, 16'd20273, 16'd22105, 16'd26864, 16'd55633, 16'd5885, 16'd46608, 16'd42829, 16'd51255, 16'd36675, 16'd17552});
	test_expansion(128'h81f785ea9e1b565eb691358b15026d7b, {16'd25321, 16'd31335, 16'd65192, 16'd24502, 16'd44534, 16'd60488, 16'd49237, 16'd36591, 16'd16667, 16'd51589, 16'd57476, 16'd43132, 16'd15136, 16'd48465, 16'd36725, 16'd58569, 16'd64684, 16'd47168, 16'd26543, 16'd40324, 16'd59173, 16'd17947, 16'd3554, 16'd42748, 16'd49407, 16'd65047});
	test_expansion(128'h6c6aa6c3c82db5cc517ce96d41fa7a3e, {16'd11765, 16'd59177, 16'd61222, 16'd23114, 16'd64851, 16'd37396, 16'd58363, 16'd27757, 16'd64818, 16'd27049, 16'd29753, 16'd1351, 16'd15279, 16'd56679, 16'd40831, 16'd24801, 16'd27900, 16'd47815, 16'd36673, 16'd20448, 16'd51005, 16'd24943, 16'd19061, 16'd23578, 16'd34274, 16'd29503});
	test_expansion(128'h55d8ae3f3a6ef2710bb6142a6604aebf, {16'd37506, 16'd13414, 16'd43640, 16'd49738, 16'd55424, 16'd7095, 16'd38772, 16'd24658, 16'd33686, 16'd38540, 16'd43965, 16'd38774, 16'd34677, 16'd2741, 16'd57238, 16'd27799, 16'd33775, 16'd8380, 16'd35927, 16'd18725, 16'd35933, 16'd40765, 16'd40564, 16'd1830, 16'd42150, 16'd10268});
	test_expansion(128'hcf16ba2919e427a26a6bfe0c20d4772c, {16'd39254, 16'd5862, 16'd41447, 16'd24753, 16'd36143, 16'd22402, 16'd33520, 16'd36370, 16'd12783, 16'd17242, 16'd29572, 16'd38481, 16'd13684, 16'd5960, 16'd18701, 16'd22601, 16'd37758, 16'd33678, 16'd14444, 16'd18151, 16'd52649, 16'd25464, 16'd57702, 16'd61474, 16'd24861, 16'd29927});
	test_expansion(128'h77e7f91c5cef7338207521babffcfc34, {16'd52800, 16'd605, 16'd872, 16'd18736, 16'd59171, 16'd9943, 16'd51462, 16'd63340, 16'd14981, 16'd25841, 16'd16709, 16'd2153, 16'd54915, 16'd52735, 16'd59411, 16'd24060, 16'd3262, 16'd58589, 16'd36243, 16'd54669, 16'd30338, 16'd34312, 16'd18524, 16'd5517, 16'd44144, 16'd64230});
	test_expansion(128'hf662e320caa60a2c3d98647a9f19448a, {16'd59791, 16'd38065, 16'd11854, 16'd60124, 16'd48915, 16'd22008, 16'd31817, 16'd13299, 16'd55094, 16'd34784, 16'd44471, 16'd21479, 16'd60926, 16'd26239, 16'd55401, 16'd63010, 16'd1331, 16'd21043, 16'd63140, 16'd22391, 16'd65108, 16'd49549, 16'd8553, 16'd27159, 16'd31838, 16'd33510});
	test_expansion(128'h318d39ce026d5423d6e2f3c34688ff32, {16'd48774, 16'd31085, 16'd46925, 16'd37470, 16'd58221, 16'd55857, 16'd48497, 16'd33716, 16'd27016, 16'd14038, 16'd36695, 16'd719, 16'd10104, 16'd43982, 16'd13843, 16'd6520, 16'd46312, 16'd36507, 16'd40280, 16'd37932, 16'd60444, 16'd6665, 16'd50873, 16'd46418, 16'd50287, 16'd61455});
	test_expansion(128'h1a6c58e4fa8f03d70ae85be553a31a51, {16'd23232, 16'd58245, 16'd39833, 16'd7984, 16'd23347, 16'd23954, 16'd2075, 16'd43686, 16'd60259, 16'd37374, 16'd18598, 16'd19090, 16'd32775, 16'd64628, 16'd8346, 16'd13169, 16'd24708, 16'd58886, 16'd37918, 16'd39796, 16'd6748, 16'd2164, 16'd46411, 16'd52837, 16'd58644, 16'd38007});
	test_expansion(128'hb28165ebcdbd3a13e96a90ca75dc223e, {16'd5114, 16'd29651, 16'd12426, 16'd33153, 16'd18805, 16'd9678, 16'd64115, 16'd63062, 16'd30919, 16'd23739, 16'd8045, 16'd33454, 16'd35240, 16'd31471, 16'd999, 16'd64223, 16'd54029, 16'd37008, 16'd57755, 16'd52090, 16'd28048, 16'd41841, 16'd31941, 16'd50381, 16'd44859, 16'd40788});
	test_expansion(128'h2cf71e9a69b1e6a548c3bb212b99dc6d, {16'd42603, 16'd34157, 16'd8558, 16'd34921, 16'd2479, 16'd5593, 16'd12798, 16'd36672, 16'd22230, 16'd50377, 16'd57148, 16'd23381, 16'd36060, 16'd43845, 16'd13774, 16'd8388, 16'd734, 16'd58013, 16'd60688, 16'd2184, 16'd53813, 16'd55980, 16'd59824, 16'd25091, 16'd23000, 16'd61262});
	test_expansion(128'h3ea59e7817b93cad41b6172c084f7428, {16'd45791, 16'd47949, 16'd30005, 16'd43566, 16'd39086, 16'd36591, 16'd27729, 16'd1777, 16'd37145, 16'd24498, 16'd28023, 16'd9211, 16'd60585, 16'd15510, 16'd10725, 16'd20800, 16'd1944, 16'd36154, 16'd52131, 16'd60531, 16'd23460, 16'd43715, 16'd39008, 16'd9934, 16'd41161, 16'd6022});
	test_expansion(128'h6801eb0566e9c388cb7db81e84ae3165, {16'd12823, 16'd50813, 16'd14052, 16'd11720, 16'd47221, 16'd49380, 16'd9265, 16'd60929, 16'd25128, 16'd53842, 16'd29802, 16'd40139, 16'd54233, 16'd40007, 16'd4491, 16'd40394, 16'd26815, 16'd29055, 16'd8387, 16'd26077, 16'd49129, 16'd18916, 16'd15786, 16'd50373, 16'd63032, 16'd25612});
	test_expansion(128'h3abcb65f920345eb3a7350b721fbf5a7, {16'd34463, 16'd47907, 16'd7183, 16'd37512, 16'd30768, 16'd29155, 16'd10291, 16'd7814, 16'd14525, 16'd13657, 16'd11531, 16'd973, 16'd45426, 16'd41379, 16'd10847, 16'd35803, 16'd24806, 16'd15331, 16'd35236, 16'd17646, 16'd35283, 16'd5130, 16'd32678, 16'd48975, 16'd57645, 16'd8822});
	test_expansion(128'hfdbe8e75d0ddf5082cb084aedf19e1c6, {16'd46919, 16'd45925, 16'd46024, 16'd34335, 16'd43816, 16'd1187, 16'd48564, 16'd2124, 16'd54449, 16'd19542, 16'd3504, 16'd35993, 16'd44038, 16'd48745, 16'd33737, 16'd61357, 16'd36827, 16'd23311, 16'd24295, 16'd15468, 16'd54118, 16'd13305, 16'd52349, 16'd6536, 16'd15805, 16'd1693});
	test_expansion(128'h96cdd13512d3a5359c8fbfe092dad954, {16'd49651, 16'd38134, 16'd7506, 16'd18467, 16'd35043, 16'd6122, 16'd26857, 16'd64647, 16'd15764, 16'd63580, 16'd37027, 16'd54575, 16'd25592, 16'd17538, 16'd3075, 16'd42076, 16'd1515, 16'd46253, 16'd50313, 16'd22326, 16'd25816, 16'd50967, 16'd44369, 16'd903, 16'd3537, 16'd11725});
	test_expansion(128'hf9fa7208d36485c334e3536d0d319b63, {16'd42595, 16'd2865, 16'd35145, 16'd51963, 16'd42093, 16'd23879, 16'd32338, 16'd21495, 16'd55425, 16'd32580, 16'd3144, 16'd27923, 16'd54356, 16'd51651, 16'd33154, 16'd57988, 16'd62330, 16'd46825, 16'd18824, 16'd55128, 16'd23134, 16'd39375, 16'd15872, 16'd20585, 16'd2964, 16'd42900});
	test_expansion(128'h8cc96356c530fddaffc3755705633d9a, {16'd8363, 16'd44956, 16'd23858, 16'd51179, 16'd6075, 16'd15978, 16'd19493, 16'd55827, 16'd30819, 16'd41947, 16'd57629, 16'd43122, 16'd51405, 16'd17109, 16'd22481, 16'd4952, 16'd22929, 16'd1993, 16'd24342, 16'd55713, 16'd2321, 16'd37138, 16'd15588, 16'd1031, 16'd33753, 16'd51785});
	test_expansion(128'h589f47ba70172eb55f04457901abfc1e, {16'd22598, 16'd58259, 16'd51992, 16'd58664, 16'd61024, 16'd3183, 16'd64904, 16'd49193, 16'd7056, 16'd8469, 16'd53843, 16'd22522, 16'd22923, 16'd50880, 16'd46602, 16'd1856, 16'd36768, 16'd4134, 16'd45405, 16'd20993, 16'd3416, 16'd62165, 16'd62656, 16'd63846, 16'd25469, 16'd20017});
	test_expansion(128'hd14af0c6c7d693445bb78220452658f7, {16'd24296, 16'd64364, 16'd25709, 16'd17774, 16'd47936, 16'd50041, 16'd26447, 16'd45164, 16'd46236, 16'd27852, 16'd16342, 16'd27093, 16'd54823, 16'd61487, 16'd17000, 16'd60213, 16'd19692, 16'd9194, 16'd3467, 16'd63799, 16'd5761, 16'd41680, 16'd2033, 16'd46752, 16'd20559, 16'd4933});
	test_expansion(128'h47c5a02fb4e5299cb511a5c34c535767, {16'd41993, 16'd63570, 16'd50544, 16'd1846, 16'd42463, 16'd23116, 16'd65111, 16'd39944, 16'd2792, 16'd24642, 16'd45620, 16'd60683, 16'd19146, 16'd60892, 16'd64520, 16'd52661, 16'd32259, 16'd54899, 16'd51874, 16'd48966, 16'd17051, 16'd13548, 16'd29925, 16'd64060, 16'd59051, 16'd21619});
	test_expansion(128'h7e00debd73115f455fcb0fdfd94d5d3c, {16'd2993, 16'd29411, 16'd2275, 16'd60900, 16'd27291, 16'd54562, 16'd38979, 16'd16750, 16'd59410, 16'd11581, 16'd35156, 16'd34182, 16'd49446, 16'd38236, 16'd38373, 16'd30282, 16'd6548, 16'd47039, 16'd31227, 16'd26442, 16'd59777, 16'd21165, 16'd1599, 16'd18822, 16'd10547, 16'd58003});
	test_expansion(128'habcc54240cb902eb0e5bb0ece75d5ca4, {16'd31407, 16'd31450, 16'd37608, 16'd55143, 16'd54685, 16'd38058, 16'd11385, 16'd30010, 16'd36799, 16'd61543, 16'd7562, 16'd18648, 16'd54290, 16'd23228, 16'd45975, 16'd12830, 16'd29444, 16'd24175, 16'd17241, 16'd15294, 16'd64155, 16'd18642, 16'd55349, 16'd55128, 16'd42012, 16'd33300});
	test_expansion(128'h1bc5cb1a9ced41ed173ec21c94fb3160, {16'd16868, 16'd18216, 16'd12852, 16'd46510, 16'd49751, 16'd35459, 16'd23359, 16'd7631, 16'd745, 16'd17456, 16'd43269, 16'd56337, 16'd55086, 16'd55504, 16'd38607, 16'd42828, 16'd16234, 16'd21858, 16'd46680, 16'd44589, 16'd5687, 16'd29299, 16'd55768, 16'd6342, 16'd19530, 16'd47696});
	test_expansion(128'h4331be74e8a7db04840e6d9768709b21, {16'd29669, 16'd49962, 16'd25748, 16'd60107, 16'd25224, 16'd1070, 16'd33237, 16'd64876, 16'd511, 16'd10247, 16'd57154, 16'd19349, 16'd49108, 16'd37576, 16'd34466, 16'd28104, 16'd9696, 16'd30299, 16'd51685, 16'd5495, 16'd4663, 16'd53931, 16'd21108, 16'd44649, 16'd13568, 16'd40759});
	test_expansion(128'hc3d091e56d89b114615feead09887206, {16'd27400, 16'd40314, 16'd9272, 16'd11481, 16'd47880, 16'd18577, 16'd23372, 16'd6986, 16'd3840, 16'd41279, 16'd9470, 16'd58116, 16'd26792, 16'd52171, 16'd48076, 16'd35798, 16'd5160, 16'd42156, 16'd3287, 16'd12566, 16'd36041, 16'd9366, 16'd35130, 16'd31827, 16'd43486, 16'd58718});
	test_expansion(128'h26b76e98c3a075c097b31a06d4f83caf, {16'd49494, 16'd51929, 16'd58833, 16'd37826, 16'd14079, 16'd19015, 16'd26823, 16'd16910, 16'd9754, 16'd30424, 16'd33654, 16'd20749, 16'd41361, 16'd54478, 16'd13006, 16'd42965, 16'd25055, 16'd59888, 16'd15657, 16'd25535, 16'd4485, 16'd19847, 16'd10447, 16'd22701, 16'd63238, 16'd13281});
	test_expansion(128'h78785809063c742b3eb2b46f3dce32d5, {16'd34629, 16'd3038, 16'd5027, 16'd40321, 16'd20515, 16'd45191, 16'd48731, 16'd11242, 16'd48677, 16'd13887, 16'd2860, 16'd43917, 16'd5528, 16'd15545, 16'd63548, 16'd14862, 16'd60397, 16'd26098, 16'd20354, 16'd11057, 16'd15867, 16'd54142, 16'd18997, 16'd23776, 16'd54580, 16'd48668});
	test_expansion(128'h2c7f56faf3f61074213dab362d1ddcc3, {16'd12280, 16'd53673, 16'd8198, 16'd23111, 16'd39374, 16'd16795, 16'd46913, 16'd34017, 16'd38133, 16'd41578, 16'd58398, 16'd35286, 16'd28293, 16'd11171, 16'd43589, 16'd54348, 16'd2436, 16'd48323, 16'd20963, 16'd56631, 16'd31059, 16'd53595, 16'd33800, 16'd22502, 16'd23962, 16'd58450});
	test_expansion(128'h014acf02b028c17568e9330527b1b141, {16'd61548, 16'd16587, 16'd5796, 16'd13432, 16'd39048, 16'd53744, 16'd14351, 16'd18126, 16'd841, 16'd30905, 16'd65166, 16'd52310, 16'd7136, 16'd30803, 16'd10651, 16'd32870, 16'd42907, 16'd46677, 16'd28601, 16'd60339, 16'd46946, 16'd42799, 16'd25984, 16'd64464, 16'd1511, 16'd28855});
	test_expansion(128'h6cf828e4e6d246b0e8133954e846de62, {16'd6186, 16'd13770, 16'd22730, 16'd32694, 16'd31742, 16'd31010, 16'd33980, 16'd45119, 16'd10165, 16'd32506, 16'd46189, 16'd35316, 16'd38717, 16'd1725, 16'd24680, 16'd42618, 16'd28561, 16'd61524, 16'd30118, 16'd23895, 16'd62671, 16'd23132, 16'd30769, 16'd52287, 16'd1764, 16'd41639});
	test_expansion(128'h0dfbb40eb69e3d87204ceabf11fd70c9, {16'd42037, 16'd59497, 16'd14116, 16'd61089, 16'd26413, 16'd47437, 16'd25822, 16'd35384, 16'd10903, 16'd1024, 16'd14178, 16'd58528, 16'd33495, 16'd10892, 16'd57299, 16'd20425, 16'd63272, 16'd37039, 16'd5053, 16'd29686, 16'd45522, 16'd49984, 16'd35267, 16'd12741, 16'd46492, 16'd37381});
	test_expansion(128'hafff817cf4c598c23c9ee40a69a9ef87, {16'd3961, 16'd31859, 16'd2412, 16'd22845, 16'd57460, 16'd29877, 16'd35113, 16'd21367, 16'd34522, 16'd19596, 16'd41248, 16'd53891, 16'd59427, 16'd51144, 16'd49987, 16'd54402, 16'd32366, 16'd22418, 16'd18448, 16'd28508, 16'd28449, 16'd4866, 16'd27673, 16'd41992, 16'd22770, 16'd61591});
	test_expansion(128'he6c3240879069ca02ce5425a19cfec51, {16'd59026, 16'd28004, 16'd59698, 16'd519, 16'd32805, 16'd36265, 16'd2125, 16'd16876, 16'd49976, 16'd57843, 16'd41811, 16'd30886, 16'd46253, 16'd11173, 16'd52767, 16'd23404, 16'd44758, 16'd47111, 16'd30827, 16'd48265, 16'd31538, 16'd37565, 16'd50778, 16'd12041, 16'd27751, 16'd31122});
	test_expansion(128'hca8e919e8904e27aceb5067ab8a59ee0, {16'd42135, 16'd40594, 16'd28418, 16'd15886, 16'd32084, 16'd44507, 16'd13263, 16'd37842, 16'd2568, 16'd25910, 16'd56239, 16'd18605, 16'd46573, 16'd45179, 16'd49512, 16'd18747, 16'd6684, 16'd20997, 16'd48878, 16'd1556, 16'd40304, 16'd9714, 16'd10654, 16'd63810, 16'd27839, 16'd1885});
	test_expansion(128'h0d622096e63bea627e2c0e083d61542c, {16'd57320, 16'd19915, 16'd10072, 16'd14613, 16'd59768, 16'd64247, 16'd7074, 16'd18631, 16'd9089, 16'd25737, 16'd20839, 16'd60240, 16'd42537, 16'd35548, 16'd41241, 16'd18847, 16'd10404, 16'd10735, 16'd39179, 16'd403, 16'd39215, 16'd12313, 16'd56201, 16'd46042, 16'd54675, 16'd28512});
	test_expansion(128'h170b3fa9679e9c3ab22f5343899f8beb, {16'd46979, 16'd51867, 16'd24854, 16'd45435, 16'd53797, 16'd11649, 16'd63772, 16'd33247, 16'd7685, 16'd18694, 16'd64723, 16'd49060, 16'd32393, 16'd8417, 16'd23302, 16'd20417, 16'd57747, 16'd26500, 16'd17371, 16'd43059, 16'd48313, 16'd26516, 16'd4336, 16'd9936, 16'd41947, 16'd54629});
	test_expansion(128'h1689c543542912626add561c75aee012, {16'd20143, 16'd51506, 16'd19019, 16'd54751, 16'd4472, 16'd37669, 16'd4643, 16'd39068, 16'd12300, 16'd25060, 16'd32371, 16'd59528, 16'd30740, 16'd20065, 16'd28426, 16'd34918, 16'd22708, 16'd44095, 16'd26755, 16'd26066, 16'd20831, 16'd31406, 16'd32931, 16'd48502, 16'd7989, 16'd13194});
	test_expansion(128'h292b98489548080a9e31d3b78d3f7c3e, {16'd31347, 16'd869, 16'd5004, 16'd49672, 16'd14811, 16'd6570, 16'd48170, 16'd49519, 16'd22417, 16'd10775, 16'd39045, 16'd62656, 16'd41015, 16'd21212, 16'd59700, 16'd46278, 16'd54442, 16'd22340, 16'd55708, 16'd62350, 16'd15582, 16'd33991, 16'd32453, 16'd35000, 16'd41969, 16'd25111});
	test_expansion(128'h8f7c1101c4514c74a779f893629b0f7e, {16'd54701, 16'd16628, 16'd33343, 16'd23853, 16'd10889, 16'd52758, 16'd8581, 16'd60754, 16'd40442, 16'd19096, 16'd49271, 16'd26874, 16'd13790, 16'd58326, 16'd55436, 16'd1222, 16'd33286, 16'd31164, 16'd40983, 16'd42853, 16'd54033, 16'd52660, 16'd26582, 16'd24250, 16'd38024, 16'd16408});
	test_expansion(128'h5323600cc881f78e7e3c6b6ec4a50174, {16'd31984, 16'd47491, 16'd3103, 16'd17108, 16'd25314, 16'd14314, 16'd30656, 16'd13690, 16'd60671, 16'd55889, 16'd8348, 16'd37207, 16'd25494, 16'd12386, 16'd41858, 16'd39086, 16'd12175, 16'd60241, 16'd4115, 16'd32827, 16'd8509, 16'd35416, 16'd61767, 16'd17734, 16'd59167, 16'd45958});
	test_expansion(128'hb28521c3a8eed2c491596ab2ec9a8338, {16'd43588, 16'd61765, 16'd63860, 16'd25384, 16'd34066, 16'd50735, 16'd24756, 16'd53777, 16'd30475, 16'd50921, 16'd24352, 16'd44344, 16'd8712, 16'd38880, 16'd52743, 16'd49281, 16'd61528, 16'd32458, 16'd10462, 16'd47202, 16'd28063, 16'd22429, 16'd3769, 16'd46481, 16'd16322, 16'd20203});
	test_expansion(128'h3253360b3a8ff90fd5473572d3b04925, {16'd45605, 16'd4451, 16'd20845, 16'd25797, 16'd55178, 16'd24407, 16'd1728, 16'd50721, 16'd57011, 16'd4157, 16'd47294, 16'd25681, 16'd32850, 16'd64380, 16'd34999, 16'd18107, 16'd6717, 16'd13018, 16'd13412, 16'd45647, 16'd34447, 16'd3362, 16'd43936, 16'd53127, 16'd62263, 16'd62474});
	test_expansion(128'h9339217b1ab367bb099fd6cd23ee3ece, {16'd1466, 16'd48154, 16'd65218, 16'd25836, 16'd64872, 16'd8820, 16'd46339, 16'd58348, 16'd57515, 16'd28252, 16'd11031, 16'd52094, 16'd3281, 16'd28841, 16'd57534, 16'd63111, 16'd40883, 16'd55773, 16'd44541, 16'd859, 16'd14626, 16'd12100, 16'd20470, 16'd55632, 16'd7243, 16'd51228});
	test_expansion(128'h86d11279b07c2787e43d60433e44c7af, {16'd18001, 16'd19758, 16'd28146, 16'd33172, 16'd44633, 16'd45123, 16'd7849, 16'd41446, 16'd21162, 16'd819, 16'd65080, 16'd12566, 16'd1982, 16'd57657, 16'd21551, 16'd39842, 16'd48829, 16'd58315, 16'd45347, 16'd65022, 16'd1103, 16'd65015, 16'd33653, 16'd59189, 16'd1187, 16'd54384});
	test_expansion(128'h013628e54e1df247d0b78c39edbabb45, {16'd5021, 16'd28244, 16'd47375, 16'd39072, 16'd56568, 16'd53669, 16'd38265, 16'd28359, 16'd15851, 16'd40538, 16'd1411, 16'd56566, 16'd35181, 16'd47211, 16'd63655, 16'd54248, 16'd1988, 16'd51979, 16'd48919, 16'd61861, 16'd5745, 16'd31247, 16'd63490, 16'd34964, 16'd10453, 16'd44268});
	test_expansion(128'h377a517ee538a5f4f17c7fac90623ec1, {16'd5427, 16'd44163, 16'd31385, 16'd58085, 16'd60327, 16'd64714, 16'd10135, 16'd30473, 16'd55576, 16'd18181, 16'd22957, 16'd28199, 16'd24254, 16'd41871, 16'd37114, 16'd32880, 16'd62242, 16'd34322, 16'd36988, 16'd29482, 16'd9770, 16'd57059, 16'd26124, 16'd53229, 16'd3222, 16'd25359});
	test_expansion(128'hf409e812763fe461e3480ae974a97f21, {16'd39651, 16'd63837, 16'd6352, 16'd64283, 16'd46024, 16'd17031, 16'd39090, 16'd12615, 16'd14283, 16'd9349, 16'd20838, 16'd36163, 16'd9251, 16'd26625, 16'd4944, 16'd25169, 16'd62759, 16'd62780, 16'd3296, 16'd20247, 16'd4953, 16'd62296, 16'd62357, 16'd54877, 16'd29456, 16'd38981});
	test_expansion(128'hda653da909285070b6859d9d29a60d80, {16'd33892, 16'd15597, 16'd10776, 16'd59266, 16'd25777, 16'd24392, 16'd36894, 16'd16149, 16'd3401, 16'd59757, 16'd29413, 16'd2150, 16'd53605, 16'd13575, 16'd47452, 16'd45974, 16'd55943, 16'd31982, 16'd2179, 16'd20405, 16'd1211, 16'd12710, 16'd1864, 16'd19552, 16'd17628, 16'd35231});
	test_expansion(128'h8e7a706f855aea2047decf684548b798, {16'd10441, 16'd50822, 16'd16635, 16'd62071, 16'd10618, 16'd24469, 16'd1345, 16'd16880, 16'd36693, 16'd30753, 16'd26460, 16'd13209, 16'd60813, 16'd9658, 16'd62808, 16'd58699, 16'd15222, 16'd41647, 16'd43350, 16'd52034, 16'd49237, 16'd35173, 16'd59588, 16'd35672, 16'd32731, 16'd2709});
	test_expansion(128'h7b6638fdd8124ec6049ab098e0d39f4a, {16'd10379, 16'd14696, 16'd58508, 16'd57068, 16'd56241, 16'd13748, 16'd59282, 16'd5097, 16'd26682, 16'd16646, 16'd25472, 16'd45765, 16'd63870, 16'd29654, 16'd14259, 16'd18848, 16'd33105, 16'd32718, 16'd20035, 16'd29994, 16'd62792, 16'd43407, 16'd19429, 16'd51936, 16'd4723, 16'd45509});
	test_expansion(128'h512bcb38b6025d1aa2c4e74bb8e20d2e, {16'd37839, 16'd12983, 16'd39931, 16'd36431, 16'd25619, 16'd20983, 16'd45602, 16'd32643, 16'd2812, 16'd39241, 16'd54796, 16'd54992, 16'd27199, 16'd16540, 16'd11984, 16'd33970, 16'd29892, 16'd6023, 16'd9437, 16'd61929, 16'd45183, 16'd26466, 16'd31, 16'd22326, 16'd43833, 16'd6021});
	test_expansion(128'h9a2003cf7f30ae4ef6d611bcc765602b, {16'd7693, 16'd64486, 16'd44326, 16'd61039, 16'd36105, 16'd44515, 16'd31604, 16'd29369, 16'd32799, 16'd58147, 16'd35904, 16'd44698, 16'd1638, 16'd24416, 16'd10132, 16'd38288, 16'd22124, 16'd54163, 16'd62867, 16'd10550, 16'd65036, 16'd4057, 16'd3090, 16'd12558, 16'd32148, 16'd64665});
	test_expansion(128'h7462cf74bc3b40bd53d4368998d77038, {16'd4089, 16'd25406, 16'd8136, 16'd22235, 16'd210, 16'd55038, 16'd58455, 16'd54862, 16'd463, 16'd62572, 16'd39782, 16'd62527, 16'd45417, 16'd39375, 16'd6604, 16'd12222, 16'd6233, 16'd56276, 16'd39229, 16'd23696, 16'd29324, 16'd39270, 16'd45761, 16'd49531, 16'd4261, 16'd24392});
	test_expansion(128'ha3e490a46176a955a4db96e296417483, {16'd5956, 16'd25376, 16'd35428, 16'd11925, 16'd41634, 16'd5458, 16'd30428, 16'd30334, 16'd44981, 16'd64355, 16'd48193, 16'd58899, 16'd50443, 16'd6446, 16'd36837, 16'd31748, 16'd58498, 16'd64317, 16'd51753, 16'd60447, 16'd36353, 16'd9677, 16'd48405, 16'd64571, 16'd32508, 16'd57396});
	test_expansion(128'h27518d4d1d24adee110dcfe7792f2ca6, {16'd45793, 16'd33795, 16'd21427, 16'd6414, 16'd16592, 16'd36683, 16'd54873, 16'd51002, 16'd13440, 16'd55898, 16'd44196, 16'd51833, 16'd39075, 16'd50987, 16'd24844, 16'd45237, 16'd21364, 16'd51085, 16'd34902, 16'd61412, 16'd40873, 16'd4307, 16'd9566, 16'd17140, 16'd44549, 16'd43726});
	test_expansion(128'h9c6480c717c1cdfadd26f104a13113ba, {16'd50356, 16'd11636, 16'd1345, 16'd56481, 16'd5366, 16'd15636, 16'd33308, 16'd13548, 16'd55518, 16'd39870, 16'd43961, 16'd34288, 16'd51725, 16'd20717, 16'd59001, 16'd27573, 16'd33635, 16'd15967, 16'd36907, 16'd26377, 16'd37071, 16'd30836, 16'd41921, 16'd35475, 16'd39353, 16'd16726});
	test_expansion(128'h6dfa98cb53717149c2aa7eb70df8a27d, {16'd27826, 16'd62844, 16'd51566, 16'd31310, 16'd9485, 16'd14610, 16'd44885, 16'd56958, 16'd25113, 16'd56991, 16'd31913, 16'd24904, 16'd21085, 16'd12810, 16'd10815, 16'd11552, 16'd64637, 16'd21396, 16'd64260, 16'd51604, 16'd32035, 16'd22741, 16'd17324, 16'd43383, 16'd55660, 16'd47005});
	test_expansion(128'h56a2bd20a837ca1c813d5f46619502c4, {16'd23458, 16'd36559, 16'd4051, 16'd20891, 16'd36834, 16'd62623, 16'd62001, 16'd24856, 16'd7749, 16'd23980, 16'd16028, 16'd51879, 16'd53568, 16'd14262, 16'd26634, 16'd25407, 16'd54995, 16'd12173, 16'd27706, 16'd23972, 16'd5421, 16'd61704, 16'd60006, 16'd40847, 16'd53699, 16'd35332});
	test_expansion(128'h22b20573de451cfcf549c0c744745f0e, {16'd16000, 16'd61400, 16'd18401, 16'd13584, 16'd13392, 16'd7123, 16'd57347, 16'd39329, 16'd32299, 16'd12057, 16'd35321, 16'd2339, 16'd3272, 16'd8544, 16'd9120, 16'd53384, 16'd45745, 16'd35712, 16'd4266, 16'd20515, 16'd12828, 16'd34601, 16'd35706, 16'd61164, 16'd45718, 16'd29425});
	test_expansion(128'hca82b09d9e00727438e7b3ab2b6902d9, {16'd54979, 16'd14939, 16'd45079, 16'd60258, 16'd48862, 16'd41865, 16'd30599, 16'd45155, 16'd21622, 16'd42416, 16'd62788, 16'd2790, 16'd42471, 16'd39235, 16'd2635, 16'd50665, 16'd61348, 16'd49012, 16'd6150, 16'd36244, 16'd48138, 16'd50954, 16'd828, 16'd27456, 16'd41795, 16'd39488});
	test_expansion(128'h7cd7f11b6ebec227ceb176bd7bd02048, {16'd34108, 16'd13953, 16'd27260, 16'd36354, 16'd42125, 16'd53518, 16'd26122, 16'd26981, 16'd38029, 16'd12353, 16'd35412, 16'd31889, 16'd63713, 16'd1873, 16'd27295, 16'd1885, 16'd33052, 16'd45313, 16'd35984, 16'd33750, 16'd59437, 16'd64317, 16'd23418, 16'd40019, 16'd59176, 16'd4205});
	test_expansion(128'ha1b54b2f9d46b06f82a657af35813e42, {16'd42270, 16'd43400, 16'd44978, 16'd28967, 16'd33642, 16'd5537, 16'd33724, 16'd41213, 16'd44791, 16'd17107, 16'd23742, 16'd12223, 16'd52029, 16'd17948, 16'd1172, 16'd34532, 16'd32455, 16'd20934, 16'd60167, 16'd18317, 16'd23777, 16'd22280, 16'd43832, 16'd263, 16'd8445, 16'd61754});
	test_expansion(128'hd8208a33219b0204058657067ab7ff76, {16'd28310, 16'd53841, 16'd9977, 16'd38199, 16'd32177, 16'd45203, 16'd57119, 16'd3541, 16'd57912, 16'd61229, 16'd46399, 16'd15646, 16'd7722, 16'd49740, 16'd51312, 16'd40818, 16'd55252, 16'd53511, 16'd60270, 16'd14522, 16'd42182, 16'd768, 16'd9043, 16'd6650, 16'd17082, 16'd44829});
	test_expansion(128'h9f86f474afa8635f91212b653ad1a3c6, {16'd15064, 16'd33482, 16'd6578, 16'd39502, 16'd32390, 16'd38108, 16'd22583, 16'd4242, 16'd16667, 16'd42919, 16'd31001, 16'd30252, 16'd57113, 16'd61313, 16'd60062, 16'd9489, 16'd13964, 16'd39796, 16'd49961, 16'd14420, 16'd36675, 16'd39735, 16'd28157, 16'd36480, 16'd21567, 16'd62341});
	test_expansion(128'h671b53d7b8e0d763acba23dd1da2196e, {16'd62516, 16'd37228, 16'd14207, 16'd8297, 16'd57480, 16'd65421, 16'd13257, 16'd24921, 16'd5642, 16'd50191, 16'd8118, 16'd23011, 16'd57120, 16'd39494, 16'd17386, 16'd9772, 16'd39885, 16'd61101, 16'd24210, 16'd25635, 16'd60094, 16'd62135, 16'd25180, 16'd2112, 16'd36722, 16'd57934});
	test_expansion(128'h4ff04db6bf53a947d222ae00a1a2acf6, {16'd6760, 16'd63378, 16'd64990, 16'd43992, 16'd40462, 16'd30578, 16'd31055, 16'd8570, 16'd14819, 16'd52493, 16'd24332, 16'd19893, 16'd49718, 16'd21254, 16'd55638, 16'd51996, 16'd7802, 16'd48590, 16'd11126, 16'd31425, 16'd20153, 16'd39468, 16'd17637, 16'd27917, 16'd41343, 16'd59835});
	test_expansion(128'h46559ae3ae9b7ccf09af796c75c1f7a4, {16'd24681, 16'd34036, 16'd11105, 16'd63828, 16'd51304, 16'd3628, 16'd17114, 16'd50863, 16'd30265, 16'd20989, 16'd20585, 16'd43210, 16'd26614, 16'd15160, 16'd2301, 16'd25772, 16'd9041, 16'd29652, 16'd37743, 16'd42005, 16'd4555, 16'd10599, 16'd42716, 16'd47434, 16'd19071, 16'd63490});
	test_expansion(128'ha3d179a6e152652ecdcc6b5b3070a93a, {16'd51729, 16'd53707, 16'd65361, 16'd33775, 16'd52191, 16'd28348, 16'd8107, 16'd22468, 16'd27290, 16'd64846, 16'd57242, 16'd6457, 16'd7471, 16'd30344, 16'd37026, 16'd19413, 16'd30775, 16'd23654, 16'd64403, 16'd56245, 16'd19191, 16'd54561, 16'd56655, 16'd60239, 16'd59286, 16'd6282});
	test_expansion(128'h72a6e532f87a937b5a0f8ccb7b9f6833, {16'd25955, 16'd10193, 16'd13824, 16'd58209, 16'd54318, 16'd44811, 16'd44193, 16'd46704, 16'd52420, 16'd36844, 16'd49775, 16'd46932, 16'd63228, 16'd10393, 16'd11685, 16'd21951, 16'd36930, 16'd40824, 16'd50634, 16'd30739, 16'd23537, 16'd51736, 16'd17607, 16'd33949, 16'd46052, 16'd45577});
	test_expansion(128'h4a2c3aba5083d08cdd26d0a6c5ecc603, {16'd46390, 16'd60986, 16'd29549, 16'd17282, 16'd15172, 16'd1100, 16'd29722, 16'd24765, 16'd32198, 16'd51182, 16'd20188, 16'd43653, 16'd3280, 16'd8973, 16'd43072, 16'd906, 16'd32874, 16'd20163, 16'd43297, 16'd41542, 16'd45164, 16'd27029, 16'd65514, 16'd11471, 16'd25941, 16'd9712});
	test_expansion(128'h062b195b22df322a6568db884dcbb348, {16'd40296, 16'd63864, 16'd7348, 16'd5746, 16'd25489, 16'd24740, 16'd42224, 16'd24945, 16'd57379, 16'd17588, 16'd14659, 16'd58385, 16'd1565, 16'd40127, 16'd22449, 16'd39677, 16'd19899, 16'd47391, 16'd23988, 16'd43860, 16'd35289, 16'd47685, 16'd19396, 16'd25004, 16'd33587, 16'd26550});
	test_expansion(128'h32d86067ef57220550fdcd99393db341, {16'd49218, 16'd35135, 16'd26977, 16'd14392, 16'd37255, 16'd54211, 16'd15924, 16'd49917, 16'd48673, 16'd65303, 16'd50029, 16'd3288, 16'd58025, 16'd17686, 16'd39797, 16'd17364, 16'd2651, 16'd13272, 16'd9652, 16'd21474, 16'd18822, 16'd31453, 16'd49966, 16'd33162, 16'd32844, 16'd56712});
	test_expansion(128'h07ef049201b2c905448f1d5e26fd341a, {16'd33369, 16'd16983, 16'd44516, 16'd48264, 16'd19543, 16'd55409, 16'd26674, 16'd35168, 16'd8129, 16'd43387, 16'd61971, 16'd5422, 16'd22925, 16'd47599, 16'd9563, 16'd62970, 16'd47009, 16'd20177, 16'd58954, 16'd44546, 16'd50443, 16'd45776, 16'd41956, 16'd55517, 16'd59329, 16'd15970});
	test_expansion(128'h7bf9d35f6634f14c9488f7753b4d67b0, {16'd1350, 16'd25494, 16'd39389, 16'd5564, 16'd21828, 16'd7286, 16'd46646, 16'd35247, 16'd64270, 16'd33579, 16'd15047, 16'd41774, 16'd5714, 16'd62161, 16'd37632, 16'd4394, 16'd23573, 16'd27973, 16'd19162, 16'd44532, 16'd61450, 16'd16633, 16'd9847, 16'd29235, 16'd34903, 16'd38670});
	test_expansion(128'h9dd98b2ed7eb5ef317cb5dbff99bcfd9, {16'd25513, 16'd38892, 16'd6000, 16'd29912, 16'd24233, 16'd17175, 16'd59722, 16'd42630, 16'd30773, 16'd16933, 16'd39110, 16'd2820, 16'd3817, 16'd1368, 16'd18743, 16'd53640, 16'd8275, 16'd19353, 16'd33205, 16'd28218, 16'd41719, 16'd40751, 16'd13984, 16'd16088, 16'd22638, 16'd23172});
	test_expansion(128'h11e6af822c2f6d4618c5ee7ee5155dce, {16'd8167, 16'd10815, 16'd35605, 16'd27222, 16'd3938, 16'd4078, 16'd4066, 16'd30013, 16'd7504, 16'd15612, 16'd50309, 16'd34997, 16'd24101, 16'd5058, 16'd21372, 16'd17744, 16'd51668, 16'd32904, 16'd65034, 16'd40051, 16'd20602, 16'd33189, 16'd56346, 16'd56553, 16'd41503, 16'd16694});
	test_expansion(128'hd581aec23a6595830a1438954f5e20a5, {16'd58884, 16'd23010, 16'd16463, 16'd35572, 16'd16670, 16'd13713, 16'd19372, 16'd7934, 16'd51151, 16'd26215, 16'd38892, 16'd31815, 16'd2146, 16'd37861, 16'd39396, 16'd42072, 16'd38303, 16'd48229, 16'd33850, 16'd12855, 16'd57988, 16'd21194, 16'd16946, 16'd44101, 16'd41223, 16'd26255});
	test_expansion(128'h576108cd9954e2a9dd781b40ce5206fe, {16'd46769, 16'd59483, 16'd53987, 16'd62820, 16'd6954, 16'd40849, 16'd31207, 16'd19384, 16'd2445, 16'd41336, 16'd38255, 16'd34214, 16'd1679, 16'd42967, 16'd33435, 16'd43776, 16'd25056, 16'd15928, 16'd9423, 16'd63827, 16'd2379, 16'd37929, 16'd30651, 16'd51771, 16'd24424, 16'd33377});
	test_expansion(128'hbf74fc3f345157eb4f2b56fdf2e6d862, {16'd19221, 16'd53706, 16'd37837, 16'd35498, 16'd6005, 16'd53842, 16'd56418, 16'd16311, 16'd58111, 16'd2450, 16'd54680, 16'd5538, 16'd54593, 16'd7357, 16'd38930, 16'd34574, 16'd61593, 16'd58498, 16'd12509, 16'd14645, 16'd54253, 16'd50065, 16'd46313, 16'd48712, 16'd20009, 16'd22351});
	test_expansion(128'h5c8ba87b0aec7e8850537e739f7b294a, {16'd13302, 16'd20645, 16'd13903, 16'd11546, 16'd27696, 16'd31492, 16'd48800, 16'd24609, 16'd13953, 16'd55174, 16'd61, 16'd61513, 16'd45498, 16'd783, 16'd20773, 16'd53909, 16'd27301, 16'd10793, 16'd64221, 16'd63282, 16'd47763, 16'd64550, 16'd24298, 16'd40836, 16'd27675, 16'd40763});
	test_expansion(128'hbae0395d91740cc3b87075b59deded4a, {16'd42686, 16'd28844, 16'd3080, 16'd1720, 16'd63677, 16'd54442, 16'd60273, 16'd22609, 16'd62867, 16'd50129, 16'd22409, 16'd31433, 16'd6914, 16'd59478, 16'd56246, 16'd11837, 16'd40464, 16'd64062, 16'd24703, 16'd37061, 16'd60425, 16'd832, 16'd36025, 16'd57910, 16'd23000, 16'd29085});
	test_expansion(128'h79fa6611f3f54cdfdb03eb9d4750cb49, {16'd23182, 16'd53688, 16'd11357, 16'd41045, 16'd54878, 16'd63071, 16'd61349, 16'd56537, 16'd9328, 16'd58721, 16'd51071, 16'd64790, 16'd17138, 16'd29512, 16'd11253, 16'd50725, 16'd31341, 16'd63175, 16'd15668, 16'd17511, 16'd19404, 16'd64966, 16'd9371, 16'd40762, 16'd59154, 16'd12495});
	test_expansion(128'ha01e93ac4f47eb33d643916d16514175, {16'd49274, 16'd24613, 16'd56612, 16'd58056, 16'd23021, 16'd4013, 16'd59077, 16'd56997, 16'd25543, 16'd1955, 16'd53932, 16'd43127, 16'd33354, 16'd4764, 16'd60742, 16'd31614, 16'd2752, 16'd60565, 16'd42485, 16'd53756, 16'd28546, 16'd14348, 16'd39477, 16'd42403, 16'd49346, 16'd52292});
	test_expansion(128'h47fbd9d705c98c479100474c9d60bc1d, {16'd29712, 16'd1946, 16'd55416, 16'd38195, 16'd51, 16'd59230, 16'd33217, 16'd54882, 16'd55349, 16'd57278, 16'd17912, 16'd4576, 16'd26397, 16'd792, 16'd53075, 16'd44554, 16'd16399, 16'd21509, 16'd18093, 16'd49495, 16'd36368, 16'd21402, 16'd16510, 16'd64274, 16'd48702, 16'd13970});
	test_expansion(128'hb80f85c8204ed03c10bd5f11a8b257e0, {16'd4379, 16'd12756, 16'd61437, 16'd29477, 16'd38424, 16'd60204, 16'd47222, 16'd21153, 16'd14807, 16'd10075, 16'd31998, 16'd29264, 16'd33339, 16'd4418, 16'd59725, 16'd9338, 16'd56002, 16'd54067, 16'd8523, 16'd18912, 16'd43481, 16'd27790, 16'd63640, 16'd20600, 16'd55861, 16'd27480});
	test_expansion(128'h984890941a42d6821c0f39281fc2da6a, {16'd62135, 16'd40746, 16'd7501, 16'd18540, 16'd48960, 16'd64626, 16'd55112, 16'd22138, 16'd2316, 16'd4190, 16'd8214, 16'd34815, 16'd30419, 16'd38701, 16'd5369, 16'd14248, 16'd7198, 16'd27833, 16'd12046, 16'd38843, 16'd19578, 16'd23424, 16'd47975, 16'd2987, 16'd18823, 16'd5991});
	test_expansion(128'h645f9f50165b761c30b4f253e0c2bb9b, {16'd52635, 16'd57594, 16'd8224, 16'd62094, 16'd62683, 16'd20182, 16'd701, 16'd44180, 16'd33106, 16'd11766, 16'd20882, 16'd54021, 16'd57144, 16'd17648, 16'd47813, 16'd28661, 16'd23102, 16'd23265, 16'd56092, 16'd17726, 16'd60228, 16'd15063, 16'd41243, 16'd37400, 16'd19613, 16'd64351});
	test_expansion(128'h1921d62ebdfb9ef37cebda0891c8ec3e, {16'd15493, 16'd49021, 16'd19524, 16'd20239, 16'd38043, 16'd42337, 16'd1224, 16'd41433, 16'd65382, 16'd60192, 16'd17921, 16'd49802, 16'd55753, 16'd5214, 16'd58575, 16'd28816, 16'd34771, 16'd53040, 16'd14111, 16'd8206, 16'd62035, 16'd1768, 16'd378, 16'd4530, 16'd8139, 16'd6443});
	test_expansion(128'hadb0ff7995702e6479c3bc5a99473bb9, {16'd46152, 16'd57812, 16'd17761, 16'd27334, 16'd33764, 16'd15433, 16'd15003, 16'd51891, 16'd5729, 16'd18517, 16'd17769, 16'd47635, 16'd62403, 16'd38102, 16'd8417, 16'd9117, 16'd25572, 16'd16124, 16'd31267, 16'd58683, 16'd1309, 16'd10524, 16'd18719, 16'd65128, 16'd17601, 16'd51898});
	test_expansion(128'hac581db6851972301420c66b4324998a, {16'd18860, 16'd9663, 16'd50157, 16'd9950, 16'd17064, 16'd25091, 16'd48339, 16'd6655, 16'd47971, 16'd65175, 16'd7066, 16'd262, 16'd9565, 16'd32727, 16'd27631, 16'd29584, 16'd37024, 16'd8463, 16'd36163, 16'd4809, 16'd34697, 16'd46695, 16'd41685, 16'd33068, 16'd89, 16'd7367});
	test_expansion(128'hb8991986bcb22d79f39eea9dc01cac81, {16'd44560, 16'd19780, 16'd49722, 16'd11642, 16'd31224, 16'd26629, 16'd40230, 16'd31816, 16'd63636, 16'd47708, 16'd28439, 16'd61266, 16'd56384, 16'd48498, 16'd18406, 16'd17202, 16'd14332, 16'd60496, 16'd45112, 16'd44022, 16'd54784, 16'd19922, 16'd52141, 16'd61446, 16'd33617, 16'd42769});
	test_expansion(128'hc27093fc4b49a6180974fe59701e3651, {16'd63952, 16'd12856, 16'd30003, 16'd51218, 16'd30418, 16'd26203, 16'd60924, 16'd2177, 16'd11128, 16'd51564, 16'd19756, 16'd61943, 16'd25707, 16'd9631, 16'd9100, 16'd27816, 16'd2999, 16'd59719, 16'd42226, 16'd31881, 16'd33963, 16'd17675, 16'd49001, 16'd21330, 16'd57420, 16'd38738});
	test_expansion(128'h5da9a3d0dff9909ffa1014d66d0cd4db, {16'd55757, 16'd17903, 16'd65209, 16'd62251, 16'd43719, 16'd41626, 16'd12264, 16'd58771, 16'd52408, 16'd59779, 16'd19542, 16'd3268, 16'd8202, 16'd18464, 16'd21417, 16'd38150, 16'd63724, 16'd1975, 16'd63748, 16'd23381, 16'd18031, 16'd3143, 16'd33240, 16'd62907, 16'd37466, 16'd50239});
	test_expansion(128'h84609d9b975cc7c88241fff8dcca7cd0, {16'd20138, 16'd51751, 16'd28071, 16'd24768, 16'd38111, 16'd39087, 16'd467, 16'd62988, 16'd38767, 16'd3679, 16'd10459, 16'd36454, 16'd4261, 16'd13521, 16'd34953, 16'd44826, 16'd13510, 16'd56174, 16'd53325, 16'd24212, 16'd11248, 16'd30701, 16'd6081, 16'd7659, 16'd10439, 16'd64391});
	test_expansion(128'hbb857c2b6264b7f93cc6e9f9ea52496d, {16'd59372, 16'd20037, 16'd25493, 16'd7611, 16'd63899, 16'd39079, 16'd15248, 16'd24301, 16'd38107, 16'd19472, 16'd60347, 16'd31631, 16'd18033, 16'd7216, 16'd8224, 16'd43660, 16'd44142, 16'd36656, 16'd52151, 16'd32190, 16'd59770, 16'd3689, 16'd43286, 16'd18259, 16'd59812, 16'd48457});
	test_expansion(128'h6b8f9909d9d913a88182230e1ff86b37, {16'd6356, 16'd21801, 16'd62485, 16'd2110, 16'd43263, 16'd7566, 16'd2519, 16'd50126, 16'd49696, 16'd10215, 16'd54511, 16'd38346, 16'd12376, 16'd26609, 16'd33481, 16'd20887, 16'd5157, 16'd60153, 16'd43712, 16'd4715, 16'd26041, 16'd42701, 16'd11753, 16'd38905, 16'd54416, 16'd35059});
	test_expansion(128'h909a9f94b7fb13388e3187c0e7ce5af2, {16'd5217, 16'd64128, 16'd39947, 16'd36716, 16'd12790, 16'd163, 16'd11200, 16'd9829, 16'd30998, 16'd41282, 16'd30089, 16'd5965, 16'd23561, 16'd623, 16'd21475, 16'd5570, 16'd60617, 16'd33238, 16'd13482, 16'd18284, 16'd44309, 16'd18770, 16'd15946, 16'd51206, 16'd4024, 16'd26494});
	test_expansion(128'hf760cc4ec755b8834092d98409bded97, {16'd3518, 16'd62902, 16'd30003, 16'd5558, 16'd41975, 16'd2350, 16'd21092, 16'd24977, 16'd25538, 16'd44927, 16'd32368, 16'd61549, 16'd57538, 16'd16057, 16'd40726, 16'd7007, 16'd2952, 16'd7445, 16'd1286, 16'd33653, 16'd8355, 16'd33594, 16'd29902, 16'd63032, 16'd58362, 16'd34200});
	test_expansion(128'h700d0016ad77ed800a41e6619a5bc8ed, {16'd65094, 16'd40595, 16'd5854, 16'd34827, 16'd9240, 16'd23985, 16'd39953, 16'd19938, 16'd16141, 16'd63224, 16'd24015, 16'd30990, 16'd39046, 16'd45823, 16'd23249, 16'd13462, 16'd46643, 16'd30792, 16'd13089, 16'd10554, 16'd26584, 16'd41883, 16'd27272, 16'd351, 16'd55418, 16'd51168});
	test_expansion(128'hd9557ff0f339fcef89c7a6f0baed40fe, {16'd16292, 16'd12006, 16'd60546, 16'd39566, 16'd32791, 16'd47304, 16'd24592, 16'd5077, 16'd4859, 16'd29162, 16'd53688, 16'd55096, 16'd8137, 16'd4675, 16'd4776, 16'd5831, 16'd25411, 16'd42333, 16'd46818, 16'd60383, 16'd14681, 16'd26992, 16'd51645, 16'd4879, 16'd10591, 16'd15540});
	test_expansion(128'h98036e4078237a78cce48975503f5e97, {16'd1357, 16'd46781, 16'd21606, 16'd55074, 16'd51875, 16'd48840, 16'd48743, 16'd40018, 16'd15210, 16'd36005, 16'd25674, 16'd26006, 16'd15534, 16'd8443, 16'd47563, 16'd58217, 16'd18510, 16'd25206, 16'd63822, 16'd15728, 16'd60117, 16'd40901, 16'd6011, 16'd32165, 16'd11778, 16'd2785});
	test_expansion(128'he744b613cae14425703042391dd86d2f, {16'd53115, 16'd13080, 16'd16072, 16'd24098, 16'd45437, 16'd30239, 16'd53271, 16'd23818, 16'd16101, 16'd28893, 16'd10034, 16'd21735, 16'd46705, 16'd20223, 16'd25940, 16'd32578, 16'd47599, 16'd14244, 16'd5372, 16'd20454, 16'd30854, 16'd57123, 16'd25482, 16'd46197, 16'd27053, 16'd12103});
	test_expansion(128'hec623c0d2aaf32a7b85a32067bb32f49, {16'd154, 16'd42096, 16'd19769, 16'd53073, 16'd62827, 16'd60064, 16'd23133, 16'd2454, 16'd50446, 16'd37124, 16'd35791, 16'd39481, 16'd28663, 16'd14347, 16'd12432, 16'd33778, 16'd58371, 16'd16655, 16'd36085, 16'd56310, 16'd27088, 16'd63925, 16'd65339, 16'd29868, 16'd11119, 16'd19432});
	test_expansion(128'h44b0b7027df25870f360c9820879da7a, {16'd55048, 16'd53499, 16'd2747, 16'd13642, 16'd14174, 16'd2363, 16'd295, 16'd9433, 16'd37193, 16'd42612, 16'd12259, 16'd16278, 16'd3398, 16'd44136, 16'd46183, 16'd62849, 16'd47430, 16'd51024, 16'd45894, 16'd25080, 16'd15927, 16'd15594, 16'd19250, 16'd2437, 16'd62678, 16'd45889});
	test_expansion(128'h9f9be13071699d0f6816cebf0975aabc, {16'd9676, 16'd12421, 16'd3395, 16'd51178, 16'd49837, 16'd11072, 16'd40909, 16'd35334, 16'd26241, 16'd59013, 16'd31361, 16'd59030, 16'd52426, 16'd5806, 16'd42238, 16'd34287, 16'd50071, 16'd45307, 16'd9149, 16'd33633, 16'd28586, 16'd26847, 16'd41979, 16'd33135, 16'd30111, 16'd53677});
	test_expansion(128'hae24da2495fc09b48c1db2cdf0dc81f7, {16'd1723, 16'd37791, 16'd9191, 16'd28199, 16'd51696, 16'd22158, 16'd34988, 16'd61643, 16'd2597, 16'd481, 16'd51341, 16'd18379, 16'd30862, 16'd33312, 16'd19793, 16'd24304, 16'd24205, 16'd8107, 16'd59579, 16'd60063, 16'd7675, 16'd1529, 16'd50577, 16'd23650, 16'd44502, 16'd65481});
	test_expansion(128'h0a9d1f33529d3dafe8e9a82257ff3aab, {16'd19688, 16'd60, 16'd42844, 16'd4235, 16'd59652, 16'd61442, 16'd39841, 16'd46758, 16'd31082, 16'd38614, 16'd29249, 16'd35773, 16'd31057, 16'd9318, 16'd16136, 16'd33402, 16'd14716, 16'd6205, 16'd42005, 16'd60103, 16'd27695, 16'd39490, 16'd59415, 16'd40921, 16'd26449, 16'd1377});
	test_expansion(128'hec904964de2135ae9bf5d512983813f5, {16'd40432, 16'd26640, 16'd38612, 16'd19177, 16'd52817, 16'd58401, 16'd25089, 16'd48492, 16'd28417, 16'd2908, 16'd21203, 16'd28965, 16'd30831, 16'd15674, 16'd55084, 16'd50924, 16'd27003, 16'd24477, 16'd4505, 16'd37496, 16'd39126, 16'd34771, 16'd48938, 16'd61927, 16'd1364, 16'd11296});
	test_expansion(128'h2703e22bd16c7e245ab98d471a1c520c, {16'd12514, 16'd56151, 16'd45340, 16'd19733, 16'd36885, 16'd57049, 16'd373, 16'd34421, 16'd30347, 16'd46391, 16'd11202, 16'd4134, 16'd12097, 16'd62726, 16'd42298, 16'd53667, 16'd39997, 16'd18855, 16'd9778, 16'd49163, 16'd32159, 16'd10927, 16'd50364, 16'd12626, 16'd53936, 16'd28765});
	test_expansion(128'h051a07d4d2ad6831a2c1ed18631f8032, {16'd35515, 16'd19437, 16'd56643, 16'd63784, 16'd26153, 16'd33878, 16'd63244, 16'd21171, 16'd6049, 16'd62667, 16'd59171, 16'd31266, 16'd43500, 16'd50860, 16'd15479, 16'd977, 16'd9477, 16'd52186, 16'd15675, 16'd20438, 16'd59885, 16'd24378, 16'd11076, 16'd57286, 16'd50028, 16'd64814});
	test_expansion(128'h1f1f6c755cd54fead13420e6f72a8bed, {16'd38402, 16'd28176, 16'd64810, 16'd59016, 16'd33061, 16'd27245, 16'd3099, 16'd44304, 16'd55987, 16'd61024, 16'd8890, 16'd50081, 16'd30503, 16'd2760, 16'd15450, 16'd31240, 16'd35590, 16'd50040, 16'd2003, 16'd14557, 16'd59744, 16'd20797, 16'd638, 16'd29926, 16'd41567, 16'd34135});
	test_expansion(128'h53deed58484210d07a38e5107129723b, {16'd33205, 16'd35596, 16'd57590, 16'd56529, 16'd50529, 16'd13248, 16'd53092, 16'd46093, 16'd6834, 16'd30441, 16'd54890, 16'd49642, 16'd11304, 16'd41410, 16'd6987, 16'd4484, 16'd14546, 16'd61400, 16'd45501, 16'd60043, 16'd51976, 16'd5312, 16'd40163, 16'd5893, 16'd51104, 16'd17969});
	test_expansion(128'h37d7e6120b3f363965f9faf7925bfc68, {16'd50175, 16'd25707, 16'd44791, 16'd54337, 16'd22070, 16'd60490, 16'd21622, 16'd6356, 16'd30982, 16'd38060, 16'd54013, 16'd34188, 16'd16242, 16'd55719, 16'd43624, 16'd62819, 16'd44561, 16'd46057, 16'd14532, 16'd11132, 16'd15089, 16'd25238, 16'd7811, 16'd26801, 16'd43096, 16'd30006});
	test_expansion(128'h2ddbc0ac7b8a1c7aa61c04cba496bee3, {16'd25711, 16'd7837, 16'd61488, 16'd49405, 16'd13553, 16'd51514, 16'd58493, 16'd62383, 16'd33069, 16'd54688, 16'd54117, 16'd56943, 16'd29681, 16'd35778, 16'd15614, 16'd20926, 16'd23242, 16'd48686, 16'd28526, 16'd7152, 16'd32000, 16'd15436, 16'd17096, 16'd36665, 16'd24632, 16'd39351});
	test_expansion(128'h741a833b648232698fe13324172a1460, {16'd29471, 16'd16775, 16'd6418, 16'd62242, 16'd14839, 16'd2593, 16'd26572, 16'd54036, 16'd55409, 16'd50853, 16'd30199, 16'd27116, 16'd43578, 16'd18751, 16'd16934, 16'd22760, 16'd28558, 16'd26528, 16'd12056, 16'd61435, 16'd3957, 16'd64340, 16'd48416, 16'd9767, 16'd39857, 16'd5795});
	test_expansion(128'h622da770c5381ebf5b717fb555174dc8, {16'd52482, 16'd14664, 16'd34111, 16'd16342, 16'd58777, 16'd50182, 16'd63996, 16'd11207, 16'd60985, 16'd24109, 16'd26770, 16'd20760, 16'd62706, 16'd60383, 16'd64840, 16'd32128, 16'd45144, 16'd50754, 16'd22069, 16'd59854, 16'd15408, 16'd8663, 16'd53045, 16'd30432, 16'd21056, 16'd59541});
	test_expansion(128'h0cdf33c0ed69477798a745be1043c85a, {16'd46218, 16'd41371, 16'd25886, 16'd221, 16'd52409, 16'd60360, 16'd64237, 16'd49240, 16'd22915, 16'd40417, 16'd49140, 16'd53944, 16'd42234, 16'd12046, 16'd25772, 16'd57292, 16'd17638, 16'd28304, 16'd45514, 16'd33879, 16'd14014, 16'd34683, 16'd15991, 16'd63787, 16'd53674, 16'd9920});
	test_expansion(128'h629b42a3ad2d966d650e318844a1514a, {16'd37963, 16'd9686, 16'd31133, 16'd55195, 16'd33893, 16'd53894, 16'd62632, 16'd29172, 16'd43605, 16'd10605, 16'd31634, 16'd25378, 16'd61807, 16'd11063, 16'd46447, 16'd58564, 16'd34061, 16'd50411, 16'd7115, 16'd14770, 16'd6538, 16'd22198, 16'd20805, 16'd58072, 16'd20994, 16'd63004});
	test_expansion(128'hd9fdd7128764dc10495d4bb2dd5aa4c7, {16'd5644, 16'd38747, 16'd46487, 16'd64636, 16'd8100, 16'd17382, 16'd30063, 16'd54233, 16'd8912, 16'd33529, 16'd55455, 16'd54502, 16'd18609, 16'd52976, 16'd25043, 16'd7685, 16'd43122, 16'd9033, 16'd63949, 16'd33766, 16'd29231, 16'd24266, 16'd15610, 16'd37887, 16'd55706, 16'd61563});
	test_expansion(128'h06633621f191e9e0103419c8a5251dba, {16'd26905, 16'd8829, 16'd61519, 16'd32143, 16'd33115, 16'd9903, 16'd15730, 16'd27626, 16'd49053, 16'd51842, 16'd42230, 16'd34970, 16'd52772, 16'd24323, 16'd19746, 16'd56518, 16'd56744, 16'd4238, 16'd28825, 16'd54855, 16'd61701, 16'd33472, 16'd20298, 16'd44003, 16'd41781, 16'd63476});
	test_expansion(128'h7af1f00f81dc4e3c769d0d174309db9a, {16'd43223, 16'd29036, 16'd25050, 16'd21110, 16'd42817, 16'd49091, 16'd5553, 16'd11750, 16'd53897, 16'd2721, 16'd20955, 16'd26720, 16'd27780, 16'd23329, 16'd3290, 16'd45170, 16'd2284, 16'd8831, 16'd11410, 16'd6397, 16'd9546, 16'd62319, 16'd56222, 16'd19553, 16'd34062, 16'd51081});
	test_expansion(128'h5af0aa5b042c494ec4663353e5d620ee, {16'd26330, 16'd15191, 16'd42729, 16'd40960, 16'd4513, 16'd27292, 16'd8218, 16'd19532, 16'd49226, 16'd51467, 16'd26147, 16'd53033, 16'd36773, 16'd21965, 16'd7546, 16'd3174, 16'd64604, 16'd50784, 16'd52496, 16'd23340, 16'd60716, 16'd8693, 16'd46745, 16'd44669, 16'd12859, 16'd13014});
	test_expansion(128'h1760f5619bf713ec2240f8966b11061f, {16'd52006, 16'd5399, 16'd14063, 16'd45178, 16'd46256, 16'd3094, 16'd49889, 16'd23298, 16'd31167, 16'd15655, 16'd51152, 16'd33851, 16'd18720, 16'd1587, 16'd20755, 16'd38232, 16'd15844, 16'd13674, 16'd52539, 16'd30624, 16'd15550, 16'd39890, 16'd34916, 16'd48876, 16'd1504, 16'd33681});
	test_expansion(128'h245c97b2e60a519c788c60e2c6b77085, {16'd26434, 16'd4283, 16'd57064, 16'd18227, 16'd54050, 16'd2835, 16'd11241, 16'd239, 16'd21204, 16'd53382, 16'd9924, 16'd63960, 16'd33874, 16'd31659, 16'd12466, 16'd53507, 16'd8425, 16'd13789, 16'd64808, 16'd40488, 16'd61359, 16'd18303, 16'd35056, 16'd39635, 16'd57981, 16'd61229});
	test_expansion(128'h7aacb9adcb7141caba39027c7b08652c, {16'd32178, 16'd17099, 16'd57589, 16'd34007, 16'd15822, 16'd39799, 16'd7065, 16'd42350, 16'd19439, 16'd11302, 16'd50001, 16'd16016, 16'd49313, 16'd12553, 16'd55380, 16'd48733, 16'd22920, 16'd9309, 16'd10690, 16'd9736, 16'd50236, 16'd6, 16'd2941, 16'd27702, 16'd36565, 16'd51354});
	test_expansion(128'h102da7c0a9eb11e21dc6449b18193ec9, {16'd29488, 16'd3306, 16'd53571, 16'd37312, 16'd59742, 16'd30206, 16'd29738, 16'd62991, 16'd8793, 16'd30651, 16'd43733, 16'd37461, 16'd3656, 16'd45660, 16'd40026, 16'd17109, 16'd17750, 16'd37050, 16'd28999, 16'd33692, 16'd43195, 16'd37478, 16'd43357, 16'd15882, 16'd7975, 16'd55458});
	test_expansion(128'h90cd2559fdbc5265c7762249f7e624a9, {16'd57682, 16'd22774, 16'd17939, 16'd60030, 16'd58499, 16'd13344, 16'd6971, 16'd62583, 16'd43519, 16'd6645, 16'd54192, 16'd47208, 16'd20832, 16'd38591, 16'd14262, 16'd6191, 16'd24389, 16'd27988, 16'd14087, 16'd7183, 16'd45102, 16'd37134, 16'd2262, 16'd50897, 16'd53906, 16'd63320});
	test_expansion(128'haca374a584a68463940bd0975217eb69, {16'd53521, 16'd25975, 16'd57993, 16'd46422, 16'd62623, 16'd54880, 16'd58161, 16'd21155, 16'd29734, 16'd543, 16'd14332, 16'd33004, 16'd15191, 16'd47931, 16'd5108, 16'd63682, 16'd11173, 16'd188, 16'd46601, 16'd23156, 16'd16796, 16'd6208, 16'd26883, 16'd14362, 16'd25183, 16'd59602});
	test_expansion(128'h8f734e9889dcf5911662a04510024a13, {16'd11000, 16'd60717, 16'd17615, 16'd57427, 16'd65115, 16'd1223, 16'd5216, 16'd53876, 16'd13731, 16'd11489, 16'd55609, 16'd62378, 16'd20138, 16'd52942, 16'd4268, 16'd47028, 16'd19520, 16'd41476, 16'd55609, 16'd24765, 16'd12860, 16'd8689, 16'd21400, 16'd11653, 16'd221, 16'd36045});
	test_expansion(128'h3cfec7806fb51abaec6f3ce084b15e47, {16'd60088, 16'd24698, 16'd11796, 16'd5174, 16'd55643, 16'd62449, 16'd57094, 16'd53257, 16'd16765, 16'd59735, 16'd16643, 16'd52195, 16'd4942, 16'd44070, 16'd49531, 16'd170, 16'd55007, 16'd42106, 16'd39809, 16'd60633, 16'd57769, 16'd49189, 16'd28915, 16'd48571, 16'd30753, 16'd61549});
	test_expansion(128'he9b1c0604de960816f3e38af49d01fdc, {16'd54917, 16'd51141, 16'd21326, 16'd37312, 16'd9814, 16'd9221, 16'd4992, 16'd13446, 16'd3772, 16'd1771, 16'd49928, 16'd43799, 16'd8784, 16'd23620, 16'd45825, 16'd18373, 16'd51853, 16'd47205, 16'd50660, 16'd49853, 16'd38809, 16'd31769, 16'd11174, 16'd33381, 16'd31294, 16'd52188});
	test_expansion(128'he92a9719c122fa7c9dfd04a4cd254e96, {16'd29212, 16'd27764, 16'd4523, 16'd54052, 16'd24648, 16'd57229, 16'd7551, 16'd50320, 16'd2373, 16'd62335, 16'd29055, 16'd40482, 16'd10585, 16'd44333, 16'd15560, 16'd26975, 16'd56365, 16'd12948, 16'd4530, 16'd4896, 16'd16875, 16'd36594, 16'd42421, 16'd51796, 16'd31471, 16'd57036});
	test_expansion(128'hbbee8f27cd38677efadfa34ed06e0626, {16'd38444, 16'd46230, 16'd25512, 16'd29151, 16'd28876, 16'd8071, 16'd47488, 16'd42366, 16'd13275, 16'd37984, 16'd59492, 16'd45926, 16'd33772, 16'd22763, 16'd23270, 16'd5019, 16'd30639, 16'd27351, 16'd1072, 16'd56622, 16'd8069, 16'd63508, 16'd27294, 16'd16400, 16'd20633, 16'd15791});
	test_expansion(128'h0d9d7a74bcac7eef54467629a82d4d52, {16'd57214, 16'd44327, 16'd8914, 16'd58287, 16'd6010, 16'd53972, 16'd2304, 16'd32261, 16'd28198, 16'd57584, 16'd8652, 16'd43060, 16'd25429, 16'd55855, 16'd41952, 16'd13073, 16'd61623, 16'd64769, 16'd2801, 16'd29536, 16'd58993, 16'd31927, 16'd47163, 16'd18357, 16'd62209, 16'd12265});
	test_expansion(128'hfd97ddc1a833d0a1c60fc930803b5d41, {16'd38692, 16'd30286, 16'd12067, 16'd52819, 16'd27757, 16'd10176, 16'd58991, 16'd59411, 16'd31171, 16'd14373, 16'd833, 16'd62253, 16'd54412, 16'd35565, 16'd30644, 16'd42732, 16'd5452, 16'd37789, 16'd7915, 16'd33890, 16'd32462, 16'd21798, 16'd60824, 16'd29711, 16'd18309, 16'd44895});
	test_expansion(128'hfb89f23365189ad7783a006ba4ff1abe, {16'd18809, 16'd17802, 16'd45384, 16'd35536, 16'd14461, 16'd38981, 16'd28017, 16'd17084, 16'd11352, 16'd39928, 16'd24410, 16'd8094, 16'd45296, 16'd61791, 16'd56271, 16'd42076, 16'd9231, 16'd57191, 16'd9257, 16'd27286, 16'd2677, 16'd47892, 16'd17849, 16'd55071, 16'd27590, 16'd36773});
	test_expansion(128'hc4a9e531b2d33ea09102d3c6a82a6c30, {16'd15375, 16'd62374, 16'd44353, 16'd32541, 16'd33575, 16'd9558, 16'd2020, 16'd6877, 16'd38163, 16'd7969, 16'd45161, 16'd26801, 16'd5710, 16'd59928, 16'd16029, 16'd56128, 16'd49352, 16'd20477, 16'd49636, 16'd51216, 16'd53931, 16'd44021, 16'd38995, 16'd20368, 16'd16876, 16'd16702});
	test_expansion(128'ha70e3099512a87b67f5622917b27ad9b, {16'd46224, 16'd56821, 16'd60182, 16'd3122, 16'd4955, 16'd24635, 16'd9004, 16'd48828, 16'd17439, 16'd61989, 16'd57336, 16'd1848, 16'd32691, 16'd53593, 16'd7669, 16'd9924, 16'd63353, 16'd27257, 16'd9479, 16'd59574, 16'd16073, 16'd686, 16'd5354, 16'd35592, 16'd11870, 16'd61991});
	test_expansion(128'hfc3a3bceae65cdf09d7115bd7130f538, {16'd48608, 16'd23982, 16'd14862, 16'd25888, 16'd21012, 16'd3607, 16'd63278, 16'd33927, 16'd65201, 16'd16774, 16'd54584, 16'd27856, 16'd21106, 16'd62169, 16'd47337, 16'd3414, 16'd14751, 16'd131, 16'd48696, 16'd27105, 16'd14141, 16'd59971, 16'd28453, 16'd51308, 16'd35559, 16'd13373});
	test_expansion(128'h336bbc28c931142d4be203b5f214de43, {16'd17809, 16'd32590, 16'd49553, 16'd38924, 16'd59704, 16'd61237, 16'd55672, 16'd38431, 16'd11833, 16'd35627, 16'd5374, 16'd22460, 16'd8215, 16'd38438, 16'd33515, 16'd19151, 16'd53202, 16'd51812, 16'd54803, 16'd26611, 16'd22457, 16'd30824, 16'd50652, 16'd10402, 16'd13333, 16'd16011});
	test_expansion(128'h48024046fc33f29a43454b7033293e14, {16'd10113, 16'd1539, 16'd47646, 16'd56093, 16'd44502, 16'd51724, 16'd48094, 16'd17678, 16'd53272, 16'd1770, 16'd51703, 16'd50352, 16'd64321, 16'd9707, 16'd27416, 16'd64215, 16'd25833, 16'd36831, 16'd45284, 16'd35900, 16'd32363, 16'd27520, 16'd30441, 16'd34907, 16'd22026, 16'd42013});
	test_expansion(128'he4ec19ff8ae2f538fbd475e956caebce, {16'd26328, 16'd49343, 16'd14060, 16'd26275, 16'd29755, 16'd41544, 16'd8282, 16'd44817, 16'd15013, 16'd62527, 16'd39056, 16'd48530, 16'd23609, 16'd8243, 16'd4624, 16'd26743, 16'd27408, 16'd49127, 16'd27699, 16'd22568, 16'd32878, 16'd21480, 16'd45605, 16'd25623, 16'd34712, 16'd51134});
	test_expansion(128'h5ce9f411484d0e7e21657f88215df3bb, {16'd59718, 16'd23232, 16'd26583, 16'd10596, 16'd56174, 16'd2605, 16'd25732, 16'd51643, 16'd16261, 16'd14307, 16'd7778, 16'd24193, 16'd10796, 16'd65177, 16'd26939, 16'd30720, 16'd36172, 16'd1322, 16'd53919, 16'd5510, 16'd4540, 16'd10059, 16'd37807, 16'd10671, 16'd50337, 16'd38318});
	test_expansion(128'hd824f0a6864d413d45624eefeade1fd9, {16'd21918, 16'd64018, 16'd54875, 16'd39442, 16'd39023, 16'd10851, 16'd571, 16'd18802, 16'd45014, 16'd28989, 16'd43409, 16'd21905, 16'd52654, 16'd32678, 16'd16441, 16'd58776, 16'd3802, 16'd63763, 16'd15255, 16'd15518, 16'd35414, 16'd58697, 16'd6379, 16'd60721, 16'd9309, 16'd64886});
	test_expansion(128'h2f1d2c35167725754d5b9d2b2135738d, {16'd20591, 16'd13433, 16'd44754, 16'd37931, 16'd58816, 16'd7984, 16'd3860, 16'd25318, 16'd44862, 16'd57159, 16'd51592, 16'd8028, 16'd8959, 16'd17318, 16'd1356, 16'd10831, 16'd22134, 16'd7808, 16'd25908, 16'd26246, 16'd41672, 16'd58114, 16'd56429, 16'd46172, 16'd7009, 16'd42225});
	test_expansion(128'h950061e9bdbe1131beae29170b17e6cf, {16'd41588, 16'd16699, 16'd55043, 16'd39348, 16'd11470, 16'd12689, 16'd43796, 16'd8165, 16'd47224, 16'd54934, 16'd24447, 16'd28736, 16'd24852, 16'd11236, 16'd36090, 16'd29030, 16'd43400, 16'd58828, 16'd44350, 16'd8578, 16'd26474, 16'd16889, 16'd46378, 16'd37692, 16'd38567, 16'd30805});
	test_expansion(128'ha082df6d69561d7280f7e19d8734f5f5, {16'd12387, 16'd16639, 16'd58253, 16'd3185, 16'd19201, 16'd40024, 16'd853, 16'd41141, 16'd28660, 16'd6168, 16'd47261, 16'd21788, 16'd50279, 16'd41046, 16'd35530, 16'd43640, 16'd59465, 16'd41397, 16'd26640, 16'd25642, 16'd16, 16'd30867, 16'd7374, 16'd50356, 16'd43754, 16'd5469});
	test_expansion(128'hc47dd0796163e618868e4005574d5ae8, {16'd57464, 16'd10012, 16'd61958, 16'd15576, 16'd26198, 16'd13179, 16'd12891, 16'd58143, 16'd58945, 16'd53952, 16'd28481, 16'd41112, 16'd59194, 16'd18426, 16'd34780, 16'd997, 16'd61181, 16'd32901, 16'd10371, 16'd59325, 16'd7851, 16'd19885, 16'd3082, 16'd14042, 16'd51207, 16'd6325});
	test_expansion(128'hbbd91540f84708f2781bb4f8ef847e92, {16'd47095, 16'd63967, 16'd42086, 16'd57471, 16'd9642, 16'd52942, 16'd18370, 16'd29999, 16'd28795, 16'd11339, 16'd28720, 16'd63173, 16'd5542, 16'd22657, 16'd46985, 16'd49842, 16'd36481, 16'd6997, 16'd3451, 16'd6231, 16'd51800, 16'd12412, 16'd51379, 16'd30521, 16'd27585, 16'd12129});
	test_expansion(128'hf0d179e64d5726b2ead24479df9f46cb, {16'd22139, 16'd7224, 16'd42489, 16'd16815, 16'd9747, 16'd64512, 16'd53571, 16'd65058, 16'd36652, 16'd52090, 16'd52126, 16'd10965, 16'd43378, 16'd42976, 16'd19617, 16'd8787, 16'd41660, 16'd30769, 16'd10544, 16'd25237, 16'd7196, 16'd33525, 16'd60295, 16'd14963, 16'd60545, 16'd1276});
	test_expansion(128'h4a67f366f7f3bd906f4ec6684036f160, {16'd11232, 16'd4580, 16'd16388, 16'd21194, 16'd50614, 16'd138, 16'd1111, 16'd4183, 16'd2152, 16'd40150, 16'd30157, 16'd43858, 16'd46082, 16'd64469, 16'd53747, 16'd50251, 16'd38821, 16'd19972, 16'd36534, 16'd10589, 16'd23440, 16'd342, 16'd51634, 16'd30742, 16'd9047, 16'd55115});
	test_expansion(128'h76c497fef724b8a6ddf88153f587af2a, {16'd12172, 16'd36428, 16'd19946, 16'd6220, 16'd42120, 16'd56070, 16'd37212, 16'd12180, 16'd44583, 16'd52546, 16'd10280, 16'd42270, 16'd31858, 16'd31832, 16'd20984, 16'd57791, 16'd26825, 16'd6287, 16'd53826, 16'd57146, 16'd23320, 16'd6522, 16'd16578, 16'd42563, 16'd42075, 16'd12037});
	test_expansion(128'he9e20cf00596d24bf3e95381d8c40cce, {16'd1843, 16'd7162, 16'd10606, 16'd481, 16'd62617, 16'd16896, 16'd42516, 16'd45618, 16'd29505, 16'd49676, 16'd26355, 16'd58750, 16'd36044, 16'd59414, 16'd25232, 16'd14896, 16'd16043, 16'd4460, 16'd59083, 16'd27779, 16'd45065, 16'd2667, 16'd41233, 16'd50905, 16'd19466, 16'd41276});
	test_expansion(128'h4ee90699a99dbb1e0724b70a208854bf, {16'd17420, 16'd40959, 16'd62265, 16'd59395, 16'd44960, 16'd56308, 16'd60171, 16'd23758, 16'd11423, 16'd29671, 16'd57186, 16'd1875, 16'd10530, 16'd46814, 16'd31995, 16'd63167, 16'd26958, 16'd23053, 16'd62824, 16'd12508, 16'd63107, 16'd43120, 16'd24316, 16'd48918, 16'd40739, 16'd46150});
	test_expansion(128'h086d96140f68e73257a826bbd199e7f6, {16'd58347, 16'd9799, 16'd11052, 16'd18548, 16'd26900, 16'd56635, 16'd9595, 16'd34953, 16'd18501, 16'd65264, 16'd57303, 16'd38434, 16'd43220, 16'd4542, 16'd57484, 16'd62243, 16'd31780, 16'd14011, 16'd41481, 16'd32225, 16'd17536, 16'd37331, 16'd4600, 16'd23934, 16'd32157, 16'd38381});
	test_expansion(128'he3e297867efcf2b302321c3fafceb2ab, {16'd52259, 16'd36240, 16'd19147, 16'd12872, 16'd19240, 16'd54390, 16'd14010, 16'd36547, 16'd39821, 16'd9456, 16'd35029, 16'd44635, 16'd12220, 16'd34795, 16'd17401, 16'd61783, 16'd24124, 16'd26331, 16'd48928, 16'd59321, 16'd48988, 16'd10456, 16'd11587, 16'd6573, 16'd63851, 16'd29068});
	test_expansion(128'h689073ef3f4c0303e07a932edecbe548, {16'd6976, 16'd32203, 16'd39238, 16'd40726, 16'd5440, 16'd62811, 16'd2401, 16'd18006, 16'd35898, 16'd37349, 16'd34657, 16'd33854, 16'd49276, 16'd55876, 16'd61162, 16'd12734, 16'd47934, 16'd16938, 16'd51153, 16'd11294, 16'd25610, 16'd3226, 16'd5943, 16'd21422, 16'd34993, 16'd61649});
	test_expansion(128'hbe16ddf65b2b5c5e8cde8022e6fe8247, {16'd9682, 16'd22739, 16'd34150, 16'd56118, 16'd53251, 16'd13443, 16'd14406, 16'd11013, 16'd7434, 16'd6792, 16'd18329, 16'd35464, 16'd24538, 16'd63801, 16'd18010, 16'd8256, 16'd64936, 16'd17384, 16'd28592, 16'd27105, 16'd43553, 16'd58958, 16'd51660, 16'd19624, 16'd41133, 16'd15021});
	test_expansion(128'hcd20277a2f33254085ac904fef58d125, {16'd39956, 16'd24588, 16'd65488, 16'd59300, 16'd53769, 16'd17934, 16'd40602, 16'd59587, 16'd47520, 16'd21993, 16'd28785, 16'd46954, 16'd37926, 16'd59930, 16'd29902, 16'd9293, 16'd53359, 16'd43771, 16'd976, 16'd29925, 16'd22180, 16'd3001, 16'd53258, 16'd45372, 16'd12829, 16'd24358});
	test_expansion(128'haa583dae3b84a56b0941eaf68655b78b, {16'd58898, 16'd10740, 16'd64324, 16'd9994, 16'd44815, 16'd34486, 16'd56618, 16'd50156, 16'd31810, 16'd31453, 16'd7000, 16'd56466, 16'd14855, 16'd20729, 16'd10300, 16'd62669, 16'd7162, 16'd28854, 16'd60788, 16'd41610, 16'd51798, 16'd63064, 16'd53825, 16'd15180, 16'd14783, 16'd24401});
	test_expansion(128'he5de307941b23d90b5e3e08a2b70dab6, {16'd5725, 16'd54805, 16'd2462, 16'd41217, 16'd1534, 16'd23730, 16'd51281, 16'd26890, 16'd35457, 16'd30578, 16'd1488, 16'd23490, 16'd63986, 16'd52730, 16'd27077, 16'd11840, 16'd52160, 16'd61287, 16'd28345, 16'd46254, 16'd61566, 16'd18516, 16'd14928, 16'd42439, 16'd29307, 16'd17585});
	test_expansion(128'h52cedeeafd28e285c8b9ce189e0cf6a6, {16'd31226, 16'd22838, 16'd19770, 16'd60565, 16'd49556, 16'd19, 16'd15128, 16'd17925, 16'd54940, 16'd49596, 16'd44403, 16'd45376, 16'd15860, 16'd60162, 16'd49090, 16'd33018, 16'd38994, 16'd7561, 16'd63695, 16'd44273, 16'd14829, 16'd38215, 16'd14786, 16'd2042, 16'd47898, 16'd31417});
	test_expansion(128'h741e7ac07049091486630f83dd12e89a, {16'd10259, 16'd16207, 16'd31927, 16'd57279, 16'd35725, 16'd36441, 16'd61786, 16'd12237, 16'd44685, 16'd64722, 16'd61948, 16'd35052, 16'd64341, 16'd30221, 16'd30833, 16'd65260, 16'd8579, 16'd13949, 16'd12, 16'd58271, 16'd29497, 16'd38109, 16'd21038, 16'd47064, 16'd25679, 16'd33391});
	test_expansion(128'hf1846acdbb80a17620bc157f62eab6ef, {16'd11065, 16'd65337, 16'd39114, 16'd52583, 16'd439, 16'd17200, 16'd58585, 16'd3975, 16'd22029, 16'd34216, 16'd45878, 16'd64655, 16'd25736, 16'd16521, 16'd59749, 16'd7767, 16'd4484, 16'd37978, 16'd46348, 16'd61690, 16'd54851, 16'd26446, 16'd38052, 16'd36528, 16'd62226, 16'd34534});
	test_expansion(128'h68ce0627038fef6d69ebe06da9ff86ff, {16'd36806, 16'd31384, 16'd43701, 16'd38882, 16'd11288, 16'd4387, 16'd41162, 16'd2348, 16'd9300, 16'd50680, 16'd51116, 16'd6040, 16'd32288, 16'd46098, 16'd2022, 16'd34692, 16'd1053, 16'd33136, 16'd7651, 16'd39265, 16'd64436, 16'd44224, 16'd14830, 16'd30450, 16'd5827, 16'd4027});
	test_expansion(128'ha31bfd125ee0ebb7de9bbb7a4fef1835, {16'd48473, 16'd58302, 16'd31080, 16'd6278, 16'd40229, 16'd29584, 16'd3478, 16'd32347, 16'd37708, 16'd593, 16'd25500, 16'd28826, 16'd11020, 16'd17844, 16'd32244, 16'd9243, 16'd46138, 16'd32645, 16'd63506, 16'd16963, 16'd3255, 16'd7809, 16'd20670, 16'd34529, 16'd51734, 16'd2274});
	test_expansion(128'h9f5a1eb8e0f077e62b0bd27231673f9a, {16'd34603, 16'd24826, 16'd45136, 16'd61068, 16'd2887, 16'd38947, 16'd28238, 16'd35243, 16'd27309, 16'd27273, 16'd53024, 16'd6283, 16'd58939, 16'd64055, 16'd30024, 16'd12523, 16'd4988, 16'd34460, 16'd52031, 16'd49661, 16'd43448, 16'd26746, 16'd54935, 16'd34683, 16'd59208, 16'd33148});
	test_expansion(128'h2a47094e7d51fd2c8fc5308c2121db1f, {16'd51682, 16'd63881, 16'd4508, 16'd6279, 16'd32389, 16'd38795, 16'd4034, 16'd8037, 16'd57449, 16'd29797, 16'd21560, 16'd350, 16'd16304, 16'd42126, 16'd47127, 16'd19138, 16'd42989, 16'd13185, 16'd58131, 16'd53782, 16'd1510, 16'd29734, 16'd17210, 16'd29969, 16'd5425, 16'd51136});
	test_expansion(128'hfc31af358579223577e902f021ad8f8c, {16'd40322, 16'd56430, 16'd24981, 16'd54472, 16'd45581, 16'd10197, 16'd60851, 16'd63547, 16'd47823, 16'd50876, 16'd59856, 16'd24081, 16'd61122, 16'd26692, 16'd29477, 16'd43670, 16'd33768, 16'd14513, 16'd36817, 16'd19029, 16'd40119, 16'd33561, 16'd53103, 16'd43345, 16'd34717, 16'd28906});
	test_expansion(128'hf9f356c7c9dc9e328375ddfc92ef7e5a, {16'd12979, 16'd9085, 16'd47217, 16'd8353, 16'd1882, 16'd60743, 16'd1575, 16'd42069, 16'd23379, 16'd16433, 16'd43681, 16'd58495, 16'd60575, 16'd7377, 16'd38956, 16'd27707, 16'd37595, 16'd62106, 16'd3707, 16'd47481, 16'd16161, 16'd11947, 16'd52176, 16'd59899, 16'd50573, 16'd48696});
	test_expansion(128'h32b5b589cbc9324071126582bfea356a, {16'd20277, 16'd23126, 16'd23969, 16'd40961, 16'd40267, 16'd63515, 16'd60898, 16'd26674, 16'd55702, 16'd10429, 16'd1607, 16'd9983, 16'd64168, 16'd8749, 16'd11355, 16'd1616, 16'd15568, 16'd60753, 16'd56636, 16'd22377, 16'd29405, 16'd11697, 16'd47580, 16'd16636, 16'd11711, 16'd21613});
	test_expansion(128'h2468d7f865f6e90c79fc79a4b9a98c4e, {16'd27700, 16'd21590, 16'd6144, 16'd58134, 16'd11043, 16'd50144, 16'd41439, 16'd8828, 16'd45570, 16'd60059, 16'd51944, 16'd56376, 16'd33501, 16'd32864, 16'd55873, 16'd19985, 16'd5363, 16'd36447, 16'd39185, 16'd24640, 16'd50593, 16'd21354, 16'd34741, 16'd44733, 16'd65416, 16'd18424});
	test_expansion(128'h39acacdb5d1352060dcd8bbe0d2591ff, {16'd669, 16'd11395, 16'd15948, 16'd43466, 16'd12188, 16'd5643, 16'd47238, 16'd11659, 16'd4539, 16'd27408, 16'd34641, 16'd7272, 16'd32409, 16'd56320, 16'd40503, 16'd2388, 16'd65060, 16'd28791, 16'd22330, 16'd47123, 16'd26765, 16'd15688, 16'd40908, 16'd23830, 16'd41607, 16'd1393});
	test_expansion(128'he213e65575a06f5f2d7141d64c1ed532, {16'd7958, 16'd65346, 16'd4857, 16'd53110, 16'd31047, 16'd40261, 16'd55648, 16'd64868, 16'd29226, 16'd4186, 16'd48868, 16'd2172, 16'd16959, 16'd44842, 16'd33193, 16'd60058, 16'd57178, 16'd61292, 16'd40756, 16'd7631, 16'd58722, 16'd54193, 16'd59827, 16'd32287, 16'd26493, 16'd25792});
	test_expansion(128'h8d897d1e597fcee6fa0b8672fbce9223, {16'd1123, 16'd33124, 16'd27831, 16'd65435, 16'd42001, 16'd40726, 16'd65461, 16'd58687, 16'd56974, 16'd23514, 16'd19755, 16'd32791, 16'd19211, 16'd61862, 16'd24313, 16'd11689, 16'd36821, 16'd62355, 16'd37751, 16'd61684, 16'd17356, 16'd20009, 16'd7972, 16'd2002, 16'd64405, 16'd31235});
	test_expansion(128'h7a971506b5e147b6283782a3c6afc38f, {16'd43251, 16'd50612, 16'd60337, 16'd61205, 16'd61661, 16'd55958, 16'd40183, 16'd61018, 16'd57730, 16'd37271, 16'd29423, 16'd15553, 16'd42086, 16'd21620, 16'd7175, 16'd48325, 16'd51608, 16'd21389, 16'd13878, 16'd17417, 16'd50571, 16'd52113, 16'd35981, 16'd49660, 16'd44419, 16'd21564});
	test_expansion(128'h20763c693cdf182e6ec2c8bb5ff1412e, {16'd28630, 16'd46194, 16'd58043, 16'd50773, 16'd27670, 16'd38637, 16'd9517, 16'd15164, 16'd53450, 16'd38335, 16'd37861, 16'd54654, 16'd5711, 16'd12386, 16'd29892, 16'd54559, 16'd22717, 16'd10423, 16'd40399, 16'd3228, 16'd17728, 16'd38125, 16'd41619, 16'd9353, 16'd23158, 16'd56042});
	test_expansion(128'h2f4506a91c3e434e98f440577af34c6f, {16'd61791, 16'd62089, 16'd49064, 16'd20374, 16'd47120, 16'd48504, 16'd19927, 16'd48345, 16'd14003, 16'd60368, 16'd31378, 16'd56165, 16'd58930, 16'd40736, 16'd40571, 16'd38796, 16'd14678, 16'd51057, 16'd56107, 16'd56824, 16'd8324, 16'd381, 16'd56311, 16'd12602, 16'd16319, 16'd37438});
	test_expansion(128'h883ce59dd28ba94581193ba23de27375, {16'd46965, 16'd26323, 16'd29388, 16'd38748, 16'd52427, 16'd9999, 16'd36324, 16'd4814, 16'd51870, 16'd7595, 16'd42656, 16'd58842, 16'd53402, 16'd4432, 16'd32735, 16'd352, 16'd12889, 16'd54844, 16'd7545, 16'd5812, 16'd29863, 16'd64806, 16'd38632, 16'd57099, 16'd39559, 16'd2761});
	test_expansion(128'h1419bec15ea9b6b887d37e66cb6720e7, {16'd43251, 16'd24695, 16'd40935, 16'd11093, 16'd4624, 16'd4611, 16'd44445, 16'd57136, 16'd48456, 16'd12167, 16'd34221, 16'd10679, 16'd12906, 16'd27550, 16'd24193, 16'd59229, 16'd50778, 16'd54807, 16'd48112, 16'd24359, 16'd24970, 16'd9320, 16'd111, 16'd41987, 16'd50018, 16'd25821});
	test_expansion(128'ha22da243422d81ac4fa184b42cfdd830, {16'd29154, 16'd6878, 16'd37734, 16'd24643, 16'd6732, 16'd22138, 16'd16939, 16'd41922, 16'd49914, 16'd60042, 16'd53065, 16'd16364, 16'd3531, 16'd40028, 16'd22597, 16'd10132, 16'd27779, 16'd51121, 16'd28342, 16'd12019, 16'd15281, 16'd58939, 16'd112, 16'd7837, 16'd12382, 16'd27203});
	test_expansion(128'hd36e6e8c54c4e6026fc9e5308f7ad370, {16'd57139, 16'd23069, 16'd15320, 16'd30233, 16'd32290, 16'd41026, 16'd48729, 16'd61176, 16'd29984, 16'd50699, 16'd65140, 16'd63205, 16'd51697, 16'd13198, 16'd6940, 16'd44237, 16'd34514, 16'd57390, 16'd42066, 16'd262, 16'd16093, 16'd6073, 16'd41290, 16'd68, 16'd26829, 16'd11297});
	test_expansion(128'h3f5e42631ec635ebc2986a2a6414af41, {16'd61029, 16'd44664, 16'd7502, 16'd8982, 16'd28588, 16'd38997, 16'd14658, 16'd63072, 16'd36656, 16'd45574, 16'd1270, 16'd16063, 16'd29301, 16'd65054, 16'd61506, 16'd23103, 16'd35641, 16'd55004, 16'd32575, 16'd19475, 16'd53347, 16'd5475, 16'd41125, 16'd11795, 16'd28469, 16'd40590});
	test_expansion(128'hce660bd48d19aa8dc95342a6653ac05a, {16'd14279, 16'd21223, 16'd30721, 16'd24454, 16'd16096, 16'd60317, 16'd9868, 16'd60118, 16'd31855, 16'd46147, 16'd58846, 16'd54280, 16'd56096, 16'd48064, 16'd28502, 16'd6992, 16'd43537, 16'd4759, 16'd9433, 16'd55798, 16'd33356, 16'd61112, 16'd21507, 16'd3624, 16'd2835, 16'd15907});
	test_expansion(128'h2abaec0d77c147e82f51553a5dbecc5d, {16'd6500, 16'd19934, 16'd9642, 16'd22377, 16'd10906, 16'd249, 16'd29034, 16'd26581, 16'd56112, 16'd19226, 16'd10575, 16'd30278, 16'd10104, 16'd24434, 16'd26998, 16'd14795, 16'd33816, 16'd38474, 16'd44154, 16'd54658, 16'd45349, 16'd9703, 16'd31424, 16'd60279, 16'd32706, 16'd903});
	test_expansion(128'h217856347a5fd00139c423acd37eead5, {16'd18600, 16'd7992, 16'd43895, 16'd10494, 16'd35743, 16'd63103, 16'd63385, 16'd31816, 16'd13360, 16'd54484, 16'd43840, 16'd41414, 16'd58993, 16'd6198, 16'd56864, 16'd57739, 16'd47301, 16'd44818, 16'd54468, 16'd33050, 16'd35547, 16'd58242, 16'd54539, 16'd52957, 16'd26194, 16'd32847});
	test_expansion(128'hf4be5b2e9f9e354ffff06e338aa7e54b, {16'd47201, 16'd20738, 16'd42502, 16'd7823, 16'd25875, 16'd12625, 16'd55128, 16'd21692, 16'd3813, 16'd51514, 16'd53803, 16'd10119, 16'd7816, 16'd16499, 16'd12857, 16'd40546, 16'd63177, 16'd35698, 16'd53705, 16'd34678, 16'd40045, 16'd6701, 16'd53433, 16'd60328, 16'd17437, 16'd13600});
	test_expansion(128'h5e11ebcd464481d3a9e04f0722f800a4, {16'd14234, 16'd16617, 16'd20599, 16'd35497, 16'd52800, 16'd61961, 16'd63090, 16'd64445, 16'd46361, 16'd4517, 16'd15061, 16'd41905, 16'd48808, 16'd63770, 16'd51981, 16'd27667, 16'd6166, 16'd30077, 16'd12401, 16'd52677, 16'd57218, 16'd49121, 16'd26380, 16'd754, 16'd46320, 16'd29653});
	test_expansion(128'hf0356d9de9782b25a555916e2828b836, {16'd63081, 16'd2723, 16'd15256, 16'd26311, 16'd18148, 16'd36607, 16'd56888, 16'd6900, 16'd50327, 16'd37301, 16'd20036, 16'd5524, 16'd7181, 16'd19168, 16'd21794, 16'd64720, 16'd45010, 16'd26061, 16'd3214, 16'd7279, 16'd59759, 16'd42077, 16'd48380, 16'd22738, 16'd59440, 16'd18839});
	test_expansion(128'h7a6b10eafc1402f4cc5f2b67ba85a9c1, {16'd1583, 16'd42909, 16'd37352, 16'd26927, 16'd14453, 16'd24706, 16'd24559, 16'd18268, 16'd9593, 16'd17015, 16'd34018, 16'd18363, 16'd6225, 16'd64970, 16'd55959, 16'd11764, 16'd2068, 16'd48455, 16'd51895, 16'd14483, 16'd13713, 16'd12734, 16'd6948, 16'd29289, 16'd4219, 16'd44868});
	test_expansion(128'hb56a3c6e83b968585a94097075b69337, {16'd16685, 16'd32284, 16'd7784, 16'd64154, 16'd18599, 16'd40285, 16'd35029, 16'd15640, 16'd10982, 16'd7146, 16'd17671, 16'd83, 16'd16586, 16'd12233, 16'd14079, 16'd46329, 16'd55404, 16'd45596, 16'd32127, 16'd4817, 16'd42257, 16'd33847, 16'd36872, 16'd55063, 16'd61542, 16'd25653});
	test_expansion(128'h5c05cd0f8c4623209ad480d282ef9903, {16'd8644, 16'd3888, 16'd7481, 16'd5833, 16'd3509, 16'd30548, 16'd55756, 16'd43203, 16'd5791, 16'd50886, 16'd18545, 16'd8814, 16'd63077, 16'd22172, 16'd47261, 16'd44253, 16'd1158, 16'd23328, 16'd57999, 16'd2531, 16'd57882, 16'd14600, 16'd55451, 16'd2498, 16'd19575, 16'd48585});
	test_expansion(128'hf6ebb0b88dbe63c58cc50471cba054a6, {16'd2468, 16'd52340, 16'd54875, 16'd4384, 16'd1933, 16'd49308, 16'd42555, 16'd35979, 16'd41972, 16'd32529, 16'd53983, 16'd63467, 16'd20543, 16'd55099, 16'd53462, 16'd11076, 16'd14419, 16'd25531, 16'd13428, 16'd17399, 16'd35467, 16'd21471, 16'd13772, 16'd59590, 16'd44763, 16'd42811});
	test_expansion(128'h8b80a23a625b2e05e3f60f63c2db79e3, {16'd58544, 16'd47787, 16'd59196, 16'd17000, 16'd49939, 16'd43613, 16'd56185, 16'd12831, 16'd34824, 16'd7594, 16'd63558, 16'd7835, 16'd544, 16'd55780, 16'd31751, 16'd42695, 16'd15250, 16'd36074, 16'd45669, 16'd106, 16'd7860, 16'd41812, 16'd9699, 16'd54998, 16'd14333, 16'd57618});
	test_expansion(128'hdbac54affdd5ff210e03acf3baba8538, {16'd14903, 16'd51486, 16'd35719, 16'd22521, 16'd3468, 16'd47882, 16'd26672, 16'd44741, 16'd21640, 16'd55383, 16'd27625, 16'd15123, 16'd36045, 16'd24294, 16'd60054, 16'd33343, 16'd5887, 16'd56315, 16'd12751, 16'd55329, 16'd47868, 16'd7866, 16'd46613, 16'd51617, 16'd43809, 16'd5652});
	test_expansion(128'h2f0ccb02d96f360a1600c75c02fc1bae, {16'd26996, 16'd54443, 16'd64155, 16'd50362, 16'd63213, 16'd38055, 16'd45007, 16'd48276, 16'd41592, 16'd7283, 16'd6280, 16'd58519, 16'd27662, 16'd9493, 16'd12116, 16'd11634, 16'd33700, 16'd15012, 16'd56007, 16'd39454, 16'd32090, 16'd19161, 16'd55599, 16'd39428, 16'd9871, 16'd29987});
	test_expansion(128'he51c459390355d8955b7e91652476fc9, {16'd8185, 16'd24373, 16'd15307, 16'd49517, 16'd19307, 16'd42344, 16'd27323, 16'd58509, 16'd20806, 16'd48202, 16'd28868, 16'd27768, 16'd3797, 16'd20223, 16'd63841, 16'd10783, 16'd16655, 16'd21941, 16'd5632, 16'd20439, 16'd55291, 16'd47226, 16'd18225, 16'd11708, 16'd8354, 16'd22648});
	test_expansion(128'hb8f538c54cd7f07d64935eac83c906ec, {16'd918, 16'd55779, 16'd49132, 16'd40895, 16'd10510, 16'd24006, 16'd14618, 16'd32803, 16'd6941, 16'd4560, 16'd24159, 16'd15876, 16'd29462, 16'd56789, 16'd3667, 16'd52112, 16'd28183, 16'd51091, 16'd45247, 16'd59761, 16'd62193, 16'd53020, 16'd28977, 16'd43123, 16'd49457, 16'd22304});
	test_expansion(128'hb112b11d05e4c0897f7a63126c355ebc, {16'd1390, 16'd42725, 16'd43880, 16'd16884, 16'd32303, 16'd63515, 16'd11779, 16'd6174, 16'd13017, 16'd55161, 16'd25727, 16'd55609, 16'd55635, 16'd14193, 16'd58255, 16'd455, 16'd7963, 16'd60256, 16'd29082, 16'd17961, 16'd64634, 16'd18857, 16'd30310, 16'd14147, 16'd45604, 16'd6435});
	test_expansion(128'hb7c798d43872a66516da4a53f922903a, {16'd16290, 16'd55217, 16'd5141, 16'd26887, 16'd55645, 16'd4488, 16'd58847, 16'd15239, 16'd10772, 16'd16244, 16'd51287, 16'd38315, 16'd30567, 16'd21632, 16'd53962, 16'd3305, 16'd17063, 16'd12998, 16'd41293, 16'd54504, 16'd52401, 16'd21936, 16'd17446, 16'd38706, 16'd52874, 16'd40640});
	test_expansion(128'hf64b2792a1034b1009b43364be2dfbb3, {16'd55906, 16'd27038, 16'd24157, 16'd42973, 16'd2745, 16'd42919, 16'd26563, 16'd62407, 16'd34819, 16'd6965, 16'd40565, 16'd4650, 16'd28256, 16'd17606, 16'd61877, 16'd38953, 16'd51380, 16'd41188, 16'd42686, 16'd13489, 16'd58282, 16'd918, 16'd22750, 16'd28778, 16'd36917, 16'd3925});
	test_expansion(128'h3b28b7293c38bf5dfcb68031912e4db3, {16'd56928, 16'd17711, 16'd11443, 16'd23293, 16'd58540, 16'd55583, 16'd10094, 16'd38162, 16'd52566, 16'd37915, 16'd2099, 16'd59851, 16'd51048, 16'd16566, 16'd63421, 16'd42225, 16'd28818, 16'd22206, 16'd47658, 16'd30046, 16'd54925, 16'd30322, 16'd51639, 16'd46862, 16'd35468, 16'd21675});
	test_expansion(128'h8d8f96552bed9c49d6d836007a9d927b, {16'd26627, 16'd35917, 16'd40071, 16'd30989, 16'd57432, 16'd34033, 16'd42135, 16'd54209, 16'd18597, 16'd13989, 16'd57183, 16'd11318, 16'd60803, 16'd14133, 16'd26115, 16'd27772, 16'd3215, 16'd43447, 16'd10603, 16'd15622, 16'd12077, 16'd32938, 16'd41465, 16'd8655, 16'd43077, 16'd46558});
	test_expansion(128'h6be11a38ec84675e5622320b37217dd4, {16'd62715, 16'd19466, 16'd14984, 16'd1399, 16'd18427, 16'd62973, 16'd32336, 16'd16728, 16'd58671, 16'd33490, 16'd45562, 16'd21894, 16'd64947, 16'd24145, 16'd43269, 16'd48034, 16'd5656, 16'd38458, 16'd28419, 16'd34356, 16'd11847, 16'd61615, 16'd60876, 16'd49843, 16'd28790, 16'd6574});
	test_expansion(128'h5199d5daa7f815576517d5d8d132966d, {16'd42606, 16'd16931, 16'd13997, 16'd13321, 16'd26857, 16'd30806, 16'd26261, 16'd62201, 16'd34640, 16'd16290, 16'd34956, 16'd41650, 16'd46325, 16'd62448, 16'd11951, 16'd28514, 16'd878, 16'd34846, 16'd7830, 16'd44006, 16'd5002, 16'd35800, 16'd12220, 16'd16042, 16'd34612, 16'd4855});
	test_expansion(128'h9519aa80075c2b578f9914ae0fc10cc8, {16'd14268, 16'd31767, 16'd5156, 16'd32814, 16'd8209, 16'd24381, 16'd7510, 16'd53565, 16'd27323, 16'd63101, 16'd7648, 16'd38018, 16'd18380, 16'd11498, 16'd57612, 16'd54417, 16'd53516, 16'd49058, 16'd12117, 16'd37779, 16'd12194, 16'd35793, 16'd13349, 16'd40234, 16'd2936, 16'd48206});
	test_expansion(128'h5b612e338fa07f24f35033fed3f6e301, {16'd5092, 16'd55084, 16'd35645, 16'd4441, 16'd18608, 16'd35325, 16'd5227, 16'd39127, 16'd29432, 16'd7526, 16'd39048, 16'd51495, 16'd58298, 16'd30367, 16'd16678, 16'd38200, 16'd18102, 16'd60534, 16'd53872, 16'd54482, 16'd40091, 16'd7134, 16'd45990, 16'd25087, 16'd13567, 16'd10085});
	test_expansion(128'h07b186ac44261de8f6784ece953057bf, {16'd32022, 16'd20018, 16'd7939, 16'd32550, 16'd60415, 16'd55179, 16'd38014, 16'd10252, 16'd7960, 16'd46872, 16'd4084, 16'd6716, 16'd27629, 16'd49241, 16'd8995, 16'd57176, 16'd19962, 16'd46761, 16'd53691, 16'd17, 16'd46444, 16'd32838, 16'd25897, 16'd8802, 16'd38619, 16'd6012});
	test_expansion(128'he654fd419c0109262ae617e8765b8ce3, {16'd10992, 16'd62016, 16'd44908, 16'd55216, 16'd19640, 16'd38770, 16'd64046, 16'd8118, 16'd37863, 16'd35350, 16'd34041, 16'd28045, 16'd60772, 16'd55196, 16'd1374, 16'd60170, 16'd51743, 16'd58237, 16'd18167, 16'd42577, 16'd45434, 16'd44842, 16'd37808, 16'd22059, 16'd53097, 16'd30272});
	test_expansion(128'he060c0026048268bcb77530914a25932, {16'd4963, 16'd63110, 16'd17213, 16'd9682, 16'd22858, 16'd32587, 16'd51025, 16'd34469, 16'd51943, 16'd59972, 16'd29423, 16'd31821, 16'd40248, 16'd38111, 16'd37230, 16'd10806, 16'd60313, 16'd23936, 16'd47405, 16'd45185, 16'd43361, 16'd19841, 16'd42579, 16'd19622, 16'd21074, 16'd27053});
	test_expansion(128'h70020d7653395a6052ff774f5f98908c, {16'd25285, 16'd17524, 16'd21103, 16'd39827, 16'd10729, 16'd11024, 16'd12221, 16'd62247, 16'd46070, 16'd63939, 16'd27570, 16'd21099, 16'd29578, 16'd39325, 16'd42830, 16'd6443, 16'd32166, 16'd48399, 16'd60651, 16'd31816, 16'd22743, 16'd33904, 16'd63841, 16'd25354, 16'd50673, 16'd62835});
	test_expansion(128'hb7f4711cf4dc289aa69bae11022a5775, {16'd49735, 16'd41926, 16'd44314, 16'd24353, 16'd61829, 16'd10898, 16'd4760, 16'd39627, 16'd5702, 16'd11510, 16'd22660, 16'd56576, 16'd27491, 16'd10676, 16'd42948, 16'd46469, 16'd27215, 16'd50835, 16'd11061, 16'd36534, 16'd41876, 16'd9451, 16'd22196, 16'd30444, 16'd50911, 16'd28826});
	test_expansion(128'h08da8e54ae1d608b4648291a136cbccf, {16'd37354, 16'd59164, 16'd30962, 16'd53691, 16'd4031, 16'd51647, 16'd53500, 16'd9059, 16'd19523, 16'd10290, 16'd55994, 16'd57992, 16'd14839, 16'd12901, 16'd27540, 16'd14296, 16'd12094, 16'd11550, 16'd7384, 16'd54944, 16'd3572, 16'd46198, 16'd55560, 16'd53013, 16'd13417, 16'd5467});
	test_expansion(128'h2b24468b2907bec29926898c3e5391d1, {16'd25818, 16'd48667, 16'd53436, 16'd29417, 16'd52197, 16'd28979, 16'd13884, 16'd29921, 16'd8036, 16'd51273, 16'd43094, 16'd63139, 16'd51551, 16'd61252, 16'd5619, 16'd25475, 16'd2719, 16'd42437, 16'd40813, 16'd38418, 16'd30738, 16'd35913, 16'd8476, 16'd12101, 16'd35391, 16'd33451});
	test_expansion(128'he101e3ab74804101fa46d7c41896c2ed, {16'd48254, 16'd42766, 16'd20154, 16'd59846, 16'd60763, 16'd7311, 16'd14605, 16'd6324, 16'd55214, 16'd62102, 16'd46325, 16'd8490, 16'd23132, 16'd32647, 16'd22436, 16'd63169, 16'd50269, 16'd57386, 16'd14037, 16'd41686, 16'd43645, 16'd37141, 16'd15389, 16'd6831, 16'd28292, 16'd18090});
	test_expansion(128'hfa3d273f408bff0a3225afbe517a14b8, {16'd7004, 16'd21837, 16'd50689, 16'd57507, 16'd4281, 16'd49446, 16'd64233, 16'd24786, 16'd47199, 16'd31422, 16'd53565, 16'd44409, 16'd20185, 16'd4535, 16'd33050, 16'd36631, 16'd58259, 16'd453, 16'd37986, 16'd36201, 16'd21498, 16'd61964, 16'd8828, 16'd62617, 16'd45330, 16'd41947});
	test_expansion(128'h667a252de9c9da750ab235ba9c89e893, {16'd15403, 16'd11476, 16'd2227, 16'd39226, 16'd34341, 16'd59217, 16'd17246, 16'd29484, 16'd10007, 16'd2076, 16'd45936, 16'd13317, 16'd11574, 16'd5707, 16'd54779, 16'd8202, 16'd18882, 16'd59108, 16'd26830, 16'd19358, 16'd37831, 16'd27254, 16'd18918, 16'd31390, 16'd44527, 16'd18073});
	test_expansion(128'h14c1f3d0e291efe1ab22a64f0223a415, {16'd13054, 16'd48280, 16'd29301, 16'd34665, 16'd32398, 16'd30747, 16'd55259, 16'd121, 16'd30626, 16'd55890, 16'd27827, 16'd57116, 16'd57013, 16'd47568, 16'd22885, 16'd44686, 16'd41698, 16'd41801, 16'd14364, 16'd61627, 16'd40572, 16'd2675, 16'd16211, 16'd850, 16'd19685, 16'd58161});
	test_expansion(128'hf65b3f6c19d669442bc8efd6a4101303, {16'd19063, 16'd51271, 16'd26529, 16'd2024, 16'd4940, 16'd23146, 16'd38503, 16'd5582, 16'd18798, 16'd35093, 16'd30717, 16'd34296, 16'd7341, 16'd65246, 16'd10083, 16'd64986, 16'd16259, 16'd27046, 16'd50566, 16'd58278, 16'd45831, 16'd906, 16'd47560, 16'd64146, 16'd34727, 16'd16419});
	test_expansion(128'h0557e7ed2408cfe41b442497d093803b, {16'd29203, 16'd65466, 16'd7145, 16'd1154, 16'd63324, 16'd16023, 16'd63078, 16'd9278, 16'd52141, 16'd23257, 16'd61947, 16'd24606, 16'd31058, 16'd18864, 16'd14346, 16'd24620, 16'd37958, 16'd55806, 16'd62642, 16'd2073, 16'd5672, 16'd29472, 16'd7876, 16'd38110, 16'd38137, 16'd45907});
	test_expansion(128'he8d880ea5e90aaa8d414c695a6985616, {16'd8659, 16'd28078, 16'd45903, 16'd7085, 16'd50075, 16'd5118, 16'd24512, 16'd34170, 16'd64314, 16'd64670, 16'd52930, 16'd9511, 16'd29796, 16'd57086, 16'd40287, 16'd12794, 16'd50666, 16'd40643, 16'd27474, 16'd20097, 16'd25676, 16'd54484, 16'd22548, 16'd8199, 16'd23319, 16'd21519});
	test_expansion(128'h35d29ff8ffb37a9c3b2e138dd30b5254, {16'd18951, 16'd22661, 16'd21122, 16'd12930, 16'd16497, 16'd13221, 16'd55905, 16'd59521, 16'd27267, 16'd14227, 16'd22032, 16'd39691, 16'd17731, 16'd51660, 16'd18265, 16'd33368, 16'd42532, 16'd45550, 16'd50690, 16'd26301, 16'd47664, 16'd59767, 16'd45634, 16'd27353, 16'd30211, 16'd46574});
	test_expansion(128'hbf8135909b7242673329af416731f845, {16'd171, 16'd17147, 16'd46627, 16'd65400, 16'd30701, 16'd53337, 16'd45151, 16'd47395, 16'd57051, 16'd58975, 16'd5214, 16'd35036, 16'd9072, 16'd35252, 16'd24238, 16'd36422, 16'd27376, 16'd64404, 16'd61995, 16'd35787, 16'd21263, 16'd64649, 16'd19984, 16'd20816, 16'd53665, 16'd13614});
	test_expansion(128'hce5ac9e5f12db777f3db7b2d77e85ad9, {16'd53776, 16'd53574, 16'd49100, 16'd16088, 16'd50421, 16'd60043, 16'd9192, 16'd41827, 16'd12586, 16'd8459, 16'd25510, 16'd26746, 16'd15764, 16'd7769, 16'd39022, 16'd33926, 16'd17051, 16'd61577, 16'd43321, 16'd41344, 16'd61370, 16'd24056, 16'd13373, 16'd61464, 16'd8171, 16'd60163});
	test_expansion(128'h6bedb1e4177f6086f44e911fad084c18, {16'd65075, 16'd49809, 16'd62029, 16'd7363, 16'd53310, 16'd50328, 16'd44989, 16'd21577, 16'd16556, 16'd51194, 16'd41002, 16'd39554, 16'd35817, 16'd3128, 16'd15255, 16'd41761, 16'd61376, 16'd30040, 16'd1279, 16'd10071, 16'd63067, 16'd21124, 16'd41770, 16'd41592, 16'd19907, 16'd33052});
	test_expansion(128'he7a238a86d01e70b9d3f1035912c5630, {16'd41031, 16'd10915, 16'd53033, 16'd55280, 16'd24267, 16'd50045, 16'd55925, 16'd18429, 16'd20315, 16'd27524, 16'd31367, 16'd11941, 16'd25662, 16'd34892, 16'd46172, 16'd19674, 16'd40239, 16'd43966, 16'd27137, 16'd23962, 16'd26047, 16'd20189, 16'd38739, 16'd102, 16'd23155, 16'd21185});
	test_expansion(128'he941b1a335a2446ee4267db00039d5fa, {16'd37733, 16'd44702, 16'd33890, 16'd31344, 16'd60406, 16'd55514, 16'd54574, 16'd45525, 16'd11713, 16'd21246, 16'd42863, 16'd41620, 16'd64841, 16'd17511, 16'd59738, 16'd58177, 16'd35132, 16'd53199, 16'd49725, 16'd1975, 16'd64035, 16'd57005, 16'd20776, 16'd22637, 16'd15602, 16'd12018});
	test_expansion(128'h840bc121dd7eca04e67a6589ed937eba, {16'd2879, 16'd60677, 16'd52740, 16'd7628, 16'd30117, 16'd18071, 16'd37677, 16'd37326, 16'd64498, 16'd31372, 16'd33003, 16'd43604, 16'd56524, 16'd38293, 16'd56587, 16'd1460, 16'd18971, 16'd54728, 16'd14574, 16'd38431, 16'd10287, 16'd64717, 16'd44769, 16'd49831, 16'd57515, 16'd9859});
	test_expansion(128'haa08fb2ee7a2fd892a9bab829a984047, {16'd64827, 16'd62051, 16'd32978, 16'd61775, 16'd23726, 16'd19596, 16'd8633, 16'd16091, 16'd2138, 16'd51964, 16'd25384, 16'd13812, 16'd61269, 16'd5065, 16'd31155, 16'd52117, 16'd43459, 16'd34781, 16'd37841, 16'd5290, 16'd56445, 16'd20004, 16'd57050, 16'd42780, 16'd40049, 16'd45944});
	test_expansion(128'hd497e8de42c52e514159b404e4d33e29, {16'd23277, 16'd52990, 16'd29591, 16'd63941, 16'd39824, 16'd36330, 16'd30692, 16'd30288, 16'd3350, 16'd4753, 16'd36869, 16'd62546, 16'd20382, 16'd51771, 16'd52250, 16'd35059, 16'd51688, 16'd65406, 16'd15345, 16'd1312, 16'd55302, 16'd24987, 16'd57351, 16'd56691, 16'd37514, 16'd13576});
	test_expansion(128'h45c1dc1ac1982882c2761256fd19132c, {16'd54555, 16'd2184, 16'd40546, 16'd26207, 16'd20983, 16'd45447, 16'd17614, 16'd46903, 16'd28693, 16'd23663, 16'd41962, 16'd8942, 16'd17708, 16'd52239, 16'd31447, 16'd27340, 16'd32980, 16'd6973, 16'd16591, 16'd14888, 16'd1075, 16'd12545, 16'd20617, 16'd24827, 16'd49819, 16'd64167});
	test_expansion(128'h693f2dceba89c64075e66a4e6279fa9c, {16'd46394, 16'd31420, 16'd65016, 16'd24477, 16'd925, 16'd11838, 16'd20165, 16'd13653, 16'd34932, 16'd28816, 16'd20956, 16'd13162, 16'd52413, 16'd38674, 16'd37533, 16'd16447, 16'd48777, 16'd4645, 16'd9299, 16'd57589, 16'd44589, 16'd50697, 16'd64690, 16'd44685, 16'd31884, 16'd31178});
	test_expansion(128'hd638ed0c30d2130e1d6c70e51a0e9181, {16'd1369, 16'd54692, 16'd30468, 16'd34150, 16'd19992, 16'd3294, 16'd50934, 16'd63810, 16'd17125, 16'd14481, 16'd12432, 16'd43780, 16'd3733, 16'd57090, 16'd7892, 16'd43923, 16'd44082, 16'd6115, 16'd47033, 16'd20341, 16'd40943, 16'd55833, 16'd9587, 16'd27160, 16'd47722, 16'd57323});
	test_expansion(128'h5d9c9078360a57d83b81edc2d73a8ea1, {16'd47823, 16'd8934, 16'd25564, 16'd45720, 16'd15998, 16'd19494, 16'd64411, 16'd3118, 16'd2643, 16'd6731, 16'd37320, 16'd17470, 16'd61948, 16'd27555, 16'd9303, 16'd6928, 16'd18734, 16'd44255, 16'd34939, 16'd30293, 16'd17789, 16'd58073, 16'd21051, 16'd35679, 16'd29425, 16'd58704});
	test_expansion(128'h29c5e6d92e70d57850b3d0fb1e72c705, {16'd43408, 16'd57219, 16'd9358, 16'd26948, 16'd45222, 16'd24899, 16'd27625, 16'd30076, 16'd6714, 16'd20123, 16'd9997, 16'd5605, 16'd60975, 16'd58731, 16'd58199, 16'd40722, 16'd64704, 16'd16655, 16'd19355, 16'd35476, 16'd48719, 16'd24360, 16'd36538, 16'd17735, 16'd18985, 16'd11792});
	test_expansion(128'h7427cf7982ddca29fcf7154d82ec4c59, {16'd405, 16'd56272, 16'd36868, 16'd45589, 16'd41128, 16'd9747, 16'd10304, 16'd65257, 16'd40444, 16'd18156, 16'd25982, 16'd53458, 16'd23787, 16'd62572, 16'd25223, 16'd4804, 16'd42717, 16'd28613, 16'd33304, 16'd61200, 16'd55412, 16'd14344, 16'd53135, 16'd44047, 16'd61471, 16'd65176});
	test_expansion(128'h03ae83b3ab9223201e87f6761280bb99, {16'd60922, 16'd23275, 16'd8841, 16'd53815, 16'd19526, 16'd34015, 16'd14740, 16'd50904, 16'd48428, 16'd10418, 16'd35275, 16'd58650, 16'd15371, 16'd1833, 16'd33665, 16'd22137, 16'd51324, 16'd15971, 16'd38433, 16'd49808, 16'd16038, 16'd32111, 16'd18139, 16'd24815, 16'd39540, 16'd36608});
	test_expansion(128'h85a15012e9385053cacb5df30f6ee17d, {16'd7264, 16'd15349, 16'd54061, 16'd52803, 16'd7000, 16'd39018, 16'd50255, 16'd40639, 16'd3349, 16'd52186, 16'd7104, 16'd10874, 16'd51841, 16'd20742, 16'd48197, 16'd21330, 16'd33733, 16'd54218, 16'd218, 16'd4219, 16'd47328, 16'd8173, 16'd32644, 16'd42576, 16'd14155, 16'd57664});
	test_expansion(128'h6d7e03eacd74b09133f2dfd6742de29d, {16'd16008, 16'd5719, 16'd41781, 16'd19182, 16'd4172, 16'd11586, 16'd37528, 16'd7976, 16'd41714, 16'd40891, 16'd4521, 16'd43188, 16'd47254, 16'd56896, 16'd24164, 16'd38890, 16'd24374, 16'd26063, 16'd4756, 16'd41538, 16'd7870, 16'd2357, 16'd53027, 16'd59367, 16'd23656, 16'd5625});
	test_expansion(128'h559a19204f996d337935bbfe97f92144, {16'd29157, 16'd37387, 16'd19628, 16'd15666, 16'd61265, 16'd60640, 16'd965, 16'd15210, 16'd7654, 16'd57931, 16'd22113, 16'd9062, 16'd55243, 16'd17847, 16'd7729, 16'd29202, 16'd13120, 16'd12156, 16'd26171, 16'd24588, 16'd62608, 16'd32712, 16'd60525, 16'd39645, 16'd54854, 16'd616});
	test_expansion(128'ha0e93ddad3729e44c415a07455f51afb, {16'd36454, 16'd31150, 16'd35231, 16'd57020, 16'd6589, 16'd26915, 16'd47331, 16'd23974, 16'd36052, 16'd52699, 16'd27018, 16'd64606, 16'd40777, 16'd33635, 16'd51684, 16'd15572, 16'd10470, 16'd40210, 16'd64780, 16'd60166, 16'd6707, 16'd22895, 16'd39949, 16'd48361, 16'd2949, 16'd47374});
	test_expansion(128'hbc1cdb8a9c25a07724922a2d882f07f0, {16'd4837, 16'd7243, 16'd7618, 16'd49384, 16'd44013, 16'd3557, 16'd34908, 16'd40959, 16'd3190, 16'd36966, 16'd2449, 16'd56914, 16'd11154, 16'd38516, 16'd64016, 16'd60019, 16'd19393, 16'd37951, 16'd50894, 16'd47342, 16'd8662, 16'd54781, 16'd39561, 16'd46698, 16'd13543, 16'd59576});
	test_expansion(128'h694c7b0b3edf62e79ae3664c708b91cc, {16'd20620, 16'd11994, 16'd56074, 16'd40365, 16'd13289, 16'd60842, 16'd10769, 16'd37186, 16'd61849, 16'd12948, 16'd30104, 16'd14112, 16'd36567, 16'd21800, 16'd31415, 16'd59596, 16'd41496, 16'd28304, 16'd24981, 16'd21209, 16'd27227, 16'd23415, 16'd27015, 16'd37723, 16'd36600, 16'd55972});
	test_expansion(128'h43fdb8494fe17adc68ba25c13dc69af2, {16'd28377, 16'd20478, 16'd62264, 16'd46166, 16'd30678, 16'd22968, 16'd5144, 16'd59458, 16'd57042, 16'd52349, 16'd55652, 16'd1059, 16'd7822, 16'd59504, 16'd38795, 16'd5145, 16'd58782, 16'd35278, 16'd59494, 16'd57933, 16'd45776, 16'd10093, 16'd39226, 16'd64878, 16'd12352, 16'd49864});
	test_expansion(128'hda5a4fcc05e6ca1b67825fdb7b1e0130, {16'd26538, 16'd33154, 16'd35196, 16'd56760, 16'd8861, 16'd2285, 16'd1665, 16'd47863, 16'd41748, 16'd1318, 16'd32041, 16'd25455, 16'd43923, 16'd32617, 16'd18137, 16'd42182, 16'd59330, 16'd44242, 16'd47882, 16'd45106, 16'd56839, 16'd44266, 16'd43406, 16'd63884, 16'd489, 16'd7122});
	test_expansion(128'h5659f3eef44f7901d7faeb721a4425d2, {16'd24450, 16'd3149, 16'd51708, 16'd54997, 16'd38431, 16'd48345, 16'd589, 16'd53979, 16'd65051, 16'd46285, 16'd48501, 16'd11399, 16'd11659, 16'd7210, 16'd65124, 16'd49807, 16'd35244, 16'd62081, 16'd58757, 16'd19750, 16'd19211, 16'd50314, 16'd17702, 16'd7554, 16'd46750, 16'd46241});
	test_expansion(128'hadb9788b1b1284a5b1b9ffa9462f1e67, {16'd61735, 16'd10054, 16'd47974, 16'd49304, 16'd53448, 16'd53001, 16'd56584, 16'd29277, 16'd56096, 16'd17573, 16'd31623, 16'd15893, 16'd34133, 16'd22211, 16'd24092, 16'd314, 16'd41279, 16'd388, 16'd42110, 16'd25395, 16'd49515, 16'd18181, 16'd33410, 16'd44878, 16'd36508, 16'd35910});
	test_expansion(128'hc9dcadf82076355d82dc4aadcba8d3c7, {16'd26970, 16'd582, 16'd65426, 16'd8422, 16'd26146, 16'd52378, 16'd61798, 16'd44860, 16'd24945, 16'd53489, 16'd56062, 16'd30637, 16'd64920, 16'd58619, 16'd17891, 16'd36250, 16'd42178, 16'd39461, 16'd27278, 16'd55216, 16'd33846, 16'd64696, 16'd21856, 16'd25877, 16'd65032, 16'd62576});
	test_expansion(128'h9ecdbc71b22fe6e3017ac8fc51e7893c, {16'd57310, 16'd14237, 16'd15695, 16'd41921, 16'd31914, 16'd50918, 16'd33774, 16'd55273, 16'd47532, 16'd27774, 16'd7025, 16'd28710, 16'd35200, 16'd39003, 16'd11372, 16'd61708, 16'd34013, 16'd26354, 16'd61599, 16'd53284, 16'd53567, 16'd17668, 16'd45620, 16'd49787, 16'd62742, 16'd48409});
	test_expansion(128'ha4fce06157b0046a26da11bfc8080510, {16'd30307, 16'd16610, 16'd32174, 16'd7201, 16'd61659, 16'd21651, 16'd26022, 16'd29987, 16'd11042, 16'd1923, 16'd54261, 16'd54302, 16'd60366, 16'd31517, 16'd4641, 16'd25194, 16'd40101, 16'd7761, 16'd25511, 16'd49690, 16'd8800, 16'd34556, 16'd59909, 16'd53011, 16'd56979, 16'd22298});
	test_expansion(128'h7e02fea5a119a74b6078ff931536b429, {16'd13704, 16'd12626, 16'd49194, 16'd28863, 16'd2662, 16'd32810, 16'd25452, 16'd31936, 16'd25738, 16'd27382, 16'd29246, 16'd51457, 16'd41976, 16'd5836, 16'd44863, 16'd21749, 16'd30597, 16'd11568, 16'd14104, 16'd10548, 16'd62220, 16'd65120, 16'd31472, 16'd38440, 16'd465, 16'd27441});
	test_expansion(128'h5b455509089c05539611ecfc67d7a1b6, {16'd29387, 16'd36164, 16'd4030, 16'd50486, 16'd9610, 16'd63181, 16'd4244, 16'd36835, 16'd25, 16'd13589, 16'd47039, 16'd23751, 16'd6912, 16'd43903, 16'd12372, 16'd2335, 16'd57384, 16'd5649, 16'd59689, 16'd16636, 16'd20649, 16'd30782, 16'd43526, 16'd31786, 16'd33286, 16'd15528});
	test_expansion(128'hc651ecbfc8055739d7b0c440e88fe2de, {16'd4941, 16'd60569, 16'd983, 16'd23706, 16'd20424, 16'd12899, 16'd57878, 16'd19584, 16'd64498, 16'd58239, 16'd9250, 16'd6692, 16'd14519, 16'd60362, 16'd8812, 16'd28496, 16'd49107, 16'd59726, 16'd26506, 16'd35222, 16'd6259, 16'd58022, 16'd32921, 16'd207, 16'd52249, 16'd50149});
	test_expansion(128'had749655f8aabcf94f67f2313eb61add, {16'd3586, 16'd65130, 16'd18520, 16'd47377, 16'd64762, 16'd11910, 16'd48783, 16'd10640, 16'd43915, 16'd35581, 16'd26781, 16'd49666, 16'd16200, 16'd59514, 16'd27228, 16'd48296, 16'd39615, 16'd58479, 16'd64783, 16'd31946, 16'd4298, 16'd24567, 16'd3304, 16'd40042, 16'd13701, 16'd43628});
	test_expansion(128'hb20552cfb6aac35a5a6ce153029aa23b, {16'd45850, 16'd50266, 16'd57902, 16'd50941, 16'd47840, 16'd54324, 16'd3558, 16'd23158, 16'd64428, 16'd40662, 16'd11063, 16'd24074, 16'd57118, 16'd63610, 16'd15067, 16'd19121, 16'd26754, 16'd28008, 16'd11580, 16'd12233, 16'd10329, 16'd62368, 16'd3330, 16'd48823, 16'd6992, 16'd26185});
	test_expansion(128'h229e1f1cf4fe01ac77af50d39546238f, {16'd56153, 16'd41521, 16'd18902, 16'd42408, 16'd48640, 16'd12544, 16'd35413, 16'd61786, 16'd46114, 16'd17028, 16'd55505, 16'd38716, 16'd36458, 16'd51085, 16'd63737, 16'd32313, 16'd55536, 16'd2997, 16'd47498, 16'd8032, 16'd52268, 16'd18252, 16'd1993, 16'd42094, 16'd28001, 16'd51575});
	test_expansion(128'hafa264c6f88cf86b4711e0b6a4bb219b, {16'd10504, 16'd52483, 16'd58932, 16'd20177, 16'd1113, 16'd22053, 16'd57620, 16'd61918, 16'd55219, 16'd9796, 16'd13286, 16'd33345, 16'd41219, 16'd17453, 16'd26848, 16'd43643, 16'd19597, 16'd12972, 16'd64948, 16'd55722, 16'd25362, 16'd28030, 16'd54449, 16'd52506, 16'd6010, 16'd23175});
	test_expansion(128'hf5fc8ae2eebe643994c513f85fe9f363, {16'd22901, 16'd18005, 16'd57951, 16'd36412, 16'd54975, 16'd25559, 16'd6344, 16'd27289, 16'd5047, 16'd57410, 16'd618, 16'd1148, 16'd44916, 16'd5536, 16'd21472, 16'd15844, 16'd3701, 16'd58676, 16'd62219, 16'd62001, 16'd43047, 16'd38539, 16'd44913, 16'd38248, 16'd9830, 16'd62416});
	test_expansion(128'hda179d9ae8f7b0970bcb55f689d8d3b5, {16'd7629, 16'd18807, 16'd25991, 16'd63274, 16'd22716, 16'd39199, 16'd60028, 16'd12505, 16'd16915, 16'd49, 16'd38864, 16'd25731, 16'd10981, 16'd4609, 16'd14124, 16'd60748, 16'd10892, 16'd35676, 16'd942, 16'd33868, 16'd54981, 16'd33619, 16'd56099, 16'd27168, 16'd29021, 16'd50025});
	test_expansion(128'h1c8b67f41aae9f91229b4e6f6e9a5c29, {16'd43689, 16'd46342, 16'd36391, 16'd36456, 16'd59669, 16'd13239, 16'd168, 16'd19591, 16'd53372, 16'd46642, 16'd29599, 16'd47926, 16'd29786, 16'd49215, 16'd2343, 16'd48822, 16'd1885, 16'd15961, 16'd56020, 16'd21094, 16'd29789, 16'd24843, 16'd48560, 16'd1620, 16'd9141, 16'd33175});
	test_expansion(128'hec3516a3b892e05a00312e324615048d, {16'd3635, 16'd25198, 16'd2523, 16'd57799, 16'd19729, 16'd45819, 16'd42215, 16'd12783, 16'd30161, 16'd57607, 16'd41700, 16'd33897, 16'd13656, 16'd10199, 16'd43112, 16'd32278, 16'd24123, 16'd52288, 16'd63812, 16'd18443, 16'd45446, 16'd18688, 16'd26833, 16'd24187, 16'd28840, 16'd49588});
	test_expansion(128'hea9d47b948a8d9e082667132c1232105, {16'd35460, 16'd47509, 16'd35164, 16'd29783, 16'd63174, 16'd44234, 16'd5065, 16'd57913, 16'd26677, 16'd1025, 16'd44882, 16'd9749, 16'd32983, 16'd22973, 16'd30672, 16'd54239, 16'd3278, 16'd58228, 16'd39007, 16'd59712, 16'd51982, 16'd1438, 16'd14233, 16'd58205, 16'd22471, 16'd45793});
	test_expansion(128'h1cfe8f89a250f604f9079d3d4d3b6a3c, {16'd45690, 16'd52999, 16'd21219, 16'd4735, 16'd64866, 16'd2260, 16'd44800, 16'd30337, 16'd53067, 16'd55515, 16'd19097, 16'd28400, 16'd18163, 16'd38175, 16'd42534, 16'd14896, 16'd15672, 16'd52909, 16'd37923, 16'd42983, 16'd47029, 16'd5711, 16'd31651, 16'd64458, 16'd57881, 16'd1990});
	test_expansion(128'he76d773d780755e42fb1d0951755c9de, {16'd26725, 16'd42948, 16'd44596, 16'd18133, 16'd1419, 16'd52740, 16'd34313, 16'd48856, 16'd1268, 16'd16180, 16'd30357, 16'd41440, 16'd64160, 16'd56804, 16'd60613, 16'd15028, 16'd10430, 16'd23891, 16'd27029, 16'd42997, 16'd20494, 16'd3696, 16'd17637, 16'd62072, 16'd31706, 16'd3600});
	test_expansion(128'h9722c6b8b1ed9f4d8f4c7bb3f62a5d37, {16'd9382, 16'd6563, 16'd49434, 16'd5242, 16'd5700, 16'd16686, 16'd62527, 16'd11290, 16'd13885, 16'd8420, 16'd228, 16'd19697, 16'd3525, 16'd51098, 16'd15141, 16'd25030, 16'd60505, 16'd58181, 16'd13414, 16'd32374, 16'd19002, 16'd33504, 16'd12790, 16'd5580, 16'd6285, 16'd40871});
	test_expansion(128'h4b19315f6c0d7a5a8918fc5f36f5caba, {16'd51154, 16'd54548, 16'd63339, 16'd28353, 16'd17215, 16'd16308, 16'd49912, 16'd28702, 16'd1587, 16'd44248, 16'd28583, 16'd58722, 16'd4448, 16'd64531, 16'd33814, 16'd17974, 16'd42333, 16'd42924, 16'd60725, 16'd25993, 16'd58319, 16'd57768, 16'd17343, 16'd11024, 16'd19080, 16'd41932});
	test_expansion(128'h69bb1675497a918f862a4dd688f8d511, {16'd38065, 16'd65123, 16'd11083, 16'd46515, 16'd49645, 16'd48807, 16'd3626, 16'd1825, 16'd27880, 16'd41802, 16'd15921, 16'd52640, 16'd38926, 16'd32134, 16'd47778, 16'd27027, 16'd17363, 16'd34827, 16'd59396, 16'd47338, 16'd31877, 16'd51504, 16'd40093, 16'd14159, 16'd61527, 16'd58841});
	test_expansion(128'h8d702f73078e096363607ab349beacf6, {16'd36491, 16'd6711, 16'd23731, 16'd26592, 16'd26795, 16'd23059, 16'd2188, 16'd59984, 16'd10671, 16'd56141, 16'd18403, 16'd40248, 16'd20855, 16'd11694, 16'd63544, 16'd54225, 16'd26081, 16'd42309, 16'd13855, 16'd37964, 16'd7212, 16'd17574, 16'd28739, 16'd43912, 16'd37582, 16'd36152});
	test_expansion(128'h7d49eac7c9c2751092e62b228a1eff08, {16'd42818, 16'd25130, 16'd53992, 16'd11447, 16'd39618, 16'd39105, 16'd14610, 16'd12461, 16'd17470, 16'd20641, 16'd23811, 16'd34082, 16'd28302, 16'd29967, 16'd13631, 16'd51230, 16'd34285, 16'd42261, 16'd19827, 16'd23399, 16'd49841, 16'd26896, 16'd9400, 16'd55153, 16'd45548, 16'd48402});
	test_expansion(128'h0df05caa44543e7055430acee0c0a4ef, {16'd2040, 16'd52764, 16'd27101, 16'd61442, 16'd18756, 16'd32266, 16'd46689, 16'd479, 16'd9842, 16'd28205, 16'd14077, 16'd10397, 16'd14355, 16'd33018, 16'd8612, 16'd64018, 16'd18951, 16'd1246, 16'd42204, 16'd32702, 16'd25410, 16'd22227, 16'd35703, 16'd44507, 16'd43435, 16'd35235});
	test_expansion(128'h9522782fd694a6bb3284ba1409ca0b46, {16'd8886, 16'd7590, 16'd24332, 16'd58027, 16'd63242, 16'd15101, 16'd2434, 16'd43903, 16'd21050, 16'd32910, 16'd42320, 16'd60620, 16'd43183, 16'd34476, 16'd18687, 16'd38451, 16'd41863, 16'd24618, 16'd3394, 16'd46611, 16'd40012, 16'd4350, 16'd62842, 16'd65001, 16'd12407, 16'd48895});
	test_expansion(128'h6ce00f666e2dd249562e3559686c3717, {16'd6532, 16'd12258, 16'd37583, 16'd35960, 16'd12208, 16'd44746, 16'd4045, 16'd28515, 16'd63963, 16'd57354, 16'd10499, 16'd13963, 16'd53445, 16'd58375, 16'd24715, 16'd18173, 16'd29308, 16'd38167, 16'd19720, 16'd57662, 16'd37416, 16'd18283, 16'd41450, 16'd38290, 16'd5408, 16'd16109});
	test_expansion(128'hdd5fec11aa4e808958dcf151d5f30716, {16'd26387, 16'd43480, 16'd62412, 16'd47565, 16'd8953, 16'd59432, 16'd16376, 16'd54292, 16'd52263, 16'd64359, 16'd30546, 16'd57647, 16'd22717, 16'd18890, 16'd18124, 16'd44850, 16'd37794, 16'd45410, 16'd56988, 16'd33135, 16'd41751, 16'd14844, 16'd37266, 16'd49746, 16'd906, 16'd16318});
	test_expansion(128'hc93b517a7c5d692bc8c2e60bf11bf504, {16'd46299, 16'd7691, 16'd59435, 16'd30916, 16'd43712, 16'd11698, 16'd28353, 16'd4624, 16'd7846, 16'd58146, 16'd2297, 16'd50922, 16'd573, 16'd50013, 16'd61456, 16'd11563, 16'd60737, 16'd64245, 16'd57575, 16'd26175, 16'd32464, 16'd16978, 16'd17224, 16'd7946, 16'd47280, 16'd30713});
	test_expansion(128'h08dbd6cb2816d964d64876189d5f7338, {16'd7973, 16'd26935, 16'd33058, 16'd39512, 16'd61607, 16'd35620, 16'd43474, 16'd33118, 16'd38066, 16'd42394, 16'd58995, 16'd28472, 16'd54177, 16'd28996, 16'd31349, 16'd22008, 16'd28363, 16'd34683, 16'd17963, 16'd36336, 16'd48091, 16'd5130, 16'd45525, 16'd49591, 16'd32995, 16'd45927});
	test_expansion(128'h4d7b6525fea32773ef6be114f7d0a795, {16'd27100, 16'd56987, 16'd57737, 16'd60112, 16'd24778, 16'd4197, 16'd52378, 16'd14287, 16'd5878, 16'd14776, 16'd29479, 16'd42908, 16'd51595, 16'd29382, 16'd45824, 16'd53904, 16'd11801, 16'd28126, 16'd33100, 16'd29493, 16'd19935, 16'd41606, 16'd31789, 16'd1286, 16'd54685, 16'd12279});
	test_expansion(128'h089b2e24a8e10d8cbae5051345c60ce6, {16'd38068, 16'd38960, 16'd23828, 16'd11460, 16'd29196, 16'd42089, 16'd33412, 16'd58751, 16'd21804, 16'd7894, 16'd35803, 16'd14886, 16'd46483, 16'd29298, 16'd21228, 16'd35385, 16'd63274, 16'd60221, 16'd64453, 16'd60506, 16'd57422, 16'd24674, 16'd19498, 16'd54674, 16'd2237, 16'd12971});
	test_expansion(128'h6e97e9e530658891632806fc86119f19, {16'd23525, 16'd37619, 16'd5006, 16'd4769, 16'd2784, 16'd54226, 16'd16529, 16'd46738, 16'd59954, 16'd22465, 16'd46744, 16'd8313, 16'd27985, 16'd41160, 16'd39873, 16'd39014, 16'd47777, 16'd13681, 16'd55797, 16'd63200, 16'd15097, 16'd12489, 16'd4750, 16'd60649, 16'd9725, 16'd27823});
	test_expansion(128'he3ef35c7aa504d79e04add5bd6ddf369, {16'd42449, 16'd1608, 16'd56283, 16'd35456, 16'd36963, 16'd50852, 16'd34165, 16'd53999, 16'd12466, 16'd5635, 16'd27300, 16'd43069, 16'd52939, 16'd32396, 16'd53427, 16'd7633, 16'd43334, 16'd54385, 16'd26537, 16'd21569, 16'd49932, 16'd39891, 16'd16454, 16'd14387, 16'd15943, 16'd42659});
	test_expansion(128'hb1e732e29d595a156cebd7386e3c0442, {16'd21741, 16'd17774, 16'd21416, 16'd20430, 16'd3470, 16'd52670, 16'd59829, 16'd36621, 16'd26616, 16'd32518, 16'd4880, 16'd37063, 16'd19331, 16'd27135, 16'd26163, 16'd5403, 16'd32898, 16'd51636, 16'd60591, 16'd44599, 16'd35743, 16'd49518, 16'd28529, 16'd26805, 16'd27303, 16'd12316});
	test_expansion(128'hdced4b07082241ff85c443f401e03bea, {16'd17724, 16'd44026, 16'd11753, 16'd22642, 16'd19082, 16'd54247, 16'd58663, 16'd42125, 16'd47630, 16'd62284, 16'd62395, 16'd19211, 16'd42436, 16'd62332, 16'd11910, 16'd49214, 16'd37839, 16'd8921, 16'd5317, 16'd51365, 16'd62937, 16'd39071, 16'd51843, 16'd318, 16'd12599, 16'd43550});
	test_expansion(128'h39ce284bd8d2852f9b3d466f2280fed7, {16'd3130, 16'd64652, 16'd19567, 16'd43042, 16'd6541, 16'd57939, 16'd59546, 16'd32144, 16'd58880, 16'd62168, 16'd42662, 16'd25038, 16'd45535, 16'd31044, 16'd62804, 16'd7352, 16'd18530, 16'd36394, 16'd45513, 16'd4930, 16'd35730, 16'd23813, 16'd26861, 16'd19959, 16'd51174, 16'd38297});
	test_expansion(128'h43fbcce23eab78929b8f089ab46a5ff1, {16'd65492, 16'd33300, 16'd47748, 16'd55959, 16'd52689, 16'd53254, 16'd39456, 16'd54758, 16'd59639, 16'd26320, 16'd56053, 16'd41933, 16'd28596, 16'd15775, 16'd19066, 16'd57251, 16'd52852, 16'd47867, 16'd64120, 16'd8871, 16'd21115, 16'd40549, 16'd57077, 16'd22872, 16'd40872, 16'd243});
	test_expansion(128'h3206577a2b52fcaa9cb8758be5984f0d, {16'd48445, 16'd1930, 16'd21866, 16'd7671, 16'd3711, 16'd36479, 16'd20191, 16'd14002, 16'd18691, 16'd17511, 16'd13251, 16'd56908, 16'd35073, 16'd22794, 16'd16532, 16'd5835, 16'd11349, 16'd57063, 16'd39103, 16'd10710, 16'd44853, 16'd31933, 16'd42962, 16'd19895, 16'd27882, 16'd25047});
	test_expansion(128'h84f21e092c7caa56ccdef7107fbbbea6, {16'd29156, 16'd40834, 16'd16318, 16'd43613, 16'd31335, 16'd58029, 16'd59190, 16'd1811, 16'd15551, 16'd49958, 16'd63000, 16'd29083, 16'd36200, 16'd10964, 16'd32898, 16'd40610, 16'd35312, 16'd14225, 16'd36255, 16'd22219, 16'd28414, 16'd33974, 16'd16174, 16'd475, 16'd44645, 16'd64295});
	test_expansion(128'he03d0e41e70810494105457b4efc85e2, {16'd33831, 16'd8058, 16'd23539, 16'd62120, 16'd18067, 16'd5170, 16'd60911, 16'd29742, 16'd57103, 16'd1227, 16'd13415, 16'd23674, 16'd57892, 16'd11049, 16'd51827, 16'd11361, 16'd998, 16'd2880, 16'd13600, 16'd26468, 16'd35866, 16'd9242, 16'd45405, 16'd15515, 16'd63593, 16'd42376});
	test_expansion(128'haefbba0ed8a502b448db954f2beed877, {16'd49434, 16'd45544, 16'd29332, 16'd27922, 16'd19745, 16'd9811, 16'd21872, 16'd15856, 16'd8101, 16'd47347, 16'd37467, 16'd37567, 16'd7512, 16'd3944, 16'd27998, 16'd57232, 16'd22134, 16'd21186, 16'd11758, 16'd14591, 16'd38820, 16'd18133, 16'd14441, 16'd45131, 16'd30280, 16'd3372});
	test_expansion(128'h7afaa36004a2671b0393a2679266d4fd, {16'd45075, 16'd62605, 16'd26170, 16'd23013, 16'd57253, 16'd46034, 16'd22327, 16'd1494, 16'd4300, 16'd51544, 16'd8646, 16'd32366, 16'd50008, 16'd63647, 16'd40680, 16'd48010, 16'd58926, 16'd42113, 16'd57994, 16'd12069, 16'd28651, 16'd59714, 16'd4726, 16'd9186, 16'd21214, 16'd29409});
	test_expansion(128'ha2ccae28a15148e5970c76f6e63c93ac, {16'd48387, 16'd30534, 16'd47638, 16'd36025, 16'd14028, 16'd25676, 16'd51966, 16'd41366, 16'd1064, 16'd64195, 16'd9578, 16'd2901, 16'd46406, 16'd63250, 16'd15098, 16'd54108, 16'd15623, 16'd61598, 16'd19192, 16'd53213, 16'd56146, 16'd55727, 16'd52123, 16'd3471, 16'd24355, 16'd25350});
	test_expansion(128'h26943ac87fe16c7bd9a0870772cec774, {16'd17636, 16'd14116, 16'd51187, 16'd32576, 16'd45371, 16'd5866, 16'd58140, 16'd51061, 16'd62015, 16'd14866, 16'd40860, 16'd13981, 16'd59124, 16'd17274, 16'd55759, 16'd47477, 16'd45505, 16'd13333, 16'd13718, 16'd36175, 16'd5869, 16'd12974, 16'd14879, 16'd14448, 16'd29668, 16'd50446});
	test_expansion(128'hc0b397ac11602b80354b86b5d1b4c4ae, {16'd26962, 16'd2279, 16'd15907, 16'd9746, 16'd61600, 16'd2213, 16'd53513, 16'd11856, 16'd59862, 16'd39010, 16'd51523, 16'd33297, 16'd48484, 16'd10221, 16'd30375, 16'd24681, 16'd25948, 16'd22934, 16'd34412, 16'd10919, 16'd2333, 16'd50349, 16'd4448, 16'd54621, 16'd20932, 16'd54119});
	test_expansion(128'he400584862cf33170aef6348f2284455, {16'd7162, 16'd6757, 16'd12438, 16'd33816, 16'd42271, 16'd6550, 16'd1716, 16'd53574, 16'd35785, 16'd4624, 16'd50530, 16'd39270, 16'd11643, 16'd27246, 16'd27894, 16'd59633, 16'd49583, 16'd12450, 16'd57800, 16'd27626, 16'd6908, 16'd29845, 16'd49589, 16'd1367, 16'd16994, 16'd57373});
	test_expansion(128'hee6d51a2d025895f7f1dafc50985d12a, {16'd9448, 16'd59057, 16'd38868, 16'd13464, 16'd16142, 16'd56437, 16'd51692, 16'd49728, 16'd55109, 16'd4534, 16'd25443, 16'd17846, 16'd64831, 16'd6216, 16'd13933, 16'd1818, 16'd46907, 16'd34304, 16'd44564, 16'd4896, 16'd3735, 16'd57078, 16'd18269, 16'd48237, 16'd55500, 16'd53609});
	test_expansion(128'h8305c7cea8c897bbf9d19094e02e2638, {16'd64831, 16'd20444, 16'd23930, 16'd54058, 16'd2454, 16'd20473, 16'd52252, 16'd41067, 16'd17834, 16'd31016, 16'd42893, 16'd5364, 16'd26481, 16'd44094, 16'd17955, 16'd62866, 16'd39329, 16'd45509, 16'd64019, 16'd14017, 16'd65109, 16'd25021, 16'd12214, 16'd54768, 16'd33742, 16'd13570});
	test_expansion(128'hf995ba1f7fa82a425b0fd41b5f4a9692, {16'd58151, 16'd22513, 16'd19497, 16'd30562, 16'd42849, 16'd38235, 16'd61556, 16'd9749, 16'd14484, 16'd65372, 16'd11193, 16'd32309, 16'd33992, 16'd59788, 16'd53277, 16'd49724, 16'd48474, 16'd19723, 16'd6812, 16'd54773, 16'd54378, 16'd14745, 16'd64786, 16'd63329, 16'd19183, 16'd11923});
	test_expansion(128'h8d7644a9b4d7face7b14a4481ef64826, {16'd7151, 16'd49785, 16'd24638, 16'd36921, 16'd33622, 16'd43666, 16'd4734, 16'd50748, 16'd45274, 16'd46443, 16'd56219, 16'd34994, 16'd13997, 16'd8536, 16'd13553, 16'd41284, 16'd40811, 16'd54422, 16'd586, 16'd35761, 16'd31659, 16'd11582, 16'd2592, 16'd14887, 16'd49152, 16'd39737});
	test_expansion(128'h1a130d1a4a4a1cbf33b2d477556f0623, {16'd16276, 16'd39426, 16'd1207, 16'd57740, 16'd45911, 16'd31011, 16'd6289, 16'd38293, 16'd23587, 16'd18755, 16'd37445, 16'd64513, 16'd33826, 16'd41773, 16'd15400, 16'd59476, 16'd32338, 16'd25902, 16'd8948, 16'd14665, 16'd28500, 16'd22238, 16'd37289, 16'd50351, 16'd44567, 16'd30218});
	test_expansion(128'h1375bc6b9596c84e076cb04ced475bc0, {16'd27890, 16'd26626, 16'd30628, 16'd5649, 16'd730, 16'd5759, 16'd12340, 16'd48408, 16'd3156, 16'd54272, 16'd49518, 16'd4081, 16'd27480, 16'd52892, 16'd4247, 16'd3439, 16'd7835, 16'd26694, 16'd3570, 16'd43578, 16'd30066, 16'd4736, 16'd37252, 16'd57557, 16'd59061, 16'd35354});
	test_expansion(128'hc91df95a8a43b5cd217e40520bda351e, {16'd59160, 16'd2074, 16'd16610, 16'd12259, 16'd27505, 16'd911, 16'd52430, 16'd62124, 16'd5548, 16'd64858, 16'd19062, 16'd24751, 16'd45745, 16'd23200, 16'd12443, 16'd11897, 16'd18324, 16'd36951, 16'd4701, 16'd40032, 16'd7780, 16'd42375, 16'd14332, 16'd22959, 16'd25568, 16'd30569});
	test_expansion(128'h3e1bfc8c80e7667108e99ea0395eafef, {16'd54760, 16'd18250, 16'd913, 16'd12388, 16'd20850, 16'd46198, 16'd29953, 16'd19516, 16'd9920, 16'd3312, 16'd23025, 16'd57163, 16'd32134, 16'd63909, 16'd11327, 16'd5745, 16'd30519, 16'd50809, 16'd50971, 16'd707, 16'd47812, 16'd65523, 16'd21871, 16'd38895, 16'd39213, 16'd48246});
	test_expansion(128'he447e889e8a5b708423064c6d655fb42, {16'd32912, 16'd65091, 16'd253, 16'd9512, 16'd2757, 16'd27306, 16'd26539, 16'd25509, 16'd45389, 16'd3481, 16'd13635, 16'd26945, 16'd49706, 16'd31803, 16'd12973, 16'd33801, 16'd738, 16'd15754, 16'd43773, 16'd58830, 16'd54865, 16'd45559, 16'd44183, 16'd30558, 16'd58348, 16'd40894});
	test_expansion(128'hc12d049429fda6ce7b95006eb4306c91, {16'd35356, 16'd19911, 16'd32995, 16'd13212, 16'd39725, 16'd48474, 16'd50470, 16'd60245, 16'd33654, 16'd52277, 16'd35454, 16'd2337, 16'd10525, 16'd49727, 16'd9891, 16'd42811, 16'd20717, 16'd4888, 16'd56431, 16'd57693, 16'd56130, 16'd7438, 16'd51410, 16'd55059, 16'd46781, 16'd18940});
	test_expansion(128'hcd3cec8c707d16d50450fafa37603930, {16'd24251, 16'd50664, 16'd58435, 16'd21833, 16'd37241, 16'd1888, 16'd54135, 16'd46182, 16'd59492, 16'd45464, 16'd5633, 16'd62582, 16'd22600, 16'd26242, 16'd35150, 16'd46069, 16'd23577, 16'd26112, 16'd22147, 16'd33022, 16'd52999, 16'd23747, 16'd33050, 16'd11626, 16'd24485, 16'd46763});
	test_expansion(128'h716f1c214e2a053ce83f484eba38ddbe, {16'd4246, 16'd52123, 16'd21937, 16'd27902, 16'd59766, 16'd13886, 16'd21724, 16'd37796, 16'd47902, 16'd21450, 16'd9121, 16'd55142, 16'd38354, 16'd22003, 16'd32230, 16'd50562, 16'd33441, 16'd60283, 16'd26051, 16'd33041, 16'd53806, 16'd31342, 16'd26208, 16'd55538, 16'd43884, 16'd53907});
	test_expansion(128'h32b334658ab2885cd57be157d1dc1944, {16'd47526, 16'd60342, 16'd50682, 16'd20635, 16'd55576, 16'd59626, 16'd850, 16'd22763, 16'd35347, 16'd270, 16'd21682, 16'd63258, 16'd59194, 16'd12921, 16'd63806, 16'd59582, 16'd31165, 16'd43148, 16'd21226, 16'd7531, 16'd58781, 16'd22246, 16'd64621, 16'd56104, 16'd36070, 16'd19328});
	test_expansion(128'h8c1973ada33331c586a59b8fd60cb298, {16'd54028, 16'd60730, 16'd44389, 16'd11014, 16'd51242, 16'd23478, 16'd39580, 16'd52813, 16'd47345, 16'd3363, 16'd21861, 16'd20657, 16'd60911, 16'd16274, 16'd16315, 16'd1402, 16'd24598, 16'd50802, 16'd7512, 16'd59981, 16'd59981, 16'd31658, 16'd8215, 16'd16765, 16'd47554, 16'd56547});
	test_expansion(128'h0fd814a5a3a7fa003ac19d786c46227a, {16'd24576, 16'd49663, 16'd1237, 16'd11843, 16'd37787, 16'd58251, 16'd8518, 16'd41540, 16'd10239, 16'd18508, 16'd29175, 16'd15630, 16'd12504, 16'd54381, 16'd64798, 16'd8241, 16'd34780, 16'd48333, 16'd22335, 16'd28911, 16'd27580, 16'd45649, 16'd19333, 16'd2522, 16'd48285, 16'd20124});
	test_expansion(128'he392850cda34901fb6d66c62c39a9d9f, {16'd16210, 16'd36687, 16'd39428, 16'd62845, 16'd26245, 16'd56800, 16'd28542, 16'd38894, 16'd894, 16'd56851, 16'd39890, 16'd40099, 16'd54614, 16'd39448, 16'd58888, 16'd25802, 16'd64913, 16'd49481, 16'd31228, 16'd48394, 16'd57239, 16'd15154, 16'd17794, 16'd30077, 16'd9418, 16'd3670});
	test_expansion(128'h99ebbf275ab1e7c7b3def1e60a866e90, {16'd3171, 16'd29285, 16'd63749, 16'd24938, 16'd35015, 16'd61058, 16'd64770, 16'd19661, 16'd18407, 16'd29184, 16'd60207, 16'd44568, 16'd27069, 16'd63573, 16'd22831, 16'd13498, 16'd57673, 16'd50993, 16'd8774, 16'd8894, 16'd33010, 16'd40895, 16'd57920, 16'd28092, 16'd55808, 16'd19817});
	test_expansion(128'h40f88cf2508f86c1e18508e909ef6f70, {16'd10891, 16'd40004, 16'd31176, 16'd111, 16'd32695, 16'd14660, 16'd50283, 16'd11443, 16'd56520, 16'd9822, 16'd1085, 16'd57934, 16'd31460, 16'd52292, 16'd46732, 16'd37427, 16'd7032, 16'd44525, 16'd46992, 16'd722, 16'd58253, 16'd51591, 16'd39468, 16'd3073, 16'd41985, 16'd42058});
	test_expansion(128'hb8d3124d564ca29684e6301322d10ef5, {16'd25296, 16'd38564, 16'd27776, 16'd18555, 16'd14100, 16'd43438, 16'd40815, 16'd1876, 16'd53909, 16'd45029, 16'd11648, 16'd28041, 16'd20901, 16'd55996, 16'd2434, 16'd43112, 16'd41968, 16'd30970, 16'd57942, 16'd18531, 16'd24069, 16'd60606, 16'd5347, 16'd29958, 16'd64399, 16'd52527});
	test_expansion(128'hba3ca2450e249252a01691ddeabe7cd4, {16'd49, 16'd46651, 16'd33586, 16'd45871, 16'd35271, 16'd59862, 16'd36381, 16'd63757, 16'd44869, 16'd53763, 16'd52928, 16'd46261, 16'd43031, 16'd15024, 16'd37844, 16'd46180, 16'd2017, 16'd56185, 16'd62056, 16'd11414, 16'd40515, 16'd28788, 16'd52318, 16'd23337, 16'd40908, 16'd11270});
	test_expansion(128'hbc042a7743b76e11d8fc09fdf75863c0, {16'd32464, 16'd34359, 16'd52474, 16'd23949, 16'd29972, 16'd41617, 16'd49762, 16'd23950, 16'd56512, 16'd45353, 16'd41449, 16'd49299, 16'd22771, 16'd58138, 16'd58502, 16'd34377, 16'd61243, 16'd35029, 16'd62716, 16'd41680, 16'd10696, 16'd16942, 16'd54918, 16'd30745, 16'd48057, 16'd27726});
	test_expansion(128'h2347f2ab78afa6d07bf2e41ef0f81e1b, {16'd173, 16'd4405, 16'd47298, 16'd9420, 16'd45718, 16'd32973, 16'd17574, 16'd42794, 16'd19265, 16'd31511, 16'd37760, 16'd43918, 16'd31560, 16'd45991, 16'd11471, 16'd26313, 16'd29257, 16'd58120, 16'd34414, 16'd37049, 16'd48144, 16'd7525, 16'd50041, 16'd58609, 16'd44388, 16'd46948});
	test_expansion(128'h9ba9a54cb86078b23c3c573ac68bafb4, {16'd63589, 16'd8103, 16'd56593, 16'd8121, 16'd32074, 16'd61654, 16'd8669, 16'd63202, 16'd36938, 16'd16099, 16'd36789, 16'd85, 16'd23332, 16'd22923, 16'd47630, 16'd44072, 16'd26189, 16'd60575, 16'd54621, 16'd59458, 16'd585, 16'd42769, 16'd11492, 16'd44635, 16'd18522, 16'd12988});
	test_expansion(128'hb4bd67ffe846235481908784ed47f4ba, {16'd61741, 16'd14531, 16'd46727, 16'd52898, 16'd2912, 16'd6992, 16'd37470, 16'd11449, 16'd10474, 16'd20406, 16'd6553, 16'd46034, 16'd27577, 16'd17993, 16'd35352, 16'd10226, 16'd10127, 16'd16094, 16'd55561, 16'd13549, 16'd26377, 16'd57768, 16'd23170, 16'd45481, 16'd12690, 16'd10237});
	test_expansion(128'hc519c38b88bb4e43601eb80d002e5313, {16'd17255, 16'd54744, 16'd3535, 16'd43221, 16'd52387, 16'd53132, 16'd31906, 16'd18591, 16'd56702, 16'd57313, 16'd48563, 16'd15481, 16'd11268, 16'd34142, 16'd39233, 16'd63018, 16'd12805, 16'd150, 16'd15871, 16'd8779, 16'd3448, 16'd12466, 16'd46100, 16'd10421, 16'd27189, 16'd1141});
	test_expansion(128'h377ad6278cf0dfa9df7766801797da48, {16'd53323, 16'd36713, 16'd5603, 16'd62816, 16'd7739, 16'd62410, 16'd221, 16'd55072, 16'd45961, 16'd15391, 16'd32511, 16'd57171, 16'd25532, 16'd11249, 16'd58090, 16'd29675, 16'd62215, 16'd61096, 16'd33914, 16'd42101, 16'd19703, 16'd16509, 16'd20085, 16'd47434, 16'd11393, 16'd48374});
	test_expansion(128'h6e733fce9d83eafa0b07e4049b375435, {16'd34099, 16'd21722, 16'd54861, 16'd47109, 16'd23418, 16'd12247, 16'd23268, 16'd61837, 16'd29685, 16'd22179, 16'd43736, 16'd3564, 16'd64356, 16'd5097, 16'd31104, 16'd51583, 16'd5918, 16'd31158, 16'd59310, 16'd64168, 16'd10853, 16'd13439, 16'd60992, 16'd11178, 16'd26374, 16'd34964});
	test_expansion(128'h50a96ae802942a8cc4114d65ea921390, {16'd36229, 16'd60569, 16'd21938, 16'd487, 16'd11448, 16'd12402, 16'd15199, 16'd14505, 16'd13629, 16'd12151, 16'd56078, 16'd44779, 16'd43647, 16'd9079, 16'd28758, 16'd48322, 16'd11455, 16'd50214, 16'd18048, 16'd3522, 16'd17980, 16'd7071, 16'd56615, 16'd39811, 16'd56970, 16'd21888});
	test_expansion(128'h9b47a2839a9f9fab99450357eafab570, {16'd45807, 16'd50520, 16'd3520, 16'd47625, 16'd16406, 16'd28672, 16'd26536, 16'd51332, 16'd11106, 16'd23960, 16'd7307, 16'd61046, 16'd9115, 16'd13083, 16'd10291, 16'd6519, 16'd57446, 16'd49369, 16'd42582, 16'd37868, 16'd3228, 16'd17355, 16'd10850, 16'd27928, 16'd54402, 16'd53382});
	test_expansion(128'h2f0356c35eee327272e17e547bfc0353, {16'd22869, 16'd25014, 16'd21358, 16'd17816, 16'd53264, 16'd7337, 16'd53258, 16'd60356, 16'd46687, 16'd49471, 16'd44541, 16'd3885, 16'd19584, 16'd38803, 16'd51892, 16'd26132, 16'd7938, 16'd53158, 16'd13245, 16'd10716, 16'd65230, 16'd5643, 16'd8654, 16'd34651, 16'd54961, 16'd58980});
	test_expansion(128'hf215b985e60a21ae810b80fd51587fbb, {16'd1686, 16'd12398, 16'd10052, 16'd51193, 16'd31665, 16'd33864, 16'd39329, 16'd35404, 16'd41035, 16'd58116, 16'd52133, 16'd18181, 16'd44047, 16'd28136, 16'd52768, 16'd3132, 16'd3430, 16'd22819, 16'd56505, 16'd13092, 16'd38959, 16'd49500, 16'd38869, 16'd218, 16'd23748, 16'd55852});
	test_expansion(128'hcb66de78a5e3238230f13659eff938e9, {16'd42717, 16'd37752, 16'd1480, 16'd41036, 16'd19269, 16'd19247, 16'd36014, 16'd34508, 16'd2284, 16'd9659, 16'd24096, 16'd6033, 16'd30507, 16'd50230, 16'd51687, 16'd41762, 16'd42960, 16'd61925, 16'd56576, 16'd46283, 16'd12551, 16'd637, 16'd48394, 16'd61355, 16'd3995, 16'd29374});
	test_expansion(128'h5018271e9b94a5e883f73b20743319fd, {16'd16553, 16'd3789, 16'd15395, 16'd39188, 16'd25650, 16'd21400, 16'd12200, 16'd52200, 16'd1781, 16'd14171, 16'd8190, 16'd17611, 16'd4847, 16'd40662, 16'd61739, 16'd12243, 16'd23022, 16'd32330, 16'd37542, 16'd6902, 16'd10494, 16'd40897, 16'd26656, 16'd35720, 16'd50518, 16'd50054});
	test_expansion(128'he2fff8961564423fd6a4c286ed524970, {16'd3212, 16'd54957, 16'd33707, 16'd50317, 16'd53991, 16'd63732, 16'd16858, 16'd42614, 16'd9275, 16'd64035, 16'd52597, 16'd2217, 16'd23257, 16'd32657, 16'd30161, 16'd24184, 16'd26051, 16'd47697, 16'd24573, 16'd11535, 16'd25117, 16'd45092, 16'd12476, 16'd2286, 16'd17808, 16'd4014});
	test_expansion(128'h0e08fe7744fe4a66c997d0e2b7bea6ec, {16'd32059, 16'd8946, 16'd28557, 16'd18322, 16'd48019, 16'd50703, 16'd54953, 16'd12382, 16'd46064, 16'd61945, 16'd11075, 16'd29617, 16'd30745, 16'd7901, 16'd24263, 16'd18963, 16'd46478, 16'd23434, 16'd27518, 16'd40176, 16'd55843, 16'd4855, 16'd53322, 16'd47787, 16'd60418, 16'd1211});
	test_expansion(128'h86aff9b62400e288ddbdadbb0009e194, {16'd36515, 16'd54688, 16'd10155, 16'd22538, 16'd44259, 16'd54479, 16'd15068, 16'd39051, 16'd43434, 16'd56921, 16'd23158, 16'd1119, 16'd27907, 16'd22465, 16'd37891, 16'd21152, 16'd40532, 16'd41117, 16'd64242, 16'd16490, 16'd15418, 16'd29110, 16'd23868, 16'd18325, 16'd27985, 16'd18715});
	test_expansion(128'h0ea9a89ecf46242431f47530635b4dd0, {16'd5580, 16'd50565, 16'd12886, 16'd22658, 16'd43326, 16'd13308, 16'd17439, 16'd2936, 16'd41896, 16'd7613, 16'd21916, 16'd28094, 16'd20498, 16'd15664, 16'd65137, 16'd39536, 16'd61698, 16'd49492, 16'd45634, 16'd22551, 16'd53556, 16'd29701, 16'd61183, 16'd36643, 16'd2347, 16'd35574});
	test_expansion(128'h25baf9f2174b26e25e411c58f6eea292, {16'd51197, 16'd12936, 16'd27380, 16'd14693, 16'd58512, 16'd240, 16'd24084, 16'd56545, 16'd46086, 16'd12878, 16'd26113, 16'd16983, 16'd43021, 16'd966, 16'd18358, 16'd22380, 16'd52354, 16'd26409, 16'd11748, 16'd46781, 16'd43113, 16'd49175, 16'd58115, 16'd56492, 16'd33493, 16'd7243});
	test_expansion(128'h689bc467d6f2bc010d52e971430c9f33, {16'd9596, 16'd17611, 16'd62852, 16'd6276, 16'd12735, 16'd19459, 16'd22673, 16'd49519, 16'd53444, 16'd61666, 16'd11456, 16'd28442, 16'd22676, 16'd583, 16'd60243, 16'd4499, 16'd55521, 16'd46618, 16'd42608, 16'd20392, 16'd15431, 16'd16476, 16'd59237, 16'd26155, 16'd4763, 16'd12103});
	test_expansion(128'he847aff02400fe95a799824a6d102fad, {16'd56343, 16'd7879, 16'd26935, 16'd59323, 16'd34980, 16'd29741, 16'd32288, 16'd38915, 16'd33315, 16'd44685, 16'd3646, 16'd17130, 16'd53825, 16'd39609, 16'd20091, 16'd45206, 16'd17989, 16'd26609, 16'd50154, 16'd23725, 16'd52791, 16'd35678, 16'd43461, 16'd24951, 16'd2069, 16'd50574});
	test_expansion(128'hcbe587b1388ea804a1f2b49da4a4a51c, {16'd60889, 16'd61191, 16'd36988, 16'd19711, 16'd7632, 16'd13194, 16'd21000, 16'd61167, 16'd6913, 16'd44308, 16'd16100, 16'd14771, 16'd62570, 16'd29269, 16'd49317, 16'd31623, 16'd53773, 16'd54101, 16'd16026, 16'd15278, 16'd51303, 16'd35241, 16'd53885, 16'd13393, 16'd49208, 16'd1083});
	test_expansion(128'h822c30034f4e0ab078c4723e73f5ed21, {16'd62814, 16'd52927, 16'd15914, 16'd61790, 16'd44364, 16'd31953, 16'd17010, 16'd8095, 16'd45123, 16'd44478, 16'd34649, 16'd44636, 16'd59644, 16'd37349, 16'd35427, 16'd18588, 16'd59455, 16'd36979, 16'd15761, 16'd42679, 16'd2510, 16'd17154, 16'd51715, 16'd21336, 16'd37375, 16'd47020});
	test_expansion(128'h5ae15340f667b97d28d468dc748ca4a5, {16'd38956, 16'd57670, 16'd17959, 16'd2400, 16'd29786, 16'd60471, 16'd6268, 16'd15469, 16'd40739, 16'd16834, 16'd36158, 16'd58434, 16'd50786, 16'd62571, 16'd35477, 16'd54893, 16'd7691, 16'd49072, 16'd53331, 16'd24700, 16'd43741, 16'd17442, 16'd22950, 16'd27983, 16'd12555, 16'd47930});
	test_expansion(128'h36d2545c5883890f7a1e147a7517a1f7, {16'd28600, 16'd32271, 16'd29457, 16'd3783, 16'd34538, 16'd8066, 16'd29095, 16'd949, 16'd63843, 16'd43539, 16'd30573, 16'd9326, 16'd35018, 16'd43311, 16'd19905, 16'd60362, 16'd64886, 16'd43676, 16'd54664, 16'd57658, 16'd21025, 16'd8372, 16'd46821, 16'd63204, 16'd50389, 16'd29504});
	test_expansion(128'h6598f05d53413ad64e7295481f19bacd, {16'd25967, 16'd25536, 16'd15402, 16'd5849, 16'd960, 16'd56180, 16'd41374, 16'd43398, 16'd59843, 16'd62784, 16'd45823, 16'd44677, 16'd40750, 16'd16339, 16'd35528, 16'd47763, 16'd29862, 16'd25123, 16'd16537, 16'd13442, 16'd34199, 16'd43702, 16'd7420, 16'd24092, 16'd62334, 16'd17016});
	test_expansion(128'hb70d250a88669c69334be02c97fd2a0a, {16'd64263, 16'd46136, 16'd35609, 16'd61241, 16'd11606, 16'd34155, 16'd412, 16'd14770, 16'd30482, 16'd12511, 16'd18040, 16'd52450, 16'd21663, 16'd58668, 16'd33076, 16'd6434, 16'd31567, 16'd65098, 16'd3296, 16'd24876, 16'd61860, 16'd8619, 16'd44102, 16'd7076, 16'd15198, 16'd33430});
	test_expansion(128'he0d61f3cdba100abeecec51b5d6a0ce6, {16'd42958, 16'd22087, 16'd62555, 16'd64205, 16'd34798, 16'd62085, 16'd37444, 16'd52919, 16'd47920, 16'd17725, 16'd19378, 16'd10963, 16'd9688, 16'd26119, 16'd1628, 16'd13054, 16'd42218, 16'd17669, 16'd8947, 16'd14359, 16'd25689, 16'd55908, 16'd2286, 16'd16798, 16'd10564, 16'd7352});
	test_expansion(128'ha05c3a9be4081fca4171925e315b29d8, {16'd14945, 16'd58990, 16'd24219, 16'd22332, 16'd36203, 16'd64635, 16'd19600, 16'd40516, 16'd26306, 16'd60385, 16'd38535, 16'd7428, 16'd15835, 16'd53278, 16'd13628, 16'd48199, 16'd15942, 16'd42873, 16'd24664, 16'd31687, 16'd25350, 16'd29722, 16'd59382, 16'd11502, 16'd40191, 16'd55377});
	test_expansion(128'hd8cfe3fbb71679d7736a0622255a10a2, {16'd62576, 16'd50870, 16'd14533, 16'd53067, 16'd38010, 16'd53075, 16'd56513, 16'd39381, 16'd61230, 16'd22276, 16'd46096, 16'd7637, 16'd63389, 16'd59683, 16'd13276, 16'd37169, 16'd43129, 16'd49201, 16'd31843, 16'd53600, 16'd3961, 16'd2569, 16'd47773, 16'd50962, 16'd62039, 16'd9155});
	test_expansion(128'h653bdd4f42d1c32dbf478b3868c5cfef, {16'd31537, 16'd65002, 16'd40133, 16'd35549, 16'd62551, 16'd17530, 16'd10401, 16'd43433, 16'd21668, 16'd60987, 16'd23163, 16'd62977, 16'd48235, 16'd20830, 16'd6053, 16'd16856, 16'd48090, 16'd27826, 16'd50384, 16'd43379, 16'd12803, 16'd47787, 16'd47926, 16'd51157, 16'd52762, 16'd6426});
	test_expansion(128'h4c274f89ba4f0630b08a8486aafef6c2, {16'd60343, 16'd12453, 16'd24436, 16'd5522, 16'd34626, 16'd60207, 16'd45903, 16'd779, 16'd24010, 16'd52610, 16'd31332, 16'd9256, 16'd39449, 16'd44938, 16'd9339, 16'd27549, 16'd20617, 16'd127, 16'd48929, 16'd4130, 16'd35867, 16'd27601, 16'd27068, 16'd52189, 16'd20872, 16'd2389});
	test_expansion(128'hbd2346cbfd3599f2a29935d64591a7cc, {16'd60778, 16'd4501, 16'd16181, 16'd33813, 16'd30407, 16'd55946, 16'd42185, 16'd17694, 16'd65491, 16'd11872, 16'd29450, 16'd7765, 16'd49589, 16'd15256, 16'd3404, 16'd33959, 16'd53282, 16'd15587, 16'd35509, 16'd37989, 16'd65094, 16'd13322, 16'd8436, 16'd35806, 16'd21714, 16'd64265});
	test_expansion(128'h70099ab5d0a0f3aec0d17ba650f2384a, {16'd6909, 16'd40003, 16'd62290, 16'd2345, 16'd27835, 16'd21111, 16'd38757, 16'd52561, 16'd11159, 16'd49693, 16'd27294, 16'd45549, 16'd61841, 16'd52228, 16'd54070, 16'd46844, 16'd19815, 16'd39973, 16'd41163, 16'd61465, 16'd16420, 16'd24076, 16'd955, 16'd4223, 16'd15452, 16'd11721});
	test_expansion(128'h17a9c67f744cc554c7e245e3637b2dd1, {16'd16192, 16'd39248, 16'd21017, 16'd3570, 16'd46696, 16'd30837, 16'd45085, 16'd1476, 16'd28419, 16'd26109, 16'd31956, 16'd46658, 16'd18247, 16'd936, 16'd51442, 16'd43210, 16'd38030, 16'd50324, 16'd57588, 16'd56177, 16'd55627, 16'd17476, 16'd25671, 16'd3262, 16'd39613, 16'd57002});
	test_expansion(128'h017cb329a63fe9ed447bb8f8a451b926, {16'd4213, 16'd6645, 16'd42429, 16'd25137, 16'd19852, 16'd15455, 16'd43664, 16'd8301, 16'd11989, 16'd24467, 16'd33352, 16'd1407, 16'd31102, 16'd51522, 16'd22060, 16'd39910, 16'd21158, 16'd14105, 16'd26278, 16'd28923, 16'd10579, 16'd25038, 16'd40748, 16'd13012, 16'd10248, 16'd26696});
	test_expansion(128'hb960097903f10b392a1a44b5af20753f, {16'd55268, 16'd60162, 16'd19659, 16'd43201, 16'd3312, 16'd15807, 16'd3324, 16'd65460, 16'd48643, 16'd9527, 16'd17937, 16'd26736, 16'd8301, 16'd50251, 16'd63063, 16'd52407, 16'd30542, 16'd31507, 16'd32636, 16'd28431, 16'd42080, 16'd48904, 16'd23221, 16'd56019, 16'd14618, 16'd46122});
	test_expansion(128'h4766dc16f5e24b9b4b21c60470e4a739, {16'd21821, 16'd2297, 16'd17335, 16'd42218, 16'd45185, 16'd4436, 16'd26111, 16'd10558, 16'd16279, 16'd59723, 16'd42516, 16'd57321, 16'd59691, 16'd17796, 16'd15831, 16'd27997, 16'd5530, 16'd40380, 16'd8604, 16'd43974, 16'd52302, 16'd63421, 16'd36343, 16'd26019, 16'd176, 16'd15110});
	test_expansion(128'ha17980e45e6881b689981e2b24bc07f2, {16'd30364, 16'd38482, 16'd58821, 16'd49243, 16'd16741, 16'd30741, 16'd30773, 16'd19918, 16'd63494, 16'd37648, 16'd23516, 16'd7153, 16'd59577, 16'd29611, 16'd3009, 16'd28207, 16'd33390, 16'd1600, 16'd32763, 16'd56724, 16'd47343, 16'd47091, 16'd33406, 16'd27006, 16'd52753, 16'd18421});
	test_expansion(128'hb3b31358fcbac464fb06389ffbc97a53, {16'd52532, 16'd43763, 16'd5333, 16'd62152, 16'd27830, 16'd47818, 16'd65114, 16'd54811, 16'd25387, 16'd8551, 16'd36715, 16'd55617, 16'd40709, 16'd47665, 16'd55258, 16'd40260, 16'd21061, 16'd21678, 16'd62582, 16'd13811, 16'd38854, 16'd53022, 16'd48431, 16'd40160, 16'd23924, 16'd20307});
	test_expansion(128'h3421cd090b52422c869993e14e93465d, {16'd29790, 16'd44151, 16'd40439, 16'd25607, 16'd18595, 16'd16151, 16'd26481, 16'd35808, 16'd14504, 16'd47624, 16'd16550, 16'd19630, 16'd46897, 16'd2684, 16'd20220, 16'd1753, 16'd20126, 16'd7575, 16'd12569, 16'd15476, 16'd48134, 16'd47094, 16'd28013, 16'd35283, 16'd8215, 16'd41817});
	test_expansion(128'h3df8f0b11d89b34b4ed5256b3e62ec5d, {16'd53509, 16'd5654, 16'd11625, 16'd9841, 16'd6198, 16'd38665, 16'd62769, 16'd20498, 16'd22800, 16'd55157, 16'd2394, 16'd34285, 16'd5674, 16'd62001, 16'd59768, 16'd34375, 16'd3718, 16'd29013, 16'd21811, 16'd32865, 16'd38510, 16'd509, 16'd39411, 16'd58451, 16'd6726, 16'd28969});
	test_expansion(128'hcee77a1cc9a1c239f87b18854cbe1f1e, {16'd59234, 16'd16263, 16'd57604, 16'd32559, 16'd1077, 16'd64987, 16'd7475, 16'd5521, 16'd21075, 16'd58071, 16'd38487, 16'd10635, 16'd45517, 16'd62497, 16'd45368, 16'd53142, 16'd41521, 16'd1998, 16'd60416, 16'd9228, 16'd5832, 16'd10430, 16'd22244, 16'd33583, 16'd53097, 16'd12384});
	test_expansion(128'h9e09368a48ba4536201192811b208dfd, {16'd37759, 16'd38519, 16'd5653, 16'd29116, 16'd54078, 16'd40863, 16'd4018, 16'd57200, 16'd28489, 16'd52176, 16'd22134, 16'd7328, 16'd19894, 16'd11928, 16'd22674, 16'd3459, 16'd48079, 16'd59000, 16'd18186, 16'd56853, 16'd20765, 16'd44687, 16'd53190, 16'd54699, 16'd51703, 16'd16296});
	test_expansion(128'h2e8a1b0c14103d3be55a0c1297dce3e9, {16'd35104, 16'd31925, 16'd12239, 16'd23477, 16'd47644, 16'd36247, 16'd54203, 16'd33055, 16'd46792, 16'd4932, 16'd33716, 16'd25549, 16'd43120, 16'd49194, 16'd55875, 16'd43673, 16'd63217, 16'd32460, 16'd48360, 16'd34302, 16'd12764, 16'd23270, 16'd6235, 16'd33428, 16'd15207, 16'd18457});
	test_expansion(128'h2a13b88ece10a68b97391d8951eb096f, {16'd16468, 16'd29896, 16'd49326, 16'd20462, 16'd23674, 16'd2847, 16'd53056, 16'd22057, 16'd3419, 16'd62197, 16'd63262, 16'd55834, 16'd59613, 16'd56417, 16'd17051, 16'd17705, 16'd1063, 16'd27830, 16'd53413, 16'd1151, 16'd60358, 16'd35712, 16'd29216, 16'd60643, 16'd6646, 16'd1881});
	test_expansion(128'h0c385b64701fa0ee54807fede017ca52, {16'd19060, 16'd56191, 16'd35807, 16'd27222, 16'd2763, 16'd10655, 16'd16842, 16'd58385, 16'd43662, 16'd27190, 16'd31764, 16'd6835, 16'd11158, 16'd31612, 16'd54541, 16'd35484, 16'd46516, 16'd8401, 16'd22367, 16'd12864, 16'd63297, 16'd29741, 16'd58779, 16'd62510, 16'd50773, 16'd23486});
	test_expansion(128'h97362991d98214f5a6fe2569b19ae21d, {16'd43678, 16'd24298, 16'd54423, 16'd14194, 16'd20691, 16'd26030, 16'd20654, 16'd65136, 16'd54997, 16'd795, 16'd47351, 16'd52905, 16'd27256, 16'd45993, 16'd18110, 16'd51296, 16'd23184, 16'd63844, 16'd50970, 16'd21797, 16'd1604, 16'd43746, 16'd60430, 16'd30882, 16'd59660, 16'd17151});
	test_expansion(128'ha82dd40fcc827683084a588c99974247, {16'd33168, 16'd48454, 16'd18472, 16'd64053, 16'd62506, 16'd43894, 16'd33473, 16'd3001, 16'd41293, 16'd57703, 16'd61460, 16'd417, 16'd14848, 16'd40483, 16'd42338, 16'd47996, 16'd21134, 16'd28299, 16'd36777, 16'd58187, 16'd7719, 16'd38311, 16'd5235, 16'd41896, 16'd13515, 16'd42777});
	test_expansion(128'h703760ddf527c303c6ea5e9921b98287, {16'd16624, 16'd51885, 16'd41864, 16'd8452, 16'd12360, 16'd15219, 16'd6661, 16'd25773, 16'd60781, 16'd60315, 16'd64178, 16'd35062, 16'd42954, 16'd12384, 16'd48235, 16'd9463, 16'd29338, 16'd435, 16'd42477, 16'd13515, 16'd60772, 16'd1782, 16'd20223, 16'd24920, 16'd64549, 16'd13430});
	test_expansion(128'hf43ec8c4530ba83e9aa233e3421c8159, {16'd51654, 16'd49156, 16'd21936, 16'd3919, 16'd22282, 16'd59084, 16'd33833, 16'd2101, 16'd59013, 16'd64443, 16'd53179, 16'd24884, 16'd37053, 16'd47926, 16'd36985, 16'd64853, 16'd49896, 16'd56204, 16'd46390, 16'd23440, 16'd19473, 16'd19717, 16'd5853, 16'd53889, 16'd40812, 16'd50276});
	test_expansion(128'hcde381f2372dd85359fc2ec3080ab9ac, {16'd10791, 16'd6460, 16'd38344, 16'd37803, 16'd46060, 16'd8093, 16'd29086, 16'd64122, 16'd24503, 16'd62591, 16'd47300, 16'd25168, 16'd3551, 16'd63841, 16'd46630, 16'd54990, 16'd22034, 16'd9543, 16'd22602, 16'd35898, 16'd8842, 16'd30322, 16'd13552, 16'd60471, 16'd50907, 16'd38930});
	test_expansion(128'h9369b780f144d11175861a9b57d3737c, {16'd7739, 16'd29124, 16'd54180, 16'd45889, 16'd43209, 16'd64626, 16'd63862, 16'd15352, 16'd9628, 16'd28171, 16'd59256, 16'd22097, 16'd619, 16'd32966, 16'd19456, 16'd61678, 16'd36049, 16'd34862, 16'd24698, 16'd53864, 16'd32741, 16'd9747, 16'd21099, 16'd33218, 16'd62269, 16'd13281});
	test_expansion(128'hf51e1853ae35d53b99911f7b06d1afbc, {16'd34939, 16'd9057, 16'd56444, 16'd58120, 16'd16676, 16'd3382, 16'd23886, 16'd52346, 16'd64736, 16'd61998, 16'd10746, 16'd9513, 16'd36331, 16'd33190, 16'd49909, 16'd48937, 16'd47382, 16'd55008, 16'd45928, 16'd24917, 16'd18046, 16'd23904, 16'd13980, 16'd58843, 16'd11316, 16'd54296});
	test_expansion(128'h1766a237dd0681de1b2f91ff75f85cc5, {16'd15262, 16'd48948, 16'd8590, 16'd44252, 16'd15843, 16'd13515, 16'd60329, 16'd61377, 16'd26720, 16'd59680, 16'd46443, 16'd19705, 16'd64541, 16'd6883, 16'd17456, 16'd55852, 16'd15517, 16'd60144, 16'd52137, 16'd51449, 16'd16019, 16'd42339, 16'd34281, 16'd10025, 16'd5894, 16'd10732});
	test_expansion(128'haa4f8f9cbc6be5b3a42649e07895a9b8, {16'd30877, 16'd13224, 16'd40955, 16'd34516, 16'd13577, 16'd19091, 16'd58346, 16'd11447, 16'd45621, 16'd65, 16'd57851, 16'd29168, 16'd44294, 16'd12638, 16'd37971, 16'd31667, 16'd5545, 16'd5722, 16'd29052, 16'd3363, 16'd29958, 16'd46074, 16'd61896, 16'd21060, 16'd61480, 16'd21269});
	test_expansion(128'h3cc6948d22ce55c799ba8f93a744077d, {16'd45381, 16'd24203, 16'd1817, 16'd59308, 16'd12903, 16'd11337, 16'd60772, 16'd6284, 16'd56721, 16'd10262, 16'd42212, 16'd51932, 16'd38571, 16'd3629, 16'd38854, 16'd55620, 16'd21646, 16'd14538, 16'd41323, 16'd11930, 16'd16804, 16'd63147, 16'd21099, 16'd55924, 16'd37350, 16'd52529});
	test_expansion(128'haedd804f96c355f5256fbe2fa80db295, {16'd63962, 16'd3705, 16'd6284, 16'd59501, 16'd46276, 16'd23859, 16'd13212, 16'd59381, 16'd45490, 16'd56842, 16'd43191, 16'd64507, 16'd11618, 16'd56697, 16'd39823, 16'd31436, 16'd54542, 16'd596, 16'd7191, 16'd2257, 16'd4708, 16'd63651, 16'd55520, 16'd33283, 16'd50401, 16'd10637});
	test_expansion(128'h3a5db1e2a47783ed26dac9a2e68dd87c, {16'd5843, 16'd47095, 16'd13307, 16'd10312, 16'd41187, 16'd32074, 16'd58129, 16'd22808, 16'd12949, 16'd48895, 16'd47889, 16'd57479, 16'd15364, 16'd7846, 16'd45103, 16'd3449, 16'd31847, 16'd60859, 16'd32852, 16'd3844, 16'd15109, 16'd27954, 16'd41518, 16'd256, 16'd63698, 16'd37781});
	test_expansion(128'h99ab955666fb52fa684b9cdeb8f86239, {16'd42054, 16'd61706, 16'd61997, 16'd7445, 16'd10164, 16'd28433, 16'd11389, 16'd59780, 16'd41791, 16'd37019, 16'd17629, 16'd22399, 16'd40258, 16'd14247, 16'd64176, 16'd22982, 16'd37930, 16'd35680, 16'd55984, 16'd17578, 16'd3943, 16'd29885, 16'd58729, 16'd42169, 16'd12011, 16'd31313});
	test_expansion(128'hc55a92c70649e6f102e013d1f4d61f22, {16'd8380, 16'd15918, 16'd51211, 16'd37312, 16'd65471, 16'd25578, 16'd10405, 16'd56706, 16'd65084, 16'd42760, 16'd12098, 16'd18689, 16'd15768, 16'd24734, 16'd19395, 16'd39355, 16'd17885, 16'd60414, 16'd33149, 16'd3952, 16'd24880, 16'd59218, 16'd59705, 16'd4443, 16'd63133, 16'd48696});
	test_expansion(128'h53142d11d009ca4556c3cac597dba485, {16'd10998, 16'd61033, 16'd16068, 16'd51174, 16'd55902, 16'd20249, 16'd60391, 16'd46008, 16'd53585, 16'd6953, 16'd20327, 16'd16700, 16'd58316, 16'd3515, 16'd1912, 16'd55018, 16'd28514, 16'd56392, 16'd24588, 16'd28535, 16'd6821, 16'd13046, 16'd6028, 16'd22335, 16'd30979, 16'd62407});
	test_expansion(128'hfce11a7413cd7b393ccbfd551a6a4557, {16'd35831, 16'd40828, 16'd14406, 16'd35858, 16'd33587, 16'd7374, 16'd41757, 16'd1343, 16'd38841, 16'd65083, 16'd53926, 16'd1793, 16'd58834, 16'd14024, 16'd8448, 16'd14061, 16'd3516, 16'd16315, 16'd30507, 16'd43533, 16'd9604, 16'd59109, 16'd62949, 16'd37054, 16'd13581, 16'd9848});
	test_expansion(128'h6ce702e2679d406cb533af28b229201c, {16'd46500, 16'd33218, 16'd15125, 16'd60717, 16'd11060, 16'd52026, 16'd19230, 16'd8691, 16'd51873, 16'd44337, 16'd20396, 16'd51428, 16'd59351, 16'd4877, 16'd54142, 16'd60728, 16'd61146, 16'd48426, 16'd45325, 16'd1542, 16'd4308, 16'd15624, 16'd51118, 16'd31231, 16'd41253, 16'd5518});
	test_expansion(128'h53697048ee3dcfa706694f53eccafdb1, {16'd55413, 16'd21139, 16'd9317, 16'd60978, 16'd31004, 16'd17525, 16'd24523, 16'd39806, 16'd396, 16'd1314, 16'd8889, 16'd12088, 16'd35913, 16'd22608, 16'd10365, 16'd59995, 16'd51599, 16'd35248, 16'd8124, 16'd63957, 16'd24904, 16'd41906, 16'd51357, 16'd22251, 16'd65383, 16'd27710});
	test_expansion(128'h61fc3394602416c8a1cc6a1b57abaaf4, {16'd6791, 16'd39468, 16'd24410, 16'd19612, 16'd33347, 16'd10373, 16'd5290, 16'd4767, 16'd40179, 16'd40682, 16'd64, 16'd806, 16'd58042, 16'd33944, 16'd21328, 16'd2541, 16'd11672, 16'd15194, 16'd31938, 16'd10000, 16'd20769, 16'd31848, 16'd62447, 16'd8506, 16'd63042, 16'd49592});
	test_expansion(128'h17314cfb71ea1008b3bbbb7c7536b5f6, {16'd60028, 16'd39542, 16'd63679, 16'd19357, 16'd65039, 16'd13136, 16'd34367, 16'd14205, 16'd52425, 16'd24279, 16'd33059, 16'd4093, 16'd16387, 16'd38429, 16'd27518, 16'd18876, 16'd331, 16'd49840, 16'd16259, 16'd32642, 16'd34600, 16'd48765, 16'd31593, 16'd22962, 16'd63066, 16'd6464});
	test_expansion(128'h993d9c8660ff4d2d22fbbaf2504d4030, {16'd9697, 16'd43088, 16'd48374, 16'd62538, 16'd57148, 16'd1172, 16'd64810, 16'd10474, 16'd27948, 16'd1349, 16'd6476, 16'd27626, 16'd5080, 16'd53593, 16'd56918, 16'd24980, 16'd40202, 16'd17118, 16'd40212, 16'd47021, 16'd31143, 16'd2653, 16'd905, 16'd2395, 16'd16453, 16'd61251});
	test_expansion(128'h086c1f7bfeb91f1f188ea2d165db2720, {16'd3957, 16'd27505, 16'd15416, 16'd4257, 16'd37119, 16'd45580, 16'd62831, 16'd51858, 16'd43806, 16'd20770, 16'd37719, 16'd51146, 16'd28723, 16'd49316, 16'd52085, 16'd50663, 16'd13454, 16'd25769, 16'd26266, 16'd63406, 16'd4586, 16'd64726, 16'd9191, 16'd21200, 16'd62706, 16'd13822});
	test_expansion(128'h5d6aaa8e9ccc12f7264cf44d69ad1cd8, {16'd63478, 16'd13767, 16'd7290, 16'd16489, 16'd7265, 16'd41602, 16'd53406, 16'd17527, 16'd36534, 16'd19759, 16'd57631, 16'd13405, 16'd13917, 16'd61674, 16'd27570, 16'd62491, 16'd11575, 16'd80, 16'd35995, 16'd5444, 16'd50715, 16'd8893, 16'd6701, 16'd1865, 16'd57150, 16'd18007});
	test_expansion(128'ha59384b18fc1a2519f33951d3e57468b, {16'd60423, 16'd45628, 16'd36831, 16'd12073, 16'd19069, 16'd61874, 16'd14433, 16'd34100, 16'd64411, 16'd25985, 16'd18542, 16'd48961, 16'd51128, 16'd52330, 16'd11548, 16'd19429, 16'd62577, 16'd39373, 16'd7057, 16'd10620, 16'd53180, 16'd46318, 16'd38416, 16'd63390, 16'd17297, 16'd38834});
	test_expansion(128'h5595d20603f076e8826c40304ccdf0a5, {16'd57575, 16'd4201, 16'd61075, 16'd21932, 16'd4275, 16'd55616, 16'd47798, 16'd14750, 16'd62654, 16'd29235, 16'd58864, 16'd13974, 16'd34975, 16'd52021, 16'd5659, 16'd19994, 16'd51404, 16'd52186, 16'd24979, 16'd27067, 16'd21892, 16'd24890, 16'd40920, 16'd60208, 16'd26558, 16'd64170});
	test_expansion(128'h5b67f15f5d671c7641421d879c509d3e, {16'd31883, 16'd30115, 16'd1852, 16'd61944, 16'd45606, 16'd37402, 16'd56044, 16'd33121, 16'd59551, 16'd37952, 16'd58532, 16'd1678, 16'd10697, 16'd46780, 16'd19336, 16'd22169, 16'd27216, 16'd56875, 16'd389, 16'd21869, 16'd63029, 16'd31173, 16'd30603, 16'd1088, 16'd36925, 16'd57017});
	test_expansion(128'h54bd83b34e01b4205b6b5915f1424f97, {16'd15281, 16'd4065, 16'd16809, 16'd20594, 16'd38048, 16'd20709, 16'd54911, 16'd64602, 16'd65414, 16'd5053, 16'd52218, 16'd30600, 16'd64208, 16'd38726, 16'd3032, 16'd57222, 16'd45601, 16'd55867, 16'd4167, 16'd50580, 16'd41608, 16'd27309, 16'd63437, 16'd50911, 16'd18517, 16'd13390});
	test_expansion(128'he8984c7fe0a770e81b12234907d90cca, {16'd28817, 16'd7289, 16'd4689, 16'd10380, 16'd1740, 16'd44469, 16'd44332, 16'd5057, 16'd55304, 16'd19811, 16'd7703, 16'd48195, 16'd54789, 16'd45618, 16'd24063, 16'd27221, 16'd28445, 16'd14837, 16'd10625, 16'd23732, 16'd49511, 16'd23736, 16'd42408, 16'd41305, 16'd54474, 16'd55207});
	test_expansion(128'he27ed4931eef91405d5d64d5d21c1d6c, {16'd25363, 16'd27670, 16'd64453, 16'd10772, 16'd34891, 16'd29452, 16'd43659, 16'd15329, 16'd44684, 16'd462, 16'd48515, 16'd52094, 16'd60782, 16'd40500, 16'd64076, 16'd59046, 16'd5375, 16'd19356, 16'd20977, 16'd3363, 16'd57678, 16'd52170, 16'd11463, 16'd29201, 16'd193, 16'd62900});
	test_expansion(128'hc4a7ee4408a1291e9311745fc3f7041e, {16'd38383, 16'd54136, 16'd30855, 16'd24846, 16'd21118, 16'd9346, 16'd24563, 16'd16069, 16'd9706, 16'd4003, 16'd41987, 16'd8712, 16'd16084, 16'd20174, 16'd35322, 16'd14917, 16'd61952, 16'd45385, 16'd22002, 16'd39206, 16'd52430, 16'd17791, 16'd20488, 16'd63551, 16'd11366, 16'd5662});
	test_expansion(128'h3d15c240c9ea678e6d8dcb03cdda1da5, {16'd29401, 16'd59042, 16'd20937, 16'd273, 16'd21127, 16'd46483, 16'd64922, 16'd54561, 16'd54219, 16'd41827, 16'd6165, 16'd9443, 16'd63771, 16'd53026, 16'd10947, 16'd43320, 16'd37204, 16'd53364, 16'd40108, 16'd44590, 16'd37745, 16'd41481, 16'd42626, 16'd21042, 16'd2302, 16'd47486});
	test_expansion(128'h0e85d2592f08cc31b104f60d4c8f34a5, {16'd37016, 16'd49980, 16'd13005, 16'd37082, 16'd65251, 16'd37115, 16'd19732, 16'd27659, 16'd25222, 16'd1189, 16'd40617, 16'd31124, 16'd2476, 16'd24486, 16'd53096, 16'd13295, 16'd38373, 16'd3822, 16'd7619, 16'd34553, 16'd35187, 16'd7196, 16'd61233, 16'd4001, 16'd8129, 16'd16336});
	test_expansion(128'h98a4071ef6fdb94a78433ed455e5bf9c, {16'd51724, 16'd41457, 16'd8342, 16'd53147, 16'd25460, 16'd5650, 16'd20065, 16'd17195, 16'd29943, 16'd4665, 16'd16760, 16'd14876, 16'd20323, 16'd17500, 16'd33490, 16'd45132, 16'd47886, 16'd46150, 16'd61435, 16'd45247, 16'd9272, 16'd13691, 16'd6420, 16'd44867, 16'd44639, 16'd35506});
	test_expansion(128'hb16806d325cf1efd93c583dcfed18eae, {16'd10915, 16'd22808, 16'd22114, 16'd60430, 16'd10004, 16'd57708, 16'd19719, 16'd18182, 16'd27699, 16'd18117, 16'd64474, 16'd43463, 16'd15859, 16'd43849, 16'd6819, 16'd49445, 16'd39567, 16'd14151, 16'd17617, 16'd3931, 16'd38306, 16'd55008, 16'd31770, 16'd5081, 16'd57363, 16'd56417});
	test_expansion(128'h9b3cc334fc5f2a97421be36f47a0498c, {16'd23369, 16'd27235, 16'd18082, 16'd44676, 16'd11000, 16'd27045, 16'd2060, 16'd33105, 16'd13335, 16'd36641, 16'd30894, 16'd28462, 16'd7300, 16'd23996, 16'd27784, 16'd6787, 16'd32321, 16'd53877, 16'd49211, 16'd23111, 16'd57871, 16'd31816, 16'd57788, 16'd63225, 16'd23586, 16'd44404});
	test_expansion(128'hf97de8fed4a9a00658c60066d94993d8, {16'd45932, 16'd29635, 16'd105, 16'd18223, 16'd36722, 16'd56058, 16'd35172, 16'd62822, 16'd5875, 16'd15982, 16'd11213, 16'd13036, 16'd32794, 16'd31862, 16'd40083, 16'd62879, 16'd54248, 16'd53092, 16'd12899, 16'd62020, 16'd62450, 16'd1889, 16'd33316, 16'd16618, 16'd18932, 16'd7933});
	test_expansion(128'hc039e227172617fde28d3e25fbab3c64, {16'd42534, 16'd18288, 16'd12391, 16'd5884, 16'd9322, 16'd45188, 16'd10708, 16'd31647, 16'd54722, 16'd19500, 16'd36139, 16'd12787, 16'd9664, 16'd20071, 16'd52680, 16'd13185, 16'd5543, 16'd7894, 16'd12139, 16'd58221, 16'd65427, 16'd40407, 16'd30031, 16'd63114, 16'd19119, 16'd24206});
	test_expansion(128'he910113469ddc7e62c0284202245fecd, {16'd45965, 16'd11214, 16'd25967, 16'd59011, 16'd10097, 16'd28397, 16'd30599, 16'd18544, 16'd39884, 16'd15522, 16'd26270, 16'd23976, 16'd26530, 16'd27479, 16'd65281, 16'd18092, 16'd44234, 16'd22566, 16'd47641, 16'd5160, 16'd31721, 16'd18014, 16'd45393, 16'd58203, 16'd26560, 16'd35162});
	test_expansion(128'h14804ed877dba04d39c0baee1abb0f31, {16'd63784, 16'd43963, 16'd38818, 16'd39790, 16'd59432, 16'd47607, 16'd13541, 16'd65522, 16'd30777, 16'd47715, 16'd8804, 16'd52508, 16'd36676, 16'd31415, 16'd35804, 16'd44977, 16'd28054, 16'd31585, 16'd7476, 16'd51033, 16'd51945, 16'd35947, 16'd22381, 16'd5549, 16'd15500, 16'd9628});
	test_expansion(128'h5317e771851b94bfc9827114bcac7449, {16'd35287, 16'd7933, 16'd37365, 16'd53227, 16'd60911, 16'd29869, 16'd7736, 16'd64183, 16'd42294, 16'd12953, 16'd27588, 16'd49808, 16'd30709, 16'd49848, 16'd59677, 16'd8868, 16'd55298, 16'd55426, 16'd56513, 16'd39975, 16'd13665, 16'd43182, 16'd42997, 16'd56952, 16'd63588, 16'd60660});
	test_expansion(128'ha07f694104aff241e3c0b637d46340e0, {16'd56767, 16'd55073, 16'd17853, 16'd36377, 16'd53790, 16'd52441, 16'd11888, 16'd26948, 16'd61581, 16'd49632, 16'd62190, 16'd1162, 16'd63482, 16'd8379, 16'd58143, 16'd54045, 16'd5198, 16'd25632, 16'd56664, 16'd64677, 16'd2643, 16'd48444, 16'd12592, 16'd53138, 16'd22355, 16'd6327});
	test_expansion(128'h512c03b87bcc1d15820208b2486953ce, {16'd1513, 16'd1859, 16'd21736, 16'd15924, 16'd3456, 16'd42191, 16'd57148, 16'd11041, 16'd47575, 16'd27946, 16'd55549, 16'd44177, 16'd38656, 16'd27390, 16'd34948, 16'd44392, 16'd4532, 16'd50183, 16'd58162, 16'd51494, 16'd2647, 16'd45011, 16'd25089, 16'd13121, 16'd6828, 16'd14155});
	test_expansion(128'h1970c2e1cb2c94bdabf089178a7b5f47, {16'd11755, 16'd11057, 16'd10305, 16'd30381, 16'd52122, 16'd5714, 16'd58435, 16'd11015, 16'd49656, 16'd40891, 16'd35426, 16'd52799, 16'd23129, 16'd3375, 16'd57565, 16'd60036, 16'd33654, 16'd57120, 16'd59145, 16'd12556, 16'd37241, 16'd2263, 16'd44339, 16'd57568, 16'd33777, 16'd17191});
	test_expansion(128'h8d66e43e7e5b0708f521ec64bb6bd103, {16'd63870, 16'd60254, 16'd17966, 16'd39910, 16'd20325, 16'd36698, 16'd6256, 16'd44830, 16'd62570, 16'd9962, 16'd19467, 16'd52996, 16'd60640, 16'd45081, 16'd21936, 16'd47010, 16'd41310, 16'd44214, 16'd47056, 16'd35024, 16'd6388, 16'd47470, 16'd56168, 16'd61254, 16'd42604, 16'd2759});
	test_expansion(128'h89927954f84c8c4a2d8931aeed5acbb9, {16'd41252, 16'd56217, 16'd46294, 16'd24210, 16'd50510, 16'd30474, 16'd65082, 16'd50878, 16'd25883, 16'd22989, 16'd8705, 16'd64197, 16'd5332, 16'd7473, 16'd55852, 16'd37552, 16'd34585, 16'd36640, 16'd51186, 16'd17640, 16'd36714, 16'd42213, 16'd49637, 16'd13251, 16'd40442, 16'd41647});
	test_expansion(128'h6477f1ff04bf77a310de3aa92f850688, {16'd51506, 16'd34028, 16'd36449, 16'd6517, 16'd9623, 16'd35216, 16'd30472, 16'd28585, 16'd21835, 16'd56524, 16'd36522, 16'd40572, 16'd31048, 16'd10907, 16'd35759, 16'd49828, 16'd23791, 16'd16380, 16'd40028, 16'd14888, 16'd44873, 16'd30426, 16'd28701, 16'd39924, 16'd6000, 16'd5789});
	test_expansion(128'h4a0706b0a931f596a51d1c0a9429c67e, {16'd3653, 16'd5170, 16'd12299, 16'd50398, 16'd4668, 16'd59059, 16'd34246, 16'd2378, 16'd55753, 16'd50598, 16'd19925, 16'd37372, 16'd49165, 16'd48240, 16'd39978, 16'd61965, 16'd21346, 16'd6706, 16'd52489, 16'd64008, 16'd24232, 16'd52595, 16'd10828, 16'd64704, 16'd41299, 16'd3650});
	test_expansion(128'hce9600897762acc34e31feb9ff722c45, {16'd63900, 16'd55322, 16'd64082, 16'd24115, 16'd12027, 16'd8567, 16'd55484, 16'd978, 16'd33299, 16'd60760, 16'd29316, 16'd58370, 16'd31443, 16'd3307, 16'd57095, 16'd17441, 16'd43616, 16'd26862, 16'd33535, 16'd63040, 16'd62050, 16'd48319, 16'd13492, 16'd52668, 16'd34763, 16'd47188});
	test_expansion(128'h4daa347d6405821b9d2e0258f639b19c, {16'd10865, 16'd58286, 16'd14923, 16'd56689, 16'd54454, 16'd44413, 16'd32371, 16'd248, 16'd63874, 16'd58512, 16'd3842, 16'd52357, 16'd33263, 16'd1007, 16'd13021, 16'd55958, 16'd63556, 16'd6847, 16'd43780, 16'd59833, 16'd32309, 16'd2448, 16'd38002, 16'd40427, 16'd47324, 16'd21294});
	test_expansion(128'h17d24e14fbf12fe96b4d225aed92bf3c, {16'd51560, 16'd28429, 16'd38408, 16'd4383, 16'd47943, 16'd24084, 16'd7496, 16'd4914, 16'd24275, 16'd21617, 16'd51204, 16'd6577, 16'd29187, 16'd43554, 16'd51525, 16'd38626, 16'd9953, 16'd31055, 16'd254, 16'd45343, 16'd326, 16'd30407, 16'd42261, 16'd52190, 16'd61467, 16'd30091});
	test_expansion(128'h9d5dffb048eb43d4ec33c3c6006a4a59, {16'd401, 16'd5029, 16'd59073, 16'd40573, 16'd8566, 16'd7505, 16'd3707, 16'd44442, 16'd22564, 16'd22126, 16'd23196, 16'd17223, 16'd8544, 16'd50207, 16'd23497, 16'd45915, 16'd44221, 16'd47375, 16'd28889, 16'd36254, 16'd20491, 16'd6600, 16'd20047, 16'd40422, 16'd34023, 16'd63118});
	test_expansion(128'h5cb0b9d4296cfb6e3049d450d90bf28e, {16'd21588, 16'd49151, 16'd37277, 16'd2061, 16'd40016, 16'd27188, 16'd7030, 16'd47220, 16'd7411, 16'd7998, 16'd21101, 16'd13200, 16'd65418, 16'd13074, 16'd16232, 16'd59724, 16'd49594, 16'd37843, 16'd37858, 16'd57954, 16'd49974, 16'd55373, 16'd15318, 16'd6005, 16'd47961, 16'd15596});
	test_expansion(128'h2d13cfd4ba6cb1f0b105399c13caa07e, {16'd43862, 16'd62479, 16'd2717, 16'd58390, 16'd31280, 16'd27492, 16'd58901, 16'd30831, 16'd48275, 16'd15256, 16'd37169, 16'd31582, 16'd56939, 16'd9445, 16'd27675, 16'd27762, 16'd40144, 16'd29959, 16'd54287, 16'd12169, 16'd5405, 16'd51495, 16'd54416, 16'd63455, 16'd44628, 16'd5054});
	test_expansion(128'h8dea537a42355999fc9fd76eafdcea95, {16'd15924, 16'd47534, 16'd8812, 16'd52972, 16'd21015, 16'd45811, 16'd54658, 16'd53295, 16'd5186, 16'd3116, 16'd33280, 16'd45667, 16'd13691, 16'd56379, 16'd61422, 16'd31606, 16'd30101, 16'd54382, 16'd31789, 16'd32718, 16'd33346, 16'd41200, 16'd27988, 16'd1904, 16'd17, 16'd41573});
	test_expansion(128'hab93b3e25de543e8019216c9aa224792, {16'd32814, 16'd18006, 16'd5890, 16'd42399, 16'd5220, 16'd26745, 16'd12157, 16'd10327, 16'd23377, 16'd4553, 16'd35363, 16'd49875, 16'd43654, 16'd27585, 16'd49810, 16'd43930, 16'd46933, 16'd19501, 16'd9665, 16'd24986, 16'd20630, 16'd65446, 16'd48338, 16'd40608, 16'd56085, 16'd28152});
	test_expansion(128'h5477d1be5bbd17fd7f4214cdb6cee88d, {16'd31247, 16'd39641, 16'd12479, 16'd53388, 16'd36294, 16'd55297, 16'd25255, 16'd24136, 16'd50090, 16'd13342, 16'd59886, 16'd13130, 16'd25369, 16'd1451, 16'd11275, 16'd18021, 16'd34585, 16'd50980, 16'd9481, 16'd51778, 16'd15245, 16'd35650, 16'd21906, 16'd41694, 16'd34526, 16'd18835});
	test_expansion(128'hf008e4eb63e33193a07ea39ac1d65279, {16'd61985, 16'd38387, 16'd41447, 16'd9932, 16'd4149, 16'd26185, 16'd31809, 16'd28340, 16'd5948, 16'd39991, 16'd62542, 16'd13651, 16'd39797, 16'd57594, 16'd52541, 16'd49374, 16'd56865, 16'd1433, 16'd28696, 16'd63093, 16'd50095, 16'd31407, 16'd17282, 16'd48948, 16'd794, 16'd65223});
	test_expansion(128'h5a887745034ec0abe2a0365d58b2dc39, {16'd1802, 16'd8741, 16'd27951, 16'd6319, 16'd31662, 16'd30176, 16'd62298, 16'd47909, 16'd5645, 16'd48405, 16'd62769, 16'd44659, 16'd24536, 16'd57736, 16'd13497, 16'd19324, 16'd23592, 16'd25474, 16'd34495, 16'd54523, 16'd43939, 16'd34553, 16'd19044, 16'd33869, 16'd16462, 16'd44565});
	test_expansion(128'h874d841b591d44a44c4964ad2c57ffad, {16'd19482, 16'd4056, 16'd40172, 16'd36554, 16'd53993, 16'd19204, 16'd53743, 16'd60919, 16'd59069, 16'd42076, 16'd12533, 16'd64951, 16'd18741, 16'd26933, 16'd54602, 16'd14165, 16'd53900, 16'd10952, 16'd43492, 16'd44547, 16'd35632, 16'd53523, 16'd65477, 16'd43605, 16'd63372, 16'd29883});
	test_expansion(128'h424b79052f43bc1c93d5c6609af5dbfc, {16'd65434, 16'd4095, 16'd12832, 16'd33289, 16'd56846, 16'd51215, 16'd47402, 16'd42545, 16'd26691, 16'd55747, 16'd58939, 16'd20224, 16'd17282, 16'd57418, 16'd22351, 16'd1193, 16'd12963, 16'd38913, 16'd19185, 16'd3291, 16'd17623, 16'd49415, 16'd5078, 16'd10664, 16'd33165, 16'd25268});
	test_expansion(128'h789870ced6979bff68b05fbc9e7fc72f, {16'd10186, 16'd10523, 16'd28048, 16'd36078, 16'd40002, 16'd9643, 16'd25910, 16'd21861, 16'd61427, 16'd59484, 16'd53972, 16'd42028, 16'd26251, 16'd25929, 16'd8717, 16'd59152, 16'd19596, 16'd35716, 16'd27132, 16'd10438, 16'd19849, 16'd40785, 16'd10740, 16'd11929, 16'd49923, 16'd1189});
	test_expansion(128'h0f8c05511b1f14f837f40ead8c2eeef9, {16'd10370, 16'd43920, 16'd17472, 16'd37629, 16'd61702, 16'd52642, 16'd28785, 16'd30426, 16'd7083, 16'd56483, 16'd22600, 16'd1175, 16'd63759, 16'd21246, 16'd64644, 16'd28359, 16'd48271, 16'd1664, 16'd38941, 16'd38193, 16'd9532, 16'd46732, 16'd41162, 16'd40401, 16'd17798, 16'd56886});
	test_expansion(128'h850ef6a1458219b3b4accf53b9933841, {16'd8861, 16'd14289, 16'd25238, 16'd32128, 16'd20857, 16'd15456, 16'd61106, 16'd35770, 16'd29427, 16'd28708, 16'd27926, 16'd6683, 16'd48916, 16'd24725, 16'd5578, 16'd38574, 16'd28649, 16'd38179, 16'd45412, 16'd62281, 16'd16484, 16'd10198, 16'd61776, 16'd22534, 16'd64753, 16'd35090});
	test_expansion(128'hfd027e66767f17029a738324c3cc0d06, {16'd36195, 16'd25707, 16'd6, 16'd34296, 16'd52967, 16'd38333, 16'd37828, 16'd12237, 16'd15890, 16'd64596, 16'd25384, 16'd12486, 16'd57931, 16'd5144, 16'd22078, 16'd6826, 16'd24029, 16'd19477, 16'd7442, 16'd1236, 16'd26742, 16'd52652, 16'd55424, 16'd24730, 16'd43680, 16'd45174});
	test_expansion(128'h0e20488d51959f633b186eb12a0e3db4, {16'd8383, 16'd18022, 16'd47729, 16'd20471, 16'd53951, 16'd22042, 16'd18981, 16'd17201, 16'd53830, 16'd47017, 16'd59105, 16'd54011, 16'd7641, 16'd50409, 16'd48278, 16'd21006, 16'd43389, 16'd16011, 16'd36871, 16'd59287, 16'd58357, 16'd12476, 16'd46748, 16'd20372, 16'd3834, 16'd25622});
	test_expansion(128'he07395efafd2e6e71f34a9ebd54b2e69, {16'd31463, 16'd28319, 16'd6405, 16'd59152, 16'd54635, 16'd6959, 16'd38915, 16'd43913, 16'd58352, 16'd47028, 16'd32209, 16'd50980, 16'd49591, 16'd25411, 16'd846, 16'd35004, 16'd44220, 16'd37223, 16'd52888, 16'd65185, 16'd31420, 16'd14347, 16'd34584, 16'd26005, 16'd6194, 16'd24037});
	test_expansion(128'hf833565a4f6a46c3b74b024136b7e543, {16'd24827, 16'd16275, 16'd47337, 16'd39900, 16'd51293, 16'd29112, 16'd25494, 16'd30183, 16'd33937, 16'd56757, 16'd60571, 16'd27392, 16'd62949, 16'd5920, 16'd9318, 16'd18977, 16'd44373, 16'd37402, 16'd30648, 16'd1312, 16'd10831, 16'd63447, 16'd54388, 16'd32350, 16'd20679, 16'd5004});
	test_expansion(128'h99f40ab41abfd06208ebe944017b2706, {16'd35683, 16'd23547, 16'd32903, 16'd16838, 16'd63452, 16'd53133, 16'd22529, 16'd56338, 16'd57077, 16'd2105, 16'd7051, 16'd46569, 16'd30977, 16'd58860, 16'd10786, 16'd47185, 16'd10713, 16'd59454, 16'd47202, 16'd62395, 16'd32851, 16'd30667, 16'd17969, 16'd59988, 16'd60090, 16'd49743});
	test_expansion(128'h43aa9244a14108e2fd560fc149a32e9f, {16'd60141, 16'd63611, 16'd64048, 16'd17763, 16'd26282, 16'd37077, 16'd18761, 16'd19911, 16'd22760, 16'd9293, 16'd41860, 16'd63221, 16'd28771, 16'd53999, 16'd20417, 16'd8392, 16'd32359, 16'd61007, 16'd52163, 16'd27462, 16'd13057, 16'd23049, 16'd47477, 16'd45821, 16'd50323, 16'd41514});
	test_expansion(128'hce29c5398418a6eed819995f51cdf2f0, {16'd65533, 16'd58028, 16'd5648, 16'd49318, 16'd1631, 16'd62219, 16'd8437, 16'd16733, 16'd54591, 16'd59662, 16'd43186, 16'd58431, 16'd12081, 16'd62730, 16'd58872, 16'd30275, 16'd3360, 16'd56188, 16'd2968, 16'd18762, 16'd27809, 16'd48645, 16'd13524, 16'd32610, 16'd36502, 16'd9384});
	test_expansion(128'h9f3059525385423f3f0136ad0ec71ccb, {16'd36172, 16'd35763, 16'd4225, 16'd60170, 16'd6921, 16'd48534, 16'd54994, 16'd25552, 16'd12631, 16'd2810, 16'd59553, 16'd48086, 16'd41776, 16'd64374, 16'd3288, 16'd61427, 16'd958, 16'd59556, 16'd19258, 16'd12992, 16'd58053, 16'd26273, 16'd50899, 16'd44278, 16'd4537, 16'd56895});
	test_expansion(128'h9ef8ce283d8ad2937a13db7bb58621df, {16'd13481, 16'd51508, 16'd25797, 16'd36050, 16'd25311, 16'd19975, 16'd10918, 16'd5625, 16'd38400, 16'd55147, 16'd63951, 16'd14463, 16'd26836, 16'd27068, 16'd6737, 16'd10800, 16'd276, 16'd64681, 16'd15145, 16'd57554, 16'd50244, 16'd12236, 16'd58584, 16'd29334, 16'd51904, 16'd44493});
	test_expansion(128'hdf7118e2d5822eeba5067d87ad98038f, {16'd40505, 16'd34511, 16'd45512, 16'd15421, 16'd15033, 16'd5809, 16'd9706, 16'd59663, 16'd15276, 16'd31277, 16'd42569, 16'd12039, 16'd24490, 16'd39217, 16'd24605, 16'd39833, 16'd53894, 16'd6524, 16'd13628, 16'd46000, 16'd29661, 16'd31518, 16'd5834, 16'd54273, 16'd30550, 16'd58126});
	test_expansion(128'h2b940907a714f3ee3658076510f11777, {16'd6019, 16'd12506, 16'd43283, 16'd57496, 16'd18482, 16'd10748, 16'd50739, 16'd50171, 16'd13363, 16'd44516, 16'd41666, 16'd42455, 16'd3175, 16'd23735, 16'd15475, 16'd58386, 16'd56597, 16'd45635, 16'd22054, 16'd35226, 16'd32659, 16'd28193, 16'd63726, 16'd58106, 16'd5115, 16'd26451});
	test_expansion(128'h292760a28edc1582c77c15da25abd45a, {16'd9226, 16'd62553, 16'd10269, 16'd10412, 16'd25705, 16'd57519, 16'd25921, 16'd8538, 16'd60389, 16'd28712, 16'd51570, 16'd23843, 16'd65387, 16'd57611, 16'd5359, 16'd12356, 16'd8788, 16'd15823, 16'd8754, 16'd14160, 16'd26176, 16'd34747, 16'd61882, 16'd36135, 16'd33374, 16'd29218});
	test_expansion(128'hf84ec004866d80816f079409ecabfbc5, {16'd60772, 16'd13862, 16'd39907, 16'd18414, 16'd39132, 16'd57206, 16'd64277, 16'd52754, 16'd60688, 16'd21141, 16'd35365, 16'd12891, 16'd7383, 16'd8460, 16'd46549, 16'd4719, 16'd49956, 16'd25255, 16'd14165, 16'd31251, 16'd29708, 16'd64685, 16'd25140, 16'd9880, 16'd10940, 16'd24848});
	test_expansion(128'ha557e321d14393bdf58f67881eea1726, {16'd27505, 16'd7581, 16'd26250, 16'd8126, 16'd62833, 16'd48966, 16'd57881, 16'd60396, 16'd39515, 16'd32903, 16'd3574, 16'd17920, 16'd22462, 16'd21402, 16'd36511, 16'd21823, 16'd14835, 16'd8661, 16'd57823, 16'd51089, 16'd55728, 16'd43026, 16'd1867, 16'd22524, 16'd14422, 16'd57076});
	test_expansion(128'hf380dc29df44fa7ead08eaff21aafe8b, {16'd27821, 16'd5190, 16'd51669, 16'd64426, 16'd38466, 16'd16831, 16'd10223, 16'd13887, 16'd55727, 16'd14812, 16'd38981, 16'd18787, 16'd41285, 16'd14261, 16'd26681, 16'd27020, 16'd55217, 16'd7531, 16'd27708, 16'd13513, 16'd5115, 16'd50936, 16'd54272, 16'd62851, 16'd37829, 16'd51868});
	test_expansion(128'h0d927369dd029d6b2d3fbbb8e0774441, {16'd26270, 16'd41485, 16'd17742, 16'd55194, 16'd28679, 16'd46532, 16'd14054, 16'd37173, 16'd777, 16'd6372, 16'd55369, 16'd29144, 16'd25646, 16'd65418, 16'd37844, 16'd16647, 16'd63007, 16'd47185, 16'd48385, 16'd1554, 16'd54077, 16'd902, 16'd46624, 16'd36652, 16'd30254, 16'd7936});
	test_expansion(128'h7b9f58502cd8e934d2a803864e1cf1cd, {16'd5138, 16'd38343, 16'd48837, 16'd49729, 16'd44372, 16'd56109, 16'd35926, 16'd27704, 16'd47023, 16'd46461, 16'd19933, 16'd33317, 16'd39555, 16'd54169, 16'd63235, 16'd37625, 16'd46331, 16'd10516, 16'd32245, 16'd37119, 16'd39425, 16'd18639, 16'd19185, 16'd29239, 16'd26763, 16'd33789});
	test_expansion(128'h001fb05775bb13c3c4cd1b9be6f76252, {16'd32850, 16'd1022, 16'd8290, 16'd44769, 16'd2956, 16'd63547, 16'd7621, 16'd12924, 16'd56793, 16'd34230, 16'd60099, 16'd52205, 16'd23210, 16'd22697, 16'd60902, 16'd38780, 16'd17016, 16'd14612, 16'd34556, 16'd62750, 16'd36348, 16'd45036, 16'd14185, 16'd60263, 16'd18885, 16'd18890});
	test_expansion(128'h5969be1f36a1d54f2ed1fa3a0d51844f, {16'd2802, 16'd36300, 16'd55574, 16'd18637, 16'd58994, 16'd32606, 16'd21808, 16'd15894, 16'd53137, 16'd34350, 16'd53693, 16'd10466, 16'd57889, 16'd30153, 16'd22124, 16'd61579, 16'd43688, 16'd64765, 16'd3738, 16'd52401, 16'd27762, 16'd50029, 16'd39394, 16'd44716, 16'd10792, 16'd39122});
	test_expansion(128'h991a01403c77f36524811c2d2ae0a5da, {16'd9915, 16'd34564, 16'd43681, 16'd54107, 16'd8681, 16'd64972, 16'd35231, 16'd8534, 16'd7432, 16'd51346, 16'd6770, 16'd50163, 16'd17239, 16'd51868, 16'd391, 16'd26190, 16'd23735, 16'd4400, 16'd49149, 16'd18572, 16'd59551, 16'd49041, 16'd31479, 16'd35877, 16'd26946, 16'd6171});
	test_expansion(128'hf7763f0da0a01dd5caa235ef2af1f6c2, {16'd18821, 16'd14035, 16'd44907, 16'd58359, 16'd54826, 16'd24827, 16'd27715, 16'd47491, 16'd12148, 16'd20467, 16'd50641, 16'd59424, 16'd43352, 16'd31314, 16'd5079, 16'd41084, 16'd11016, 16'd64192, 16'd62261, 16'd59891, 16'd20801, 16'd35168, 16'd37585, 16'd63969, 16'd4731, 16'd60095});
	test_expansion(128'h34cd2813a2ef44953fd93ec1477814b2, {16'd24672, 16'd56633, 16'd56811, 16'd23616, 16'd36082, 16'd14410, 16'd64950, 16'd37595, 16'd33282, 16'd58218, 16'd17475, 16'd51799, 16'd27960, 16'd31054, 16'd39894, 16'd63027, 16'd33719, 16'd29904, 16'd17631, 16'd28646, 16'd41839, 16'd19580, 16'd47881, 16'd6375, 16'd65062, 16'd44342});
	test_expansion(128'h74a880dba5d0d55adc58b3e9aaf5dc71, {16'd21175, 16'd55394, 16'd2458, 16'd55153, 16'd4322, 16'd4652, 16'd38809, 16'd60636, 16'd48644, 16'd61567, 16'd48907, 16'd47244, 16'd30424, 16'd27715, 16'd46758, 16'd21782, 16'd28169, 16'd31911, 16'd3729, 16'd19750, 16'd40775, 16'd54723, 16'd23343, 16'd46704, 16'd37078, 16'd53933});
	test_expansion(128'h2e1360967c8eb432475772b4064fa2e8, {16'd30900, 16'd26311, 16'd56903, 16'd16407, 16'd20129, 16'd21153, 16'd62737, 16'd27848, 16'd23618, 16'd46286, 16'd27787, 16'd2765, 16'd42294, 16'd2849, 16'd16692, 16'd26499, 16'd38452, 16'd10354, 16'd63411, 16'd3481, 16'd39960, 16'd24837, 16'd30875, 16'd54355, 16'd34506, 16'd12702});
	test_expansion(128'h703ffe223ab62264238d58515e32cd07, {16'd28324, 16'd17861, 16'd46985, 16'd34909, 16'd43405, 16'd25808, 16'd27169, 16'd30997, 16'd18344, 16'd294, 16'd34848, 16'd52343, 16'd21041, 16'd47841, 16'd53892, 16'd13045, 16'd51785, 16'd9300, 16'd60183, 16'd42904, 16'd24557, 16'd30073, 16'd14439, 16'd2849, 16'd49641, 16'd7633});
	test_expansion(128'ha464e385c6d373301cab6facbe428255, {16'd53078, 16'd43538, 16'd2244, 16'd24714, 16'd49992, 16'd47115, 16'd39789, 16'd65474, 16'd37399, 16'd18651, 16'd35625, 16'd55340, 16'd6996, 16'd58500, 16'd27707, 16'd20791, 16'd46481, 16'd41085, 16'd63523, 16'd19, 16'd11119, 16'd44816, 16'd54005, 16'd38631, 16'd35686, 16'd12312});
	test_expansion(128'ha520552ecbe0ddf2fe291078e4e0117c, {16'd35334, 16'd28002, 16'd6699, 16'd43515, 16'd48480, 16'd13502, 16'd32423, 16'd8504, 16'd60292, 16'd49876, 16'd16653, 16'd38884, 16'd22375, 16'd7952, 16'd9145, 16'd19616, 16'd3146, 16'd23372, 16'd22154, 16'd690, 16'd11190, 16'd33822, 16'd1994, 16'd661, 16'd17228, 16'd46548});
	test_expansion(128'h1954645b195113e4262673bc52a79c67, {16'd22108, 16'd7453, 16'd64338, 16'd36389, 16'd11158, 16'd17011, 16'd37314, 16'd4043, 16'd53793, 16'd49010, 16'd11765, 16'd39047, 16'd56899, 16'd41400, 16'd56444, 16'd35893, 16'd465, 16'd31443, 16'd47767, 16'd7158, 16'd41146, 16'd58214, 16'd45501, 16'd47993, 16'd23283, 16'd63219});
	test_expansion(128'h2bf5f9b739d6c3703c5507578503e803, {16'd25198, 16'd55369, 16'd32063, 16'd54634, 16'd8415, 16'd7587, 16'd58735, 16'd27709, 16'd25867, 16'd42887, 16'd46402, 16'd19269, 16'd43455, 16'd11368, 16'd45219, 16'd62248, 16'd51502, 16'd32766, 16'd45148, 16'd45742, 16'd38047, 16'd18275, 16'd1213, 16'd28426, 16'd26286, 16'd22153});
	test_expansion(128'hb0f38b4a2f7942ec05fa501bff40019a, {16'd6513, 16'd7672, 16'd18785, 16'd58642, 16'd18977, 16'd42771, 16'd52476, 16'd35635, 16'd11193, 16'd17650, 16'd26172, 16'd51281, 16'd38010, 16'd62762, 16'd32097, 16'd31431, 16'd25884, 16'd56116, 16'd17886, 16'd7197, 16'd32533, 16'd11473, 16'd60524, 16'd12382, 16'd51285, 16'd37574});
	test_expansion(128'h3635c58bd594690b46ef0f8e3340ee14, {16'd54596, 16'd14937, 16'd49471, 16'd64307, 16'd21518, 16'd41175, 16'd54387, 16'd61195, 16'd3013, 16'd21176, 16'd25112, 16'd29317, 16'd10821, 16'd21348, 16'd44606, 16'd33296, 16'd15224, 16'd41612, 16'd63599, 16'd63850, 16'd4891, 16'd13285, 16'd37217, 16'd59753, 16'd5526, 16'd33160});
	test_expansion(128'h8865e0567caf77300550d686b7e1692a, {16'd31194, 16'd42569, 16'd6406, 16'd56510, 16'd35124, 16'd291, 16'd52702, 16'd36704, 16'd53442, 16'd24636, 16'd20724, 16'd5755, 16'd48834, 16'd4690, 16'd27448, 16'd14484, 16'd31865, 16'd28858, 16'd39922, 16'd20083, 16'd8373, 16'd12676, 16'd29820, 16'd62010, 16'd29263, 16'd33247});
	test_expansion(128'h273d07d8679b9c11558b9011154857b0, {16'd33523, 16'd57530, 16'd21207, 16'd35949, 16'd60290, 16'd615, 16'd23903, 16'd44370, 16'd62945, 16'd58352, 16'd5532, 16'd18677, 16'd57644, 16'd39704, 16'd61164, 16'd3461, 16'd34437, 16'd56854, 16'd8929, 16'd27131, 16'd4256, 16'd33493, 16'd39329, 16'd35426, 16'd30993, 16'd56484});
	test_expansion(128'h7bfccff25d5fe6d732a71c779822a2c2, {16'd48640, 16'd62003, 16'd40992, 16'd52515, 16'd51878, 16'd36350, 16'd47350, 16'd21633, 16'd42433, 16'd3558, 16'd26837, 16'd3122, 16'd46087, 16'd50549, 16'd41806, 16'd49687, 16'd4192, 16'd45780, 16'd54457, 16'd62298, 16'd10805, 16'd57475, 16'd20740, 16'd26187, 16'd55378, 16'd58213});
	test_expansion(128'hb6c9959f0d5ef59a71423c9460757c31, {16'd40491, 16'd56302, 16'd55383, 16'd39926, 16'd59976, 16'd47552, 16'd55983, 16'd38693, 16'd51734, 16'd38908, 16'd42093, 16'd47085, 16'd38625, 16'd45328, 16'd21226, 16'd35002, 16'd10792, 16'd56609, 16'd33280, 16'd32823, 16'd24056, 16'd30523, 16'd23298, 16'd57333, 16'd44183, 16'd63568});
	test_expansion(128'h018d424a0036a4d0a7309a536c788516, {16'd18286, 16'd2393, 16'd9120, 16'd1206, 16'd54453, 16'd29118, 16'd12055, 16'd9952, 16'd16788, 16'd35534, 16'd40714, 16'd41329, 16'd42417, 16'd40435, 16'd53220, 16'd59674, 16'd7990, 16'd16772, 16'd23937, 16'd28863, 16'd8731, 16'd21722, 16'd11375, 16'd45028, 16'd44128, 16'd10751});
	test_expansion(128'h82d14e2247d5be9b2f75b09401cd088a, {16'd7376, 16'd55810, 16'd58538, 16'd56526, 16'd16337, 16'd23677, 16'd34715, 16'd4738, 16'd22719, 16'd18608, 16'd23583, 16'd35772, 16'd37326, 16'd40784, 16'd13035, 16'd21591, 16'd44372, 16'd12898, 16'd62430, 16'd35630, 16'd17832, 16'd42807, 16'd48708, 16'd7581, 16'd8631, 16'd29698});
	test_expansion(128'h62081ec135aa0100e126667559b1ec74, {16'd16814, 16'd32379, 16'd64598, 16'd38301, 16'd13926, 16'd2744, 16'd16550, 16'd4814, 16'd33477, 16'd65266, 16'd9306, 16'd28658, 16'd28928, 16'd14075, 16'd62302, 16'd607, 16'd2227, 16'd57491, 16'd59198, 16'd34544, 16'd57546, 16'd45242, 16'd24042, 16'd58694, 16'd26421, 16'd35276});
	test_expansion(128'h0a3d575578fed61e62ab442d10322ef9, {16'd44079, 16'd54378, 16'd50921, 16'd63867, 16'd35730, 16'd28122, 16'd43599, 16'd7701, 16'd37277, 16'd60061, 16'd56162, 16'd9920, 16'd22855, 16'd17953, 16'd25264, 16'd29896, 16'd11907, 16'd19323, 16'd37775, 16'd44717, 16'd30327, 16'd32391, 16'd37554, 16'd7562, 16'd63830, 16'd7133});
	test_expansion(128'h6a51c8ee142f46343f4692e29d4a17d4, {16'd15376, 16'd20630, 16'd55443, 16'd3680, 16'd54707, 16'd36389, 16'd40855, 16'd21293, 16'd29345, 16'd31868, 16'd62855, 16'd38641, 16'd50061, 16'd33372, 16'd17210, 16'd21527, 16'd39700, 16'd14702, 16'd48637, 16'd52220, 16'd19869, 16'd18677, 16'd30561, 16'd10135, 16'd16302, 16'd26852});
	test_expansion(128'h3006e6ca491ed327e39909d7c9fe27c3, {16'd5397, 16'd2379, 16'd34810, 16'd65387, 16'd27193, 16'd29093, 16'd36569, 16'd32417, 16'd45599, 16'd26124, 16'd32952, 16'd56245, 16'd51923, 16'd45167, 16'd34043, 16'd2194, 16'd1334, 16'd54421, 16'd24620, 16'd26501, 16'd32603, 16'd28980, 16'd16471, 16'd22569, 16'd23765, 16'd22430});
	test_expansion(128'h5e1560c765ed0d3eb172d9ecb05d5658, {16'd22701, 16'd18880, 16'd35783, 16'd46822, 16'd20809, 16'd41800, 16'd32898, 16'd24856, 16'd62442, 16'd47267, 16'd39779, 16'd14128, 16'd29843, 16'd56036, 16'd55316, 16'd44108, 16'd35176, 16'd54982, 16'd33414, 16'd56461, 16'd54016, 16'd59693, 16'd16571, 16'd37912, 16'd62638, 16'd44663});
	test_expansion(128'h9579d25771d8d2828f97b94a3c5e4958, {16'd52103, 16'd46643, 16'd29587, 16'd34283, 16'd38, 16'd44357, 16'd27133, 16'd33486, 16'd64150, 16'd44599, 16'd27264, 16'd58514, 16'd48509, 16'd52631, 16'd31535, 16'd4612, 16'd44750, 16'd40692, 16'd34886, 16'd40015, 16'd50383, 16'd31780, 16'd55044, 16'd45515, 16'd20258, 16'd63432});
	test_expansion(128'hc01700786a024c26a9c88148e4d62912, {16'd5882, 16'd47851, 16'd49389, 16'd46983, 16'd54247, 16'd2766, 16'd38721, 16'd43324, 16'd31542, 16'd37697, 16'd10043, 16'd16247, 16'd65459, 16'd56960, 16'd36963, 16'd39690, 16'd41377, 16'd63814, 16'd20130, 16'd32165, 16'd54143, 16'd60923, 16'd44133, 16'd30269, 16'd27117, 16'd1473});
	test_expansion(128'hf74c6fc5c8299f656140223a0797ede8, {16'd40359, 16'd41157, 16'd13660, 16'd40578, 16'd25581, 16'd22641, 16'd5224, 16'd49711, 16'd23112, 16'd61, 16'd3409, 16'd55642, 16'd5963, 16'd51635, 16'd58598, 16'd4430, 16'd34422, 16'd53447, 16'd47706, 16'd26807, 16'd23557, 16'd2743, 16'd42637, 16'd17286, 16'd54818, 16'd396});
	test_expansion(128'hb992c880f6d1b3db19e81701dc7533b1, {16'd20003, 16'd7939, 16'd26336, 16'd20789, 16'd56895, 16'd16886, 16'd33886, 16'd55634, 16'd15026, 16'd42870, 16'd20288, 16'd15983, 16'd44776, 16'd24936, 16'd60949, 16'd53150, 16'd23217, 16'd52448, 16'd22815, 16'd58774, 16'd9897, 16'd25388, 16'd62931, 16'd29986, 16'd61687, 16'd24397});
	test_expansion(128'h352843d0d63c469504b5cd3310bf3277, {16'd37725, 16'd1032, 16'd10459, 16'd56478, 16'd6969, 16'd50875, 16'd3786, 16'd58970, 16'd4448, 16'd16852, 16'd42583, 16'd54120, 16'd298, 16'd60635, 16'd57429, 16'd12786, 16'd62554, 16'd56683, 16'd16983, 16'd13394, 16'd58443, 16'd32244, 16'd15897, 16'd31931, 16'd48735, 16'd7426});
	test_expansion(128'h8c4ee630edb7c52c2b006e60a15fbd58, {16'd36265, 16'd27260, 16'd63895, 16'd50993, 16'd50359, 16'd38939, 16'd47415, 16'd18463, 16'd31684, 16'd21019, 16'd59735, 16'd48331, 16'd25943, 16'd19368, 16'd35147, 16'd3086, 16'd25902, 16'd58266, 16'd7185, 16'd30795, 16'd43125, 16'd51785, 16'd38414, 16'd15621, 16'd62845, 16'd27636});
	test_expansion(128'hde3d4e98cd4715b491ee256bde4c350a, {16'd65013, 16'd29435, 16'd6088, 16'd16155, 16'd11520, 16'd5290, 16'd41295, 16'd44829, 16'd7188, 16'd62155, 16'd48034, 16'd23639, 16'd34066, 16'd11669, 16'd28712, 16'd62798, 16'd31425, 16'd39656, 16'd7552, 16'd43588, 16'd11479, 16'd60465, 16'd63864, 16'd57594, 16'd17006, 16'd56960});
	test_expansion(128'he54d72384801f60cbf810f9b0e34551f, {16'd18644, 16'd49921, 16'd62583, 16'd36119, 16'd60237, 16'd2161, 16'd16353, 16'd61754, 16'd37112, 16'd61622, 16'd47951, 16'd35324, 16'd31229, 16'd25342, 16'd65407, 16'd56679, 16'd36310, 16'd50679, 16'd13884, 16'd17312, 16'd48690, 16'd31311, 16'd6193, 16'd26491, 16'd52353, 16'd42861});
	test_expansion(128'hb94b9effa081e3c8f8bf6c1bfa97445c, {16'd29860, 16'd53866, 16'd2400, 16'd34591, 16'd36883, 16'd17470, 16'd59941, 16'd40439, 16'd41425, 16'd14843, 16'd49720, 16'd12223, 16'd46446, 16'd26401, 16'd40283, 16'd1623, 16'd2658, 16'd14263, 16'd50323, 16'd58630, 16'd26254, 16'd15169, 16'd6182, 16'd54732, 16'd46329, 16'd17947});
	test_expansion(128'he8ec094b78f792b520f79c8875db5944, {16'd2156, 16'd36173, 16'd64886, 16'd16899, 16'd54795, 16'd3862, 16'd50363, 16'd37671, 16'd8696, 16'd31400, 16'd1303, 16'd28539, 16'd19177, 16'd57578, 16'd61175, 16'd42146, 16'd112, 16'd32194, 16'd32714, 16'd59092, 16'd25659, 16'd36339, 16'd40347, 16'd14447, 16'd5850, 16'd38177});
	test_expansion(128'h6b76af9955487d71a1850b5588ebc063, {16'd43141, 16'd17811, 16'd17039, 16'd19614, 16'd9139, 16'd61309, 16'd62995, 16'd17413, 16'd30857, 16'd25038, 16'd44287, 16'd4993, 16'd34246, 16'd58770, 16'd1452, 16'd38729, 16'd23701, 16'd12540, 16'd47328, 16'd42976, 16'd29846, 16'd42490, 16'd33627, 16'd7479, 16'd50289, 16'd17855});
	test_expansion(128'h0421871b0203c2999fdaaf6b2c649fc2, {16'd44319, 16'd59791, 16'd54720, 16'd4787, 16'd7919, 16'd51556, 16'd37475, 16'd35762, 16'd23865, 16'd41542, 16'd52203, 16'd13249, 16'd55744, 16'd14444, 16'd60728, 16'd43186, 16'd11991, 16'd19899, 16'd48761, 16'd52195, 16'd24751, 16'd655, 16'd23089, 16'd28644, 16'd15871, 16'd47613});
	test_expansion(128'hdc2af203218c487cd77f373a138c853c, {16'd13186, 16'd35396, 16'd58959, 16'd48391, 16'd35982, 16'd37780, 16'd36411, 16'd46528, 16'd52136, 16'd41667, 16'd21800, 16'd49672, 16'd3722, 16'd46620, 16'd25200, 16'd63083, 16'd48836, 16'd50562, 16'd39631, 16'd21600, 16'd16237, 16'd42628, 16'd21563, 16'd50718, 16'd11564, 16'd57099});
	test_expansion(128'hdb01edd3cabe869491231fe886eceaf5, {16'd32660, 16'd52063, 16'd62525, 16'd15708, 16'd60716, 16'd50098, 16'd25360, 16'd61167, 16'd53599, 16'd2407, 16'd29043, 16'd30641, 16'd55480, 16'd56664, 16'd21272, 16'd19152, 16'd42360, 16'd25456, 16'd48047, 16'd19074, 16'd19397, 16'd54446, 16'd17636, 16'd52572, 16'd28084, 16'd60178});
	test_expansion(128'h02c928f0be1c1a4ad1fa53622f892e00, {16'd36016, 16'd23108, 16'd2357, 16'd13055, 16'd8646, 16'd39112, 16'd20468, 16'd22000, 16'd38355, 16'd34841, 16'd45616, 16'd64533, 16'd34507, 16'd10492, 16'd6227, 16'd3803, 16'd37703, 16'd52009, 16'd7231, 16'd19565, 16'd9378, 16'd6515, 16'd13118, 16'd9344, 16'd29115, 16'd54687});
	test_expansion(128'hb3982fa977803f85987a672a6250a389, {16'd58540, 16'd46476, 16'd15997, 16'd15751, 16'd40667, 16'd55676, 16'd56882, 16'd16832, 16'd35493, 16'd42517, 16'd10024, 16'd22382, 16'd32000, 16'd62651, 16'd24319, 16'd42939, 16'd56879, 16'd40694, 16'd19384, 16'd52223, 16'd24823, 16'd21833, 16'd61631, 16'd13932, 16'd27454, 16'd3560});
	test_expansion(128'h8470b379d741b7946dec307d2a83d047, {16'd3557, 16'd6463, 16'd61841, 16'd17241, 16'd58977, 16'd8858, 16'd38730, 16'd15575, 16'd47480, 16'd2360, 16'd38408, 16'd16002, 16'd29828, 16'd5097, 16'd3361, 16'd8690, 16'd45221, 16'd16209, 16'd47520, 16'd44282, 16'd57861, 16'd35001, 16'd31622, 16'd26592, 16'd33667, 16'd43867});
	test_expansion(128'h5037f4d76d705448a2f6ee41c6d87b53, {16'd41586, 16'd28887, 16'd51656, 16'd16913, 16'd38169, 16'd8979, 16'd23914, 16'd48226, 16'd12826, 16'd19817, 16'd40949, 16'd14761, 16'd1571, 16'd59930, 16'd35126, 16'd17266, 16'd49487, 16'd6130, 16'd18787, 16'd19804, 16'd40795, 16'd10971, 16'd55737, 16'd40267, 16'd32361, 16'd42519});
	test_expansion(128'h013cb97c4adcd922b7ffcb0153013871, {16'd10593, 16'd62436, 16'd55627, 16'd55091, 16'd44051, 16'd57292, 16'd6671, 16'd15507, 16'd36521, 16'd22988, 16'd24984, 16'd20458, 16'd25614, 16'd18438, 16'd816, 16'd56902, 16'd52834, 16'd7300, 16'd22614, 16'd58803, 16'd32141, 16'd993, 16'd59257, 16'd35447, 16'd62521, 16'd27790});
	test_expansion(128'h087037eae04a1cf7b5449ffadd9f37cb, {16'd34733, 16'd63262, 16'd57926, 16'd10730, 16'd45127, 16'd28105, 16'd30525, 16'd30280, 16'd34290, 16'd7998, 16'd30294, 16'd48219, 16'd11864, 16'd48040, 16'd37090, 16'd7201, 16'd3642, 16'd56008, 16'd19903, 16'd33683, 16'd965, 16'd59783, 16'd7700, 16'd38729, 16'd37199, 16'd57074});
	test_expansion(128'hd1688b10ec971cf3ec2eea00bbdbd831, {16'd4537, 16'd50851, 16'd5032, 16'd14348, 16'd38325, 16'd49815, 16'd20275, 16'd15611, 16'd37801, 16'd42876, 16'd29809, 16'd29911, 16'd23759, 16'd10285, 16'd20064, 16'd44368, 16'd5967, 16'd14106, 16'd7362, 16'd53828, 16'd38687, 16'd64590, 16'd22049, 16'd27237, 16'd42616, 16'd41032});
	test_expansion(128'h5b9ea5978682156810bc0afaddd0e184, {16'd40366, 16'd53897, 16'd18874, 16'd30314, 16'd34632, 16'd5528, 16'd37715, 16'd10479, 16'd9944, 16'd8203, 16'd48943, 16'd57500, 16'd53212, 16'd34355, 16'd51970, 16'd63541, 16'd46943, 16'd27435, 16'd5276, 16'd38608, 16'd40229, 16'd35263, 16'd24894, 16'd52215, 16'd29032, 16'd30019});
	test_expansion(128'hd8311ea1e8a379d59c3f454fa63ef7df, {16'd292, 16'd36375, 16'd60804, 16'd16335, 16'd46600, 16'd37789, 16'd13866, 16'd51456, 16'd9921, 16'd22166, 16'd46607, 16'd12784, 16'd23314, 16'd62804, 16'd40745, 16'd61371, 16'd45985, 16'd49252, 16'd55442, 16'd19688, 16'd45172, 16'd13807, 16'd13277, 16'd61672, 16'd41994, 16'd23186});
	test_expansion(128'h97ad2ea3fead5474c2357575e1837be3, {16'd26882, 16'd9465, 16'd55310, 16'd34630, 16'd45942, 16'd22989, 16'd16913, 16'd48478, 16'd31979, 16'd38011, 16'd47548, 16'd10791, 16'd7716, 16'd53245, 16'd683, 16'd12813, 16'd52540, 16'd51241, 16'd22893, 16'd26053, 16'd35060, 16'd21988, 16'd7223, 16'd29614, 16'd63317, 16'd4848});
	test_expansion(128'hfba3238bca5d8d3d87cebda523ba3a3f, {16'd55527, 16'd38270, 16'd58966, 16'd52463, 16'd33667, 16'd21481, 16'd27221, 16'd43906, 16'd13537, 16'd1660, 16'd41444, 16'd48866, 16'd584, 16'd19995, 16'd34216, 16'd58633, 16'd9877, 16'd51199, 16'd59038, 16'd42222, 16'd57993, 16'd14619, 16'd18010, 16'd32322, 16'd47042, 16'd20638});
	test_expansion(128'h95949ef2229e87be3b7d2898abdaef77, {16'd4031, 16'd30315, 16'd43738, 16'd19158, 16'd15878, 16'd21868, 16'd53365, 16'd41272, 16'd58537, 16'd34014, 16'd8719, 16'd35084, 16'd22093, 16'd7364, 16'd11981, 16'd31075, 16'd32374, 16'd35657, 16'd46088, 16'd14886, 16'd32095, 16'd14831, 16'd17504, 16'd19728, 16'd55105, 16'd43860});
	test_expansion(128'h3af16b68d9fd8274e5359b02a38a141c, {16'd20558, 16'd611, 16'd37452, 16'd28370, 16'd44178, 16'd9023, 16'd47574, 16'd17214, 16'd47551, 16'd38339, 16'd27544, 16'd51221, 16'd53647, 16'd7428, 16'd32102, 16'd12270, 16'd37112, 16'd62050, 16'd13441, 16'd37994, 16'd61706, 16'd12823, 16'd10977, 16'd28589, 16'd51394, 16'd43551});
	test_expansion(128'h648a6e6b5a3aea2a0e7544d8d32e1940, {16'd41378, 16'd42666, 16'd24398, 16'd24101, 16'd526, 16'd32402, 16'd38257, 16'd20604, 16'd20853, 16'd14874, 16'd56196, 16'd37590, 16'd41178, 16'd18372, 16'd15780, 16'd18094, 16'd9172, 16'd15990, 16'd15194, 16'd22502, 16'd40502, 16'd41608, 16'd8485, 16'd4642, 16'd42081, 16'd55286});
	test_expansion(128'h03828481bb1392f5758fbca60adf2135, {16'd62396, 16'd19971, 16'd14459, 16'd23581, 16'd26938, 16'd49107, 16'd45479, 16'd40798, 16'd40070, 16'd20622, 16'd24964, 16'd14562, 16'd43517, 16'd64059, 16'd12227, 16'd37309, 16'd51961, 16'd10001, 16'd22589, 16'd30822, 16'd6727, 16'd6090, 16'd45018, 16'd53889, 16'd36532, 16'd59466});
	test_expansion(128'h9702052a03b8efc5519aaabb771e1001, {16'd55146, 16'd63476, 16'd24762, 16'd43118, 16'd48166, 16'd35178, 16'd51126, 16'd34674, 16'd46160, 16'd50425, 16'd20814, 16'd24815, 16'd17859, 16'd12410, 16'd51743, 16'd5964, 16'd49177, 16'd42658, 16'd51347, 16'd22041, 16'd62359, 16'd2556, 16'd8384, 16'd23951, 16'd29709, 16'd6198});
	test_expansion(128'h4b0ddc3d296d92de3c8884ef542d9f85, {16'd31894, 16'd15653, 16'd38210, 16'd9815, 16'd2014, 16'd23052, 16'd22272, 16'd16462, 16'd49282, 16'd59441, 16'd32341, 16'd36100, 16'd52399, 16'd1863, 16'd63457, 16'd63518, 16'd61643, 16'd62081, 16'd6556, 16'd12189, 16'd30712, 16'd55120, 16'd13976, 16'd20421, 16'd51591, 16'd3082});
	test_expansion(128'h5f750492540e2e4e5fe7c16839a75107, {16'd52970, 16'd6465, 16'd61803, 16'd47969, 16'd39580, 16'd11664, 16'd17633, 16'd39892, 16'd37631, 16'd39510, 16'd23164, 16'd58955, 16'd36325, 16'd41011, 16'd27778, 16'd4058, 16'd57940, 16'd18483, 16'd29746, 16'd15141, 16'd59445, 16'd55480, 16'd64107, 16'd54318, 16'd22470, 16'd28291});
	test_expansion(128'h259a3fb3b3cdd619a569fe90b59e6c77, {16'd64537, 16'd15041, 16'd12959, 16'd59570, 16'd63145, 16'd41861, 16'd15082, 16'd43113, 16'd47489, 16'd35713, 16'd40575, 16'd15494, 16'd7367, 16'd29272, 16'd38709, 16'd23602, 16'd41398, 16'd42731, 16'd22823, 16'd64466, 16'd49984, 16'd40268, 16'd31083, 16'd2483, 16'd40315, 16'd56376});
	test_expansion(128'h8417188b98d78741a57fe23ff18f6fbf, {16'd10926, 16'd8703, 16'd102, 16'd10144, 16'd45226, 16'd39954, 16'd58114, 16'd29212, 16'd17039, 16'd45755, 16'd1913, 16'd33884, 16'd43713, 16'd45017, 16'd54032, 16'd5785, 16'd56992, 16'd39971, 16'd42148, 16'd2878, 16'd20673, 16'd37282, 16'd28968, 16'd37576, 16'd17631, 16'd58762});
	test_expansion(128'h6c47b6239c1854b8dafdbe00a9ca8bda, {16'd10629, 16'd15880, 16'd38914, 16'd44773, 16'd55839, 16'd44696, 16'd8064, 16'd33257, 16'd16682, 16'd10594, 16'd17511, 16'd694, 16'd62024, 16'd57128, 16'd21219, 16'd13453, 16'd49531, 16'd57619, 16'd41404, 16'd31224, 16'd42432, 16'd33400, 16'd27176, 16'd64916, 16'd58697, 16'd64209});
	test_expansion(128'hf6bf1dd634c34c2ac2eb0a06f4992409, {16'd17126, 16'd55770, 16'd59989, 16'd55764, 16'd31042, 16'd21236, 16'd29392, 16'd65505, 16'd35582, 16'd30570, 16'd35603, 16'd45445, 16'd48537, 16'd33681, 16'd31485, 16'd41304, 16'd29469, 16'd32895, 16'd20600, 16'd21583, 16'd15257, 16'd6577, 16'd51995, 16'd17973, 16'd6093, 16'd15458});
	test_expansion(128'h0c106c38652d52b5e8454abc3a2814ce, {16'd33817, 16'd3507, 16'd6929, 16'd39985, 16'd2287, 16'd64336, 16'd32574, 16'd29205, 16'd4750, 16'd34484, 16'd12185, 16'd62909, 16'd27742, 16'd34524, 16'd59564, 16'd55892, 16'd42075, 16'd37507, 16'd45029, 16'd48903, 16'd37381, 16'd46520, 16'd51894, 16'd8881, 16'd46163, 16'd36029});
	test_expansion(128'h31796c3ec8ed8c116fe8c710bca41924, {16'd40645, 16'd47468, 16'd52628, 16'd2086, 16'd54396, 16'd34670, 16'd45565, 16'd15829, 16'd33131, 16'd41005, 16'd62862, 16'd56691, 16'd63025, 16'd16478, 16'd64775, 16'd6225, 16'd34813, 16'd56181, 16'd29852, 16'd24855, 16'd32490, 16'd1619, 16'd9171, 16'd15316, 16'd5279, 16'd14416});
	test_expansion(128'he8b63b0c8fb9a19b1fae559ff32d7703, {16'd32620, 16'd20039, 16'd64246, 16'd45717, 16'd9939, 16'd39282, 16'd20409, 16'd36609, 16'd20694, 16'd43063, 16'd59877, 16'd18345, 16'd14339, 16'd15576, 16'd58381, 16'd26946, 16'd20921, 16'd25233, 16'd14235, 16'd55586, 16'd30724, 16'd22538, 16'd57990, 16'd54906, 16'd37541, 16'd41487});
	test_expansion(128'h7a97e56aea60ed89c8f24511614b42fd, {16'd3563, 16'd39208, 16'd63908, 16'd45049, 16'd59029, 16'd8011, 16'd35181, 16'd13441, 16'd23618, 16'd56084, 16'd58703, 16'd1481, 16'd3916, 16'd24987, 16'd43740, 16'd9078, 16'd6054, 16'd8281, 16'd39281, 16'd59084, 16'd14608, 16'd46268, 16'd63441, 16'd4161, 16'd65394, 16'd48282});
	test_expansion(128'h9bbd06a4a9e123ca1e604e885d3acf80, {16'd42239, 16'd24537, 16'd19356, 16'd10261, 16'd30112, 16'd7817, 16'd7911, 16'd16124, 16'd61412, 16'd19179, 16'd11428, 16'd30013, 16'd52599, 16'd51684, 16'd11195, 16'd40098, 16'd15834, 16'd7705, 16'd43351, 16'd38790, 16'd6251, 16'd63777, 16'd4170, 16'd30780, 16'd7377, 16'd18699});
	test_expansion(128'h12132bd438115f459a8b48ef25598834, {16'd48142, 16'd2584, 16'd30936, 16'd40083, 16'd51891, 16'd44981, 16'd25510, 16'd11070, 16'd58488, 16'd27958, 16'd17732, 16'd50684, 16'd30992, 16'd37912, 16'd25033, 16'd58699, 16'd13402, 16'd28816, 16'd13136, 16'd30000, 16'd31887, 16'd21120, 16'd43109, 16'd38607, 16'd63318, 16'd30914});
	test_expansion(128'hbb15afc32d3f241afc144dd020d75098, {16'd17224, 16'd30633, 16'd53685, 16'd4884, 16'd57592, 16'd9926, 16'd5089, 16'd3250, 16'd13376, 16'd38064, 16'd50268, 16'd35581, 16'd63185, 16'd24402, 16'd19896, 16'd38924, 16'd42542, 16'd51539, 16'd10800, 16'd1173, 16'd58137, 16'd16354, 16'd55144, 16'd33835, 16'd437, 16'd27033});
	test_expansion(128'hb4d8ccd986f354b2952108070661d422, {16'd41786, 16'd12929, 16'd65109, 16'd22703, 16'd47722, 16'd57300, 16'd4777, 16'd49519, 16'd63352, 16'd46836, 16'd29921, 16'd42143, 16'd62552, 16'd25485, 16'd26992, 16'd5180, 16'd18891, 16'd12358, 16'd4990, 16'd57488, 16'd28357, 16'd28497, 16'd7607, 16'd50144, 16'd33092, 16'd17661});
	test_expansion(128'h466eb3bdb68573264613c1abbb16ae0d, {16'd46809, 16'd25661, 16'd53459, 16'd50628, 16'd16775, 16'd5078, 16'd41264, 16'd29610, 16'd11579, 16'd8489, 16'd40825, 16'd6739, 16'd63645, 16'd30368, 16'd25028, 16'd45079, 16'd46483, 16'd37378, 16'd17105, 16'd6361, 16'd49268, 16'd22110, 16'd54195, 16'd22693, 16'd24247, 16'd40752});
	test_expansion(128'he1f894701e5d2d85690fbcc4b2d965a3, {16'd47442, 16'd20423, 16'd21802, 16'd32274, 16'd42567, 16'd26026, 16'd46014, 16'd18287, 16'd50233, 16'd10418, 16'd35602, 16'd37393, 16'd51344, 16'd36394, 16'd52973, 16'd36215, 16'd48532, 16'd2994, 16'd64000, 16'd24613, 16'd24648, 16'd37492, 16'd4972, 16'd59027, 16'd29310, 16'd3262});
	test_expansion(128'h6668b62d20a9bb824ab2dc42bdafc7fd, {16'd51544, 16'd57900, 16'd33855, 16'd15633, 16'd35641, 16'd16318, 16'd12133, 16'd53262, 16'd3551, 16'd54621, 16'd19529, 16'd55101, 16'd49490, 16'd21564, 16'd15938, 16'd11590, 16'd56717, 16'd22016, 16'd19540, 16'd60262, 16'd4758, 16'd51901, 16'd12731, 16'd12326, 16'd25173, 16'd43951});
	test_expansion(128'h742c981da54ace05133435e76e756063, {16'd31981, 16'd44635, 16'd11978, 16'd55412, 16'd57524, 16'd43868, 16'd45623, 16'd9115, 16'd30427, 16'd64045, 16'd40173, 16'd30118, 16'd65010, 16'd22527, 16'd65149, 16'd14275, 16'd49771, 16'd21397, 16'd43669, 16'd57830, 16'd11195, 16'd38952, 16'd28098, 16'd9950, 16'd39133, 16'd58886});
	test_expansion(128'hedbcc3026b29e55478c8cfbb4ec82a28, {16'd34264, 16'd37519, 16'd11099, 16'd18578, 16'd63401, 16'd57600, 16'd11306, 16'd58129, 16'd28874, 16'd40806, 16'd417, 16'd48029, 16'd20898, 16'd50925, 16'd14671, 16'd47275, 16'd47447, 16'd61784, 16'd15928, 16'd44250, 16'd3702, 16'd55675, 16'd54667, 16'd38834, 16'd42874, 16'd7070});
	test_expansion(128'h001bc284782f20cb282e882b456669e8, {16'd34149, 16'd108, 16'd7928, 16'd31057, 16'd11746, 16'd60985, 16'd64568, 16'd9190, 16'd13297, 16'd22078, 16'd28055, 16'd3061, 16'd40504, 16'd10965, 16'd29121, 16'd58086, 16'd24404, 16'd12769, 16'd6451, 16'd17560, 16'd54199, 16'd9358, 16'd48570, 16'd7752, 16'd60608, 16'd35411});
	test_expansion(128'h78108a1533fa8bab162e88c19633249d, {16'd1654, 16'd36278, 16'd54158, 16'd1968, 16'd35318, 16'd59598, 16'd61432, 16'd6215, 16'd35864, 16'd44937, 16'd37224, 16'd35788, 16'd16889, 16'd31261, 16'd27567, 16'd37290, 16'd54611, 16'd5762, 16'd43731, 16'd22267, 16'd32769, 16'd31321, 16'd20952, 16'd56815, 16'd55769, 16'd16869});
	test_expansion(128'h7c429370c630e72458e36ffc9600a9f6, {16'd45143, 16'd19722, 16'd48865, 16'd23556, 16'd25531, 16'd1180, 16'd5082, 16'd1570, 16'd21866, 16'd5941, 16'd20121, 16'd61105, 16'd55622, 16'd49348, 16'd14416, 16'd30403, 16'd52991, 16'd61059, 16'd63629, 16'd30500, 16'd4440, 16'd57146, 16'd16417, 16'd5402, 16'd53369, 16'd61465});
	test_expansion(128'h6cccfc0fa9f4670b4aa8cbf559972fee, {16'd59361, 16'd41987, 16'd53413, 16'd33474, 16'd45023, 16'd2400, 16'd32033, 16'd28157, 16'd49516, 16'd38959, 16'd61012, 16'd24027, 16'd61276, 16'd29185, 16'd63497, 16'd45750, 16'd49812, 16'd36018, 16'd41476, 16'd61898, 16'd49077, 16'd9791, 16'd42971, 16'd59497, 16'd48930, 16'd22636});
	test_expansion(128'hd32d46f65c97de286f0727a669128cb4, {16'd57200, 16'd4296, 16'd22475, 16'd56309, 16'd59993, 16'd59701, 16'd19256, 16'd40065, 16'd45109, 16'd17579, 16'd32196, 16'd16580, 16'd13260, 16'd9420, 16'd18200, 16'd22887, 16'd63014, 16'd46157, 16'd56135, 16'd18, 16'd43595, 16'd42862, 16'd30878, 16'd20214, 16'd14132, 16'd18860});
	test_expansion(128'h43ad0b3834a959e106a502aad2861f2e, {16'd30623, 16'd55190, 16'd34982, 16'd62225, 16'd30705, 16'd39242, 16'd22937, 16'd51117, 16'd16023, 16'd42948, 16'd39864, 16'd33991, 16'd21340, 16'd63526, 16'd52406, 16'd34174, 16'd60206, 16'd17519, 16'd13466, 16'd47896, 16'd32032, 16'd9212, 16'd26598, 16'd65523, 16'd39050, 16'd28400});
	test_expansion(128'hc6dfa531a7c6ce259d4188975b449103, {16'd30913, 16'd52713, 16'd1117, 16'd61387, 16'd63087, 16'd2209, 16'd63219, 16'd38040, 16'd19406, 16'd59102, 16'd11322, 16'd52894, 16'd47141, 16'd11916, 16'd45728, 16'd4036, 16'd36727, 16'd41515, 16'd13431, 16'd47938, 16'd46194, 16'd33395, 16'd17015, 16'd38803, 16'd56928, 16'd4737});
	test_expansion(128'hac272c204168602cf5787c2271b3d625, {16'd37419, 16'd21340, 16'd36361, 16'd48959, 16'd50258, 16'd44349, 16'd27713, 16'd12003, 16'd16146, 16'd42407, 16'd58056, 16'd48711, 16'd7292, 16'd55719, 16'd33295, 16'd46165, 16'd212, 16'd56255, 16'd41064, 16'd56473, 16'd28311, 16'd52850, 16'd43778, 16'd41784, 16'd16276, 16'd61787});
	test_expansion(128'hfc7bbfb60a0a5606eb5716636139868b, {16'd10096, 16'd47758, 16'd32201, 16'd32991, 16'd63685, 16'd57322, 16'd27211, 16'd2904, 16'd21930, 16'd14970, 16'd20595, 16'd53642, 16'd17468, 16'd14166, 16'd11995, 16'd50559, 16'd18966, 16'd14043, 16'd51521, 16'd52525, 16'd54223, 16'd8408, 16'd35421, 16'd21517, 16'd57884, 16'd40550});
	test_expansion(128'hd1797c753a05ef2363f4d21713ce35ff, {16'd19815, 16'd34249, 16'd21065, 16'd27989, 16'd8169, 16'd36712, 16'd46471, 16'd55395, 16'd18439, 16'd8806, 16'd8018, 16'd41740, 16'd44331, 16'd21371, 16'd35625, 16'd54570, 16'd4089, 16'd35222, 16'd22100, 16'd12020, 16'd11795, 16'd21324, 16'd42106, 16'd31052, 16'd27488, 16'd5936});
	test_expansion(128'hba4e9292aa8abb8dc2dabcabb523bef8, {16'd58739, 16'd20615, 16'd50175, 16'd33787, 16'd7787, 16'd40033, 16'd52418, 16'd12291, 16'd26001, 16'd9557, 16'd21999, 16'd15996, 16'd14664, 16'd5280, 16'd43681, 16'd55547, 16'd60023, 16'd5367, 16'd52147, 16'd35887, 16'd8, 16'd9568, 16'd50002, 16'd39672, 16'd38887, 16'd26515});
	test_expansion(128'hecc3981983fde6f26930f77bda7591e7, {16'd44632, 16'd28016, 16'd20994, 16'd42768, 16'd7320, 16'd26003, 16'd3300, 16'd15102, 16'd62716, 16'd63963, 16'd35033, 16'd7465, 16'd32289, 16'd14051, 16'd15948, 16'd29900, 16'd24417, 16'd24406, 16'd36458, 16'd42769, 16'd54892, 16'd57995, 16'd39408, 16'd1688, 16'd21548, 16'd51335});
	test_expansion(128'hec0a5faf710a849331b5ec6ef19c3ad0, {16'd51706, 16'd48053, 16'd20154, 16'd18542, 16'd64290, 16'd13477, 16'd26753, 16'd26422, 16'd43706, 16'd49657, 16'd19080, 16'd16229, 16'd18808, 16'd35797, 16'd25904, 16'd41433, 16'd6820, 16'd24300, 16'd13493, 16'd23820, 16'd24990, 16'd5591, 16'd25588, 16'd1435, 16'd10732, 16'd23612});
	test_expansion(128'hf2e6b8eb642b5275660d11e7d0fdb8fd, {16'd282, 16'd46644, 16'd25533, 16'd64543, 16'd32224, 16'd32180, 16'd51976, 16'd27719, 16'd29227, 16'd19133, 16'd24718, 16'd43659, 16'd36242, 16'd35287, 16'd64303, 16'd44734, 16'd60648, 16'd10717, 16'd53983, 16'd22263, 16'd19665, 16'd24348, 16'd44340, 16'd32978, 16'd25326, 16'd21920});
	test_expansion(128'h19506b8c94e226a5aefc4bec2a7f6bb7, {16'd22679, 16'd60330, 16'd10602, 16'd37951, 16'd16288, 16'd54158, 16'd58910, 16'd26786, 16'd23955, 16'd33222, 16'd57331, 16'd26817, 16'd14873, 16'd21516, 16'd6015, 16'd62181, 16'd44188, 16'd25641, 16'd37264, 16'd54544, 16'd31060, 16'd53738, 16'd60553, 16'd46084, 16'd43652, 16'd23504});
	test_expansion(128'hf77e7ae0fa84ff1bf8a95b4d9876b504, {16'd4405, 16'd64728, 16'd38692, 16'd51904, 16'd20133, 16'd38430, 16'd51664, 16'd8121, 16'd55270, 16'd64871, 16'd39775, 16'd6896, 16'd50364, 16'd57470, 16'd11610, 16'd27377, 16'd62035, 16'd26987, 16'd29821, 16'd706, 16'd22136, 16'd20119, 16'd18705, 16'd65186, 16'd1629, 16'd55151});
	test_expansion(128'h5ea6035b0d44619630facc8143176afb, {16'd129, 16'd54226, 16'd15927, 16'd41998, 16'd22625, 16'd2324, 16'd36853, 16'd4997, 16'd7171, 16'd64720, 16'd3416, 16'd14943, 16'd35481, 16'd46563, 16'd61223, 16'd51786, 16'd30935, 16'd22807, 16'd19115, 16'd35228, 16'd29169, 16'd26647, 16'd51232, 16'd14147, 16'd5915, 16'd56160});
	test_expansion(128'h57f1a233fd29ac03fd10f1f2f9419068, {16'd28488, 16'd46945, 16'd25292, 16'd55068, 16'd60222, 16'd27665, 16'd27333, 16'd22198, 16'd52767, 16'd24453, 16'd12043, 16'd14030, 16'd46202, 16'd49967, 16'd48825, 16'd29285, 16'd40668, 16'd3168, 16'd46720, 16'd16182, 16'd3557, 16'd38177, 16'd62915, 16'd24999, 16'd2529, 16'd14028});
	test_expansion(128'h0b2f44dffef3ce1cd10c10241f13dc62, {16'd32643, 16'd19269, 16'd43506, 16'd22177, 16'd47456, 16'd51184, 16'd9251, 16'd36241, 16'd47859, 16'd1469, 16'd54960, 16'd40831, 16'd1051, 16'd52810, 16'd55709, 16'd31981, 16'd43644, 16'd38428, 16'd63722, 16'd34960, 16'd37154, 16'd11466, 16'd26247, 16'd4793, 16'd50654, 16'd2752});
	test_expansion(128'hf0be852caa71a7c769d0f9db03a9b985, {16'd18999, 16'd22773, 16'd64928, 16'd17399, 16'd56950, 16'd40081, 16'd24839, 16'd17225, 16'd18021, 16'd38985, 16'd63571, 16'd27430, 16'd12693, 16'd29381, 16'd49846, 16'd65238, 16'd18690, 16'd53909, 16'd19516, 16'd58298, 16'd59401, 16'd9733, 16'd395, 16'd51911, 16'd53039, 16'd55201});
	test_expansion(128'ha17ad8f8f6576a714f3121f77c0886ac, {16'd21665, 16'd60312, 16'd45853, 16'd17729, 16'd61153, 16'd10412, 16'd33901, 16'd60914, 16'd2156, 16'd23993, 16'd22027, 16'd33454, 16'd38792, 16'd37559, 16'd10226, 16'd51116, 16'd15896, 16'd33347, 16'd8990, 16'd319, 16'd8357, 16'd63050, 16'd9633, 16'd3395, 16'd998, 16'd43159});
	test_expansion(128'he60dd2fc2823b86be3e6a8ca28cc586b, {16'd51494, 16'd39242, 16'd51243, 16'd50008, 16'd53037, 16'd28355, 16'd17674, 16'd17121, 16'd24917, 16'd61027, 16'd4893, 16'd2462, 16'd51758, 16'd34535, 16'd58464, 16'd1140, 16'd36337, 16'd63697, 16'd56100, 16'd61025, 16'd46617, 16'd29598, 16'd51917, 16'd37210, 16'd33972, 16'd40401});
	test_expansion(128'h4d5ff4fe3aff87f30de0a30de2cc8941, {16'd31456, 16'd38736, 16'd3867, 16'd20151, 16'd2052, 16'd388, 16'd54690, 16'd29089, 16'd31539, 16'd58240, 16'd41723, 16'd7350, 16'd22782, 16'd57005, 16'd13775, 16'd11041, 16'd15934, 16'd46499, 16'd52673, 16'd2127, 16'd6855, 16'd65411, 16'd13492, 16'd58499, 16'd7784, 16'd6935});
	test_expansion(128'h41339a45245229bf314dc27c2482ef26, {16'd19260, 16'd35731, 16'd39413, 16'd35134, 16'd36799, 16'd11759, 16'd56661, 16'd55718, 16'd43559, 16'd20658, 16'd24969, 16'd4845, 16'd46991, 16'd45309, 16'd31089, 16'd41162, 16'd65406, 16'd62870, 16'd10168, 16'd64993, 16'd17671, 16'd35715, 16'd5156, 16'd52422, 16'd18221, 16'd33277});
	test_expansion(128'h0bf9eed8d5ba50bb4fa5bfb004a03a63, {16'd37363, 16'd56541, 16'd26124, 16'd23954, 16'd28197, 16'd4623, 16'd22659, 16'd25693, 16'd27381, 16'd4392, 16'd5475, 16'd12210, 16'd3097, 16'd18874, 16'd29581, 16'd45525, 16'd34103, 16'd37213, 16'd29503, 16'd22797, 16'd26048, 16'd11695, 16'd23169, 16'd20874, 16'd43620, 16'd43832});
	test_expansion(128'h14ee8fd226192caad7336452e19b577c, {16'd21407, 16'd49620, 16'd2694, 16'd54636, 16'd52513, 16'd22190, 16'd37498, 16'd16621, 16'd49785, 16'd47331, 16'd61961, 16'd61758, 16'd33440, 16'd59908, 16'd63749, 16'd693, 16'd40144, 16'd43844, 16'd37078, 16'd40047, 16'd52239, 16'd32192, 16'd39010, 16'd25974, 16'd33644, 16'd27322});
	test_expansion(128'h116e50abaa6906f49254a9f0df585a0a, {16'd42634, 16'd27610, 16'd62368, 16'd38734, 16'd28621, 16'd31772, 16'd62738, 16'd12372, 16'd41143, 16'd3837, 16'd52519, 16'd42631, 16'd8214, 16'd23947, 16'd7889, 16'd51770, 16'd58744, 16'd41517, 16'd61277, 16'd6370, 16'd14842, 16'd60476, 16'd44158, 16'd30360, 16'd14386, 16'd64510});
	test_expansion(128'hc1824ab53e30d83b6bcd240755cf98ad, {16'd17825, 16'd55211, 16'd12790, 16'd30657, 16'd19280, 16'd27581, 16'd38856, 16'd6476, 16'd35144, 16'd59772, 16'd24670, 16'd44786, 16'd6363, 16'd34513, 16'd17751, 16'd30081, 16'd32871, 16'd38680, 16'd31411, 16'd46262, 16'd62116, 16'd35203, 16'd37467, 16'd12698, 16'd9436, 16'd24138});
	test_expansion(128'h797683f55ae457aad1446713f7d446fd, {16'd15880, 16'd21423, 16'd53158, 16'd57911, 16'd23850, 16'd22452, 16'd9101, 16'd31888, 16'd14574, 16'd24812, 16'd43132, 16'd49222, 16'd31749, 16'd36882, 16'd34348, 16'd30471, 16'd33994, 16'd448, 16'd51508, 16'd23049, 16'd21286, 16'd33319, 16'd2408, 16'd54427, 16'd24105, 16'd4599});
	test_expansion(128'heaa26b0ac90646f7598b0734b449a9a0, {16'd2706, 16'd5733, 16'd27291, 16'd12339, 16'd30537, 16'd39501, 16'd58879, 16'd27714, 16'd712, 16'd28193, 16'd6457, 16'd23793, 16'd3290, 16'd52240, 16'd14540, 16'd63575, 16'd51278, 16'd3136, 16'd51948, 16'd64744, 16'd19535, 16'd10468, 16'd26625, 16'd17960, 16'd7109, 16'd51166});
	test_expansion(128'h79e34dc0d8dec2da43872ff9407b82c2, {16'd6249, 16'd22031, 16'd41089, 16'd47380, 16'd45270, 16'd46065, 16'd15799, 16'd6469, 16'd61894, 16'd44633, 16'd5618, 16'd11792, 16'd25979, 16'd53126, 16'd8499, 16'd23642, 16'd51408, 16'd12771, 16'd40433, 16'd43803, 16'd40313, 16'd26833, 16'd18522, 16'd28952, 16'd37257, 16'd9068});
	test_expansion(128'haf1f4a659de341649752aee1bfb73a35, {16'd34906, 16'd9585, 16'd54965, 16'd25079, 16'd33727, 16'd23145, 16'd5098, 16'd46117, 16'd11107, 16'd2703, 16'd25739, 16'd32420, 16'd47859, 16'd38410, 16'd58318, 16'd34176, 16'd8334, 16'd30851, 16'd4469, 16'd19864, 16'd9082, 16'd39988, 16'd40733, 16'd10080, 16'd40741, 16'd29115});
	test_expansion(128'h1d5e34837369d7f557c1dc6645b2f0db, {16'd16690, 16'd30085, 16'd17856, 16'd56839, 16'd20932, 16'd21225, 16'd18015, 16'd57317, 16'd25992, 16'd29795, 16'd61875, 16'd48507, 16'd51246, 16'd22370, 16'd32538, 16'd30352, 16'd1576, 16'd57167, 16'd52579, 16'd8136, 16'd17554, 16'd32267, 16'd23169, 16'd49736, 16'd24233, 16'd11049});
	test_expansion(128'ha23d893b48d8ac48a7467ce1dcb5fb9b, {16'd56631, 16'd63098, 16'd41502, 16'd44369, 16'd21073, 16'd28080, 16'd44553, 16'd64401, 16'd47082, 16'd59421, 16'd29498, 16'd35519, 16'd26098, 16'd61964, 16'd4512, 16'd53814, 16'd31249, 16'd21797, 16'd46500, 16'd55562, 16'd54505, 16'd14696, 16'd13691, 16'd25766, 16'd47583, 16'd56082});
	test_expansion(128'he841d59bdafed87e5dfea6c204d91aad, {16'd33846, 16'd51587, 16'd44516, 16'd4556, 16'd51627, 16'd52519, 16'd18823, 16'd19767, 16'd12897, 16'd10529, 16'd63019, 16'd10129, 16'd35033, 16'd30606, 16'd7674, 16'd25582, 16'd13559, 16'd44100, 16'd45744, 16'd26391, 16'd14332, 16'd39373, 16'd59544, 16'd8204, 16'd53487, 16'd51267});
	test_expansion(128'h20dc8700f7245c3565d75e1a8ce50ecb, {16'd582, 16'd40056, 16'd50706, 16'd23113, 16'd37261, 16'd46109, 16'd50010, 16'd43110, 16'd35945, 16'd42169, 16'd16228, 16'd39592, 16'd36178, 16'd45077, 16'd2170, 16'd31671, 16'd7673, 16'd7628, 16'd36736, 16'd61508, 16'd46717, 16'd5656, 16'd34608, 16'd61267, 16'd37477, 16'd43574});
	test_expansion(128'hea75bcb471d9adfe4b4cbe0de1f8194e, {16'd55470, 16'd64854, 16'd54195, 16'd9284, 16'd13784, 16'd59840, 16'd25096, 16'd52699, 16'd849, 16'd13320, 16'd62779, 16'd15131, 16'd52027, 16'd62867, 16'd44263, 16'd55855, 16'd29891, 16'd10652, 16'd41748, 16'd49270, 16'd58971, 16'd61897, 16'd16641, 16'd16517, 16'd3712, 16'd36466});
	test_expansion(128'h7a9f6245ea1abd444c20e57eda992c63, {16'd43333, 16'd32708, 16'd38514, 16'd3066, 16'd42841, 16'd16412, 16'd59105, 16'd58935, 16'd48425, 16'd34396, 16'd42787, 16'd13790, 16'd28423, 16'd15447, 16'd64624, 16'd4056, 16'd59845, 16'd44157, 16'd9700, 16'd2986, 16'd37860, 16'd12361, 16'd24000, 16'd49451, 16'd37504, 16'd13457});
	test_expansion(128'h224f97ab6ff9b116810c41b283221106, {16'd40978, 16'd33763, 16'd48200, 16'd62652, 16'd51616, 16'd35212, 16'd41542, 16'd1859, 16'd50993, 16'd44674, 16'd19769, 16'd20758, 16'd30248, 16'd45748, 16'd604, 16'd41905, 16'd56610, 16'd51442, 16'd29714, 16'd21492, 16'd18785, 16'd13907, 16'd59688, 16'd34426, 16'd33162, 16'd12274});
	test_expansion(128'h5feb74b221cd592beeb8f13191ce3a44, {16'd36956, 16'd64651, 16'd23573, 16'd25522, 16'd24588, 16'd13518, 16'd36912, 16'd9956, 16'd15975, 16'd33979, 16'd17653, 16'd48036, 16'd22434, 16'd57205, 16'd25903, 16'd26760, 16'd38930, 16'd54159, 16'd17882, 16'd7888, 16'd36501, 16'd20111, 16'd51632, 16'd65234, 16'd49671, 16'd46298});
	test_expansion(128'h824aefa1bc07d62608ff57da9661ef35, {16'd45496, 16'd12697, 16'd45578, 16'd55822, 16'd57853, 16'd37130, 16'd45518, 16'd32554, 16'd16515, 16'd41230, 16'd26097, 16'd35378, 16'd5908, 16'd28216, 16'd19533, 16'd54625, 16'd18090, 16'd55392, 16'd12344, 16'd37938, 16'd7567, 16'd40762, 16'd59374, 16'd4401, 16'd18707, 16'd36857});
	test_expansion(128'h7c8702f5caa0146b75f27f6ef6ceffa7, {16'd26321, 16'd47213, 16'd38598, 16'd45665, 16'd24701, 16'd37471, 16'd61348, 16'd2213, 16'd56228, 16'd42619, 16'd47220, 16'd37686, 16'd11406, 16'd20941, 16'd50683, 16'd57759, 16'd18998, 16'd39474, 16'd29629, 16'd57408, 16'd59192, 16'd28746, 16'd37141, 16'd44634, 16'd8667, 16'd5824});
	test_expansion(128'haff6510855454f732da634fa1094b4b8, {16'd36749, 16'd18016, 16'd40777, 16'd36516, 16'd59856, 16'd25591, 16'd42436, 16'd2744, 16'd4396, 16'd35664, 16'd18534, 16'd2597, 16'd20357, 16'd44318, 16'd57283, 16'd16568, 16'd687, 16'd54473, 16'd17835, 16'd40433, 16'd1970, 16'd27101, 16'd41659, 16'd19482, 16'd12158, 16'd31977});
	test_expansion(128'h13a66e0f78d673c1c3a6225da4853273, {16'd53684, 16'd46806, 16'd1784, 16'd62502, 16'd3189, 16'd5970, 16'd28753, 16'd38292, 16'd19537, 16'd22417, 16'd57077, 16'd25966, 16'd45723, 16'd58881, 16'd58092, 16'd3878, 16'd3638, 16'd58321, 16'd36998, 16'd27926, 16'd65338, 16'd58796, 16'd63569, 16'd8334, 16'd11377, 16'd55477});
	test_expansion(128'h691909bf4f5f6b8ca0a456187d7d7d44, {16'd23533, 16'd25273, 16'd25255, 16'd9737, 16'd41048, 16'd48922, 16'd37712, 16'd40175, 16'd36835, 16'd50141, 16'd27597, 16'd15773, 16'd61407, 16'd25326, 16'd48277, 16'd62390, 16'd5493, 16'd12455, 16'd63071, 16'd59260, 16'd19874, 16'd31490, 16'd56450, 16'd11405, 16'd18693, 16'd27892});
	test_expansion(128'h40a6e56f1079f035cea87b4edd33475b, {16'd59469, 16'd7080, 16'd45335, 16'd10340, 16'd19311, 16'd56509, 16'd21357, 16'd12517, 16'd4395, 16'd61785, 16'd29000, 16'd24068, 16'd23432, 16'd40241, 16'd34810, 16'd30311, 16'd14965, 16'd39771, 16'd49834, 16'd60075, 16'd22967, 16'd29718, 16'd54298, 16'd45919, 16'd56681, 16'd29604});
	test_expansion(128'hbabd4eb62e9f25de992ea4ed9e773c6e, {16'd25539, 16'd26650, 16'd57219, 16'd62238, 16'd36317, 16'd63136, 16'd43881, 16'd16994, 16'd614, 16'd33323, 16'd39429, 16'd17915, 16'd12564, 16'd31393, 16'd48641, 16'd32113, 16'd7152, 16'd34212, 16'd60607, 16'd52029, 16'd41794, 16'd34920, 16'd26559, 16'd56131, 16'd16880, 16'd9446});
	test_expansion(128'hc28ac7326489ea65bb1f80a18ae563a2, {16'd42608, 16'd53162, 16'd5024, 16'd43426, 16'd62232, 16'd33299, 16'd50476, 16'd8890, 16'd28477, 16'd19528, 16'd3526, 16'd64709, 16'd39803, 16'd14078, 16'd7036, 16'd34391, 16'd31876, 16'd31004, 16'd56804, 16'd36628, 16'd930, 16'd44842, 16'd133, 16'd24168, 16'd59617, 16'd922});
	test_expansion(128'h3f1488d385eb18cc10de000daf3c8662, {16'd60000, 16'd55211, 16'd37567, 16'd36647, 16'd13077, 16'd42940, 16'd20044, 16'd31789, 16'd29906, 16'd1589, 16'd3941, 16'd46126, 16'd14483, 16'd57967, 16'd54337, 16'd52577, 16'd40140, 16'd40702, 16'd27341, 16'd63478, 16'd35800, 16'd32330, 16'd9032, 16'd20239, 16'd12527, 16'd28925});
	test_expansion(128'h51c086383f19004b285ce1e2b4d6f4cc, {16'd18047, 16'd33167, 16'd53535, 16'd49341, 16'd36528, 16'd19718, 16'd38378, 16'd52617, 16'd34655, 16'd48570, 16'd36980, 16'd64444, 16'd5373, 16'd40272, 16'd26560, 16'd41789, 16'd49106, 16'd51063, 16'd22000, 16'd12036, 16'd39341, 16'd58644, 16'd13685, 16'd52769, 16'd63251, 16'd64719});
	test_expansion(128'h807944f6a6255cb3101bef2d1db8f403, {16'd50791, 16'd64073, 16'd1250, 16'd39841, 16'd20441, 16'd24803, 16'd64590, 16'd18014, 16'd10282, 16'd7965, 16'd1365, 16'd64076, 16'd59410, 16'd61019, 16'd32761, 16'd42019, 16'd50921, 16'd19508, 16'd9994, 16'd27726, 16'd8417, 16'd5572, 16'd33048, 16'd60782, 16'd36223, 16'd25473});
	test_expansion(128'h973942cfc2cfcb7c4bf771ecf7c03653, {16'd11033, 16'd64552, 16'd26627, 16'd18763, 16'd57602, 16'd40177, 16'd34998, 16'd11482, 16'd32880, 16'd53319, 16'd40576, 16'd56086, 16'd43616, 16'd18515, 16'd22688, 16'd5063, 16'd44731, 16'd2608, 16'd40362, 16'd42601, 16'd17390, 16'd6204, 16'd5253, 16'd29171, 16'd18970, 16'd43092});
	test_expansion(128'h61b9c971cdd99c987c1a7e72d7f6cc70, {16'd63540, 16'd8794, 16'd22117, 16'd29695, 16'd9092, 16'd41491, 16'd4166, 16'd62752, 16'd1956, 16'd49978, 16'd15360, 16'd12743, 16'd48501, 16'd47107, 16'd27061, 16'd63534, 16'd56154, 16'd32368, 16'd53410, 16'd8411, 16'd7400, 16'd54684, 16'd46530, 16'd40695, 16'd6703, 16'd36415});
	test_expansion(128'hd13311f83219b2e07ca907d2e958c67d, {16'd4707, 16'd23417, 16'd7833, 16'd37836, 16'd25834, 16'd56858, 16'd10086, 16'd15667, 16'd41518, 16'd55306, 16'd37609, 16'd248, 16'd10344, 16'd30297, 16'd9959, 16'd61308, 16'd50460, 16'd34825, 16'd22460, 16'd51824, 16'd37293, 16'd41276, 16'd17737, 16'd56186, 16'd9847, 16'd25930});
	test_expansion(128'h06c1bee88eff0d403eed140275bee580, {16'd42925, 16'd18106, 16'd61378, 16'd59140, 16'd7066, 16'd34318, 16'd38670, 16'd36817, 16'd9148, 16'd23633, 16'd60498, 16'd11993, 16'd63396, 16'd12782, 16'd44216, 16'd56197, 16'd9014, 16'd24778, 16'd48848, 16'd44865, 16'd27162, 16'd50806, 16'd1610, 16'd30938, 16'd57172, 16'd13597});
	test_expansion(128'he0e474e2806a8d848bd0083cfe7d6def, {16'd59739, 16'd56699, 16'd2221, 16'd42073, 16'd49639, 16'd41195, 16'd55552, 16'd18158, 16'd48610, 16'd57637, 16'd4544, 16'd15264, 16'd20454, 16'd37998, 16'd50958, 16'd58, 16'd4948, 16'd44105, 16'd44830, 16'd14099, 16'd1359, 16'd28578, 16'd39624, 16'd59338, 16'd44389, 16'd26559});
	test_expansion(128'hc2572a0fc974fa8df504983f173c73db, {16'd17282, 16'd57997, 16'd10115, 16'd41981, 16'd20625, 16'd54815, 16'd52961, 16'd15273, 16'd34462, 16'd62328, 16'd32528, 16'd61391, 16'd56009, 16'd36856, 16'd23324, 16'd2022, 16'd1174, 16'd39353, 16'd16113, 16'd6003, 16'd57432, 16'd55438, 16'd23046, 16'd12447, 16'd44588, 16'd42661});
	test_expansion(128'h408c8c900c1ea043c93253a26e9576c3, {16'd26195, 16'd50056, 16'd47250, 16'd20017, 16'd45122, 16'd53476, 16'd9986, 16'd38499, 16'd9881, 16'd32316, 16'd7068, 16'd19542, 16'd37487, 16'd47893, 16'd19928, 16'd17138, 16'd34093, 16'd18153, 16'd20389, 16'd34004, 16'd46136, 16'd26285, 16'd34511, 16'd34411, 16'd60011, 16'd5183});
	test_expansion(128'h29b7f9c6bccaf35bd6847ca802c8bc41, {16'd52242, 16'd61137, 16'd12953, 16'd5234, 16'd11166, 16'd38401, 16'd39576, 16'd23909, 16'd11737, 16'd4427, 16'd50808, 16'd39707, 16'd12264, 16'd15721, 16'd19104, 16'd31612, 16'd42433, 16'd52989, 16'd34797, 16'd46992, 16'd20617, 16'd36320, 16'd59759, 16'd32564, 16'd32323, 16'd41652});
	test_expansion(128'h8ed3bea9ad07671829dccf4cf0b33043, {16'd23032, 16'd64715, 16'd47210, 16'd4010, 16'd12044, 16'd16345, 16'd29777, 16'd56569, 16'd1376, 16'd39995, 16'd35985, 16'd9006, 16'd20394, 16'd9122, 16'd43346, 16'd65364, 16'd44981, 16'd63025, 16'd19510, 16'd5523, 16'd29125, 16'd13945, 16'd37865, 16'd59382, 16'd44620, 16'd21114});
	test_expansion(128'h4a19f26f9cfde6fdda0f8a756483dc5f, {16'd4090, 16'd54755, 16'd24476, 16'd35577, 16'd40198, 16'd31738, 16'd47741, 16'd33546, 16'd13299, 16'd52605, 16'd54877, 16'd64000, 16'd42089, 16'd55102, 16'd21315, 16'd33332, 16'd25952, 16'd15150, 16'd61419, 16'd63054, 16'd53505, 16'd35764, 16'd22607, 16'd40848, 16'd8556, 16'd52725});
	test_expansion(128'hb054e87ced4f5bc88bd9d803d753687b, {16'd3270, 16'd33864, 16'd730, 16'd43892, 16'd27552, 16'd40470, 16'd59848, 16'd33644, 16'd61079, 16'd61704, 16'd7263, 16'd31315, 16'd25228, 16'd9789, 16'd43220, 16'd4890, 16'd43497, 16'd48918, 16'd38065, 16'd47409, 16'd51146, 16'd13935, 16'd1694, 16'd16201, 16'd59520, 16'd20117});
	test_expansion(128'h4c517cfdd4391db31bf738f6550b3caa, {16'd35937, 16'd31676, 16'd58857, 16'd61304, 16'd56383, 16'd23032, 16'd42132, 16'd47241, 16'd18437, 16'd55080, 16'd22644, 16'd35068, 16'd10751, 16'd53007, 16'd54742, 16'd41709, 16'd22473, 16'd8697, 16'd22100, 16'd23626, 16'd25665, 16'd62326, 16'd17743, 16'd26933, 16'd10583, 16'd29121});
	test_expansion(128'h1e88ee9150662b8e7e1c556bcfff09d9, {16'd31526, 16'd51215, 16'd47995, 16'd54792, 16'd12262, 16'd65386, 16'd2875, 16'd4536, 16'd53271, 16'd3696, 16'd40003, 16'd2143, 16'd40251, 16'd48025, 16'd46397, 16'd27654, 16'd37974, 16'd8965, 16'd13812, 16'd27410, 16'd16083, 16'd19966, 16'd65507, 16'd49806, 16'd49648, 16'd20453});
	test_expansion(128'hccf37acd483017884c1a5c5574dc6a95, {16'd7496, 16'd18189, 16'd54009, 16'd16854, 16'd62328, 16'd23799, 16'd41564, 16'd30621, 16'd24307, 16'd25379, 16'd23637, 16'd39768, 16'd40399, 16'd59702, 16'd62911, 16'd20230, 16'd15414, 16'd55547, 16'd22732, 16'd21414, 16'd46152, 16'd52890, 16'd37090, 16'd38096, 16'd29517, 16'd57012});
	test_expansion(128'h318bdf69554529ef3acfe1a0a40ba734, {16'd9334, 16'd19755, 16'd1343, 16'd2718, 16'd11083, 16'd14664, 16'd64433, 16'd5640, 16'd12577, 16'd1942, 16'd12414, 16'd12729, 16'd13309, 16'd18324, 16'd61450, 16'd46535, 16'd36998, 16'd52428, 16'd4702, 16'd2877, 16'd9435, 16'd24429, 16'd26615, 16'd1382, 16'd33416, 16'd6920});
	test_expansion(128'hce0aa181e902bf4e2f562845cb976d6f, {16'd16241, 16'd31224, 16'd18037, 16'd3038, 16'd11760, 16'd43154, 16'd47101, 16'd50808, 16'd17, 16'd4734, 16'd26918, 16'd54384, 16'd21454, 16'd27657, 16'd59868, 16'd57258, 16'd33021, 16'd45195, 16'd18120, 16'd7854, 16'd19316, 16'd5648, 16'd630, 16'd41787, 16'd28522, 16'd49942});
	test_expansion(128'hdc2021cbe377c3ecaec0b6aa912b7be3, {16'd36848, 16'd1522, 16'd44879, 16'd41666, 16'd56004, 16'd1613, 16'd41937, 16'd57849, 16'd25278, 16'd56417, 16'd44336, 16'd28639, 16'd3495, 16'd30385, 16'd56919, 16'd21204, 16'd45105, 16'd3893, 16'd52498, 16'd31953, 16'd30294, 16'd14636, 16'd24916, 16'd28356, 16'd40347, 16'd60288});
	test_expansion(128'hbb522f5263eb1056b66539431141c545, {16'd1406, 16'd11096, 16'd62623, 16'd33752, 16'd52135, 16'd49756, 16'd23330, 16'd32362, 16'd29519, 16'd21281, 16'd4492, 16'd46471, 16'd48118, 16'd30607, 16'd39535, 16'd27806, 16'd244, 16'd48207, 16'd4529, 16'd45447, 16'd7634, 16'd13421, 16'd39214, 16'd21509, 16'd15388, 16'd58669});
	test_expansion(128'h633aa0d0644f8fcbf005f362fbeaff37, {16'd52398, 16'd24917, 16'd57531, 16'd61848, 16'd36545, 16'd43771, 16'd64992, 16'd21820, 16'd2536, 16'd7333, 16'd61547, 16'd41675, 16'd58508, 16'd43958, 16'd2658, 16'd23662, 16'd9504, 16'd41941, 16'd24095, 16'd22920, 16'd58254, 16'd2155, 16'd8415, 16'd40282, 16'd21646, 16'd58714});
	test_expansion(128'h9e318bcff51c29d76b5dc05ebbafa9e1, {16'd21224, 16'd40916, 16'd60052, 16'd55098, 16'd3882, 16'd44078, 16'd29016, 16'd9283, 16'd14401, 16'd37910, 16'd31133, 16'd1583, 16'd63314, 16'd39442, 16'd52691, 16'd58735, 16'd34285, 16'd47715, 16'd9714, 16'd60801, 16'd41338, 16'd43422, 16'd450, 16'd17367, 16'd58244, 16'd11623});
	test_expansion(128'h23d2ece3eefeddcd2be7124526cf4e24, {16'd128, 16'd63598, 16'd2999, 16'd40288, 16'd36296, 16'd29055, 16'd56957, 16'd21632, 16'd64548, 16'd27989, 16'd47075, 16'd48503, 16'd13842, 16'd47053, 16'd37795, 16'd60758, 16'd20718, 16'd9393, 16'd9380, 16'd1540, 16'd15352, 16'd12435, 16'd17739, 16'd24059, 16'd26281, 16'd59618});
	test_expansion(128'hd5ec6aa05f75874ae5a1a361f84eea93, {16'd52298, 16'd30354, 16'd22991, 16'd21589, 16'd34837, 16'd40138, 16'd21793, 16'd61349, 16'd41758, 16'd3156, 16'd5643, 16'd55812, 16'd62353, 16'd51541, 16'd12973, 16'd20921, 16'd49627, 16'd18152, 16'd55347, 16'd18796, 16'd23305, 16'd6526, 16'd30908, 16'd22921, 16'd5391, 16'd58237});
	test_expansion(128'h2c9b941b2af7b608898362820c4d3325, {16'd22437, 16'd3526, 16'd62229, 16'd59378, 16'd2094, 16'd19427, 16'd14130, 16'd20588, 16'd61878, 16'd11667, 16'd48531, 16'd62724, 16'd31579, 16'd50755, 16'd571, 16'd26113, 16'd55793, 16'd47962, 16'd9540, 16'd41141, 16'd59972, 16'd62368, 16'd58817, 16'd56142, 16'd38385, 16'd60588});
	test_expansion(128'hc4f4b05dd2104ae9fd5f48dc7e134c12, {16'd62853, 16'd44303, 16'd37165, 16'd4262, 16'd43865, 16'd49225, 16'd9407, 16'd18300, 16'd31234, 16'd16779, 16'd32576, 16'd52004, 16'd2976, 16'd65298, 16'd39582, 16'd46065, 16'd4565, 16'd36078, 16'd18981, 16'd38272, 16'd62270, 16'd3192, 16'd14746, 16'd53133, 16'd46028, 16'd9197});
	test_expansion(128'hd8ee86751bd1af50f7dc0d5dafe3b290, {16'd5107, 16'd31293, 16'd62254, 16'd31799, 16'd63357, 16'd34159, 16'd37177, 16'd33473, 16'd26247, 16'd28271, 16'd5364, 16'd55515, 16'd20832, 16'd34609, 16'd22231, 16'd34573, 16'd56317, 16'd53474, 16'd8924, 16'd65036, 16'd32244, 16'd24731, 16'd14506, 16'd13976, 16'd33323, 16'd5312});
	test_expansion(128'h8643213558108da08a6992b10fd3a64f, {16'd22432, 16'd42744, 16'd35218, 16'd22676, 16'd31734, 16'd47131, 16'd21151, 16'd19217, 16'd56562, 16'd161, 16'd48120, 16'd17804, 16'd40370, 16'd37862, 16'd56929, 16'd9220, 16'd21630, 16'd1674, 16'd18195, 16'd15464, 16'd34716, 16'd54825, 16'd35028, 16'd45471, 16'd64710, 16'd59791});
	test_expansion(128'h50b75fb0fc3932876e5b9cc92168ba4d, {16'd4024, 16'd14177, 16'd16806, 16'd64784, 16'd24084, 16'd32053, 16'd29649, 16'd4251, 16'd25945, 16'd8945, 16'd28152, 16'd15044, 16'd2696, 16'd12622, 16'd39709, 16'd12942, 16'd50041, 16'd33960, 16'd42702, 16'd62424, 16'd35125, 16'd49095, 16'd12293, 16'd3353, 16'd20384, 16'd41745});
	test_expansion(128'h527e795e4a70fb482309c9ceb84c470e, {16'd20226, 16'd3819, 16'd20070, 16'd42388, 16'd9062, 16'd47405, 16'd1955, 16'd25198, 16'd5911, 16'd1678, 16'd46951, 16'd65015, 16'd57060, 16'd3036, 16'd26950, 16'd33892, 16'd15281, 16'd4550, 16'd55279, 16'd60586, 16'd41492, 16'd18956, 16'd8276, 16'd63072, 16'd61889, 16'd62603});
	test_expansion(128'h28dd6b35c15febda25ecd01291c6bf90, {16'd3588, 16'd38957, 16'd56115, 16'd25712, 16'd37466, 16'd5683, 16'd11603, 16'd10542, 16'd33995, 16'd38995, 16'd57061, 16'd13090, 16'd25368, 16'd26741, 16'd62542, 16'd46895, 16'd40065, 16'd62592, 16'd60903, 16'd24549, 16'd3944, 16'd15533, 16'd5639, 16'd63636, 16'd44019, 16'd16360});
	test_expansion(128'h78a32eea8f2ddbcdc584830fb1e41006, {16'd62838, 16'd41998, 16'd361, 16'd11195, 16'd44710, 16'd62770, 16'd28569, 16'd28823, 16'd22079, 16'd32116, 16'd20899, 16'd58140, 16'd44741, 16'd31596, 16'd1537, 16'd12745, 16'd50080, 16'd28419, 16'd45566, 16'd50967, 16'd64101, 16'd34261, 16'd16279, 16'd60966, 16'd30471, 16'd15149});
	test_expansion(128'h5866e39d4033ac5db1cd6acf87e0164a, {16'd51741, 16'd51867, 16'd61844, 16'd11581, 16'd37736, 16'd64604, 16'd1054, 16'd55460, 16'd29606, 16'd5097, 16'd7861, 16'd13423, 16'd35015, 16'd8326, 16'd41537, 16'd22271, 16'd9471, 16'd40735, 16'd27847, 16'd36344, 16'd8464, 16'd55569, 16'd7131, 16'd20564, 16'd22404, 16'd12867});
	test_expansion(128'h52a761cc65d28cd19575058ad377d496, {16'd27683, 16'd35522, 16'd2865, 16'd64939, 16'd28315, 16'd35948, 16'd56771, 16'd10900, 16'd14734, 16'd13025, 16'd16628, 16'd21576, 16'd12627, 16'd12533, 16'd27371, 16'd4868, 16'd53601, 16'd55592, 16'd44438, 16'd57293, 16'd25239, 16'd51196, 16'd7035, 16'd9089, 16'd19843, 16'd3274});
	test_expansion(128'h5bc8960c810bba675800553a5ba72fb3, {16'd21607, 16'd44166, 16'd62735, 16'd24264, 16'd26231, 16'd20691, 16'd14312, 16'd8278, 16'd17389, 16'd4657, 16'd20798, 16'd22201, 16'd51107, 16'd44883, 16'd4587, 16'd58308, 16'd39025, 16'd12681, 16'd36405, 16'd8171, 16'd17786, 16'd47948, 16'd23067, 16'd55726, 16'd45944, 16'd59249});
	test_expansion(128'h5dd1c08fb011677fd5fb5077e8273493, {16'd52989, 16'd26208, 16'd37595, 16'd47505, 16'd18610, 16'd2070, 16'd23813, 16'd44872, 16'd62675, 16'd44008, 16'd25695, 16'd24964, 16'd31255, 16'd38031, 16'd51105, 16'd29530, 16'd18124, 16'd60180, 16'd21517, 16'd47817, 16'd38192, 16'd40771, 16'd10637, 16'd9215, 16'd46518, 16'd8757});
	test_expansion(128'h7ce10ae45ab2c16c02f24bed3a0f0d38, {16'd19789, 16'd15261, 16'd52612, 16'd23986, 16'd63909, 16'd43164, 16'd21766, 16'd39076, 16'd23287, 16'd60526, 16'd42655, 16'd20248, 16'd59761, 16'd26339, 16'd29843, 16'd40401, 16'd32301, 16'd31204, 16'd1733, 16'd23379, 16'd32297, 16'd18926, 16'd13174, 16'd62539, 16'd34704, 16'd19702});
	test_expansion(128'h9c1c17214e0834ac7e23001179b72cae, {16'd15198, 16'd5995, 16'd60880, 16'd25278, 16'd9568, 16'd27702, 16'd18391, 16'd3147, 16'd6755, 16'd2011, 16'd18482, 16'd49565, 16'd48643, 16'd61694, 16'd51562, 16'd43752, 16'd40230, 16'd40549, 16'd9950, 16'd31702, 16'd40995, 16'd41182, 16'd40470, 16'd52920, 16'd24442, 16'd15838});
	test_expansion(128'hf5a26325a5d5aca0c5b46008af5d34f2, {16'd59329, 16'd2384, 16'd9979, 16'd57001, 16'd47577, 16'd5826, 16'd40413, 16'd55879, 16'd25126, 16'd48472, 16'd41818, 16'd40229, 16'd32242, 16'd25400, 16'd197, 16'd58425, 16'd50094, 16'd49583, 16'd48032, 16'd41158, 16'd54171, 16'd55263, 16'd59678, 16'd12986, 16'd44506, 16'd30110});
	test_expansion(128'hd144dcd0a83fbbf1adb010fdb737b26e, {16'd24628, 16'd30857, 16'd9655, 16'd60384, 16'd38371, 16'd43234, 16'd19199, 16'd2232, 16'd30923, 16'd19823, 16'd43777, 16'd63213, 16'd34693, 16'd30266, 16'd46133, 16'd47963, 16'd37233, 16'd2261, 16'd57380, 16'd691, 16'd44877, 16'd51610, 16'd60320, 16'd51874, 16'd53384, 16'd60016});
	test_expansion(128'h3fbc48008da8557c0423b8f80cd9a0af, {16'd30931, 16'd54114, 16'd59456, 16'd5308, 16'd59402, 16'd43950, 16'd25542, 16'd53022, 16'd755, 16'd39220, 16'd43153, 16'd41902, 16'd16524, 16'd22636, 16'd28423, 16'd730, 16'd27747, 16'd3837, 16'd38741, 16'd61494, 16'd51296, 16'd7754, 16'd18839, 16'd51996, 16'd10024, 16'd33734});
	test_expansion(128'h5497c931e372f3007e36878f581e150f, {16'd47328, 16'd3466, 16'd49760, 16'd56108, 16'd17921, 16'd6114, 16'd39952, 16'd22332, 16'd59866, 16'd3122, 16'd46697, 16'd25292, 16'd39722, 16'd27255, 16'd7820, 16'd28492, 16'd24016, 16'd48390, 16'd28308, 16'd50617, 16'd12865, 16'd25227, 16'd38108, 16'd5140, 16'd53511, 16'd11896});
	test_expansion(128'hd57989926a262b4d50731f8b08a5de4f, {16'd10909, 16'd11195, 16'd50317, 16'd52373, 16'd26861, 16'd61848, 16'd40215, 16'd23355, 16'd14721, 16'd65183, 16'd51008, 16'd44576, 16'd63436, 16'd32044, 16'd2458, 16'd59514, 16'd34040, 16'd48046, 16'd2511, 16'd35573, 16'd34040, 16'd2577, 16'd53340, 16'd5838, 16'd20103, 16'd2562});
	test_expansion(128'h04b6f44bddd5a60943b94e5a314c8606, {16'd35892, 16'd62770, 16'd56989, 16'd31696, 16'd52567, 16'd12021, 16'd24603, 16'd32106, 16'd46625, 16'd60433, 16'd74, 16'd6236, 16'd60124, 16'd52282, 16'd16865, 16'd17238, 16'd41174, 16'd51396, 16'd49208, 16'd6718, 16'd17932, 16'd15363, 16'd38869, 16'd979, 16'd27820, 16'd46964});
	test_expansion(128'h51861b9fc05e9fa5590508dafddf91fb, {16'd59968, 16'd45813, 16'd24185, 16'd28464, 16'd39864, 16'd29788, 16'd2324, 16'd34718, 16'd55327, 16'd48336, 16'd3380, 16'd20413, 16'd14460, 16'd26646, 16'd10466, 16'd37291, 16'd40087, 16'd56547, 16'd24831, 16'd58130, 16'd34698, 16'd24300, 16'd6121, 16'd15443, 16'd11333, 16'd20494});
	test_expansion(128'h40991b00936b4b3fded1d9a88dfd3554, {16'd60149, 16'd20766, 16'd27165, 16'd11684, 16'd9548, 16'd37575, 16'd8511, 16'd62422, 16'd40694, 16'd44119, 16'd13347, 16'd62209, 16'd7345, 16'd16965, 16'd49983, 16'd480, 16'd28818, 16'd47057, 16'd18791, 16'd58662, 16'd51059, 16'd28013, 16'd12309, 16'd51562, 16'd63188, 16'd33033});
	test_expansion(128'hf9fbbc666063c2a42615a99c0a7901ff, {16'd60686, 16'd29325, 16'd23559, 16'd57043, 16'd14143, 16'd18339, 16'd33804, 16'd31932, 16'd46361, 16'd1044, 16'd12659, 16'd27772, 16'd53198, 16'd57556, 16'd50306, 16'd15723, 16'd27562, 16'd60972, 16'd23975, 16'd63475, 16'd49113, 16'd60489, 16'd10912, 16'd49410, 16'd63110, 16'd5221});
	test_expansion(128'hc429e25121925039143e8eb3501aa680, {16'd41177, 16'd43914, 16'd11194, 16'd55599, 16'd52531, 16'd22695, 16'd32410, 16'd14674, 16'd30213, 16'd48012, 16'd63019, 16'd4532, 16'd5777, 16'd48238, 16'd31214, 16'd59526, 16'd11044, 16'd58419, 16'd10603, 16'd17655, 16'd47838, 16'd31300, 16'd32921, 16'd44829, 16'd9731, 16'd23490});
	test_expansion(128'h8a01705b3eaad4f1e947e9bdea579f75, {16'd34408, 16'd37161, 16'd8564, 16'd19926, 16'd21731, 16'd64055, 16'd22753, 16'd27953, 16'd2497, 16'd946, 16'd7922, 16'd47532, 16'd11390, 16'd9532, 16'd11591, 16'd13476, 16'd49410, 16'd40847, 16'd51356, 16'd27173, 16'd50179, 16'd45952, 16'd57481, 16'd30796, 16'd10824, 16'd63178});
	test_expansion(128'hb13ce6dc8268ae9950a003a83e9d960b, {16'd57177, 16'd32376, 16'd44156, 16'd51102, 16'd25693, 16'd36704, 16'd6109, 16'd36136, 16'd26607, 16'd21170, 16'd30530, 16'd53068, 16'd24305, 16'd50213, 16'd10859, 16'd4512, 16'd11323, 16'd21067, 16'd23078, 16'd1276, 16'd58044, 16'd61165, 16'd784, 16'd44608, 16'd62456, 16'd60773});
	test_expansion(128'h18a3bf15bd65ede0ab86997a851a7a20, {16'd26552, 16'd64007, 16'd9655, 16'd44095, 16'd26631, 16'd23480, 16'd6287, 16'd13882, 16'd31697, 16'd44318, 16'd60825, 16'd13969, 16'd37019, 16'd36656, 16'd28849, 16'd41710, 16'd10121, 16'd57919, 16'd1457, 16'd19755, 16'd28540, 16'd38373, 16'd33821, 16'd7339, 16'd41559, 16'd28875});
	test_expansion(128'h9969f90414583680fd34f3c364304650, {16'd42519, 16'd7129, 16'd14124, 16'd41346, 16'd5101, 16'd54180, 16'd27855, 16'd48330, 16'd56402, 16'd12102, 16'd36681, 16'd37210, 16'd3879, 16'd3519, 16'd65133, 16'd3609, 16'd55237, 16'd64863, 16'd34662, 16'd49315, 16'd40267, 16'd44336, 16'd46505, 16'd58088, 16'd55121, 16'd4204});
	test_expansion(128'hb396b5c4a036fb77117058525069d6c3, {16'd20968, 16'd63310, 16'd32766, 16'd45617, 16'd8336, 16'd36896, 16'd46633, 16'd47539, 16'd17967, 16'd22928, 16'd44016, 16'd52462, 16'd55311, 16'd28259, 16'd61240, 16'd21363, 16'd21762, 16'd54641, 16'd40524, 16'd37655, 16'd59282, 16'd28363, 16'd517, 16'd64200, 16'd60278, 16'd4466});
	test_expansion(128'he1e56e10f669b4c53741a11f86b5d4b8, {16'd42653, 16'd52977, 16'd24413, 16'd58695, 16'd44278, 16'd12519, 16'd33553, 16'd51382, 16'd58730, 16'd16420, 16'd32101, 16'd58475, 16'd26384, 16'd10342, 16'd56623, 16'd43405, 16'd46949, 16'd26950, 16'd60615, 16'd47415, 16'd55820, 16'd1351, 16'd35573, 16'd47994, 16'd4605, 16'd30468});
	test_expansion(128'h4a992b276104ea760711fec31670a322, {16'd12248, 16'd29733, 16'd57116, 16'd65405, 16'd41612, 16'd57458, 16'd14786, 16'd46406, 16'd61433, 16'd54251, 16'd46301, 16'd55657, 16'd12509, 16'd47066, 16'd38594, 16'd27834, 16'd36398, 16'd38036, 16'd5197, 16'd38312, 16'd46995, 16'd10251, 16'd23607, 16'd1259, 16'd11279, 16'd29799});
	test_expansion(128'h5e7fa40dd0763d23b33c596982626a10, {16'd12345, 16'd46358, 16'd6180, 16'd47348, 16'd54963, 16'd14058, 16'd62633, 16'd37909, 16'd13474, 16'd48994, 16'd33533, 16'd33860, 16'd33725, 16'd14908, 16'd51156, 16'd118, 16'd10547, 16'd62350, 16'd45757, 16'd37333, 16'd6678, 16'd20656, 16'd48178, 16'd616, 16'd38573, 16'd60457});
	test_expansion(128'hba00fb93e78ca464538bd9662b095d7b, {16'd39100, 16'd18004, 16'd7193, 16'd49420, 16'd23224, 16'd63135, 16'd26576, 16'd62625, 16'd38158, 16'd57132, 16'd52005, 16'd46497, 16'd56739, 16'd33344, 16'd39520, 16'd1046, 16'd64420, 16'd11404, 16'd29414, 16'd22256, 16'd42073, 16'd49892, 16'd52602, 16'd12059, 16'd49291, 16'd45680});
	test_expansion(128'he0c42ecd0e102bbe63210beddd29d64f, {16'd14375, 16'd47179, 16'd42367, 16'd43024, 16'd54873, 16'd10743, 16'd18014, 16'd9736, 16'd63405, 16'd21958, 16'd58114, 16'd59208, 16'd39854, 16'd58988, 16'd33216, 16'd12374, 16'd46744, 16'd46533, 16'd39103, 16'd48446, 16'd9742, 16'd14724, 16'd32381, 16'd23003, 16'd17876, 16'd49266});
	test_expansion(128'hc4ec5d8374de0b45a65685069c644993, {16'd33206, 16'd29619, 16'd30293, 16'd6667, 16'd55817, 16'd58780, 16'd22673, 16'd26319, 16'd37997, 16'd61228, 16'd39112, 16'd35784, 16'd8814, 16'd59355, 16'd30638, 16'd62786, 16'd19198, 16'd48789, 16'd4156, 16'd2210, 16'd27304, 16'd4606, 16'd63753, 16'd18177, 16'd45348, 16'd55189});
	test_expansion(128'hb839a61a819750322b598fa2b6ee3d44, {16'd57852, 16'd49290, 16'd41502, 16'd12964, 16'd11634, 16'd20509, 16'd51862, 16'd64145, 16'd49223, 16'd51842, 16'd45831, 16'd18781, 16'd20968, 16'd38990, 16'd53565, 16'd28222, 16'd53019, 16'd63797, 16'd8078, 16'd1810, 16'd19726, 16'd33735, 16'd17635, 16'd9017, 16'd48035, 16'd29879});
	test_expansion(128'hf569eb0908e61899f9f151c8f490321b, {16'd36233, 16'd43544, 16'd43879, 16'd28420, 16'd10807, 16'd63289, 16'd8027, 16'd27554, 16'd35402, 16'd48642, 16'd47513, 16'd45150, 16'd14851, 16'd6320, 16'd40347, 16'd55428, 16'd17286, 16'd50081, 16'd39430, 16'd35614, 16'd44500, 16'd16425, 16'd8509, 16'd38958, 16'd42567, 16'd57829});
	test_expansion(128'h1051449b152dd77a8f74a7ca4b1a4d8b, {16'd3061, 16'd6418, 16'd48300, 16'd4542, 16'd13083, 16'd32132, 16'd57484, 16'd31703, 16'd34229, 16'd20639, 16'd12312, 16'd45386, 16'd48635, 16'd13962, 16'd47429, 16'd30928, 16'd49144, 16'd65347, 16'd50382, 16'd9726, 16'd40871, 16'd43824, 16'd22914, 16'd27455, 16'd35981, 16'd15569});
	test_expansion(128'h15903b59529c5c6d76e4aaa4d2409c28, {16'd37826, 16'd49458, 16'd29134, 16'd44984, 16'd4189, 16'd52143, 16'd46834, 16'd37804, 16'd6511, 16'd57760, 16'd63407, 16'd61437, 16'd55139, 16'd59841, 16'd51242, 16'd19497, 16'd52546, 16'd28179, 16'd3574, 16'd18331, 16'd28298, 16'd27361, 16'd5967, 16'd19770, 16'd56514, 16'd13999});
	test_expansion(128'h199d6b84d2787fa955df3d86c4d48a3c, {16'd37432, 16'd22912, 16'd40197, 16'd5209, 16'd3366, 16'd46048, 16'd3954, 16'd5766, 16'd8435, 16'd8254, 16'd42499, 16'd9969, 16'd21983, 16'd59984, 16'd52977, 16'd17248, 16'd1568, 16'd54192, 16'd28229, 16'd42476, 16'd62234, 16'd25137, 16'd1505, 16'd62934, 16'd40158, 16'd54370});
	test_expansion(128'h2d875fade6e92ab194f820ebdfebf466, {16'd23888, 16'd60653, 16'd1986, 16'd3352, 16'd30846, 16'd21108, 16'd10034, 16'd61315, 16'd45545, 16'd55249, 16'd41926, 16'd35996, 16'd23678, 16'd23522, 16'd24552, 16'd64376, 16'd39136, 16'd65013, 16'd52690, 16'd20820, 16'd33896, 16'd57061, 16'd131, 16'd4220, 16'd52613, 16'd5480});
	test_expansion(128'ha817c34865bec23e124fbebe4f870abe, {16'd59401, 16'd13382, 16'd42466, 16'd28418, 16'd46786, 16'd26429, 16'd31085, 16'd29469, 16'd44412, 16'd8861, 16'd63056, 16'd8372, 16'd44403, 16'd55473, 16'd15320, 16'd5457, 16'd15241, 16'd11689, 16'd34403, 16'd46346, 16'd57652, 16'd41696, 16'd45757, 16'd30466, 16'd3980, 16'd40736});
	test_expansion(128'h6f0938377790093bb331d2d969f8e51d, {16'd21019, 16'd52109, 16'd53396, 16'd56104, 16'd50415, 16'd16030, 16'd20176, 16'd61116, 16'd10539, 16'd42452, 16'd41618, 16'd57113, 16'd31452, 16'd47125, 16'd12760, 16'd28315, 16'd36343, 16'd42916, 16'd15990, 16'd36829, 16'd57867, 16'd53043, 16'd64050, 16'd32917, 16'd29505, 16'd34968});
	test_expansion(128'h298a4fd0b0374b56c2c12b6df97ccca4, {16'd63588, 16'd35217, 16'd47718, 16'd3727, 16'd29371, 16'd25673, 16'd53297, 16'd10259, 16'd9100, 16'd37585, 16'd343, 16'd22966, 16'd26032, 16'd44695, 16'd33615, 16'd49440, 16'd6291, 16'd29059, 16'd40469, 16'd1195, 16'd14390, 16'd17955, 16'd59307, 16'd57990, 16'd17251, 16'd60484});
	test_expansion(128'hbf641167b551f9a4ee0b1a7eb98ed36b, {16'd31426, 16'd31612, 16'd7840, 16'd50475, 16'd30449, 16'd8502, 16'd33781, 16'd62936, 16'd47802, 16'd44972, 16'd9524, 16'd51526, 16'd51040, 16'd59359, 16'd35231, 16'd61442, 16'd21035, 16'd45344, 16'd52427, 16'd4033, 16'd11757, 16'd35824, 16'd25608, 16'd17687, 16'd8414, 16'd45217});
	test_expansion(128'h98c0e943d523422978efc59798798bd1, {16'd16233, 16'd55371, 16'd51034, 16'd20837, 16'd2465, 16'd20592, 16'd62240, 16'd26083, 16'd15619, 16'd60929, 16'd2581, 16'd46755, 16'd41992, 16'd13355, 16'd23866, 16'd1053, 16'd58709, 16'd46645, 16'd51370, 16'd40991, 16'd61405, 16'd53837, 16'd10580, 16'd6654, 16'd63932, 16'd4201});
	test_expansion(128'h98864f271055a981f8903fede136a681, {16'd16061, 16'd3140, 16'd10123, 16'd62470, 16'd28600, 16'd16235, 16'd61161, 16'd62221, 16'd31523, 16'd17659, 16'd61894, 16'd22786, 16'd12850, 16'd28821, 16'd53427, 16'd58988, 16'd19365, 16'd5554, 16'd48623, 16'd16392, 16'd61429, 16'd48199, 16'd44377, 16'd971, 16'd56368, 16'd15206});
	test_expansion(128'h1a2d1a9cfbb747a399240c8a407a24a4, {16'd61904, 16'd34903, 16'd34219, 16'd28818, 16'd45779, 16'd35505, 16'd35652, 16'd38320, 16'd11556, 16'd8944, 16'd10010, 16'd65087, 16'd25586, 16'd20219, 16'd2063, 16'd37826, 16'd6202, 16'd26281, 16'd43442, 16'd56151, 16'd59830, 16'd54397, 16'd17466, 16'd39234, 16'd10295, 16'd1757});
	test_expansion(128'h69d33f24a7896d8934c3da0a1a3d082b, {16'd29801, 16'd39289, 16'd65309, 16'd33258, 16'd23067, 16'd62502, 16'd17071, 16'd11166, 16'd63438, 16'd43052, 16'd28643, 16'd30669, 16'd9935, 16'd54899, 16'd31624, 16'd44195, 16'd5093, 16'd19675, 16'd5105, 16'd29336, 16'd32249, 16'd62124, 16'd22806, 16'd10317, 16'd2473, 16'd24999});
	test_expansion(128'h5145d6850c6eabb7c378ca36bb159e7d, {16'd47448, 16'd8446, 16'd53074, 16'd49752, 16'd62625, 16'd51386, 16'd18348, 16'd15432, 16'd9365, 16'd21638, 16'd53633, 16'd56144, 16'd49717, 16'd49094, 16'd42900, 16'd12918, 16'd22659, 16'd64135, 16'd5278, 16'd20880, 16'd14832, 16'd50291, 16'd48490, 16'd3069, 16'd32715, 16'd25613});
	test_expansion(128'hbbefcd48f3d29e658c2a92de2d6f7268, {16'd6999, 16'd46205, 16'd52502, 16'd22676, 16'd4942, 16'd407, 16'd44331, 16'd40609, 16'd27148, 16'd36197, 16'd42639, 16'd52802, 16'd3566, 16'd46995, 16'd28093, 16'd10620, 16'd42149, 16'd54821, 16'd59740, 16'd49604, 16'd52023, 16'd3050, 16'd59849, 16'd45301, 16'd61196, 16'd29476});
	test_expansion(128'h924054694ce4157f54463942645bc4dd, {16'd61599, 16'd53201, 16'd49550, 16'd8133, 16'd15816, 16'd31695, 16'd29591, 16'd58531, 16'd4384, 16'd33519, 16'd11822, 16'd1067, 16'd13954, 16'd22936, 16'd31878, 16'd14031, 16'd2518, 16'd147, 16'd19964, 16'd15077, 16'd35042, 16'd9995, 16'd41545, 16'd51710, 16'd42502, 16'd43445});
	test_expansion(128'h478fa1acf735e4f868360f3db727c7c1, {16'd26267, 16'd38279, 16'd15227, 16'd25937, 16'd56217, 16'd44686, 16'd40205, 16'd49592, 16'd46970, 16'd49440, 16'd51202, 16'd27777, 16'd32499, 16'd42421, 16'd35595, 16'd4543, 16'd46104, 16'd54100, 16'd62038, 16'd46322, 16'd38619, 16'd11239, 16'd62652, 16'd53935, 16'd44417, 16'd64497});
	test_expansion(128'h1e19bd4b313593372ecebc724c48a894, {16'd31719, 16'd43427, 16'd10756, 16'd32550, 16'd40400, 16'd57596, 16'd15594, 16'd16381, 16'd51120, 16'd48372, 16'd45586, 16'd793, 16'd5226, 16'd5518, 16'd26124, 16'd35395, 16'd47671, 16'd36927, 16'd24802, 16'd39628, 16'd3411, 16'd53298, 16'd54397, 16'd53915, 16'd25991, 16'd40435});
	test_expansion(128'h99d4a169a74708bbc9556b9361268d2c, {16'd28001, 16'd64656, 16'd33401, 16'd22666, 16'd8837, 16'd37887, 16'd56415, 16'd12204, 16'd2203, 16'd24760, 16'd57064, 16'd56115, 16'd21806, 16'd51218, 16'd48087, 16'd11797, 16'd31826, 16'd52140, 16'd2159, 16'd26077, 16'd56204, 16'd47900, 16'd40799, 16'd22668, 16'd20015, 16'd11750});
	test_expansion(128'hbc0177769215e051c879d1e470f6614f, {16'd20044, 16'd21363, 16'd14169, 16'd22587, 16'd34661, 16'd40674, 16'd52968, 16'd8091, 16'd22727, 16'd11136, 16'd44759, 16'd38349, 16'd37277, 16'd38134, 16'd21471, 16'd48389, 16'd31660, 16'd40594, 16'd17793, 16'd29106, 16'd25387, 16'd49239, 16'd63811, 16'd15969, 16'd24183, 16'd14544});
	test_expansion(128'h963a7143cca2b573e3a1692b0b72bb08, {16'd13403, 16'd52693, 16'd47432, 16'd50622, 16'd49486, 16'd13979, 16'd23758, 16'd45164, 16'd41126, 16'd64792, 16'd891, 16'd58289, 16'd1771, 16'd62904, 16'd52179, 16'd18139, 16'd14525, 16'd40652, 16'd31707, 16'd54573, 16'd48097, 16'd360, 16'd54444, 16'd16234, 16'd6329, 16'd34499});
	test_expansion(128'h97fa386ffb2530dcad141834e45757a6, {16'd59498, 16'd14755, 16'd25323, 16'd41060, 16'd49887, 16'd55316, 16'd14515, 16'd46049, 16'd18883, 16'd36540, 16'd46784, 16'd14408, 16'd30011, 16'd63046, 16'd40406, 16'd39628, 16'd52169, 16'd13301, 16'd25469, 16'd59843, 16'd22217, 16'd15616, 16'd4672, 16'd39323, 16'd10403, 16'd48125});
	test_expansion(128'h2fdb0490e68af04fc47b4f6432d04004, {16'd4311, 16'd4374, 16'd13814, 16'd33367, 16'd47949, 16'd24927, 16'd35283, 16'd52855, 16'd63715, 16'd35045, 16'd1056, 16'd8729, 16'd4008, 16'd38912, 16'd24913, 16'd30064, 16'd26654, 16'd56054, 16'd30953, 16'd46598, 16'd13909, 16'd16958, 16'd54336, 16'd65429, 16'd49456, 16'd52853});
	test_expansion(128'h54500d38800f9119e25ae1f0bb8fe381, {16'd49505, 16'd27343, 16'd31057, 16'd62561, 16'd32534, 16'd9993, 16'd3436, 16'd12129, 16'd39455, 16'd28066, 16'd52129, 16'd18206, 16'd51474, 16'd5753, 16'd19224, 16'd49374, 16'd6721, 16'd52417, 16'd25649, 16'd30749, 16'd23492, 16'd29309, 16'd52837, 16'd24074, 16'd4560, 16'd12094});
	test_expansion(128'h4ca899725c5ebe8a5baead6c6fafedb4, {16'd8767, 16'd8325, 16'd2255, 16'd59123, 16'd51674, 16'd53241, 16'd43858, 16'd37319, 16'd39368, 16'd16530, 16'd44475, 16'd34506, 16'd20309, 16'd1386, 16'd20747, 16'd41422, 16'd25462, 16'd4170, 16'd38909, 16'd40989, 16'd7828, 16'd28390, 16'd10371, 16'd55417, 16'd34438, 16'd57658});
	test_expansion(128'h335bcb062586809349a724912082b85b, {16'd6005, 16'd65339, 16'd47048, 16'd44773, 16'd38725, 16'd63211, 16'd10944, 16'd46861, 16'd25753, 16'd35449, 16'd48655, 16'd17623, 16'd56025, 16'd64103, 16'd51226, 16'd8032, 16'd36261, 16'd43608, 16'd22540, 16'd11639, 16'd61262, 16'd46835, 16'd8414, 16'd43817, 16'd39106, 16'd65228});
	test_expansion(128'h7e260bfeb257caf1bf70621db541a8b7, {16'd24398, 16'd31471, 16'd17698, 16'd3207, 16'd2783, 16'd47870, 16'd32303, 16'd10627, 16'd10268, 16'd8513, 16'd59925, 16'd35986, 16'd19407, 16'd60168, 16'd4845, 16'd31355, 16'd26571, 16'd29482, 16'd40282, 16'd58915, 16'd56663, 16'd29564, 16'd59858, 16'd39304, 16'd11349, 16'd17637});
	test_expansion(128'h803b70e6c788e3a8cd0d72b23585f5d9, {16'd10682, 16'd64124, 16'd34452, 16'd33773, 16'd57893, 16'd47267, 16'd42629, 16'd9799, 16'd15449, 16'd46176, 16'd50744, 16'd63446, 16'd41326, 16'd43911, 16'd38462, 16'd30157, 16'd55292, 16'd13747, 16'd11774, 16'd19400, 16'd55335, 16'd21265, 16'd38259, 16'd10588, 16'd7041, 16'd7573});
	test_expansion(128'hef546bda49be3265431bf35a3574fc65, {16'd47391, 16'd57263, 16'd24326, 16'd29912, 16'd10891, 16'd22437, 16'd51837, 16'd64014, 16'd28835, 16'd20969, 16'd16861, 16'd45591, 16'd56541, 16'd47985, 16'd40747, 16'd17328, 16'd30848, 16'd42968, 16'd55294, 16'd62738, 16'd24104, 16'd37213, 16'd1021, 16'd3746, 16'd48138, 16'd49394});
	test_expansion(128'h4b770b0c54bee9e564c20cb297198615, {16'd29571, 16'd33570, 16'd51475, 16'd19427, 16'd46589, 16'd48036, 16'd2454, 16'd4441, 16'd61235, 16'd23256, 16'd27409, 16'd25913, 16'd9631, 16'd22641, 16'd42792, 16'd38290, 16'd17258, 16'd1339, 16'd10140, 16'd8320, 16'd60775, 16'd9580, 16'd27265, 16'd15729, 16'd65379, 16'd60517});
	test_expansion(128'hc0abad9dd8e197e79ce300214954e40e, {16'd24454, 16'd52805, 16'd1401, 16'd10685, 16'd7601, 16'd56722, 16'd45497, 16'd65301, 16'd31659, 16'd54112, 16'd33484, 16'd16006, 16'd23927, 16'd56128, 16'd15131, 16'd30360, 16'd46067, 16'd61119, 16'd48711, 16'd23366, 16'd28677, 16'd49472, 16'd63945, 16'd50270, 16'd50858, 16'd34771});
	test_expansion(128'h61a0d9b13bf9b70281dbc6472763a6a9, {16'd52940, 16'd4132, 16'd40545, 16'd48334, 16'd36552, 16'd48025, 16'd58429, 16'd35580, 16'd7485, 16'd37320, 16'd47467, 16'd64098, 16'd45095, 16'd25550, 16'd2298, 16'd53692, 16'd10801, 16'd42982, 16'd57785, 16'd43366, 16'd63823, 16'd56758, 16'd31192, 16'd35703, 16'd9826, 16'd40516});
	test_expansion(128'h42d4cc8c3fe7bf04bdfce84b622cfe64, {16'd17720, 16'd63193, 16'd58143, 16'd2611, 16'd33886, 16'd53337, 16'd46989, 16'd65338, 16'd15922, 16'd13964, 16'd21342, 16'd37583, 16'd42017, 16'd8587, 16'd15393, 16'd24790, 16'd358, 16'd34837, 16'd62898, 16'd54874, 16'd49423, 16'd35307, 16'd24260, 16'd45391, 16'd38561, 16'd61618});
	test_expansion(128'haba224ceb7cd42953b96aab7ef86ff0b, {16'd36940, 16'd30082, 16'd44807, 16'd10794, 16'd44542, 16'd406, 16'd13850, 16'd26913, 16'd26624, 16'd51097, 16'd6318, 16'd62366, 16'd21790, 16'd51618, 16'd8931, 16'd48982, 16'd41744, 16'd61524, 16'd22183, 16'd6009, 16'd61378, 16'd46110, 16'd15357, 16'd57146, 16'd58163, 16'd40687});
	test_expansion(128'h5eb1c59286b1ddc33832d7e27fddaa1a, {16'd19156, 16'd33961, 16'd51918, 16'd32330, 16'd26649, 16'd17438, 16'd58625, 16'd57773, 16'd6443, 16'd49962, 16'd32255, 16'd5855, 16'd63085, 16'd44574, 16'd50867, 16'd32817, 16'd31482, 16'd9262, 16'd28027, 16'd55980, 16'd19798, 16'd16378, 16'd56477, 16'd49962, 16'd30212, 16'd19986});
	test_expansion(128'h09005eb8b30f38347b2d2029e80713e4, {16'd35822, 16'd5533, 16'd57646, 16'd35043, 16'd45352, 16'd3572, 16'd26076, 16'd18260, 16'd46543, 16'd57140, 16'd28841, 16'd21522, 16'd60759, 16'd1359, 16'd65024, 16'd43855, 16'd20915, 16'd62658, 16'd6088, 16'd44292, 16'd37381, 16'd45983, 16'd61270, 16'd22747, 16'd21743, 16'd31830});
	test_expansion(128'h669bae11b26db6507edb2b835c4c06f8, {16'd4274, 16'd904, 16'd10476, 16'd12826, 16'd27264, 16'd59256, 16'd38001, 16'd56938, 16'd4386, 16'd18652, 16'd61373, 16'd60956, 16'd36225, 16'd14881, 16'd60316, 16'd65036, 16'd61284, 16'd61124, 16'd39608, 16'd21157, 16'd28111, 16'd24656, 16'd49390, 16'd27133, 16'd22689, 16'd50979});
	test_expansion(128'hde76ea90c8aa4f39fb1705bbe11471e4, {16'd6493, 16'd59964, 16'd33254, 16'd7468, 16'd21753, 16'd37912, 16'd19257, 16'd47271, 16'd3493, 16'd34377, 16'd41973, 16'd35981, 16'd604, 16'd60712, 16'd7035, 16'd27749, 16'd51337, 16'd4875, 16'd42825, 16'd22541, 16'd36333, 16'd35994, 16'd54133, 16'd26164, 16'd6623, 16'd44476});
	test_expansion(128'h372bad30a70b0983ccd41a43d1612f62, {16'd43483, 16'd27863, 16'd47485, 16'd65263, 16'd56394, 16'd60201, 16'd46441, 16'd61078, 16'd62026, 16'd51231, 16'd52014, 16'd47130, 16'd3739, 16'd3363, 16'd11871, 16'd39055, 16'd13327, 16'd64293, 16'd6733, 16'd62797, 16'd30023, 16'd52496, 16'd51811, 16'd43436, 16'd29705, 16'd20702});
	test_expansion(128'h329fb4f41ee028d551ced6bce12c2a07, {16'd57724, 16'd22850, 16'd57540, 16'd15735, 16'd37922, 16'd30083, 16'd3024, 16'd17342, 16'd2408, 16'd10159, 16'd56045, 16'd57986, 16'd21424, 16'd39070, 16'd825, 16'd41736, 16'd10426, 16'd55260, 16'd32049, 16'd26951, 16'd26437, 16'd1101, 16'd22467, 16'd6001, 16'd52511, 16'd237});
	test_expansion(128'h1e68552806a65abef32499745004e880, {16'd6608, 16'd7718, 16'd50685, 16'd16495, 16'd33182, 16'd31680, 16'd53278, 16'd21270, 16'd51377, 16'd7709, 16'd61602, 16'd35415, 16'd64491, 16'd56576, 16'd43548, 16'd5222, 16'd9960, 16'd2127, 16'd61447, 16'd29305, 16'd1077, 16'd36698, 16'd59826, 16'd29289, 16'd27225, 16'd26351});
	test_expansion(128'h280bc687c893e9222e26b399975338f1, {16'd22664, 16'd6250, 16'd48233, 16'd38801, 16'd44921, 16'd44279, 16'd39322, 16'd54295, 16'd27385, 16'd197, 16'd38507, 16'd44259, 16'd45786, 16'd9006, 16'd1616, 16'd10387, 16'd4339, 16'd58703, 16'd32055, 16'd65185, 16'd39596, 16'd60691, 16'd42086, 16'd63266, 16'd12808, 16'd3193});
	test_expansion(128'h63c754e8105bb37d627165cc16b8dd2a, {16'd15285, 16'd37660, 16'd2753, 16'd59111, 16'd4303, 16'd30519, 16'd37098, 16'd52834, 16'd49122, 16'd59891, 16'd23812, 16'd50684, 16'd41305, 16'd20360, 16'd11373, 16'd25316, 16'd35628, 16'd42077, 16'd43943, 16'd57014, 16'd42854, 16'd43760, 16'd17844, 16'd58297, 16'd12543, 16'd53161});
	test_expansion(128'h1812850b344a0eef0c11c77f5a5c58aa, {16'd43378, 16'd27172, 16'd56877, 16'd58165, 16'd57332, 16'd41539, 16'd48532, 16'd57187, 16'd49393, 16'd41077, 16'd64297, 16'd63563, 16'd23635, 16'd6351, 16'd31852, 16'd63946, 16'd2453, 16'd50382, 16'd18160, 16'd42422, 16'd31322, 16'd33630, 16'd25702, 16'd13705, 16'd61604, 16'd10702});
	test_expansion(128'h757dd87e59d811aea5b41d84caa8c8bb, {16'd37713, 16'd8111, 16'd39722, 16'd33000, 16'd31028, 16'd63508, 16'd31528, 16'd12626, 16'd33036, 16'd25897, 16'd2959, 16'd7449, 16'd28243, 16'd17623, 16'd33886, 16'd8524, 16'd50572, 16'd27204, 16'd61495, 16'd27440, 16'd14464, 16'd33469, 16'd40334, 16'd8376, 16'd47688, 16'd4545});
	test_expansion(128'h1b16724cdf3e0a630cae3babc66afeb8, {16'd30922, 16'd3402, 16'd1646, 16'd30433, 16'd11806, 16'd13332, 16'd42608, 16'd64663, 16'd42490, 16'd58302, 16'd2326, 16'd15732, 16'd12496, 16'd62683, 16'd1984, 16'd23979, 16'd17628, 16'd2136, 16'd21558, 16'd60608, 16'd47211, 16'd51378, 16'd52871, 16'd9903, 16'd20383, 16'd17820});
	test_expansion(128'h93647d02938bff52cb6a9b9022c60e02, {16'd51745, 16'd65410, 16'd28006, 16'd50483, 16'd25797, 16'd22453, 16'd4930, 16'd2423, 16'd29811, 16'd15935, 16'd18496, 16'd59138, 16'd6531, 16'd9545, 16'd16469, 16'd27498, 16'd26221, 16'd30033, 16'd17569, 16'd20487, 16'd46467, 16'd61457, 16'd43626, 16'd63555, 16'd1535, 16'd50272});
	test_expansion(128'hcad61186668697802df2de7ba0cda6fe, {16'd44112, 16'd53536, 16'd16614, 16'd6491, 16'd48109, 16'd34387, 16'd54695, 16'd43626, 16'd19768, 16'd25889, 16'd47496, 16'd25592, 16'd15406, 16'd2401, 16'd11985, 16'd6133, 16'd24130, 16'd1704, 16'd23038, 16'd23340, 16'd23383, 16'd22329, 16'd29390, 16'd3884, 16'd57378, 16'd52766});
	test_expansion(128'hf310b04005bb98bc25372790e02e64b2, {16'd10294, 16'd5540, 16'd44064, 16'd29162, 16'd49684, 16'd55999, 16'd12465, 16'd38847, 16'd61228, 16'd24824, 16'd12458, 16'd21298, 16'd32315, 16'd43470, 16'd54164, 16'd32908, 16'd48317, 16'd18678, 16'd41323, 16'd44227, 16'd62547, 16'd16071, 16'd47107, 16'd19128, 16'd61018, 16'd4587});
	test_expansion(128'he048f9a5f1bdeb03f54543492377384e, {16'd27370, 16'd50241, 16'd40774, 16'd63482, 16'd15070, 16'd55775, 16'd12209, 16'd58209, 16'd37279, 16'd6353, 16'd50178, 16'd8207, 16'd42922, 16'd49326, 16'd46395, 16'd32416, 16'd40064, 16'd10338, 16'd34615, 16'd41185, 16'd37456, 16'd49786, 16'd2897, 16'd21497, 16'd5294, 16'd29295});
	test_expansion(128'h9607ccc1aadff08e8a53ad3ef6c84b62, {16'd62720, 16'd55604, 16'd48793, 16'd21950, 16'd7510, 16'd23007, 16'd9572, 16'd21645, 16'd18595, 16'd18196, 16'd7553, 16'd25294, 16'd37089, 16'd44698, 16'd44173, 16'd13008, 16'd14471, 16'd14012, 16'd238, 16'd50448, 16'd41238, 16'd46526, 16'd54358, 16'd47832, 16'd4891, 16'd22979});
	test_expansion(128'h719ffe8bc28cdb68a8644bbb40665981, {16'd32338, 16'd64983, 16'd54231, 16'd22626, 16'd54439, 16'd36740, 16'd3258, 16'd40584, 16'd30472, 16'd4069, 16'd22167, 16'd13285, 16'd52285, 16'd17143, 16'd32060, 16'd64867, 16'd60383, 16'd232, 16'd18170, 16'd49173, 16'd41591, 16'd49616, 16'd22731, 16'd13943, 16'd592, 16'd55124});
	test_expansion(128'h77c08d8cba7b54b7d84f855858a99abf, {16'd45156, 16'd60602, 16'd59791, 16'd11163, 16'd46359, 16'd19492, 16'd7172, 16'd31727, 16'd18491, 16'd25864, 16'd20287, 16'd13691, 16'd55326, 16'd34925, 16'd37232, 16'd49855, 16'd16498, 16'd2876, 16'd28928, 16'd39794, 16'd48005, 16'd15323, 16'd31728, 16'd16755, 16'd62180, 16'd41940});
	test_expansion(128'h5cc0b5c3843c8620c7e40f7fb04c7b52, {16'd64251, 16'd21302, 16'd21244, 16'd39814, 16'd10481, 16'd39074, 16'd26960, 16'd50352, 16'd43433, 16'd15212, 16'd40529, 16'd29540, 16'd40007, 16'd63907, 16'd54393, 16'd19297, 16'd44273, 16'd60809, 16'd30198, 16'd58584, 16'd14805, 16'd63234, 16'd35171, 16'd45884, 16'd50762, 16'd8457});
	test_expansion(128'hb9cdbe8ce24059b34786b5969f1b4b8d, {16'd5341, 16'd14569, 16'd2023, 16'd29717, 16'd9294, 16'd40163, 16'd61564, 16'd58650, 16'd58434, 16'd1479, 16'd26448, 16'd35070, 16'd58784, 16'd40727, 16'd35203, 16'd58496, 16'd47702, 16'd28444, 16'd37982, 16'd44772, 16'd18478, 16'd17461, 16'd53217, 16'd9202, 16'd24309, 16'd63050});
	test_expansion(128'hac81728cdd85017b6001a00e502d4a05, {16'd35167, 16'd36772, 16'd32563, 16'd1576, 16'd49316, 16'd29945, 16'd33649, 16'd28601, 16'd10802, 16'd64110, 16'd10687, 16'd18626, 16'd35319, 16'd54520, 16'd14758, 16'd35286, 16'd36408, 16'd29192, 16'd9122, 16'd30163, 16'd62418, 16'd9991, 16'd62158, 16'd34896, 16'd18619, 16'd59551});
	test_expansion(128'h67d5cfde6ce3cfbc0a00d031101cd267, {16'd61895, 16'd52193, 16'd41280, 16'd57052, 16'd45772, 16'd33547, 16'd58481, 16'd44776, 16'd47978, 16'd51870, 16'd60579, 16'd18679, 16'd25236, 16'd61993, 16'd30145, 16'd62186, 16'd1058, 16'd15237, 16'd37464, 16'd21037, 16'd56343, 16'd831, 16'd47468, 16'd36032, 16'd42029, 16'd27156});
	test_expansion(128'h7f1f049d037c5dc3aac1956d7694e1e7, {16'd34539, 16'd55818, 16'd42444, 16'd22672, 16'd26413, 16'd27852, 16'd37185, 16'd21824, 16'd56862, 16'd22818, 16'd42539, 16'd36531, 16'd33315, 16'd57759, 16'd39669, 16'd33925, 16'd60104, 16'd6563, 16'd33146, 16'd33825, 16'd44726, 16'd56143, 16'd63673, 16'd48908, 16'd46011, 16'd29817});
	test_expansion(128'h84677d8891c034712077732b80cf4921, {16'd45552, 16'd42172, 16'd34208, 16'd49002, 16'd45604, 16'd1969, 16'd57139, 16'd9828, 16'd23634, 16'd42349, 16'd9643, 16'd63789, 16'd43248, 16'd12371, 16'd4803, 16'd32598, 16'd4408, 16'd41532, 16'd52818, 16'd30092, 16'd20201, 16'd53619, 16'd32179, 16'd59996, 16'd23880, 16'd53713});
	test_expansion(128'h695a35804ae023b762b5a24d9da78b3c, {16'd44467, 16'd36977, 16'd27432, 16'd53370, 16'd9834, 16'd42657, 16'd42600, 16'd59717, 16'd36815, 16'd46499, 16'd58610, 16'd43995, 16'd54854, 16'd28852, 16'd60005, 16'd30138, 16'd53157, 16'd30076, 16'd25384, 16'd5891, 16'd14310, 16'd4899, 16'd19010, 16'd36979, 16'd39478, 16'd42411});
	test_expansion(128'h9f29df01b747e82e6d90e61ac8798f8d, {16'd38324, 16'd64001, 16'd17530, 16'd10876, 16'd59701, 16'd29676, 16'd60508, 16'd18535, 16'd47759, 16'd20624, 16'd224, 16'd29278, 16'd43911, 16'd59175, 16'd14067, 16'd11261, 16'd62789, 16'd47584, 16'd44485, 16'd3222, 16'd26566, 16'd6241, 16'd37114, 16'd20426, 16'd61646, 16'd33007});
	test_expansion(128'h9d375e15743029f76e654d7591515677, {16'd61648, 16'd16128, 16'd52876, 16'd28744, 16'd35086, 16'd22986, 16'd52532, 16'd60919, 16'd34052, 16'd27889, 16'd44273, 16'd45440, 16'd16312, 16'd55266, 16'd31318, 16'd46261, 16'd40308, 16'd45156, 16'd1699, 16'd42426, 16'd17200, 16'd16899, 16'd25995, 16'd8535, 16'd34852, 16'd15631});
	test_expansion(128'hdbfe5bcc49b6b79457ed2f5efb8de8e0, {16'd29121, 16'd30432, 16'd30914, 16'd49457, 16'd47349, 16'd64595, 16'd20586, 16'd39703, 16'd1854, 16'd17129, 16'd56195, 16'd10407, 16'd59804, 16'd32156, 16'd54531, 16'd31588, 16'd38463, 16'd3887, 16'd8295, 16'd57946, 16'd22701, 16'd4292, 16'd29595, 16'd57456, 16'd41679, 16'd19943});
	test_expansion(128'ha33ce777c71d720f74b36268adb76b6e, {16'd19423, 16'd38217, 16'd33767, 16'd17935, 16'd64195, 16'd28201, 16'd53237, 16'd46689, 16'd43702, 16'd52027, 16'd4795, 16'd55318, 16'd37318, 16'd23652, 16'd41053, 16'd22163, 16'd49223, 16'd16837, 16'd39887, 16'd39528, 16'd47495, 16'd32382, 16'd44140, 16'd10801, 16'd29292, 16'd37865});
	test_expansion(128'h51ceffc7a82d8241d41f037e6e0e330d, {16'd37661, 16'd64227, 16'd63212, 16'd51764, 16'd15277, 16'd62446, 16'd19167, 16'd53147, 16'd52240, 16'd27703, 16'd42254, 16'd138, 16'd11689, 16'd25746, 16'd44508, 16'd22574, 16'd12701, 16'd1623, 16'd26294, 16'd26844, 16'd35610, 16'd1000, 16'd53061, 16'd37373, 16'd65167, 16'd20977});
	test_expansion(128'he074b58124d1e5b9c9682fcc9e1165a9, {16'd55318, 16'd62988, 16'd6607, 16'd32195, 16'd27289, 16'd54334, 16'd50028, 16'd44215, 16'd43313, 16'd53721, 16'd19344, 16'd43951, 16'd37927, 16'd28553, 16'd38519, 16'd632, 16'd27051, 16'd60502, 16'd3727, 16'd6620, 16'd30366, 16'd13190, 16'd14010, 16'd63435, 16'd47460, 16'd12963});
	test_expansion(128'h180cdf4227b097d6e16dbaa0072decaf, {16'd2077, 16'd13258, 16'd1141, 16'd8613, 16'd14586, 16'd58209, 16'd5104, 16'd64289, 16'd18831, 16'd41711, 16'd54629, 16'd20050, 16'd15259, 16'd59617, 16'd44214, 16'd43606, 16'd55373, 16'd62107, 16'd18424, 16'd39977, 16'd17895, 16'd62610, 16'd43856, 16'd54454, 16'd34585, 16'd50540});
	test_expansion(128'h352a416debf83dd86862e438aa36337d, {16'd47830, 16'd545, 16'd60526, 16'd9949, 16'd8447, 16'd46042, 16'd41915, 16'd4900, 16'd47975, 16'd10753, 16'd62532, 16'd7658, 16'd30314, 16'd54970, 16'd30422, 16'd7569, 16'd44250, 16'd57262, 16'd40492, 16'd21526, 16'd8593, 16'd17537, 16'd15525, 16'd9323, 16'd47431, 16'd9914});
	test_expansion(128'hef88bd0922e489b0875bf4e9f267fbbc, {16'd61616, 16'd50020, 16'd64736, 16'd234, 16'd57814, 16'd43299, 16'd7784, 16'd46069, 16'd21317, 16'd51215, 16'd42501, 16'd17689, 16'd15244, 16'd14296, 16'd59341, 16'd60624, 16'd53788, 16'd46952, 16'd25469, 16'd9897, 16'd57048, 16'd57025, 16'd34614, 16'd57418, 16'd5389, 16'd9061});
	test_expansion(128'hd9441caa1024cdb2309bda8748f54522, {16'd2434, 16'd58005, 16'd59989, 16'd35735, 16'd39692, 16'd10063, 16'd41814, 16'd5750, 16'd36165, 16'd41443, 16'd9043, 16'd29076, 16'd54338, 16'd32962, 16'd20836, 16'd46085, 16'd57029, 16'd49388, 16'd25107, 16'd33338, 16'd8553, 16'd38399, 16'd51772, 16'd26924, 16'd17729, 16'd28790});
	test_expansion(128'hd3877467457d5c641b9e81337a8c44bd, {16'd53021, 16'd60168, 16'd8157, 16'd56236, 16'd57044, 16'd19994, 16'd3125, 16'd14044, 16'd17699, 16'd58340, 16'd45777, 16'd57576, 16'd21151, 16'd40404, 16'd47898, 16'd30367, 16'd47157, 16'd31482, 16'd36415, 16'd22518, 16'd52306, 16'd41738, 16'd17067, 16'd43564, 16'd5599, 16'd17131});
	test_expansion(128'h030b2417ebfefb7a73a1e4703e58a54f, {16'd64952, 16'd49427, 16'd5979, 16'd48096, 16'd44470, 16'd44892, 16'd12289, 16'd43180, 16'd47119, 16'd36628, 16'd36119, 16'd15794, 16'd36857, 16'd961, 16'd34454, 16'd14760, 16'd18493, 16'd10433, 16'd54106, 16'd36111, 16'd19706, 16'd53393, 16'd52182, 16'd18508, 16'd13124, 16'd12987});
	test_expansion(128'hf49d29ea27321141d58f6edb156a8269, {16'd50872, 16'd61566, 16'd20233, 16'd10189, 16'd5640, 16'd29941, 16'd60089, 16'd60592, 16'd21765, 16'd6421, 16'd5541, 16'd28115, 16'd64481, 16'd62907, 16'd22593, 16'd47228, 16'd27587, 16'd57824, 16'd45121, 16'd7880, 16'd6573, 16'd26030, 16'd59019, 16'd21853, 16'd61636, 16'd60369});
	test_expansion(128'h440f65fc1c3b301f1937b22f2572e3a8, {16'd26636, 16'd1503, 16'd10500, 16'd60811, 16'd55955, 16'd40793, 16'd15897, 16'd61427, 16'd23928, 16'd24619, 16'd57669, 16'd4865, 16'd9580, 16'd27918, 16'd62649, 16'd51547, 16'd35647, 16'd14671, 16'd60627, 16'd6955, 16'd24889, 16'd37919, 16'd18809, 16'd5303, 16'd1037, 16'd11288});
	test_expansion(128'h7e8244e9efac63dff3705bcfa2eded58, {16'd22833, 16'd29666, 16'd31527, 16'd39527, 16'd20989, 16'd31841, 16'd50044, 16'd42821, 16'd46636, 16'd40266, 16'd2710, 16'd53045, 16'd3842, 16'd14340, 16'd8089, 16'd52662, 16'd38618, 16'd25187, 16'd24196, 16'd15039, 16'd14620, 16'd39804, 16'd24078, 16'd64314, 16'd63087, 16'd36250});
	test_expansion(128'h20b994f8fe6b9ce1dbfe6d4424e9a20a, {16'd17017, 16'd29760, 16'd48418, 16'd59128, 16'd4529, 16'd58968, 16'd60458, 16'd63498, 16'd19699, 16'd21876, 16'd6721, 16'd11687, 16'd27715, 16'd49199, 16'd28319, 16'd4471, 16'd7415, 16'd50199, 16'd19394, 16'd19329, 16'd38681, 16'd396, 16'd2963, 16'd33016, 16'd19525, 16'd42862});
	test_expansion(128'h257bbbbd246d86c02b2554adba5282d0, {16'd14259, 16'd49505, 16'd21550, 16'd15848, 16'd4444, 16'd54467, 16'd39977, 16'd22403, 16'd30269, 16'd16887, 16'd8764, 16'd1451, 16'd58218, 16'd36431, 16'd47987, 16'd1676, 16'd11442, 16'd58353, 16'd60388, 16'd5957, 16'd30352, 16'd43579, 16'd54646, 16'd9004, 16'd51286, 16'd20512});
	test_expansion(128'h6b45937a51a7ba7380959f68191b1c31, {16'd63609, 16'd62155, 16'd1122, 16'd59714, 16'd64684, 16'd18041, 16'd44939, 16'd4097, 16'd16913, 16'd164, 16'd25944, 16'd6367, 16'd13085, 16'd48778, 16'd28496, 16'd47517, 16'd32364, 16'd1868, 16'd35103, 16'd63954, 16'd7394, 16'd36937, 16'd44201, 16'd17291, 16'd47567, 16'd61789});
	test_expansion(128'h57560e82af9751cb522769ab6145f0f1, {16'd33180, 16'd43308, 16'd56072, 16'd30451, 16'd55352, 16'd6860, 16'd27806, 16'd58687, 16'd32114, 16'd16676, 16'd35483, 16'd20671, 16'd25835, 16'd58325, 16'd50536, 16'd46393, 16'd45262, 16'd27012, 16'd48922, 16'd59365, 16'd30852, 16'd65400, 16'd53803, 16'd39685, 16'd32611, 16'd46045});
	test_expansion(128'ha60146cf6a5442854e931f7e21db58b4, {16'd18626, 16'd11322, 16'd39939, 16'd46436, 16'd39478, 16'd39467, 16'd59273, 16'd55348, 16'd4369, 16'd17176, 16'd8588, 16'd60766, 16'd27537, 16'd22395, 16'd56038, 16'd13306, 16'd11779, 16'd64992, 16'd48215, 16'd57672, 16'd46012, 16'd4817, 16'd3386, 16'd19886, 16'd51378, 16'd1262});
	test_expansion(128'hf2e7ab5d272f12dc738dbba765d9c27d, {16'd4815, 16'd25485, 16'd33659, 16'd26695, 16'd29947, 16'd58862, 16'd8926, 16'd59983, 16'd22163, 16'd60570, 16'd4609, 16'd46887, 16'd52748, 16'd30475, 16'd8294, 16'd16165, 16'd38897, 16'd19377, 16'd59734, 16'd36189, 16'd20352, 16'd30018, 16'd22937, 16'd57768, 16'd10549, 16'd19731});
	test_expansion(128'h9e65b85af88fb84fddf76ef8696fc841, {16'd9610, 16'd17396, 16'd42757, 16'd13697, 16'd43253, 16'd62928, 16'd43402, 16'd52516, 16'd43638, 16'd63825, 16'd64556, 16'd4004, 16'd36197, 16'd17260, 16'd7625, 16'd52389, 16'd13436, 16'd4873, 16'd56417, 16'd50086, 16'd45022, 16'd56258, 16'd56905, 16'd42551, 16'd44953, 16'd34011});
	test_expansion(128'he1beeeab7d04f928796407f92c9a9196, {16'd8029, 16'd59438, 16'd56930, 16'd56597, 16'd60573, 16'd13453, 16'd41368, 16'd23613, 16'd56687, 16'd31427, 16'd36606, 16'd1661, 16'd19601, 16'd60358, 16'd56279, 16'd17227, 16'd45199, 16'd49217, 16'd27902, 16'd60807, 16'd2149, 16'd5557, 16'd46437, 16'd53790, 16'd59804, 16'd6362});
	test_expansion(128'hdf549613fb03e8f728753757c97b5baf, {16'd65505, 16'd41238, 16'd57850, 16'd5166, 16'd29527, 16'd41968, 16'd10474, 16'd63973, 16'd31615, 16'd4152, 16'd1117, 16'd75, 16'd9080, 16'd35632, 16'd29393, 16'd23180, 16'd19002, 16'd64905, 16'd63343, 16'd52326, 16'd43627, 16'd8659, 16'd3277, 16'd15224, 16'd27901, 16'd44840});
	test_expansion(128'h609444854b1f940a613845de589bc3a5, {16'd34673, 16'd6837, 16'd63196, 16'd5056, 16'd59841, 16'd51720, 16'd43013, 16'd44078, 16'd57004, 16'd50119, 16'd62017, 16'd60871, 16'd9230, 16'd49909, 16'd8506, 16'd33838, 16'd46374, 16'd39315, 16'd14044, 16'd15698, 16'd57509, 16'd26019, 16'd16753, 16'd2066, 16'd12936, 16'd7509});
	test_expansion(128'h10d9572b0fa124c6e321fa19a3f11114, {16'd60210, 16'd23936, 16'd10726, 16'd13848, 16'd47562, 16'd36609, 16'd23455, 16'd19109, 16'd14468, 16'd10804, 16'd58367, 16'd38385, 16'd9844, 16'd45069, 16'd30192, 16'd62587, 16'd16854, 16'd23602, 16'd35228, 16'd2682, 16'd36647, 16'd64705, 16'd54604, 16'd31961, 16'd20815, 16'd51282});
	test_expansion(128'h8d1abdaf6aa23e7322019aca3415e0de, {16'd58396, 16'd12444, 16'd21982, 16'd10161, 16'd21629, 16'd50992, 16'd16098, 16'd60646, 16'd63559, 16'd54349, 16'd52397, 16'd13015, 16'd12690, 16'd8718, 16'd13853, 16'd4678, 16'd37144, 16'd17149, 16'd3781, 16'd35034, 16'd5958, 16'd24185, 16'd19745, 16'd65086, 16'd45341, 16'd5551});
	test_expansion(128'h78152a89f9529de54f5cf225fa9e223b, {16'd35788, 16'd62472, 16'd39402, 16'd53074, 16'd63075, 16'd64139, 16'd62071, 16'd35219, 16'd39459, 16'd27634, 16'd56408, 16'd26694, 16'd31521, 16'd25346, 16'd64934, 16'd24464, 16'd24613, 16'd24633, 16'd36245, 16'd24349, 16'd27250, 16'd7484, 16'd35464, 16'd52595, 16'd24668, 16'd62543});
	test_expansion(128'ha6534ccadee4bb8b2618e0fce6f24bea, {16'd31259, 16'd7473, 16'd6488, 16'd11367, 16'd47469, 16'd55546, 16'd63623, 16'd45940, 16'd61472, 16'd29434, 16'd15115, 16'd39373, 16'd34126, 16'd13057, 16'd47707, 16'd10938, 16'd17765, 16'd18274, 16'd29257, 16'd24595, 16'd62271, 16'd50650, 16'd11666, 16'd59247, 16'd30667, 16'd49562});
	test_expansion(128'h221a2925d61ee4963e144a5ab9c46632, {16'd48208, 16'd22639, 16'd16878, 16'd35408, 16'd33461, 16'd13885, 16'd51988, 16'd26368, 16'd53927, 16'd50569, 16'd20301, 16'd11690, 16'd32980, 16'd12151, 16'd26019, 16'd42963, 16'd18035, 16'd94, 16'd8782, 16'd10529, 16'd52186, 16'd17316, 16'd8776, 16'd7756, 16'd25655, 16'd48817});
	test_expansion(128'hf71da05b45307c8b4bcaabbb8758a8f8, {16'd14122, 16'd7982, 16'd42491, 16'd18168, 16'd54825, 16'd13472, 16'd25798, 16'd55427, 16'd17552, 16'd15579, 16'd4715, 16'd38202, 16'd40814, 16'd4379, 16'd60768, 16'd56981, 16'd58953, 16'd63430, 16'd59190, 16'd53368, 16'd51686, 16'd10928, 16'd47613, 16'd35204, 16'd14404, 16'd34992});
	test_expansion(128'h74c9fd385a615d86fcfe3c288c203edb, {16'd46881, 16'd14291, 16'd30889, 16'd44670, 16'd30864, 16'd48401, 16'd21703, 16'd62059, 16'd30997, 16'd46213, 16'd64005, 16'd54727, 16'd26532, 16'd56786, 16'd20093, 16'd4562, 16'd21033, 16'd5842, 16'd9674, 16'd60172, 16'd36743, 16'd64012, 16'd56113, 16'd62930, 16'd60771, 16'd29256});
	test_expansion(128'h59e3a01a252cf3e4e1279770066869e4, {16'd34569, 16'd3061, 16'd43563, 16'd32757, 16'd60613, 16'd62295, 16'd36760, 16'd43070, 16'd17825, 16'd30790, 16'd51856, 16'd63300, 16'd31284, 16'd2930, 16'd49435, 16'd58772, 16'd38469, 16'd15949, 16'd44980, 16'd26281, 16'd1589, 16'd6031, 16'd39446, 16'd34123, 16'd62770, 16'd57244});
	test_expansion(128'ha0ea9d65b278bbbf1378808949f2708b, {16'd5319, 16'd38660, 16'd46822, 16'd57278, 16'd38776, 16'd7565, 16'd59681, 16'd27891, 16'd54598, 16'd50099, 16'd59978, 16'd60820, 16'd50684, 16'd58120, 16'd8346, 16'd10901, 16'd39161, 16'd13210, 16'd20676, 16'd54514, 16'd57023, 16'd52147, 16'd56650, 16'd52945, 16'd3165, 16'd53589});
	test_expansion(128'hbf9149653eb6d418de38da05a2ca495f, {16'd2603, 16'd55599, 16'd6781, 16'd61877, 16'd55805, 16'd6475, 16'd29955, 16'd35054, 16'd24424, 16'd50248, 16'd12247, 16'd29892, 16'd5083, 16'd16712, 16'd7650, 16'd33515, 16'd18762, 16'd36826, 16'd54204, 16'd22624, 16'd26397, 16'd27340, 16'd43310, 16'd57524, 16'd13351, 16'd39957});
	test_expansion(128'h749f021128ae4355ff564f251523edda, {16'd53580, 16'd32801, 16'd8342, 16'd16865, 16'd25700, 16'd12760, 16'd25325, 16'd57319, 16'd7072, 16'd33164, 16'd12487, 16'd44794, 16'd37543, 16'd21730, 16'd59104, 16'd2207, 16'd43372, 16'd14740, 16'd57757, 16'd34054, 16'd28045, 16'd33478, 16'd33658, 16'd55834, 16'd1664, 16'd46961});
	test_expansion(128'h9de5da10ad514dfbf6379eaae300678c, {16'd52177, 16'd64889, 16'd11577, 16'd28009, 16'd7229, 16'd9357, 16'd40280, 16'd39635, 16'd41506, 16'd20917, 16'd39049, 16'd8057, 16'd58234, 16'd62929, 16'd56472, 16'd60568, 16'd35724, 16'd53741, 16'd7802, 16'd55304, 16'd119, 16'd58847, 16'd59401, 16'd5189, 16'd49820, 16'd2123});
	test_expansion(128'h449793dacf995ec6d3bfe32d58871b81, {16'd13324, 16'd61036, 16'd47780, 16'd12293, 16'd63712, 16'd24492, 16'd689, 16'd65390, 16'd19321, 16'd61877, 16'd19273, 16'd19539, 16'd47148, 16'd38671, 16'd63713, 16'd27268, 16'd63052, 16'd4481, 16'd12808, 16'd36511, 16'd49241, 16'd34603, 16'd25337, 16'd24287, 16'd2588, 16'd5933});
	test_expansion(128'haad68a3fd606e977ddcbbeef0bd5a47a, {16'd24586, 16'd59371, 16'd28455, 16'd30604, 16'd8503, 16'd8217, 16'd16925, 16'd26370, 16'd27483, 16'd64189, 16'd10206, 16'd54447, 16'd48801, 16'd56419, 16'd14056, 16'd41585, 16'd42948, 16'd30345, 16'd37681, 16'd10323, 16'd1464, 16'd16070, 16'd47937, 16'd1065, 16'd59595, 16'd50413});
	test_expansion(128'h42f7575a2cfb1ab8910c7b1f8aec9017, {16'd33142, 16'd62712, 16'd43221, 16'd43063, 16'd12985, 16'd28861, 16'd53285, 16'd65369, 16'd31970, 16'd38094, 16'd9101, 16'd62119, 16'd57062, 16'd44434, 16'd51531, 16'd10223, 16'd17151, 16'd1814, 16'd41463, 16'd16840, 16'd53039, 16'd10250, 16'd42630, 16'd50211, 16'd9752, 16'd43990});
	test_expansion(128'h4715bc6f5bb43ef2507dcf394a2e3274, {16'd35008, 16'd44815, 16'd34323, 16'd44385, 16'd22084, 16'd40270, 16'd49337, 16'd49754, 16'd39542, 16'd7604, 16'd64597, 16'd53368, 16'd2625, 16'd39064, 16'd50833, 16'd58398, 16'd17169, 16'd18605, 16'd33307, 16'd30844, 16'd1297, 16'd24214, 16'd12824, 16'd17001, 16'd53485, 16'd28388});
	test_expansion(128'h9b3cc35e2562f688add2f972fafc8dcd, {16'd37644, 16'd2164, 16'd3369, 16'd8999, 16'd52894, 16'd31752, 16'd50226, 16'd28580, 16'd36256, 16'd12583, 16'd25440, 16'd41589, 16'd29118, 16'd34099, 16'd59839, 16'd35996, 16'd10312, 16'd15968, 16'd28848, 16'd44431, 16'd23017, 16'd54849, 16'd34431, 16'd45073, 16'd32364, 16'd56278});
	test_expansion(128'h3226900c88f3f9293150704a06f24930, {16'd51847, 16'd54345, 16'd29778, 16'd47241, 16'd277, 16'd35898, 16'd16196, 16'd34964, 16'd2748, 16'd53386, 16'd42980, 16'd52285, 16'd55406, 16'd241, 16'd28688, 16'd34090, 16'd58658, 16'd31754, 16'd9262, 16'd45053, 16'd28727, 16'd47376, 16'd35365, 16'd40658, 16'd38514, 16'd42089});
	test_expansion(128'h07d01f18723e04389cf6f1f410a7726d, {16'd61970, 16'd55725, 16'd29681, 16'd65371, 16'd44074, 16'd22702, 16'd47837, 16'd38020, 16'd58643, 16'd51911, 16'd23911, 16'd11233, 16'd47813, 16'd35889, 16'd29948, 16'd13348, 16'd16895, 16'd65073, 16'd10362, 16'd22734, 16'd21978, 16'd22158, 16'd13039, 16'd6629, 16'd26378, 16'd42232});
	test_expansion(128'h201ed9dc68808d5970b1ce9fde5ab70d, {16'd40582, 16'd45184, 16'd38659, 16'd43892, 16'd22808, 16'd44639, 16'd39954, 16'd9977, 16'd52862, 16'd21610, 16'd28844, 16'd31568, 16'd34244, 16'd53722, 16'd28023, 16'd61551, 16'd38404, 16'd26159, 16'd16304, 16'd10315, 16'd45765, 16'd28000, 16'd15253, 16'd62946, 16'd4083, 16'd5175});
	test_expansion(128'h6c0776db9a53814883add48fcc2f3f40, {16'd14183, 16'd1214, 16'd30435, 16'd17420, 16'd25252, 16'd1320, 16'd14134, 16'd17393, 16'd62429, 16'd44204, 16'd23797, 16'd38403, 16'd7254, 16'd5497, 16'd25210, 16'd7984, 16'd14778, 16'd31176, 16'd46279, 16'd23717, 16'd11293, 16'd52541, 16'd11424, 16'd51088, 16'd59693, 16'd26900});
	test_expansion(128'h9543d8f572ea7ae342b60ec5e017c6a0, {16'd2303, 16'd59997, 16'd52349, 16'd64835, 16'd38195, 16'd59016, 16'd12860, 16'd28468, 16'd21396, 16'd42084, 16'd8707, 16'd35104, 16'd12968, 16'd13453, 16'd27295, 16'd13574, 16'd33055, 16'd16703, 16'd44931, 16'd7815, 16'd62862, 16'd52461, 16'd52056, 16'd41708, 16'd1187, 16'd40094});
	test_expansion(128'ha8d9b8c03e16c001066082c9b3375643, {16'd33788, 16'd27637, 16'd23225, 16'd55320, 16'd10766, 16'd33616, 16'd32669, 16'd31367, 16'd57452, 16'd26629, 16'd27015, 16'd6483, 16'd50074, 16'd39831, 16'd38822, 16'd26753, 16'd64111, 16'd7258, 16'd16443, 16'd42637, 16'd58236, 16'd56016, 16'd35723, 16'd26312, 16'd50915, 16'd64387});
	test_expansion(128'h7c0911ed5a06e5cc95b73564d8f62e63, {16'd38392, 16'd52143, 16'd9006, 16'd58317, 16'd5391, 16'd37897, 16'd35299, 16'd46201, 16'd61531, 16'd33753, 16'd14417, 16'd8278, 16'd18512, 16'd52634, 16'd13179, 16'd42793, 16'd47032, 16'd49862, 16'd47817, 16'd9674, 16'd21103, 16'd31602, 16'd4965, 16'd31938, 16'd37053, 16'd3563});
	test_expansion(128'hc0375e777752e3850a9f6d193bb3bca3, {16'd42921, 16'd63230, 16'd19610, 16'd48613, 16'd28228, 16'd14483, 16'd3548, 16'd38356, 16'd5795, 16'd15596, 16'd11951, 16'd41654, 16'd40933, 16'd5777, 16'd59242, 16'd29940, 16'd11262, 16'd1251, 16'd38812, 16'd23180, 16'd12410, 16'd19993, 16'd31310, 16'd62464, 16'd40792, 16'd30178});
	test_expansion(128'h498ed5243ceb099dbe3a5b379a92ecd0, {16'd20798, 16'd14670, 16'd17647, 16'd11087, 16'd17849, 16'd20348, 16'd23282, 16'd48475, 16'd25897, 16'd38152, 16'd61605, 16'd43284, 16'd3993, 16'd6120, 16'd18266, 16'd25756, 16'd194, 16'd50913, 16'd46959, 16'd11134, 16'd61784, 16'd48847, 16'd14687, 16'd19266, 16'd35589, 16'd56704});
	test_expansion(128'h66a6f0025890c32c7111758f3323c64c, {16'd44733, 16'd64308, 16'd60830, 16'd50441, 16'd45903, 16'd23431, 16'd52097, 16'd43368, 16'd12571, 16'd56971, 16'd29837, 16'd18368, 16'd17090, 16'd41769, 16'd57267, 16'd61945, 16'd30953, 16'd34734, 16'd18670, 16'd13266, 16'd53000, 16'd59779, 16'd9273, 16'd52842, 16'd14170, 16'd38023});
	test_expansion(128'h0dc7dae33c0d44c4187103a271f9aa8b, {16'd17156, 16'd43868, 16'd54942, 16'd3738, 16'd3044, 16'd23979, 16'd43117, 16'd49751, 16'd21126, 16'd48218, 16'd13374, 16'd12168, 16'd19256, 16'd28970, 16'd7571, 16'd1521, 16'd14772, 16'd54945, 16'd58968, 16'd28914, 16'd10062, 16'd43894, 16'd17910, 16'd9790, 16'd26216, 16'd30214});
	test_expansion(128'hd1529f509f99366047c2c557ce27ba6e, {16'd42563, 16'd22632, 16'd54389, 16'd2015, 16'd2592, 16'd1479, 16'd41217, 16'd44201, 16'd31856, 16'd7172, 16'd11007, 16'd3957, 16'd62547, 16'd11023, 16'd14765, 16'd38595, 16'd1351, 16'd27100, 16'd19895, 16'd58251, 16'd9665, 16'd50633, 16'd62553, 16'd41009, 16'd47808, 16'd49038});
	test_expansion(128'hf702ae19880eef70d368596969785459, {16'd30328, 16'd48594, 16'd54530, 16'd49743, 16'd6819, 16'd9964, 16'd60701, 16'd21785, 16'd50470, 16'd39238, 16'd48982, 16'd11738, 16'd57944, 16'd35027, 16'd61193, 16'd33208, 16'd38025, 16'd50154, 16'd29405, 16'd10857, 16'd30839, 16'd29196, 16'd12075, 16'd19384, 16'd60142, 16'd18159});
	test_expansion(128'he1cee51871d352aa7b295cd4e39a50d3, {16'd21664, 16'd7507, 16'd15161, 16'd25785, 16'd16526, 16'd48504, 16'd40447, 16'd29262, 16'd47684, 16'd42792, 16'd26733, 16'd51099, 16'd21910, 16'd51337, 16'd41114, 16'd40658, 16'd3776, 16'd5851, 16'd17630, 16'd4152, 16'd8338, 16'd56611, 16'd39797, 16'd59979, 16'd3026, 16'd30351});
	test_expansion(128'h5d0530986647225ba8644238c2721776, {16'd14858, 16'd58756, 16'd46205, 16'd2003, 16'd35703, 16'd49422, 16'd36563, 16'd21549, 16'd41268, 16'd7902, 16'd16140, 16'd39300, 16'd54989, 16'd7198, 16'd23381, 16'd5504, 16'd62384, 16'd44687, 16'd63419, 16'd23058, 16'd8905, 16'd18416, 16'd45380, 16'd63621, 16'd49618, 16'd11554});
	test_expansion(128'h710eab9fec74141c12d3309e0d14bee6, {16'd54835, 16'd60982, 16'd54723, 16'd42467, 16'd5173, 16'd5569, 16'd22655, 16'd41088, 16'd7892, 16'd43235, 16'd17690, 16'd16172, 16'd59857, 16'd51650, 16'd35949, 16'd12376, 16'd25761, 16'd45846, 16'd29969, 16'd31201, 16'd49817, 16'd25868, 16'd39373, 16'd51079, 16'd31033, 16'd48789});
	test_expansion(128'h79cdddb8d5ee5d067f4389c70e844f38, {16'd20600, 16'd64139, 16'd46703, 16'd33694, 16'd45310, 16'd59987, 16'd38144, 16'd62883, 16'd23657, 16'd41982, 16'd12701, 16'd44455, 16'd44722, 16'd28699, 16'd24678, 16'd30982, 16'd64176, 16'd11163, 16'd25656, 16'd46121, 16'd14366, 16'd43029, 16'd4263, 16'd7307, 16'd20820, 16'd60669});
	test_expansion(128'h4abe0d9492c6f48fb9f0ab2009ffa969, {16'd15487, 16'd14738, 16'd5017, 16'd17812, 16'd40885, 16'd37451, 16'd53094, 16'd5440, 16'd20062, 16'd43597, 16'd50221, 16'd42642, 16'd46628, 16'd46711, 16'd3821, 16'd8939, 16'd58892, 16'd8671, 16'd40403, 16'd31559, 16'd62452, 16'd28663, 16'd25237, 16'd39647, 16'd49934, 16'd25740});
	test_expansion(128'h4afc626c2d64eb28fe53e2a6e5cb0230, {16'd56665, 16'd4548, 16'd49128, 16'd31922, 16'd15219, 16'd60101, 16'd19039, 16'd12560, 16'd41562, 16'd984, 16'd8302, 16'd55318, 16'd30094, 16'd6203, 16'd23009, 16'd23003, 16'd17755, 16'd31697, 16'd46468, 16'd47387, 16'd31924, 16'd64233, 16'd25487, 16'd41569, 16'd29216, 16'd6563});
	test_expansion(128'h486dadc5bd8847f9641264a9add53bf4, {16'd16997, 16'd32454, 16'd60535, 16'd62633, 16'd64820, 16'd7392, 16'd42857, 16'd5477, 16'd11921, 16'd42853, 16'd28688, 16'd19578, 16'd65467, 16'd22048, 16'd16743, 16'd18911, 16'd49898, 16'd23430, 16'd38286, 16'd23008, 16'd23838, 16'd57730, 16'd4381, 16'd48382, 16'd10397, 16'd58399});
	test_expansion(128'heff290b94ca4e4eaecb8738aae5e09a5, {16'd45264, 16'd22218, 16'd51313, 16'd25749, 16'd57921, 16'd45144, 16'd64717, 16'd3290, 16'd54423, 16'd20960, 16'd27466, 16'd27376, 16'd28674, 16'd16693, 16'd26283, 16'd31165, 16'd18166, 16'd61161, 16'd61292, 16'd48147, 16'd26755, 16'd15071, 16'd34541, 16'd48546, 16'd61674, 16'd55684});
	test_expansion(128'he3ccbc5401af410095baf90c745ccdc4, {16'd17423, 16'd28454, 16'd13033, 16'd10451, 16'd6198, 16'd25551, 16'd24169, 16'd23749, 16'd63226, 16'd29037, 16'd4522, 16'd47440, 16'd55973, 16'd46878, 16'd40686, 16'd48463, 16'd44170, 16'd6758, 16'd18228, 16'd34519, 16'd6395, 16'd26612, 16'd28676, 16'd23932, 16'd49905, 16'd63808});
	test_expansion(128'h91955b5a154fe50dce1571338abe4e14, {16'd35019, 16'd32342, 16'd27998, 16'd30480, 16'd61046, 16'd29301, 16'd44405, 16'd27465, 16'd12007, 16'd26554, 16'd59633, 16'd56562, 16'd11758, 16'd30833, 16'd9595, 16'd24636, 16'd41219, 16'd14561, 16'd37799, 16'd53821, 16'd46974, 16'd25259, 16'd24168, 16'd6733, 16'd48683, 16'd26883});
	test_expansion(128'h9ebaf34ddeb179e96ddeb1330af1011a, {16'd62539, 16'd12177, 16'd34805, 16'd62417, 16'd22148, 16'd22456, 16'd35871, 16'd23592, 16'd49185, 16'd37778, 16'd17712, 16'd14449, 16'd35988, 16'd2479, 16'd11870, 16'd20373, 16'd6584, 16'd47191, 16'd52518, 16'd2858, 16'd52803, 16'd30112, 16'd38128, 16'd16889, 16'd16688, 16'd54234});
	test_expansion(128'he7a6dc5ef5120ae8ff38413619327b59, {16'd62188, 16'd13992, 16'd37450, 16'd50910, 16'd60686, 16'd33473, 16'd19102, 16'd13849, 16'd24298, 16'd64037, 16'd55531, 16'd32215, 16'd20369, 16'd42496, 16'd50346, 16'd36408, 16'd4842, 16'd38762, 16'd45041, 16'd21948, 16'd49024, 16'd6905, 16'd52411, 16'd31141, 16'd41945, 16'd48080});
	test_expansion(128'he40c787b80858dd5eb5ddd7b6692628c, {16'd60095, 16'd52218, 16'd6831, 16'd60452, 16'd19325, 16'd8778, 16'd51477, 16'd64100, 16'd5162, 16'd1648, 16'd2343, 16'd47848, 16'd40692, 16'd23562, 16'd47005, 16'd52988, 16'd49103, 16'd20432, 16'd36796, 16'd16156, 16'd24185, 16'd9338, 16'd37036, 16'd56213, 16'd50541, 16'd40393});
	test_expansion(128'h435dc9371979b1bfa0487062b11d2df4, {16'd33276, 16'd4175, 16'd64897, 16'd24875, 16'd6251, 16'd8762, 16'd30754, 16'd20462, 16'd40232, 16'd9374, 16'd53194, 16'd31801, 16'd16058, 16'd17901, 16'd31034, 16'd16190, 16'd2646, 16'd10448, 16'd31677, 16'd62534, 16'd27148, 16'd6603, 16'd5721, 16'd8834, 16'd32916, 16'd253});
	test_expansion(128'h4ccee84ffd42f805e1a4a5f38518c939, {16'd18308, 16'd15148, 16'd40396, 16'd49266, 16'd39489, 16'd29152, 16'd60670, 16'd21539, 16'd18948, 16'd51933, 16'd25659, 16'd49828, 16'd62629, 16'd26657, 16'd9119, 16'd58493, 16'd64921, 16'd45841, 16'd63997, 16'd65024, 16'd55483, 16'd23503, 16'd13813, 16'd20248, 16'd2659, 16'd54735});
	test_expansion(128'he84b5991270cce4dbb8daed925f52ef4, {16'd16857, 16'd61205, 16'd63864, 16'd50269, 16'd55472, 16'd15533, 16'd49975, 16'd36614, 16'd31609, 16'd58674, 16'd40914, 16'd7672, 16'd47667, 16'd54728, 16'd26540, 16'd7950, 16'd60222, 16'd26194, 16'd51707, 16'd61730, 16'd57395, 16'd13434, 16'd34545, 16'd41351, 16'd40166, 16'd26018});
	test_expansion(128'h5edd29d401ae52c6b673fe54ed1dfe9a, {16'd7749, 16'd31263, 16'd27601, 16'd56506, 16'd10040, 16'd17777, 16'd21894, 16'd61963, 16'd37298, 16'd11409, 16'd24062, 16'd63494, 16'd51092, 16'd47607, 16'd14769, 16'd64370, 16'd12711, 16'd7959, 16'd16288, 16'd26455, 16'd57978, 16'd2885, 16'd11896, 16'd30150, 16'd29974, 16'd54284});
	test_expansion(128'h9c2fb07875b9a3a4e9b6bc4c6951f2c2, {16'd26320, 16'd38226, 16'd54327, 16'd21125, 16'd43579, 16'd52359, 16'd52121, 16'd49198, 16'd34165, 16'd43421, 16'd50944, 16'd17135, 16'd13665, 16'd7128, 16'd53979, 16'd47684, 16'd7854, 16'd13458, 16'd49472, 16'd3842, 16'd5147, 16'd36645, 16'd47920, 16'd23759, 16'd63442, 16'd29331});
	test_expansion(128'h27e612fb20dd3c714acd73a5d69a466c, {16'd44304, 16'd18630, 16'd5620, 16'd63477, 16'd43707, 16'd583, 16'd41982, 16'd51095, 16'd38189, 16'd60398, 16'd20029, 16'd55325, 16'd9012, 16'd31018, 16'd3853, 16'd4217, 16'd14761, 16'd25260, 16'd64112, 16'd55894, 16'd42764, 16'd25059, 16'd38557, 16'd17666, 16'd40626, 16'd18586});
	test_expansion(128'h22d1c22ea43f8586f62231f1cc27cf33, {16'd49663, 16'd41637, 16'd3839, 16'd53447, 16'd8586, 16'd43727, 16'd22370, 16'd48448, 16'd39971, 16'd18305, 16'd12852, 16'd32032, 16'd18428, 16'd5821, 16'd25810, 16'd9798, 16'd43157, 16'd34877, 16'd1925, 16'd63364, 16'd48755, 16'd56651, 16'd47076, 16'd38678, 16'd38434, 16'd9443});
	test_expansion(128'h7def3e652a678bf6a4f0e5dcf0a59fcc, {16'd58660, 16'd64734, 16'd54648, 16'd49177, 16'd63733, 16'd46511, 16'd27762, 16'd12509, 16'd15711, 16'd13583, 16'd32524, 16'd41601, 16'd32064, 16'd45957, 16'd51230, 16'd62312, 16'd55319, 16'd39038, 16'd40150, 16'd60944, 16'd36670, 16'd34467, 16'd57832, 16'd57643, 16'd36132, 16'd16891});
	test_expansion(128'h97d74acb7cf1fea6d2deb83ab90c58eb, {16'd35905, 16'd34361, 16'd52110, 16'd9253, 16'd58351, 16'd13168, 16'd64824, 16'd6071, 16'd57766, 16'd40874, 16'd26824, 16'd62814, 16'd53138, 16'd41718, 16'd47937, 16'd36658, 16'd26510, 16'd20609, 16'd46361, 16'd43004, 16'd22475, 16'd40885, 16'd63401, 16'd54362, 16'd42870, 16'd58705});
	test_expansion(128'hc6a6bac2c799003f3c318a691e0f1a6a, {16'd64497, 16'd2469, 16'd64278, 16'd60666, 16'd18600, 16'd33679, 16'd64060, 16'd49235, 16'd3333, 16'd52794, 16'd25404, 16'd18952, 16'd35373, 16'd3017, 16'd3587, 16'd12075, 16'd24594, 16'd8378, 16'd17307, 16'd1669, 16'd43144, 16'd54114, 16'd28777, 16'd47436, 16'd28729, 16'd30541});
	test_expansion(128'hbf103940447ad25dcc0c1b924ae84aed, {16'd31141, 16'd37851, 16'd563, 16'd10984, 16'd49757, 16'd21106, 16'd28315, 16'd25023, 16'd64480, 16'd27759, 16'd15429, 16'd49794, 16'd11555, 16'd32422, 16'd26824, 16'd51011, 16'd37803, 16'd227, 16'd48519, 16'd13862, 16'd11603, 16'd16105, 16'd24204, 16'd618, 16'd4854, 16'd36181});
	test_expansion(128'h673d2b2b45d227c15da01d2ee708201f, {16'd10382, 16'd30018, 16'd43822, 16'd42139, 16'd36355, 16'd36324, 16'd44586, 16'd47964, 16'd43083, 16'd44129, 16'd43747, 16'd55833, 16'd63271, 16'd42282, 16'd58104, 16'd42584, 16'd16690, 16'd32824, 16'd61758, 16'd58669, 16'd60504, 16'd48489, 16'd41722, 16'd40958, 16'd30737, 16'd21527});
	test_expansion(128'he7f2d47bb36e023c4277f2c2c462670b, {16'd11096, 16'd10767, 16'd42732, 16'd19692, 16'd54235, 16'd58711, 16'd18055, 16'd15385, 16'd60847, 16'd49820, 16'd8901, 16'd39578, 16'd64678, 16'd55314, 16'd6608, 16'd48516, 16'd45228, 16'd18520, 16'd19890, 16'd33280, 16'd13364, 16'd15736, 16'd41285, 16'd53355, 16'd59122, 16'd19473});
	test_expansion(128'hc14b03488f78c821bcc21bdab0b8b05f, {16'd59127, 16'd37506, 16'd29636, 16'd44087, 16'd55278, 16'd11531, 16'd51027, 16'd5152, 16'd32285, 16'd58480, 16'd38291, 16'd59934, 16'd63631, 16'd16511, 16'd14870, 16'd40337, 16'd4408, 16'd8284, 16'd40691, 16'd46288, 16'd35790, 16'd13757, 16'd37337, 16'd22052, 16'd41315, 16'd23686});
	test_expansion(128'h997a2c9e41a2f95f368b15e30497d93d, {16'd40213, 16'd29266, 16'd15352, 16'd34068, 16'd36817, 16'd63577, 16'd14561, 16'd20127, 16'd15871, 16'd23365, 16'd20250, 16'd28600, 16'd2428, 16'd489, 16'd5788, 16'd43315, 16'd41048, 16'd16744, 16'd23818, 16'd9633, 16'd61213, 16'd23906, 16'd43928, 16'd32531, 16'd21571, 16'd60442});
	test_expansion(128'hb50be1a19c58bc8bd1f3002c30f92e1b, {16'd931, 16'd37647, 16'd48828, 16'd44177, 16'd14252, 16'd36026, 16'd53389, 16'd23058, 16'd57807, 16'd25766, 16'd961, 16'd9434, 16'd13162, 16'd42797, 16'd15242, 16'd30287, 16'd44813, 16'd23739, 16'd28647, 16'd48610, 16'd9407, 16'd53847, 16'd42210, 16'd37013, 16'd61584, 16'd16225});
	test_expansion(128'hb2986a511513405d87496a7720af07f4, {16'd46608, 16'd21608, 16'd28928, 16'd2466, 16'd61178, 16'd4122, 16'd60655, 16'd16300, 16'd4809, 16'd47544, 16'd41976, 16'd13641, 16'd33295, 16'd22868, 16'd59305, 16'd12777, 16'd40113, 16'd11605, 16'd5222, 16'd10860, 16'd6258, 16'd36671, 16'd14544, 16'd5505, 16'd13338, 16'd14571});
	test_expansion(128'hfb5397fdb62a3e96237a649e8f368394, {16'd38172, 16'd19361, 16'd24957, 16'd37919, 16'd23838, 16'd45750, 16'd28911, 16'd150, 16'd60244, 16'd23530, 16'd22542, 16'd19152, 16'd48641, 16'd48589, 16'd26219, 16'd28709, 16'd47833, 16'd35779, 16'd50691, 16'd53424, 16'd33050, 16'd18377, 16'd43991, 16'd61667, 16'd45169, 16'd36924});
	test_expansion(128'h15b0adc21eb1890373e428be25f4de13, {16'd61827, 16'd22186, 16'd6302, 16'd24740, 16'd29738, 16'd65434, 16'd7236, 16'd43479, 16'd21631, 16'd40567, 16'd34556, 16'd45822, 16'd64632, 16'd54782, 16'd28359, 16'd21553, 16'd11430, 16'd56375, 16'd60383, 16'd54221, 16'd44089, 16'd22797, 16'd36275, 16'd65236, 16'd57935, 16'd58858});
	test_expansion(128'h1652c2138538052a93b9fdd3baec5a4d, {16'd42882, 16'd53780, 16'd9261, 16'd27103, 16'd63159, 16'd14923, 16'd63627, 16'd43256, 16'd1952, 16'd55618, 16'd44964, 16'd40428, 16'd59972, 16'd47607, 16'd63369, 16'd39276, 16'd59034, 16'd35685, 16'd41437, 16'd55749, 16'd22135, 16'd5374, 16'd57900, 16'd13839, 16'd48472, 16'd52059});
	test_expansion(128'h8995a8b757fc66e1ceb38706f12f0311, {16'd26410, 16'd60651, 16'd61891, 16'd21999, 16'd39617, 16'd44296, 16'd8874, 16'd2008, 16'd352, 16'd12180, 16'd43155, 16'd8479, 16'd32309, 16'd60473, 16'd19667, 16'd58432, 16'd48697, 16'd45572, 16'd26438, 16'd56834, 16'd61753, 16'd18722, 16'd42989, 16'd63315, 16'd30453, 16'd19829});
	test_expansion(128'hceef9bdb93760d14ae4d95a3c7ab3d05, {16'd56404, 16'd15701, 16'd49715, 16'd57024, 16'd22702, 16'd25019, 16'd8216, 16'd37923, 16'd61319, 16'd41597, 16'd44013, 16'd24145, 16'd58978, 16'd37350, 16'd32191, 16'd26402, 16'd46393, 16'd38773, 16'd24015, 16'd24833, 16'd9916, 16'd35901, 16'd18182, 16'd9823, 16'd19291, 16'd20977});
	test_expansion(128'h526d3125b2eb3d4ef4c94f4ca0741e1f, {16'd1780, 16'd51529, 16'd3422, 16'd15209, 16'd41375, 16'd29781, 16'd8190, 16'd35541, 16'd8737, 16'd61163, 16'd22645, 16'd47307, 16'd38367, 16'd51495, 16'd8871, 16'd52949, 16'd26040, 16'd47298, 16'd47923, 16'd40242, 16'd2217, 16'd42050, 16'd63555, 16'd13500, 16'd14089, 16'd62182});
	test_expansion(128'h03f2361ed2edff0c0da63bdd7ee2e6c4, {16'd34491, 16'd58342, 16'd1013, 16'd19828, 16'd9535, 16'd26746, 16'd62808, 16'd16370, 16'd5733, 16'd22597, 16'd25673, 16'd16201, 16'd61742, 16'd61339, 16'd21069, 16'd51100, 16'd46965, 16'd3489, 16'd31666, 16'd25331, 16'd50771, 16'd35571, 16'd18363, 16'd41195, 16'd19536, 16'd32016});
	test_expansion(128'h8b3f871b1e38abaa8b30ca4e0caa187b, {16'd8673, 16'd40316, 16'd41761, 16'd50066, 16'd62669, 16'd31628, 16'd48146, 16'd32199, 16'd42516, 16'd24866, 16'd2014, 16'd39626, 16'd20919, 16'd19482, 16'd53173, 16'd51480, 16'd25979, 16'd4143, 16'd48180, 16'd59037, 16'd58366, 16'd46647, 16'd28744, 16'd24545, 16'd50480, 16'd42285});
	test_expansion(128'h8013f0d72882ca393364f5dced26c078, {16'd28768, 16'd63831, 16'd37042, 16'd19251, 16'd29840, 16'd38807, 16'd8084, 16'd41958, 16'd20861, 16'd53103, 16'd17366, 16'd4526, 16'd31335, 16'd738, 16'd65467, 16'd928, 16'd929, 16'd49997, 16'd18443, 16'd47959, 16'd10664, 16'd4204, 16'd27275, 16'd19206, 16'd23922, 16'd50864});
	test_expansion(128'h67fd70e7807de6fa84bc84ae3e92646f, {16'd22230, 16'd47609, 16'd32652, 16'd20446, 16'd52393, 16'd23041, 16'd22265, 16'd41926, 16'd34057, 16'd15338, 16'd20092, 16'd63796, 16'd50319, 16'd40800, 16'd1360, 16'd11015, 16'd47826, 16'd31448, 16'd58275, 16'd59541, 16'd19901, 16'd44580, 16'd54245, 16'd63657, 16'd15061, 16'd12442});
	test_expansion(128'he5653ddb68c8c92c2ad1c4f4e28d1d91, {16'd48675, 16'd17354, 16'd50556, 16'd15780, 16'd57895, 16'd3679, 16'd59884, 16'd63256, 16'd64893, 16'd49053, 16'd57858, 16'd31053, 16'd61769, 16'd21325, 16'd34266, 16'd52343, 16'd40652, 16'd31129, 16'd15756, 16'd57403, 16'd14375, 16'd57252, 16'd38541, 16'd5643, 16'd52804, 16'd21498});
	test_expansion(128'h800a478004abe501941611362cd2db28, {16'd22522, 16'd22720, 16'd60501, 16'd38642, 16'd31844, 16'd25365, 16'd52712, 16'd29126, 16'd30386, 16'd26931, 16'd60649, 16'd60116, 16'd52555, 16'd45217, 16'd37420, 16'd14374, 16'd46588, 16'd53578, 16'd19697, 16'd40912, 16'd49861, 16'd60268, 16'd44829, 16'd2415, 16'd3537, 16'd59762});
	test_expansion(128'h41f3de0950c1778194b17cc3466818b9, {16'd32714, 16'd19065, 16'd64439, 16'd51931, 16'd46190, 16'd5635, 16'd58422, 16'd60433, 16'd33447, 16'd65308, 16'd59327, 16'd39005, 16'd4581, 16'd30423, 16'd31445, 16'd51742, 16'd60279, 16'd15115, 16'd25221, 16'd23511, 16'd48890, 16'd15950, 16'd37631, 16'd14099, 16'd41927, 16'd63512});
	test_expansion(128'h06750c71e943cabf0282253c76da5c82, {16'd61004, 16'd61066, 16'd1388, 16'd60276, 16'd5832, 16'd35078, 16'd19266, 16'd40977, 16'd17215, 16'd34408, 16'd21948, 16'd35903, 16'd43149, 16'd33171, 16'd35584, 16'd1563, 16'd44242, 16'd16846, 16'd16517, 16'd34676, 16'd10351, 16'd36983, 16'd53468, 16'd58796, 16'd15174, 16'd35834});
	test_expansion(128'h3b9b6cadf15a79010c526bc82407b998, {16'd34444, 16'd35606, 16'd20948, 16'd54009, 16'd3742, 16'd4813, 16'd40854, 16'd5508, 16'd58459, 16'd8992, 16'd64278, 16'd22113, 16'd26034, 16'd36138, 16'd53613, 16'd64433, 16'd45688, 16'd11330, 16'd41961, 16'd2452, 16'd61726, 16'd23400, 16'd25123, 16'd54075, 16'd58834, 16'd4713});
	test_expansion(128'hc86bf96bc8e6440829e9be58115462da, {16'd38417, 16'd64815, 16'd44299, 16'd10489, 16'd15482, 16'd23670, 16'd40443, 16'd42843, 16'd34545, 16'd37508, 16'd22915, 16'd37341, 16'd19949, 16'd18468, 16'd10022, 16'd43020, 16'd48080, 16'd23634, 16'd57290, 16'd5518, 16'd63245, 16'd55255, 16'd45748, 16'd36043, 16'd59628, 16'd56960});
	test_expansion(128'hfc9c09c07a6c5b0bedf12f2991996a5e, {16'd13359, 16'd58325, 16'd34051, 16'd64455, 16'd25247, 16'd55674, 16'd27831, 16'd31795, 16'd26781, 16'd45272, 16'd29525, 16'd51485, 16'd62353, 16'd65429, 16'd55140, 16'd10794, 16'd27974, 16'd18905, 16'd7042, 16'd59196, 16'd27124, 16'd57746, 16'd5409, 16'd24907, 16'd6775, 16'd43426});
	test_expansion(128'h5cf30abf8b0578cbb2e7268ec9157e47, {16'd49490, 16'd39841, 16'd8399, 16'd48112, 16'd54589, 16'd50648, 16'd36028, 16'd39552, 16'd26234, 16'd45577, 16'd43696, 16'd6204, 16'd65043, 16'd7748, 16'd47167, 16'd45634, 16'd12971, 16'd61368, 16'd39681, 16'd19168, 16'd55798, 16'd34876, 16'd40693, 16'd14990, 16'd50318, 16'd23930});
	test_expansion(128'h241a68d5c163cd4d9f448773ce2b0b81, {16'd32926, 16'd2751, 16'd43245, 16'd8316, 16'd352, 16'd60818, 16'd17066, 16'd10909, 16'd990, 16'd46338, 16'd49505, 16'd8657, 16'd19750, 16'd39247, 16'd35632, 16'd8542, 16'd32376, 16'd25694, 16'd1326, 16'd63403, 16'd2544, 16'd4008, 16'd60745, 16'd24830, 16'd51835, 16'd2484});
	test_expansion(128'h84e68e6fb7184a57c7460eedfe6f3d5d, {16'd14887, 16'd147, 16'd61082, 16'd56152, 16'd51152, 16'd28756, 16'd59010, 16'd57838, 16'd38715, 16'd24338, 16'd24627, 16'd24089, 16'd41607, 16'd10439, 16'd36884, 16'd29758, 16'd9586, 16'd64790, 16'd36609, 16'd18334, 16'd3833, 16'd8940, 16'd19731, 16'd10572, 16'd2934, 16'd59390});
	test_expansion(128'h324579ee6d80cfe52dc4d3e18ba48d3d, {16'd15090, 16'd24198, 16'd13466, 16'd37746, 16'd31358, 16'd62702, 16'd29781, 16'd21467, 16'd10002, 16'd18664, 16'd59168, 16'd26340, 16'd1660, 16'd20121, 16'd52730, 16'd37813, 16'd30444, 16'd37053, 16'd48836, 16'd50818, 16'd34419, 16'd61479, 16'd259, 16'd56475, 16'd10745, 16'd40284});
	test_expansion(128'hdd65207c4c8093edfe54d04eeb8193a4, {16'd49497, 16'd43856, 16'd48476, 16'd10201, 16'd57099, 16'd35223, 16'd25254, 16'd1354, 16'd426, 16'd50283, 16'd61256, 16'd13171, 16'd54990, 16'd39625, 16'd56029, 16'd54142, 16'd42215, 16'd20739, 16'd8719, 16'd64074, 16'd19154, 16'd29933, 16'd41477, 16'd10679, 16'd44523, 16'd57415});
	test_expansion(128'h967574ecf2b49ac92d34b63e86259dd5, {16'd59197, 16'd4397, 16'd21533, 16'd53366, 16'd19156, 16'd60340, 16'd37075, 16'd4629, 16'd19117, 16'd52162, 16'd37414, 16'd54760, 16'd60611, 16'd35209, 16'd15377, 16'd40891, 16'd2537, 16'd51469, 16'd21859, 16'd16945, 16'd61348, 16'd28955, 16'd46654, 16'd28542, 16'd39897, 16'd19911});
	test_expansion(128'h304f97cee8cfe7da05fecc0c647e2565, {16'd4708, 16'd6341, 16'd39730, 16'd6743, 16'd31051, 16'd53110, 16'd22535, 16'd65379, 16'd61323, 16'd14207, 16'd65508, 16'd26720, 16'd58240, 16'd5608, 16'd46282, 16'd32448, 16'd42545, 16'd55108, 16'd10201, 16'd26915, 16'd23189, 16'd394, 16'd28546, 16'd21520, 16'd57134, 16'd28139});
	test_expansion(128'h6278c1f908f649a0d1994123d35d0acd, {16'd13654, 16'd32061, 16'd50265, 16'd17120, 16'd24886, 16'd46146, 16'd2161, 16'd51710, 16'd10343, 16'd26700, 16'd58813, 16'd53768, 16'd13772, 16'd61498, 16'd58661, 16'd34638, 16'd24737, 16'd11851, 16'd32319, 16'd25105, 16'd37846, 16'd57998, 16'd64806, 16'd63430, 16'd20097, 16'd27903});
	test_expansion(128'h7b36e57f0a762c1b809b87b6e79c0a1f, {16'd29875, 16'd28580, 16'd8996, 16'd4359, 16'd9636, 16'd62980, 16'd62689, 16'd49617, 16'd58721, 16'd37222, 16'd44889, 16'd5508, 16'd47870, 16'd10251, 16'd3337, 16'd3037, 16'd19577, 16'd10018, 16'd63271, 16'd22602, 16'd54701, 16'd3414, 16'd2621, 16'd47423, 16'd49268, 16'd27132});
	test_expansion(128'hb9da1172f740c25a65ebc73c117eeb82, {16'd62803, 16'd517, 16'd20597, 16'd4567, 16'd48516, 16'd22500, 16'd26386, 16'd3585, 16'd15701, 16'd38409, 16'd929, 16'd38087, 16'd20335, 16'd60468, 16'd33696, 16'd52903, 16'd23919, 16'd52042, 16'd59629, 16'd6711, 16'd33558, 16'd12757, 16'd54136, 16'd23700, 16'd19190, 16'd63090});
	test_expansion(128'hbe32b79e0f8f2d26158903900cc3ceee, {16'd57353, 16'd44731, 16'd13316, 16'd57421, 16'd3603, 16'd5400, 16'd6573, 16'd42331, 16'd15925, 16'd40866, 16'd54955, 16'd56101, 16'd6107, 16'd5637, 16'd24958, 16'd44905, 16'd20753, 16'd34794, 16'd4587, 16'd48850, 16'd38128, 16'd40992, 16'd58741, 16'd2410, 16'd30658, 16'd30118});
	test_expansion(128'h88fd86573cfc801459d8f059f0ed20ff, {16'd50591, 16'd18405, 16'd5418, 16'd27433, 16'd15941, 16'd33041, 16'd8834, 16'd63159, 16'd28457, 16'd45911, 16'd48065, 16'd40336, 16'd60555, 16'd61367, 16'd18248, 16'd46068, 16'd65335, 16'd11931, 16'd37782, 16'd19206, 16'd62546, 16'd22159, 16'd49640, 16'd12128, 16'd18014, 16'd6161});
	test_expansion(128'h5bd26c7b80d2b502f9bac513c9f52c04, {16'd8973, 16'd48058, 16'd23841, 16'd64559, 16'd21674, 16'd55208, 16'd21886, 16'd31225, 16'd56961, 16'd38107, 16'd22491, 16'd62251, 16'd43998, 16'd51966, 16'd26637, 16'd17303, 16'd17490, 16'd62176, 16'd2736, 16'd55811, 16'd22722, 16'd19233, 16'd9830, 16'd65383, 16'd23708, 16'd24100});
	test_expansion(128'h0f446a4d06f470d6c8d9e7af4c7901de, {16'd21411, 16'd49521, 16'd53456, 16'd62476, 16'd54548, 16'd309, 16'd35067, 16'd3450, 16'd35862, 16'd48122, 16'd54364, 16'd3355, 16'd11612, 16'd38776, 16'd21535, 16'd13595, 16'd15274, 16'd618, 16'd35053, 16'd42762, 16'd28762, 16'd24103, 16'd43846, 16'd46014, 16'd24440, 16'd41233});
	test_expansion(128'h5ad275fb301bae6d01365d2f1d9d57df, {16'd42648, 16'd19540, 16'd607, 16'd40203, 16'd15225, 16'd58590, 16'd41559, 16'd46742, 16'd49268, 16'd43234, 16'd30226, 16'd51001, 16'd19063, 16'd56006, 16'd36553, 16'd8943, 16'd7704, 16'd5847, 16'd35111, 16'd8722, 16'd11034, 16'd11974, 16'd26845, 16'd14865, 16'd56681, 16'd27573});
	test_expansion(128'hed5e897ee946b7a4cd8be2bb9b94230f, {16'd44711, 16'd47489, 16'd17960, 16'd52782, 16'd47108, 16'd48153, 16'd5192, 16'd42680, 16'd31940, 16'd47587, 16'd22857, 16'd52481, 16'd45969, 16'd11004, 16'd46970, 16'd6260, 16'd59128, 16'd43150, 16'd62735, 16'd28150, 16'd56669, 16'd23469, 16'd13649, 16'd26124, 16'd46103, 16'd35482});
	test_expansion(128'h64989944be2685bdbe34db1e9b882a92, {16'd4225, 16'd33854, 16'd10817, 16'd30071, 16'd21487, 16'd51368, 16'd36849, 16'd9948, 16'd1649, 16'd64197, 16'd23521, 16'd24467, 16'd38613, 16'd45882, 16'd48820, 16'd21832, 16'd4282, 16'd43725, 16'd51758, 16'd39708, 16'd26358, 16'd20584, 16'd41848, 16'd22894, 16'd15348, 16'd25456});
	test_expansion(128'h0b23174e422c6ddc790c0a1add6d38c5, {16'd40059, 16'd17333, 16'd39246, 16'd46623, 16'd52878, 16'd351, 16'd13305, 16'd42977, 16'd2270, 16'd7580, 16'd27980, 16'd25862, 16'd36497, 16'd38833, 16'd38461, 16'd58447, 16'd26028, 16'd35269, 16'd61098, 16'd56720, 16'd52729, 16'd41423, 16'd39234, 16'd37408, 16'd45855, 16'd58625});
	test_expansion(128'h0006fe872a5e10a1349f33880eed9b07, {16'd29606, 16'd48406, 16'd22076, 16'd10844, 16'd8218, 16'd55111, 16'd17520, 16'd19697, 16'd16612, 16'd46126, 16'd41247, 16'd12974, 16'd18306, 16'd59421, 16'd42869, 16'd38022, 16'd32432, 16'd30597, 16'd5787, 16'd12397, 16'd3419, 16'd46753, 16'd12314, 16'd32293, 16'd7311, 16'd11766});
	test_expansion(128'hb883116db25603984b69dcd5cdd80b1b, {16'd14400, 16'd292, 16'd40607, 16'd55815, 16'd23864, 16'd28597, 16'd57272, 16'd4048, 16'd13470, 16'd39126, 16'd37955, 16'd54677, 16'd33304, 16'd53286, 16'd11963, 16'd63604, 16'd45078, 16'd35151, 16'd16340, 16'd61702, 16'd38006, 16'd11830, 16'd11090, 16'd49493, 16'd43620, 16'd61546});
	test_expansion(128'h4aa613939ddb24ceeb36f3ed4d8c1a10, {16'd57977, 16'd12844, 16'd34132, 16'd28382, 16'd62305, 16'd6770, 16'd14809, 16'd44996, 16'd36067, 16'd18211, 16'd11225, 16'd64872, 16'd46828, 16'd14873, 16'd58289, 16'd33209, 16'd46114, 16'd601, 16'd60492, 16'd34722, 16'd60419, 16'd57925, 16'd7211, 16'd30139, 16'd31815, 16'd47779});
	test_expansion(128'h7a44864d3906eca46b8a71d75e5a17fe, {16'd42840, 16'd64565, 16'd15671, 16'd13512, 16'd5897, 16'd47593, 16'd14206, 16'd64803, 16'd11987, 16'd60140, 16'd6116, 16'd19404, 16'd30819, 16'd21156, 16'd46943, 16'd40982, 16'd22109, 16'd44131, 16'd41388, 16'd30871, 16'd35260, 16'd38949, 16'd53457, 16'd51348, 16'd8130, 16'd62289});
	test_expansion(128'h30d9fe4f88e9cdb3254a6c31fbf615b7, {16'd47587, 16'd45594, 16'd20160, 16'd16412, 16'd38628, 16'd46322, 16'd35592, 16'd35790, 16'd1290, 16'd12001, 16'd52457, 16'd47532, 16'd37952, 16'd6103, 16'd39504, 16'd45301, 16'd40302, 16'd36196, 16'd39080, 16'd40329, 16'd1070, 16'd51667, 16'd41055, 16'd11058, 16'd2283, 16'd35683});
	test_expansion(128'hebe43a74ee58dc5a7e1990cfa5ae8091, {16'd56071, 16'd11495, 16'd52977, 16'd7978, 16'd50335, 16'd11655, 16'd45712, 16'd17706, 16'd53813, 16'd27452, 16'd48484, 16'd31332, 16'd43336, 16'd44210, 16'd37586, 16'd25313, 16'd18775, 16'd41616, 16'd19901, 16'd11356, 16'd11908, 16'd10062, 16'd63424, 16'd54127, 16'd29361, 16'd7521});
	test_expansion(128'h833b1807e4874bca27a256688477e616, {16'd33782, 16'd49352, 16'd48662, 16'd49806, 16'd47072, 16'd59894, 16'd9150, 16'd28886, 16'd14223, 16'd42147, 16'd49970, 16'd62615, 16'd59497, 16'd22540, 16'd24403, 16'd52930, 16'd26778, 16'd25968, 16'd856, 16'd61233, 16'd8993, 16'd38727, 16'd37230, 16'd37702, 16'd10190, 16'd8496});
	test_expansion(128'haea1f5f751617f9820a7f17046e9770e, {16'd42235, 16'd27979, 16'd22632, 16'd48816, 16'd58798, 16'd2304, 16'd38015, 16'd53315, 16'd33910, 16'd54858, 16'd63280, 16'd62023, 16'd12877, 16'd7271, 16'd18663, 16'd26127, 16'd55119, 16'd18737, 16'd32593, 16'd6001, 16'd11431, 16'd41825, 16'd14989, 16'd40864, 16'd36284, 16'd24641});
	test_expansion(128'h783f5b6444754ba1487ea21034d31f60, {16'd1167, 16'd48825, 16'd64556, 16'd20315, 16'd40763, 16'd56249, 16'd44988, 16'd14004, 16'd61602, 16'd33505, 16'd6039, 16'd3322, 16'd14964, 16'd30588, 16'd38490, 16'd5651, 16'd3358, 16'd30891, 16'd6788, 16'd25892, 16'd6765, 16'd12671, 16'd59139, 16'd6115, 16'd11839, 16'd63090});
	test_expansion(128'hbf689e615e1ebee5527022bca5739fe7, {16'd24060, 16'd18116, 16'd38215, 16'd36529, 16'd18980, 16'd56355, 16'd1637, 16'd18149, 16'd50869, 16'd59607, 16'd23729, 16'd55947, 16'd7552, 16'd6519, 16'd9537, 16'd54291, 16'd33161, 16'd15456, 16'd20513, 16'd45834, 16'd31796, 16'd1589, 16'd49002, 16'd43465, 16'd29314, 16'd1713});
	test_expansion(128'h4b14635f4440f6d0af581abd6fd343fa, {16'd14587, 16'd24710, 16'd57676, 16'd5517, 16'd59834, 16'd18961, 16'd52430, 16'd18509, 16'd18914, 16'd32764, 16'd12079, 16'd56161, 16'd50558, 16'd17013, 16'd62250, 16'd16323, 16'd3290, 16'd27269, 16'd36837, 16'd65403, 16'd38336, 16'd60417, 16'd46723, 16'd53219, 16'd45069, 16'd11719});
	test_expansion(128'h27968a6d6f19a276dbd58502cc9b1d55, {16'd25051, 16'd13389, 16'd35665, 16'd49786, 16'd38599, 16'd38904, 16'd16829, 16'd39790, 16'd18684, 16'd50554, 16'd16387, 16'd29211, 16'd21758, 16'd61365, 16'd63797, 16'd5027, 16'd2730, 16'd12175, 16'd41021, 16'd7193, 16'd29080, 16'd7743, 16'd19131, 16'd62686, 16'd65089, 16'd55090});
	test_expansion(128'hb40d4183de82c0dfe96bd80e35b8aa97, {16'd34030, 16'd13696, 16'd7808, 16'd47917, 16'd41141, 16'd9364, 16'd59275, 16'd47259, 16'd3096, 16'd34517, 16'd55720, 16'd54627, 16'd20201, 16'd15484, 16'd21102, 16'd48272, 16'd42676, 16'd31011, 16'd25454, 16'd17844, 16'd9392, 16'd61917, 16'd18488, 16'd9555, 16'd34204, 16'd51694});
	test_expansion(128'hee90864a7606dd827300e76c3636f597, {16'd44758, 16'd15078, 16'd6267, 16'd29351, 16'd18312, 16'd35812, 16'd50526, 16'd55030, 16'd58472, 16'd21919, 16'd26992, 16'd42527, 16'd15181, 16'd7149, 16'd8124, 16'd26896, 16'd16089, 16'd475, 16'd12146, 16'd32822, 16'd39300, 16'd19269, 16'd14077, 16'd17173, 16'd25950, 16'd7535});
	test_expansion(128'hb57df22c273603ad1571d55d0b81e89b, {16'd35680, 16'd30801, 16'd10325, 16'd57690, 16'd39696, 16'd46912, 16'd36122, 16'd42302, 16'd63418, 16'd65449, 16'd36146, 16'd14322, 16'd61389, 16'd26139, 16'd7896, 16'd19792, 16'd58537, 16'd26647, 16'd2336, 16'd11488, 16'd47075, 16'd63677, 16'd46264, 16'd18845, 16'd6050, 16'd17094});
	test_expansion(128'hdca040be5b0af644e503bfe2f67b9be5, {16'd8737, 16'd40252, 16'd62393, 16'd8941, 16'd9219, 16'd20863, 16'd29587, 16'd13086, 16'd26422, 16'd32437, 16'd7698, 16'd28320, 16'd12382, 16'd13524, 16'd17213, 16'd6897, 16'd58930, 16'd46508, 16'd42806, 16'd22984, 16'd62256, 16'd21463, 16'd48507, 16'd31083, 16'd51250, 16'd22800});
	test_expansion(128'h17cd85f9aa1edd757a1613631fc16751, {16'd8375, 16'd31921, 16'd64260, 16'd24437, 16'd14726, 16'd34976, 16'd51771, 16'd43689, 16'd8583, 16'd53964, 16'd43125, 16'd7141, 16'd1035, 16'd6018, 16'd45112, 16'd21463, 16'd19803, 16'd25495, 16'd50928, 16'd43117, 16'd45763, 16'd35801, 16'd37039, 16'd14720, 16'd18303, 16'd6106});
	test_expansion(128'h7c7edbd0f8f003719741f09b63a50a2b, {16'd62369, 16'd12409, 16'd13999, 16'd21266, 16'd41259, 16'd33064, 16'd52511, 16'd30823, 16'd65031, 16'd25546, 16'd59102, 16'd56464, 16'd29918, 16'd60883, 16'd35358, 16'd34793, 16'd43609, 16'd60529, 16'd57502, 16'd12634, 16'd54390, 16'd37307, 16'd6888, 16'd3966, 16'd38150, 16'd19694});
	test_expansion(128'hd09f1b808a0db909fd017ee83ff0e7e2, {16'd35095, 16'd27154, 16'd33648, 16'd24094, 16'd40589, 16'd19458, 16'd18831, 16'd49183, 16'd23634, 16'd29210, 16'd4294, 16'd24529, 16'd31481, 16'd21672, 16'd37203, 16'd21094, 16'd50280, 16'd11009, 16'd14449, 16'd57440, 16'd25237, 16'd46168, 16'd19792, 16'd3481, 16'd64933, 16'd63711});
	test_expansion(128'h1752853b8a10fd14b1a800cf566e43e3, {16'd3795, 16'd28635, 16'd13631, 16'd38085, 16'd48160, 16'd33037, 16'd44757, 16'd33988, 16'd5098, 16'd40700, 16'd9848, 16'd39285, 16'd54641, 16'd21516, 16'd11047, 16'd1334, 16'd8712, 16'd15011, 16'd25176, 16'd54510, 16'd10501, 16'd51397, 16'd27959, 16'd51327, 16'd46055, 16'd50334});
	test_expansion(128'h100601035ff14d8b837368f394eb7546, {16'd15940, 16'd2785, 16'd64215, 16'd57373, 16'd19248, 16'd9796, 16'd36415, 16'd5875, 16'd47131, 16'd5408, 16'd14218, 16'd25611, 16'd17413, 16'd24257, 16'd27193, 16'd58443, 16'd36296, 16'd52445, 16'd886, 16'd48019, 16'd11556, 16'd41921, 16'd24979, 16'd46059, 16'd13656, 16'd13167});
	test_expansion(128'h4a02fd078b5e7e1b03658055cc014d5e, {16'd36150, 16'd48640, 16'd4939, 16'd63201, 16'd43899, 16'd39089, 16'd25849, 16'd42675, 16'd6977, 16'd10082, 16'd221, 16'd60016, 16'd25560, 16'd45686, 16'd5166, 16'd58729, 16'd43820, 16'd48759, 16'd365, 16'd63619, 16'd17303, 16'd16096, 16'd17097, 16'd6610, 16'd62105, 16'd20921});
	test_expansion(128'h9b7a79248b6c39eb92a77540b3367b4e, {16'd34418, 16'd41914, 16'd12491, 16'd2670, 16'd63390, 16'd53447, 16'd62163, 16'd44082, 16'd32930, 16'd62535, 16'd22137, 16'd23809, 16'd39433, 16'd14627, 16'd6843, 16'd18251, 16'd59493, 16'd18984, 16'd12623, 16'd45242, 16'd4377, 16'd28742, 16'd998, 16'd49649, 16'd14897, 16'd24773});
	test_expansion(128'h839aa51afa82d4cf7172035866e0fb95, {16'd28770, 16'd59311, 16'd8152, 16'd54583, 16'd18586, 16'd40738, 16'd27630, 16'd18221, 16'd22952, 16'd55871, 16'd47793, 16'd50207, 16'd55388, 16'd43367, 16'd28978, 16'd56187, 16'd48577, 16'd65319, 16'd27027, 16'd15636, 16'd54995, 16'd59757, 16'd39406, 16'd6779, 16'd3081, 16'd1039});
	test_expansion(128'he777e7c7bffb309f9e6be884325dc1d3, {16'd32088, 16'd36502, 16'd37266, 16'd18576, 16'd36086, 16'd30395, 16'd10369, 16'd5126, 16'd36857, 16'd32573, 16'd51231, 16'd25864, 16'd26594, 16'd8693, 16'd52878, 16'd47844, 16'd21140, 16'd28097, 16'd3175, 16'd46952, 16'd45162, 16'd57719, 16'd11263, 16'd32562, 16'd10852, 16'd4149});
	test_expansion(128'h5f8ef0c811ad2204ea7cbb0b5bc48236, {16'd17203, 16'd50069, 16'd36502, 16'd40079, 16'd9302, 16'd36350, 16'd22223, 16'd37641, 16'd56390, 16'd12001, 16'd37354, 16'd32715, 16'd14496, 16'd37357, 16'd27667, 16'd49492, 16'd18877, 16'd1152, 16'd17617, 16'd58997, 16'd24364, 16'd22354, 16'd36562, 16'd41312, 16'd38593, 16'd24850});
	test_expansion(128'he53eb6c1a213f69bc6ebc724c47636a7, {16'd63026, 16'd61334, 16'd31617, 16'd33740, 16'd62517, 16'd24289, 16'd5915, 16'd11750, 16'd38909, 16'd17492, 16'd5532, 16'd45955, 16'd26876, 16'd41996, 16'd50223, 16'd1207, 16'd63134, 16'd9684, 16'd22559, 16'd3733, 16'd9943, 16'd25704, 16'd28477, 16'd41215, 16'd63093, 16'd62211});
	test_expansion(128'h67d47b80f0dc3a810a2b971e8852dd9c, {16'd64253, 16'd11553, 16'd20771, 16'd14581, 16'd46275, 16'd34538, 16'd4108, 16'd12378, 16'd21059, 16'd46194, 16'd11195, 16'd5668, 16'd53154, 16'd53674, 16'd62711, 16'd44007, 16'd28406, 16'd54485, 16'd32237, 16'd26782, 16'd24485, 16'd64254, 16'd6987, 16'd10931, 16'd22111, 16'd65338});
	test_expansion(128'he7b74ea0232353d351d705ee2bbd5b84, {16'd4139, 16'd44439, 16'd18804, 16'd20449, 16'd31255, 16'd26715, 16'd40643, 16'd25542, 16'd22944, 16'd34492, 16'd36841, 16'd28669, 16'd60233, 16'd13551, 16'd49057, 16'd47904, 16'd15195, 16'd37092, 16'd18813, 16'd52066, 16'd50946, 16'd24854, 16'd20444, 16'd10545, 16'd9864, 16'd53169});
	test_expansion(128'ha3d0dc79ebae6ccfeb6aae7bdfc9b3e1, {16'd36400, 16'd25480, 16'd28715, 16'd15388, 16'd26687, 16'd4775, 16'd53384, 16'd39706, 16'd34967, 16'd21254, 16'd22180, 16'd58752, 16'd4351, 16'd9475, 16'd38236, 16'd44340, 16'd34632, 16'd8055, 16'd61863, 16'd43174, 16'd18299, 16'd64869, 16'd62530, 16'd60205, 16'd30610, 16'd42224});
	test_expansion(128'hcfbdd98f3a69870290cce7219d8ff0a3, {16'd23460, 16'd41503, 16'd1639, 16'd53048, 16'd54631, 16'd34401, 16'd46384, 16'd23460, 16'd49759, 16'd3395, 16'd4811, 16'd45536, 16'd29865, 16'd43392, 16'd12798, 16'd19374, 16'd9775, 16'd16960, 16'd48875, 16'd56480, 16'd1696, 16'd64525, 16'd44298, 16'd996, 16'd51522, 16'd62428});
	test_expansion(128'hbd1c0b07fdab0c0243681725296c1dd4, {16'd31684, 16'd3940, 16'd19574, 16'd33935, 16'd38323, 16'd62737, 16'd34653, 16'd49904, 16'd56523, 16'd46711, 16'd32311, 16'd53302, 16'd27375, 16'd35474, 16'd31101, 16'd53339, 16'd15273, 16'd49156, 16'd52895, 16'd45187, 16'd48757, 16'd42156, 16'd43211, 16'd25290, 16'd26853, 16'd12284});
	test_expansion(128'hbbfac3d926df6a51aa70517073f7042b, {16'd36667, 16'd42819, 16'd33673, 16'd45520, 16'd11529, 16'd52260, 16'd20152, 16'd56776, 16'd49360, 16'd27473, 16'd22935, 16'd39218, 16'd17629, 16'd61024, 16'd24726, 16'd44756, 16'd55137, 16'd46747, 16'd41055, 16'd40753, 16'd9435, 16'd55135, 16'd16120, 16'd42994, 16'd45484, 16'd62914});
	test_expansion(128'hd257b2c426fb13ce8ced9897aff5ab29, {16'd55536, 16'd21015, 16'd45571, 16'd41322, 16'd61580, 16'd63065, 16'd30253, 16'd42016, 16'd42942, 16'd13236, 16'd23830, 16'd51854, 16'd58831, 16'd29356, 16'd47276, 16'd25192, 16'd51403, 16'd14333, 16'd4297, 16'd51474, 16'd34270, 16'd26536, 16'd54356, 16'd27454, 16'd2350, 16'd37617});
	test_expansion(128'h0878a2040289313b706c3ea8a734fc51, {16'd52118, 16'd15420, 16'd35072, 16'd32307, 16'd7493, 16'd61420, 16'd6278, 16'd7494, 16'd55199, 16'd28299, 16'd10392, 16'd38660, 16'd2047, 16'd28557, 16'd49257, 16'd29390, 16'd24189, 16'd30429, 16'd36395, 16'd62661, 16'd61909, 16'd36705, 16'd45733, 16'd10961, 16'd51410, 16'd42577});
	test_expansion(128'hcb95c1b3f0b32bcabb5d762da519d4b4, {16'd64637, 16'd20344, 16'd8935, 16'd38426, 16'd38131, 16'd39761, 16'd38223, 16'd33609, 16'd56880, 16'd27598, 16'd20064, 16'd31093, 16'd27937, 16'd24725, 16'd30143, 16'd28405, 16'd39682, 16'd42308, 16'd62791, 16'd65250, 16'd24445, 16'd58848, 16'd42490, 16'd52248, 16'd52519, 16'd15587});
	test_expansion(128'h7df43ae5bae4621163ef97b0d5b8d93a, {16'd11751, 16'd24470, 16'd43357, 16'd60308, 16'd5224, 16'd34616, 16'd23656, 16'd65111, 16'd26755, 16'd52129, 16'd25124, 16'd31532, 16'd57007, 16'd27748, 16'd21236, 16'd52167, 16'd6692, 16'd2295, 16'd15169, 16'd27360, 16'd61308, 16'd52041, 16'd28315, 16'd27641, 16'd54928, 16'd8144});
	test_expansion(128'hc20fd75fca3fbcb466b5d02b750dc835, {16'd63003, 16'd25951, 16'd34083, 16'd36380, 16'd45023, 16'd45637, 16'd51802, 16'd37626, 16'd54899, 16'd34886, 16'd34425, 16'd52935, 16'd7279, 16'd11852, 16'd23478, 16'd38583, 16'd24059, 16'd35115, 16'd42435, 16'd52199, 16'd46626, 16'd33076, 16'd44913, 16'd38244, 16'd17130, 16'd49413});
	test_expansion(128'ha72183d828dd7b05b6d426dfd94053a1, {16'd11844, 16'd21963, 16'd51870, 16'd20674, 16'd1780, 16'd10545, 16'd17531, 16'd32868, 16'd43262, 16'd29083, 16'd7387, 16'd59740, 16'd26082, 16'd25290, 16'd32269, 16'd29085, 16'd26000, 16'd12876, 16'd30278, 16'd11884, 16'd52728, 16'd55932, 16'd2789, 16'd27994, 16'd4915, 16'd13028});
	test_expansion(128'hca43242ec258221ce099838e7ab20784, {16'd39967, 16'd22715, 16'd41142, 16'd7220, 16'd32919, 16'd2241, 16'd58080, 16'd9695, 16'd51621, 16'd53605, 16'd30860, 16'd24911, 16'd37555, 16'd43019, 16'd13887, 16'd10542, 16'd5589, 16'd46232, 16'd23966, 16'd62049, 16'd9827, 16'd11848, 16'd24996, 16'd13249, 16'd44159, 16'd57085});
	test_expansion(128'h28c0f07a2cfbdc78b46f86905a451248, {16'd46170, 16'd10967, 16'd12364, 16'd15400, 16'd31744, 16'd788, 16'd19204, 16'd33169, 16'd28950, 16'd55361, 16'd59097, 16'd29647, 16'd15674, 16'd8776, 16'd19368, 16'd6964, 16'd22124, 16'd35143, 16'd47485, 16'd47944, 16'd55961, 16'd46393, 16'd19915, 16'd17773, 16'd42858, 16'd54886});
	test_expansion(128'h1c502fbff5b18eb93635100441e092f6, {16'd46961, 16'd58692, 16'd45640, 16'd47326, 16'd62169, 16'd21171, 16'd60519, 16'd54621, 16'd30084, 16'd4476, 16'd32145, 16'd37739, 16'd17564, 16'd17842, 16'd12140, 16'd3426, 16'd44320, 16'd24457, 16'd62696, 16'd36285, 16'd61839, 16'd24137, 16'd32072, 16'd19287, 16'd1832, 16'd41153});
	test_expansion(128'hca26dfed932633ae1d651c1ffcb0130c, {16'd7649, 16'd46020, 16'd3427, 16'd49222, 16'd16818, 16'd16309, 16'd12664, 16'd47809, 16'd18770, 16'd6783, 16'd30996, 16'd52649, 16'd10812, 16'd35275, 16'd30722, 16'd20801, 16'd19530, 16'd18470, 16'd25486, 16'd15773, 16'd55541, 16'd53038, 16'd32597, 16'd9342, 16'd16386, 16'd53556});
	test_expansion(128'h94bd694396fc17e4e594b1f7f657bb21, {16'd5082, 16'd65277, 16'd31567, 16'd10487, 16'd34998, 16'd42379, 16'd63558, 16'd5719, 16'd16425, 16'd651, 16'd9769, 16'd8018, 16'd1545, 16'd36830, 16'd59814, 16'd10306, 16'd47487, 16'd50265, 16'd25313, 16'd51692, 16'd59937, 16'd23967, 16'd2334, 16'd37244, 16'd41680, 16'd59994});
	test_expansion(128'hcb2c98b3336f0221063cfe5cebab1926, {16'd14115, 16'd37133, 16'd37820, 16'd19387, 16'd18244, 16'd12316, 16'd33473, 16'd54383, 16'd18982, 16'd40076, 16'd7009, 16'd3677, 16'd54440, 16'd31310, 16'd48900, 16'd26175, 16'd58551, 16'd20610, 16'd4512, 16'd56282, 16'd37829, 16'd43628, 16'd53983, 16'd14688, 16'd6929, 16'd33884});
	test_expansion(128'h73af43cb1d88ea8c65f99322b0a4c7ff, {16'd1279, 16'd41156, 16'd53820, 16'd22152, 16'd50765, 16'd4026, 16'd56167, 16'd9443, 16'd59063, 16'd12076, 16'd46737, 16'd63749, 16'd61839, 16'd30477, 16'd893, 16'd18768, 16'd17627, 16'd8351, 16'd3761, 16'd57170, 16'd28330, 16'd42475, 16'd1337, 16'd51428, 16'd12093, 16'd27185});
	test_expansion(128'hb451568234a20ab8c6893b656cd8ef2f, {16'd11694, 16'd44249, 16'd64896, 16'd12672, 16'd4846, 16'd53218, 16'd53005, 16'd21675, 16'd24148, 16'd22914, 16'd41365, 16'd2545, 16'd48938, 16'd32418, 16'd9850, 16'd41213, 16'd60711, 16'd31987, 16'd20765, 16'd4724, 16'd31753, 16'd21843, 16'd61935, 16'd29091, 16'd51991, 16'd16189});
	test_expansion(128'h82df7df595bb16b52bbbcd5b83b5c80c, {16'd4408, 16'd2963, 16'd2095, 16'd16289, 16'd59753, 16'd1562, 16'd13332, 16'd55308, 16'd20647, 16'd2865, 16'd377, 16'd46260, 16'd28854, 16'd21902, 16'd6527, 16'd54867, 16'd17622, 16'd5705, 16'd22770, 16'd17997, 16'd64645, 16'd8005, 16'd30120, 16'd55455, 16'd40064, 16'd5233});
	test_expansion(128'hef2b3db4a43925613b1e241857eaf054, {16'd14949, 16'd43728, 16'd5327, 16'd4263, 16'd1530, 16'd30900, 16'd8755, 16'd19467, 16'd8162, 16'd62346, 16'd31347, 16'd2924, 16'd28903, 16'd25683, 16'd54380, 16'd24587, 16'd6166, 16'd49454, 16'd30662, 16'd6581, 16'd23406, 16'd54524, 16'd30434, 16'd42734, 16'd45005, 16'd1007});
	test_expansion(128'hb8b031b2b3b80a7a53d5dd085144e8d3, {16'd61386, 16'd32311, 16'd27586, 16'd43562, 16'd27027, 16'd42057, 16'd45923, 16'd43070, 16'd27236, 16'd19278, 16'd5810, 16'd35095, 16'd11310, 16'd35757, 16'd20092, 16'd47914, 16'd13130, 16'd14410, 16'd36719, 16'd20256, 16'd30798, 16'd34316, 16'd14382, 16'd24922, 16'd18734, 16'd44033});
	test_expansion(128'h460affe8e75ca0ebed8c002328104bc1, {16'd8394, 16'd33817, 16'd20185, 16'd23222, 16'd49849, 16'd52101, 16'd2250, 16'd59347, 16'd35363, 16'd59636, 16'd30066, 16'd41602, 16'd29326, 16'd25587, 16'd18225, 16'd19707, 16'd52577, 16'd7927, 16'd36927, 16'd20837, 16'd56331, 16'd46960, 16'd64528, 16'd28609, 16'd28194, 16'd64115});
	test_expansion(128'hf78774e51f97f3e500cd8232c32633f2, {16'd1271, 16'd18775, 16'd3223, 16'd62293, 16'd9370, 16'd16138, 16'd51708, 16'd26821, 16'd3738, 16'd55404, 16'd60226, 16'd24396, 16'd34445, 16'd57448, 16'd45494, 16'd64744, 16'd25316, 16'd5393, 16'd33841, 16'd16456, 16'd18176, 16'd27075, 16'd30670, 16'd11822, 16'd9448, 16'd1200});
	test_expansion(128'hec457ae6a245eef9e507bde1834b0307, {16'd2835, 16'd37304, 16'd58826, 16'd30295, 16'd9728, 16'd36066, 16'd19162, 16'd12943, 16'd40567, 16'd24114, 16'd19420, 16'd20166, 16'd9462, 16'd49705, 16'd18637, 16'd38787, 16'd13556, 16'd20747, 16'd17390, 16'd13173, 16'd30620, 16'd46093, 16'd5206, 16'd56967, 16'd25399, 16'd19716});
	test_expansion(128'hc92b7ce9ed7769180ce3209a5069de25, {16'd9849, 16'd1495, 16'd37154, 16'd46186, 16'd51131, 16'd1517, 16'd120, 16'd2417, 16'd27074, 16'd15140, 16'd35973, 16'd45921, 16'd37744, 16'd29371, 16'd50108, 16'd26549, 16'd37996, 16'd53585, 16'd14645, 16'd34198, 16'd56672, 16'd48985, 16'd768, 16'd16712, 16'd16225, 16'd37563});
	test_expansion(128'h8acc21c994feadfb4c6edbdb4c825359, {16'd59701, 16'd27402, 16'd38037, 16'd22809, 16'd65009, 16'd50562, 16'd51671, 16'd59087, 16'd34983, 16'd62023, 16'd58547, 16'd9755, 16'd39354, 16'd7171, 16'd863, 16'd1004, 16'd6934, 16'd25900, 16'd49539, 16'd5129, 16'd2676, 16'd44373, 16'd33397, 16'd20160, 16'd12743, 16'd36851});
	test_expansion(128'h9478ece113b91aec014c8fa64fe7746f, {16'd34885, 16'd10987, 16'd18182, 16'd10695, 16'd3002, 16'd43413, 16'd18266, 16'd17159, 16'd17450, 16'd10281, 16'd5411, 16'd36290, 16'd8290, 16'd5734, 16'd63519, 16'd32161, 16'd10637, 16'd59753, 16'd47110, 16'd34291, 16'd29524, 16'd22948, 16'd56596, 16'd13014, 16'd25761, 16'd40097});
	test_expansion(128'ha263f888af1cee4979d89da874a3a6b3, {16'd19838, 16'd57695, 16'd29257, 16'd42557, 16'd12096, 16'd59670, 16'd40617, 16'd52375, 16'd42822, 16'd44825, 16'd31709, 16'd10043, 16'd57805, 16'd24710, 16'd50403, 16'd53777, 16'd64567, 16'd16957, 16'd580, 16'd5768, 16'd52812, 16'd39861, 16'd20512, 16'd65460, 16'd49530, 16'd3749});
	test_expansion(128'h92e2216272a420fa1985d72d6ce40f31, {16'd44822, 16'd37211, 16'd35920, 16'd48853, 16'd40796, 16'd61058, 16'd25065, 16'd7711, 16'd38668, 16'd40428, 16'd30903, 16'd42055, 16'd17163, 16'd49962, 16'd52383, 16'd50074, 16'd41801, 16'd61346, 16'd36427, 16'd39492, 16'd35848, 16'd19451, 16'd8817, 16'd30744, 16'd15319, 16'd21506});
	test_expansion(128'he68d370a1002df892c2b2d13c6af5001, {16'd24230, 16'd11091, 16'd45901, 16'd39888, 16'd52053, 16'd43743, 16'd9249, 16'd27466, 16'd20821, 16'd25371, 16'd59394, 16'd8600, 16'd24246, 16'd61214, 16'd23186, 16'd1997, 16'd15074, 16'd25677, 16'd40498, 16'd29672, 16'd14132, 16'd23108, 16'd14013, 16'd25383, 16'd41033, 16'd22533});
	test_expansion(128'h43074b106e9ba7efcab3dd478fb6b055, {16'd40304, 16'd51756, 16'd6982, 16'd33674, 16'd16117, 16'd55016, 16'd8949, 16'd50561, 16'd43844, 16'd42560, 16'd32965, 16'd20155, 16'd887, 16'd44868, 16'd17656, 16'd37646, 16'd40244, 16'd46512, 16'd51736, 16'd4976, 16'd18855, 16'd61835, 16'd6037, 16'd30963, 16'd12086, 16'd13705});
	test_expansion(128'h42d7ca72dd24449d5d7e96074e93010a, {16'd59977, 16'd45602, 16'd37650, 16'd8307, 16'd20230, 16'd56325, 16'd48759, 16'd2110, 16'd44678, 16'd153, 16'd27093, 16'd43790, 16'd50250, 16'd64593, 16'd2291, 16'd54294, 16'd28069, 16'd32253, 16'd383, 16'd50099, 16'd36355, 16'd62146, 16'd34139, 16'd61678, 16'd14378, 16'd4999});
	test_expansion(128'h7d1b8cbc90b536e93af0a072ad267862, {16'd3568, 16'd39971, 16'd55533, 16'd44962, 16'd14344, 16'd60700, 16'd7223, 16'd797, 16'd38822, 16'd4651, 16'd63553, 16'd64889, 16'd53414, 16'd21733, 16'd35808, 16'd16059, 16'd22895, 16'd22396, 16'd58152, 16'd2104, 16'd53775, 16'd44666, 16'd36898, 16'd19336, 16'd53870, 16'd48403});
	test_expansion(128'hde526807efc72140f4983e860cca29f9, {16'd25816, 16'd40989, 16'd11638, 16'd45366, 16'd51399, 16'd23624, 16'd56959, 16'd36026, 16'd62577, 16'd61489, 16'd10584, 16'd20464, 16'd13335, 16'd35865, 16'd61697, 16'd3517, 16'd60983, 16'd9352, 16'd32511, 16'd21658, 16'd61824, 16'd39150, 16'd20803, 16'd55854, 16'd56359, 16'd58187});
	test_expansion(128'h2687ceee6aca3aef1239deba5c228397, {16'd60259, 16'd59537, 16'd54806, 16'd40806, 16'd29109, 16'd59016, 16'd45899, 16'd44476, 16'd39473, 16'd1094, 16'd50772, 16'd60242, 16'd22975, 16'd64307, 16'd5584, 16'd44104, 16'd32650, 16'd59657, 16'd11519, 16'd27943, 16'd50455, 16'd24358, 16'd28620, 16'd30818, 16'd19213, 16'd37472});
	test_expansion(128'h644c975ad6d0c80dcfb637baa36b4c0c, {16'd32765, 16'd1235, 16'd29685, 16'd60265, 16'd56268, 16'd32895, 16'd4768, 16'd4782, 16'd8758, 16'd48930, 16'd4387, 16'd39012, 16'd17360, 16'd43183, 16'd6214, 16'd47035, 16'd8510, 16'd31604, 16'd39712, 16'd21381, 16'd1416, 16'd56123, 16'd10317, 16'd57255, 16'd10862, 16'd12556});
	test_expansion(128'ha5fbaf8036ad693e8e399214fc4d9025, {16'd38769, 16'd23415, 16'd4898, 16'd42097, 16'd23939, 16'd19803, 16'd37290, 16'd27096, 16'd45795, 16'd21037, 16'd26588, 16'd43969, 16'd10905, 16'd37749, 16'd23014, 16'd48403, 16'd28573, 16'd17170, 16'd48480, 16'd27091, 16'd39690, 16'd6103, 16'd54876, 16'd59339, 16'd48658, 16'd49307});
	test_expansion(128'he9563d916c41657cbb3305ab30d581bb, {16'd27092, 16'd33772, 16'd20745, 16'd36695, 16'd52703, 16'd26538, 16'd3068, 16'd30244, 16'd48776, 16'd40457, 16'd57856, 16'd13262, 16'd23106, 16'd19620, 16'd44936, 16'd10666, 16'd48970, 16'd28219, 16'd63240, 16'd36015, 16'd56812, 16'd42648, 16'd53111, 16'd6783, 16'd16158, 16'd44484});
	test_expansion(128'hb9e6b8d93159aa095d3c8704714dda8a, {16'd22154, 16'd52519, 16'd8939, 16'd40926, 16'd8301, 16'd47330, 16'd2675, 16'd46389, 16'd10716, 16'd61021, 16'd43898, 16'd29849, 16'd25195, 16'd6685, 16'd13056, 16'd29939, 16'd64326, 16'd59805, 16'd62471, 16'd14900, 16'd50757, 16'd14223, 16'd41964, 16'd58459, 16'd61042, 16'd40245});
	test_expansion(128'h06cd98f81f67966a51e7815b4b603eb9, {16'd1970, 16'd49035, 16'd59681, 16'd57327, 16'd32720, 16'd31942, 16'd17754, 16'd16755, 16'd34109, 16'd25239, 16'd62619, 16'd33301, 16'd62044, 16'd5459, 16'd34376, 16'd57860, 16'd20146, 16'd16441, 16'd5838, 16'd45422, 16'd57973, 16'd23681, 16'd2569, 16'd63131, 16'd19436, 16'd64729});
	test_expansion(128'hdfbbabe1b6bf569f67f44160751d541a, {16'd44825, 16'd17675, 16'd16738, 16'd41494, 16'd12649, 16'd61458, 16'd48276, 16'd19809, 16'd52717, 16'd18938, 16'd19656, 16'd28649, 16'd64907, 16'd25035, 16'd20028, 16'd51584, 16'd29123, 16'd50969, 16'd8178, 16'd12083, 16'd40954, 16'd7659, 16'd63223, 16'd16837, 16'd22344, 16'd53481});
	test_expansion(128'ha7c7906eb82f22fef90952ac16f8d8bc, {16'd65295, 16'd38257, 16'd50283, 16'd41597, 16'd61962, 16'd28841, 16'd18550, 16'd21424, 16'd46908, 16'd13036, 16'd12228, 16'd45958, 16'd46001, 16'd21684, 16'd30603, 16'd60674, 16'd39730, 16'd25172, 16'd37355, 16'd50568, 16'd1056, 16'd15257, 16'd25080, 16'd21955, 16'd31005, 16'd44782});
	test_expansion(128'hbf331734b1b0c5609b87f0d88e53faf1, {16'd50672, 16'd8954, 16'd41397, 16'd47797, 16'd34500, 16'd47883, 16'd10826, 16'd16183, 16'd4014, 16'd49895, 16'd35717, 16'd24356, 16'd26507, 16'd32784, 16'd130, 16'd56637, 16'd41066, 16'd38349, 16'd12481, 16'd14682, 16'd62920, 16'd46553, 16'd37676, 16'd49562, 16'd11228, 16'd38711});
	test_expansion(128'h9c14c19f24601a599c478b51689740db, {16'd11166, 16'd26879, 16'd33978, 16'd47547, 16'd60427, 16'd39572, 16'd13233, 16'd3652, 16'd44785, 16'd39388, 16'd12999, 16'd1381, 16'd11817, 16'd1719, 16'd58202, 16'd23388, 16'd49754, 16'd37941, 16'd537, 16'd43729, 16'd27733, 16'd6432, 16'd37066, 16'd40802, 16'd49915, 16'd15920});
	test_expansion(128'hf8409533413ee6220cc1d6fc03396fc3, {16'd62943, 16'd45367, 16'd4895, 16'd5140, 16'd13593, 16'd31025, 16'd26274, 16'd33551, 16'd49334, 16'd27669, 16'd29644, 16'd20461, 16'd18983, 16'd29906, 16'd55629, 16'd37396, 16'd19370, 16'd57504, 16'd63206, 16'd42263, 16'd38334, 16'd45905, 16'd39857, 16'd13424, 16'd6369, 16'd45114});
	test_expansion(128'h1f98c556fd7ff37f5995cd029a03c1e3, {16'd55350, 16'd56625, 16'd43862, 16'd32024, 16'd21557, 16'd47813, 16'd51617, 16'd44943, 16'd35907, 16'd5265, 16'd4703, 16'd9587, 16'd21598, 16'd42626, 16'd22054, 16'd57842, 16'd39517, 16'd59629, 16'd45737, 16'd11725, 16'd47275, 16'd26827, 16'd4775, 16'd39124, 16'd35440, 16'd25047});
	test_expansion(128'h52afb9cb90c6f0953890f40b4c17a2d0, {16'd5671, 16'd38089, 16'd25249, 16'd7654, 16'd19278, 16'd12822, 16'd2498, 16'd5510, 16'd10281, 16'd39420, 16'd6098, 16'd29919, 16'd58658, 16'd12244, 16'd51214, 16'd14728, 16'd28522, 16'd32858, 16'd47602, 16'd61049, 16'd28576, 16'd14429, 16'd11974, 16'd1770, 16'd57307, 16'd65135});
	test_expansion(128'hf394b82acf4d8fddd3a80d1e3f5df4cb, {16'd48803, 16'd64956, 16'd58740, 16'd33281, 16'd11325, 16'd4486, 16'd51888, 16'd9680, 16'd10083, 16'd60128, 16'd40952, 16'd34727, 16'd16106, 16'd39082, 16'd44926, 16'd45297, 16'd28787, 16'd33625, 16'd27394, 16'd54440, 16'd35045, 16'd31169, 16'd3578, 16'd44711, 16'd48416, 16'd6442});
	test_expansion(128'h9ec63fa0d6356f0e45ec5d610e82fd40, {16'd22944, 16'd6469, 16'd60583, 16'd30027, 16'd16320, 16'd13830, 16'd12519, 16'd20002, 16'd31135, 16'd59432, 16'd62612, 16'd5441, 16'd64473, 16'd56529, 16'd5991, 16'd41222, 16'd16935, 16'd2436, 16'd42280, 16'd54080, 16'd38663, 16'd53721, 16'd55942, 16'd41674, 16'd11729, 16'd12664});
	test_expansion(128'h67035ca5e31ea3a51b45753bb229e312, {16'd52725, 16'd64703, 16'd53627, 16'd53810, 16'd83, 16'd37384, 16'd2073, 16'd5261, 16'd56556, 16'd31972, 16'd39509, 16'd48889, 16'd2516, 16'd38017, 16'd54087, 16'd48330, 16'd39940, 16'd13702, 16'd64185, 16'd62186, 16'd3533, 16'd54730, 16'd4478, 16'd54591, 16'd19729, 16'd18658});
	test_expansion(128'h36d82f984b7711a92558d4f6237f2de5, {16'd8001, 16'd44479, 16'd4246, 16'd681, 16'd25118, 16'd3430, 16'd421, 16'd19856, 16'd10009, 16'd31029, 16'd6529, 16'd16556, 16'd28888, 16'd7605, 16'd58267, 16'd58707, 16'd38511, 16'd52510, 16'd32003, 16'd64781, 16'd40280, 16'd46639, 16'd24509, 16'd58817, 16'd41218, 16'd64790});
	test_expansion(128'hc3a02e147ce4ff41ae435a7ce38da209, {16'd413, 16'd37559, 16'd54602, 16'd42702, 16'd60632, 16'd40479, 16'd40811, 16'd21457, 16'd34986, 16'd8769, 16'd27463, 16'd48696, 16'd8710, 16'd24337, 16'd62845, 16'd2837, 16'd7713, 16'd63130, 16'd1798, 16'd40885, 16'd33608, 16'd5683, 16'd65427, 16'd10558, 16'd46177, 16'd36426});
	test_expansion(128'h113ada98081e322e2062963b056e08da, {16'd57716, 16'd64747, 16'd63021, 16'd11950, 16'd714, 16'd30989, 16'd57728, 16'd47056, 16'd27090, 16'd16539, 16'd9198, 16'd56224, 16'd40837, 16'd49163, 16'd40315, 16'd5042, 16'd49610, 16'd20124, 16'd58681, 16'd47079, 16'd613, 16'd1038, 16'd14618, 16'd59771, 16'd10083, 16'd24568});
	test_expansion(128'hcec06b01c63f493205808a300e4f08ce, {16'd64944, 16'd27964, 16'd18170, 16'd39437, 16'd17464, 16'd35611, 16'd27333, 16'd34928, 16'd12174, 16'd10927, 16'd41705, 16'd28216, 16'd26993, 16'd259, 16'd16905, 16'd9380, 16'd56451, 16'd30709, 16'd24372, 16'd52394, 16'd19919, 16'd12481, 16'd3363, 16'd33614, 16'd34779, 16'd34608});
	test_expansion(128'h64e5e2fc8e615ed0483fc8221d929e93, {16'd8442, 16'd39733, 16'd10031, 16'd27623, 16'd2796, 16'd8372, 16'd32489, 16'd46366, 16'd8138, 16'd37234, 16'd62937, 16'd8856, 16'd27362, 16'd27030, 16'd58219, 16'd44024, 16'd3907, 16'd53264, 16'd3622, 16'd39699, 16'd53361, 16'd17963, 16'd44815, 16'd21422, 16'd59529, 16'd8810});
	test_expansion(128'h39cfb04ba4dd66851f1da1fb953e6544, {16'd9559, 16'd18041, 16'd41130, 16'd31401, 16'd20261, 16'd34721, 16'd26593, 16'd30812, 16'd46549, 16'd52756, 16'd14857, 16'd21704, 16'd57678, 16'd855, 16'd6629, 16'd36581, 16'd42735, 16'd56509, 16'd13328, 16'd3303, 16'd1055, 16'd26994, 16'd16620, 16'd22586, 16'd23110, 16'd48865});
	test_expansion(128'h9715cbb02016885a60de250b2f39d057, {16'd31388, 16'd21887, 16'd33307, 16'd13039, 16'd18378, 16'd63771, 16'd19044, 16'd42192, 16'd39756, 16'd30311, 16'd32688, 16'd4562, 16'd22195, 16'd53903, 16'd20335, 16'd989, 16'd9800, 16'd59656, 16'd9023, 16'd30581, 16'd11053, 16'd9218, 16'd41146, 16'd60498, 16'd32631, 16'd13123});
	test_expansion(128'h8fc92248a21b97d229d7db199c933a58, {16'd44609, 16'd4670, 16'd22300, 16'd61500, 16'd53676, 16'd25367, 16'd59412, 16'd26951, 16'd51513, 16'd34670, 16'd41743, 16'd62650, 16'd18516, 16'd12021, 16'd17253, 16'd16785, 16'd12502, 16'd15213, 16'd4315, 16'd64101, 16'd19366, 16'd65, 16'd22476, 16'd48716, 16'd14345, 16'd57672});
	test_expansion(128'h499be4b47fec83a3c4fbffd5140d8e0b, {16'd49430, 16'd34803, 16'd25321, 16'd21103, 16'd64231, 16'd18596, 16'd56982, 16'd172, 16'd62917, 16'd61757, 16'd43359, 16'd14405, 16'd28112, 16'd15893, 16'd3040, 16'd61562, 16'd50576, 16'd1329, 16'd46677, 16'd38788, 16'd11319, 16'd64225, 16'd23922, 16'd44614, 16'd30292, 16'd17765});
	test_expansion(128'h6e5967f048150cafbfc06fa5bff02b66, {16'd32156, 16'd55783, 16'd35938, 16'd49862, 16'd54272, 16'd18157, 16'd4120, 16'd31137, 16'd61110, 16'd10406, 16'd24665, 16'd45541, 16'd63668, 16'd14388, 16'd57484, 16'd28487, 16'd6056, 16'd57594, 16'd34056, 16'd26081, 16'd310, 16'd23077, 16'd54939, 16'd37655, 16'd15440, 16'd6131});
	test_expansion(128'h34a3769e5dee6eac26bb24d03d27053e, {16'd30661, 16'd24540, 16'd65261, 16'd34494, 16'd28880, 16'd24837, 16'd18231, 16'd45256, 16'd61150, 16'd42448, 16'd18271, 16'd24792, 16'd49941, 16'd53646, 16'd60376, 16'd43028, 16'd9082, 16'd39545, 16'd36151, 16'd44197, 16'd12089, 16'd55280, 16'd60816, 16'd4323, 16'd35731, 16'd64419});
	test_expansion(128'hfb2dd163f02f55b9d141762039c1b970, {16'd65058, 16'd40643, 16'd58108, 16'd32194, 16'd21001, 16'd21127, 16'd32271, 16'd64218, 16'd37127, 16'd50622, 16'd41495, 16'd53254, 16'd22288, 16'd29533, 16'd16524, 16'd49168, 16'd41598, 16'd13778, 16'd17427, 16'd38177, 16'd49514, 16'd12840, 16'd61916, 16'd34241, 16'd62981, 16'd4354});
	test_expansion(128'h259a5a4ed1b30978b69ff1b68024c9b2, {16'd8734, 16'd51994, 16'd52354, 16'd14654, 16'd742, 16'd64882, 16'd36847, 16'd12617, 16'd29560, 16'd12101, 16'd16801, 16'd196, 16'd63706, 16'd17437, 16'd59183, 16'd42986, 16'd57595, 16'd39019, 16'd61335, 16'd3095, 16'd48229, 16'd58452, 16'd11832, 16'd60132, 16'd46059, 16'd2902});
	test_expansion(128'h33f57fd02cb0201df8884e0c90aaa2c0, {16'd33473, 16'd44802, 16'd23524, 16'd7117, 16'd25902, 16'd14518, 16'd48917, 16'd53858, 16'd60280, 16'd38135, 16'd32863, 16'd52855, 16'd38757, 16'd15977, 16'd21190, 16'd22240, 16'd41834, 16'd49292, 16'd44684, 16'd21218, 16'd32818, 16'd2748, 16'd31465, 16'd60780, 16'd25984, 16'd44679});
	test_expansion(128'h0777c354beedb1a648e39f8f7a3044f5, {16'd21089, 16'd40645, 16'd6969, 16'd26789, 16'd4017, 16'd57135, 16'd62877, 16'd46675, 16'd44025, 16'd2292, 16'd57849, 16'd27367, 16'd59504, 16'd36166, 16'd26600, 16'd32243, 16'd24046, 16'd25663, 16'd43198, 16'd24966, 16'd44066, 16'd45852, 16'd23067, 16'd4635, 16'd17509, 16'd24208});
	test_expansion(128'ha83c7215761cd5fd13161ee1236b0629, {16'd32677, 16'd45105, 16'd25439, 16'd20257, 16'd14316, 16'd506, 16'd49020, 16'd8884, 16'd45113, 16'd876, 16'd29776, 16'd58696, 16'd41265, 16'd16497, 16'd61898, 16'd30718, 16'd16241, 16'd1578, 16'd44877, 16'd13137, 16'd54954, 16'd42239, 16'd28233, 16'd56114, 16'd10075, 16'd38849});
	test_expansion(128'hdf2f7a3abaf9eed5d1b736e8301629e9, {16'd3010, 16'd55895, 16'd58497, 16'd18969, 16'd48133, 16'd26197, 16'd47399, 16'd30033, 16'd36352, 16'd15569, 16'd1871, 16'd54435, 16'd40650, 16'd4798, 16'd65135, 16'd14917, 16'd42474, 16'd28890, 16'd64239, 16'd5695, 16'd790, 16'd5041, 16'd16843, 16'd41809, 16'd38064, 16'd30704});
	test_expansion(128'hb6335a666c204175d1f27efc0edb828d, {16'd45337, 16'd27233, 16'd54250, 16'd56811, 16'd3665, 16'd47885, 16'd29559, 16'd20591, 16'd5793, 16'd9898, 16'd64198, 16'd26437, 16'd51280, 16'd33004, 16'd61213, 16'd52457, 16'd60449, 16'd58251, 16'd15634, 16'd45752, 16'd14739, 16'd18652, 16'd34592, 16'd38340, 16'd815, 16'd20885});
	test_expansion(128'hb3ff1594eff4ee4bf01cd3d64a531ea5, {16'd63764, 16'd6274, 16'd5882, 16'd62540, 16'd18973, 16'd35301, 16'd10761, 16'd61213, 16'd49739, 16'd8570, 16'd1314, 16'd20010, 16'd32824, 16'd2588, 16'd57487, 16'd50168, 16'd13973, 16'd17907, 16'd45223, 16'd9846, 16'd57215, 16'd62026, 16'd38765, 16'd53433, 16'd29279, 16'd3804});
	test_expansion(128'h2b9380b08d97619f07be571b15c17346, {16'd26100, 16'd62013, 16'd33779, 16'd29266, 16'd2935, 16'd11904, 16'd28833, 16'd58800, 16'd25588, 16'd9565, 16'd44492, 16'd47408, 16'd20642, 16'd47294, 16'd1905, 16'd57690, 16'd21583, 16'd20809, 16'd6505, 16'd47190, 16'd50309, 16'd60132, 16'd60140, 16'd10143, 16'd14747, 16'd10970});
	test_expansion(128'h900a29767248e8e926fdb4a21df99b73, {16'd27774, 16'd19941, 16'd28608, 16'd61025, 16'd17659, 16'd48011, 16'd850, 16'd24700, 16'd25175, 16'd24613, 16'd12723, 16'd13584, 16'd9656, 16'd36863, 16'd28779, 16'd48566, 16'd7518, 16'd556, 16'd49908, 16'd15203, 16'd42497, 16'd45570, 16'd64481, 16'd24853, 16'd46707, 16'd43638});
	test_expansion(128'hd7f5f6ddba6c36b8f3c9a19a5b32d4e0, {16'd3107, 16'd15147, 16'd41601, 16'd33163, 16'd42167, 16'd43246, 16'd65151, 16'd49297, 16'd18395, 16'd46819, 16'd60465, 16'd476, 16'd65421, 16'd26879, 16'd55640, 16'd39215, 16'd15746, 16'd54505, 16'd33132, 16'd30604, 16'd28654, 16'd63250, 16'd21148, 16'd10050, 16'd2817, 16'd50060});
	test_expansion(128'ha3fc824327c539c0f68742509f6bcca3, {16'd58613, 16'd47641, 16'd51864, 16'd54259, 16'd7826, 16'd5433, 16'd44230, 16'd40743, 16'd27624, 16'd33927, 16'd22546, 16'd22265, 16'd50930, 16'd4934, 16'd45945, 16'd38003, 16'd49658, 16'd57015, 16'd4974, 16'd52461, 16'd35050, 16'd16340, 16'd40174, 16'd15807, 16'd39428, 16'd14034});
	test_expansion(128'h2ab51bd257643060979074a0606fc33e, {16'd18501, 16'd35191, 16'd11205, 16'd16591, 16'd41601, 16'd43131, 16'd6998, 16'd6654, 16'd2063, 16'd39398, 16'd32088, 16'd14883, 16'd28083, 16'd35998, 16'd2755, 16'd46622, 16'd54768, 16'd3954, 16'd51647, 16'd59737, 16'd1032, 16'd9328, 16'd40716, 16'd29563, 16'd65188, 16'd18545});
	test_expansion(128'hf668da9a3c7f86d71bb2068815c28654, {16'd62775, 16'd49727, 16'd19410, 16'd56523, 16'd64008, 16'd63951, 16'd15376, 16'd49329, 16'd16447, 16'd61595, 16'd39849, 16'd35769, 16'd50093, 16'd11581, 16'd24012, 16'd62632, 16'd46722, 16'd38748, 16'd416, 16'd23682, 16'd19382, 16'd32496, 16'd21698, 16'd64379, 16'd43104, 16'd9759});
	test_expansion(128'h6283c11ea8afc114dc62df4c49877744, {16'd52755, 16'd10459, 16'd22449, 16'd22998, 16'd49221, 16'd49698, 16'd48566, 16'd55953, 16'd58847, 16'd2969, 16'd7846, 16'd11621, 16'd25876, 16'd11110, 16'd49767, 16'd33952, 16'd54180, 16'd32842, 16'd32755, 16'd20322, 16'd5466, 16'd61081, 16'd19956, 16'd17967, 16'd52838, 16'd8034});
	test_expansion(128'hf72f6c5c24451be3e16f5c000a12756b, {16'd11443, 16'd20931, 16'd32683, 16'd16155, 16'd49951, 16'd12533, 16'd23954, 16'd51114, 16'd62692, 16'd24775, 16'd5149, 16'd26784, 16'd30133, 16'd12165, 16'd9557, 16'd11028, 16'd1674, 16'd55864, 16'd10916, 16'd60801, 16'd48715, 16'd38550, 16'd16257, 16'd664, 16'd55323, 16'd47477});
	test_expansion(128'h0200e138026c7fbed6915fe6ede9642d, {16'd48891, 16'd7539, 16'd48710, 16'd12451, 16'd4909, 16'd47806, 16'd2084, 16'd23485, 16'd51479, 16'd31483, 16'd64665, 16'd52719, 16'd47529, 16'd20778, 16'd22871, 16'd34058, 16'd17156, 16'd56977, 16'd25596, 16'd15420, 16'd30196, 16'd7889, 16'd20734, 16'd28396, 16'd15764, 16'd59728});
	test_expansion(128'h7f816faad4ca3995ef306d36eb328a1b, {16'd25169, 16'd5611, 16'd63031, 16'd8790, 16'd32667, 16'd30000, 16'd28557, 16'd54800, 16'd10122, 16'd47432, 16'd54152, 16'd25157, 16'd13032, 16'd34980, 16'd33781, 16'd57351, 16'd44441, 16'd45478, 16'd34294, 16'd23409, 16'd43671, 16'd42213, 16'd14536, 16'd2240, 16'd4162, 16'd16492});
	test_expansion(128'h10720de9cd22d59054aa0c5469a0a0e8, {16'd61316, 16'd52686, 16'd62386, 16'd49781, 16'd45377, 16'd872, 16'd11010, 16'd32781, 16'd2644, 16'd17373, 16'd36961, 16'd41835, 16'd40692, 16'd21816, 16'd7734, 16'd57353, 16'd6033, 16'd25363, 16'd55714, 16'd40683, 16'd17906, 16'd54406, 16'd52131, 16'd46670, 16'd34968, 16'd19401});
	test_expansion(128'h168793054b3812a3a9aa5be116049f99, {16'd49810, 16'd59955, 16'd19405, 16'd51349, 16'd28975, 16'd48116, 16'd48875, 16'd21260, 16'd28491, 16'd31413, 16'd62086, 16'd53848, 16'd47999, 16'd2515, 16'd4486, 16'd15086, 16'd36520, 16'd31090, 16'd59729, 16'd26126, 16'd24380, 16'd34131, 16'd41539, 16'd32302, 16'd36036, 16'd5451});
	test_expansion(128'h2221e728745f1e9fe3e1a40c823226ed, {16'd6101, 16'd37697, 16'd46662, 16'd65469, 16'd7096, 16'd8597, 16'd35409, 16'd27734, 16'd9224, 16'd32517, 16'd43981, 16'd22928, 16'd16458, 16'd62154, 16'd64975, 16'd50850, 16'd11891, 16'd34474, 16'd14318, 16'd5202, 16'd50583, 16'd36970, 16'd4406, 16'd16197, 16'd12599, 16'd22360});
	test_expansion(128'h209387ccde34446b4b7e84a9a9c91e64, {16'd58715, 16'd54918, 16'd45583, 16'd4463, 16'd29468, 16'd14575, 16'd57630, 16'd24886, 16'd40363, 16'd29766, 16'd29963, 16'd1327, 16'd19410, 16'd43670, 16'd44446, 16'd60086, 16'd35610, 16'd44367, 16'd54364, 16'd23520, 16'd35424, 16'd26387, 16'd9222, 16'd31476, 16'd47400, 16'd3207});
	test_expansion(128'h5377ad45219234c370b2c2c2d2ed1a40, {16'd64322, 16'd45284, 16'd29805, 16'd55278, 16'd35738, 16'd2181, 16'd15412, 16'd7935, 16'd29795, 16'd54436, 16'd39695, 16'd14665, 16'd12734, 16'd60735, 16'd28439, 16'd62198, 16'd61078, 16'd57059, 16'd22371, 16'd60305, 16'd51577, 16'd19127, 16'd42312, 16'd2351, 16'd35568, 16'd45524});
	test_expansion(128'hf8fc8c60db7409ca439181e1ab5822b2, {16'd9336, 16'd45006, 16'd62034, 16'd25790, 16'd63293, 16'd59872, 16'd2757, 16'd28700, 16'd24450, 16'd46198, 16'd28354, 16'd31135, 16'd30392, 16'd20237, 16'd48234, 16'd59280, 16'd34779, 16'd43746, 16'd52589, 16'd58978, 16'd28546, 16'd4243, 16'd13146, 16'd24999, 16'd2785, 16'd53707});
	test_expansion(128'h05c9c7cddac0f330c69a18ee88b80ff3, {16'd52295, 16'd31005, 16'd18661, 16'd18660, 16'd16298, 16'd20644, 16'd55224, 16'd980, 16'd9456, 16'd47287, 16'd3835, 16'd31500, 16'd62115, 16'd31340, 16'd8532, 16'd3970, 16'd15294, 16'd46443, 16'd61420, 16'd20219, 16'd8964, 16'd16137, 16'd10811, 16'd35884, 16'd1202, 16'd52878});
	test_expansion(128'h957eaf2b4fd986f1993624d1c030292b, {16'd45532, 16'd57050, 16'd51264, 16'd25618, 16'd46847, 16'd31563, 16'd21355, 16'd2609, 16'd43653, 16'd51782, 16'd31337, 16'd33877, 16'd44101, 16'd14490, 16'd21302, 16'd39231, 16'd13251, 16'd22196, 16'd6388, 16'd50164, 16'd21834, 16'd39965, 16'd41683, 16'd27887, 16'd29568, 16'd11584});
	test_expansion(128'hedc067f190b0e69eb770079d4f492925, {16'd12706, 16'd20122, 16'd2039, 16'd60289, 16'd31917, 16'd51581, 16'd13316, 16'd16360, 16'd30933, 16'd38860, 16'd19015, 16'd57192, 16'd55457, 16'd34143, 16'd22301, 16'd10581, 16'd9151, 16'd50396, 16'd40376, 16'd34540, 16'd46375, 16'd18477, 16'd37249, 16'd57494, 16'd41618, 16'd55153});
	test_expansion(128'hdc1812ab9309048f014147f38107c870, {16'd12054, 16'd9639, 16'd48625, 16'd24874, 16'd28287, 16'd17483, 16'd26410, 16'd26620, 16'd38412, 16'd57056, 16'd61577, 16'd65145, 16'd26493, 16'd5023, 16'd8101, 16'd58372, 16'd2408, 16'd48298, 16'd26263, 16'd609, 16'd43591, 16'd24288, 16'd38363, 16'd738, 16'd61896, 16'd31165});
	test_expansion(128'h890b54fd46ece356838eb486b655e955, {16'd9617, 16'd1710, 16'd51769, 16'd21180, 16'd50324, 16'd15866, 16'd31438, 16'd44758, 16'd1721, 16'd56616, 16'd387, 16'd63556, 16'd60408, 16'd15625, 16'd40567, 16'd27765, 16'd42046, 16'd9627, 16'd58056, 16'd17348, 16'd23820, 16'd26526, 16'd39675, 16'd10431, 16'd23410, 16'd361});
	test_expansion(128'hb56d345cea52618c915c42dfc15167e6, {16'd57649, 16'd33732, 16'd10128, 16'd65225, 16'd40635, 16'd21192, 16'd802, 16'd11553, 16'd60171, 16'd31069, 16'd14037, 16'd18759, 16'd34260, 16'd22339, 16'd27582, 16'd2566, 16'd20078, 16'd50905, 16'd14995, 16'd32585, 16'd65113, 16'd48455, 16'd28348, 16'd33433, 16'd11132, 16'd34298});
	test_expansion(128'hf71f0350767d5f11c954ea236835dfcc, {16'd45626, 16'd12082, 16'd47209, 16'd17253, 16'd49444, 16'd19956, 16'd53754, 16'd56584, 16'd17202, 16'd6278, 16'd32902, 16'd25535, 16'd44688, 16'd18242, 16'd19891, 16'd48427, 16'd35280, 16'd27841, 16'd31139, 16'd33007, 16'd61630, 16'd49793, 16'd36555, 16'd17364, 16'd34118, 16'd16293});
	test_expansion(128'hda26216ef088288cce2ab9c5e823d68b, {16'd36770, 16'd6812, 16'd41821, 16'd20962, 16'd14744, 16'd62030, 16'd58818, 16'd18849, 16'd48396, 16'd43835, 16'd53454, 16'd22291, 16'd29861, 16'd50715, 16'd28249, 16'd13683, 16'd30463, 16'd6537, 16'd20468, 16'd37776, 16'd39327, 16'd48906, 16'd6537, 16'd22132, 16'd40177, 16'd39031});
	test_expansion(128'h65aaec081eece7aac1aa2bc4be4943f2, {16'd13681, 16'd34910, 16'd27325, 16'd17641, 16'd65125, 16'd28026, 16'd41150, 16'd33286, 16'd22419, 16'd44388, 16'd39385, 16'd25642, 16'd35889, 16'd52767, 16'd16642, 16'd49796, 16'd54067, 16'd33504, 16'd12910, 16'd16927, 16'd56085, 16'd31281, 16'd31754, 16'd20902, 16'd40422, 16'd35661});
	test_expansion(128'h9a3a629b0f62497881c2d61a83b98ec4, {16'd991, 16'd26966, 16'd26434, 16'd31588, 16'd23565, 16'd45940, 16'd18762, 16'd29563, 16'd51096, 16'd50869, 16'd41444, 16'd63535, 16'd41993, 16'd10514, 16'd6206, 16'd60479, 16'd8073, 16'd42990, 16'd59830, 16'd56692, 16'd47060, 16'd20552, 16'd17206, 16'd59311, 16'd6346, 16'd34496});
	test_expansion(128'h15e7d7406c47f16e3e0b794f91ac45fd, {16'd54177, 16'd36548, 16'd7576, 16'd60947, 16'd23737, 16'd18342, 16'd22533, 16'd5208, 16'd41684, 16'd32808, 16'd15657, 16'd56882, 16'd35904, 16'd21929, 16'd30805, 16'd53153, 16'd28182, 16'd4041, 16'd41317, 16'd18206, 16'd58616, 16'd58513, 16'd51148, 16'd57782, 16'd24440, 16'd22450});
	test_expansion(128'h05becf7d9a574f83a282232252fd9894, {16'd49017, 16'd39354, 16'd23788, 16'd60451, 16'd14483, 16'd9169, 16'd33304, 16'd60226, 16'd57222, 16'd65238, 16'd1130, 16'd39899, 16'd34370, 16'd9213, 16'd51476, 16'd9498, 16'd21075, 16'd63775, 16'd31568, 16'd34969, 16'd42498, 16'd11608, 16'd41293, 16'd57101, 16'd59850, 16'd55911});
	test_expansion(128'hdcfd9c453ed4ccfbd54d08d6f53e2685, {16'd61146, 16'd51618, 16'd62690, 16'd37175, 16'd20913, 16'd60437, 16'd6675, 16'd19361, 16'd5045, 16'd23549, 16'd38657, 16'd3426, 16'd62531, 16'd41379, 16'd21995, 16'd55046, 16'd35050, 16'd2382, 16'd5240, 16'd29713, 16'd7735, 16'd60442, 16'd48169, 16'd10442, 16'd58246, 16'd3678});
	test_expansion(128'ha575a8dd64bc866ae62d1d5e20eba0d0, {16'd56861, 16'd6366, 16'd28068, 16'd57677, 16'd8848, 16'd29600, 16'd26738, 16'd17170, 16'd43948, 16'd24454, 16'd15407, 16'd42564, 16'd40606, 16'd62058, 16'd17497, 16'd46174, 16'd500, 16'd46526, 16'd49783, 16'd23873, 16'd37488, 16'd37185, 16'd19034, 16'd37219, 16'd9499, 16'd27909});
	test_expansion(128'h409bb0e5357636dab5049a960008dacb, {16'd50778, 16'd37184, 16'd37724, 16'd10439, 16'd39420, 16'd52732, 16'd8240, 16'd43205, 16'd23810, 16'd8702, 16'd5578, 16'd55128, 16'd59238, 16'd5580, 16'd42593, 16'd14365, 16'd40730, 16'd39930, 16'd3578, 16'd14049, 16'd53660, 16'd39855, 16'd11237, 16'd31860, 16'd36390, 16'd62230});
	test_expansion(128'h7e4cf360fcbc85b7eddefc05d4f9debd, {16'd31266, 16'd44428, 16'd47174, 16'd26182, 16'd29320, 16'd39790, 16'd22077, 16'd1631, 16'd50187, 16'd46408, 16'd28329, 16'd61459, 16'd8600, 16'd28391, 16'd46699, 16'd65451, 16'd56035, 16'd61581, 16'd4631, 16'd10028, 16'd42315, 16'd47714, 16'd64533, 16'd3497, 16'd43787, 16'd9842});
	test_expansion(128'hb30c9f06038ed18a10c2f893c6293576, {16'd50540, 16'd54407, 16'd57240, 16'd35669, 16'd36500, 16'd52781, 16'd25241, 16'd59726, 16'd42390, 16'd10443, 16'd40837, 16'd36635, 16'd5747, 16'd24317, 16'd2952, 16'd28802, 16'd5891, 16'd2681, 16'd28741, 16'd59149, 16'd22406, 16'd45330, 16'd17450, 16'd19045, 16'd20116, 16'd5676});
	test_expansion(128'ha4374c1acd2327b6b874cc3188f1326f, {16'd44551, 16'd13964, 16'd50648, 16'd45382, 16'd49855, 16'd35172, 16'd27458, 16'd59087, 16'd56009, 16'd22328, 16'd3545, 16'd48376, 16'd29391, 16'd56325, 16'd8683, 16'd40580, 16'd8068, 16'd38290, 16'd44562, 16'd64711, 16'd19847, 16'd7240, 16'd8924, 16'd20644, 16'd31730, 16'd35401});
	test_expansion(128'h366f5e99ea44b24caaa28594da870191, {16'd475, 16'd22151, 16'd22217, 16'd35215, 16'd26049, 16'd19133, 16'd31213, 16'd55254, 16'd25204, 16'd5993, 16'd21925, 16'd23164, 16'd27757, 16'd11101, 16'd393, 16'd41479, 16'd11226, 16'd20244, 16'd31035, 16'd44190, 16'd15418, 16'd27570, 16'd57197, 16'd29711, 16'd59474, 16'd34219});
	test_expansion(128'h8d8d6e15a6699694fa22b9ef8fefe861, {16'd63597, 16'd4045, 16'd45086, 16'd44748, 16'd7536, 16'd6993, 16'd32146, 16'd55601, 16'd20803, 16'd57594, 16'd33727, 16'd64163, 16'd27306, 16'd3639, 16'd5159, 16'd1684, 16'd53464, 16'd40833, 16'd40569, 16'd13409, 16'd62, 16'd39266, 16'd63983, 16'd16578, 16'd6950, 16'd11325});
	test_expansion(128'h6bf02b04d18c30dbb88944fed6d4d9a8, {16'd53805, 16'd6539, 16'd2566, 16'd265, 16'd23536, 16'd10890, 16'd47170, 16'd5763, 16'd46748, 16'd21727, 16'd19605, 16'd25854, 16'd52403, 16'd23370, 16'd53228, 16'd15642, 16'd6333, 16'd18937, 16'd49504, 16'd45112, 16'd42464, 16'd3476, 16'd46191, 16'd23473, 16'd34872, 16'd61888});
	test_expansion(128'h4837722032d43c4f5ac882b7f743d9ad, {16'd2168, 16'd60843, 16'd10388, 16'd36148, 16'd16325, 16'd2324, 16'd55981, 16'd2801, 16'd20662, 16'd20306, 16'd6634, 16'd39571, 16'd34409, 16'd18818, 16'd10678, 16'd55170, 16'd56887, 16'd37887, 16'd2110, 16'd36052, 16'd34562, 16'd7704, 16'd6575, 16'd34479, 16'd35646, 16'd4376});
	test_expansion(128'h1b5c0811336beb7a4494181d4c19f865, {16'd13589, 16'd30715, 16'd19923, 16'd34509, 16'd61146, 16'd63631, 16'd32286, 16'd5939, 16'd12515, 16'd55800, 16'd21608, 16'd64750, 16'd5898, 16'd14953, 16'd44719, 16'd50260, 16'd53887, 16'd33622, 16'd25165, 16'd29791, 16'd24534, 16'd16653, 16'd64799, 16'd35761, 16'd23140, 16'd22731});
	test_expansion(128'he47684f5055704167540ff1ad93b7c33, {16'd24808, 16'd34747, 16'd31245, 16'd28739, 16'd13345, 16'd35850, 16'd23616, 16'd38641, 16'd30906, 16'd48369, 16'd63520, 16'd29650, 16'd33918, 16'd27573, 16'd49448, 16'd45421, 16'd55924, 16'd9092, 16'd55646, 16'd37953, 16'd45257, 16'd13528, 16'd24442, 16'd61867, 16'd59696, 16'd27860});
	test_expansion(128'h32723838d8ee188a92864d88571084f2, {16'd54770, 16'd35942, 16'd42266, 16'd37350, 16'd24470, 16'd49491, 16'd3238, 16'd2560, 16'd44392, 16'd29782, 16'd53660, 16'd37057, 16'd8745, 16'd40973, 16'd45449, 16'd45012, 16'd64388, 16'd8804, 16'd61404, 16'd60643, 16'd16152, 16'd56748, 16'd43572, 16'd63324, 16'd35079, 16'd37348});
	test_expansion(128'h9dc498a6cb62aa1fc0e7a4e822cd4583, {16'd33265, 16'd19817, 16'd48842, 16'd40045, 16'd15605, 16'd17451, 16'd57456, 16'd12300, 16'd36415, 16'd29941, 16'd26421, 16'd39140, 16'd58915, 16'd23206, 16'd44806, 16'd8221, 16'd12103, 16'd55626, 16'd30952, 16'd47435, 16'd60980, 16'd25580, 16'd27866, 16'd9436, 16'd13905, 16'd65318});
	test_expansion(128'hc3c40d274a130efc4daaf623b85b400d, {16'd53800, 16'd38273, 16'd58557, 16'd51797, 16'd12032, 16'd46151, 16'd62340, 16'd28065, 16'd31272, 16'd63984, 16'd21066, 16'd16356, 16'd5644, 16'd11214, 16'd48462, 16'd27662, 16'd52565, 16'd24543, 16'd9008, 16'd15204, 16'd62185, 16'd40054, 16'd55444, 16'd17728, 16'd38400, 16'd13688});
	test_expansion(128'ha4e6a2e1620d8351ba3baa15152d06b0, {16'd28863, 16'd64986, 16'd32576, 16'd17528, 16'd51068, 16'd14976, 16'd13926, 16'd49962, 16'd20314, 16'd9790, 16'd39046, 16'd51292, 16'd27426, 16'd22006, 16'd56247, 16'd43676, 16'd12871, 16'd61139, 16'd17695, 16'd30614, 16'd7594, 16'd20733, 16'd24080, 16'd3396, 16'd49445, 16'd11553});
	test_expansion(128'haadafbbfb1e23dfb4b1b74ea23b50f94, {16'd1222, 16'd36021, 16'd6791, 16'd15242, 16'd2043, 16'd55810, 16'd55714, 16'd3840, 16'd5499, 16'd16325, 16'd36127, 16'd57475, 16'd41425, 16'd48196, 16'd53816, 16'd40380, 16'd7226, 16'd65074, 16'd15779, 16'd32219, 16'd53550, 16'd17812, 16'd60544, 16'd31271, 16'd34953, 16'd12777});
	test_expansion(128'h19a888de54b4e61d7238ca2582cc9232, {16'd51203, 16'd42569, 16'd37788, 16'd49487, 16'd57035, 16'd24627, 16'd402, 16'd30223, 16'd38923, 16'd47287, 16'd60741, 16'd18603, 16'd11350, 16'd53272, 16'd10113, 16'd10604, 16'd15688, 16'd28424, 16'd49731, 16'd13663, 16'd18560, 16'd6891, 16'd13797, 16'd39796, 16'd48167, 16'd52263});
	test_expansion(128'heb4d572d1d1aa297b1c32ec55c500600, {16'd44773, 16'd64855, 16'd44428, 16'd25464, 16'd40509, 16'd23444, 16'd16087, 16'd27352, 16'd5254, 16'd1402, 16'd16641, 16'd46577, 16'd62990, 16'd64726, 16'd14553, 16'd61380, 16'd56996, 16'd13934, 16'd56880, 16'd41867, 16'd62456, 16'd17421, 16'd60325, 16'd36487, 16'd41444, 16'd28278});
	test_expansion(128'h08e98703b40c1c7c522da2b821cca219, {16'd64074, 16'd58051, 16'd43174, 16'd64727, 16'd52682, 16'd9957, 16'd19263, 16'd27072, 16'd42710, 16'd58969, 16'd46880, 16'd62204, 16'd62786, 16'd40988, 16'd36283, 16'd18696, 16'd24225, 16'd7164, 16'd58916, 16'd43018, 16'd2050, 16'd39943, 16'd50401, 16'd26317, 16'd8951, 16'd44550});
	test_expansion(128'h063717995d1f6eaec63c13f2b0e59ae2, {16'd54641, 16'd41963, 16'd65468, 16'd50394, 16'd44582, 16'd40461, 16'd20314, 16'd52018, 16'd17006, 16'd63739, 16'd5260, 16'd51074, 16'd64551, 16'd10561, 16'd8560, 16'd5250, 16'd28324, 16'd22599, 16'd2622, 16'd10593, 16'd37867, 16'd65465, 16'd43625, 16'd24070, 16'd27746, 16'd19974});
	test_expansion(128'hc6395e4088c3c51b9d821a32380e95a3, {16'd39790, 16'd13625, 16'd55884, 16'd53279, 16'd33758, 16'd39581, 16'd21502, 16'd24773, 16'd7659, 16'd23854, 16'd41970, 16'd47586, 16'd5775, 16'd21193, 16'd33405, 16'd24546, 16'd3474, 16'd42602, 16'd32932, 16'd59543, 16'd48519, 16'd18177, 16'd36965, 16'd14602, 16'd37440, 16'd21412});
	test_expansion(128'hfb11f90a3f45ca99f469ed8bd29a6f26, {16'd64991, 16'd42435, 16'd24111, 16'd1536, 16'd35613, 16'd60627, 16'd6173, 16'd19499, 16'd35648, 16'd51093, 16'd19399, 16'd52098, 16'd56431, 16'd28061, 16'd3330, 16'd37958, 16'd46182, 16'd15422, 16'd27638, 16'd14693, 16'd48469, 16'd54181, 16'd58081, 16'd10119, 16'd39454, 16'd57975});
	test_expansion(128'h3f2f8ba5b154194c59348fce5bc895dd, {16'd34293, 16'd23950, 16'd44378, 16'd20552, 16'd7121, 16'd47492, 16'd10648, 16'd24989, 16'd21552, 16'd44555, 16'd55459, 16'd9540, 16'd7032, 16'd45044, 16'd21680, 16'd31529, 16'd33986, 16'd8375, 16'd36539, 16'd48440, 16'd60299, 16'd42091, 16'd31256, 16'd53637, 16'd1416, 16'd55809});
	test_expansion(128'h129180e1414ca16c28c1b582596ddca8, {16'd63911, 16'd7609, 16'd64800, 16'd41169, 16'd31046, 16'd40740, 16'd31964, 16'd22710, 16'd49100, 16'd48511, 16'd51442, 16'd40331, 16'd19624, 16'd48259, 16'd23335, 16'd32578, 16'd46586, 16'd11348, 16'd16083, 16'd53439, 16'd17032, 16'd40025, 16'd6466, 16'd62556, 16'd22488, 16'd49902});
	test_expansion(128'h1d7754fa4c315d3a93eec246aabb44ef, {16'd5409, 16'd15988, 16'd59072, 16'd24532, 16'd34133, 16'd24721, 16'd4963, 16'd43979, 16'd36738, 16'd55940, 16'd22263, 16'd55135, 16'd35608, 16'd19849, 16'd47180, 16'd28977, 16'd43097, 16'd39625, 16'd7824, 16'd23563, 16'd10536, 16'd2912, 16'd15803, 16'd12531, 16'd50553, 16'd5338});
	test_expansion(128'h7bcb4a516ab13184fb4dd2a60ecb87e1, {16'd23763, 16'd46566, 16'd6461, 16'd31420, 16'd60478, 16'd2648, 16'd27749, 16'd4787, 16'd15535, 16'd4287, 16'd7367, 16'd19778, 16'd60387, 16'd33737, 16'd32167, 16'd57510, 16'd13257, 16'd7634, 16'd53757, 16'd58876, 16'd5529, 16'd16822, 16'd31383, 16'd4033, 16'd24475, 16'd56057});
	test_expansion(128'hb5f3689112a1f0fb42a4b2e445dc85a9, {16'd47303, 16'd43919, 16'd65309, 16'd25470, 16'd28574, 16'd33702, 16'd27612, 16'd24994, 16'd23936, 16'd30650, 16'd22735, 16'd64310, 16'd10662, 16'd32733, 16'd4285, 16'd31612, 16'd23114, 16'd18236, 16'd22640, 16'd47198, 16'd2501, 16'd38764, 16'd59948, 16'd29031, 16'd31980, 16'd58519});
	test_expansion(128'ha11ff0b5bbb8f265d1f9b3ebf40666b7, {16'd35452, 16'd38844, 16'd27138, 16'd9295, 16'd35979, 16'd5482, 16'd38555, 16'd44580, 16'd61026, 16'd33376, 16'd18864, 16'd30367, 16'd18807, 16'd21974, 16'd27418, 16'd64866, 16'd36990, 16'd46188, 16'd52452, 16'd56998, 16'd61247, 16'd13207, 16'd2584, 16'd15262, 16'd26698, 16'd8198});
	test_expansion(128'h21c95b4af73b1031b3e237f29c984cb9, {16'd47579, 16'd65333, 16'd57015, 16'd31104, 16'd12825, 16'd16103, 16'd60048, 16'd52988, 16'd24121, 16'd21156, 16'd1963, 16'd12837, 16'd60100, 16'd60395, 16'd24921, 16'd58798, 16'd59088, 16'd60341, 16'd44612, 16'd2537, 16'd29667, 16'd37311, 16'd53149, 16'd48169, 16'd59234, 16'd62344});
	test_expansion(128'ha9d95ee3ba2b8551c48b01596f7e64a2, {16'd17109, 16'd59937, 16'd20403, 16'd57962, 16'd12528, 16'd8511, 16'd22025, 16'd17256, 16'd44611, 16'd6013, 16'd44303, 16'd63865, 16'd57210, 16'd58540, 16'd3793, 16'd29451, 16'd17997, 16'd2011, 16'd48724, 16'd6697, 16'd55510, 16'd42914, 16'd2279, 16'd22540, 16'd35401, 16'd13871});
	test_expansion(128'h4db7c2d6c97da7fa7473b73d4c9d86a7, {16'd41335, 16'd17471, 16'd60478, 16'd64386, 16'd28504, 16'd29402, 16'd15904, 16'd40873, 16'd26361, 16'd9361, 16'd20229, 16'd64727, 16'd23764, 16'd46242, 16'd6843, 16'd43019, 16'd11822, 16'd25976, 16'd9743, 16'd18468, 16'd47878, 16'd34482, 16'd3094, 16'd5641, 16'd49061, 16'd59016});
	test_expansion(128'h69e349ec9463848c7e92d2232d21b1d3, {16'd5060, 16'd49506, 16'd21453, 16'd27229, 16'd6804, 16'd58715, 16'd35584, 16'd38454, 16'd54995, 16'd7164, 16'd23648, 16'd53965, 16'd523, 16'd26679, 16'd9956, 16'd31899, 16'd59015, 16'd17784, 16'd1677, 16'd666, 16'd62466, 16'd51677, 16'd2203, 16'd51247, 16'd37317, 16'd35901});
	test_expansion(128'he22268bb3d17cc25b59d8db1cee51eef, {16'd8359, 16'd4283, 16'd17719, 16'd36059, 16'd63423, 16'd53174, 16'd31547, 16'd49246, 16'd62921, 16'd21952, 16'd20143, 16'd5193, 16'd11662, 16'd51470, 16'd23315, 16'd6668, 16'd58866, 16'd33427, 16'd26987, 16'd52278, 16'd45873, 16'd17017, 16'd43885, 16'd30361, 16'd12120, 16'd28491});
	test_expansion(128'hcdff1c4a613ebbd8908833705497300a, {16'd41541, 16'd33605, 16'd47745, 16'd62902, 16'd22703, 16'd24281, 16'd27556, 16'd6489, 16'd29253, 16'd49142, 16'd57165, 16'd39392, 16'd10531, 16'd15674, 16'd20723, 16'd32416, 16'd572, 16'd43455, 16'd60757, 16'd6848, 16'd20588, 16'd19925, 16'd57327, 16'd3742, 16'd25350, 16'd20151});
	test_expansion(128'h105f1b1a8e383894f8c2438be5630d88, {16'd18333, 16'd58587, 16'd63137, 16'd34176, 16'd37163, 16'd44712, 16'd29028, 16'd31194, 16'd63993, 16'd18236, 16'd23107, 16'd3265, 16'd22415, 16'd61117, 16'd60326, 16'd44396, 16'd12758, 16'd48650, 16'd31186, 16'd53220, 16'd47943, 16'd21096, 16'd56169, 16'd54908, 16'd62915, 16'd34887});
	test_expansion(128'he15a166dffe3c0effc65000af15fd1c1, {16'd19378, 16'd41465, 16'd24811, 16'd64609, 16'd28272, 16'd24796, 16'd40393, 16'd56997, 16'd11646, 16'd48127, 16'd58240, 16'd46303, 16'd21135, 16'd43719, 16'd46043, 16'd21488, 16'd10189, 16'd62188, 16'd50982, 16'd23375, 16'd26968, 16'd1712, 16'd27797, 16'd49525, 16'd63089, 16'd19898});
	test_expansion(128'hed1584e2ffd638b1961c3e099c03106e, {16'd4846, 16'd32849, 16'd3211, 16'd41840, 16'd564, 16'd26564, 16'd17956, 16'd63239, 16'd40251, 16'd59639, 16'd25583, 16'd47879, 16'd30535, 16'd33583, 16'd62572, 16'd40913, 16'd48739, 16'd52463, 16'd18893, 16'd6982, 16'd40178, 16'd54099, 16'd18031, 16'd41385, 16'd43430, 16'd58979});
	test_expansion(128'h675912f3c55f88458c2be018f98f1b77, {16'd5670, 16'd23564, 16'd8214, 16'd21626, 16'd55382, 16'd1312, 16'd1549, 16'd50731, 16'd65424, 16'd36778, 16'd25874, 16'd51367, 16'd53501, 16'd7110, 16'd42142, 16'd32162, 16'd9030, 16'd58054, 16'd21593, 16'd38825, 16'd38124, 16'd37464, 16'd15465, 16'd41034, 16'd43923, 16'd23429});
	test_expansion(128'hc6cd06cb6b994d510a0aa13a7a612fd7, {16'd23144, 16'd24167, 16'd42452, 16'd39008, 16'd5250, 16'd28555, 16'd21841, 16'd38188, 16'd21640, 16'd12433, 16'd58703, 16'd59254, 16'd30965, 16'd23429, 16'd62782, 16'd49102, 16'd54821, 16'd55076, 16'd24534, 16'd21650, 16'd7520, 16'd13118, 16'd21241, 16'd56693, 16'd43159, 16'd52611});
	test_expansion(128'h95cc49260d76a72b65b1855045858f36, {16'd4968, 16'd28760, 16'd620, 16'd924, 16'd500, 16'd48327, 16'd25973, 16'd8466, 16'd40171, 16'd5830, 16'd15324, 16'd63248, 16'd41256, 16'd8235, 16'd969, 16'd51357, 16'd22034, 16'd64030, 16'd44098, 16'd23790, 16'd14911, 16'd14882, 16'd16490, 16'd22548, 16'd36779, 16'd40765});
	test_expansion(128'h20ac3c7dc752519ef385412f907b0b09, {16'd44447, 16'd59198, 16'd8856, 16'd30717, 16'd28973, 16'd62339, 16'd40912, 16'd9450, 16'd47205, 16'd598, 16'd63846, 16'd7764, 16'd26918, 16'd22358, 16'd61352, 16'd11044, 16'd46821, 16'd38037, 16'd45639, 16'd1792, 16'd62311, 16'd13532, 16'd29035, 16'd28302, 16'd22180, 16'd37439});
	test_expansion(128'h9be27b006b87cdaf5e54322b81855b29, {16'd29842, 16'd38180, 16'd30816, 16'd26769, 16'd5883, 16'd57669, 16'd24432, 16'd20113, 16'd18935, 16'd54358, 16'd18404, 16'd20313, 16'd35212, 16'd31019, 16'd38416, 16'd30234, 16'd14105, 16'd48839, 16'd49783, 16'd51282, 16'd45444, 16'd3639, 16'd22990, 16'd18357, 16'd13552, 16'd48003});
	test_expansion(128'h75f2a58b22d21e6e21ab4a7e36830c1e, {16'd59222, 16'd9464, 16'd6413, 16'd25873, 16'd45158, 16'd49313, 16'd46540, 16'd21635, 16'd34933, 16'd15686, 16'd53785, 16'd55252, 16'd59898, 16'd46569, 16'd14180, 16'd30480, 16'd7916, 16'd12809, 16'd12117, 16'd33122, 16'd28894, 16'd18668, 16'd52609, 16'd11143, 16'd57273, 16'd10934});
	test_expansion(128'h90b84c7e8eecf01abb78778502ff02a0, {16'd50843, 16'd59735, 16'd19100, 16'd22981, 16'd13730, 16'd65483, 16'd15246, 16'd20352, 16'd14710, 16'd36368, 16'd39018, 16'd14337, 16'd30879, 16'd38893, 16'd24500, 16'd51435, 16'd63932, 16'd46420, 16'd37172, 16'd134, 16'd18194, 16'd16202, 16'd46983, 16'd44542, 16'd15992, 16'd23115});
	test_expansion(128'hb5c2526b89e2e792e5246b70e13b7d97, {16'd59008, 16'd26488, 16'd21538, 16'd7750, 16'd12016, 16'd38149, 16'd50969, 16'd57499, 16'd46524, 16'd54389, 16'd1791, 16'd51928, 16'd915, 16'd41592, 16'd48052, 16'd33571, 16'd12866, 16'd49848, 16'd36612, 16'd37952, 16'd55389, 16'd33905, 16'd52576, 16'd46540, 16'd739, 16'd44895});
	test_expansion(128'hd8d95c019448519713072f68f45bdc05, {16'd3214, 16'd44660, 16'd17487, 16'd31977, 16'd35703, 16'd57327, 16'd53100, 16'd65338, 16'd24383, 16'd44076, 16'd24747, 16'd55586, 16'd31228, 16'd5644, 16'd58019, 16'd57416, 16'd10371, 16'd961, 16'd51521, 16'd49048, 16'd11099, 16'd7004, 16'd20661, 16'd49647, 16'd35609, 16'd57231});
	test_expansion(128'hf4a89f55f032a95bf450e682d34c1963, {16'd5586, 16'd16785, 16'd14809, 16'd20770, 16'd59965, 16'd13311, 16'd55322, 16'd21474, 16'd40235, 16'd20401, 16'd30239, 16'd52636, 16'd28942, 16'd16957, 16'd31628, 16'd57281, 16'd41024, 16'd10806, 16'd14070, 16'd30546, 16'd42757, 16'd5549, 16'd63149, 16'd5564, 16'd10837, 16'd399});
	test_expansion(128'h7c1feb6c3421856ac7d021d302411b41, {16'd7589, 16'd16426, 16'd62137, 16'd41075, 16'd29394, 16'd38875, 16'd13864, 16'd614, 16'd27811, 16'd61556, 16'd30217, 16'd1620, 16'd37083, 16'd26634, 16'd24066, 16'd3388, 16'd87, 16'd19203, 16'd41514, 16'd58956, 16'd17288, 16'd57309, 16'd42125, 16'd63830, 16'd52346, 16'd20809});
	test_expansion(128'ha1774564a12e767d291e4cc43eaa2f8c, {16'd59214, 16'd18498, 16'd17884, 16'd44916, 16'd14851, 16'd15565, 16'd28299, 16'd7894, 16'd55986, 16'd55604, 16'd11494, 16'd17168, 16'd51265, 16'd8843, 16'd22087, 16'd17839, 16'd53087, 16'd27392, 16'd37001, 16'd33458, 16'd9294, 16'd4202, 16'd37626, 16'd60927, 16'd34855, 16'd38169});
	test_expansion(128'hb3b0d979e907d55cb9a32a86f4a9c655, {16'd35915, 16'd20282, 16'd50994, 16'd57115, 16'd31042, 16'd19402, 16'd2258, 16'd25098, 16'd59993, 16'd11043, 16'd44228, 16'd28404, 16'd16432, 16'd39054, 16'd25798, 16'd7970, 16'd58693, 16'd61838, 16'd40604, 16'd6769, 16'd29182, 16'd33965, 16'd50490, 16'd26279, 16'd43551, 16'd42394});
	test_expansion(128'h3eb58dcde9d181345dcbcb8dd4e86291, {16'd24861, 16'd40424, 16'd31511, 16'd62459, 16'd56637, 16'd26061, 16'd35695, 16'd17749, 16'd51217, 16'd57540, 16'd5109, 16'd54557, 16'd13317, 16'd33611, 16'd63238, 16'd45898, 16'd30443, 16'd36133, 16'd15561, 16'd48282, 16'd10001, 16'd28490, 16'd58000, 16'd3332, 16'd58750, 16'd22100});
	test_expansion(128'hb9e35cab48441ed3d428cf61bb7ee527, {16'd9498, 16'd18237, 16'd33841, 16'd1936, 16'd2779, 16'd27559, 16'd23087, 16'd44960, 16'd64730, 16'd44727, 16'd58751, 16'd64699, 16'd5271, 16'd62036, 16'd63380, 16'd19486, 16'd34527, 16'd56000, 16'd18911, 16'd20557, 16'd1160, 16'd36349, 16'd60597, 16'd60619, 16'd41891, 16'd55847});
	test_expansion(128'h216057a4f2d3868cab5587398b727f96, {16'd47709, 16'd37907, 16'd42629, 16'd3404, 16'd42889, 16'd62886, 16'd41592, 16'd45283, 16'd1656, 16'd40887, 16'd19182, 16'd8231, 16'd22421, 16'd15203, 16'd25187, 16'd58964, 16'd16995, 16'd16676, 16'd43616, 16'd10636, 16'd57319, 16'd54766, 16'd4935, 16'd7384, 16'd34460, 16'd47375});
	test_expansion(128'hef529e04ea69b4cce56ba9a670a6cc3e, {16'd43709, 16'd63311, 16'd29140, 16'd25004, 16'd18888, 16'd5677, 16'd36858, 16'd59633, 16'd77, 16'd55064, 16'd32517, 16'd26693, 16'd59370, 16'd45364, 16'd47196, 16'd51873, 16'd41984, 16'd15745, 16'd2248, 16'd8930, 16'd3028, 16'd23688, 16'd55863, 16'd1613, 16'd27750, 16'd64103});
	test_expansion(128'hb7fc1e9a311e0f539d53d56f3fc96a6d, {16'd38529, 16'd57853, 16'd49584, 16'd39010, 16'd50205, 16'd64662, 16'd59341, 16'd57358, 16'd27616, 16'd24492, 16'd27606, 16'd43579, 16'd3316, 16'd25585, 16'd46072, 16'd44515, 16'd41309, 16'd62908, 16'd41186, 16'd10171, 16'd27406, 16'd32420, 16'd111, 16'd22838, 16'd46748, 16'd6221});
	test_expansion(128'h21850b1a937e93842d0550af72dde5df, {16'd47034, 16'd61867, 16'd17232, 16'd40933, 16'd52128, 16'd46326, 16'd61903, 16'd58291, 16'd21123, 16'd32083, 16'd33658, 16'd485, 16'd61759, 16'd2691, 16'd6927, 16'd22674, 16'd25576, 16'd50824, 16'd16444, 16'd37553, 16'd54264, 16'd6399, 16'd59469, 16'd30930, 16'd25226, 16'd16136});
	test_expansion(128'h570a47b0f451e9705403e957f36a841b, {16'd55856, 16'd36258, 16'd51520, 16'd25434, 16'd3621, 16'd52985, 16'd48013, 16'd59270, 16'd29845, 16'd36579, 16'd10043, 16'd17293, 16'd4390, 16'd57762, 16'd27115, 16'd32391, 16'd46714, 16'd35047, 16'd22040, 16'd36972, 16'd45096, 16'd51650, 16'd18188, 16'd15623, 16'd27349, 16'd1549});
	test_expansion(128'h87990a0d2c040751f065c3f57dccfbbf, {16'd18102, 16'd47554, 16'd12023, 16'd2219, 16'd60361, 16'd2334, 16'd61986, 16'd3799, 16'd54080, 16'd27251, 16'd57189, 16'd57483, 16'd38346, 16'd41761, 16'd414, 16'd23063, 16'd8811, 16'd12625, 16'd32990, 16'd29445, 16'd48076, 16'd55267, 16'd36530, 16'd39993, 16'd56939, 16'd33721});
	test_expansion(128'h6d515c8fb03deb52dad52ac0485e8cd4, {16'd64566, 16'd19282, 16'd53279, 16'd59780, 16'd25178, 16'd62250, 16'd49161, 16'd12003, 16'd5798, 16'd55612, 16'd3788, 16'd645, 16'd37262, 16'd16660, 16'd25629, 16'd4355, 16'd15950, 16'd60782, 16'd57078, 16'd15989, 16'd10642, 16'd43716, 16'd9976, 16'd28897, 16'd47081, 16'd49794});
	test_expansion(128'hbfff0d2f2be63e3769cd106dd96ce2ca, {16'd41531, 16'd50989, 16'd48829, 16'd63716, 16'd38854, 16'd38652, 16'd60813, 16'd23360, 16'd1620, 16'd39950, 16'd35213, 16'd36570, 16'd25738, 16'd27903, 16'd28041, 16'd12803, 16'd41170, 16'd24849, 16'd49766, 16'd64853, 16'd49788, 16'd4532, 16'd1075, 16'd596, 16'd11355, 16'd10101});
	test_expansion(128'h99b6407f839f3e44144fc487f87e0a75, {16'd25371, 16'd37228, 16'd26851, 16'd65443, 16'd42814, 16'd62079, 16'd51471, 16'd10863, 16'd60085, 16'd837, 16'd23914, 16'd29533, 16'd53463, 16'd56393, 16'd21598, 16'd47339, 16'd40603, 16'd40205, 16'd20914, 16'd50707, 16'd46489, 16'd44758, 16'd17269, 16'd35586, 16'd39166, 16'd1271});
	test_expansion(128'h0483ccdad222e339510bc7081c7e0fc9, {16'd44920, 16'd49941, 16'd45480, 16'd44634, 16'd55561, 16'd6454, 16'd20980, 16'd65475, 16'd46532, 16'd44422, 16'd8706, 16'd31097, 16'd37107, 16'd63882, 16'd37187, 16'd44093, 16'd44855, 16'd44903, 16'd27872, 16'd29378, 16'd28423, 16'd29243, 16'd30864, 16'd36917, 16'd41310, 16'd65249});
	test_expansion(128'h4d7fb832d4b72b36a65740b86d2c7dbb, {16'd10358, 16'd17873, 16'd31404, 16'd52073, 16'd48964, 16'd50503, 16'd37098, 16'd39095, 16'd52368, 16'd52026, 16'd24718, 16'd4229, 16'd53562, 16'd58139, 16'd48324, 16'd11451, 16'd10567, 16'd34213, 16'd31009, 16'd50379, 16'd62200, 16'd51746, 16'd21487, 16'd18650, 16'd39736, 16'd9406});
	test_expansion(128'h9a3607c12d5836d8d6d03e18f44ecaa1, {16'd8245, 16'd49795, 16'd59048, 16'd21317, 16'd32626, 16'd53979, 16'd3345, 16'd50668, 16'd42778, 16'd44831, 16'd21451, 16'd24386, 16'd20400, 16'd39245, 16'd51229, 16'd42432, 16'd23246, 16'd45989, 16'd53956, 16'd50055, 16'd24759, 16'd39481, 16'd60407, 16'd50306, 16'd10953, 16'd33665});
	test_expansion(128'h6c5a3f0acb2ec3c8ff03586d3ae2024a, {16'd22753, 16'd30776, 16'd17636, 16'd5674, 16'd52651, 16'd58431, 16'd47875, 16'd43417, 16'd35586, 16'd20973, 16'd57181, 16'd50879, 16'd26920, 16'd60162, 16'd45047, 16'd856, 16'd26344, 16'd58008, 16'd33881, 16'd35387, 16'd53422, 16'd63496, 16'd19261, 16'd22831, 16'd62468, 16'd44728});
	test_expansion(128'he4d2c1278031b06ea984edb6080beba5, {16'd63700, 16'd48870, 16'd13423, 16'd41497, 16'd24151, 16'd19258, 16'd55933, 16'd10179, 16'd17724, 16'd27317, 16'd52547, 16'd24323, 16'd58408, 16'd27269, 16'd52890, 16'd2970, 16'd61227, 16'd19467, 16'd4912, 16'd21879, 16'd44986, 16'd467, 16'd15819, 16'd14990, 16'd41983, 16'd20795});
	test_expansion(128'h2bb6330aae144951e48354d88859a787, {16'd2880, 16'd29006, 16'd63655, 16'd4309, 16'd49015, 16'd22460, 16'd56060, 16'd24512, 16'd5794, 16'd24094, 16'd37215, 16'd55266, 16'd26686, 16'd16670, 16'd61711, 16'd13257, 16'd32204, 16'd42348, 16'd46571, 16'd7581, 16'd46458, 16'd34518, 16'd24666, 16'd45916, 16'd63927, 16'd23297});
	test_expansion(128'hba6750824e829a99ffd8e40759bf185a, {16'd3639, 16'd58075, 16'd49892, 16'd54940, 16'd65169, 16'd51145, 16'd9816, 16'd49320, 16'd2158, 16'd45947, 16'd56089, 16'd59518, 16'd34534, 16'd42079, 16'd45030, 16'd9995, 16'd7332, 16'd13104, 16'd29560, 16'd8796, 16'd55390, 16'd5684, 16'd13628, 16'd45769, 16'd36855, 16'd40607});
	test_expansion(128'h1a545a36071f5fc8b3852b3c6244730d, {16'd29049, 16'd1361, 16'd33431, 16'd46459, 16'd4975, 16'd56018, 16'd34648, 16'd32519, 16'd39266, 16'd18843, 16'd55865, 16'd19306, 16'd1225, 16'd48824, 16'd10974, 16'd45170, 16'd34470, 16'd37627, 16'd63063, 16'd37455, 16'd655, 16'd44620, 16'd11738, 16'd50612, 16'd29027, 16'd48968});
	test_expansion(128'h347207d96d3f5e48dc1fcb2e389e8152, {16'd35144, 16'd14371, 16'd10943, 16'd887, 16'd1176, 16'd41897, 16'd19061, 16'd27914, 16'd41792, 16'd3122, 16'd49021, 16'd22927, 16'd26940, 16'd60670, 16'd11559, 16'd28005, 16'd44560, 16'd51193, 16'd27755, 16'd58224, 16'd34009, 16'd37785, 16'd35840, 16'd18302, 16'd12510, 16'd442});
	test_expansion(128'h4232f0a167b21b7e6c9a17a14651e2b7, {16'd50113, 16'd62739, 16'd54415, 16'd39723, 16'd16657, 16'd51155, 16'd7035, 16'd24139, 16'd28067, 16'd60056, 16'd34573, 16'd49443, 16'd1200, 16'd36244, 16'd19028, 16'd40348, 16'd21246, 16'd11399, 16'd29514, 16'd61236, 16'd49531, 16'd3740, 16'd32111, 16'd52623, 16'd33319, 16'd31275});
	test_expansion(128'h6bf0fb7b186651be9a5f0d16dea285ac, {16'd23280, 16'd4186, 16'd36168, 16'd33750, 16'd58151, 16'd16758, 16'd19281, 16'd11566, 16'd21673, 16'd58074, 16'd9894, 16'd9740, 16'd12726, 16'd13213, 16'd28153, 16'd57834, 16'd55975, 16'd62333, 16'd17929, 16'd40975, 16'd60264, 16'd25801, 16'd17221, 16'd57183, 16'd42417, 16'd42327});
	test_expansion(128'h68df387e8f4e5d8dcef60de90bcb911f, {16'd14714, 16'd22086, 16'd8525, 16'd22796, 16'd22493, 16'd4363, 16'd59770, 16'd9526, 16'd48579, 16'd51216, 16'd57855, 16'd4861, 16'd65315, 16'd12645, 16'd52188, 16'd40979, 16'd35450, 16'd18052, 16'd4549, 16'd61064, 16'd53638, 16'd54339, 16'd29655, 16'd42631, 16'd26918, 16'd16789});
	test_expansion(128'hdf26b4c614252479882302fd2d341933, {16'd13886, 16'd12565, 16'd31582, 16'd49505, 16'd10599, 16'd52613, 16'd30670, 16'd35822, 16'd23295, 16'd49217, 16'd42059, 16'd18200, 16'd60750, 16'd14760, 16'd11251, 16'd39826, 16'd6226, 16'd57256, 16'd50677, 16'd55703, 16'd5266, 16'd25331, 16'd10967, 16'd1171, 16'd11985, 16'd40286});
	test_expansion(128'h364fdb4098f9a4fad536a51cb192eea3, {16'd38914, 16'd21911, 16'd18642, 16'd58890, 16'd49485, 16'd33448, 16'd21180, 16'd39244, 16'd54602, 16'd61649, 16'd47522, 16'd56342, 16'd43425, 16'd8643, 16'd38155, 16'd41466, 16'd30525, 16'd45716, 16'd18737, 16'd30048, 16'd29927, 16'd31522, 16'd20279, 16'd18721, 16'd38283, 16'd17680});
	test_expansion(128'h9735e3ec19b760b977811ce5cbb17d0e, {16'd4150, 16'd33095, 16'd37958, 16'd11927, 16'd50698, 16'd45709, 16'd2581, 16'd1730, 16'd4528, 16'd14092, 16'd58150, 16'd56871, 16'd23245, 16'd50880, 16'd26005, 16'd54724, 16'd60805, 16'd62182, 16'd58386, 16'd15390, 16'd18328, 16'd65357, 16'd26926, 16'd50309, 16'd40605, 16'd61808});
	test_expansion(128'h1c90539590bddba5b5140c8db2b7b9df, {16'd54979, 16'd16965, 16'd27580, 16'd15352, 16'd15205, 16'd23533, 16'd20541, 16'd17409, 16'd31363, 16'd31586, 16'd1534, 16'd46311, 16'd61216, 16'd58660, 16'd15889, 16'd51734, 16'd63076, 16'd38091, 16'd14823, 16'd899, 16'd37905, 16'd565, 16'd8087, 16'd32346, 16'd56976, 16'd56869});
	test_expansion(128'h6dacb94765ffb5d5eca84acb7f522c03, {16'd51911, 16'd21921, 16'd363, 16'd12203, 16'd20789, 16'd34467, 16'd12488, 16'd29703, 16'd40855, 16'd6045, 16'd47970, 16'd64067, 16'd50207, 16'd48063, 16'd4967, 16'd43322, 16'd14450, 16'd7707, 16'd30959, 16'd44466, 16'd49037, 16'd40120, 16'd21736, 16'd17562, 16'd53546, 16'd26347});
	test_expansion(128'hcf17d7652c30d8aec49fb8b6d55dea5a, {16'd39848, 16'd1923, 16'd14865, 16'd38266, 16'd41563, 16'd28011, 16'd37566, 16'd13176, 16'd59183, 16'd48374, 16'd11009, 16'd53243, 16'd47319, 16'd37867, 16'd37247, 16'd45685, 16'd4040, 16'd29735, 16'd38809, 16'd61714, 16'd3003, 16'd37055, 16'd8490, 16'd13619, 16'd46927, 16'd20694});
	test_expansion(128'h362ca52e985691b3cb8054f01b0d50a9, {16'd47544, 16'd11399, 16'd55589, 16'd32598, 16'd48569, 16'd41838, 16'd33265, 16'd52728, 16'd44250, 16'd34809, 16'd9616, 16'd7744, 16'd63642, 16'd55185, 16'd4533, 16'd7745, 16'd36241, 16'd3454, 16'd19146, 16'd1095, 16'd58010, 16'd50791, 16'd48368, 16'd10803, 16'd25008, 16'd43858});
	test_expansion(128'h70d382f74edd6e698fdaf8903482ae4d, {16'd42377, 16'd22998, 16'd60438, 16'd31963, 16'd64739, 16'd31886, 16'd57078, 16'd49257, 16'd63850, 16'd58002, 16'd46902, 16'd38179, 16'd31778, 16'd4834, 16'd51323, 16'd107, 16'd41944, 16'd21702, 16'd25845, 16'd15472, 16'd10920, 16'd14240, 16'd7262, 16'd31001, 16'd43021, 16'd33902});
	test_expansion(128'hcc918ea89c9fc04f8e8989a4df7a3cc2, {16'd7063, 16'd57700, 16'd45263, 16'd29309, 16'd47044, 16'd54127, 16'd63733, 16'd20938, 16'd37050, 16'd38607, 16'd21303, 16'd57905, 16'd11950, 16'd12744, 16'd7818, 16'd30188, 16'd60596, 16'd2472, 16'd7039, 16'd31519, 16'd42124, 16'd9540, 16'd14695, 16'd46770, 16'd18441, 16'd28368});
	test_expansion(128'h500b8619b8f6297f41f8c4996edcd9ad, {16'd2320, 16'd61016, 16'd47458, 16'd23853, 16'd27491, 16'd35065, 16'd61800, 16'd40315, 16'd16574, 16'd29604, 16'd41826, 16'd59567, 16'd61932, 16'd24924, 16'd55025, 16'd53681, 16'd45721, 16'd50234, 16'd57809, 16'd62924, 16'd47028, 16'd24064, 16'd44193, 16'd42927, 16'd11963, 16'd54079});
	test_expansion(128'hec5cb52a5d6e4428c3a42ead134c2214, {16'd19929, 16'd13313, 16'd4310, 16'd35089, 16'd53876, 16'd4556, 16'd40922, 16'd40422, 16'd40154, 16'd11236, 16'd8870, 16'd45909, 16'd28634, 16'd48218, 16'd60993, 16'd59301, 16'd15043, 16'd53141, 16'd45168, 16'd45090, 16'd44624, 16'd37909, 16'd38795, 16'd17842, 16'd34294, 16'd36981});
	test_expansion(128'hd611e4d57d886bec538f79c63a46b797, {16'd42604, 16'd24437, 16'd37895, 16'd40726, 16'd5438, 16'd54750, 16'd7923, 16'd54938, 16'd21762, 16'd16047, 16'd62450, 16'd6362, 16'd58821, 16'd58980, 16'd33866, 16'd62669, 16'd42559, 16'd63018, 16'd13798, 16'd7814, 16'd15132, 16'd19234, 16'd43052, 16'd55536, 16'd36896, 16'd63044});
	test_expansion(128'hbc50de48290e341dbc520082463f077f, {16'd9570, 16'd6551, 16'd5482, 16'd49857, 16'd38861, 16'd55381, 16'd22749, 16'd45803, 16'd57544, 16'd878, 16'd8367, 16'd32778, 16'd45038, 16'd53379, 16'd6227, 16'd39046, 16'd14646, 16'd55966, 16'd26288, 16'd29943, 16'd21607, 16'd49088, 16'd37748, 16'd6863, 16'd13598, 16'd54149});
	test_expansion(128'hefa19de6590fea25ee9178e532b315e0, {16'd52944, 16'd2362, 16'd46965, 16'd14670, 16'd10636, 16'd40394, 16'd46347, 16'd35063, 16'd2158, 16'd43314, 16'd17260, 16'd21218, 16'd183, 16'd7615, 16'd44905, 16'd23390, 16'd28945, 16'd44299, 16'd59066, 16'd53137, 16'd63921, 16'd58164, 16'd60035, 16'd11616, 16'd34525, 16'd25450});
	test_expansion(128'h58cfe2ac85e8f0549dc0ff46c0d93213, {16'd1906, 16'd15316, 16'd40365, 16'd61565, 16'd22322, 16'd21089, 16'd27658, 16'd16320, 16'd30260, 16'd61610, 16'd57330, 16'd12550, 16'd28191, 16'd20052, 16'd50611, 16'd49344, 16'd18424, 16'd30439, 16'd38885, 16'd47736, 16'd40160, 16'd58457, 16'd38392, 16'd6908, 16'd61014, 16'd59472});
	test_expansion(128'h609d56caf04da9315693e6e1a4e2793b, {16'd38700, 16'd19422, 16'd11472, 16'd18865, 16'd30991, 16'd19188, 16'd42119, 16'd31786, 16'd23803, 16'd9351, 16'd43725, 16'd18956, 16'd9153, 16'd63387, 16'd44250, 16'd49624, 16'd31875, 16'd20121, 16'd34491, 16'd11088, 16'd52464, 16'd11443, 16'd22487, 16'd22990, 16'd10314, 16'd44003});
	test_expansion(128'h110a9c16846f68be80921248a67dbc61, {16'd4979, 16'd55739, 16'd42623, 16'd55108, 16'd37828, 16'd8779, 16'd27416, 16'd14571, 16'd48871, 16'd22730, 16'd41111, 16'd65418, 16'd21625, 16'd4296, 16'd5259, 16'd24759, 16'd543, 16'd19378, 16'd24384, 16'd10630, 16'd38545, 16'd36664, 16'd33950, 16'd53207, 16'd25725, 16'd15169});
	test_expansion(128'h4366dff56cec3f4f07e9321340b4ee73, {16'd51425, 16'd65453, 16'd26823, 16'd36345, 16'd41758, 16'd46114, 16'd41113, 16'd59692, 16'd10034, 16'd55498, 16'd38561, 16'd58687, 16'd46059, 16'd35270, 16'd25723, 16'd59901, 16'd38570, 16'd1951, 16'd47454, 16'd43208, 16'd64156, 16'd20442, 16'd52619, 16'd28521, 16'd40551, 16'd36082});
	test_expansion(128'h3e1b7888328dc883d11553305ca05d89, {16'd18819, 16'd55014, 16'd1566, 16'd31789, 16'd43068, 16'd24608, 16'd23322, 16'd59412, 16'd23074, 16'd9808, 16'd14015, 16'd60011, 16'd40406, 16'd16295, 16'd64645, 16'd32497, 16'd38027, 16'd1262, 16'd44009, 16'd53883, 16'd5549, 16'd28813, 16'd50745, 16'd386, 16'd43617, 16'd29594});
	test_expansion(128'h4cb2b1c934c10e9724435a1d7bec8b49, {16'd29237, 16'd40795, 16'd55985, 16'd50793, 16'd63065, 16'd29269, 16'd60691, 16'd38572, 16'd27933, 16'd13470, 16'd52477, 16'd64186, 16'd50511, 16'd12573, 16'd25099, 16'd24830, 16'd25633, 16'd22073, 16'd34738, 16'd16244, 16'd42968, 16'd58937, 16'd46127, 16'd25264, 16'd65463, 16'd7015});
	test_expansion(128'h896d78e2a303b78177cef1ec358c18ea, {16'd60830, 16'd32264, 16'd56184, 16'd14146, 16'd30336, 16'd6808, 16'd15618, 16'd31634, 16'd52125, 16'd9278, 16'd42452, 16'd10743, 16'd59221, 16'd48177, 16'd20767, 16'd20066, 16'd28330, 16'd46334, 16'd53334, 16'd13924, 16'd18217, 16'd61986, 16'd34323, 16'd62980, 16'd46912, 16'd17397});
	test_expansion(128'he0b67ec5da5ad8dd7bf221ae8a852afc, {16'd59336, 16'd54779, 16'd10803, 16'd16846, 16'd46787, 16'd39339, 16'd58482, 16'd39088, 16'd5439, 16'd52112, 16'd20288, 16'd54039, 16'd56063, 16'd13088, 16'd45797, 16'd14190, 16'd37647, 16'd48150, 16'd46267, 16'd32964, 16'd40677, 16'd58834, 16'd54021, 16'd59508, 16'd47945, 16'd25575});
	test_expansion(128'h1e440aa39c9981d92c6e9ad0ffdaa475, {16'd50250, 16'd18245, 16'd22945, 16'd16585, 16'd22842, 16'd8216, 16'd12660, 16'd47815, 16'd51757, 16'd60176, 16'd885, 16'd22172, 16'd16544, 16'd63133, 16'd48128, 16'd34934, 16'd59715, 16'd28481, 16'd41659, 16'd59380, 16'd7286, 16'd33546, 16'd34765, 16'd21706, 16'd40694, 16'd54277});
	test_expansion(128'ha9acd1e6c3a95009bcd9f6942324ae2f, {16'd18383, 16'd6847, 16'd11042, 16'd22625, 16'd47961, 16'd1001, 16'd7070, 16'd27324, 16'd44148, 16'd19194, 16'd57228, 16'd47437, 16'd11346, 16'd53863, 16'd8103, 16'd43285, 16'd18423, 16'd55462, 16'd55790, 16'd26572, 16'd24815, 16'd37578, 16'd4601, 16'd56478, 16'd41297, 16'd61985});
	test_expansion(128'he993d88213d6a07645783476d9359248, {16'd40840, 16'd49890, 16'd2077, 16'd24243, 16'd53944, 16'd59225, 16'd55501, 16'd17337, 16'd64161, 16'd37077, 16'd12029, 16'd51358, 16'd24795, 16'd5357, 16'd33972, 16'd32110, 16'd6705, 16'd45604, 16'd34319, 16'd19162, 16'd48258, 16'd24980, 16'd41177, 16'd50173, 16'd63208, 16'd9204});
	test_expansion(128'h783016695a5f57f6761fa79a612d921b, {16'd55328, 16'd51147, 16'd6392, 16'd37737, 16'd49907, 16'd56838, 16'd40475, 16'd42285, 16'd28090, 16'd25816, 16'd25992, 16'd13839, 16'd19722, 16'd8797, 16'd37635, 16'd58006, 16'd47129, 16'd11099, 16'd17935, 16'd7638, 16'd17600, 16'd23027, 16'd56818, 16'd36452, 16'd61454, 16'd55699});
	test_expansion(128'h0ece14da50a315d7397d24a672effb7e, {16'd63860, 16'd23504, 16'd434, 16'd11723, 16'd62257, 16'd23185, 16'd59277, 16'd58856, 16'd61978, 16'd63221, 16'd28334, 16'd45907, 16'd10786, 16'd61434, 16'd25837, 16'd13658, 16'd33226, 16'd24732, 16'd51643, 16'd40753, 16'd5502, 16'd2481, 16'd10089, 16'd54283, 16'd3842, 16'd4851});
	test_expansion(128'h7e6dbb55a8328cd2516d16f2fabcb05e, {16'd15893, 16'd22102, 16'd44776, 16'd35982, 16'd31982, 16'd10716, 16'd16679, 16'd53190, 16'd52959, 16'd26169, 16'd30453, 16'd30334, 16'd12414, 16'd63219, 16'd17587, 16'd58725, 16'd39528, 16'd12679, 16'd21750, 16'd16891, 16'd42764, 16'd13197, 16'd12462, 16'd47818, 16'd18058, 16'd5957});
	test_expansion(128'hd7f8464bb5fcb0afed4d7675419d1aa2, {16'd53846, 16'd1871, 16'd63776, 16'd11728, 16'd64091, 16'd20581, 16'd9048, 16'd43548, 16'd65298, 16'd4910, 16'd32350, 16'd27791, 16'd26569, 16'd59352, 16'd13534, 16'd54404, 16'd23338, 16'd42452, 16'd54564, 16'd62214, 16'd6149, 16'd60712, 16'd5567, 16'd6209, 16'd57402, 16'd38948});
	test_expansion(128'h7671748c273bcd4fb5a98e01ffa4c0a0, {16'd40283, 16'd21207, 16'd26163, 16'd29996, 16'd26339, 16'd50478, 16'd26456, 16'd30109, 16'd2846, 16'd47344, 16'd23346, 16'd55921, 16'd37661, 16'd23836, 16'd54882, 16'd59855, 16'd27003, 16'd23136, 16'd27949, 16'd48109, 16'd25889, 16'd27758, 16'd52929, 16'd2919, 16'd19885, 16'd64511});
	test_expansion(128'hcea1ddc4ef825947641dac2fef595f96, {16'd7025, 16'd53427, 16'd17741, 16'd61206, 16'd64978, 16'd63834, 16'd57383, 16'd33708, 16'd53421, 16'd13224, 16'd54308, 16'd12866, 16'd65209, 16'd27962, 16'd36711, 16'd32786, 16'd23305, 16'd4885, 16'd57441, 16'd4385, 16'd33975, 16'd38181, 16'd58954, 16'd4295, 16'd54431, 16'd50850});
	test_expansion(128'h65721943be21676ab461cf296a615db5, {16'd19130, 16'd40310, 16'd35446, 16'd1675, 16'd61860, 16'd6387, 16'd2731, 16'd48931, 16'd61499, 16'd54713, 16'd18040, 16'd32367, 16'd19771, 16'd43456, 16'd31862, 16'd27986, 16'd39389, 16'd10038, 16'd1618, 16'd60828, 16'd11736, 16'd4156, 16'd62509, 16'd48949, 16'd46038, 16'd31604});
	test_expansion(128'h64ac103cb53809eb79e4b72459da36f4, {16'd156, 16'd35922, 16'd45868, 16'd42085, 16'd60311, 16'd10579, 16'd37483, 16'd32614, 16'd29631, 16'd64309, 16'd38811, 16'd3745, 16'd50257, 16'd62684, 16'd32021, 16'd46539, 16'd30961, 16'd61512, 16'd42254, 16'd4997, 16'd29366, 16'd11288, 16'd19731, 16'd26333, 16'd45491, 16'd41235});
	test_expansion(128'h376e0e90ece4b709fbcb6512c9dd4ffe, {16'd36944, 16'd49083, 16'd58456, 16'd44267, 16'd40000, 16'd52128, 16'd48436, 16'd5910, 16'd47023, 16'd25215, 16'd27565, 16'd9296, 16'd26722, 16'd52987, 16'd37429, 16'd8671, 16'd42161, 16'd25762, 16'd38499, 16'd34477, 16'd17529, 16'd46441, 16'd18884, 16'd10807, 16'd6579, 16'd28568});
	test_expansion(128'h5c6951cf97d6d92138dd07bf5c7a557e, {16'd50008, 16'd47812, 16'd35808, 16'd49048, 16'd3496, 16'd49812, 16'd2695, 16'd37529, 16'd56282, 16'd30162, 16'd3386, 16'd4755, 16'd12996, 16'd28357, 16'd59117, 16'd43821, 16'd2371, 16'd33512, 16'd61037, 16'd31929, 16'd18092, 16'd39726, 16'd65471, 16'd10885, 16'd17691, 16'd52220});
	test_expansion(128'hde3818b568d15dbd338c6c82b9f75ae7, {16'd54473, 16'd52441, 16'd45070, 16'd7405, 16'd58899, 16'd55966, 16'd22810, 16'd5066, 16'd29205, 16'd36046, 16'd24914, 16'd27132, 16'd6841, 16'd1062, 16'd7949, 16'd25634, 16'd60644, 16'd34807, 16'd30205, 16'd13462, 16'd1371, 16'd9306, 16'd15377, 16'd31051, 16'd65311, 16'd60836});
	test_expansion(128'h7335f6fddedb7db6932744563c4b7cc2, {16'd36325, 16'd30881, 16'd59658, 16'd43255, 16'd7904, 16'd21438, 16'd10061, 16'd21734, 16'd3210, 16'd9335, 16'd24605, 16'd8539, 16'd22539, 16'd5930, 16'd50087, 16'd38021, 16'd47964, 16'd64072, 16'd53808, 16'd48971, 16'd3212, 16'd1157, 16'd43263, 16'd6478, 16'd3368, 16'd20534});
	test_expansion(128'h1ac3c48fbb4de0c093cc796ff832077f, {16'd44387, 16'd952, 16'd39316, 16'd27716, 16'd5562, 16'd38179, 16'd31576, 16'd47045, 16'd13250, 16'd37239, 16'd40076, 16'd24079, 16'd47142, 16'd43794, 16'd60206, 16'd54701, 16'd64209, 16'd34742, 16'd815, 16'd61120, 16'd8364, 16'd12707, 16'd8798, 16'd4674, 16'd14848, 16'd53503});
	test_expansion(128'h1c03b31a90a6071c3a9e9758ab33fc7a, {16'd29892, 16'd3460, 16'd25666, 16'd59604, 16'd47559, 16'd28619, 16'd21958, 16'd16587, 16'd56295, 16'd49935, 16'd37674, 16'd24391, 16'd29521, 16'd4785, 16'd14482, 16'd4587, 16'd53497, 16'd39432, 16'd46474, 16'd8656, 16'd25938, 16'd39233, 16'd11127, 16'd27822, 16'd49799, 16'd37596});
	test_expansion(128'hbed3a051ec043028e4b0a752f3e8049c, {16'd36572, 16'd32518, 16'd47012, 16'd57538, 16'd18232, 16'd36149, 16'd47698, 16'd7985, 16'd22913, 16'd54477, 16'd156, 16'd46792, 16'd61410, 16'd2869, 16'd28468, 16'd2443, 16'd27111, 16'd26641, 16'd27548, 16'd42735, 16'd30938, 16'd20415, 16'd51416, 16'd30149, 16'd3949, 16'd36888});
	test_expansion(128'hb5e796a25c6dd73b096e8ff9aed0b1f1, {16'd36729, 16'd44455, 16'd56120, 16'd44217, 16'd58506, 16'd59525, 16'd25747, 16'd64781, 16'd14240, 16'd52700, 16'd35818, 16'd12968, 16'd1987, 16'd44982, 16'd41155, 16'd6108, 16'd3177, 16'd11680, 16'd29938, 16'd23729, 16'd17543, 16'd5982, 16'd6958, 16'd54781, 16'd41998, 16'd14297});
	test_expansion(128'h14f2f6f8bb5f433ae59d97bcb02c2ffd, {16'd55471, 16'd21759, 16'd3843, 16'd55744, 16'd569, 16'd18344, 16'd28869, 16'd6353, 16'd48700, 16'd8149, 16'd28084, 16'd13054, 16'd9804, 16'd25406, 16'd38711, 16'd43590, 16'd49225, 16'd1717, 16'd61470, 16'd64514, 16'd27186, 16'd12485, 16'd58336, 16'd63873, 16'd5040, 16'd43321});
	test_expansion(128'h28e50ecfc882771b70460a2c934023a0, {16'd2997, 16'd42779, 16'd42719, 16'd35239, 16'd41482, 16'd39218, 16'd6912, 16'd12488, 16'd24407, 16'd17749, 16'd18575, 16'd44063, 16'd50854, 16'd28357, 16'd18803, 16'd38305, 16'd22000, 16'd20461, 16'd20642, 16'd50046, 16'd31218, 16'd16728, 16'd45255, 16'd14910, 16'd39611, 16'd19336});
	test_expansion(128'hd13eac3c27f5d38714e8f29a5835d8e3, {16'd6651, 16'd54086, 16'd50680, 16'd47558, 16'd24774, 16'd60821, 16'd52950, 16'd13792, 16'd47991, 16'd64714, 16'd5364, 16'd31128, 16'd30118, 16'd55462, 16'd55043, 16'd39232, 16'd37186, 16'd52379, 16'd53322, 16'd5755, 16'd51335, 16'd25168, 16'd57804, 16'd59666, 16'd8461, 16'd43582});
	test_expansion(128'ha048d1e584608cbcb6a71c4bf3372771, {16'd55146, 16'd7349, 16'd65146, 16'd2821, 16'd51203, 16'd4215, 16'd1552, 16'd12240, 16'd60526, 16'd25060, 16'd5014, 16'd56610, 16'd24962, 16'd6923, 16'd56980, 16'd19421, 16'd25560, 16'd55181, 16'd64772, 16'd33335, 16'd10704, 16'd8267, 16'd34693, 16'd53736, 16'd42676, 16'd35715});
	test_expansion(128'h84893612a38948aacf006969ecb1fbf4, {16'd35062, 16'd52419, 16'd20721, 16'd30823, 16'd10862, 16'd48799, 16'd55276, 16'd32749, 16'd36575, 16'd50295, 16'd57027, 16'd255, 16'd43379, 16'd26478, 16'd46083, 16'd51931, 16'd23641, 16'd55082, 16'd40252, 16'd16375, 16'd3191, 16'd11115, 16'd22994, 16'd8202, 16'd56289, 16'd52022});
	test_expansion(128'h9f7cdd7fb96c17e5d1c7a904251d99ea, {16'd16102, 16'd854, 16'd48374, 16'd14184, 16'd477, 16'd13678, 16'd53270, 16'd51219, 16'd39835, 16'd53968, 16'd40027, 16'd2601, 16'd64839, 16'd30965, 16'd19080, 16'd725, 16'd38209, 16'd23529, 16'd27718, 16'd51802, 16'd54714, 16'd12153, 16'd18009, 16'd58907, 16'd17690, 16'd42926});
	test_expansion(128'h163220465b35d1c3a64ec8ed3e56de2c, {16'd10379, 16'd9050, 16'd10906, 16'd37040, 16'd38518, 16'd56226, 16'd20127, 16'd7225, 16'd44414, 16'd59417, 16'd19956, 16'd25242, 16'd51122, 16'd57345, 16'd53355, 16'd51784, 16'd52983, 16'd26257, 16'd26844, 16'd60734, 16'd57409, 16'd33475, 16'd24947, 16'd38116, 16'd35967, 16'd64598});
	test_expansion(128'h660b44ee42722a10733a29dc2db0227b, {16'd28619, 16'd7122, 16'd2492, 16'd58713, 16'd1399, 16'd65512, 16'd31977, 16'd60162, 16'd33833, 16'd34948, 16'd9301, 16'd27339, 16'd12808, 16'd38914, 16'd16894, 16'd57380, 16'd29900, 16'd58879, 16'd2978, 16'd33735, 16'd24256, 16'd22019, 16'd6215, 16'd11211, 16'd24091, 16'd48810});
	test_expansion(128'h813c6f51bdc0152e02089f44b33cf104, {16'd49501, 16'd41823, 16'd25654, 16'd44571, 16'd8833, 16'd32985, 16'd4426, 16'd540, 16'd14044, 16'd32604, 16'd41142, 16'd51047, 16'd17724, 16'd56198, 16'd40974, 16'd51574, 16'd48896, 16'd47908, 16'd39089, 16'd18232, 16'd32544, 16'd53646, 16'd19764, 16'd25219, 16'd23111, 16'd45288});
	test_expansion(128'hf6fd8dcbccd2b4927c412befaf8f155b, {16'd64799, 16'd19404, 16'd65074, 16'd50416, 16'd56144, 16'd39906, 16'd6622, 16'd33029, 16'd32923, 16'd5687, 16'd30186, 16'd27363, 16'd4874, 16'd46718, 16'd44955, 16'd63511, 16'd47062, 16'd43507, 16'd40460, 16'd27119, 16'd64719, 16'd64557, 16'd39488, 16'd54419, 16'd45646, 16'd7087});
	test_expansion(128'hdc2d80d1410c3bd4ab2427fe34ecc477, {16'd11325, 16'd45006, 16'd48290, 16'd48416, 16'd46928, 16'd23980, 16'd18434, 16'd24233, 16'd26327, 16'd11950, 16'd15026, 16'd54492, 16'd7457, 16'd8166, 16'd55469, 16'd19097, 16'd8643, 16'd10190, 16'd57640, 16'd21302, 16'd1608, 16'd63164, 16'd61735, 16'd62650, 16'd21516, 16'd5801});
	test_expansion(128'hdc1289929fea52b7988822310e533400, {16'd21853, 16'd3802, 16'd10686, 16'd62144, 16'd23130, 16'd20744, 16'd14350, 16'd14709, 16'd22243, 16'd51792, 16'd45055, 16'd18705, 16'd53807, 16'd33186, 16'd59149, 16'd10077, 16'd19979, 16'd34234, 16'd20576, 16'd63106, 16'd19965, 16'd14400, 16'd58105, 16'd11020, 16'd42899, 16'd35579});
	test_expansion(128'h8d3d01ce932fc9d29ebf83d9f5db7405, {16'd15212, 16'd29357, 16'd4228, 16'd59236, 16'd59981, 16'd644, 16'd5447, 16'd40325, 16'd64243, 16'd13802, 16'd30008, 16'd45032, 16'd58442, 16'd53527, 16'd33475, 16'd34941, 16'd42011, 16'd54976, 16'd40337, 16'd13064, 16'd31132, 16'd26016, 16'd46000, 16'd32989, 16'd33325, 16'd6473});
	test_expansion(128'h47b7e1be32395671fe772cb6d083bf29, {16'd58375, 16'd54948, 16'd57157, 16'd28078, 16'd30465, 16'd2202, 16'd57879, 16'd9414, 16'd56006, 16'd31194, 16'd47518, 16'd18832, 16'd21345, 16'd3680, 16'd56308, 16'd49649, 16'd27995, 16'd59416, 16'd4509, 16'd7178, 16'd30341, 16'd64096, 16'd54229, 16'd12807, 16'd43054, 16'd10331});
	test_expansion(128'h03300f454f2be5aec59c745c3a43169e, {16'd42111, 16'd52626, 16'd2015, 16'd45598, 16'd27414, 16'd50949, 16'd63574, 16'd47643, 16'd40400, 16'd32680, 16'd31650, 16'd812, 16'd17843, 16'd45377, 16'd35464, 16'd25491, 16'd49851, 16'd53687, 16'd10876, 16'd35490, 16'd50347, 16'd2785, 16'd37407, 16'd62753, 16'd63763, 16'd48900});
	test_expansion(128'hbae5ca2969470051fbd165b3100b7c40, {16'd15723, 16'd6093, 16'd51073, 16'd48975, 16'd919, 16'd59975, 16'd20392, 16'd61236, 16'd20888, 16'd34286, 16'd15662, 16'd31101, 16'd56128, 16'd64356, 16'd41976, 16'd13392, 16'd28270, 16'd559, 16'd42878, 16'd13979, 16'd59520, 16'd28090, 16'd48366, 16'd9398, 16'd53517, 16'd7087});
	test_expansion(128'h3466fa3d533bf1533bb000fcdc4a51f4, {16'd35231, 16'd52503, 16'd49618, 16'd35073, 16'd57062, 16'd32523, 16'd27557, 16'd16262, 16'd4783, 16'd40746, 16'd16744, 16'd40943, 16'd48156, 16'd13543, 16'd37957, 16'd55806, 16'd57780, 16'd14199, 16'd19341, 16'd48242, 16'd19875, 16'd64322, 16'd37492, 16'd5351, 16'd60513, 16'd19467});
	test_expansion(128'h37bb21fa06081f430cbcbcdd62adf637, {16'd13141, 16'd62532, 16'd39603, 16'd54704, 16'd43957, 16'd7270, 16'd19053, 16'd63015, 16'd39978, 16'd16693, 16'd2676, 16'd17781, 16'd4718, 16'd6609, 16'd52939, 16'd60471, 16'd15647, 16'd7633, 16'd32981, 16'd44593, 16'd2191, 16'd2035, 16'd1959, 16'd16747, 16'd26106, 16'd41955});
	test_expansion(128'h0b08891ae4188bba177d94b780421be8, {16'd13961, 16'd29212, 16'd38518, 16'd17090, 16'd9177, 16'd38356, 16'd48363, 16'd9729, 16'd11925, 16'd18634, 16'd56706, 16'd24484, 16'd16288, 16'd4240, 16'd61685, 16'd6234, 16'd25520, 16'd51741, 16'd64063, 16'd34036, 16'd21496, 16'd28335, 16'd28268, 16'd64587, 16'd2537, 16'd5255});
	test_expansion(128'h6945e5284fadc4d11cae50c83df2f9d2, {16'd38455, 16'd35854, 16'd14691, 16'd30531, 16'd21697, 16'd48205, 16'd62336, 16'd55646, 16'd21395, 16'd35231, 16'd30523, 16'd33690, 16'd14839, 16'd26466, 16'd55307, 16'd3624, 16'd23666, 16'd57025, 16'd2522, 16'd3699, 16'd30063, 16'd63767, 16'd32905, 16'd12582, 16'd11830, 16'd31361});
	test_expansion(128'h340450d4e8eda79dd265774cf43d2042, {16'd7345, 16'd23042, 16'd61416, 16'd45374, 16'd20201, 16'd21198, 16'd11828, 16'd47941, 16'd62840, 16'd29145, 16'd60766, 16'd52209, 16'd33517, 16'd3790, 16'd20760, 16'd62908, 16'd47930, 16'd18508, 16'd2497, 16'd38342, 16'd21617, 16'd55724, 16'd28911, 16'd6114, 16'd43340, 16'd17797});
	test_expansion(128'h4ca21ef36c46aefebe1bef94d7d7e015, {16'd24894, 16'd2756, 16'd57163, 16'd58485, 16'd15132, 16'd6306, 16'd40349, 16'd5610, 16'd45345, 16'd14236, 16'd29104, 16'd49350, 16'd5601, 16'd63635, 16'd32802, 16'd18062, 16'd58702, 16'd18101, 16'd25728, 16'd30011, 16'd52001, 16'd61534, 16'd47206, 16'd37363, 16'd19225, 16'd30617});
	test_expansion(128'h9675a6878de0ffe0b65aa0bb6a2ab4e6, {16'd31502, 16'd29000, 16'd24485, 16'd48847, 16'd49404, 16'd20788, 16'd43067, 16'd37187, 16'd6240, 16'd56164, 16'd53029, 16'd28500, 16'd1737, 16'd7483, 16'd17984, 16'd37745, 16'd54095, 16'd2946, 16'd12369, 16'd28250, 16'd17748, 16'd54767, 16'd61318, 16'd54125, 16'd12959, 16'd17304});
	test_expansion(128'h8a5447f1d8eea428f531307cf4f55d5c, {16'd50736, 16'd5035, 16'd54182, 16'd43654, 16'd19940, 16'd16189, 16'd15833, 16'd35191, 16'd645, 16'd10962, 16'd37892, 16'd63382, 16'd41435, 16'd28325, 16'd60366, 16'd9409, 16'd42950, 16'd23617, 16'd62306, 16'd55805, 16'd51971, 16'd59360, 16'd38481, 16'd25017, 16'd42312, 16'd35622});
	test_expansion(128'h261478ae2a06f6fffe9f74107ef6d856, {16'd55057, 16'd58960, 16'd29253, 16'd14643, 16'd36632, 16'd20231, 16'd4410, 16'd4544, 16'd25001, 16'd4466, 16'd51651, 16'd42254, 16'd47622, 16'd53176, 16'd11533, 16'd29159, 16'd62946, 16'd33188, 16'd52226, 16'd240, 16'd14292, 16'd2412, 16'd26769, 16'd57533, 16'd4109, 16'd5812});
	test_expansion(128'h75cbcbf547761ac8a90c9b39aa56bd05, {16'd58982, 16'd35334, 16'd19993, 16'd4928, 16'd33221, 16'd53473, 16'd23923, 16'd37265, 16'd17143, 16'd65008, 16'd34341, 16'd36363, 16'd52755, 16'd53463, 16'd25678, 16'd3950, 16'd37508, 16'd28694, 16'd52887, 16'd59702, 16'd63609, 16'd467, 16'd17357, 16'd7133, 16'd24645, 16'd43517});
	test_expansion(128'hff7f9bb83bdc188054403838c17650f9, {16'd35487, 16'd5136, 16'd38730, 16'd61573, 16'd36376, 16'd32973, 16'd61817, 16'd881, 16'd63151, 16'd41973, 16'd8581, 16'd11945, 16'd18255, 16'd26397, 16'd43132, 16'd29494, 16'd21263, 16'd65341, 16'd62639, 16'd17017, 16'd44827, 16'd50896, 16'd35849, 16'd64035, 16'd22255, 16'd12155});
	test_expansion(128'h9ec7524b391b819f5dac618371afc5d7, {16'd3943, 16'd5268, 16'd18054, 16'd54822, 16'd36683, 16'd57101, 16'd60626, 16'd28725, 16'd12021, 16'd64233, 16'd33291, 16'd26880, 16'd60807, 16'd36704, 16'd27874, 16'd50189, 16'd22341, 16'd58377, 16'd55008, 16'd60412, 16'd27015, 16'd35342, 16'd28796, 16'd17079, 16'd41389, 16'd27635});
	test_expansion(128'ha6533d461b9c265ddab485bafdeaf314, {16'd59097, 16'd54060, 16'd45534, 16'd7039, 16'd26671, 16'd10320, 16'd26556, 16'd58072, 16'd35818, 16'd55337, 16'd32626, 16'd52977, 16'd17287, 16'd59530, 16'd10993, 16'd25620, 16'd45897, 16'd21968, 16'd45467, 16'd40508, 16'd34493, 16'd48206, 16'd28025, 16'd1118, 16'd20104, 16'd50396});
	test_expansion(128'h495215934897bfba9f7ff8329b9aa8ce, {16'd32727, 16'd65232, 16'd56151, 16'd14669, 16'd1607, 16'd37964, 16'd48, 16'd33336, 16'd32992, 16'd9013, 16'd58900, 16'd31917, 16'd23519, 16'd61121, 16'd29559, 16'd30905, 16'd27163, 16'd39164, 16'd47210, 16'd33574, 16'd48646, 16'd54219, 16'd47822, 16'd27604, 16'd65484, 16'd38759});
	test_expansion(128'hae3b72c8e304222040050e224d70ebe1, {16'd45751, 16'd24703, 16'd52379, 16'd56125, 16'd6092, 16'd31780, 16'd29093, 16'd55152, 16'd16968, 16'd28904, 16'd47249, 16'd15351, 16'd64040, 16'd63546, 16'd19452, 16'd58266, 16'd21606, 16'd62836, 16'd33513, 16'd54836, 16'd23397, 16'd45366, 16'd15864, 16'd39798, 16'd19497, 16'd1076});
	test_expansion(128'h9193f02be35b86cb0f9183591ce8c065, {16'd21696, 16'd14487, 16'd333, 16'd29270, 16'd395, 16'd6394, 16'd38909, 16'd2005, 16'd13272, 16'd17515, 16'd59343, 16'd18255, 16'd39156, 16'd37802, 16'd5757, 16'd18665, 16'd61753, 16'd7594, 16'd45622, 16'd11873, 16'd60843, 16'd35288, 16'd17694, 16'd744, 16'd36333, 16'd2476});
	test_expansion(128'h1443d68513a2ddb5a23b15a563a03c57, {16'd13329, 16'd18960, 16'd61542, 16'd16899, 16'd52826, 16'd10538, 16'd64350, 16'd32615, 16'd4945, 16'd63262, 16'd9796, 16'd28725, 16'd3917, 16'd4089, 16'd24238, 16'd15616, 16'd51792, 16'd60118, 16'd38083, 16'd57340, 16'd4459, 16'd52841, 16'd88, 16'd55999, 16'd20178, 16'd20064});
	test_expansion(128'h8f0859bd5d5700a1b7064d6e213110b5, {16'd39285, 16'd12486, 16'd52749, 16'd28760, 16'd38464, 16'd8378, 16'd41089, 16'd44061, 16'd20645, 16'd6359, 16'd38940, 16'd21617, 16'd63383, 16'd48998, 16'd2256, 16'd841, 16'd20878, 16'd1074, 16'd11948, 16'd28815, 16'd10224, 16'd6333, 16'd31809, 16'd5507, 16'd47248, 16'd40085});
	test_expansion(128'h656640ba551e13fb4ec5c8200602a7c0, {16'd4624, 16'd48756, 16'd46398, 16'd7294, 16'd49806, 16'd47022, 16'd46520, 16'd23494, 16'd2497, 16'd31497, 16'd56024, 16'd57735, 16'd16109, 16'd48102, 16'd10846, 16'd20182, 16'd10207, 16'd17140, 16'd10509, 16'd26817, 16'd42177, 16'd50427, 16'd9749, 16'd40592, 16'd12938, 16'd39315});
	test_expansion(128'h75d0826aaea05e45c30a51a182458194, {16'd14382, 16'd31004, 16'd14531, 16'd61080, 16'd29357, 16'd39925, 16'd31719, 16'd5792, 16'd34260, 16'd11273, 16'd1807, 16'd54998, 16'd39789, 16'd9753, 16'd7482, 16'd26598, 16'd36124, 16'd7756, 16'd55754, 16'd23019, 16'd24998, 16'd59856, 16'd39735, 16'd41929, 16'd27346, 16'd37807});
	test_expansion(128'h3211a58d9b4b9faf455b2b38e05ef577, {16'd54646, 16'd18373, 16'd637, 16'd62135, 16'd64740, 16'd20679, 16'd49885, 16'd41522, 16'd44718, 16'd12916, 16'd27377, 16'd787, 16'd21497, 16'd12277, 16'd25066, 16'd24517, 16'd44069, 16'd8536, 16'd7825, 16'd60490, 16'd5757, 16'd39276, 16'd42457, 16'd34195, 16'd64724, 16'd9963});
	test_expansion(128'haaec50e9b71e56a9efdf3923798e2a49, {16'd42747, 16'd23514, 16'd39906, 16'd4194, 16'd18008, 16'd62126, 16'd59288, 16'd33597, 16'd46978, 16'd16775, 16'd43185, 16'd31977, 16'd9772, 16'd60717, 16'd60530, 16'd37170, 16'd6860, 16'd17384, 16'd63358, 16'd51827, 16'd33491, 16'd38813, 16'd56613, 16'd17353, 16'd25931, 16'd62803});
	test_expansion(128'h24a9097718238a0d511ace63f3823d40, {16'd37627, 16'd63834, 16'd43148, 16'd31366, 16'd11287, 16'd48367, 16'd8747, 16'd35607, 16'd36673, 16'd38709, 16'd21181, 16'd6206, 16'd15283, 16'd24643, 16'd35549, 16'd57770, 16'd12637, 16'd61430, 16'd50339, 16'd11678, 16'd26496, 16'd22168, 16'd12570, 16'd36307, 16'd23609, 16'd55698});
	test_expansion(128'h1c37d7ecd760c009468cc48e8d1c6978, {16'd38807, 16'd52033, 16'd47007, 16'd57061, 16'd44957, 16'd631, 16'd34456, 16'd53991, 16'd24597, 16'd40916, 16'd26401, 16'd47441, 16'd14965, 16'd20536, 16'd22002, 16'd51895, 16'd49276, 16'd301, 16'd14432, 16'd48515, 16'd1891, 16'd209, 16'd3168, 16'd42729, 16'd29285, 16'd9130});
	test_expansion(128'h820524c70aa13b44c3e17958fc8b005a, {16'd46521, 16'd56720, 16'd44284, 16'd7915, 16'd60563, 16'd35120, 16'd40923, 16'd40069, 16'd44617, 16'd5761, 16'd17408, 16'd55963, 16'd58460, 16'd21793, 16'd49906, 16'd19178, 16'd17232, 16'd59713, 16'd42881, 16'd59892, 16'd64371, 16'd3350, 16'd59048, 16'd47975, 16'd40982, 16'd22311});
	test_expansion(128'h02a1f82da0b8acc7df50f9747f471832, {16'd40968, 16'd56161, 16'd38418, 16'd64090, 16'd24500, 16'd30288, 16'd16125, 16'd27532, 16'd15067, 16'd24414, 16'd42111, 16'd64306, 16'd29507, 16'd16647, 16'd49214, 16'd49612, 16'd47509, 16'd41012, 16'd55445, 16'd3446, 16'd59084, 16'd18207, 16'd29902, 16'd8676, 16'd23963, 16'd49733});
	test_expansion(128'h7f5e7a1790b006628cafe64498594ba5, {16'd38218, 16'd12528, 16'd38198, 16'd36819, 16'd32109, 16'd32106, 16'd2292, 16'd20037, 16'd46687, 16'd46046, 16'd38064, 16'd10993, 16'd38820, 16'd43397, 16'd40068, 16'd41662, 16'd26837, 16'd36882, 16'd13, 16'd30865, 16'd12538, 16'd7400, 16'd18685, 16'd23865, 16'd58850, 16'd54151});
	test_expansion(128'h7803828751067d0e4e6b110f2a51ff4d, {16'd42964, 16'd2875, 16'd38772, 16'd47505, 16'd60869, 16'd27497, 16'd10700, 16'd7539, 16'd23811, 16'd34315, 16'd60957, 16'd55129, 16'd1395, 16'd23242, 16'd40976, 16'd40387, 16'd20426, 16'd57086, 16'd32232, 16'd12637, 16'd572, 16'd9919, 16'd23782, 16'd54566, 16'd46981, 16'd56863});
	test_expansion(128'h98b058d65dba6d9f84bfb9a8a48fd7a8, {16'd52583, 16'd43903, 16'd36117, 16'd9550, 16'd65403, 16'd13934, 16'd52715, 16'd38133, 16'd56919, 16'd28918, 16'd7275, 16'd63922, 16'd17029, 16'd33038, 16'd42527, 16'd52811, 16'd11810, 16'd55550, 16'd62406, 16'd24185, 16'd60129, 16'd9274, 16'd12850, 16'd7223, 16'd62774, 16'd12676});
	test_expansion(128'hdda3c662d65fc086a8f5aea3985b3d7a, {16'd53987, 16'd18553, 16'd59508, 16'd16176, 16'd30019, 16'd40811, 16'd61182, 16'd26350, 16'd23341, 16'd36260, 16'd63903, 16'd63912, 16'd27741, 16'd28078, 16'd9848, 16'd14681, 16'd21161, 16'd16921, 16'd9955, 16'd43522, 16'd58806, 16'd11792, 16'd37429, 16'd63400, 16'd42080, 16'd12239});
	test_expansion(128'h66f3948073cf1de3ea612903cb21f9c3, {16'd17706, 16'd6973, 16'd14822, 16'd1203, 16'd51901, 16'd10795, 16'd21892, 16'd43591, 16'd58341, 16'd40767, 16'd30790, 16'd44719, 16'd13050, 16'd24221, 16'd19867, 16'd36230, 16'd41598, 16'd31925, 16'd62469, 16'd56178, 16'd62209, 16'd13102, 16'd21181, 16'd56060, 16'd44683, 16'd38303});
	test_expansion(128'he34c2040ed287181a717a1a3ae286318, {16'd29048, 16'd21879, 16'd43110, 16'd54632, 16'd37458, 16'd38619, 16'd59397, 16'd34627, 16'd49026, 16'd33728, 16'd15871, 16'd31386, 16'd21262, 16'd14366, 16'd21986, 16'd62919, 16'd9902, 16'd25062, 16'd7233, 16'd50208, 16'd2429, 16'd6703, 16'd36927, 16'd8405, 16'd45267, 16'd61707});
	test_expansion(128'h7c92f225910450f2e29626a694a9b558, {16'd47876, 16'd45284, 16'd13592, 16'd57623, 16'd44767, 16'd24323, 16'd48348, 16'd36691, 16'd11924, 16'd6068, 16'd10962, 16'd57508, 16'd15363, 16'd14190, 16'd56679, 16'd60894, 16'd52497, 16'd44765, 16'd36586, 16'd47443, 16'd40999, 16'd8118, 16'd19523, 16'd53652, 16'd27564, 16'd47926});
	test_expansion(128'h85ce9ab852ed1a2d1984b739d536f634, {16'd23341, 16'd11122, 16'd42850, 16'd59954, 16'd18435, 16'd15078, 16'd30919, 16'd52964, 16'd15541, 16'd34999, 16'd38202, 16'd35911, 16'd26012, 16'd12947, 16'd18158, 16'd46061, 16'd30184, 16'd50078, 16'd55875, 16'd33978, 16'd54840, 16'd46801, 16'd12003, 16'd39376, 16'd2883, 16'd54252});
	test_expansion(128'h24b8875b062db8c17ecb5a832539450d, {16'd46472, 16'd4581, 16'd30811, 16'd56016, 16'd64887, 16'd1628, 16'd61107, 16'd21065, 16'd49877, 16'd47437, 16'd4936, 16'd49788, 16'd50829, 16'd59451, 16'd38257, 16'd8609, 16'd46941, 16'd59105, 16'd14660, 16'd31177, 16'd60749, 16'd28406, 16'd24873, 16'd5980, 16'd41369, 16'd64738});
	test_expansion(128'h9b5fe26e40a392c446ff955ecfbdd45f, {16'd1677, 16'd53501, 16'd22297, 16'd19563, 16'd27144, 16'd55078, 16'd13993, 16'd13834, 16'd23552, 16'd27921, 16'd20331, 16'd43984, 16'd42107, 16'd30149, 16'd34459, 16'd12590, 16'd38380, 16'd37041, 16'd14545, 16'd20777, 16'd43803, 16'd34913, 16'd55556, 16'd60164, 16'd36749, 16'd5799});
	test_expansion(128'h4d471159c4f9ef3a28aeae88c08e6851, {16'd25247, 16'd65089, 16'd53563, 16'd35617, 16'd56783, 16'd49592, 16'd46649, 16'd21077, 16'd56026, 16'd62699, 16'd13424, 16'd15207, 16'd10448, 16'd43444, 16'd4701, 16'd62116, 16'd12880, 16'd44821, 16'd58862, 16'd26840, 16'd54622, 16'd937, 16'd53994, 16'd13602, 16'd65013, 16'd7270});
	test_expansion(128'h0307edb3ab22a4f4a546d4b53a81e220, {16'd12239, 16'd56113, 16'd43250, 16'd23661, 16'd47666, 16'd65324, 16'd51805, 16'd62132, 16'd12884, 16'd24959, 16'd4536, 16'd10887, 16'd53532, 16'd34913, 16'd12963, 16'd34461, 16'd60414, 16'd16272, 16'd21019, 16'd6448, 16'd30659, 16'd33605, 16'd16020, 16'd21550, 16'd56487, 16'd12188});
	test_expansion(128'he770932cef59fee2951386c3da247812, {16'd25197, 16'd57811, 16'd524, 16'd41627, 16'd14528, 16'd24565, 16'd7722, 16'd58457, 16'd45788, 16'd21487, 16'd12011, 16'd32882, 16'd51020, 16'd65477, 16'd27274, 16'd3272, 16'd2835, 16'd30298, 16'd35593, 16'd42574, 16'd23827, 16'd36968, 16'd46910, 16'd5685, 16'd30087, 16'd12583});
	test_expansion(128'hd0c840ecd21fb8053933e12d304bfb92, {16'd25036, 16'd62931, 16'd35028, 16'd32039, 16'd6987, 16'd53187, 16'd27769, 16'd61041, 16'd10477, 16'd3066, 16'd4812, 16'd26717, 16'd21924, 16'd47837, 16'd53108, 16'd58532, 16'd29647, 16'd64343, 16'd31075, 16'd1768, 16'd60805, 16'd22200, 16'd18303, 16'd65242, 16'd35551, 16'd45489});
	test_expansion(128'h29b692097afa157d4037ae0f1e87e80a, {16'd48317, 16'd13523, 16'd41269, 16'd38764, 16'd57671, 16'd30313, 16'd54019, 16'd1735, 16'd56543, 16'd39240, 16'd55623, 16'd34128, 16'd63362, 16'd2121, 16'd62495, 16'd35013, 16'd47227, 16'd38749, 16'd64026, 16'd28418, 16'd46825, 16'd21375, 16'd27682, 16'd5771, 16'd5047, 16'd17724});
	test_expansion(128'ha75711dd23d7d5b039b4fa611e728fd3, {16'd27354, 16'd25673, 16'd49087, 16'd56446, 16'd58010, 16'd3868, 16'd48749, 16'd40081, 16'd47058, 16'd55484, 16'd15210, 16'd59906, 16'd49765, 16'd36826, 16'd23391, 16'd64910, 16'd34766, 16'd53290, 16'd45278, 16'd35294, 16'd16429, 16'd53726, 16'd45169, 16'd42641, 16'd50330, 16'd45554});
	test_expansion(128'h5073208d0dd410a371b85dd15f5ae9d7, {16'd23811, 16'd56334, 16'd17025, 16'd16922, 16'd33968, 16'd3892, 16'd57260, 16'd28964, 16'd19714, 16'd30290, 16'd35937, 16'd26947, 16'd12489, 16'd13924, 16'd36471, 16'd10892, 16'd50832, 16'd10588, 16'd54400, 16'd41872, 16'd45378, 16'd6142, 16'd10181, 16'd38726, 16'd27788, 16'd19807});
	test_expansion(128'h4e73d999d4f4772dc5e554e10f8a3eae, {16'd26696, 16'd25714, 16'd50325, 16'd5957, 16'd47236, 16'd2804, 16'd17568, 16'd44634, 16'd18701, 16'd12591, 16'd29945, 16'd33733, 16'd15707, 16'd27585, 16'd25892, 16'd6743, 16'd46728, 16'd38269, 16'd54679, 16'd13015, 16'd10625, 16'd17600, 16'd59266, 16'd762, 16'd8595, 16'd35756});
	test_expansion(128'hbc7f09b965ad1035ebd380d8e7b76c00, {16'd51597, 16'd29520, 16'd58620, 16'd27116, 16'd21432, 16'd37192, 16'd38043, 16'd33918, 16'd64018, 16'd36666, 16'd63138, 16'd62378, 16'd41293, 16'd52542, 16'd3751, 16'd37202, 16'd64095, 16'd64761, 16'd45534, 16'd57419, 16'd48501, 16'd826, 16'd56841, 16'd5926, 16'd25586, 16'd26286});
	test_expansion(128'h73a6a084fd3f6b48b8fb793aeb791e07, {16'd7964, 16'd32002, 16'd62564, 16'd17086, 16'd11429, 16'd28962, 16'd220, 16'd6621, 16'd48083, 16'd20279, 16'd15919, 16'd55272, 16'd12812, 16'd9602, 16'd49256, 16'd21895, 16'd22212, 16'd63116, 16'd44251, 16'd54259, 16'd25364, 16'd24060, 16'd4997, 16'd42678, 16'd37990, 16'd19401});
	test_expansion(128'h85e7d325686da8a2980f7df1cda70505, {16'd18015, 16'd39293, 16'd31673, 16'd15940, 16'd15649, 16'd27219, 16'd33403, 16'd42104, 16'd58510, 16'd39905, 16'd28784, 16'd26987, 16'd43461, 16'd40604, 16'd1619, 16'd59211, 16'd49023, 16'd30852, 16'd63449, 16'd21819, 16'd24807, 16'd2291, 16'd20227, 16'd39209, 16'd47081, 16'd30955});
	test_expansion(128'h7d9850ac343e768813ff298641924e1c, {16'd9818, 16'd21015, 16'd49544, 16'd1533, 16'd21446, 16'd59680, 16'd11588, 16'd51633, 16'd5131, 16'd57920, 16'd35179, 16'd64772, 16'd3069, 16'd18818, 16'd18459, 16'd34481, 16'd25910, 16'd32823, 16'd44894, 16'd3933, 16'd11150, 16'd4729, 16'd16254, 16'd51900, 16'd11804, 16'd29260});
	test_expansion(128'hbee91c14cb7ede8d9b2583ed18ab5b36, {16'd23446, 16'd11214, 16'd36640, 16'd23183, 16'd52931, 16'd12148, 16'd64650, 16'd40944, 16'd40028, 16'd61143, 16'd30635, 16'd41208, 16'd6980, 16'd64793, 16'd25883, 16'd10030, 16'd53907, 16'd2332, 16'd4024, 16'd24585, 16'd18362, 16'd20349, 16'd15403, 16'd27923, 16'd55961, 16'd63774});
	test_expansion(128'hf36aa88cece3b0d7599aac8fe3c37978, {16'd51440, 16'd33431, 16'd22629, 16'd56643, 16'd59366, 16'd56751, 16'd41143, 16'd59142, 16'd63671, 16'd26524, 16'd25589, 16'd14879, 16'd24529, 16'd18764, 16'd42300, 16'd16773, 16'd35751, 16'd45858, 16'd32848, 16'd37740, 16'd59074, 16'd31992, 16'd62650, 16'd45752, 16'd17001, 16'd64426});
	test_expansion(128'h362ec603c358a996448882278b037822, {16'd5388, 16'd43931, 16'd523, 16'd59676, 16'd43594, 16'd44971, 16'd26469, 16'd41791, 16'd12488, 16'd8035, 16'd23122, 16'd37300, 16'd47824, 16'd1605, 16'd29271, 16'd55942, 16'd20737, 16'd33097, 16'd1711, 16'd5930, 16'd46538, 16'd61021, 16'd1068, 16'd24285, 16'd38444, 16'd18537});
	test_expansion(128'hd6de7dbbb4d4cf79997ded8e64dc8955, {16'd51068, 16'd12071, 16'd25264, 16'd14470, 16'd59817, 16'd10085, 16'd5872, 16'd51537, 16'd47027, 16'd53730, 16'd7380, 16'd26296, 16'd4552, 16'd45490, 16'd41739, 16'd13326, 16'd29874, 16'd61720, 16'd29920, 16'd29090, 16'd16282, 16'd60913, 16'd54382, 16'd47297, 16'd10236, 16'd9751});
	test_expansion(128'h0aba7ef50735d9695d894790c34be2c0, {16'd19055, 16'd62882, 16'd60214, 16'd26388, 16'd8775, 16'd15249, 16'd60880, 16'd55983, 16'd30525, 16'd61771, 16'd20170, 16'd51124, 16'd8992, 16'd32232, 16'd10818, 16'd26469, 16'd23961, 16'd10303, 16'd17054, 16'd32053, 16'd28040, 16'd53807, 16'd47786, 16'd24265, 16'd12113, 16'd61409});
	test_expansion(128'h8753b40d340fcac14e7db1a5c456a877, {16'd3077, 16'd64637, 16'd62544, 16'd43627, 16'd13563, 16'd29770, 16'd35389, 16'd1023, 16'd6122, 16'd64319, 16'd54687, 16'd64554, 16'd35230, 16'd9138, 16'd3825, 16'd441, 16'd38713, 16'd5165, 16'd4226, 16'd12351, 16'd46213, 16'd45044, 16'd48884, 16'd34260, 16'd53236, 16'd25714});
	test_expansion(128'hce90f0a77a8bbfc204eb9db7910747bd, {16'd51728, 16'd2520, 16'd54805, 16'd37826, 16'd39305, 16'd23450, 16'd64848, 16'd46397, 16'd39950, 16'd11380, 16'd46894, 16'd28482, 16'd51436, 16'd25046, 16'd51052, 16'd57301, 16'd23319, 16'd54895, 16'd16869, 16'd22221, 16'd36341, 16'd41278, 16'd26964, 16'd48214, 16'd12612, 16'd50847});
	test_expansion(128'hecfa6690573543acf591d67a9c355015, {16'd41200, 16'd15979, 16'd12074, 16'd44735, 16'd11002, 16'd60899, 16'd4275, 16'd6436, 16'd38970, 16'd64766, 16'd51522, 16'd51538, 16'd2502, 16'd63291, 16'd52195, 16'd44807, 16'd43684, 16'd58014, 16'd3117, 16'd2241, 16'd33898, 16'd36186, 16'd24041, 16'd30433, 16'd65369, 16'd45783});
	test_expansion(128'hee0c363184ffa337467de78610b800e4, {16'd47142, 16'd48466, 16'd33648, 16'd45785, 16'd54732, 16'd18179, 16'd5039, 16'd23645, 16'd57568, 16'd61878, 16'd44164, 16'd4975, 16'd42009, 16'd35691, 16'd51499, 16'd19927, 16'd4295, 16'd50276, 16'd8959, 16'd57102, 16'd11068, 16'd59031, 16'd21552, 16'd55349, 16'd64714, 16'd60292});
	test_expansion(128'hc85429194a52ebda2fa10efd4522bf1f, {16'd25209, 16'd28130, 16'd21246, 16'd8462, 16'd49219, 16'd39795, 16'd24006, 16'd1371, 16'd38240, 16'd58875, 16'd41870, 16'd63131, 16'd3216, 16'd45316, 16'd3765, 16'd36175, 16'd57719, 16'd9909, 16'd60177, 16'd32220, 16'd24075, 16'd29832, 16'd39742, 16'd43069, 16'd44608, 16'd35066});
	test_expansion(128'h8ae52f6243f0bbe124fd452a9502f0cb, {16'd31005, 16'd35057, 16'd4058, 16'd1478, 16'd1884, 16'd32698, 16'd18734, 16'd13587, 16'd35294, 16'd46586, 16'd59785, 16'd23768, 16'd9657, 16'd27136, 16'd42701, 16'd9900, 16'd24429, 16'd8281, 16'd27066, 16'd50059, 16'd29164, 16'd4238, 16'd18291, 16'd45430, 16'd52224, 16'd611});
	test_expansion(128'hc26383b709bfff6194b5859583da1303, {16'd52455, 16'd20224, 16'd11477, 16'd51499, 16'd45014, 16'd33360, 16'd59865, 16'd30572, 16'd50303, 16'd26816, 16'd43397, 16'd14708, 16'd912, 16'd27251, 16'd25663, 16'd28072, 16'd58282, 16'd29410, 16'd43688, 16'd6982, 16'd64771, 16'd27843, 16'd33800, 16'd51369, 16'd35512, 16'd16160});
	test_expansion(128'h51cb81c95000636e371b2a91d48932b5, {16'd46851, 16'd15469, 16'd34592, 16'd33147, 16'd45069, 16'd249, 16'd50875, 16'd50845, 16'd29221, 16'd26461, 16'd33958, 16'd6574, 16'd8046, 16'd54013, 16'd59972, 16'd27723, 16'd16234, 16'd7295, 16'd41613, 16'd36820, 16'd26576, 16'd28850, 16'd48161, 16'd46490, 16'd60030, 16'd9279});
	test_expansion(128'h0f53cafdbb389b13e8423621b5a6d584, {16'd15400, 16'd30833, 16'd9846, 16'd17019, 16'd42435, 16'd60209, 16'd63596, 16'd1738, 16'd29305, 16'd30272, 16'd4724, 16'd21343, 16'd18415, 16'd607, 16'd2414, 16'd13492, 16'd43347, 16'd49679, 16'd51933, 16'd64522, 16'd6215, 16'd47196, 16'd19601, 16'd17983, 16'd28499, 16'd24771});
	test_expansion(128'hfb0e7a180735711eb736fd7e6a60a569, {16'd32870, 16'd41913, 16'd18421, 16'd39950, 16'd5145, 16'd31899, 16'd6506, 16'd19029, 16'd2490, 16'd29740, 16'd29370, 16'd24296, 16'd11551, 16'd43000, 16'd11841, 16'd10661, 16'd53913, 16'd16980, 16'd46973, 16'd51327, 16'd42417, 16'd51380, 16'd5274, 16'd59525, 16'd60504, 16'd34346});
	test_expansion(128'hfdb97c2771d01c00ab207caabfe6a1d0, {16'd27890, 16'd2610, 16'd43738, 16'd64419, 16'd37128, 16'd18157, 16'd21486, 16'd36172, 16'd45754, 16'd14451, 16'd35797, 16'd45731, 16'd44159, 16'd21150, 16'd30213, 16'd4602, 16'd22065, 16'd57955, 16'd44424, 16'd311, 16'd17856, 16'd12555, 16'd12046, 16'd28792, 16'd6473, 16'd14318});
	test_expansion(128'h9cb6199b5bc631da6063b1df36653085, {16'd35880, 16'd20377, 16'd31483, 16'd55536, 16'd35676, 16'd17455, 16'd6750, 16'd63566, 16'd62380, 16'd49445, 16'd52244, 16'd4382, 16'd16101, 16'd36785, 16'd26278, 16'd7376, 16'd21132, 16'd65088, 16'd48759, 16'd7161, 16'd24631, 16'd18575, 16'd26984, 16'd33729, 16'd3594, 16'd46306});
	test_expansion(128'hbc1b39df1a16fc46e415b41160b2f0cb, {16'd47143, 16'd42705, 16'd47873, 16'd24211, 16'd12110, 16'd24736, 16'd900, 16'd27927, 16'd54690, 16'd13347, 16'd62491, 16'd56810, 16'd14690, 16'd18689, 16'd35311, 16'd38875, 16'd27081, 16'd48582, 16'd55536, 16'd63286, 16'd50712, 16'd13153, 16'd37277, 16'd46160, 16'd17313, 16'd31980});
	test_expansion(128'ha9a83f1ecd55cba1f1e0df44eab16770, {16'd41097, 16'd37230, 16'd48892, 16'd64838, 16'd34051, 16'd65053, 16'd63591, 16'd32706, 16'd46872, 16'd42455, 16'd47618, 16'd12490, 16'd60097, 16'd40631, 16'd23267, 16'd22476, 16'd33181, 16'd61482, 16'd29524, 16'd63747, 16'd54849, 16'd49742, 16'd49558, 16'd38623, 16'd10690, 16'd62792});
	test_expansion(128'h5ddfa4444250f330661d2083c8313a8e, {16'd15787, 16'd37059, 16'd27942, 16'd53400, 16'd27742, 16'd9675, 16'd29088, 16'd48057, 16'd26488, 16'd60232, 16'd47579, 16'd11369, 16'd1605, 16'd2065, 16'd18119, 16'd46504, 16'd30509, 16'd46585, 16'd47675, 16'd57122, 16'd2965, 16'd56860, 16'd8182, 16'd53003, 16'd48573, 16'd4757});
	test_expansion(128'h77122eb35abaf75eae3bf062b5370241, {16'd16225, 16'd24649, 16'd23294, 16'd27706, 16'd41217, 16'd11112, 16'd61756, 16'd26713, 16'd28647, 16'd41344, 16'd24549, 16'd35601, 16'd12444, 16'd11414, 16'd35958, 16'd19796, 16'd23488, 16'd28113, 16'd7794, 16'd44507, 16'd32208, 16'd41064, 16'd38646, 16'd1332, 16'd7526, 16'd37125});
	test_expansion(128'he7fef8c55139ecd576d9aa530b917597, {16'd22816, 16'd63227, 16'd59682, 16'd17065, 16'd3259, 16'd61410, 16'd16628, 16'd24479, 16'd6549, 16'd51312, 16'd39596, 16'd20546, 16'd42858, 16'd15212, 16'd51486, 16'd34515, 16'd15748, 16'd6680, 16'd53694, 16'd10727, 16'd31624, 16'd28252, 16'd17097, 16'd3006, 16'd18692, 16'd60005});
	test_expansion(128'he4fa7f3413e395c81d6bbc6dd2012b1c, {16'd1765, 16'd50406, 16'd21393, 16'd36116, 16'd56806, 16'd55957, 16'd48844, 16'd13237, 16'd33825, 16'd15770, 16'd63577, 16'd43930, 16'd45325, 16'd13111, 16'd6420, 16'd35844, 16'd18055, 16'd12028, 16'd53541, 16'd21151, 16'd45168, 16'd60165, 16'd20046, 16'd63885, 16'd65025, 16'd2455});
	test_expansion(128'haf5640eed773e94a673b52843cd7af3c, {16'd57182, 16'd36451, 16'd47813, 16'd30917, 16'd55759, 16'd56048, 16'd35104, 16'd52914, 16'd65124, 16'd12685, 16'd45531, 16'd7810, 16'd20449, 16'd39659, 16'd13708, 16'd15854, 16'd42922, 16'd12667, 16'd25392, 16'd31009, 16'd3847, 16'd15535, 16'd65221, 16'd35366, 16'd33546, 16'd51348});
	test_expansion(128'hf4e58d14de07a9105be942d11ad27646, {16'd3720, 16'd36521, 16'd23917, 16'd30258, 16'd25876, 16'd22635, 16'd44100, 16'd31904, 16'd14270, 16'd13366, 16'd29807, 16'd44221, 16'd20593, 16'd1590, 16'd32732, 16'd53386, 16'd14189, 16'd18613, 16'd4931, 16'd43120, 16'd59415, 16'd47980, 16'd6712, 16'd20577, 16'd17601, 16'd49284});
	test_expansion(128'h0f1b53796a9696a08e3774497294d5f8, {16'd45460, 16'd40292, 16'd44840, 16'd34442, 16'd4962, 16'd14972, 16'd59260, 16'd20076, 16'd10043, 16'd26216, 16'd39356, 16'd26695, 16'd46437, 16'd40258, 16'd36851, 16'd6557, 16'd30210, 16'd23311, 16'd19284, 16'd63769, 16'd63503, 16'd1545, 16'd16324, 16'd10379, 16'd46580, 16'd28634});
	test_expansion(128'ha9c54e9698a58068b22a6314aa9bdfbb, {16'd56544, 16'd21671, 16'd45319, 16'd44737, 16'd18696, 16'd12973, 16'd41716, 16'd7710, 16'd49343, 16'd55540, 16'd45307, 16'd13945, 16'd54611, 16'd58252, 16'd53042, 16'd20795, 16'd29500, 16'd30390, 16'd3903, 16'd62217, 16'd42127, 16'd65384, 16'd37027, 16'd34716, 16'd18308, 16'd30258});
	test_expansion(128'hf0f812754e5ca151951160a598378ebd, {16'd35176, 16'd65042, 16'd29273, 16'd51758, 16'd32672, 16'd62365, 16'd62763, 16'd5111, 16'd43861, 16'd12404, 16'd10758, 16'd51346, 16'd32137, 16'd50838, 16'd27905, 16'd58645, 16'd32618, 16'd48920, 16'd44822, 16'd52611, 16'd25168, 16'd25125, 16'd13845, 16'd19444, 16'd5268, 16'd45535});
	test_expansion(128'h67117a94f0c29e54f55cc70ee2c626b9, {16'd25539, 16'd2826, 16'd21431, 16'd26494, 16'd43329, 16'd51149, 16'd29785, 16'd29544, 16'd25598, 16'd47868, 16'd17723, 16'd24175, 16'd29630, 16'd8689, 16'd59179, 16'd37128, 16'd37528, 16'd15354, 16'd56997, 16'd52118, 16'd23023, 16'd6507, 16'd50163, 16'd52141, 16'd55946, 16'd53611});
	test_expansion(128'h6f3a2f704640c27165e77e747125affa, {16'd52749, 16'd15312, 16'd60358, 16'd59047, 16'd24178, 16'd11433, 16'd39792, 16'd61043, 16'd25500, 16'd15969, 16'd16306, 16'd15517, 16'd56298, 16'd9064, 16'd57371, 16'd36991, 16'd18090, 16'd32111, 16'd54837, 16'd54570, 16'd27600, 16'd31785, 16'd28038, 16'd52210, 16'd4461, 16'd55182});
	test_expansion(128'hd4540b9699e877cfa9b8e1ce62680e6d, {16'd15609, 16'd4822, 16'd339, 16'd6240, 16'd4931, 16'd53574, 16'd54714, 16'd62808, 16'd33595, 16'd43316, 16'd17051, 16'd28808, 16'd17850, 16'd44736, 16'd60968, 16'd8766, 16'd10741, 16'd59565, 16'd32451, 16'd14812, 16'd62828, 16'd53052, 16'd42146, 16'd28531, 16'd6422, 16'd50490});
	test_expansion(128'h28af78e01c4dba1e62d3e7c57c49070c, {16'd59100, 16'd41495, 16'd36884, 16'd53290, 16'd47995, 16'd43554, 16'd10741, 16'd40325, 16'd23764, 16'd58073, 16'd59291, 16'd56526, 16'd47879, 16'd513, 16'd60466, 16'd34304, 16'd36755, 16'd1698, 16'd54342, 16'd22882, 16'd13150, 16'd42479, 16'd62399, 16'd26687, 16'd9960, 16'd61528});
	test_expansion(128'hf952b4e7994245f1126bbba9c9ce58dd, {16'd49388, 16'd1591, 16'd54888, 16'd54046, 16'd45938, 16'd37119, 16'd11621, 16'd27481, 16'd16440, 16'd1108, 16'd54327, 16'd64473, 16'd17299, 16'd17975, 16'd48500, 16'd21926, 16'd54197, 16'd55022, 16'd19293, 16'd31624, 16'd16308, 16'd36456, 16'd20428, 16'd17180, 16'd41671, 16'd6962});
	test_expansion(128'h4ba9d06a91f2f8b34992b6544c8b9d74, {16'd60134, 16'd38514, 16'd45831, 16'd40437, 16'd35808, 16'd50583, 16'd24338, 16'd52792, 16'd27856, 16'd2802, 16'd39143, 16'd14906, 16'd29966, 16'd63963, 16'd38973, 16'd64110, 16'd8035, 16'd38400, 16'd1402, 16'd22685, 16'd7713, 16'd42179, 16'd1511, 16'd5782, 16'd32962, 16'd28987});
	test_expansion(128'h1b5a9d7d2764f5367609fd7e2000543b, {16'd5921, 16'd5065, 16'd37707, 16'd36757, 16'd35995, 16'd64341, 16'd49074, 16'd59287, 16'd48559, 16'd60695, 16'd20284, 16'd51362, 16'd46726, 16'd27322, 16'd10960, 16'd24445, 16'd38756, 16'd8798, 16'd21102, 16'd131, 16'd10753, 16'd47958, 16'd524, 16'd49497, 16'd38342, 16'd4879});
	test_expansion(128'h10f958486142eca45c8900558baa5265, {16'd15500, 16'd19685, 16'd64991, 16'd2696, 16'd29338, 16'd11113, 16'd41725, 16'd19186, 16'd4963, 16'd13973, 16'd12134, 16'd57276, 16'd6747, 16'd5698, 16'd57506, 16'd59924, 16'd20756, 16'd37342, 16'd25234, 16'd28250, 16'd22921, 16'd63787, 16'd37536, 16'd2155, 16'd6041, 16'd6620});
	test_expansion(128'hcff61ffa7c41dbae8ce595acd047cd81, {16'd40516, 16'd20739, 16'd1576, 16'd11795, 16'd59143, 16'd9632, 16'd64293, 16'd30436, 16'd26996, 16'd15342, 16'd45106, 16'd45092, 16'd1867, 16'd64429, 16'd29524, 16'd53053, 16'd60548, 16'd2949, 16'd6768, 16'd55739, 16'd40940, 16'd25146, 16'd39743, 16'd61514, 16'd23981, 16'd1838});
	test_expansion(128'h860706894a780c0215871e496979ee7a, {16'd59817, 16'd3831, 16'd23134, 16'd58649, 16'd26495, 16'd51839, 16'd33503, 16'd57518, 16'd13514, 16'd34328, 16'd19213, 16'd53112, 16'd9027, 16'd24891, 16'd46455, 16'd42251, 16'd32648, 16'd28018, 16'd61864, 16'd58461, 16'd55173, 16'd6488, 16'd30808, 16'd37747, 16'd33049, 16'd40334});
	test_expansion(128'hf85390fb8d33ac2f5291cc6c8320f386, {16'd30871, 16'd2834, 16'd44459, 16'd52436, 16'd30421, 16'd11202, 16'd12251, 16'd29050, 16'd14196, 16'd62245, 16'd15784, 16'd55765, 16'd64986, 16'd29151, 16'd15885, 16'd333, 16'd41389, 16'd45551, 16'd2459, 16'd58716, 16'd30876, 16'd40220, 16'd41841, 16'd28283, 16'd2333, 16'd48719});
	test_expansion(128'hf9b2d9c0aca3190551105b6fa8013137, {16'd19744, 16'd38933, 16'd745, 16'd920, 16'd65137, 16'd36828, 16'd53828, 16'd28712, 16'd18122, 16'd48202, 16'd59540, 16'd25336, 16'd60264, 16'd21582, 16'd54, 16'd16143, 16'd10159, 16'd62851, 16'd64257, 16'd64386, 16'd4804, 16'd8404, 16'd64889, 16'd26877, 16'd54527, 16'd56474});
	test_expansion(128'h511b509fa0253b1177d1976d35755b95, {16'd19582, 16'd32320, 16'd61751, 16'd44604, 16'd17968, 16'd55989, 16'd11014, 16'd46206, 16'd2117, 16'd49530, 16'd5658, 16'd65374, 16'd34257, 16'd42786, 16'd39042, 16'd51637, 16'd2227, 16'd28781, 16'd25567, 16'd27254, 16'd41596, 16'd52690, 16'd40072, 16'd15028, 16'd27293, 16'd3906});
	test_expansion(128'hb77544597881d988f9a49efb58fd9928, {16'd37325, 16'd50682, 16'd34409, 16'd1736, 16'd11195, 16'd17158, 16'd1399, 16'd17461, 16'd26750, 16'd10109, 16'd32940, 16'd57902, 16'd34125, 16'd20522, 16'd59876, 16'd47345, 16'd24478, 16'd5351, 16'd47641, 16'd38726, 16'd23726, 16'd59850, 16'd40682, 16'd62889, 16'd26176, 16'd24225});
	test_expansion(128'hd5bee86c16e52fb763bcf86970bf0987, {16'd29180, 16'd39550, 16'd30244, 16'd30118, 16'd59395, 16'd59564, 16'd57925, 16'd33283, 16'd1234, 16'd42305, 16'd17728, 16'd52337, 16'd61986, 16'd16125, 16'd13094, 16'd29878, 16'd50669, 16'd27554, 16'd53003, 16'd5775, 16'd40875, 16'd18068, 16'd17131, 16'd4983, 16'd32449, 16'd1702});
	test_expansion(128'h9c7334507e7c9eff23589fc96c4b86cd, {16'd42629, 16'd47194, 16'd22593, 16'd48496, 16'd45695, 16'd14523, 16'd41069, 16'd56209, 16'd5296, 16'd52308, 16'd57019, 16'd11068, 16'd38840, 16'd4875, 16'd51111, 16'd42939, 16'd63241, 16'd61031, 16'd14114, 16'd35842, 16'd61746, 16'd29841, 16'd30145, 16'd46148, 16'd47033, 16'd56254});
	test_expansion(128'hf947f3d6a0e68c26be386a21f63e180e, {16'd53707, 16'd17531, 16'd22616, 16'd6279, 16'd2995, 16'd63123, 16'd60034, 16'd26311, 16'd1173, 16'd25129, 16'd22540, 16'd2909, 16'd36050, 16'd44402, 16'd11785, 16'd52364, 16'd60029, 16'd63228, 16'd16111, 16'd8912, 16'd58645, 16'd56964, 16'd51180, 16'd5293, 16'd33154, 16'd43883});
	test_expansion(128'h51bf4e78259f53b5716cf5b2982ec59c, {16'd26086, 16'd2918, 16'd20909, 16'd63042, 16'd25462, 16'd36165, 16'd17233, 16'd43033, 16'd9289, 16'd46057, 16'd62919, 16'd61241, 16'd1723, 16'd37253, 16'd62297, 16'd55689, 16'd46907, 16'd1130, 16'd15914, 16'd64442, 16'd43405, 16'd20604, 16'd58327, 16'd12522, 16'd52839, 16'd53780});
	test_expansion(128'hd8b337a5e4f289a009abac8c817bf454, {16'd919, 16'd15971, 16'd7038, 16'd61185, 16'd21115, 16'd65377, 16'd38411, 16'd50771, 16'd29242, 16'd9807, 16'd46542, 16'd59260, 16'd31434, 16'd44540, 16'd56544, 16'd58403, 16'd4499, 16'd7941, 16'd5585, 16'd13591, 16'd30872, 16'd25176, 16'd37478, 16'd8685, 16'd38485, 16'd28727});
	test_expansion(128'h1ed895239ea5729c7038c9de23d8f515, {16'd49885, 16'd31611, 16'd22906, 16'd2525, 16'd217, 16'd30486, 16'd40333, 16'd27217, 16'd39580, 16'd4916, 16'd39716, 16'd4282, 16'd19696, 16'd57426, 16'd27718, 16'd11558, 16'd24886, 16'd38717, 16'd17463, 16'd46487, 16'd55042, 16'd41674, 16'd40042, 16'd47256, 16'd21311, 16'd8049});
	test_expansion(128'he6d4b69e614c73b4405828682786348d, {16'd3359, 16'd33371, 16'd18213, 16'd58341, 16'd46217, 16'd59060, 16'd46206, 16'd7255, 16'd61939, 16'd1352, 16'd52930, 16'd44204, 16'd37244, 16'd57410, 16'd27556, 16'd55667, 16'd57186, 16'd10601, 16'd57404, 16'd35439, 16'd60395, 16'd12287, 16'd20528, 16'd10352, 16'd52016, 16'd8434});
	test_expansion(128'h727df3d9292091fd09b0d660015d5f5a, {16'd51070, 16'd56874, 16'd65204, 16'd47183, 16'd9600, 16'd11776, 16'd12057, 16'd58350, 16'd18620, 16'd41753, 16'd22700, 16'd16608, 16'd51748, 16'd38615, 16'd5091, 16'd33876, 16'd30884, 16'd52005, 16'd27914, 16'd3520, 16'd753, 16'd29718, 16'd54774, 16'd57742, 16'd63160, 16'd6098});
	test_expansion(128'h9e7f7c4b3826290c6d648d458f61860f, {16'd45992, 16'd30398, 16'd60198, 16'd59850, 16'd34241, 16'd24923, 16'd44460, 16'd27777, 16'd34025, 16'd1642, 16'd10909, 16'd2903, 16'd34748, 16'd23737, 16'd62167, 16'd53479, 16'd18693, 16'd61331, 16'd12812, 16'd19470, 16'd15975, 16'd8862, 16'd55927, 16'd23736, 16'd51762, 16'd43042});
	test_expansion(128'h507b4dc9d32e916067f81503f1c8e6a3, {16'd49804, 16'd46386, 16'd6098, 16'd64178, 16'd3757, 16'd59757, 16'd36752, 16'd19327, 16'd61360, 16'd35913, 16'd1655, 16'd58455, 16'd57462, 16'd57569, 16'd27727, 16'd47847, 16'd65102, 16'd34683, 16'd46083, 16'd64129, 16'd40150, 16'd30576, 16'd65343, 16'd35327, 16'd18184, 16'd12165});
	test_expansion(128'hd3a0cbe59ff8f407924a60c58c5c62fc, {16'd64285, 16'd34634, 16'd44664, 16'd47095, 16'd48, 16'd48252, 16'd32030, 16'd6606, 16'd45693, 16'd37116, 16'd2744, 16'd33094, 16'd18034, 16'd47755, 16'd13389, 16'd4590, 16'd13279, 16'd11418, 16'd49975, 16'd16306, 16'd44381, 16'd8125, 16'd63578, 16'd19592, 16'd24309, 16'd22166});
	test_expansion(128'hb30878906931e7a509a087db88b0a23c, {16'd22013, 16'd49322, 16'd51641, 16'd39122, 16'd23484, 16'd57150, 16'd57770, 16'd50697, 16'd37399, 16'd44669, 16'd24436, 16'd15364, 16'd51819, 16'd3064, 16'd60277, 16'd38196, 16'd4010, 16'd50332, 16'd27048, 16'd31953, 16'd38445, 16'd19871, 16'd61688, 16'd36229, 16'd21068, 16'd28160});
	test_expansion(128'hf2acb9d3d8d6fe268466003a0901e969, {16'd9768, 16'd55770, 16'd15816, 16'd61018, 16'd11927, 16'd36512, 16'd9970, 16'd10434, 16'd39367, 16'd47188, 16'd35485, 16'd55831, 16'd60588, 16'd62908, 16'd58507, 16'd38410, 16'd28967, 16'd49427, 16'd2270, 16'd64536, 16'd46794, 16'd13482, 16'd37043, 16'd6416, 16'd29764, 16'd30616});
	test_expansion(128'h037e36699f721248f19918b5d2f8666a, {16'd13180, 16'd52249, 16'd32130, 16'd38418, 16'd25367, 16'd21314, 16'd59435, 16'd37658, 16'd56625, 16'd4648, 16'd38386, 16'd64180, 16'd16685, 16'd16215, 16'd34658, 16'd15050, 16'd19159, 16'd38936, 16'd47820, 16'd25163, 16'd2528, 16'd9508, 16'd43488, 16'd59484, 16'd62453, 16'd65072});
	test_expansion(128'h08f4872437e55262f7e0c00b86cee16c, {16'd50115, 16'd63005, 16'd53394, 16'd57395, 16'd33323, 16'd7471, 16'd57510, 16'd52841, 16'd8367, 16'd50493, 16'd7940, 16'd49113, 16'd57665, 16'd11820, 16'd33465, 16'd54646, 16'd32756, 16'd65196, 16'd22723, 16'd14357, 16'd7211, 16'd5445, 16'd37656, 16'd35514, 16'd15316, 16'd64723});
	test_expansion(128'h9f64603a1ed6003ba2c201dfc723b0e7, {16'd27269, 16'd43940, 16'd13311, 16'd60242, 16'd61961, 16'd57514, 16'd64976, 16'd41445, 16'd12113, 16'd36482, 16'd38196, 16'd60842, 16'd23581, 16'd59343, 16'd14134, 16'd40529, 16'd17592, 16'd2907, 16'd25734, 16'd21693, 16'd18674, 16'd21901, 16'd26824, 16'd36665, 16'd17573, 16'd24757});
	test_expansion(128'hcd49470bd3ca61a87b2495a20ea14b0b, {16'd64923, 16'd51561, 16'd36492, 16'd49697, 16'd25315, 16'd33020, 16'd44293, 16'd21834, 16'd38257, 16'd11631, 16'd40929, 16'd47457, 16'd44040, 16'd50981, 16'd64845, 16'd18145, 16'd31126, 16'd24161, 16'd23376, 16'd47749, 16'd32995, 16'd56635, 16'd21345, 16'd48379, 16'd3106, 16'd21190});
	test_expansion(128'h3ed03987b277ade1c2fe257c68fad73e, {16'd39297, 16'd910, 16'd51177, 16'd45795, 16'd60731, 16'd35643, 16'd15936, 16'd22088, 16'd20104, 16'd16429, 16'd26154, 16'd19518, 16'd52899, 16'd48399, 16'd49238, 16'd48066, 16'd28040, 16'd10782, 16'd57518, 16'd15851, 16'd42647, 16'd7029, 16'd22759, 16'd18601, 16'd5668, 16'd63828});
	test_expansion(128'hb25fe80a4a1da229eecbb467a4baa4f6, {16'd37535, 16'd24315, 16'd29077, 16'd15072, 16'd3769, 16'd27756, 16'd29204, 16'd14838, 16'd48228, 16'd27392, 16'd13657, 16'd13906, 16'd64689, 16'd56802, 16'd7383, 16'd40696, 16'd16401, 16'd7053, 16'd214, 16'd62122, 16'd4322, 16'd11407, 16'd542, 16'd19859, 16'd24810, 16'd52732});
	test_expansion(128'he312330e54ba870dace49e25fb968d7f, {16'd63792, 16'd3098, 16'd27166, 16'd30366, 16'd3612, 16'd2403, 16'd40587, 16'd50119, 16'd48878, 16'd1184, 16'd57693, 16'd14567, 16'd32086, 16'd12387, 16'd26792, 16'd17221, 16'd59776, 16'd37087, 16'd2858, 16'd14843, 16'd37353, 16'd63605, 16'd1874, 16'd48670, 16'd29776, 16'd61248});
	test_expansion(128'hd93c977a3a4edf9eb4a4eb3c29ac8105, {16'd60273, 16'd52577, 16'd50764, 16'd62565, 16'd37452, 16'd65321, 16'd38142, 16'd51820, 16'd51060, 16'd34746, 16'd17738, 16'd28426, 16'd14871, 16'd40315, 16'd64963, 16'd19822, 16'd50533, 16'd51037, 16'd62004, 16'd21806, 16'd41801, 16'd9970, 16'd45381, 16'd59934, 16'd17219, 16'd29943});
	test_expansion(128'hb59288188fde959218a7bc6275b7c5fd, {16'd31988, 16'd64481, 16'd43083, 16'd64400, 16'd19885, 16'd50754, 16'd16303, 16'd28627, 16'd53506, 16'd44963, 16'd2059, 16'd27264, 16'd8819, 16'd43039, 16'd23866, 16'd30976, 16'd6165, 16'd54689, 16'd40145, 16'd4513, 16'd13039, 16'd56881, 16'd31512, 16'd31428, 16'd24402, 16'd36020});
	test_expansion(128'h7640e836611d100181353b1ffa28baee, {16'd31508, 16'd46845, 16'd46726, 16'd60569, 16'd5340, 16'd21799, 16'd49431, 16'd433, 16'd38386, 16'd63932, 16'd32358, 16'd9908, 16'd1909, 16'd52938, 16'd4254, 16'd25987, 16'd21774, 16'd32931, 16'd4721, 16'd51113, 16'd44759, 16'd49228, 16'd22564, 16'd61319, 16'd9194, 16'd54780});
	test_expansion(128'h2c662b4ff2a300d9a061833bd9441645, {16'd53596, 16'd15865, 16'd18956, 16'd25864, 16'd39772, 16'd4877, 16'd23346, 16'd23662, 16'd7306, 16'd25526, 16'd16448, 16'd42798, 16'd11043, 16'd24598, 16'd19748, 16'd46073, 16'd34844, 16'd20136, 16'd50029, 16'd21460, 16'd40973, 16'd13580, 16'd53492, 16'd14183, 16'd26915, 16'd20462});
	test_expansion(128'heae77ecca19af2a6739cc17d1bbb7e80, {16'd38473, 16'd58932, 16'd25207, 16'd21229, 16'd30242, 16'd40626, 16'd56963, 16'd58248, 16'd40469, 16'd36579, 16'd37185, 16'd8685, 16'd55919, 16'd58426, 16'd30808, 16'd3708, 16'd37005, 16'd38506, 16'd22089, 16'd50260, 16'd2745, 16'd14394, 16'd62661, 16'd29224, 16'd4882, 16'd16462});
	test_expansion(128'h92a25faac781a6d25801250417e1640f, {16'd43393, 16'd10599, 16'd56809, 16'd3681, 16'd32631, 16'd32358, 16'd18712, 16'd42494, 16'd17202, 16'd418, 16'd39716, 16'd19097, 16'd5289, 16'd23912, 16'd63464, 16'd7785, 16'd483, 16'd54766, 16'd38638, 16'd19097, 16'd35475, 16'd48799, 16'd24173, 16'd18549, 16'd18549, 16'd50553});
	test_expansion(128'h5cc75a3fbd8bcb84da6d6916b01f3d10, {16'd22314, 16'd51202, 16'd2151, 16'd30599, 16'd41972, 16'd57616, 16'd26259, 16'd1128, 16'd24154, 16'd56853, 16'd24146, 16'd23313, 16'd31821, 16'd41443, 16'd31055, 16'd38398, 16'd9159, 16'd61166, 16'd38086, 16'd8980, 16'd39267, 16'd31948, 16'd28151, 16'd15990, 16'd33472, 16'd46233});
	test_expansion(128'h1d780ffefed7f097f6dc38c063601801, {16'd52360, 16'd12190, 16'd11477, 16'd553, 16'd63750, 16'd23855, 16'd37796, 16'd5487, 16'd37464, 16'd57450, 16'd17628, 16'd53660, 16'd44963, 16'd28958, 16'd36, 16'd25140, 16'd6552, 16'd1720, 16'd43878, 16'd5322, 16'd23383, 16'd42275, 16'd42439, 16'd16247, 16'd39213, 16'd47711});
	test_expansion(128'hd4d31b8a88bdabd1521d2967ecf6e47e, {16'd26483, 16'd15181, 16'd1658, 16'd34430, 16'd60087, 16'd47622, 16'd20897, 16'd1730, 16'd63158, 16'd51555, 16'd31608, 16'd9897, 16'd30515, 16'd45621, 16'd59618, 16'd45120, 16'd49128, 16'd30507, 16'd24679, 16'd49502, 16'd36978, 16'd63633, 16'd31565, 16'd38313, 16'd41532, 16'd53717});
	test_expansion(128'h94c89dbd10c0291d119746a2b27ce4d2, {16'd29030, 16'd61044, 16'd24638, 16'd35167, 16'd61312, 16'd64025, 16'd50336, 16'd54429, 16'd64550, 16'd19920, 16'd61577, 16'd37868, 16'd15674, 16'd30408, 16'd14314, 16'd30052, 16'd17583, 16'd5066, 16'd52785, 16'd52981, 16'd60873, 16'd15065, 16'd23989, 16'd22014, 16'd14520, 16'd28375});
	test_expansion(128'hca7c4dcce2b656899a3951db111b7191, {16'd30640, 16'd28123, 16'd56930, 16'd19644, 16'd27721, 16'd47283, 16'd39606, 16'd30998, 16'd17697, 16'd53873, 16'd24090, 16'd28345, 16'd10031, 16'd61793, 16'd24345, 16'd26787, 16'd36876, 16'd43679, 16'd40499, 16'd60471, 16'd22345, 16'd50521, 16'd45321, 16'd5892, 16'd26542, 16'd10566});
	test_expansion(128'h498760c4d3b3cbdc7cb75b8c1f52245d, {16'd1924, 16'd54777, 16'd60486, 16'd4306, 16'd17899, 16'd59040, 16'd40325, 16'd41028, 16'd7143, 16'd58579, 16'd53360, 16'd60163, 16'd44689, 16'd59758, 16'd41896, 16'd46592, 16'd51586, 16'd37586, 16'd64142, 16'd10295, 16'd22779, 16'd48005, 16'd60026, 16'd24044, 16'd41022, 16'd1326});
	test_expansion(128'h46a92125fc243577abda3e361ea46468, {16'd52352, 16'd45153, 16'd5843, 16'd46573, 16'd11592, 16'd23209, 16'd63671, 16'd39278, 16'd46888, 16'd29454, 16'd39345, 16'd28716, 16'd29324, 16'd60009, 16'd13063, 16'd32244, 16'd324, 16'd53402, 16'd17182, 16'd38991, 16'd4045, 16'd38733, 16'd39560, 16'd25846, 16'd34302, 16'd46368});
	test_expansion(128'had0367de8c63db7729bca34bc5f5dab0, {16'd49251, 16'd49319, 16'd43018, 16'd50348, 16'd64190, 16'd55436, 16'd13367, 16'd52909, 16'd65389, 16'd26329, 16'd12081, 16'd31929, 16'd8062, 16'd7279, 16'd24424, 16'd31435, 16'd10321, 16'd53305, 16'd31134, 16'd12273, 16'd44865, 16'd19708, 16'd45667, 16'd32026, 16'd62935, 16'd6851});
	test_expansion(128'h806775c1ee190513b83155b18b920433, {16'd29135, 16'd7480, 16'd39204, 16'd5738, 16'd4136, 16'd40699, 16'd63544, 16'd56495, 16'd18787, 16'd46782, 16'd17469, 16'd65109, 16'd51293, 16'd57249, 16'd64729, 16'd32099, 16'd40554, 16'd36903, 16'd56435, 16'd3026, 16'd48910, 16'd56955, 16'd63323, 16'd61032, 16'd20941, 16'd5672});
	test_expansion(128'h51569c3c0d7fb1fb953f743bf75a8f21, {16'd56233, 16'd31666, 16'd28872, 16'd22495, 16'd61651, 16'd64812, 16'd62836, 16'd49189, 16'd23535, 16'd4191, 16'd35676, 16'd40598, 16'd45475, 16'd56243, 16'd10586, 16'd13302, 16'd8876, 16'd28027, 16'd26801, 16'd4189, 16'd49651, 16'd38102, 16'd60260, 16'd24690, 16'd50008, 16'd36746});
	test_expansion(128'hc49b6b061acf1375fda709b2fb32a6ac, {16'd15174, 16'd58122, 16'd6881, 16'd19866, 16'd62614, 16'd52155, 16'd20845, 16'd58751, 16'd60890, 16'd5821, 16'd28290, 16'd17743, 16'd60848, 16'd13832, 16'd39411, 16'd20541, 16'd53094, 16'd16217, 16'd32819, 16'd39575, 16'd31244, 16'd20088, 16'd55907, 16'd41317, 16'd40069, 16'd35679});
	test_expansion(128'h1dbc93902c3f7dcbf36bc60cb59833b5, {16'd23248, 16'd46309, 16'd1315, 16'd37850, 16'd31137, 16'd52957, 16'd6786, 16'd42288, 16'd44049, 16'd2775, 16'd56183, 16'd9636, 16'd33353, 16'd36645, 16'd21569, 16'd52067, 16'd28601, 16'd3602, 16'd38856, 16'd47967, 16'd7734, 16'd45671, 16'd54157, 16'd57799, 16'd32127, 16'd62114});
	test_expansion(128'h9234b864fecd69e8c3210b33c624412a, {16'd54117, 16'd25759, 16'd39670, 16'd42687, 16'd56671, 16'd7209, 16'd6066, 16'd51739, 16'd7212, 16'd31875, 16'd58778, 16'd23009, 16'd27162, 16'd59973, 16'd3186, 16'd6037, 16'd19487, 16'd55881, 16'd40518, 16'd6291, 16'd62477, 16'd35642, 16'd52604, 16'd3111, 16'd48224, 16'd40490});
	test_expansion(128'hc2cc17e8434bf63fb1a52dd225fd9bf6, {16'd53457, 16'd51358, 16'd5162, 16'd56811, 16'd9478, 16'd26857, 16'd44794, 16'd42922, 16'd38628, 16'd14578, 16'd10078, 16'd25525, 16'd40612, 16'd65159, 16'd43623, 16'd16545, 16'd49072, 16'd47714, 16'd64631, 16'd10207, 16'd34133, 16'd3545, 16'd35199, 16'd51268, 16'd64050, 16'd3989});
	test_expansion(128'hd2180bc74f87afb988a0071757a5c462, {16'd11867, 16'd34634, 16'd41034, 16'd45612, 16'd19128, 16'd54441, 16'd20285, 16'd50332, 16'd36325, 16'd60413, 16'd63396, 16'd48313, 16'd223, 16'd61724, 16'd61764, 16'd36763, 16'd3428, 16'd11408, 16'd5412, 16'd7196, 16'd43851, 16'd9550, 16'd37527, 16'd29187, 16'd19218, 16'd14805});
	test_expansion(128'h3608489a4671b54ec8bb1d64af3793fd, {16'd49301, 16'd18136, 16'd196, 16'd60323, 16'd37374, 16'd46722, 16'd50801, 16'd52248, 16'd13985, 16'd4745, 16'd9888, 16'd12981, 16'd29790, 16'd44624, 16'd9528, 16'd21644, 16'd19165, 16'd28403, 16'd54771, 16'd60587, 16'd34019, 16'd703, 16'd38977, 16'd16189, 16'd62963, 16'd13684});
	test_expansion(128'h955f3c0a6d2d5b87ea5b0fd69a4ffc2c, {16'd25673, 16'd42376, 16'd32600, 16'd64454, 16'd17311, 16'd63944, 16'd63222, 16'd478, 16'd58682, 16'd35631, 16'd21883, 16'd30260, 16'd30894, 16'd35717, 16'd15771, 16'd29023, 16'd56048, 16'd31247, 16'd21579, 16'd31642, 16'd52504, 16'd24765, 16'd58191, 16'd1421, 16'd1002, 16'd48450});
	test_expansion(128'h567db4ca39c53d058b37df8cb29019d3, {16'd52761, 16'd37206, 16'd37038, 16'd34264, 16'd57198, 16'd37928, 16'd24158, 16'd37111, 16'd55711, 16'd59287, 16'd25728, 16'd10928, 16'd16707, 16'd27722, 16'd30871, 16'd51599, 16'd51223, 16'd53868, 16'd32348, 16'd38297, 16'd60896, 16'd29658, 16'd56052, 16'd52374, 16'd16504, 16'd7042});
	test_expansion(128'hdc9bbc27293a1f58ec4306267ad48556, {16'd47669, 16'd47550, 16'd39773, 16'd49027, 16'd32997, 16'd26878, 16'd15498, 16'd36556, 16'd2871, 16'd21299, 16'd14557, 16'd36033, 16'd21477, 16'd1135, 16'd28615, 16'd7683, 16'd47166, 16'd26781, 16'd30999, 16'd22110, 16'd10580, 16'd45106, 16'd3417, 16'd58043, 16'd27852, 16'd58997});
	test_expansion(128'hc2cfa9be773d86f98688dd1cdfcdb075, {16'd33471, 16'd9680, 16'd6973, 16'd31268, 16'd25863, 16'd10151, 16'd3218, 16'd55091, 16'd25511, 16'd41062, 16'd18662, 16'd60269, 16'd27024, 16'd44830, 16'd51650, 16'd39889, 16'd56189, 16'd48959, 16'd41872, 16'd14557, 16'd27880, 16'd50515, 16'd32777, 16'd2827, 16'd23661, 16'd16268});
	test_expansion(128'h1fdf020848ab3f5978ac970a0538951a, {16'd35269, 16'd41002, 16'd64306, 16'd55385, 16'd30916, 16'd43022, 16'd17824, 16'd48375, 16'd26863, 16'd58265, 16'd53035, 16'd46357, 16'd55920, 16'd26756, 16'd5300, 16'd49694, 16'd26942, 16'd8548, 16'd50257, 16'd40923, 16'd28594, 16'd6382, 16'd41540, 16'd62446, 16'd31456, 16'd41708});
	test_expansion(128'h36559e506b553d00cbea7cf9d88fc3b1, {16'd36418, 16'd15125, 16'd4510, 16'd31001, 16'd8143, 16'd8277, 16'd63854, 16'd63804, 16'd56767, 16'd6984, 16'd13792, 16'd46767, 16'd52966, 16'd48807, 16'd26548, 16'd60401, 16'd3090, 16'd13506, 16'd15310, 16'd15221, 16'd43440, 16'd45095, 16'd14872, 16'd64315, 16'd9664, 16'd14951});
	test_expansion(128'hcccee7d55c9cfb07ede4475bd639fdda, {16'd40800, 16'd32507, 16'd18040, 16'd28888, 16'd44004, 16'd38421, 16'd36762, 16'd54549, 16'd28723, 16'd20464, 16'd3463, 16'd19750, 16'd51116, 16'd33616, 16'd29971, 16'd2344, 16'd23496, 16'd53491, 16'd16408, 16'd41764, 16'd2213, 16'd29874, 16'd56933, 16'd38605, 16'd11295, 16'd1983});
	test_expansion(128'he96be4c4236ee90f177cd21434eb1858, {16'd11472, 16'd9570, 16'd40690, 16'd53137, 16'd11512, 16'd62835, 16'd33679, 16'd56306, 16'd6447, 16'd33946, 16'd5793, 16'd14603, 16'd23584, 16'd36247, 16'd27552, 16'd57745, 16'd59883, 16'd63734, 16'd2417, 16'd64362, 16'd19295, 16'd58262, 16'd833, 16'd51087, 16'd60500, 16'd44721});
	test_expansion(128'hc02a29c51a0dff77d8564047ed685b86, {16'd35766, 16'd32309, 16'd61385, 16'd61166, 16'd41329, 16'd28514, 16'd16716, 16'd37517, 16'd27940, 16'd32332, 16'd35158, 16'd23213, 16'd23148, 16'd27422, 16'd51476, 16'd50689, 16'd22626, 16'd27183, 16'd51085, 16'd7758, 16'd24728, 16'd46375, 16'd28678, 16'd34725, 16'd36205, 16'd45329});
	test_expansion(128'h7b7c2fc3c9c9aa82de88462388575e6f, {16'd58526, 16'd9555, 16'd6921, 16'd54263, 16'd9750, 16'd18510, 16'd26301, 16'd171, 16'd43414, 16'd61890, 16'd53404, 16'd65461, 16'd53609, 16'd36454, 16'd51457, 16'd4724, 16'd17831, 16'd16396, 16'd64685, 16'd1996, 16'd12627, 16'd64679, 16'd209, 16'd49260, 16'd4075, 16'd6049});
	test_expansion(128'hc887580d0a395998a1527174d09a58c9, {16'd41721, 16'd43547, 16'd26083, 16'd34788, 16'd6824, 16'd13708, 16'd11440, 16'd59649, 16'd58033, 16'd20216, 16'd12999, 16'd51237, 16'd37499, 16'd26521, 16'd22377, 16'd4382, 16'd37266, 16'd7315, 16'd28181, 16'd59501, 16'd37305, 16'd15124, 16'd1300, 16'd33991, 16'd657, 16'd34511});
	test_expansion(128'h0cd6e06f3d1f684309b72dbfd7a7d0ce, {16'd26203, 16'd11068, 16'd9526, 16'd65286, 16'd41506, 16'd8964, 16'd18421, 16'd17868, 16'd53389, 16'd62052, 16'd17135, 16'd58455, 16'd28819, 16'd27030, 16'd44591, 16'd14248, 16'd12184, 16'd54831, 16'd314, 16'd61640, 16'd22457, 16'd56654, 16'd25125, 16'd3297, 16'd60678, 16'd38424});
	test_expansion(128'h994a06c57efd550b285d6e79ef952c40, {16'd17578, 16'd35664, 16'd9527, 16'd8347, 16'd51736, 16'd44572, 16'd21834, 16'd24005, 16'd31583, 16'd6171, 16'd40757, 16'd28460, 16'd10767, 16'd45487, 16'd4, 16'd15384, 16'd52374, 16'd60147, 16'd60327, 16'd14790, 16'd36842, 16'd4140, 16'd13785, 16'd34155, 16'd54818, 16'd58462});
	test_expansion(128'h757aa5c0f7c9822af8dab3aa5710b76c, {16'd48728, 16'd14785, 16'd10393, 16'd11942, 16'd26886, 16'd61843, 16'd43159, 16'd27497, 16'd32951, 16'd48275, 16'd34699, 16'd11505, 16'd30266, 16'd23480, 16'd53175, 16'd47932, 16'd29338, 16'd34616, 16'd25801, 16'd52962, 16'd11664, 16'd55789, 16'd15422, 16'd51202, 16'd23746, 16'd40932});
	test_expansion(128'h013cf429a0bef5cad025609bcca7008d, {16'd50661, 16'd59808, 16'd29613, 16'd64504, 16'd4255, 16'd5839, 16'd31164, 16'd24296, 16'd33809, 16'd6468, 16'd18202, 16'd15758, 16'd866, 16'd374, 16'd13014, 16'd26808, 16'd62622, 16'd35460, 16'd10430, 16'd16442, 16'd20747, 16'd6606, 16'd47445, 16'd35176, 16'd23690, 16'd3843});
	test_expansion(128'h7001f4e7aed7b77eb00faab0453d0542, {16'd23586, 16'd31160, 16'd44513, 16'd13492, 16'd59930, 16'd54018, 16'd53555, 16'd57536, 16'd59172, 16'd53130, 16'd50393, 16'd20574, 16'd51915, 16'd53467, 16'd22846, 16'd10278, 16'd22519, 16'd48707, 16'd24296, 16'd2421, 16'd54033, 16'd3854, 16'd7363, 16'd59866, 16'd7808, 16'd32874});
	test_expansion(128'he0e12083d583bd9166d6e74d9d975004, {16'd54237, 16'd5711, 16'd29905, 16'd711, 16'd6525, 16'd9661, 16'd59678, 16'd18502, 16'd55424, 16'd64553, 16'd15053, 16'd8288, 16'd40305, 16'd50953, 16'd59397, 16'd34437, 16'd44215, 16'd23275, 16'd55722, 16'd4049, 16'd9118, 16'd64807, 16'd6934, 16'd23613, 16'd27838, 16'd18756});
	test_expansion(128'h9b72407d9407fa37e6ea52e5c1e43e1b, {16'd25904, 16'd18682, 16'd5856, 16'd30193, 16'd27717, 16'd39387, 16'd20375, 16'd50018, 16'd23552, 16'd38967, 16'd25153, 16'd13054, 16'd10063, 16'd37302, 16'd14023, 16'd20728, 16'd48888, 16'd47533, 16'd28988, 16'd65269, 16'd44406, 16'd15047, 16'd52147, 16'd39936, 16'd24089, 16'd11390});
	test_expansion(128'hbe5dcc84bca38b58cebc9e66b903f513, {16'd34864, 16'd52190, 16'd6831, 16'd13044, 16'd35748, 16'd7931, 16'd29767, 16'd17154, 16'd62476, 16'd59908, 16'd38825, 16'd57602, 16'd21729, 16'd51423, 16'd18285, 16'd9081, 16'd48850, 16'd26754, 16'd56907, 16'd22023, 16'd25097, 16'd54428, 16'd64278, 16'd25529, 16'd58077, 16'd56305});
	test_expansion(128'hf7ea165a0e71eaa431b8b084e0a5da1d, {16'd45513, 16'd11749, 16'd47193, 16'd12418, 16'd62934, 16'd24396, 16'd45509, 16'd20849, 16'd43321, 16'd35874, 16'd8793, 16'd23413, 16'd27369, 16'd34920, 16'd42343, 16'd20977, 16'd47156, 16'd54773, 16'd6924, 16'd52346, 16'd17676, 16'd1421, 16'd18563, 16'd52122, 16'd37433, 16'd41239});
	test_expansion(128'hb7672c2cf96849c141d67d5a410e38ac, {16'd63141, 16'd54298, 16'd26583, 16'd33535, 16'd9157, 16'd31172, 16'd15140, 16'd44542, 16'd60783, 16'd60709, 16'd36767, 16'd25849, 16'd58722, 16'd33865, 16'd50615, 16'd8884, 16'd14223, 16'd23825, 16'd53231, 16'd44895, 16'd26765, 16'd61707, 16'd38664, 16'd43943, 16'd40322, 16'd48632});
	test_expansion(128'h9243e8a76cc68b37824ee0b4f49d7c26, {16'd4704, 16'd12850, 16'd32109, 16'd57633, 16'd44008, 16'd21141, 16'd18550, 16'd57271, 16'd36947, 16'd62809, 16'd6561, 16'd13081, 16'd43434, 16'd64162, 16'd34361, 16'd51258, 16'd29732, 16'd43184, 16'd49239, 16'd57265, 16'd19212, 16'd19712, 16'd13802, 16'd61996, 16'd36460, 16'd55078});
	test_expansion(128'haed3a60586251c80b39e23b5c069583e, {16'd54251, 16'd62450, 16'd58349, 16'd17417, 16'd6435, 16'd64238, 16'd36884, 16'd48707, 16'd3111, 16'd27612, 16'd5980, 16'd22984, 16'd52388, 16'd7881, 16'd24515, 16'd26184, 16'd34864, 16'd52778, 16'd53435, 16'd35336, 16'd34791, 16'd4845, 16'd5690, 16'd7713, 16'd41874, 16'd47613});
	test_expansion(128'h763c1c063fde500f9e4766e9622f3f21, {16'd2233, 16'd13566, 16'd8774, 16'd34112, 16'd15301, 16'd7850, 16'd19556, 16'd23819, 16'd14390, 16'd59237, 16'd7729, 16'd25445, 16'd26109, 16'd40245, 16'd25271, 16'd44172, 16'd8078, 16'd8904, 16'd51623, 16'd12680, 16'd65468, 16'd14229, 16'd4633, 16'd45578, 16'd6944, 16'd62326});
	test_expansion(128'ha3fc62da1499243fed97b4ed2fcd6a67, {16'd48393, 16'd42538, 16'd25298, 16'd9617, 16'd53240, 16'd17001, 16'd9252, 16'd39060, 16'd55899, 16'd14772, 16'd36124, 16'd44359, 16'd16274, 16'd51971, 16'd20815, 16'd27565, 16'd35259, 16'd20656, 16'd31247, 16'd57006, 16'd39342, 16'd41508, 16'd7511, 16'd46996, 16'd31869, 16'd20426});
	test_expansion(128'h97f1b1bec651b34b8d2293f7a19cf4c3, {16'd1691, 16'd25176, 16'd63198, 16'd37466, 16'd29010, 16'd39527, 16'd37180, 16'd11132, 16'd28005, 16'd29787, 16'd30987, 16'd53757, 16'd31751, 16'd26660, 16'd59573, 16'd63352, 16'd62995, 16'd9130, 16'd1498, 16'd15082, 16'd60666, 16'd43571, 16'd64437, 16'd49932, 16'd61355, 16'd25374});
	test_expansion(128'h1aa87f7211ace23955fc6808a52ae140, {16'd38349, 16'd28604, 16'd64107, 16'd65301, 16'd40796, 16'd35988, 16'd31438, 16'd8542, 16'd37610, 16'd36329, 16'd51639, 16'd33281, 16'd30262, 16'd61680, 16'd35063, 16'd41, 16'd56152, 16'd49432, 16'd8152, 16'd35988, 16'd23864, 16'd25723, 16'd49468, 16'd63809, 16'd35169, 16'd20003});
	test_expansion(128'h251ff19dd4abadf8367407ae2525cf85, {16'd37194, 16'd5107, 16'd48719, 16'd23692, 16'd36384, 16'd28048, 16'd36861, 16'd39979, 16'd51977, 16'd54349, 16'd52485, 16'd49562, 16'd2785, 16'd56984, 16'd21028, 16'd44672, 16'd60583, 16'd7680, 16'd4906, 16'd39451, 16'd1956, 16'd41210, 16'd11368, 16'd23365, 16'd38147, 16'd40393});
	test_expansion(128'hb46c0e2ef3ccde602827f9f54b1c9981, {16'd42456, 16'd36581, 16'd3887, 16'd2455, 16'd11267, 16'd47446, 16'd11798, 16'd58320, 16'd34898, 16'd19509, 16'd25277, 16'd21270, 16'd49964, 16'd6519, 16'd54155, 16'd59199, 16'd24340, 16'd61970, 16'd6431, 16'd26476, 16'd23073, 16'd58655, 16'd60210, 16'd17723, 16'd18022, 16'd61155});
	test_expansion(128'h0654d6790ccd551ac5c57f6f96367656, {16'd39300, 16'd46444, 16'd6418, 16'd58239, 16'd16278, 16'd58372, 16'd38328, 16'd44630, 16'd6751, 16'd19765, 16'd10407, 16'd11996, 16'd60540, 16'd21829, 16'd41725, 16'd45692, 16'd58412, 16'd44094, 16'd18290, 16'd1844, 16'd5576, 16'd11312, 16'd12177, 16'd14547, 16'd37682, 16'd44365});
	test_expansion(128'h396415c7a5946bbffa2b55c313169df2, {16'd61407, 16'd47767, 16'd2165, 16'd35386, 16'd58120, 16'd46828, 16'd34456, 16'd11139, 16'd63600, 16'd44841, 16'd36660, 16'd17015, 16'd22721, 16'd52133, 16'd45693, 16'd16646, 16'd30407, 16'd58808, 16'd58147, 16'd607, 16'd4151, 16'd6042, 16'd47973, 16'd31235, 16'd14027, 16'd38841});
	test_expansion(128'h98b131fb99d0d4a7397d9f1dc7fca8b0, {16'd58153, 16'd49212, 16'd19236, 16'd61843, 16'd34072, 16'd157, 16'd50379, 16'd41942, 16'd65484, 16'd46693, 16'd38172, 16'd24403, 16'd5630, 16'd4906, 16'd39577, 16'd32549, 16'd61962, 16'd10579, 16'd64024, 16'd46762, 16'd23454, 16'd57130, 16'd25236, 16'd12225, 16'd54591, 16'd22715});
	test_expansion(128'hd42bf106ffcc3f0a9cb053d4bb5cada6, {16'd48450, 16'd19799, 16'd45640, 16'd42076, 16'd44747, 16'd7062, 16'd44463, 16'd65121, 16'd32294, 16'd47302, 16'd23686, 16'd45247, 16'd7399, 16'd44932, 16'd25957, 16'd44541, 16'd50818, 16'd24388, 16'd54195, 16'd53527, 16'd27864, 16'd12289, 16'd53655, 16'd52030, 16'd37477, 16'd15562});
	test_expansion(128'h727fff633f5a6a8d25b82fb9e3890496, {16'd32571, 16'd7372, 16'd15119, 16'd25977, 16'd26918, 16'd47939, 16'd7284, 16'd21957, 16'd59651, 16'd28994, 16'd54583, 16'd40544, 16'd31018, 16'd35736, 16'd55219, 16'd10507, 16'd30957, 16'd56158, 16'd16360, 16'd64777, 16'd50866, 16'd61780, 16'd748, 16'd64039, 16'd22931, 16'd18481});
	test_expansion(128'h5da1234a946c85f55fa247d95ca933a6, {16'd28686, 16'd14539, 16'd43654, 16'd21758, 16'd6982, 16'd33822, 16'd23587, 16'd47352, 16'd41859, 16'd26820, 16'd32584, 16'd18033, 16'd895, 16'd16124, 16'd13639, 16'd60713, 16'd63834, 16'd25143, 16'd33856, 16'd10977, 16'd64578, 16'd59606, 16'd29266, 16'd27978, 16'd53228, 16'd10258});
	test_expansion(128'hd49da8fcaa97ede440e2be7d3581b2ee, {16'd5260, 16'd12320, 16'd8742, 16'd60098, 16'd6938, 16'd26782, 16'd12017, 16'd21448, 16'd25143, 16'd7006, 16'd11336, 16'd38555, 16'd44343, 16'd13576, 16'd53761, 16'd13542, 16'd23569, 16'd6946, 16'd42561, 16'd52594, 16'd14313, 16'd51266, 16'd9790, 16'd14312, 16'd52535, 16'd63964});
	test_expansion(128'hebcfccaec5b484023496c5d5fb3b8e1a, {16'd3657, 16'd54152, 16'd49593, 16'd3393, 16'd39308, 16'd6350, 16'd40916, 16'd16819, 16'd16588, 16'd45709, 16'd44868, 16'd39708, 16'd38431, 16'd60162, 16'd47499, 16'd5174, 16'd34128, 16'd22867, 16'd50926, 16'd21354, 16'd40638, 16'd15031, 16'd60828, 16'd47201, 16'd27149, 16'd47758});
	test_expansion(128'hbfbd19cf8fee67e931aa77dc9f01ef35, {16'd43166, 16'd58432, 16'd52697, 16'd58111, 16'd38455, 16'd609, 16'd59454, 16'd41534, 16'd59953, 16'd296, 16'd29832, 16'd2977, 16'd20949, 16'd11252, 16'd1150, 16'd38037, 16'd62843, 16'd37399, 16'd46469, 16'd1192, 16'd29200, 16'd24299, 16'd20708, 16'd64171, 16'd12109, 16'd7541});
	test_expansion(128'h612b7fac1f698a5d3af887126f243e2a, {16'd34471, 16'd43330, 16'd40217, 16'd30197, 16'd2273, 16'd33435, 16'd25275, 16'd50295, 16'd42388, 16'd13449, 16'd63700, 16'd35602, 16'd2097, 16'd11604, 16'd4747, 16'd30787, 16'd64144, 16'd38178, 16'd49784, 16'd17445, 16'd21008, 16'd13872, 16'd19817, 16'd45265, 16'd33966, 16'd10620});
	test_expansion(128'hb912b17ce5d459cd671d35b455c86226, {16'd54122, 16'd20788, 16'd6205, 16'd39713, 16'd9989, 16'd42727, 16'd52890, 16'd14246, 16'd8828, 16'd52030, 16'd37536, 16'd18692, 16'd44707, 16'd17581, 16'd24217, 16'd32948, 16'd13290, 16'd40474, 16'd61713, 16'd62517, 16'd16437, 16'd11908, 16'd24572, 16'd11567, 16'd26507, 16'd23822});
	test_expansion(128'hc5ca3df0edf2f652f5eebb55c03ff34c, {16'd1829, 16'd3928, 16'd32476, 16'd10751, 16'd31566, 16'd44726, 16'd16796, 16'd39856, 16'd46349, 16'd20420, 16'd32627, 16'd35925, 16'd16896, 16'd16307, 16'd34558, 16'd58658, 16'd6012, 16'd28293, 16'd38983, 16'd40248, 16'd14857, 16'd60164, 16'd3925, 16'd49649, 16'd58949, 16'd2536});
	test_expansion(128'hf0151b125719412f5977b31cf145d026, {16'd13687, 16'd63993, 16'd37899, 16'd1591, 16'd7280, 16'd39100, 16'd47429, 16'd41986, 16'd22119, 16'd55359, 16'd62511, 16'd6823, 16'd35899, 16'd32440, 16'd54627, 16'd34077, 16'd1795, 16'd34244, 16'd4122, 16'd9517, 16'd52981, 16'd27906, 16'd32596, 16'd15672, 16'd52958, 16'd12390});
	test_expansion(128'h1f77aee62d46f71eb2c2a4ebf858e5ef, {16'd45043, 16'd10747, 16'd9850, 16'd39439, 16'd40981, 16'd16322, 16'd56048, 16'd59939, 16'd61629, 16'd49702, 16'd43434, 16'd20268, 16'd48232, 16'd28607, 16'd59323, 16'd27719, 16'd14313, 16'd36061, 16'd28875, 16'd48539, 16'd47353, 16'd20612, 16'd42675, 16'd19329, 16'd10577, 16'd57735});
	test_expansion(128'h1eeaf697bde6be9d6c76d46135f492da, {16'd26096, 16'd5357, 16'd56778, 16'd42904, 16'd3641, 16'd36424, 16'd15254, 16'd44161, 16'd36436, 16'd50658, 16'd43573, 16'd32901, 16'd18178, 16'd8413, 16'd30433, 16'd33415, 16'd26052, 16'd11149, 16'd6982, 16'd10991, 16'd15480, 16'd21304, 16'd42590, 16'd7155, 16'd44690, 16'd24188});
	test_expansion(128'h3e5f70d1060b2a78a1b59cdec9b8e4b3, {16'd23870, 16'd37821, 16'd61137, 16'd64557, 16'd34986, 16'd49434, 16'd14355, 16'd607, 16'd35634, 16'd62262, 16'd38522, 16'd41499, 16'd51682, 16'd26824, 16'd4380, 16'd22703, 16'd290, 16'd27197, 16'd21171, 16'd17448, 16'd38504, 16'd58589, 16'd19418, 16'd36261, 16'd20236, 16'd8975});
	test_expansion(128'h1a66c22e42653622001a6eecb2fcc082, {16'd55383, 16'd62132, 16'd25607, 16'd16359, 16'd18714, 16'd43935, 16'd40041, 16'd24014, 16'd39846, 16'd50172, 16'd42640, 16'd56544, 16'd23248, 16'd41387, 16'd19806, 16'd45103, 16'd59464, 16'd28945, 16'd13281, 16'd1519, 16'd35503, 16'd61953, 16'd8340, 16'd47382, 16'd48710, 16'd40530});
	test_expansion(128'h31612c63e03cdbe51b7da5dcdafc1820, {16'd44430, 16'd25089, 16'd24601, 16'd53783, 16'd41775, 16'd193, 16'd50635, 16'd11316, 16'd42846, 16'd5657, 16'd60259, 16'd53716, 16'd3877, 16'd29374, 16'd27816, 16'd2590, 16'd64103, 16'd28585, 16'd28284, 16'd33946, 16'd41695, 16'd32728, 16'd54871, 16'd34923, 16'd36339, 16'd52351});
	test_expansion(128'hebd8aaca934b4604efeed7ab47d6f28a, {16'd38224, 16'd663, 16'd35703, 16'd5302, 16'd51876, 16'd36365, 16'd33966, 16'd38384, 16'd37639, 16'd3776, 16'd30321, 16'd21078, 16'd35776, 16'd61097, 16'd1841, 16'd60075, 16'd13170, 16'd63360, 16'd25414, 16'd17340, 16'd36943, 16'd24589, 16'd53743, 16'd61617, 16'd18813, 16'd10722});
	test_expansion(128'h1f1306407aacb053ac5d2e5ab15d653b, {16'd9445, 16'd60792, 16'd32189, 16'd47011, 16'd6097, 16'd64716, 16'd37689, 16'd7001, 16'd49518, 16'd50334, 16'd16150, 16'd21420, 16'd29371, 16'd65234, 16'd15380, 16'd12062, 16'd26604, 16'd15955, 16'd36947, 16'd44586, 16'd38560, 16'd6106, 16'd31471, 16'd516, 16'd32323, 16'd33323});
	test_expansion(128'hd6afa847152f8b6db25b0c4d821dcb40, {16'd20577, 16'd780, 16'd10274, 16'd33955, 16'd30741, 16'd61296, 16'd52620, 16'd9619, 16'd31275, 16'd53274, 16'd23709, 16'd18323, 16'd65053, 16'd53581, 16'd35107, 16'd14371, 16'd8247, 16'd16198, 16'd17917, 16'd47975, 16'd58507, 16'd21953, 16'd61309, 16'd48617, 16'd36339, 16'd31631});
	test_expansion(128'hbc5447efa6e8b688b4f625ede63b4312, {16'd57752, 16'd49887, 16'd17789, 16'd19668, 16'd6334, 16'd34266, 16'd1160, 16'd6306, 16'd39194, 16'd33237, 16'd47518, 16'd43691, 16'd5648, 16'd6412, 16'd35533, 16'd29821, 16'd15681, 16'd30383, 16'd53120, 16'd41250, 16'd48900, 16'd1389, 16'd12205, 16'd41596, 16'd54723, 16'd38501});
	test_expansion(128'h2704612e9b716abb45e679bfa2bb39c9, {16'd4580, 16'd62308, 16'd15959, 16'd18383, 16'd50818, 16'd61874, 16'd57639, 16'd18760, 16'd57259, 16'd32793, 16'd9885, 16'd57253, 16'd59587, 16'd35756, 16'd5325, 16'd12584, 16'd60256, 16'd8598, 16'd42344, 16'd19521, 16'd46849, 16'd24008, 16'd31489, 16'd63713, 16'd22185, 16'd41542});
	test_expansion(128'hf195091268a6dfb9f07c902213b5198c, {16'd22344, 16'd47869, 16'd59593, 16'd31566, 16'd15742, 16'd45090, 16'd40576, 16'd54859, 16'd58840, 16'd38674, 16'd29220, 16'd13606, 16'd22757, 16'd21462, 16'd40746, 16'd26179, 16'd9880, 16'd59768, 16'd27077, 16'd44709, 16'd44272, 16'd36949, 16'd26634, 16'd18842, 16'd51838, 16'd56014});
	test_expansion(128'h5e2e4f9d5ac993571b15fdd28a55dd8b, {16'd56367, 16'd14390, 16'd59308, 16'd57073, 16'd23102, 16'd13813, 16'd37141, 16'd55773, 16'd6788, 16'd34554, 16'd54264, 16'd20560, 16'd30388, 16'd62802, 16'd24589, 16'd13632, 16'd54897, 16'd4021, 16'd2094, 16'd39541, 16'd64320, 16'd49479, 16'd32390, 16'd17241, 16'd4980, 16'd46964});
	test_expansion(128'h2ba0872512939e936a3c158def5e2163, {16'd21740, 16'd25950, 16'd35542, 16'd37622, 16'd59270, 16'd62014, 16'd12516, 16'd37505, 16'd6058, 16'd9951, 16'd22265, 16'd24249, 16'd55782, 16'd41924, 16'd17758, 16'd8458, 16'd10323, 16'd30806, 16'd11461, 16'd48625, 16'd7705, 16'd63137, 16'd45226, 16'd54048, 16'd40701, 16'd20455});
	test_expansion(128'hadf6b0191111efb22363775ea3653ee4, {16'd11007, 16'd44711, 16'd2633, 16'd30061, 16'd53215, 16'd16164, 16'd40123, 16'd59966, 16'd58367, 16'd25599, 16'd15130, 16'd36484, 16'd39484, 16'd7769, 16'd20876, 16'd65069, 16'd28173, 16'd29296, 16'd64214, 16'd30898, 16'd26471, 16'd14497, 16'd36445, 16'd50603, 16'd24056, 16'd51133});
	test_expansion(128'h3737bc097d79aee82465f2d6bb45eae8, {16'd64519, 16'd49543, 16'd63021, 16'd33400, 16'd45223, 16'd23052, 16'd17901, 16'd15447, 16'd17458, 16'd22359, 16'd43320, 16'd60980, 16'd13162, 16'd21712, 16'd33474, 16'd13898, 16'd33004, 16'd37991, 16'd51036, 16'd40219, 16'd56888, 16'd12995, 16'd5700, 16'd60465, 16'd37094, 16'd5862});
	test_expansion(128'h40028ae3a81b2637da0083f115bc8626, {16'd8819, 16'd19874, 16'd16078, 16'd10184, 16'd8400, 16'd38121, 16'd6455, 16'd59377, 16'd39618, 16'd36474, 16'd52639, 16'd53071, 16'd24070, 16'd37615, 16'd42546, 16'd57486, 16'd48561, 16'd29210, 16'd3404, 16'd26280, 16'd41782, 16'd41512, 16'd65384, 16'd24555, 16'd245, 16'd13262});
	test_expansion(128'hc53b779d440871efb1d723f934820e76, {16'd2072, 16'd17202, 16'd53738, 16'd29694, 16'd25727, 16'd60840, 16'd65373, 16'd5072, 16'd2499, 16'd11641, 16'd24218, 16'd14121, 16'd21717, 16'd52790, 16'd24979, 16'd47681, 16'd47756, 16'd47823, 16'd45518, 16'd45281, 16'd41750, 16'd63647, 16'd5754, 16'd2039, 16'd51467, 16'd44665});
	test_expansion(128'ha03372f4f3496ade1ccb7e4fbd6af890, {16'd8523, 16'd26220, 16'd60324, 16'd22849, 16'd36440, 16'd47252, 16'd19927, 16'd14450, 16'd54423, 16'd38566, 16'd9772, 16'd50788, 16'd13030, 16'd63889, 16'd32786, 16'd4634, 16'd41688, 16'd38601, 16'd20060, 16'd27238, 16'd10961, 16'd48367, 16'd11014, 16'd49180, 16'd46965, 16'd28190});
	test_expansion(128'h56b2cb6929a21e48cd63780bf85d4f14, {16'd8410, 16'd10436, 16'd64895, 16'd16543, 16'd3987, 16'd12473, 16'd29459, 16'd18015, 16'd42667, 16'd65162, 16'd34523, 16'd31411, 16'd53291, 16'd27480, 16'd22804, 16'd13197, 16'd28380, 16'd2800, 16'd45140, 16'd58043, 16'd60610, 16'd43528, 16'd1198, 16'd29015, 16'd42927, 16'd49812});
	test_expansion(128'h4851d5280bf3494c8918ae07dec8a17a, {16'd37866, 16'd48122, 16'd50563, 16'd42963, 16'd24497, 16'd49952, 16'd17744, 16'd25541, 16'd8606, 16'd9512, 16'd8959, 16'd42330, 16'd50463, 16'd8912, 16'd2861, 16'd55983, 16'd32390, 16'd56344, 16'd16479, 16'd9627, 16'd2931, 16'd49976, 16'd58517, 16'd36708, 16'd13820, 16'd34095});
	test_expansion(128'h96810a3af80c48737e604bc72d4c04ae, {16'd56028, 16'd40218, 16'd41700, 16'd60612, 16'd23724, 16'd28718, 16'd52238, 16'd61810, 16'd24980, 16'd34356, 16'd50720, 16'd4410, 16'd37029, 16'd7476, 16'd15032, 16'd20372, 16'd44224, 16'd35185, 16'd5010, 16'd33890, 16'd46393, 16'd51701, 16'd32968, 16'd33347, 16'd15527, 16'd27944});
	test_expansion(128'h5c09fd7cec6b1e554009ec3eca99fbd2, {16'd22561, 16'd1725, 16'd5360, 16'd30501, 16'd40063, 16'd15317, 16'd4440, 16'd5661, 16'd63484, 16'd56396, 16'd22361, 16'd47954, 16'd49649, 16'd15377, 16'd57043, 16'd5163, 16'd37224, 16'd15936, 16'd26721, 16'd20900, 16'd41155, 16'd13569, 16'd57806, 16'd20540, 16'd65522, 16'd31714});
	test_expansion(128'hdd0926bde5f4939760105f148c2222ee, {16'd13037, 16'd4174, 16'd7841, 16'd19282, 16'd58746, 16'd64091, 16'd43181, 16'd9472, 16'd59459, 16'd2854, 16'd63822, 16'd22482, 16'd26457, 16'd39594, 16'd26159, 16'd45718, 16'd26171, 16'd39268, 16'd11253, 16'd48382, 16'd13323, 16'd53486, 16'd39095, 16'd14441, 16'd32569, 16'd34289});
	test_expansion(128'h974a80eb320041dfebe1dd6ac2bcf0a4, {16'd39032, 16'd10883, 16'd28427, 16'd5906, 16'd55445, 16'd23244, 16'd40616, 16'd15066, 16'd8239, 16'd46619, 16'd25849, 16'd28314, 16'd2329, 16'd64696, 16'd31643, 16'd8907, 16'd18848, 16'd41182, 16'd14723, 16'd7766, 16'd50276, 16'd36738, 16'd6786, 16'd17161, 16'd34095, 16'd495});
	test_expansion(128'h860dc1d80b2f146bcbeb5dde125c22bf, {16'd41346, 16'd43091, 16'd36639, 16'd51663, 16'd57684, 16'd52358, 16'd23497, 16'd6228, 16'd49685, 16'd35112, 16'd23397, 16'd26288, 16'd785, 16'd62398, 16'd18134, 16'd2480, 16'd7401, 16'd59812, 16'd20764, 16'd64708, 16'd5679, 16'd14287, 16'd62456, 16'd5009, 16'd24078, 16'd42623});
	test_expansion(128'h0a034c729905109154c63591a791b23c, {16'd32227, 16'd44105, 16'd18515, 16'd50032, 16'd53471, 16'd46176, 16'd45248, 16'd41301, 16'd42595, 16'd64571, 16'd63877, 16'd33378, 16'd10544, 16'd15693, 16'd38891, 16'd64063, 16'd62890, 16'd34375, 16'd61186, 16'd59901, 16'd27102, 16'd5245, 16'd29493, 16'd44470, 16'd15037, 16'd8846});
	test_expansion(128'h21606679c2f390fa618d0a54686fa5ba, {16'd27685, 16'd17734, 16'd44249, 16'd16482, 16'd58123, 16'd64436, 16'd60498, 16'd44934, 16'd50374, 16'd58398, 16'd33452, 16'd36628, 16'd8388, 16'd9824, 16'd48789, 16'd605, 16'd48786, 16'd52422, 16'd28723, 16'd16563, 16'd29042, 16'd8940, 16'd60986, 16'd58767, 16'd64958, 16'd15253});
	test_expansion(128'h36c5e7cacb695263982c7f4897af7bae, {16'd33517, 16'd51194, 16'd18709, 16'd15779, 16'd23896, 16'd48120, 16'd55409, 16'd45239, 16'd57819, 16'd55695, 16'd28813, 16'd49280, 16'd5267, 16'd16439, 16'd2674, 16'd18141, 16'd35696, 16'd6689, 16'd14628, 16'd64742, 16'd6660, 16'd62266, 16'd24619, 16'd47523, 16'd19729, 16'd61556});
	test_expansion(128'h408e43aec598d2bf2b1033cfd45743ad, {16'd30175, 16'd18347, 16'd29457, 16'd50888, 16'd59900, 16'd46264, 16'd41587, 16'd21247, 16'd51539, 16'd2885, 16'd31401, 16'd15253, 16'd50457, 16'd58006, 16'd30130, 16'd41183, 16'd56010, 16'd55170, 16'd7687, 16'd12010, 16'd30913, 16'd4615, 16'd35068, 16'd55680, 16'd27328, 16'd19099});
	test_expansion(128'h2b6347246a19d758df868a5f93520df9, {16'd50057, 16'd2327, 16'd36053, 16'd1403, 16'd58708, 16'd4909, 16'd44333, 16'd53650, 16'd40789, 16'd979, 16'd44219, 16'd49119, 16'd25182, 16'd51975, 16'd36045, 16'd3332, 16'd33920, 16'd22894, 16'd35186, 16'd19855, 16'd30922, 16'd10628, 16'd30262, 16'd7500, 16'd59524, 16'd17273});
	test_expansion(128'h0b23adf400dcad51e5174f6790461505, {16'd33331, 16'd61192, 16'd61154, 16'd38050, 16'd54771, 16'd57099, 16'd51609, 16'd27564, 16'd54675, 16'd13484, 16'd1720, 16'd22662, 16'd45552, 16'd49155, 16'd2800, 16'd43152, 16'd39231, 16'd40982, 16'd25962, 16'd2941, 16'd24287, 16'd13409, 16'd1903, 16'd20141, 16'd33327, 16'd25212});
	test_expansion(128'h24705c1de61a4c3dad5529c2ed25358c, {16'd5670, 16'd9639, 16'd31888, 16'd17544, 16'd8916, 16'd22168, 16'd64546, 16'd9060, 16'd64141, 16'd12808, 16'd23371, 16'd523, 16'd25133, 16'd18933, 16'd51660, 16'd15693, 16'd12972, 16'd40067, 16'd61668, 16'd62603, 16'd19508, 16'd54134, 16'd26376, 16'd37259, 16'd30535, 16'd28920});
	test_expansion(128'hf01d2f9c015917e48dd21282d59123d0, {16'd10261, 16'd43627, 16'd32024, 16'd26055, 16'd14236, 16'd28395, 16'd47705, 16'd39747, 16'd10563, 16'd23062, 16'd6445, 16'd57362, 16'd18601, 16'd31747, 16'd1211, 16'd32986, 16'd20699, 16'd9363, 16'd10012, 16'd52444, 16'd3185, 16'd52652, 16'd36642, 16'd8838, 16'd34836, 16'd59304});
	test_expansion(128'ha3873e9d0acb11bcbaab82fcc212dd8e, {16'd56007, 16'd62779, 16'd10403, 16'd29930, 16'd57453, 16'd23643, 16'd12529, 16'd6611, 16'd24637, 16'd6321, 16'd18327, 16'd58622, 16'd42884, 16'd9630, 16'd13467, 16'd36291, 16'd28322, 16'd27130, 16'd46237, 16'd32615, 16'd25567, 16'd60209, 16'd54910, 16'd44290, 16'd42744, 16'd22634});
	test_expansion(128'h7d798b6fb2a24be7314bfc43204b2e9f, {16'd8548, 16'd47376, 16'd19994, 16'd4686, 16'd36252, 16'd21236, 16'd54935, 16'd38461, 16'd65285, 16'd16581, 16'd53413, 16'd7109, 16'd24025, 16'd5171, 16'd30675, 16'd40413, 16'd15636, 16'd9398, 16'd10890, 16'd14610, 16'd36614, 16'd36631, 16'd26367, 16'd24187, 16'd36537, 16'd11658});
	test_expansion(128'h08e30f709b2afedf018cb7e479492f55, {16'd54217, 16'd50041, 16'd55435, 16'd29198, 16'd54010, 16'd46322, 16'd30180, 16'd390, 16'd40565, 16'd64365, 16'd245, 16'd2220, 16'd60165, 16'd48368, 16'd13061, 16'd7146, 16'd4252, 16'd48613, 16'd39880, 16'd59025, 16'd30526, 16'd52728, 16'd57617, 16'd55775, 16'd20436, 16'd40826});
	test_expansion(128'h43059992e1e488e5727f836e60369201, {16'd21862, 16'd3517, 16'd14549, 16'd43164, 16'd39377, 16'd20982, 16'd62373, 16'd7343, 16'd14580, 16'd46482, 16'd32644, 16'd238, 16'd6994, 16'd27484, 16'd35307, 16'd5412, 16'd42713, 16'd47470, 16'd46341, 16'd42264, 16'd26409, 16'd7057, 16'd6739, 16'd11601, 16'd41256, 16'd27037});
	test_expansion(128'h0e252231c2f54e51052c46c767b6792a, {16'd48953, 16'd20683, 16'd40815, 16'd46490, 16'd39788, 16'd51980, 16'd65177, 16'd60191, 16'd9383, 16'd29774, 16'd16048, 16'd27561, 16'd55900, 16'd62387, 16'd62202, 16'd19040, 16'd61135, 16'd23243, 16'd55109, 16'd32409, 16'd40121, 16'd9942, 16'd13942, 16'd19201, 16'd12682, 16'd58360});
	test_expansion(128'h7d2f6b13bc69b1cc87fb4315835c06fa, {16'd45135, 16'd24880, 16'd9585, 16'd51393, 16'd33214, 16'd45008, 16'd41316, 16'd15045, 16'd25605, 16'd4442, 16'd28899, 16'd48165, 16'd40000, 16'd1043, 16'd6391, 16'd9686, 16'd5216, 16'd52810, 16'd62176, 16'd35192, 16'd60112, 16'd45946, 16'd55449, 16'd23267, 16'd61191, 16'd38072});
	test_expansion(128'h5c7fa7561156346a8d7a44d541e19854, {16'd31716, 16'd23031, 16'd55043, 16'd37128, 16'd30126, 16'd60034, 16'd41393, 16'd18794, 16'd55054, 16'd29084, 16'd62591, 16'd37625, 16'd49102, 16'd39847, 16'd25632, 16'd52580, 16'd31259, 16'd52914, 16'd36974, 16'd37686, 16'd19563, 16'd26771, 16'd25660, 16'd5335, 16'd50473, 16'd54808});
	test_expansion(128'h5c1ee8881743c12b23946a7425fd9cd0, {16'd34629, 16'd62294, 16'd35180, 16'd34510, 16'd6829, 16'd5445, 16'd62978, 16'd36145, 16'd37024, 16'd22348, 16'd29618, 16'd60024, 16'd25728, 16'd31710, 16'd31163, 16'd46424, 16'd6169, 16'd37256, 16'd56184, 16'd6557, 16'd20832, 16'd25772, 16'd52266, 16'd6727, 16'd8695, 16'd36611});
	test_expansion(128'h8409cd7a7b4a7ff4d04dac93d5b92665, {16'd55864, 16'd41052, 16'd18146, 16'd62753, 16'd60616, 16'd15135, 16'd34250, 16'd7870, 16'd9853, 16'd38115, 16'd27040, 16'd11574, 16'd30226, 16'd52102, 16'd33414, 16'd20144, 16'd17237, 16'd10560, 16'd3653, 16'd54158, 16'd21675, 16'd28480, 16'd29455, 16'd6299, 16'd9850, 16'd7610});
	test_expansion(128'h6035eed76eda8ba24c022aa9d944bfda, {16'd60733, 16'd52065, 16'd25723, 16'd51015, 16'd45063, 16'd2310, 16'd36815, 16'd39496, 16'd9594, 16'd53271, 16'd28968, 16'd62804, 16'd50827, 16'd59034, 16'd33964, 16'd43579, 16'd56620, 16'd3797, 16'd40057, 16'd19214, 16'd6782, 16'd7102, 16'd30557, 16'd14073, 16'd5775, 16'd57812});
	test_expansion(128'hbfb6c4e4902817c98d85e23f44a56988, {16'd55202, 16'd22546, 16'd32266, 16'd60942, 16'd18774, 16'd12946, 16'd13539, 16'd28334, 16'd31941, 16'd3267, 16'd59474, 16'd64252, 16'd40279, 16'd60700, 16'd2030, 16'd6261, 16'd39227, 16'd17919, 16'd8076, 16'd41670, 16'd20242, 16'd46403, 16'd38957, 16'd19668, 16'd39898, 16'd29044});
	test_expansion(128'h556302df145e100c62780bb782ec54a3, {16'd38923, 16'd4597, 16'd50998, 16'd25384, 16'd33427, 16'd3753, 16'd59569, 16'd31431, 16'd11177, 16'd2445, 16'd19857, 16'd25438, 16'd19531, 16'd16647, 16'd51672, 16'd21323, 16'd57307, 16'd41501, 16'd52652, 16'd5368, 16'd40990, 16'd40377, 16'd49908, 16'd28219, 16'd24379, 16'd9337});
	test_expansion(128'ha4ea4f1796644822bc2bc758994efaaf, {16'd65177, 16'd63743, 16'd38714, 16'd9584, 16'd54548, 16'd30018, 16'd50706, 16'd6891, 16'd24394, 16'd1656, 16'd13781, 16'd20645, 16'd44401, 16'd10421, 16'd17042, 16'd4199, 16'd43937, 16'd6081, 16'd57068, 16'd19107, 16'd27344, 16'd62943, 16'd60292, 16'd33105, 16'd22820, 16'd44250});
	test_expansion(128'h33ec797abde98231f7454432d3b3d741, {16'd31646, 16'd4496, 16'd27102, 16'd22621, 16'd64877, 16'd3778, 16'd22818, 16'd41575, 16'd5936, 16'd50149, 16'd383, 16'd56803, 16'd12129, 16'd18357, 16'd47772, 16'd55877, 16'd54575, 16'd17424, 16'd11632, 16'd46921, 16'd42412, 16'd27424, 16'd2545, 16'd23338, 16'd57784, 16'd39880});
	test_expansion(128'h46b46f2f889e83284a2b07da6898561a, {16'd21471, 16'd54058, 16'd39091, 16'd15588, 16'd60285, 16'd56650, 16'd57271, 16'd27689, 16'd4176, 16'd11416, 16'd48884, 16'd57038, 16'd6171, 16'd37718, 16'd43668, 16'd50877, 16'd43505, 16'd32266, 16'd40909, 16'd52264, 16'd1914, 16'd14818, 16'd511, 16'd1726, 16'd28036, 16'd47993});
	test_expansion(128'h76607a9bcb872539075cc88cb10e5264, {16'd52881, 16'd25787, 16'd13751, 16'd1482, 16'd33780, 16'd21447, 16'd44014, 16'd59813, 16'd44410, 16'd41791, 16'd6775, 16'd12265, 16'd43534, 16'd40612, 16'd64027, 16'd1124, 16'd49593, 16'd18358, 16'd21126, 16'd17820, 16'd49361, 16'd56233, 16'd22706, 16'd41239, 16'd35062, 16'd50179});
	test_expansion(128'h3869697f37a0cf4f4514ed5b2ef2f05e, {16'd63858, 16'd19523, 16'd6812, 16'd43255, 16'd8977, 16'd31504, 16'd16101, 16'd39114, 16'd21263, 16'd14654, 16'd24483, 16'd60656, 16'd41178, 16'd55816, 16'd14385, 16'd4379, 16'd49637, 16'd36677, 16'd47729, 16'd60433, 16'd2667, 16'd46271, 16'd30514, 16'd5142, 16'd51240, 16'd11339});
	test_expansion(128'hd5d60d7356e7618915e3c0237a922e5c, {16'd27945, 16'd61481, 16'd5218, 16'd33867, 16'd14752, 16'd25525, 16'd41923, 16'd55509, 16'd36460, 16'd46532, 16'd31350, 16'd40140, 16'd62938, 16'd27335, 16'd8204, 16'd33272, 16'd42950, 16'd53186, 16'd56406, 16'd48560, 16'd39287, 16'd13359, 16'd52054, 16'd12142, 16'd14555, 16'd26834});
	test_expansion(128'hc49a44928595e1d10e3e184cfb6ec83d, {16'd36894, 16'd36969, 16'd8286, 16'd47786, 16'd18819, 16'd29268, 16'd62204, 16'd3542, 16'd51148, 16'd58607, 16'd37917, 16'd9789, 16'd22456, 16'd60439, 16'd14925, 16'd22696, 16'd6750, 16'd11807, 16'd34704, 16'd51636, 16'd28825, 16'd25605, 16'd21195, 16'd48752, 16'd51760, 16'd47628});
	test_expansion(128'h025695e818668c873e45db8ba70f26d1, {16'd40153, 16'd8306, 16'd27484, 16'd40819, 16'd54001, 16'd45049, 16'd55341, 16'd29173, 16'd37829, 16'd22943, 16'd19293, 16'd9178, 16'd1587, 16'd53333, 16'd1764, 16'd59691, 16'd8025, 16'd45867, 16'd53628, 16'd43888, 16'd43447, 16'd42246, 16'd26267, 16'd9497, 16'd52452, 16'd42637});
	test_expansion(128'hd33f631c4ea220dd3183f20f263b666c, {16'd44510, 16'd5703, 16'd57955, 16'd2252, 16'd45914, 16'd7712, 16'd8020, 16'd54535, 16'd34552, 16'd40380, 16'd42057, 16'd29181, 16'd46847, 16'd17621, 16'd46402, 16'd17091, 16'd25145, 16'd2806, 16'd1906, 16'd52410, 16'd33664, 16'd28878, 16'd55144, 16'd57018, 16'd59283, 16'd2095});
	test_expansion(128'hde3daa62b53af3597ea4027cf5b5a1da, {16'd34378, 16'd30374, 16'd30610, 16'd23611, 16'd31898, 16'd48472, 16'd6063, 16'd33935, 16'd57167, 16'd45033, 16'd11497, 16'd13613, 16'd48295, 16'd16548, 16'd60550, 16'd27596, 16'd49134, 16'd14279, 16'd5904, 16'd55168, 16'd43800, 16'd63786, 16'd9559, 16'd20156, 16'd41298, 16'd61203});
	test_expansion(128'h4754037889d03dc0915efbb66e8976bc, {16'd39809, 16'd9530, 16'd44729, 16'd21201, 16'd64188, 16'd41564, 16'd18324, 16'd8177, 16'd17172, 16'd41906, 16'd28059, 16'd7402, 16'd32491, 16'd20876, 16'd19437, 16'd51178, 16'd19124, 16'd20164, 16'd3194, 16'd27280, 16'd63059, 16'd16634, 16'd59626, 16'd8818, 16'd51639, 16'd49775});
	test_expansion(128'h331aaaa3ef2bb04447b28c41836e9029, {16'd31077, 16'd33791, 16'd5763, 16'd8035, 16'd58058, 16'd936, 16'd34219, 16'd27554, 16'd49578, 16'd55207, 16'd25664, 16'd23621, 16'd6753, 16'd48862, 16'd3973, 16'd9214, 16'd53660, 16'd44232, 16'd51529, 16'd27795, 16'd35950, 16'd4233, 16'd17035, 16'd46722, 16'd50774, 16'd44914});
	test_expansion(128'hb327d056bfba1be70d10e8109c7c7980, {16'd25535, 16'd32857, 16'd38106, 16'd17901, 16'd11750, 16'd8818, 16'd23718, 16'd45439, 16'd9770, 16'd57172, 16'd61347, 16'd48825, 16'd25133, 16'd1390, 16'd64920, 16'd53959, 16'd37958, 16'd48421, 16'd9832, 16'd15885, 16'd50165, 16'd47120, 16'd23174, 16'd14264, 16'd17484, 16'd25837});
	test_expansion(128'hadcfb80d7e1dd66184efbfea4416949c, {16'd44962, 16'd4491, 16'd54084, 16'd61740, 16'd1036, 16'd8868, 16'd36520, 16'd24881, 16'd50443, 16'd16572, 16'd60597, 16'd63041, 16'd27034, 16'd40745, 16'd60615, 16'd33041, 16'd63605, 16'd36272, 16'd24114, 16'd19670, 16'd19599, 16'd41198, 16'd53539, 16'd22864, 16'd7363, 16'd7171});
	test_expansion(128'h446e694ad9880b8c01ee9166c935f9e8, {16'd56096, 16'd21583, 16'd6049, 16'd48090, 16'd11165, 16'd62234, 16'd37158, 16'd20496, 16'd26944, 16'd29671, 16'd8473, 16'd59212, 16'd16388, 16'd54350, 16'd45762, 16'd53883, 16'd43719, 16'd60967, 16'd37103, 16'd11363, 16'd27187, 16'd61932, 16'd35720, 16'd1620, 16'd28900, 16'd7052});
	test_expansion(128'ha52cc7cf42ed2646ccb508e259076021, {16'd6855, 16'd5315, 16'd20521, 16'd28978, 16'd38242, 16'd36025, 16'd24163, 16'd63368, 16'd32431, 16'd2482, 16'd8372, 16'd7216, 16'd11348, 16'd46566, 16'd23775, 16'd32343, 16'd47449, 16'd33296, 16'd17369, 16'd4086, 16'd32630, 16'd39357, 16'd40928, 16'd32877, 16'd27086, 16'd65026});
	test_expansion(128'he359fefaa5895325583ba6bc9da097b0, {16'd34886, 16'd60624, 16'd31777, 16'd15500, 16'd63207, 16'd8452, 16'd23088, 16'd46496, 16'd47771, 16'd50338, 16'd44278, 16'd1487, 16'd15642, 16'd6891, 16'd64229, 16'd15766, 16'd56404, 16'd45400, 16'd45989, 16'd1865, 16'd11736, 16'd13678, 16'd8542, 16'd62108, 16'd20379, 16'd28161});
	test_expansion(128'h372be1379a86ccabae7b6964ba9b7ad4, {16'd673, 16'd52079, 16'd61746, 16'd28896, 16'd32379, 16'd42312, 16'd45969, 16'd8906, 16'd3050, 16'd54134, 16'd44821, 16'd63356, 16'd64825, 16'd9814, 16'd17362, 16'd12491, 16'd34809, 16'd1590, 16'd821, 16'd5233, 16'd47138, 16'd6821, 16'd13297, 16'd48331, 16'd44690, 16'd7023});
	test_expansion(128'h21a2848bc0ab5bb362e5de6e1d02e968, {16'd17051, 16'd54659, 16'd63216, 16'd38117, 16'd11741, 16'd49143, 16'd65279, 16'd45849, 16'd2505, 16'd34253, 16'd13521, 16'd32613, 16'd39194, 16'd27158, 16'd13457, 16'd19090, 16'd14420, 16'd53143, 16'd24140, 16'd14120, 16'd22121, 16'd36714, 16'd50318, 16'd57903, 16'd10140, 16'd53373});
	test_expansion(128'h7b0195302cb00863b02e34ac99490d06, {16'd8708, 16'd54440, 16'd29520, 16'd59324, 16'd40563, 16'd29836, 16'd38398, 16'd57878, 16'd39066, 16'd58419, 16'd14535, 16'd13119, 16'd7978, 16'd42765, 16'd9541, 16'd32197, 16'd19029, 16'd40590, 16'd53004, 16'd34318, 16'd43239, 16'd21139, 16'd42095, 16'd8807, 16'd18389, 16'd39551});
	test_expansion(128'h9377db74029369f9982386f302e7b81f, {16'd5936, 16'd28117, 16'd57276, 16'd11618, 16'd14930, 16'd33360, 16'd24532, 16'd11045, 16'd42979, 16'd407, 16'd7078, 16'd30798, 16'd22292, 16'd50596, 16'd10579, 16'd39055, 16'd33150, 16'd60361, 16'd10001, 16'd6270, 16'd20442, 16'd39331, 16'd55255, 16'd48000, 16'd62198, 16'd22686});
	test_expansion(128'h9498a013f1bacc10d8fd8ff445273635, {16'd33586, 16'd4289, 16'd30113, 16'd36052, 16'd10811, 16'd27089, 16'd46129, 16'd7815, 16'd12645, 16'd5528, 16'd19235, 16'd4553, 16'd56496, 16'd16278, 16'd28463, 16'd36813, 16'd22634, 16'd34556, 16'd43441, 16'd53017, 16'd31951, 16'd34940, 16'd53819, 16'd8575, 16'd31942, 16'd2923});
	test_expansion(128'h045a17ca28e027e08efdd3b5dcf323d4, {16'd60104, 16'd3895, 16'd60481, 16'd26936, 16'd5354, 16'd20654, 16'd30000, 16'd41777, 16'd64119, 16'd39492, 16'd31285, 16'd37197, 16'd34307, 16'd5431, 16'd5742, 16'd11340, 16'd25688, 16'd57844, 16'd60351, 16'd63670, 16'd18719, 16'd54206, 16'd11123, 16'd12767, 16'd57772, 16'd46999});
	test_expansion(128'h0c8f8b5ef16e87cfa7a70ed7a576baad, {16'd35833, 16'd50303, 16'd16364, 16'd23612, 16'd45453, 16'd28086, 16'd16844, 16'd64047, 16'd46739, 16'd25649, 16'd62037, 16'd24790, 16'd10093, 16'd24339, 16'd18229, 16'd34224, 16'd26737, 16'd62143, 16'd63706, 16'd34805, 16'd39762, 16'd17367, 16'd28891, 16'd23879, 16'd47346, 16'd19558});
	test_expansion(128'hd95a9ac239e26ee5515931f31986aeb3, {16'd31856, 16'd24836, 16'd39583, 16'd72, 16'd40140, 16'd14493, 16'd44182, 16'd17699, 16'd10953, 16'd10001, 16'd43817, 16'd29065, 16'd29429, 16'd56456, 16'd38052, 16'd43010, 16'd60377, 16'd47152, 16'd12092, 16'd41929, 16'd11337, 16'd7899, 16'd16970, 16'd31163, 16'd48603, 16'd56314});
	test_expansion(128'he771b90c5ee9f6016127312675893dcc, {16'd19604, 16'd9835, 16'd32309, 16'd48065, 16'd58440, 16'd5216, 16'd38940, 16'd28112, 16'd3261, 16'd41669, 16'd34281, 16'd62953, 16'd42510, 16'd58571, 16'd57812, 16'd47763, 16'd50077, 16'd11092, 16'd40062, 16'd32763, 16'd29729, 16'd38266, 16'd56708, 16'd37601, 16'd9484, 16'd38864});
	test_expansion(128'h4a56377d903ebd3b1f2187db2690e03c, {16'd54801, 16'd13380, 16'd56789, 16'd56827, 16'd7031, 16'd19059, 16'd54619, 16'd6665, 16'd26178, 16'd5677, 16'd6751, 16'd25790, 16'd10041, 16'd5850, 16'd10411, 16'd33389, 16'd29862, 16'd2776, 16'd55143, 16'd50390, 16'd43118, 16'd26297, 16'd38150, 16'd9461, 16'd42532, 16'd35179});
	test_expansion(128'h41d0d5f0bdd64bccc96a0663f4c9d584, {16'd11725, 16'd21894, 16'd14803, 16'd17185, 16'd45421, 16'd17896, 16'd51534, 16'd20860, 16'd53787, 16'd12592, 16'd2557, 16'd53997, 16'd54166, 16'd25155, 16'd57661, 16'd57352, 16'd57201, 16'd48258, 16'd37407, 16'd16935, 16'd3499, 16'd27896, 16'd12840, 16'd7841, 16'd58496, 16'd47209});
	test_expansion(128'h9c218067f0fab0531b4b2d499c6b4ab9, {16'd7903, 16'd64684, 16'd59838, 16'd21817, 16'd6154, 16'd62890, 16'd46368, 16'd10265, 16'd24277, 16'd3376, 16'd41849, 16'd15546, 16'd59439, 16'd55387, 16'd32254, 16'd7270, 16'd41534, 16'd7214, 16'd25825, 16'd4888, 16'd27434, 16'd5312, 16'd20162, 16'd5276, 16'd53711, 16'd23622});
	test_expansion(128'h48148dbbdf70a7ad3ba9d2c8bc424f02, {16'd3442, 16'd63852, 16'd52424, 16'd5583, 16'd18513, 16'd1498, 16'd4112, 16'd49989, 16'd59139, 16'd48200, 16'd5248, 16'd6846, 16'd2940, 16'd50661, 16'd39771, 16'd2492, 16'd3217, 16'd50193, 16'd54358, 16'd13603, 16'd64718, 16'd27019, 16'd24038, 16'd19963, 16'd54770, 16'd13232});
	test_expansion(128'hd24380cd4956a9e7dc527646d3be2291, {16'd63975, 16'd57753, 16'd25572, 16'd57592, 16'd16358, 16'd9395, 16'd23605, 16'd54787, 16'd44058, 16'd59956, 16'd29899, 16'd24687, 16'd19643, 16'd6273, 16'd57191, 16'd15416, 16'd39279, 16'd59646, 16'd31760, 16'd4507, 16'd47996, 16'd9018, 16'd4928, 16'd22187, 16'd51001, 16'd60588});
	test_expansion(128'hfcdd7cbba787d6c458b4c8c8b51cf79a, {16'd30313, 16'd57651, 16'd5951, 16'd39371, 16'd52258, 16'd51085, 16'd50173, 16'd58401, 16'd51754, 16'd4056, 16'd63179, 16'd53835, 16'd7015, 16'd34961, 16'd3537, 16'd51693, 16'd20979, 16'd1931, 16'd60025, 16'd60236, 16'd58753, 16'd56380, 16'd62250, 16'd52594, 16'd46167, 16'd21482});
	test_expansion(128'hbc1916a26cdf3f2452e2661ff99c737c, {16'd37657, 16'd58600, 16'd7633, 16'd3550, 16'd43410, 16'd47350, 16'd34951, 16'd24586, 16'd60892, 16'd7302, 16'd14080, 16'd61803, 16'd27234, 16'd48466, 16'd9228, 16'd10699, 16'd6223, 16'd36028, 16'd9375, 16'd30253, 16'd25260, 16'd7902, 16'd61881, 16'd25227, 16'd38098, 16'd60849});
	test_expansion(128'h7dc0df4ab55a515fb0d1464e9623a792, {16'd7233, 16'd9147, 16'd55746, 16'd4046, 16'd5399, 16'd25829, 16'd59104, 16'd28534, 16'd36461, 16'd25442, 16'd61272, 16'd6171, 16'd37283, 16'd38779, 16'd35526, 16'd19539, 16'd55813, 16'd56059, 16'd54822, 16'd2059, 16'd21810, 16'd7998, 16'd64760, 16'd11151, 16'd31820, 16'd62252});
	test_expansion(128'hb8a18ed043b3dd3b985062ec74ac4eb6, {16'd29959, 16'd44029, 16'd4465, 16'd27720, 16'd59439, 16'd60038, 16'd21983, 16'd386, 16'd26275, 16'd63797, 16'd623, 16'd36866, 16'd5090, 16'd51687, 16'd6851, 16'd8387, 16'd15305, 16'd48163, 16'd5409, 16'd51782, 16'd5109, 16'd17023, 16'd2104, 16'd12185, 16'd57469, 16'd60677});
	test_expansion(128'h8961f437a3f5de1a5042bd2227e336d6, {16'd24058, 16'd36495, 16'd45851, 16'd59934, 16'd48138, 16'd22657, 16'd42969, 16'd48088, 16'd46811, 16'd39702, 16'd30343, 16'd34721, 16'd48621, 16'd6863, 16'd56466, 16'd53233, 16'd44409, 16'd58479, 16'd53148, 16'd55938, 16'd63769, 16'd28941, 16'd31090, 16'd51696, 16'd266, 16'd51180});
	test_expansion(128'h1a8ae18afa7a085b8711d48608180200, {16'd24956, 16'd23537, 16'd27490, 16'd24921, 16'd2693, 16'd34173, 16'd60864, 16'd14689, 16'd45993, 16'd30103, 16'd52188, 16'd7371, 16'd54718, 16'd4475, 16'd13984, 16'd710, 16'd29243, 16'd54501, 16'd25113, 16'd29500, 16'd58871, 16'd26041, 16'd53216, 16'd14309, 16'd22384, 16'd55802});
	test_expansion(128'hf1d0e3758e4016e254a4d8f9d8204af1, {16'd10962, 16'd15616, 16'd32239, 16'd41296, 16'd26011, 16'd11388, 16'd50152, 16'd65514, 16'd11233, 16'd26628, 16'd37841, 16'd5769, 16'd5958, 16'd41016, 16'd55643, 16'd27022, 16'd49722, 16'd15847, 16'd17530, 16'd39112, 16'd20999, 16'd47802, 16'd12380, 16'd61038, 16'd10063, 16'd23281});
	test_expansion(128'h66d8bb4751f3c6a5b7ea2fcd434d0c0c, {16'd10486, 16'd30470, 16'd30593, 16'd21126, 16'd34207, 16'd49005, 16'd44232, 16'd3602, 16'd13781, 16'd49047, 16'd9871, 16'd32843, 16'd42982, 16'd62248, 16'd59206, 16'd19019, 16'd50767, 16'd38933, 16'd53746, 16'd50935, 16'd9490, 16'd48765, 16'd9467, 16'd57865, 16'd5914, 16'd8859});
	test_expansion(128'h98a1097b20c045dc8cde6d198bb193c7, {16'd44676, 16'd22859, 16'd39189, 16'd14507, 16'd39783, 16'd23531, 16'd65263, 16'd4386, 16'd45129, 16'd53409, 16'd38359, 16'd8889, 16'd33629, 16'd16640, 16'd21844, 16'd1763, 16'd53550, 16'd9348, 16'd53962, 16'd13171, 16'd5597, 16'd23722, 16'd13712, 16'd5551, 16'd20634, 16'd41727});
	test_expansion(128'he5b3198fac8de7f11f0d683cb3185e2f, {16'd61239, 16'd64221, 16'd62225, 16'd50162, 16'd27399, 16'd31390, 16'd5536, 16'd58507, 16'd55350, 16'd8538, 16'd32210, 16'd5110, 16'd30739, 16'd50790, 16'd28335, 16'd3713, 16'd8930, 16'd22863, 16'd38562, 16'd45259, 16'd34831, 16'd28814, 16'd9043, 16'd44600, 16'd10013, 16'd16719});
	test_expansion(128'h052e5769558d421d38e523aa38dd12a1, {16'd25976, 16'd29766, 16'd60586, 16'd34882, 16'd48938, 16'd40067, 16'd37408, 16'd33278, 16'd31882, 16'd14452, 16'd6101, 16'd53601, 16'd32741, 16'd43960, 16'd53199, 16'd42266, 16'd1168, 16'd23433, 16'd47418, 16'd36250, 16'd62274, 16'd16242, 16'd9820, 16'd6722, 16'd45167, 16'd20604});
	test_expansion(128'h8029ee22cec617996afe9faa65579578, {16'd46889, 16'd27042, 16'd56822, 16'd1491, 16'd12523, 16'd23687, 16'd14415, 16'd16508, 16'd11893, 16'd25537, 16'd28098, 16'd492, 16'd15650, 16'd8219, 16'd16444, 16'd59595, 16'd26045, 16'd9766, 16'd54831, 16'd40984, 16'd35682, 16'd16535, 16'd18423, 16'd223, 16'd27188, 16'd41183});
	test_expansion(128'h267c5a253a9dbd015de653a17ba57230, {16'd27938, 16'd18035, 16'd44426, 16'd40596, 16'd31497, 16'd14239, 16'd39868, 16'd56334, 16'd34010, 16'd29744, 16'd56289, 16'd17526, 16'd58397, 16'd43009, 16'd39894, 16'd8302, 16'd42676, 16'd60056, 16'd15945, 16'd16352, 16'd59213, 16'd13301, 16'd14519, 16'd61418, 16'd11653, 16'd62134});
	test_expansion(128'hc653c840893718e47f382fcd855382e3, {16'd49365, 16'd35095, 16'd7570, 16'd14521, 16'd26697, 16'd23719, 16'd7791, 16'd15650, 16'd4302, 16'd56925, 16'd50995, 16'd20283, 16'd33887, 16'd11227, 16'd12839, 16'd49076, 16'd19854, 16'd3146, 16'd32739, 16'd37100, 16'd53047, 16'd5791, 16'd64778, 16'd36882, 16'd53830, 16'd54797});
	test_expansion(128'h7b7776ffe4cbe3333b219b90d6b043a6, {16'd6081, 16'd20892, 16'd12378, 16'd29469, 16'd8786, 16'd11308, 16'd23961, 16'd24405, 16'd21371, 16'd18376, 16'd45669, 16'd3197, 16'd50336, 16'd37334, 16'd36940, 16'd3016, 16'd20413, 16'd53971, 16'd37070, 16'd49267, 16'd8752, 16'd44135, 16'd49245, 16'd31126, 16'd19536, 16'd46807});
	test_expansion(128'h1b0391532f9ff02e01a120cd4babc963, {16'd48683, 16'd11355, 16'd9467, 16'd55688, 16'd1529, 16'd9554, 16'd33581, 16'd48717, 16'd32659, 16'd6551, 16'd27308, 16'd57262, 16'd48947, 16'd43427, 16'd7611, 16'd25865, 16'd27132, 16'd60963, 16'd37936, 16'd45839, 16'd1749, 16'd58653, 16'd28643, 16'd35966, 16'd28496, 16'd7783});
	test_expansion(128'h7667e4c7ef65a00bbfa4e5b9a87918ae, {16'd1824, 16'd3052, 16'd10284, 16'd13924, 16'd30675, 16'd28764, 16'd17840, 16'd35248, 16'd21214, 16'd33529, 16'd35068, 16'd51856, 16'd58201, 16'd53520, 16'd56986, 16'd21589, 16'd44132, 16'd39136, 16'd39225, 16'd55800, 16'd11337, 16'd40583, 16'd44786, 16'd45700, 16'd57468, 16'd8615});
	test_expansion(128'h4a9adf07a980112f84017c4437a7a848, {16'd55773, 16'd62657, 16'd60155, 16'd8508, 16'd51894, 16'd5620, 16'd46837, 16'd12413, 16'd5251, 16'd13267, 16'd11210, 16'd6142, 16'd51738, 16'd26913, 16'd35488, 16'd2805, 16'd1109, 16'd45980, 16'd5467, 16'd41528, 16'd5782, 16'd48380, 16'd1853, 16'd55005, 16'd48623, 16'd36657});
	test_expansion(128'ha9b71cc3ab8bd2dcd1682231b208a08c, {16'd49868, 16'd52025, 16'd29303, 16'd40337, 16'd39593, 16'd47997, 16'd58733, 16'd30962, 16'd56260, 16'd62841, 16'd32084, 16'd54731, 16'd27726, 16'd3888, 16'd54182, 16'd63182, 16'd39016, 16'd12309, 16'd3876, 16'd46413, 16'd49034, 16'd15915, 16'd50361, 16'd37882, 16'd36674, 16'd58800});
	test_expansion(128'h4318e7daaecbd9510611ba8c4ca3e67e, {16'd22417, 16'd53708, 16'd15967, 16'd51889, 16'd30420, 16'd60113, 16'd8512, 16'd60682, 16'd50082, 16'd62511, 16'd50262, 16'd46934, 16'd15687, 16'd27026, 16'd46319, 16'd57419, 16'd45319, 16'd32660, 16'd34642, 16'd12221, 16'd46436, 16'd43819, 16'd33727, 16'd55557, 16'd26165, 16'd18033});
	test_expansion(128'h05383cb8770f4c9311b5f426717f3b17, {16'd38563, 16'd56931, 16'd8715, 16'd29002, 16'd2362, 16'd62244, 16'd2070, 16'd34937, 16'd44370, 16'd2690, 16'd49352, 16'd32515, 16'd47300, 16'd46182, 16'd26876, 16'd43047, 16'd48727, 16'd60981, 16'd33243, 16'd20553, 16'd24631, 16'd10814, 16'd35445, 16'd1678, 16'd9102, 16'd642});
	test_expansion(128'hd305c1f1a8ba3ac35db9a33de0c1324e, {16'd4129, 16'd33140, 16'd1084, 16'd6444, 16'd31280, 16'd62580, 16'd35417, 16'd31074, 16'd55302, 16'd46583, 16'd37274, 16'd12592, 16'd31755, 16'd14081, 16'd52257, 16'd41729, 16'd50669, 16'd45338, 16'd42827, 16'd45551, 16'd11338, 16'd15327, 16'd39398, 16'd9153, 16'd5123, 16'd42249});
	test_expansion(128'he7b13bb37fa2200dfab9543e210af01b, {16'd48095, 16'd35008, 16'd57697, 16'd41971, 16'd19079, 16'd33651, 16'd26501, 16'd42223, 16'd12576, 16'd41527, 16'd7160, 16'd58913, 16'd57916, 16'd54590, 16'd54480, 16'd22068, 16'd29856, 16'd32801, 16'd39740, 16'd60051, 16'd2326, 16'd56587, 16'd57592, 16'd44798, 16'd22900, 16'd53840});
	test_expansion(128'hb391ba36d50068fdc78e5beef82926f3, {16'd59734, 16'd24057, 16'd24738, 16'd3024, 16'd30307, 16'd28826, 16'd40969, 16'd20511, 16'd53138, 16'd57086, 16'd14977, 16'd45429, 16'd26733, 16'd4018, 16'd47621, 16'd65518, 16'd55650, 16'd23281, 16'd41144, 16'd23308, 16'd23293, 16'd44434, 16'd930, 16'd8914, 16'd25280, 16'd33325});
	test_expansion(128'hccc0fba32681926c633e90daa23d410d, {16'd34578, 16'd48620, 16'd7084, 16'd33713, 16'd42747, 16'd50753, 16'd36251, 16'd53215, 16'd23748, 16'd28789, 16'd6768, 16'd29335, 16'd6614, 16'd43731, 16'd34474, 16'd6838, 16'd21456, 16'd57987, 16'd49561, 16'd23519, 16'd16339, 16'd24981, 16'd32536, 16'd10825, 16'd41911, 16'd60969});
	test_expansion(128'h490a76f3d32ec0e9cec23a3ab7138ae9, {16'd61403, 16'd31732, 16'd34957, 16'd1863, 16'd39186, 16'd14276, 16'd57540, 16'd56826, 16'd18565, 16'd64693, 16'd35910, 16'd56255, 16'd18356, 16'd54073, 16'd9218, 16'd46307, 16'd1164, 16'd35334, 16'd13100, 16'd17359, 16'd29605, 16'd58592, 16'd50666, 16'd21708, 16'd16905, 16'd24674});
	test_expansion(128'hc3a176ff0397212fcb12f37815919993, {16'd17372, 16'd9334, 16'd43805, 16'd27511, 16'd11090, 16'd24438, 16'd38012, 16'd63884, 16'd45116, 16'd24764, 16'd17157, 16'd14, 16'd63415, 16'd21107, 16'd2517, 16'd56363, 16'd54515, 16'd64892, 16'd23414, 16'd25794, 16'd65365, 16'd6815, 16'd58876, 16'd11939, 16'd15985, 16'd9687});
	test_expansion(128'h980b5e4b5240cf23777b735d84b0af61, {16'd800, 16'd10900, 16'd15725, 16'd21716, 16'd12667, 16'd51074, 16'd33332, 16'd56815, 16'd59311, 16'd61288, 16'd43333, 16'd4525, 16'd14302, 16'd48763, 16'd28345, 16'd34936, 16'd39695, 16'd57495, 16'd2808, 16'd50909, 16'd43121, 16'd12856, 16'd46083, 16'd31584, 16'd37730, 16'd18424});
	test_expansion(128'h9c8176a8c3cb051081bf9d22ea13cb6a, {16'd24973, 16'd21627, 16'd64442, 16'd33944, 16'd19461, 16'd51393, 16'd10116, 16'd1472, 16'd476, 16'd36206, 16'd28716, 16'd1701, 16'd26431, 16'd13802, 16'd62444, 16'd37006, 16'd47944, 16'd47338, 16'd41243, 16'd61163, 16'd8410, 16'd22018, 16'd13198, 16'd8062, 16'd29754, 16'd59120});
	test_expansion(128'h51c9f9ba56e1d3716d3886d386648952, {16'd27682, 16'd4366, 16'd43999, 16'd60368, 16'd36147, 16'd39115, 16'd35053, 16'd14965, 16'd16065, 16'd33201, 16'd47922, 16'd16985, 16'd25077, 16'd7432, 16'd41694, 16'd28796, 16'd56386, 16'd63120, 16'd59773, 16'd23675, 16'd48807, 16'd56058, 16'd54668, 16'd53511, 16'd58444, 16'd24266});
	test_expansion(128'hc7125e603ffc0ba2c62789b1ce6dc47a, {16'd30584, 16'd51921, 16'd62054, 16'd6403, 16'd29552, 16'd18781, 16'd56739, 16'd12160, 16'd8725, 16'd28057, 16'd23664, 16'd13736, 16'd33994, 16'd20879, 16'd40588, 16'd19533, 16'd65211, 16'd484, 16'd36061, 16'd26247, 16'd46625, 16'd50399, 16'd64902, 16'd11258, 16'd44321, 16'd39752});
	test_expansion(128'h7d7e4dd04f07fac092a5344a28238554, {16'd48950, 16'd14296, 16'd37234, 16'd4456, 16'd9238, 16'd25836, 16'd32989, 16'd47001, 16'd28546, 16'd63279, 16'd15645, 16'd6706, 16'd20667, 16'd44175, 16'd11871, 16'd42620, 16'd24, 16'd40385, 16'd34120, 16'd62330, 16'd3581, 16'd57518, 16'd47953, 16'd61805, 16'd12667, 16'd61478});
	test_expansion(128'hb74cdbc0211674f3ad29839ad5c97c36, {16'd16355, 16'd12020, 16'd8259, 16'd49069, 16'd48142, 16'd599, 16'd20858, 16'd36518, 16'd62061, 16'd8602, 16'd25426, 16'd9627, 16'd16317, 16'd1674, 16'd45362, 16'd49611, 16'd28098, 16'd33485, 16'd51012, 16'd49075, 16'd48655, 16'd5545, 16'd11314, 16'd52474, 16'd64882, 16'd62660});
	test_expansion(128'h642a641becbc6ae824c70518a5d490c5, {16'd45893, 16'd30383, 16'd31632, 16'd19331, 16'd3028, 16'd19438, 16'd43932, 16'd55972, 16'd42646, 16'd6051, 16'd51479, 16'd29661, 16'd22568, 16'd2185, 16'd6543, 16'd39965, 16'd32641, 16'd39432, 16'd39173, 16'd7888, 16'd63707, 16'd19031, 16'd55134, 16'd61367, 16'd34524, 16'd41736});
	test_expansion(128'hdbe5f62f0940f5c6e024e5b471d0d178, {16'd32524, 16'd60513, 16'd46627, 16'd8833, 16'd20587, 16'd41828, 16'd12235, 16'd37595, 16'd6716, 16'd11402, 16'd59602, 16'd55894, 16'd48640, 16'd5824, 16'd24790, 16'd27304, 16'd40420, 16'd37617, 16'd16853, 16'd43701, 16'd34463, 16'd15809, 16'd63468, 16'd22348, 16'd50068, 16'd49072});
	test_expansion(128'h31aa9ab39dd903c0825b549445b048ee, {16'd6765, 16'd45391, 16'd18294, 16'd1420, 16'd11523, 16'd7645, 16'd16284, 16'd61685, 16'd27407, 16'd62876, 16'd48344, 16'd37478, 16'd63247, 16'd22206, 16'd4463, 16'd32262, 16'd56415, 16'd47439, 16'd4071, 16'd52465, 16'd51996, 16'd3510, 16'd38581, 16'd9677, 16'd65346, 16'd1261});
	test_expansion(128'h24fefa853991192350951e290ca78ad2, {16'd19574, 16'd48435, 16'd31039, 16'd59723, 16'd7665, 16'd5434, 16'd60271, 16'd34080, 16'd814, 16'd29925, 16'd15569, 16'd3873, 16'd40586, 16'd50806, 16'd32468, 16'd50054, 16'd13842, 16'd28274, 16'd62852, 16'd15471, 16'd55479, 16'd10501, 16'd9665, 16'd44736, 16'd53048, 16'd49829});
	test_expansion(128'h89b890559b93c8c73c4419373fbae81b, {16'd21411, 16'd35292, 16'd39543, 16'd25050, 16'd4088, 16'd32173, 16'd44503, 16'd30334, 16'd48525, 16'd41107, 16'd23874, 16'd42146, 16'd64721, 16'd30639, 16'd50083, 16'd4346, 16'd54802, 16'd13852, 16'd33399, 16'd40715, 16'd53605, 16'd10592, 16'd65199, 16'd24300, 16'd63060, 16'd8125});
	test_expansion(128'h647afeed2683413121524f15f263aa0e, {16'd58059, 16'd36002, 16'd23886, 16'd36018, 16'd7551, 16'd37103, 16'd4538, 16'd11105, 16'd60274, 16'd17779, 16'd25060, 16'd46093, 16'd58721, 16'd15135, 16'd56123, 16'd61305, 16'd5442, 16'd57766, 16'd30087, 16'd3923, 16'd23042, 16'd46428, 16'd59284, 16'd54017, 16'd13533, 16'd55763});
	test_expansion(128'h74462755a7a91f962ac50f3cf03b0efd, {16'd35643, 16'd22068, 16'd24682, 16'd4708, 16'd46005, 16'd46920, 16'd56897, 16'd262, 16'd55132, 16'd63007, 16'd21075, 16'd40874, 16'd20785, 16'd28030, 16'd45687, 16'd63882, 16'd65483, 16'd41317, 16'd1408, 16'd16442, 16'd36258, 16'd19397, 16'd15270, 16'd9283, 16'd51616, 16'd59085});
	test_expansion(128'h24aa65774179c91d01706de61b5a30eb, {16'd12533, 16'd61606, 16'd47965, 16'd14440, 16'd33276, 16'd62444, 16'd22218, 16'd28467, 16'd52268, 16'd4199, 16'd61885, 16'd60725, 16'd20376, 16'd31236, 16'd64775, 16'd15596, 16'd25224, 16'd34561, 16'd3097, 16'd44102, 16'd58137, 16'd40130, 16'd4730, 16'd45223, 16'd43767, 16'd2230});
	test_expansion(128'ha695964ccc79eb02661dab8b52e8c6ab, {16'd11855, 16'd23752, 16'd5112, 16'd37657, 16'd51348, 16'd52050, 16'd43833, 16'd33891, 16'd46516, 16'd39849, 16'd63344, 16'd22956, 16'd48393, 16'd46220, 16'd46203, 16'd8077, 16'd50424, 16'd46018, 16'd38042, 16'd49506, 16'd22370, 16'd7262, 16'd10299, 16'd47694, 16'd16156, 16'd47057});
	test_expansion(128'h6d5d9a29c98dc0d818e2f8f8cd3891b2, {16'd56109, 16'd16842, 16'd13527, 16'd55852, 16'd33803, 16'd39745, 16'd4917, 16'd5225, 16'd48557, 16'd6825, 16'd57978, 16'd24677, 16'd43337, 16'd7136, 16'd58823, 16'd62729, 16'd38987, 16'd28882, 16'd24406, 16'd19799, 16'd62399, 16'd56882, 16'd64353, 16'd19503, 16'd6849, 16'd21802});
	test_expansion(128'hf334d5cfd193f8057913d050a0a3fa44, {16'd31097, 16'd17227, 16'd26374, 16'd34260, 16'd21358, 16'd42679, 16'd6273, 16'd60385, 16'd9974, 16'd15597, 16'd48699, 16'd6922, 16'd45345, 16'd55389, 16'd24859, 16'd5757, 16'd30176, 16'd58354, 16'd60859, 16'd40434, 16'd32900, 16'd5035, 16'd41078, 16'd21575, 16'd58096, 16'd15024});
	test_expansion(128'hca3f1faaf79d4ab2afd141d39cbc2536, {16'd50209, 16'd15254, 16'd52473, 16'd35117, 16'd39168, 16'd18233, 16'd60941, 16'd44911, 16'd39890, 16'd2929, 16'd54134, 16'd17995, 16'd21954, 16'd61821, 16'd6953, 16'd56726, 16'd6402, 16'd18782, 16'd13461, 16'd57312, 16'd62909, 16'd57648, 16'd47975, 16'd3751, 16'd47023, 16'd24820});
	test_expansion(128'he93c7c3f462f1a1feeff78d6ca8883b5, {16'd27269, 16'd35190, 16'd32797, 16'd13003, 16'd1607, 16'd34493, 16'd53503, 16'd54194, 16'd6156, 16'd47517, 16'd17179, 16'd64180, 16'd36736, 16'd21531, 16'd19176, 16'd18674, 16'd52472, 16'd15161, 16'd56913, 16'd34, 16'd46459, 16'd13706, 16'd22736, 16'd49955, 16'd43669, 16'd40964});
	test_expansion(128'h8e1c0caeb679aeacabe2f7d1140a98ae, {16'd8302, 16'd62241, 16'd60681, 16'd33497, 16'd40406, 16'd63784, 16'd35780, 16'd39581, 16'd6534, 16'd43133, 16'd34040, 16'd12371, 16'd55227, 16'd24814, 16'd33368, 16'd25794, 16'd26847, 16'd49329, 16'd52159, 16'd10436, 16'd30753, 16'd55730, 16'd26380, 16'd64525, 16'd47315, 16'd40116});
	test_expansion(128'h2854f048f8613ea7374c7765f07f9757, {16'd60276, 16'd52955, 16'd2360, 16'd22462, 16'd64847, 16'd55429, 16'd33908, 16'd42075, 16'd47506, 16'd58747, 16'd42546, 16'd54021, 16'd23681, 16'd64735, 16'd21008, 16'd6100, 16'd53113, 16'd55227, 16'd9225, 16'd49502, 16'd25695, 16'd11625, 16'd31274, 16'd7244, 16'd39414, 16'd26491});
	test_expansion(128'hc6ce36a19e822ac95658e599268ee18b, {16'd3042, 16'd17715, 16'd46374, 16'd19506, 16'd65053, 16'd43360, 16'd34871, 16'd31444, 16'd29123, 16'd12512, 16'd7840, 16'd64798, 16'd37081, 16'd60104, 16'd48428, 16'd10276, 16'd48641, 16'd33462, 16'd38381, 16'd213, 16'd29215, 16'd10490, 16'd59565, 16'd22151, 16'd14897, 16'd53933});
	test_expansion(128'ha0c40f51f39e6d4015c46371cea5f975, {16'd37290, 16'd50023, 16'd44644, 16'd54473, 16'd59083, 16'd6354, 16'd58081, 16'd19791, 16'd34649, 16'd41222, 16'd59643, 16'd42152, 16'd47143, 16'd53945, 16'd11078, 16'd42003, 16'd13643, 16'd54946, 16'd58052, 16'd46488, 16'd34122, 16'd36270, 16'd24337, 16'd38496, 16'd45035, 16'd26387});
	test_expansion(128'hbbf3348560392f9dae6e3a9f2fefed2a, {16'd15192, 16'd37752, 16'd7941, 16'd41285, 16'd22272, 16'd16708, 16'd42808, 16'd14815, 16'd64439, 16'd1960, 16'd29815, 16'd59431, 16'd11543, 16'd42520, 16'd56424, 16'd46352, 16'd37197, 16'd27221, 16'd58224, 16'd8073, 16'd63518, 16'd11980, 16'd27971, 16'd4378, 16'd48983, 16'd40723});
	test_expansion(128'h3e0043024743b383693490ff65d492b6, {16'd57402, 16'd21603, 16'd29925, 16'd63376, 16'd32950, 16'd21731, 16'd34647, 16'd26223, 16'd61084, 16'd3058, 16'd34248, 16'd743, 16'd60273, 16'd49837, 16'd7000, 16'd21187, 16'd53382, 16'd53367, 16'd48090, 16'd12642, 16'd7745, 16'd35499, 16'd10496, 16'd44323, 16'd41512, 16'd41972});
	test_expansion(128'h58e12c9521b6100ee38ccc28f0c503da, {16'd31580, 16'd39325, 16'd3874, 16'd63178, 16'd33807, 16'd53258, 16'd48222, 16'd6722, 16'd4410, 16'd35938, 16'd41405, 16'd52784, 16'd5773, 16'd5210, 16'd53503, 16'd3317, 16'd61250, 16'd63319, 16'd57946, 16'd7362, 16'd5789, 16'd54782, 16'd60800, 16'd60140, 16'd39013, 16'd35826});
	test_expansion(128'hd0c9eb97e824d8b8dd98dc5697e2e9fc, {16'd25656, 16'd2412, 16'd36096, 16'd23687, 16'd35564, 16'd30719, 16'd8484, 16'd16940, 16'd3127, 16'd345, 16'd46855, 16'd42531, 16'd34901, 16'd36568, 16'd54205, 16'd50462, 16'd36972, 16'd41480, 16'd3277, 16'd16204, 16'd55260, 16'd24369, 16'd26985, 16'd18512, 16'd37658, 16'd21911});
	test_expansion(128'he406fe9e3178e18d208a8305d38e5362, {16'd53188, 16'd51936, 16'd3228, 16'd47544, 16'd31013, 16'd37706, 16'd9646, 16'd48677, 16'd8215, 16'd45936, 16'd9780, 16'd41854, 16'd51592, 16'd13092, 16'd49564, 16'd10314, 16'd13060, 16'd40469, 16'd59437, 16'd8387, 16'd30185, 16'd39027, 16'd62052, 16'd32239, 16'd47187, 16'd26445});
	test_expansion(128'hcd9d7f4d6fc22db620aed7e96e79228e, {16'd43157, 16'd36794, 16'd38801, 16'd45720, 16'd36009, 16'd51145, 16'd11181, 16'd59297, 16'd13011, 16'd20406, 16'd6808, 16'd38385, 16'd18415, 16'd56562, 16'd20196, 16'd64503, 16'd16577, 16'd17290, 16'd11739, 16'd4001, 16'd21793, 16'd5244, 16'd13372, 16'd57075, 16'd11361, 16'd33439});
	test_expansion(128'hff9b18b0a0e0f90bcf15e7d001d410c0, {16'd49311, 16'd54286, 16'd36157, 16'd3447, 16'd285, 16'd61487, 16'd62787, 16'd130, 16'd32316, 16'd6866, 16'd14802, 16'd42897, 16'd61185, 16'd49822, 16'd35185, 16'd56422, 16'd56400, 16'd38529, 16'd404, 16'd62381, 16'd13555, 16'd26542, 16'd35191, 16'd62052, 16'd8128, 16'd39800});
	test_expansion(128'h5a503ddcd44b647645fa00a26a9f6033, {16'd41591, 16'd41611, 16'd9140, 16'd18926, 16'd17530, 16'd42118, 16'd25576, 16'd61390, 16'd65193, 16'd33050, 16'd32420, 16'd15141, 16'd23554, 16'd48097, 16'd26387, 16'd33155, 16'd10436, 16'd61885, 16'd20338, 16'd2891, 16'd7712, 16'd61246, 16'd35789, 16'd21029, 16'd37964, 16'd43983});
	test_expansion(128'hea2d843c4ddf4b0ea164801e4a396494, {16'd30660, 16'd22377, 16'd27039, 16'd41657, 16'd3832, 16'd19354, 16'd58788, 16'd32748, 16'd30655, 16'd47267, 16'd2675, 16'd64641, 16'd42020, 16'd60443, 16'd24180, 16'd24512, 16'd43372, 16'd15890, 16'd34867, 16'd16929, 16'd61263, 16'd24658, 16'd3737, 16'd22168, 16'd40524, 16'd12787});
	test_expansion(128'h1857ed54e9c36a1350b7743b467fa8fd, {16'd46557, 16'd42111, 16'd48452, 16'd32235, 16'd50955, 16'd13634, 16'd13256, 16'd15197, 16'd32095, 16'd8097, 16'd6554, 16'd36810, 16'd34991, 16'd34580, 16'd30927, 16'd3521, 16'd9994, 16'd43129, 16'd53896, 16'd20131, 16'd59654, 16'd49189, 16'd13877, 16'd23851, 16'd16943, 16'd54060});
	test_expansion(128'hff75e9e66951906f4f587fab048ad80f, {16'd32803, 16'd55968, 16'd39794, 16'd61314, 16'd64891, 16'd59027, 16'd61662, 16'd53568, 16'd5075, 16'd35942, 16'd17446, 16'd21412, 16'd18683, 16'd62760, 16'd51590, 16'd55664, 16'd32239, 16'd48859, 16'd467, 16'd50372, 16'd30174, 16'd35702, 16'd5572, 16'd47327, 16'd23358, 16'd47017});
	test_expansion(128'h7fc0cd7aa89b969115351bdfc7105e98, {16'd23725, 16'd55633, 16'd6790, 16'd49065, 16'd9716, 16'd20520, 16'd34274, 16'd21700, 16'd60007, 16'd24034, 16'd21384, 16'd62602, 16'd11568, 16'd62048, 16'd57071, 16'd8032, 16'd49481, 16'd49009, 16'd57433, 16'd24576, 16'd20278, 16'd47886, 16'd16016, 16'd35121, 16'd57000, 16'd3885});
	test_expansion(128'h3ac9dc8d0429b77f9edc0d4b811282b4, {16'd47736, 16'd7181, 16'd27937, 16'd6896, 16'd6266, 16'd32081, 16'd20372, 16'd35463, 16'd30118, 16'd5402, 16'd59363, 16'd30233, 16'd46148, 16'd36278, 16'd5694, 16'd30392, 16'd38495, 16'd16851, 16'd13982, 16'd50220, 16'd51555, 16'd3703, 16'd62643, 16'd49737, 16'd64648, 16'd63216});
	test_expansion(128'h7be534d7fee3aaac053caf3b45ac6c4b, {16'd43142, 16'd15576, 16'd38598, 16'd9078, 16'd1779, 16'd39521, 16'd12015, 16'd50321, 16'd20483, 16'd11639, 16'd13227, 16'd60827, 16'd40513, 16'd21534, 16'd60506, 16'd24539, 16'd17976, 16'd50830, 16'd55649, 16'd30126, 16'd481, 16'd27088, 16'd31121, 16'd914, 16'd36849, 16'd57595});
	test_expansion(128'h97fa2aa0ab4363f912acc18a1909340c, {16'd62024, 16'd31829, 16'd48931, 16'd10358, 16'd45084, 16'd35340, 16'd30488, 16'd26968, 16'd63184, 16'd12203, 16'd22708, 16'd53731, 16'd46767, 16'd61123, 16'd54830, 16'd20677, 16'd14525, 16'd26401, 16'd36892, 16'd57379, 16'd8051, 16'd63611, 16'd53975, 16'd8422, 16'd2394, 16'd36485});
	test_expansion(128'hd08560c66e875700ed53a89b4cd34ba8, {16'd11701, 16'd65437, 16'd29448, 16'd3677, 16'd41132, 16'd42651, 16'd23594, 16'd11826, 16'd63153, 16'd35758, 16'd51969, 16'd25974, 16'd25349, 16'd36159, 16'd41676, 16'd33512, 16'd31972, 16'd58291, 16'd63457, 16'd49464, 16'd49037, 16'd50603, 16'd5689, 16'd22983, 16'd48079, 16'd54577});
	test_expansion(128'hdd9cf950dcb33867e87968ce213fcb47, {16'd39567, 16'd42666, 16'd12873, 16'd32973, 16'd59069, 16'd18900, 16'd60665, 16'd16828, 16'd24424, 16'd40999, 16'd59739, 16'd32191, 16'd29195, 16'd7816, 16'd38779, 16'd51933, 16'd18415, 16'd14290, 16'd49985, 16'd43062, 16'd10554, 16'd56838, 16'd129, 16'd31980, 16'd27693, 16'd13938});
	test_expansion(128'h2434e680398c605437b3c77aad672032, {16'd38401, 16'd53598, 16'd8922, 16'd12195, 16'd58958, 16'd54055, 16'd6102, 16'd50010, 16'd29766, 16'd50168, 16'd26081, 16'd19850, 16'd41735, 16'd34788, 16'd62179, 16'd5251, 16'd27392, 16'd19242, 16'd7429, 16'd61791, 16'd39299, 16'd31317, 16'd11572, 16'd1030, 16'd28467, 16'd57071});
	test_expansion(128'h2e8c2c8888fe495b6b944986ef7580e7, {16'd40577, 16'd28918, 16'd9039, 16'd54694, 16'd920, 16'd4674, 16'd57788, 16'd19959, 16'd52378, 16'd20046, 16'd32035, 16'd17412, 16'd61645, 16'd51300, 16'd16593, 16'd29585, 16'd48905, 16'd54911, 16'd19188, 16'd56156, 16'd55865, 16'd26002, 16'd11799, 16'd6504, 16'd4618, 16'd38415});
	test_expansion(128'h97257037fa6c57f5566bbea8e60c356f, {16'd59193, 16'd34009, 16'd10309, 16'd38565, 16'd45460, 16'd57868, 16'd65497, 16'd16808, 16'd20752, 16'd42437, 16'd38248, 16'd12969, 16'd2586, 16'd60581, 16'd44833, 16'd43201, 16'd35755, 16'd9068, 16'd1861, 16'd39664, 16'd19667, 16'd42979, 16'd9946, 16'd63105, 16'd46549, 16'd34495});
	test_expansion(128'hcd2c09814aa310a6bb4f061a4535ab55, {16'd43084, 16'd18876, 16'd61649, 16'd64007, 16'd34532, 16'd10299, 16'd11298, 16'd15590, 16'd50616, 16'd8891, 16'd34956, 16'd22846, 16'd50768, 16'd56151, 16'd45746, 16'd22476, 16'd8458, 16'd55753, 16'd9956, 16'd20113, 16'd57327, 16'd64884, 16'd12235, 16'd8835, 16'd55795, 16'd11638});
	test_expansion(128'hfca21e50c3d2617d8a52d955cb0c60e2, {16'd32669, 16'd14211, 16'd60260, 16'd9302, 16'd46937, 16'd12865, 16'd23672, 16'd533, 16'd21076, 16'd20612, 16'd60378, 16'd54750, 16'd9988, 16'd22957, 16'd62494, 16'd48811, 16'd40083, 16'd50401, 16'd44038, 16'd30824, 16'd4820, 16'd58120, 16'd30639, 16'd18679, 16'd33574, 16'd59066});
	test_expansion(128'h9647d63b413cb2babbd69022cda02bbc, {16'd60729, 16'd48793, 16'd58757, 16'd61038, 16'd27535, 16'd1043, 16'd57204, 16'd24432, 16'd21660, 16'd14045, 16'd6298, 16'd15100, 16'd38088, 16'd59020, 16'd62883, 16'd9156, 16'd12985, 16'd58263, 16'd33155, 16'd8409, 16'd24558, 16'd18583, 16'd39112, 16'd4547, 16'd65346, 16'd36642});
	test_expansion(128'h441b74c0ea00936b9c2b03e136d069a1, {16'd8213, 16'd46308, 16'd12794, 16'd54627, 16'd38952, 16'd65231, 16'd33673, 16'd53043, 16'd6931, 16'd39555, 16'd11452, 16'd40199, 16'd34715, 16'd20540, 16'd54688, 16'd96, 16'd14043, 16'd9529, 16'd30807, 16'd62241, 16'd62635, 16'd63600, 16'd19619, 16'd13560, 16'd28157, 16'd7484});
	test_expansion(128'h6bf5d0e13bde95dd98f045c874696106, {16'd45021, 16'd14757, 16'd339, 16'd52111, 16'd17279, 16'd2480, 16'd4162, 16'd44778, 16'd20628, 16'd58142, 16'd25400, 16'd2739, 16'd38765, 16'd40415, 16'd40723, 16'd19417, 16'd58060, 16'd7362, 16'd29551, 16'd18551, 16'd12655, 16'd48096, 16'd39874, 16'd14747, 16'd7158, 16'd34462});
	test_expansion(128'hd1c97e55b48735074335b999dd68da4f, {16'd52005, 16'd13334, 16'd45500, 16'd31395, 16'd2821, 16'd20040, 16'd50628, 16'd59564, 16'd49524, 16'd51147, 16'd41944, 16'd47107, 16'd18335, 16'd61693, 16'd47913, 16'd3148, 16'd42247, 16'd15523, 16'd24486, 16'd18211, 16'd4284, 16'd46291, 16'd55851, 16'd34022, 16'd43630, 16'd32394});
	test_expansion(128'h498c08403b6565350b3e453f95f52453, {16'd18646, 16'd39432, 16'd28876, 16'd41293, 16'd50224, 16'd64799, 16'd14761, 16'd56632, 16'd25544, 16'd39630, 16'd34517, 16'd46106, 16'd32959, 16'd44738, 16'd33397, 16'd63152, 16'd48994, 16'd27586, 16'd60595, 16'd4514, 16'd19862, 16'd51404, 16'd4671, 16'd30464, 16'd65265, 16'd4154});
	test_expansion(128'h15859d87470c9ec05a6546729131f60c, {16'd13266, 16'd53707, 16'd8808, 16'd68, 16'd27293, 16'd6505, 16'd37933, 16'd26830, 16'd44746, 16'd48353, 16'd17834, 16'd11322, 16'd5970, 16'd15907, 16'd53878, 16'd25693, 16'd48198, 16'd54714, 16'd52535, 16'd61479, 16'd43764, 16'd6187, 16'd54959, 16'd25400, 16'd18187, 16'd64558});
	test_expansion(128'h5ab02d0f2133b71a3aa56de2dc5d8bdc, {16'd53341, 16'd29567, 16'd17212, 16'd7548, 16'd49347, 16'd55386, 16'd46855, 16'd50247, 16'd12430, 16'd44503, 16'd31940, 16'd34984, 16'd55543, 16'd7277, 16'd13753, 16'd60450, 16'd41584, 16'd28548, 16'd46973, 16'd15671, 16'd13303, 16'd58046, 16'd35192, 16'd33352, 16'd57389, 16'd57126});
	test_expansion(128'hba1a6deca940636ba6240e9fca9d9e40, {16'd56147, 16'd8054, 16'd48821, 16'd31192, 16'd54996, 16'd36443, 16'd3602, 16'd23394, 16'd60754, 16'd34848, 16'd7829, 16'd37010, 16'd53680, 16'd48142, 16'd13761, 16'd56612, 16'd44331, 16'd23, 16'd40042, 16'd42353, 16'd35155, 16'd50500, 16'd40366, 16'd29411, 16'd27246, 16'd29561});
	test_expansion(128'hbcbd3c1a8306afdb7ded8527f51bbd4e, {16'd24064, 16'd55447, 16'd56667, 16'd43269, 16'd24369, 16'd8041, 16'd55255, 16'd13974, 16'd111, 16'd22156, 16'd13930, 16'd49218, 16'd1397, 16'd34151, 16'd37766, 16'd36241, 16'd12578, 16'd41667, 16'd57697, 16'd9685, 16'd24635, 16'd35577, 16'd59815, 16'd58621, 16'd32676, 16'd7865});
	test_expansion(128'he27be58545dcb88b50ad5be5bd58a74d, {16'd15771, 16'd36882, 16'd17502, 16'd2124, 16'd5655, 16'd6194, 16'd16714, 16'd51193, 16'd41328, 16'd21388, 16'd8632, 16'd11748, 16'd12662, 16'd54807, 16'd11142, 16'd64326, 16'd37302, 16'd23392, 16'd6802, 16'd6632, 16'd3454, 16'd42036, 16'd64078, 16'd21169, 16'd32957, 16'd40642});
	test_expansion(128'h4bbd17df95d1cb08aa6c252ea79b0ab7, {16'd49072, 16'd41753, 16'd12552, 16'd28716, 16'd30773, 16'd24846, 16'd51784, 16'd37472, 16'd49906, 16'd64331, 16'd10790, 16'd55138, 16'd39947, 16'd15518, 16'd7388, 16'd49320, 16'd1924, 16'd43688, 16'd5651, 16'd45549, 16'd14679, 16'd58282, 16'd34194, 16'd9047, 16'd51665, 16'd37261});
	test_expansion(128'hd167541133056367f0c0073c3a8d6af7, {16'd32316, 16'd39584, 16'd40009, 16'd19689, 16'd19928, 16'd20236, 16'd50400, 16'd32817, 16'd20345, 16'd53304, 16'd54045, 16'd53915, 16'd3285, 16'd59626, 16'd18308, 16'd57391, 16'd25260, 16'd272, 16'd7919, 16'd57341, 16'd59504, 16'd53459, 16'd38578, 16'd52016, 16'd46692, 16'd53860});
	test_expansion(128'h71ea94180479a4d9dc0c1d7acc301747, {16'd57542, 16'd45854, 16'd16460, 16'd59765, 16'd61802, 16'd47388, 16'd36862, 16'd18785, 16'd3405, 16'd17587, 16'd38235, 16'd56440, 16'd45397, 16'd31407, 16'd31365, 16'd29397, 16'd18226, 16'd275, 16'd19512, 16'd37244, 16'd41222, 16'd63795, 16'd13650, 16'd60665, 16'd48570, 16'd34020});
	test_expansion(128'h271c1e0879f34d3931864c60f99ff092, {16'd63343, 16'd33900, 16'd64951, 16'd55245, 16'd12767, 16'd48994, 16'd27620, 16'd30404, 16'd43653, 16'd33543, 16'd58023, 16'd32042, 16'd65296, 16'd44164, 16'd49339, 16'd2453, 16'd41361, 16'd32086, 16'd28549, 16'd50740, 16'd32640, 16'd63006, 16'd46635, 16'd490, 16'd32719, 16'd60861});
	test_expansion(128'h3a20950e175b8fb9594c5c03563bd19e, {16'd17021, 16'd51582, 16'd64624, 16'd13361, 16'd6561, 16'd2259, 16'd25624, 16'd22300, 16'd15761, 16'd35827, 16'd35457, 16'd22924, 16'd39906, 16'd15325, 16'd64531, 16'd51312, 16'd65295, 16'd23849, 16'd65155, 16'd18314, 16'd38408, 16'd6210, 16'd59391, 16'd45791, 16'd41122, 16'd7555});
	test_expansion(128'he2ab3d6d87ce3f2366785b5a4cde9d30, {16'd775, 16'd13774, 16'd31045, 16'd36841, 16'd14052, 16'd46825, 16'd44618, 16'd18688, 16'd26105, 16'd4918, 16'd60884, 16'd47444, 16'd32915, 16'd33477, 16'd54746, 16'd40522, 16'd45416, 16'd53311, 16'd11800, 16'd59305, 16'd53717, 16'd23445, 16'd39020, 16'd24968, 16'd57444, 16'd11693});
	test_expansion(128'hcb26b1fc1c39418de7990bb1d86e968f, {16'd16455, 16'd43188, 16'd46844, 16'd36520, 16'd53509, 16'd11032, 16'd42894, 16'd3140, 16'd55550, 16'd22929, 16'd48494, 16'd40486, 16'd44366, 16'd4732, 16'd44255, 16'd39704, 16'd34123, 16'd45820, 16'd4508, 16'd13879, 16'd9283, 16'd2061, 16'd64183, 16'd31310, 16'd21285, 16'd39398});
	test_expansion(128'hbd81561bb8c9cc687d6fb0fd76373f68, {16'd42873, 16'd42602, 16'd27313, 16'd44947, 16'd3428, 16'd41162, 16'd55032, 16'd11111, 16'd40350, 16'd37305, 16'd23555, 16'd48544, 16'd15965, 16'd17912, 16'd26933, 16'd49772, 16'd12583, 16'd37475, 16'd61211, 16'd37674, 16'd53616, 16'd2181, 16'd31480, 16'd58014, 16'd51904, 16'd62782});
	test_expansion(128'h88de69b80b0b7ee4b740f2a894519569, {16'd64239, 16'd57628, 16'd2021, 16'd17144, 16'd5946, 16'd6665, 16'd27287, 16'd17399, 16'd50962, 16'd53290, 16'd2274, 16'd31605, 16'd11089, 16'd33992, 16'd17710, 16'd60554, 16'd21988, 16'd29115, 16'd58225, 16'd42402, 16'd8427, 16'd474, 16'd8089, 16'd62257, 16'd6064, 16'd58899});
	test_expansion(128'h7e6e34060d6e7264e15c9f8f4559dbe1, {16'd53039, 16'd38253, 16'd45395, 16'd16674, 16'd1048, 16'd61986, 16'd21416, 16'd28985, 16'd56175, 16'd12446, 16'd26353, 16'd15652, 16'd60252, 16'd57084, 16'd42382, 16'd14283, 16'd40269, 16'd15581, 16'd54874, 16'd21082, 16'd13336, 16'd25112, 16'd13570, 16'd16028, 16'd33138, 16'd31750});
	test_expansion(128'h8a9fd194adc4b332311e4dcd8c5c0314, {16'd31869, 16'd869, 16'd50108, 16'd60906, 16'd18629, 16'd2, 16'd59249, 16'd35519, 16'd40626, 16'd20084, 16'd17665, 16'd34037, 16'd50728, 16'd35984, 16'd54397, 16'd29966, 16'd64490, 16'd58962, 16'd64480, 16'd25384, 16'd50549, 16'd21702, 16'd54822, 16'd995, 16'd56742, 16'd2984});
	test_expansion(128'hcd6cc19ead2fd8b908d2930c50072110, {16'd4742, 16'd56351, 16'd36075, 16'd9692, 16'd58481, 16'd27014, 16'd37400, 16'd46734, 16'd47684, 16'd28376, 16'd63678, 16'd29414, 16'd60945, 16'd37031, 16'd42413, 16'd7197, 16'd26525, 16'd31880, 16'd44885, 16'd62800, 16'd17682, 16'd40710, 16'd27695, 16'd62411, 16'd60172, 16'd17091});
	test_expansion(128'h4c5b41f4dc65441f405a77286668be15, {16'd25012, 16'd14951, 16'd26467, 16'd56864, 16'd20604, 16'd64107, 16'd50730, 16'd8371, 16'd39762, 16'd52678, 16'd47253, 16'd63412, 16'd37466, 16'd54469, 16'd44906, 16'd36616, 16'd28013, 16'd62102, 16'd44576, 16'd51641, 16'd15734, 16'd38662, 16'd42208, 16'd25686, 16'd41681, 16'd2107});
	test_expansion(128'h57244a18ec1ba189ce151795687b122a, {16'd50263, 16'd35830, 16'd44281, 16'd55018, 16'd34542, 16'd54094, 16'd22844, 16'd22327, 16'd37815, 16'd52696, 16'd9478, 16'd13754, 16'd17840, 16'd22843, 16'd20975, 16'd56928, 16'd6523, 16'd47094, 16'd59286, 16'd55888, 16'd2305, 16'd20137, 16'd9142, 16'd58412, 16'd10058, 16'd21174});
	test_expansion(128'h2068b6e312475da9f41bf2f3364cc24a, {16'd49107, 16'd5826, 16'd49798, 16'd59738, 16'd19497, 16'd56347, 16'd6430, 16'd29660, 16'd20497, 16'd21314, 16'd63639, 16'd25188, 16'd30377, 16'd7016, 16'd23787, 16'd60065, 16'd33699, 16'd42451, 16'd8036, 16'd63243, 16'd4951, 16'd1193, 16'd25279, 16'd22597, 16'd36615, 16'd15919});
	test_expansion(128'hfc0060eb38f576f5246624ca8214319d, {16'd20090, 16'd25180, 16'd6614, 16'd39518, 16'd31512, 16'd15313, 16'd42992, 16'd43189, 16'd47386, 16'd57731, 16'd8934, 16'd42384, 16'd51914, 16'd17851, 16'd37528, 16'd17047, 16'd63482, 16'd38831, 16'd54356, 16'd55478, 16'd19964, 16'd3271, 16'd22781, 16'd24645, 16'd6045, 16'd18364});
	test_expansion(128'h124ebe37ff3c6228c96693b632c35f28, {16'd47999, 16'd5865, 16'd27521, 16'd42158, 16'd10772, 16'd58239, 16'd61474, 16'd51635, 16'd40777, 16'd13072, 16'd9633, 16'd1081, 16'd12282, 16'd25554, 16'd21334, 16'd18451, 16'd48260, 16'd24520, 16'd2533, 16'd33440, 16'd4535, 16'd35256, 16'd48961, 16'd17116, 16'd47319, 16'd54871});
	test_expansion(128'h891cfd479a8428b9c6b494da70d92b14, {16'd32072, 16'd35434, 16'd36862, 16'd56006, 16'd65472, 16'd33836, 16'd38214, 16'd66, 16'd12285, 16'd8959, 16'd17326, 16'd17112, 16'd65126, 16'd1140, 16'd11662, 16'd2771, 16'd36997, 16'd21299, 16'd32877, 16'd7352, 16'd46219, 16'd56565, 16'd19692, 16'd18796, 16'd48527, 16'd44694});
	test_expansion(128'h98c4b6eee32031c2ddc496bf748ddf84, {16'd50404, 16'd54538, 16'd43589, 16'd45661, 16'd7310, 16'd24591, 16'd57170, 16'd50410, 16'd12206, 16'd21186, 16'd12685, 16'd53507, 16'd41992, 16'd3970, 16'd59355, 16'd1248, 16'd35898, 16'd39406, 16'd22476, 16'd48992, 16'd15720, 16'd55453, 16'd12174, 16'd23606, 16'd26091, 16'd53000});
	test_expansion(128'h44d7e17cbadd86157f0af7c83edb3885, {16'd26980, 16'd25340, 16'd38015, 16'd38371, 16'd17349, 16'd61623, 16'd18397, 16'd10086, 16'd33549, 16'd7700, 16'd47571, 16'd45885, 16'd26006, 16'd19450, 16'd1382, 16'd56529, 16'd63776, 16'd37640, 16'd25461, 16'd5522, 16'd23915, 16'd31758, 16'd21436, 16'd49468, 16'd64691, 16'd17577});
	test_expansion(128'hf5631d6d9111cef83314874a2b1d7e2d, {16'd25440, 16'd57902, 16'd24371, 16'd61388, 16'd15392, 16'd8618, 16'd6085, 16'd54553, 16'd29620, 16'd6305, 16'd36365, 16'd22586, 16'd50236, 16'd1045, 16'd26116, 16'd46189, 16'd29749, 16'd54390, 16'd5375, 16'd31549, 16'd25852, 16'd58028, 16'd4540, 16'd8243, 16'd62732, 16'd11309});
	test_expansion(128'h738af51437ba03435604c76e308f50aa, {16'd50912, 16'd61074, 16'd50347, 16'd23751, 16'd10795, 16'd39520, 16'd32270, 16'd36225, 16'd34725, 16'd15730, 16'd53651, 16'd1959, 16'd40245, 16'd64229, 16'd26730, 16'd2235, 16'd14568, 16'd15619, 16'd10222, 16'd24499, 16'd15223, 16'd5634, 16'd10750, 16'd62351, 16'd61207, 16'd41501});
	test_expansion(128'h384a6da4da116d3f77bb61baa5ec1103, {16'd55384, 16'd19372, 16'd18122, 16'd58624, 16'd2405, 16'd21823, 16'd52253, 16'd53249, 16'd63068, 16'd2822, 16'd7673, 16'd19273, 16'd2429, 16'd42538, 16'd41233, 16'd27574, 16'd9671, 16'd33668, 16'd857, 16'd25531, 16'd47148, 16'd21533, 16'd12542, 16'd18704, 16'd23022, 16'd54196});
	test_expansion(128'h24b79ac284692101261f7ba65bb6e8ea, {16'd20519, 16'd6303, 16'd24765, 16'd20537, 16'd2265, 16'd63932, 16'd51933, 16'd29194, 16'd53291, 16'd31172, 16'd41828, 16'd40822, 16'd39678, 16'd20827, 16'd11967, 16'd13003, 16'd26300, 16'd7980, 16'd8431, 16'd56523, 16'd10151, 16'd58477, 16'd57180, 16'd53423, 16'd43235, 16'd41318});
	test_expansion(128'habb31d8d218f5d8d6c14f7e59a95419b, {16'd4520, 16'd55380, 16'd57128, 16'd17715, 16'd22572, 16'd14638, 16'd54899, 16'd29997, 16'd56396, 16'd4081, 16'd55444, 16'd55399, 16'd50649, 16'd8572, 16'd32802, 16'd48109, 16'd58632, 16'd34996, 16'd11631, 16'd21360, 16'd36449, 16'd54485, 16'd51303, 16'd4635, 16'd7752, 16'd22692});
	test_expansion(128'hde20867c8f1581339e10746220e8e774, {16'd44518, 16'd56134, 16'd60745, 16'd5961, 16'd37336, 16'd6339, 16'd53234, 16'd24538, 16'd33778, 16'd13373, 16'd38704, 16'd33791, 16'd35532, 16'd20240, 16'd38700, 16'd61621, 16'd34212, 16'd29903, 16'd43623, 16'd4902, 16'd50175, 16'd33278, 16'd55779, 16'd56922, 16'd42412, 16'd44151});
	test_expansion(128'hc694af964b75b79abdc1b02538c6d116, {16'd44044, 16'd12652, 16'd42203, 16'd17698, 16'd12423, 16'd18889, 16'd41059, 16'd58290, 16'd3757, 16'd22155, 16'd15731, 16'd64236, 16'd2312, 16'd59459, 16'd61654, 16'd43055, 16'd20332, 16'd55771, 16'd12375, 16'd50626, 16'd63458, 16'd41058, 16'd42613, 16'd19433, 16'd59843, 16'd52671});
	test_expansion(128'h3f64e08ed604bffbacb686d98f4de14f, {16'd11250, 16'd4245, 16'd28004, 16'd35603, 16'd55477, 16'd46352, 16'd27631, 16'd10839, 16'd34846, 16'd24489, 16'd14124, 16'd43233, 16'd35541, 16'd12090, 16'd3823, 16'd65420, 16'd39235, 16'd13557, 16'd39031, 16'd21960, 16'd30132, 16'd518, 16'd25743, 16'd46584, 16'd50749, 16'd6639});
	test_expansion(128'he888c3af1b183b278e62062521824c04, {16'd50335, 16'd50228, 16'd29526, 16'd49671, 16'd63172, 16'd14353, 16'd46825, 16'd1489, 16'd46622, 16'd49337, 16'd62426, 16'd12576, 16'd2834, 16'd36310, 16'd7544, 16'd14811, 16'd62594, 16'd19778, 16'd65503, 16'd253, 16'd58162, 16'd39667, 16'd42814, 16'd57315, 16'd61561, 16'd34970});
	test_expansion(128'h43b85b7b57da279b1a057513b3ab5bac, {16'd41243, 16'd7988, 16'd15537, 16'd32734, 16'd24821, 16'd8053, 16'd43119, 16'd30841, 16'd12218, 16'd32502, 16'd21208, 16'd13900, 16'd12972, 16'd48098, 16'd59991, 16'd14747, 16'd25905, 16'd300, 16'd794, 16'd43250, 16'd49331, 16'd31021, 16'd29443, 16'd26465, 16'd32089, 16'd7227});
	test_expansion(128'he0f0ee681e4903e4755f0b713f3e7343, {16'd19667, 16'd45162, 16'd44720, 16'd15477, 16'd22533, 16'd21862, 16'd58943, 16'd33255, 16'd64477, 16'd18590, 16'd38641, 16'd54983, 16'd18973, 16'd7724, 16'd23302, 16'd14967, 16'd37498, 16'd46618, 16'd30769, 16'd32000, 16'd28486, 16'd62481, 16'd6281, 16'd8134, 16'd49250, 16'd43155});
	test_expansion(128'h82a8e55c83e167e543a9c3e14bf7ca36, {16'd35093, 16'd23782, 16'd24569, 16'd16924, 16'd39891, 16'd24955, 16'd59651, 16'd6800, 16'd21748, 16'd14851, 16'd60965, 16'd35863, 16'd22103, 16'd7511, 16'd37801, 16'd8214, 16'd37101, 16'd35114, 16'd40510, 16'd63878, 16'd38749, 16'd53346, 16'd40471, 16'd58667, 16'd60883, 16'd4852});
	test_expansion(128'h27555d4d85f4fce357af6550be447ded, {16'd25032, 16'd18566, 16'd6163, 16'd59607, 16'd4417, 16'd44982, 16'd55633, 16'd36385, 16'd54243, 16'd17066, 16'd25160, 16'd36085, 16'd54624, 16'd65376, 16'd63169, 16'd53804, 16'd12375, 16'd33108, 16'd61532, 16'd30065, 16'd685, 16'd52541, 16'd58312, 16'd34667, 16'd57051, 16'd24519});


	`endif

    $display("SUCCESS :: FINISH CALLED FROM END OF FILE!");
    $finish;

end


endmodule

