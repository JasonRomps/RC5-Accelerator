
`timescale 1ns / 1ps
module rotl_tb;

logic clk;
logic [15:0] data, shifted, n_shifts;

rotl ROTL(
    .data_i(data),
    .n_i(n_shifts),
    .data_o(shifted)
);

task test_shift(input logic [15:0] test_data, input logic [15:0] n, input logic [15:0] correct);
    data <= test_data;
    n_shifts <= n;
    #2;

    assert(shifted == correct)
        else begin
            $error("Bad Shift: 0x%x << 0x%x: 0x%x, Needed: 0x%x", data, n_shifts, shifted, correct);
            $finish;
        end
endtask


always begin
    clk = 1'b0;
    #1;
    clk = 1'b1;
    #1;
end


initial begin
    $fsdbDumpfile("dump.fsdb");
	$fsdbDumpvars(0, "+all");
    data = 16'b0;

    #2;

	test_shift(16'b1110000011111011, 16'd114, 16'b1000001111101111);
	test_shift(16'b1010010011111111, 16'd22691, 16'b0010011111111101);
	test_shift(16'b0001010100001111, 16'd52790, 16'b0100001111000101);
	test_shift(16'b1001110111011101, 16'd15586, 16'b0111011101110110);
	test_shift(16'b1010010010111111, 16'd62182, 16'b0010111111101001);
	test_shift(16'b0011101011000100, 16'd39083, 16'b0010000111010110);
	test_shift(16'b1001000010100110, 16'd16294, 16'b0010100110100100);
	test_shift(16'b1010111001100000, 16'd48372, 16'b1110011000001010);
	test_shift(16'b0110110100001110, 16'd62653, 16'b1100110110100001);
	test_shift(16'b0110110001100100, 16'd61796, 16'b1100011001000110);
	test_shift(16'b0010111010010111, 16'd37686, 16'b1010010111001011);
	test_shift(16'b1100010010110001, 16'd42599, 16'b0101100011100010);
	test_shift(16'b0110111010010001, 16'd37610, 16'b0100010110111010);
	test_shift(16'b1100110111111100, 16'd21632, 16'b1100110111111100);
	test_shift(16'b0010011100110000, 16'd58587, 16'b1000000100111001);
	test_shift(16'b1100000110101110, 16'd44157, 16'b1101100000110101);
	test_shift(16'b0010011101111001, 16'd47717, 16'b1110111100100100);
	test_shift(16'b0110011101011110, 16'd22029, 16'b1100110011101011);
	test_shift(16'b1111000010011101, 16'd371, 16'b1000010011101111);
	test_shift(16'b1010111110100001, 16'd53350, 16'b1110100001101011);
	test_shift(16'b0111101101001111, 16'd29649, 16'b1111011010011110);
	test_shift(16'b1000110111110001, 16'd32958, 16'b0110001101111100);
	test_shift(16'b0001000001111110, 16'd51509, 16'b0000111111000010);
	test_shift(16'b1110010100000110, 16'd2756, 16'b0101000001101110);
	test_shift(16'b1011001010011100, 16'd14162, 16'b1100101001110010);
	test_shift(16'b1111010010111101, 16'd38467, 16'b1010010111101111);
	test_shift(16'b1110001101110101, 16'd61085, 16'b1011110001101110);
	test_shift(16'b0110010001000000, 16'd15104, 16'b0110010001000000);
	test_shift(16'b0000111111100110, 16'd28919, 16'b1111001100000111);
	test_shift(16'b0011011111111101, 16'd35868, 16'b1101001101111111);
	test_shift(16'b0101100001010101, 16'd8854, 16'b0001010101010110);
	test_shift(16'b1111110110000100, 16'd11052, 16'b0100111111011000);
	test_shift(16'b1011010011011011, 16'd2033, 16'b0110100110110111);
	test_shift(16'b0001100011110100, 16'd49294, 16'b0000011000111101);
	test_shift(16'b1001101100111111, 16'd29756, 16'b1111100110110011);
	test_shift(16'b1100000101110110, 16'd26484, 16'b0001011101101100);
	test_shift(16'b0101000111010110, 16'd23161, 16'b1010110010100011);
	test_shift(16'b1110010010101001, 16'd64541, 16'b0011110010010101);
	test_shift(16'b0100011010111110, 16'd60765, 16'b1100100011010111);
	test_shift(16'b1101111111100000, 16'd55447, 16'b1111000001101111);
	test_shift(16'b0010111000000010, 16'd47327, 16'b0001011100000001);
	test_shift(16'b0001010011100101, 16'd43906, 16'b0101001110010100);
	test_shift(16'b1010101100110110, 16'd46003, 16'b0101100110110101);
	test_shift(16'b0001000001000000, 16'd56763, 16'b0000000010000010);
	test_shift(16'b1111001011100000, 16'd28599, 16'b0111000001111001);
	test_shift(16'b0010001000011011, 16'd30682, 16'b0110110010001000);
	test_shift(16'b1111010001000000, 16'd9754, 16'b0000001111010001);
	test_shift(16'b1100110111000011, 16'd30569, 16'b1000011110011011);
	test_shift(16'b0111011100100011, 16'd57069, 16'b0110111011100100);
	test_shift(16'b1110101010100101, 16'd1797, 16'b0101010010111101);
	test_shift(16'b0110100111000101, 16'd43485, 16'b1010110100111000);
	test_shift(16'b0000110011101101, 16'd53362, 16'b0011001110110100);
	test_shift(16'b1001001000011110, 16'd54007, 16'b0000111101001001);
	test_shift(16'b1011001010001100, 16'd12522, 16'b0011001011001010);
	test_shift(16'b0011001101110000, 16'd28267, 16'b1000000110011011);
	test_shift(16'b0110001010010111, 16'd1437, 16'b1110110001010010);
	test_shift(16'b1111000110000001, 16'd15546, 16'b0000011111000110);
	test_shift(16'b0101100111110010, 16'd52695, 16'b1111100100101100);
	test_shift(16'b1100110101111000, 16'd19485, 16'b0001100110101111);
	test_shift(16'b0101100101010110, 16'd44016, 16'b0101100101010110);
	test_shift(16'b1001100100100000, 16'd18732, 16'b0000100110010010);
	test_shift(16'b0101011110001010, 16'd470, 16'b1110001010010101);
	test_shift(16'b0110011011001111, 16'd18539, 16'b0111101100110110);
	test_shift(16'b1110100101000101, 16'd7321, 16'b1000101111010010);
	test_shift(16'b0100111000111010, 16'd56259, 16'b0111000111010010);
	test_shift(16'b1110011011101000, 16'd25921, 16'b1100110111010001);
	test_shift(16'b1010010111001111, 16'd16544, 16'b1010010111001111);
	test_shift(16'b0100010011110011, 16'd15589, 16'b1001111001101000);
	test_shift(16'b0100001001100010, 16'd51206, 16'b1001100010010000);
	test_shift(16'b1110101001000000, 16'd42375, 16'b0010000001110101);
	test_shift(16'b0100111101110011, 16'd19250, 16'b0011110111001101);
	test_shift(16'b1111101010101101, 16'd7922, 16'b1110101010110111);
	test_shift(16'b1011101111111011, 16'd64527, 16'b1101110111111101);
	test_shift(16'b1111110101100010, 16'd28903, 16'b1011000101111110);
	test_shift(16'b0010101100101110, 16'd9322, 16'b1011100010101100);
	test_shift(16'b0011011111010001, 16'd15485, 16'b0010011011111010);
	test_shift(16'b0000101011011100, 16'd39808, 16'b0000101011011100);
	test_shift(16'b1000111101001100, 16'd46158, 16'b0010001111010011);
	test_shift(16'b0111110101101110, 16'd38168, 16'b0110111001111101);
	test_shift(16'b1011011110001101, 16'd39614, 16'b0110110111100011);
	test_shift(16'b0000111101000101, 16'd55844, 16'b1111010001010000);
	test_shift(16'b0000000110010010, 16'd25382, 16'b0110010010000000);
	test_shift(16'b1011111101010001, 16'd61367, 16'b1010100011011111);
	test_shift(16'b0001011110101011, 16'd33670, 16'b1110101011000101);
	test_shift(16'b0100011000111101, 16'd7521, 16'b1000110001111010);
	test_shift(16'b0111111001100101, 16'd57714, 16'b1111100110010101);
	test_shift(16'b1001010111111010, 16'd9434, 16'b1110101001010111);
	test_shift(16'b1011101000000111, 16'd7484, 16'b0111101110100000);
	test_shift(16'b0110010111111011, 16'd11112, 16'b1111101101100101);
	test_shift(16'b1010000000101011, 16'd9877, 16'b0000010101110100);
	test_shift(16'b1010000011011110, 16'd50514, 16'b1000001101111010);
	test_shift(16'b1011011001101001, 16'd57490, 16'b1101100110100110);
	test_shift(16'b0100000111011101, 16'd58820, 16'b0001110111010100);
	test_shift(16'b1101001111011100, 16'd40798, 16'b0011010011110111);
	test_shift(16'b0001001111110101, 16'd13762, 16'b0100111111010100);
	test_shift(16'b1101110110111111, 16'd37631, 16'b1110111011011111);
	test_shift(16'b0011000111001001, 16'd26632, 16'b1100100100110001);
	test_shift(16'b0110100111100100, 16'd48136, 16'b1110010001101001);
	test_shift(16'b1110110001110100, 16'd13819, 16'b1010011101100011);
	test_shift(16'b0110101110001100, 16'd27900, 16'b1100011010111000);
	test_shift(16'b1010001001111000, 16'd63500, 16'b1000101000100111);
	test_shift(16'b0100111111100111, 16'd26438, 16'b1111100111010011);
	test_shift(16'b1101011011110000, 16'd41270, 16'b1011110000110101);
	test_shift(16'b0011000110110100, 16'd6545, 16'b0110001101101000);
	test_shift(16'b0111111001111000, 16'd38993, 16'b1111110011110000);
	test_shift(16'b1100101010000001, 16'd48387, 16'b0101010000001110);
	test_shift(16'b1011010011111011, 16'd7230, 16'b1110110100111110);
	test_shift(16'b0100000000100011, 16'd54721, 16'b1000000001000110);
	test_shift(16'b0110111111100110, 16'd27807, 16'b0011011111110011);
	test_shift(16'b1111110000100010, 16'd41836, 16'b0010111111000010);
	test_shift(16'b1000101000000001, 16'd31231, 16'b1100010100000000);
	test_shift(16'b1000000100010111, 16'd44078, 16'b1110000001000101);
	test_shift(16'b1110010101101001, 16'd42515, 16'b0010101101001111);
	test_shift(16'b0010011110010100, 16'd1083, 16'b1010000100111100);
	test_shift(16'b1111100010100000, 16'd6012, 16'b0000111110001010);
	test_shift(16'b1110101111011101, 16'd46702, 16'b0111101011110111);
	test_shift(16'b0111001111011111, 16'd11345, 16'b1110011110111110);
	test_shift(16'b1011011011001110, 16'd54728, 16'b1100111010110110);
	test_shift(16'b1000111111100011, 16'd57952, 16'b1000111111100011);
	test_shift(16'b1000001101101000, 16'd33503, 16'b0100000110110100);
	test_shift(16'b0010000101010100, 16'd34921, 16'b1010100001000010);
	test_shift(16'b1101011011101010, 16'd1128, 16'b1110101011010110);
	test_shift(16'b0010010101100111, 16'd17970, 16'b1001010110011100);
	test_shift(16'b0000110011101101, 16'd5369, 16'b1101101000011001);
	test_shift(16'b1111010100100011, 16'd46140, 16'b0011111101010010);
	test_shift(16'b0001110111110101, 16'd53358, 16'b0100011101111101);
	test_shift(16'b0000011100011001, 16'd1237, 16'b1110001100100000);
	test_shift(16'b0011010100011001, 16'd44568, 16'b0001100100110101);
	test_shift(16'b0100011000000010, 16'd6372, 16'b0110000000100100);
	test_shift(16'b1110100000101110, 16'd50030, 16'b1011101000001011);
	test_shift(16'b1101110011101001, 16'd42732, 16'b1001110111001110);
	test_shift(16'b1100101011100111, 16'd25769, 16'b1100111110010101);
	test_shift(16'b1011110010001001, 16'd29183, 16'b1101111001000100);
	test_shift(16'b1111100001101010, 16'd50214, 16'b0001101010111110);
	test_shift(16'b0110011110010111, 16'd8293, 16'b1111001011101100);
	test_shift(16'b0010101001010000, 16'd5172, 16'b1010010100000010);
	test_shift(16'b1100101101101111, 16'd36007, 16'b1011011111100101);
	test_shift(16'b0101010101000011, 16'd37995, 16'b0001101010101010);
	test_shift(16'b0110100111100111, 16'd55893, 16'b0011110011101101);
	test_shift(16'b1000010000011000, 16'd3541, 16'b1000001100010000);
	test_shift(16'b0010000001011001, 16'd61304, 16'b0101100100100000);
	test_shift(16'b1010100100111010, 16'd13411, 16'b0100100111010101);
	test_shift(16'b1000110111110101, 16'd27458, 16'b0011011111010110);
	test_shift(16'b0110010010100000, 16'd14504, 16'b1010000001100100);
	test_shift(16'b1010010010010101, 16'd11159, 16'b0100101011010010);
	test_shift(16'b0110100110111010, 16'd11872, 16'b0110100110111010);
	test_shift(16'b1000010111010010, 16'd10591, 16'b0100001011101001);
	test_shift(16'b1110001000010100, 16'd57925, 16'b0100001010011100);
	test_shift(16'b0110000111010101, 16'd61178, 16'b0101010110000111);
	test_shift(16'b1100110001001111, 16'd34177, 16'b1001100010011111);
	test_shift(16'b1000111000000110, 16'd52614, 16'b1000000110100011);
	test_shift(16'b0101011001111011, 16'd14173, 16'b0110101011001111);
	test_shift(16'b1001011010011010, 16'd21323, 16'b1101010010110100);
	test_shift(16'b0001000110110111, 16'd64430, 16'b1100010001101101);
	test_shift(16'b1010111101100011, 16'd17841, 16'b0101111011000111);
	test_shift(16'b0100000000010100, 16'd59951, 16'b0010000000001010);
	test_shift(16'b1000111011111001, 16'd59060, 16'b1110111110011000);
	test_shift(16'b0111000101010000, 16'd47315, 16'b1000101010000011);
	test_shift(16'b0011100011100010, 16'd12330, 16'b1000100011100011);
	test_shift(16'b0110001010101000, 16'd23985, 16'b1100010101010000);
	test_shift(16'b0001000111111110, 16'd50184, 16'b1111111000010001);
	test_shift(16'b1010011000100000, 16'd33410, 16'b1001100010000010);
	test_shift(16'b1100001000000001, 16'd5081, 16'b0000001110000100);
	test_shift(16'b0000100011111010, 16'd29080, 16'b1111101000001000);
	test_shift(16'b0111000110110111, 16'd1218, 16'b1100011011011101);
	test_shift(16'b0110101011011110, 16'd6423, 16'b0110111100110101);
	test_shift(16'b1110110110100101, 16'd39443, 16'b0110110100101111);
	test_shift(16'b1110110000100010, 16'd19735, 16'b0001000101110110);
	test_shift(16'b1001000101000101, 16'd28109, 16'b1011001000101000);
	test_shift(16'b0001101010010000, 16'd14733, 16'b0000001101010010);
	test_shift(16'b0111111010011101, 16'd15068, 16'b1101011111101001);
	test_shift(16'b0000011100111000, 16'd44984, 16'b0011100000000111);
	test_shift(16'b1111001111111011, 16'd38285, 16'b0111111001111111);
	test_shift(16'b1010111111010111, 16'd62881, 16'b0101111110101111);
	test_shift(16'b1100001001111101, 16'd34078, 16'b0111000010011111);
	test_shift(16'b0110000111110001, 16'd7209, 16'b1110001011000011);
	test_shift(16'b1110111000010011, 16'd2270, 16'b1111101110000100);
	test_shift(16'b1111001000000010, 16'd17600, 16'b1111001000000010);
	test_shift(16'b0101100111100110, 16'd1121, 16'b1011001111001100);
	test_shift(16'b0100000000110111, 16'd41340, 16'b0111010000000011);
	test_shift(16'b0010000110000111, 16'd12145, 16'b0100001100001110);
	test_shift(16'b0000010001110000, 16'd10634, 16'b1100000000010001);
	test_shift(16'b0011001001000010, 16'd54690, 16'b1100100100001000);
	test_shift(16'b0010110110101101, 16'd59586, 16'b1011011010110100);
	test_shift(16'b0011001011110011, 16'd63992, 16'b1111001100110010);
	test_shift(16'b0011000110011101, 16'd48178, 16'b1100011001110100);
	test_shift(16'b0000101011100011, 16'd5604, 16'b1010111000110000);
	test_shift(16'b0101100000011110, 16'd32659, 16'b1100000011110010);
	test_shift(16'b1100110001010110, 16'd8472, 16'b0101011011001100);
	test_shift(16'b1000000001000000, 16'd216, 16'b0100000010000000);
	test_shift(16'b1000010100011110, 16'd45399, 16'b1000111101000010);
	test_shift(16'b1101101001000010, 16'd301, 16'b0101101101001000);
	test_shift(16'b0101010001111000, 16'd64820, 16'b0100011110000101);
	test_shift(16'b0111011110111001, 16'd48787, 16'b1011110111001011);
	test_shift(16'b0110100100011001, 16'd47473, 16'b1101001000110010);
	test_shift(16'b0011100100101001, 16'd1159, 16'b1001010010011100);
	test_shift(16'b1000000110010010, 16'd61695, 16'b0100000011001001);
	test_shift(16'b1100101100010101, 16'd63183, 16'b1110010110001010);
	test_shift(16'b0101001011101000, 16'd28830, 16'b0001010010111010);
	test_shift(16'b1100000100010001, 16'd32946, 16'b0000010001000111);
	test_shift(16'b0011111000011001, 16'd13296, 16'b0011111000011001);
	test_shift(16'b1010111111110000, 16'd18890, 16'b1100001010111111);
	test_shift(16'b0100111000010111, 16'd6421, 16'b1100001011101001);
	test_shift(16'b0100001101011010, 16'd57478, 16'b1101011010010000);
	test_shift(16'b0000011100001110, 16'd13546, 16'b0011100000011100);
	test_shift(16'b1110000010001000, 16'd6018, 16'b1000001000100011);
	test_shift(16'b1110001011111010, 16'd19325, 16'b0101110001011111);
	test_shift(16'b1101110011010110, 16'd33658, 16'b0101101101110011);
	test_shift(16'b0001010100101100, 16'd14050, 16'b0101010010110000);
	test_shift(16'b0100110110110000, 16'd43705, 16'b0110000010011011);
	test_shift(16'b1000000001010101, 16'd25032, 16'b0101010110000000);
	test_shift(16'b1000101011001000, 16'd36627, 16'b0101011001000100);
	test_shift(16'b1001011111001110, 16'd33716, 16'b0111110011101001);
	test_shift(16'b0110011001000000, 16'd13865, 16'b1000000011001100);
	test_shift(16'b1100011011111011, 16'd35334, 16'b1011111011110001);
	test_shift(16'b1011101111010000, 16'd46244, 16'b1011110100001011);
	test_shift(16'b1000111100101110, 16'd7700, 16'b1111001011101000);
	test_shift(16'b1111110101111110, 16'd53842, 16'b1111010111111011);
	test_shift(16'b1101111111110010, 16'd64353, 16'b1011111111100101);
	test_shift(16'b0011111100001100, 16'd44141, 16'b1000011111100001);
	test_shift(16'b0000001000001010, 16'd35979, 16'b0101000000010000);
	test_shift(16'b1101111101110101, 16'd23808, 16'b1101111101110101);
	test_shift(16'b0010111111010000, 16'd16741, 16'b1111101000000101);
	test_shift(16'b0010011101110011, 16'd43474, 16'b1001110111001100);
	test_shift(16'b0110110110101010, 16'd42461, 16'b0100110110110101);
	test_shift(16'b1001101111111101, 16'd41212, 16'b1101100110111111);
	test_shift(16'b1000011001101110, 16'd19161, 16'b1101110100001100);
	test_shift(16'b0010000000000101, 16'd37924, 16'b0000000001010010);
	test_shift(16'b1100100010100001, 16'd29416, 16'b1010000111001000);
	test_shift(16'b0010100000111011, 16'd20804, 16'b1000001110110010);
	test_shift(16'b1101000001001110, 16'd35708, 16'b1110110100000100);
	test_shift(16'b1101110111100001, 16'd52782, 16'b0111011101111000);
	test_shift(16'b1001100100000010, 16'd15443, 16'b1100100000010100);
	test_shift(16'b0010000100110110, 16'd57432, 16'b0011011000100001);
	test_shift(16'b0111001100111110, 16'd15925, 16'b0110011111001110);
	test_shift(16'b1110101000110101, 16'd50106, 16'b1101011110101000);
	test_shift(16'b0010010111011001, 16'd15896, 16'b1101100100100101);
	test_shift(16'b0011001010010110, 16'd46091, 16'b1011000110010100);
	test_shift(16'b0101100011001100, 16'd54256, 16'b0101100011001100);
	test_shift(16'b0110101010011100, 16'd37775, 16'b0011010101001110);
	test_shift(16'b0001110000100001, 16'd50912, 16'b0001110000100001);
	test_shift(16'b1001011101010001, 16'd53785, 16'b1010001100101110);
	test_shift(16'b1011000001100111, 16'd1842, 16'b1100000110011110);
	test_shift(16'b0100010011011100, 16'd32171, 16'b1110001000100110);
	test_shift(16'b1110001100011111, 16'd38311, 16'b1000111111110001);
	test_shift(16'b1101011111110100, 16'd52229, 16'b1111111010011010);
	test_shift(16'b0100010111111011, 16'd33361, 16'b1000101111110110);
	test_shift(16'b1001001000010100, 16'd27579, 16'b1010010010010000);
	test_shift(16'b0010011010101001, 16'd47357, 16'b0010010011010101);
	test_shift(16'b0110010010101101, 16'd13205, 16'b1001010110101100);
	test_shift(16'b0011110010110011, 16'd24562, 16'b1111001011001100);
	test_shift(16'b1110011111110111, 16'd26863, 16'b1111001111111011);
	test_shift(16'b0010100110010000, 16'd9456, 16'b0010100110010000);
	test_shift(16'b0011000110110010, 16'd9202, 16'b1100011011001000);
	test_shift(16'b1011010001011100, 16'd7730, 16'b1101000101110010);
	test_shift(16'b0010110110101001, 16'd874, 16'b1010010010110110);
	test_shift(16'b1010110011101110, 16'd42957, 16'b1101010110011101);
	test_shift(16'b1010010111101100, 16'd21320, 16'b1110110010100101);
	test_shift(16'b0011111111011111, 16'd45786, 16'b0111110011111111);
	test_shift(16'b0110000010011101, 16'd43332, 16'b0000100111010110);
	test_shift(16'b1100000001111111, 16'd53698, 16'b0000000111111111);
	test_shift(16'b0101100010101110, 16'd27454, 16'b1001011000101011);
	test_shift(16'b1001110001010010, 16'd3356, 16'b0010100111000101);
	test_shift(16'b0101111011010101, 16'd54381, 16'b1010101111011010);
	test_shift(16'b0010100100001001, 16'd52714, 16'b0010010010100100);
	test_shift(16'b1011011111100000, 16'd9557, 16'b1111110000010110);
	test_shift(16'b0101000111011100, 16'd60125, 16'b1000101000111011);
	test_shift(16'b0100000110110100, 16'd18669, 16'b1000100000110110);
	test_shift(16'b0101011011011100, 16'd22708, 16'b0110110111000101);
	test_shift(16'b1001101111110010, 16'd56849, 16'b0011011111100101);
	test_shift(16'b0010111010000000, 16'd593, 16'b0101110100000000);
	test_shift(16'b1000110001101001, 16'd48245, 16'b1000110100110001);
	test_shift(16'b1111101000110101, 16'd62916, 16'b1010001101011111);
	test_shift(16'b1001111001001111, 16'd44645, 16'b1100100111110011);
	test_shift(16'b1001110111010010, 16'd20455, 16'b1110100101001110);
	test_shift(16'b0011101110100001, 16'd42607, 16'b1001110111010000);
	test_shift(16'b1010011011111011, 16'd18759, 16'b0111110111010011);
	test_shift(16'b1010011111001100, 16'd41652, 16'b0111110011001010);
	test_shift(16'b1010101100111110, 16'd47093, 16'b0110011111010101);
	test_shift(16'b1110001101010011, 16'd6238, 16'b1111100011010100);
	test_shift(16'b0011101011100010, 16'd51283, 16'b1101011100010001);
	test_shift(16'b0110000101000001, 16'd12994, 16'b1000010100000101);
	test_shift(16'b0011010101101110, 16'd45813, 16'b1010110111000110);
	test_shift(16'b1000000001110110, 16'd44234, 16'b1101101000000001);
	test_shift(16'b0000111101011100, 16'd39543, 16'b1010111000000111);
	test_shift(16'b0011001111011001, 16'd40303, 16'b1001100111101100);
	test_shift(16'b0001110100010101, 16'd30209, 16'b0011101000101010);
	test_shift(16'b0000010011111110, 16'd61291, 16'b1111000000100111);
	test_shift(16'b1000111110010111, 16'd18543, 16'b1100011111001011);
	test_shift(16'b0011110001010111, 16'd62954, 16'b0101110011110001);
	test_shift(16'b0010100010111101, 16'd22566, 16'b0010111101001010);
	test_shift(16'b0011010010001001, 16'd29513, 16'b0001001001101001);
	test_shift(16'b0011000111110001, 16'd53543, 16'b1111100010011000);
	test_shift(16'b1101110111100100, 16'd31304, 16'b1110010011011101);
	test_shift(16'b1100101010101111, 16'd41712, 16'b1100101010101111);
	test_shift(16'b0011000101111010, 16'd61857, 16'b0110001011110100);
	test_shift(16'b0110111000101011, 16'd63507, 16'b0111000101011011);
	test_shift(16'b0001010010110011, 16'd10005, 16'b1001011001100010);
	test_shift(16'b0001001001100111, 16'd22916, 16'b0010011001110001);
	test_shift(16'b0000010100101011, 16'd43393, 16'b0000101001010110);
	test_shift(16'b1110111010001101, 16'd35691, 16'b0110111101110100);
	test_shift(16'b0110110110111010, 16'd36844, 16'b1010011011011011);
	test_shift(16'b0000000000111110, 16'd17605, 16'b0000011111000000);
	test_shift(16'b1111001000001000, 16'd931, 16'b1001000001000111);
	test_shift(16'b1000111100100010, 16'd43420, 16'b0010100011110010);
	test_shift(16'b0000110101000010, 16'd8270, 16'b1000001101010000);
	test_shift(16'b1101000111001111, 16'd22143, 16'b1110100011100111);
	test_shift(16'b0011100101100010, 16'd4441, 16'b1100010001110010);
	test_shift(16'b0010000001010100, 16'd78, 16'b0000100000010101);
	test_shift(16'b1110001100001000, 16'd5720, 16'b0000100011100011);
	test_shift(16'b1110110110111000, 16'd16952, 16'b1011100011101101);
	test_shift(16'b1101010101010101, 16'd10787, 16'b1010101010101110);
	test_shift(16'b0101001011010001, 16'd2565, 16'b0101101000101010);
	test_shift(16'b1100110100000010, 16'd53509, 16'b1010000001011001);
	test_shift(16'b0000100011101011, 16'd31397, 16'b0001110101100001);
	test_shift(16'b0001110010110000, 16'd32427, 16'b1000000011100101);
	test_shift(16'b1000011010001100, 16'd40306, 16'b0001101000110010);
	test_shift(16'b1001000100000101, 16'd428, 16'b0101100100010000);
	test_shift(16'b0010100110100100, 16'd27099, 16'b0010000101001101);
	test_shift(16'b0000100111011001, 16'd20345, 16'b1011001000010011);
	test_shift(16'b0010010000101011, 16'd41264, 16'b0010010000101011);
	test_shift(16'b1111011011111101, 16'd7022, 16'b0111110110111111);
	test_shift(16'b0100000001001011, 16'd8972, 16'b1011010000000100);
	test_shift(16'b0111101101001100, 16'd38229, 16'b0110100110001111);
	test_shift(16'b0010001010101011, 16'd15105, 16'b0100010101010110);
	test_shift(16'b0100100000110110, 16'd1770, 16'b1101100100100000);
	test_shift(16'b1011011011100000, 16'd4507, 16'b0000010110110111);
	test_shift(16'b1100100100100001, 16'd45832, 16'b0010000111001001);
	test_shift(16'b1011000001001100, 16'd42660, 16'b0000010011001011);
	test_shift(16'b0010000110001110, 16'd49635, 16'b0000110001110001);
	test_shift(16'b1101001000011011, 16'd60878, 16'b1111010010000110);
	test_shift(16'b1010110011001110, 16'd8391, 16'b0110011101010110);
	test_shift(16'b0111110111011111, 16'd4262, 16'b0111011111011111);
	test_shift(16'b1000111111110111, 16'd34452, 16'b1111111101111000);
	test_shift(16'b1100011111100110, 16'd44115, 16'b0011111100110110);
	test_shift(16'b1111011010111011, 16'd34187, 16'b1101111110110101);
	test_shift(16'b0111101100010011, 16'd16577, 16'b1111011000100110);
	test_shift(16'b1111001100010010, 16'd60712, 16'b0001001011110011);
	test_shift(16'b1111101001011010, 16'd36987, 16'b1101011111010010);
	test_shift(16'b1100100100011110, 16'd46579, 16'b0100100011110110);
	test_shift(16'b1100110101101100, 16'd4285, 16'b1001100110101101);
	test_shift(16'b1111011100110101, 16'd6612, 16'b0111001101011111);
	test_shift(16'b1001010100011100, 16'd44980, 16'b0101000111001001);
	test_shift(16'b1111000101011110, 16'd20803, 16'b1000101011110111);
	test_shift(16'b1100111010011100, 16'd53676, 16'b1100110011101001);
	test_shift(16'b0110011001000111, 16'd14315, 16'b0011101100110010);
	test_shift(16'b0100110110111001, 16'd45961, 16'b0111001010011011);
	test_shift(16'b0011110001001011, 16'd28851, 16'b1110001001011001);
	test_shift(16'b1111101110001001, 16'd38243, 16'b1101110001001111);
	test_shift(16'b1011111001001010, 16'd12322, 16'b1111100100101010);
	test_shift(16'b0111110000011001, 16'd29958, 16'b0000011001011111);
	test_shift(16'b1011010010001111, 16'd25941, 16'b1001000111110110);
	test_shift(16'b0011000100100100, 16'd31131, 16'b0010000110001001);
	test_shift(16'b0110101100000001, 16'd12181, 16'b0110000000101101);
	test_shift(16'b1011101011110001, 16'd52676, 16'b1010111100011011);
	test_shift(16'b1100001101000111, 16'd17834, 16'b0001111100001101);
	test_shift(16'b1101100001100010, 16'd19530, 16'b1000101101100001);
	test_shift(16'b1001101011010111, 16'd38028, 16'b0111100110101101);
	test_shift(16'b0111001001110110, 16'd7868, 16'b0110011100100111);
	test_shift(16'b1001001100011111, 16'd47303, 16'b1000111111001001);
	test_shift(16'b0100111011100101, 16'd38504, 16'b1110010101001110);
	test_shift(16'b0101011110011101, 16'd33883, 16'b1110101010111100);
	test_shift(16'b0000010010010011, 16'd50988, 16'b0011000001001001);
	test_shift(16'b1110110100011011, 16'd31599, 16'b1111011010001101);
	test_shift(16'b1110101011000101, 16'd57947, 16'b0010111101010110);
	test_shift(16'b0000101001111011, 16'd191, 16'b1000010100111101);
	test_shift(16'b0111110001001110, 16'd29712, 16'b0111110001001110);
	test_shift(16'b0001100110110101, 16'd30302, 16'b0100011001101101);
	test_shift(16'b0101001010110101, 16'd17942, 16'b1010110101010100);
	test_shift(16'b0000101011010000, 16'd11463, 16'b0110100000000101);
	test_shift(16'b0110100001001000, 16'd54272, 16'b0110100001001000);
	test_shift(16'b1011110001010101, 16'd53457, 16'b0111100010101011);
	test_shift(16'b0010110110001011, 16'd10086, 16'b0110001011001011);
	test_shift(16'b0010010000111000, 16'd22492, 16'b1000001001000011);
	test_shift(16'b1001010100100110, 16'd47444, 16'b0101001001101001);
	test_shift(16'b1001110000010000, 16'd41333, 16'b1000001000010011);
	test_shift(16'b1000110101001110, 16'd65366, 16'b0101001110100011);
	test_shift(16'b0000110010001100, 16'd20999, 16'b0100011000000110);
	test_shift(16'b1000101011101101, 16'd3254, 16'b1011101101100010);
	test_shift(16'b1101101110100010, 16'd5320, 16'b1010001011011011);
	test_shift(16'b0100100100000011, 16'd53966, 16'b1101001001000000);
	test_shift(16'b0101100011000100, 16'd47386, 16'b0001000101100011);
	test_shift(16'b1010011110011110, 16'd29848, 16'b1001111010100111);
	test_shift(16'b1101001100000011, 16'd7588, 16'b0011000000111101);
	test_shift(16'b1011101110010111, 16'd6890, 16'b0101111011101110);
	test_shift(16'b0111101001110011, 16'd54959, 16'b1011110100111001);
	test_shift(16'b1100100010000011, 16'd16050, 16'b0010001000001111);
	test_shift(16'b1010001011111110, 16'd57565, 16'b1101010001011111);
	test_shift(16'b1100110000000000, 16'd25926, 16'b0000000000110011);
	test_shift(16'b1001010110100110, 16'd62839, 16'b1101001101001010);
	test_shift(16'b1011110111000010, 16'd47843, 16'b1110111000010101);
	test_shift(16'b0011011111000001, 16'd34617, 16'b1000001001101111);
	test_shift(16'b0000000111001101, 16'd10593, 16'b0000001110011010);
	test_shift(16'b0100111100101110, 16'd26470, 16'b1100101110010011);
	test_shift(16'b0010110000011011, 16'd53195, 16'b1101100101100000);
	test_shift(16'b0010111010110111, 16'd52087, 16'b0101101110010111);
	test_shift(16'b1101100111100010, 16'd41586, 16'b0110011110001011);
	test_shift(16'b1000110011000111, 16'd27488, 16'b1000110011000111);
	test_shift(16'b0011100010011010, 16'd21618, 16'b1110001001101000);
	test_shift(16'b1110101110001010, 16'd19024, 16'b1110101110001010);
	test_shift(16'b1001100100101100, 16'd58201, 16'b0101100100110010);
	test_shift(16'b1101011011011111, 16'd47815, 16'b0110111111101011);
	test_shift(16'b0111110001100101, 16'd54773, 16'b1000110010101111);
	test_shift(16'b1111110011101010, 16'd28585, 16'b1101010111111001);
	test_shift(16'b1010010000111000, 16'd55539, 16'b0010000111000101);
	test_shift(16'b0111010000000000, 16'd58088, 16'b0000000001110100);
	test_shift(16'b1011010100011100, 16'd15672, 16'b0001110010110101);
	test_shift(16'b1111011110111001, 16'd19541, 16'b1111011100111110);
	test_shift(16'b1011010111010110, 16'd30252, 16'b0110101101011101);
	test_shift(16'b1001010010111100, 16'd15580, 16'b1100100101001011);
	test_shift(16'b0111011011100001, 16'd12150, 16'b1011100001011101);
	test_shift(16'b1010111010000010, 16'd23235, 16'b0111010000010101);
	test_shift(16'b1100011011011010, 16'd46596, 16'b0110110110101100);
	test_shift(16'b0111010110101000, 16'd45869, 16'b0000111010110101);
	test_shift(16'b0010011100101110, 16'd22845, 16'b1100010011100101);
	test_shift(16'b0010000101010001, 16'd15299, 16'b0000101010001001);
	test_shift(16'b0000111100101010, 16'd1602, 16'b0011110010101000);
	test_shift(16'b1001101001010011, 16'd63250, 16'b0110100101001110);
	test_shift(16'b0010010011010111, 16'd23260, 16'b0111001001001101);
	test_shift(16'b0111011011101110, 16'd58999, 16'b0111011100111011);
	test_shift(16'b1100100010101000, 16'd51261, 16'b0001100100010101);
	test_shift(16'b0011100101100000, 16'd26647, 16'b1011000000011100);
	test_shift(16'b0101101100110011, 16'd11421, 16'b0110101101100110);
	test_shift(16'b0000100001101000, 16'd25770, 16'b1010000000100001);
	test_shift(16'b0100100111001111, 16'd1830, 16'b0111001111010010);
	test_shift(16'b0101111110001111, 16'd52658, 16'b0111111000111101);
	test_shift(16'b1100000001001110, 16'd55157, 16'b0000100111011000);
	test_shift(16'b1100111101100011, 16'd2085, 16'b1110110001111001);
	test_shift(16'b0011010111110001, 16'd21860, 16'b0101111100010011);
	test_shift(16'b0111000100111101, 16'd46895, 16'b1011100010011110);
	test_shift(16'b1001011101010111, 16'd64102, 16'b1101010111100101);
	test_shift(16'b1110111000011010, 16'd58695, 16'b0000110101110111);
	test_shift(16'b1001110001011011, 16'd31278, 16'b1110011100010110);
	test_shift(16'b0101100111110110, 16'd29267, 16'b1100111110110010);
	test_shift(16'b0010110010111100, 16'd48720, 16'b0010110010111100);
	test_shift(16'b0100001000111111, 16'd53560, 16'b0011111101000010);
	test_shift(16'b1101100110011011, 16'd44984, 16'b1001101111011001);
	test_shift(16'b0010001011100011, 16'd60633, 16'b1100011001000101);
	test_shift(16'b1000011110110111, 16'd36879, 16'b1100001111011011);
	test_shift(16'b1100111011100101, 16'd32328, 16'b1110010111001110);
	test_shift(16'b1110110000111010, 16'd28556, 16'b1010111011000011);
	test_shift(16'b0011101010110110, 16'd1313, 16'b0111010101101100);
	test_shift(16'b0111010111100111, 16'd22961, 16'b1110101111001110);
	test_shift(16'b1001010010001010, 16'd41952, 16'b1001010010001010);
	test_shift(16'b1101001001111111, 16'd6332, 16'b1111110100100111);
	test_shift(16'b1010000011110110, 16'd32432, 16'b1010000011110110);
	test_shift(16'b1101111101011001, 16'd17300, 16'b1111010110011101);
	test_shift(16'b0001111001010010, 16'd38750, 16'b1000011110010100);
	test_shift(16'b1101000100000101, 16'd53222, 16'b0100000101110100);
	test_shift(16'b0000010110010100, 16'd38188, 16'b0100000001011001);
	test_shift(16'b0011101101010011, 16'd59910, 16'b1101010011001110);
	test_shift(16'b0000101101111000, 16'd39481, 16'b1111000000010110);
	test_shift(16'b1001110101011110, 16'd49020, 16'b1110100111010101);
	test_shift(16'b0110110101010000, 16'd33350, 16'b0101010000011011);
	test_shift(16'b1001101101111010, 16'd8244, 16'b1011011110101001);
	test_shift(16'b1010111001001111, 16'd9492, 16'b1110010011111010);
	test_shift(16'b1000000010001001, 16'd57695, 16'b1100000001000100);
	test_shift(16'b1110110010000010, 16'd42299, 16'b0001011101100100);
	test_shift(16'b1101001000010000, 16'd12297, 16'b0010000110100100);
	test_shift(16'b1111011010111100, 16'd15696, 16'b1111011010111100);
	test_shift(16'b0101001110101110, 16'd61037, 16'b1100101001110101);
	test_shift(16'b1011110110101000, 16'd6512, 16'b1011110110101000);
	test_shift(16'b0011011000010101, 16'd11820, 16'b0101001101100001);
	test_shift(16'b0010011100000100, 16'd54961, 16'b0100111000001000);
	test_shift(16'b0100001110010010, 16'd24898, 16'b0000111001001001);
	test_shift(16'b0000101001000011, 16'd8655, 16'b1000010100100001);
	test_shift(16'b1100101100110000, 16'd58287, 16'b0110010110011000);
	test_shift(16'b1001001011101010, 16'd35171, 16'b1001011101010100);
	test_shift(16'b1011011100000000, 16'd65345, 16'b0110111000000001);
	test_shift(16'b0010001010010001, 16'd38728, 16'b1001000100100010);
	test_shift(16'b1100001101001001, 16'd51395, 16'b0001101001001110);
	test_shift(16'b1100100000001101, 16'd27108, 16'b1000000011011100);
	test_shift(16'b0001000111110001, 16'd26094, 16'b0100010001111100);
	test_shift(16'b0010000010010000, 16'd63003, 16'b1000000100000100);
	test_shift(16'b0111001100100100, 16'd54605, 16'b1000111001100100);
	test_shift(16'b1110100111000010, 16'd32691, 16'b0100111000010111);
	test_shift(16'b0101001101101101, 16'd63217, 16'b1010011011011010);
	test_shift(16'b0110001100010100, 16'd57693, 16'b1000110001100010);
	test_shift(16'b1111111011010000, 16'd50002, 16'b1111101101000011);
	test_shift(16'b0001011010110001, 16'd52266, 16'b1100010001011010);
	test_shift(16'b1000111100111000, 16'd9668, 16'b1111001110001000);
	test_shift(16'b0001101001110001, 16'd62268, 16'b0001000110100111);
	test_shift(16'b1001000111000011, 16'd45313, 16'b0010001110000111);
	test_shift(16'b1111100110111000, 16'd60551, 16'b1101110001111100);
	test_shift(16'b1001001001100001, 16'd43081, 16'b1100001100100100);
	test_shift(16'b1111110010111010, 16'd55183, 16'b0111111001011101);
	test_shift(16'b0011111100001100, 16'd16656, 16'b0011111100001100);
	test_shift(16'b0010001100101010, 16'd26316, 16'b1010001000110010);
	test_shift(16'b1100101110010110, 16'd23851, 16'b1011011001011100);
	test_shift(16'b1001000111100010, 16'd57649, 16'b0010001111000101);
	test_shift(16'b1101010100101111, 16'd63630, 16'b1111010101001011);
	test_shift(16'b0101001011110111, 16'd45742, 16'b1101010010111101);
	test_shift(16'b0010011101001000, 16'd43693, 16'b0000010011101001);
	test_shift(16'b1111101101010110, 16'd18141, 16'b1101111101101010);
	test_shift(16'b0010000100001110, 16'd19642, 16'b0011100010000100);
	test_shift(16'b0101110010100100, 16'd48560, 16'b0101110010100100);
	test_shift(16'b0100100100111111, 16'd44116, 16'b1001001111110100);
	test_shift(16'b0000000011000110, 16'd33747, 16'b0000011000110000);
	test_shift(16'b1010111111000100, 16'd52890, 16'b0001001010111111);
	test_shift(16'b0101111100111110, 16'd59345, 16'b1011111001111100);
	test_shift(16'b1001010100101111, 16'd29485, 16'b1111001010100101);
	test_shift(16'b0001101000100101, 16'd14702, 16'b0100011010001001);
	test_shift(16'b0110111001101101, 16'd44799, 16'b1011011100110110);
	test_shift(16'b1000011100110001, 16'd15291, 16'b1000110000111001);
	test_shift(16'b0100111000010110, 16'd14022, 16'b1000010110010011);
	test_shift(16'b0000010100000000, 16'd59666, 16'b0001010000000000);
	test_shift(16'b1000100110000011, 16'd51479, 16'b1100000111000100);
	test_shift(16'b0111010010101000, 16'd45205, 16'b1001010100001110);
	test_shift(16'b0101100111100001, 16'd63055, 16'b1010110011110000);
	test_shift(16'b0100011101101111, 16'd51806, 16'b1101000111011011);
	test_shift(16'b1110110010000011, 16'd7065, 16'b0000011111011001);
	test_shift(16'b1100100000110000, 16'd27007, 16'b0110010000011000);
	test_shift(16'b1111001101100010, 16'd8971, 16'b0001011110011011);
	test_shift(16'b0010101110100100, 16'd17087, 16'b0001010111010010);
	test_shift(16'b1001011001010111, 16'd14639, 16'b1100101100101011);
	test_shift(16'b1011101001111111, 16'd28115, 16'b1101001111111101);
	test_shift(16'b1000100110010110, 16'd7648, 16'b1000100110010110);
	test_shift(16'b1101001010101100, 16'd31200, 16'b1101001010101100);
	test_shift(16'b1011110101101000, 16'd54595, 16'b1110101101000101);
	test_shift(16'b1111010101001101, 16'd64467, 16'b1010101001101111);
	test_shift(16'b0111111011110010, 16'd56475, 16'b1001001111110111);
	test_shift(16'b0111110100010100, 16'd27713, 16'b1111101000101000);
	test_shift(16'b1101001010110001, 16'd28137, 16'b0110001110100101);
	test_shift(16'b0101110000010010, 16'd37341, 16'b0100101110000010);
	test_shift(16'b0001111001010111, 16'd37835, 16'b1011100011110010);
	test_shift(16'b0000011001110110, 16'd27311, 16'b0000001100111011);
	test_shift(16'b0111010001100001, 16'd40318, 16'b0101110100011000);
	test_shift(16'b0100011100000001, 16'd56836, 16'b0111000000010100);
	test_shift(16'b1111001110110001, 16'd53757, 16'b0011111001110110);
	test_shift(16'b1011101100100100, 16'd2125, 16'b1001011101100100);
	test_shift(16'b0111100101011110, 16'd24452, 16'b1001010111100111);
	test_shift(16'b0000000001010000, 16'd40473, 16'b1010000000000000);
	test_shift(16'b0001101100001110, 16'd44244, 16'b1011000011100001);
	test_shift(16'b1110011011011111, 16'd2705, 16'b1100110110111111);
	test_shift(16'b1100101101010111, 16'd40508, 16'b0111110010110101);
	test_shift(16'b1000110011010011, 16'd2215, 16'b0110100111000110);
	test_shift(16'b1111000001100100, 16'd24571, 16'b0010011110000011);
	test_shift(16'b1011100010000011, 16'd22095, 16'b1101110001000001);
	test_shift(16'b0010010110110001, 16'd57403, 16'b1000100100101101);
	test_shift(16'b1001000101110011, 16'd23686, 16'b0101110011100100);
	test_shift(16'b0001000111011010, 16'd61539, 16'b1000111011010000);
	test_shift(16'b0100111011101101, 16'd26740, 16'b1110111011010100);
	test_shift(16'b1010001001101111, 16'd13485, 16'b1111010001001101);
	test_shift(16'b0000101011100111, 16'd4977, 16'b0001010111001110);
	test_shift(16'b0000101010110100, 16'd42977, 16'b0001010101101000);
	test_shift(16'b0001001110101110, 16'd56661, 16'b0111010111000010);
	test_shift(16'b1001011000110101, 16'd9206, 16'b1000110101100101);
	test_shift(16'b0000011010110101, 16'd64833, 16'b0000110101101010);
	test_shift(16'b1011101000110100, 16'd27800, 16'b0011010010111010);
	test_shift(16'b1110101011100100, 16'd55137, 16'b1101010111001001);
	test_shift(16'b0001011000100011, 16'd21074, 16'b0101100010001100);
	test_shift(16'b0001011100011010, 16'd18058, 16'b0110100001011100);
	test_shift(16'b0111110000010001, 16'd56324, 16'b1100000100010111);
	test_shift(16'b1001000110101111, 16'd44524, 16'b1111100100011010);
	test_shift(16'b1011101010111111, 16'd31525, 16'b0101011111110111);
	test_shift(16'b0111111110010000, 16'd65391, 16'b0011111111001000);
	test_shift(16'b1011000000101010, 16'd34021, 16'b0000010101010110);
	test_shift(16'b0011101010100100, 16'd44914, 16'b1110101010010000);
	test_shift(16'b1010010010110101, 16'd26821, 16'b1001011010110100);
	test_shift(16'b0011011011000110, 16'd40031, 16'b0001101101100011);
	test_shift(16'b0111101101101111, 16'd581, 16'b0110110111101111);
	test_shift(16'b1110011001000010, 16'd28280, 16'b0100001011100110);
	test_shift(16'b0110011011001000, 16'd9500, 16'b1000011001101100);
	test_shift(16'b0111000000000011, 16'd32555, 16'b0001101110000000);
	test_shift(16'b0011110011110110, 16'd10185, 16'b1110110001111001);
	test_shift(16'b1010001000010101, 16'd3614, 16'b0110100010000101);
	test_shift(16'b1111101000010011, 16'd63530, 16'b0100111111101000);
	test_shift(16'b1100111101000001, 16'd12129, 16'b1001111010000011);
	test_shift(16'b0011011101100001, 16'd38130, 16'b1101110110000100);
	test_shift(16'b1011111110100101, 16'd25433, 16'b0100101101111111);
	test_shift(16'b1000110100110010, 16'd53737, 16'b0110010100011010);
	test_shift(16'b1010111001110111, 16'd40537, 16'b1110111101011100);
	test_shift(16'b1111101001101001, 16'd64522, 16'b1010011111101001);
	test_shift(16'b0110011101100101, 16'd36595, 16'b0011101100101011);
	test_shift(16'b1101110011001001, 16'd28777, 16'b1001001110111001);
	test_shift(16'b1100010000110111, 16'd43639, 16'b0001101111100010);
	test_shift(16'b1111110110101010, 16'd27018, 16'b1010101111110110);
	test_shift(16'b1011001010001101, 16'd39788, 16'b1101101100101000);
	test_shift(16'b0011010000110101, 16'd54076, 16'b0101001101000011);
	test_shift(16'b1101001110111100, 16'd57805, 16'b1001101001110111);
	test_shift(16'b0000100010001010, 16'd52818, 16'b0010001000101000);
	test_shift(16'b1110110000010001, 16'd9994, 16'b0100011110110000);
	test_shift(16'b0111010101110011, 16'd20594, 16'b1101010111001101);
	test_shift(16'b0111011011011110, 16'd521, 16'b1011110011101101);
	test_shift(16'b0110111100101111, 16'd34511, 16'b1011011110010111);
	test_shift(16'b0110110111011110, 16'd47141, 16'b1011101111001101);
	test_shift(16'b0111000011101010, 16'd48087, 16'b0111010100111000);
	test_shift(16'b0001000011101110, 16'd16958, 16'b1000010000111011);
	test_shift(16'b1100001111011100, 16'd512, 16'b1100001111011100);
	test_shift(16'b0001001000100001, 16'd14530, 16'b0100100010000100);
	test_shift(16'b1000101101001110, 16'd60857, 16'b1001110100010110);
	test_shift(16'b1100001000011010, 16'd56604, 16'b1010110000100001);
	test_shift(16'b0001110011000100, 16'd22645, 16'b1001100010000011);
	test_shift(16'b0111010110001110, 16'd62359, 16'b1100011100111010);
	test_shift(16'b0010001010110010, 16'd35945, 16'b0110010001000101);
	test_shift(16'b0110111111001111, 16'd31866, 16'b0011110110111111);
	test_shift(16'b1111101001011111, 16'd38184, 16'b0101111111111010);
	test_shift(16'b0101001010010000, 16'd25959, 16'b0100100000101001);
	test_shift(16'b0111111000100011, 16'd37021, 16'b0110111111000100);
	test_shift(16'b0101011011101011, 16'd23314, 16'b0101101110101101);
	test_shift(16'b0010111110110011, 16'd63746, 16'b1011111011001100);
	test_shift(16'b0100110111110011, 16'd61874, 16'b0011011111001101);
	test_shift(16'b1001010000010011, 16'd13626, 16'b0100111001010000);
	test_shift(16'b0001111110001011, 16'd8219, 16'b0101100011111100);
	test_shift(16'b1001100011001011, 16'd61382, 16'b0011001011100110);
	test_shift(16'b0011000001100101, 16'd64960, 16'b0011000001100101);
	test_shift(16'b0001100101010011, 16'd10634, 16'b0100110001100101);
	test_shift(16'b1001010101110100, 16'd34331, 16'b1010010010101011);
	test_shift(16'b0011010100110011, 16'd23779, 16'b1010100110011001);
	test_shift(16'b1011000010100001, 16'd1963, 16'b0000110110000101);
	test_shift(16'b0100000010010111, 16'd61882, 16'b0101110100000010);
	test_shift(16'b1111110111110110, 16'd37320, 16'b1111011011111101);
	test_shift(16'b0101010001000111, 16'd43297, 16'b1010100010001110);
	test_shift(16'b0111100001000011, 16'd1971, 16'b1100001000011011);
	test_shift(16'b0011011010010000, 16'd64210, 16'b1101101001000000);
	test_shift(16'b0011001001110000, 16'd14310, 16'b1001110000001100);
	test_shift(16'b1101010101000111, 16'd63922, 16'b0101010100011111);
	test_shift(16'b1010101000000011, 16'd18258, 16'b1010100000001110);
	test_shift(16'b0110010000001011, 16'd65445, 16'b1000000101101100);
	test_shift(16'b0110001111111110, 16'd1608, 16'b1111111001100011);
	test_shift(16'b1101001011010010, 16'd33652, 16'b0010110100101101);
	test_shift(16'b0111110100011011, 16'd27193, 16'b0011011011111010);
	test_shift(16'b0110000010100000, 16'd63898, 16'b1000000110000010);
	test_shift(16'b0011111111111010, 16'd21549, 16'b0100011111111111);
	test_shift(16'b0101010011010111, 16'd51364, 16'b0100110101110101);
	test_shift(16'b1010110110110011, 16'd8975, 16'b1101011011011001);
	test_shift(16'b0111111011001000, 16'd1903, 16'b0011111101100100);
	test_shift(16'b1101010110011010, 16'd5177, 16'b0011010110101011);
	test_shift(16'b1100010101101010, 16'd12117, 16'b1010110101011000);
	test_shift(16'b0111101001010110, 16'd4768, 16'b0111101001010110);
	test_shift(16'b0101011111111001, 16'd30828, 16'b1001010101111111);
	test_shift(16'b1000000110101111, 16'd49065, 16'b0101111100000011);
	test_shift(16'b0111011100010011, 16'd22038, 16'b1100010011011101);
	test_shift(16'b0001011100110011, 16'd34737, 16'b0010111001100110);
	test_shift(16'b1010000101010001, 16'd44421, 16'b0010101000110100);
	test_shift(16'b0001001100011011, 16'd61922, 16'b0100110001101100);
	test_shift(16'b0111111101001001, 16'd2449, 16'b1111111010010010);
	test_shift(16'b1100101010000101, 16'd26238, 16'b0111001010100001);
	test_shift(16'b1100000010101000, 16'd28065, 16'b1000000101010001);
	test_shift(16'b0100000110111101, 16'd9715, 16'b0000110111101010);
	test_shift(16'b1111010001101011, 16'd55919, 16'b1111101000110101);
	test_shift(16'b0100100111000101, 16'd33199, 16'b1010010011100010);
	test_shift(16'b1100100001001111, 16'd13657, 16'b1001111110010000);
	test_shift(16'b1010110001001110, 16'd10172, 16'b1110101011000100);
	test_shift(16'b0000111011101101, 16'd35981, 16'b1010000111011101);
	test_shift(16'b0110100010110111, 16'd50232, 16'b1011011101101000);
	test_shift(16'b0110001101101110, 16'd63104, 16'b0110001101101110);
	test_shift(16'b1010001000101111, 16'd40834, 16'b1000100010111110);
	test_shift(16'b0101110001101010, 16'd62416, 16'b0101110001101010);
	test_shift(16'b1001101111000110, 16'd18370, 16'b0110111100011010);
	test_shift(16'b1101010011100110, 16'd18234, 16'b1001101101010011);
	test_shift(16'b0010000011000101, 16'd10452, 16'b0000110001010010);
	test_shift(16'b0100001101111110, 16'd26211, 16'b0001101111110010);
	test_shift(16'b1111011000101110, 16'd17470, 16'b1011110110001011);
	test_shift(16'b1100010000110001, 16'd9560, 16'b0011000111000100);
	test_shift(16'b0101011101101100, 16'd14324, 16'b0111011011000101);
	test_shift(16'b0011000111001111, 16'd9855, 16'b1001100011100111);
	test_shift(16'b0110010010110110, 16'd40410, 16'b1101100110010010);
	test_shift(16'b1110100000100101, 16'd15412, 16'b1000001001011110);
	test_shift(16'b0010000000010000, 16'd36184, 16'b0001000000100000);
	test_shift(16'b1011001000001001, 16'd27756, 16'b1001101100100000);
	test_shift(16'b1110110001110001, 16'd15824, 16'b1110110001110001);
	test_shift(16'b1001101100001110, 16'd2130, 16'b0110110000111010);
	test_shift(16'b0101110101111111, 16'd49827, 16'b1110101111111010);
	test_shift(16'b1010010111110000, 16'd50395, 16'b1000010100101111);
	test_shift(16'b0000010110101001, 16'd6170, 16'b1010010000010110);
	test_shift(16'b1110001110000110, 16'd40174, 16'b1011100011100001);
	test_shift(16'b0011100000011010, 16'd31756, 16'b1010001110000001);
	test_shift(16'b1111011100001111, 16'd30196, 16'b0111000011111111);
	test_shift(16'b1010101001100110, 16'd39366, 16'b1001100110101010);
	test_shift(16'b1101101001000000, 16'd59168, 16'b1101101001000000);
	test_shift(16'b0100110001001101, 16'd3045, 16'b1000100110101001);
	test_shift(16'b1111000110111101, 16'd53749, 16'b0011011110111110);
	test_shift(16'b0000010010110101, 16'd13337, 16'b0110101000001001);
	test_shift(16'b1001010001000101, 16'd57183, 16'b1100101000100010);
	test_shift(16'b1000110010110111, 16'd35023, 16'b1100011001011011);
	test_shift(16'b0111101111110011, 16'd15679, 16'b1011110111111001);
	test_shift(16'b1010101001001010, 16'd15711, 16'b0101010100100101);
	test_shift(16'b0100011100011100, 16'd58455, 16'b1000111000100011);
	test_shift(16'b1100101000101100, 16'd15366, 16'b1000101100110010);
	test_shift(16'b0001111111001000, 16'd48386, 16'b0111111100100000);
	test_shift(16'b1000110000100000, 16'd60924, 16'b0000100011000010);
	test_shift(16'b1011110011101101, 16'd22307, 16'b1110011101101101);
	test_shift(16'b1000011111000110, 16'd29916, 16'b0110100001111100);
	test_shift(16'b0101011001010000, 16'd46724, 16'b0110010100000101);
	test_shift(16'b0001101110101000, 16'd32940, 16'b1000000110111010);
	test_shift(16'b0110011010000101, 16'd43953, 16'b1100110100001010);
	test_shift(16'b1110101001011001, 16'd21624, 16'b0101100111101010);
	test_shift(16'b1010000100010110, 16'd51859, 16'b0000100010110101);
	test_shift(16'b1010000000000110, 16'd8144, 16'b1010000000000110);
	test_shift(16'b1111000111000111, 16'd30223, 16'b1111100011100011);
	test_shift(16'b1101000000101110, 16'd62178, 16'b0100000010111011);
	test_shift(16'b0011100010011001, 16'd241, 16'b0111000100110010);
	test_shift(16'b0110001100000011, 16'd40746, 16'b0000110110001100);
	test_shift(16'b1000100010010101, 16'd43941, 16'b0001001010110001);
	test_shift(16'b1011111011111111, 16'd35509, 16'b1101111111110111);
	test_shift(16'b1001011000000000, 16'd31137, 16'b0010110000000001);
	test_shift(16'b0010001011101010, 16'd52910, 16'b1000100010111010);
	test_shift(16'b1111010001101000, 16'd31573, 16'b1000110100011110);
	test_shift(16'b1001110011101001, 16'd20131, 16'b1110011101001100);
	test_shift(16'b0101000001010010, 16'd12303, 16'b0010100000101001);
	test_shift(16'b0101011001011010, 16'd58709, 16'b1100101101001010);
	test_shift(16'b1001110111001111, 16'd18343, 16'b1110011111001110);
	test_shift(16'b1001011100000100, 16'd39919, 16'b0100101110000010);
	test_shift(16'b0100111000101110, 16'd47643, 16'b0111001001110001);
	test_shift(16'b1111110100010111, 16'd3693, 16'b1111111110100010);
	test_shift(16'b1011111001011001, 16'd56426, 16'b0110011011111001);
	test_shift(16'b1111100111100110, 16'd45993, 16'b1100110111110011);
	test_shift(16'b1011001001011110, 16'd26298, 16'b0111101011001001);
	test_shift(16'b1100000000001011, 16'd49872, 16'b1100000000001011);
	test_shift(16'b0101010010011110, 16'd22160, 16'b0101010010011110);
	test_shift(16'b1000101101001101, 16'd3742, 16'b0110001011010011);
	test_shift(16'b0100010011001110, 16'd29721, 16'b1001110010001001);
	test_shift(16'b1111100010010000, 16'd41516, 16'b0000111110001001);
	test_shift(16'b1111011010000000, 16'd36098, 16'b1101101000000011);
	test_shift(16'b1000001011100101, 16'd9304, 16'b1110010110000010);
	test_shift(16'b0101010100100011, 16'd54658, 16'b0101010010001101);
	test_shift(16'b0100000101111010, 16'd62424, 16'b0111101001000001);
	test_shift(16'b0010000101100110, 16'd25115, 16'b0011000100001011);
	test_shift(16'b0001100110010011, 16'd7620, 16'b1001100100110001);
	test_shift(16'b0010111100011100, 16'd55891, 16'b0111100011100001);
	test_shift(16'b0001011000100000, 16'd11552, 16'b0001011000100000);
	test_shift(16'b1001100010101101, 16'd30756, 16'b1000101011011001);
	test_shift(16'b0010000010001011, 16'd48609, 16'b0100000100010110);
	test_shift(16'b0001010101111111, 16'd16994, 16'b0101010111111100);
	test_shift(16'b1001011010011010, 16'd55746, 16'b0101101001101010);
	test_shift(16'b1111111000011111, 16'd4950, 16'b1000011111111111);
	test_shift(16'b1110000110111111, 16'd23170, 16'b1000011011111111);
	test_shift(16'b0010000111101010, 16'd22597, 16'b0011110101000100);
	test_shift(16'b0110001101000001, 16'd30786, 16'b1000110100000101);
	test_shift(16'b0110000101010001, 16'd28363, 16'b1000101100001010);
	test_shift(16'b1001000000000101, 16'd56794, 16'b0001011001000000);
	test_shift(16'b0100011111000110, 16'd53806, 16'b1001000111110001);
	test_shift(16'b1011000100011000, 16'd45064, 16'b0001100010110001);
	test_shift(16'b0101010010011010, 16'd10868, 16'b0100100110100101);
	test_shift(16'b1101010101001100, 16'd9938, 16'b0101010100110011);
	test_shift(16'b0010010100110010, 16'd54408, 16'b0011001000100101);
	test_shift(16'b0001110010100100, 16'd1636, 16'b1100101001000001);
	test_shift(16'b1011101100011101, 16'd45155, 16'b1101100011101101);
	test_shift(16'b1010110011011010, 16'd49748, 16'b1100110110101010);
	test_shift(16'b0110011100110010, 16'd18891, 16'b1001001100111001);
	test_shift(16'b0100011101000011, 16'd28437, 16'b1110100001101000);
	test_shift(16'b1110101011010011, 16'd16082, 16'b1010101101001111);
	test_shift(16'b1101110000010010, 16'd3861, 16'b1000001001011011);
	test_shift(16'b1101011010001011, 16'd29521, 16'b1010110100010111);
	test_shift(16'b0100001111010011, 16'd720, 16'b0100001111010011);
	test_shift(16'b0101000001011011, 16'd34714, 16'b0110110101000001);
	test_shift(16'b0101110000100010, 16'd25631, 16'b0010111000010001);
	test_shift(16'b1101101110101000, 16'd57852, 16'b1000110110111010);
	test_shift(16'b0100001101001011, 16'd58329, 16'b1001011010000110);
	test_shift(16'b0100010111000110, 16'd45956, 16'b0101110001100100);
	test_shift(16'b0011000111111001, 16'd22035, 16'b1000111111001001);
	test_shift(16'b0101111010101000, 16'd47848, 16'b1010100001011110);
	test_shift(16'b1000001100001000, 16'd65368, 16'b0000100010000011);
	test_shift(16'b1000110011101111, 16'd36149, 16'b1001110111110001);
	test_shift(16'b0000011100010110, 16'd42808, 16'b0001011000000111);
	test_shift(16'b0110010110010111, 16'd57209, 16'b0010111011001011);
	test_shift(16'b0000110010000000, 16'd55103, 16'b0000011001000000);
	test_shift(16'b1111011000001100, 16'd933, 16'b1100000110011110);
	test_shift(16'b1011110010111001, 16'd37876, 16'b1100101110011011);
	test_shift(16'b1111110100101000, 16'd54024, 16'b0010100011111101);
	test_shift(16'b1101001010101110, 16'd27868, 16'b1110110100101010);
	test_shift(16'b1110101110001001, 16'd50284, 16'b1001111010111000);
	test_shift(16'b1000000001100010, 16'd39781, 16'b0000110001010000);
	test_shift(16'b1001011111111001, 16'd5757, 16'b0011001011111111);
	test_shift(16'b0001000001001101, 16'd48829, 16'b1010001000001001);
	test_shift(16'b0011011111001100, 16'd53200, 16'b0011011111001100);
	test_shift(16'b0111000100111111, 16'd13133, 16'b1110111000100111);
	test_shift(16'b0100111011011110, 16'd47418, 16'b0111100100111011);
	test_shift(16'b1011101101000111, 16'd12699, 16'b0011110111011010);
	test_shift(16'b0011000111010110, 16'd12509, 16'b1100011000111010);
	test_shift(16'b1111110011010101, 16'd41850, 16'b0101011111110011);
	test_shift(16'b0100000011000110, 16'd60505, 16'b1000110010000001);
	test_shift(16'b0111111101000111, 16'd25614, 16'b1101111111010001);
	test_shift(16'b1101111110101100, 16'd34710, 16'b1110101100110111);
	test_shift(16'b1001110101010111, 16'd15038, 16'b1110011101010101);
	test_shift(16'b0100000111000011, 16'd708, 16'b0001110000110100);
	test_shift(16'b0011110111101110, 16'd26570, 16'b1011100011110111);
	test_shift(16'b0100010110110010, 16'd22642, 16'b0001011011001001);
	test_shift(16'b1001101000001011, 16'd22643, 16'b1101000001011100);
	test_shift(16'b0011100000011010, 16'd46414, 16'b1000111000000110);
	test_shift(16'b0010101110110001, 16'd46264, 16'b1011000100101011);
	test_shift(16'b1011010000100001, 16'd13703, 16'b0001000011011010);
	test_shift(16'b0110010100011010, 16'd26851, 16'b0010100011010011);
	test_shift(16'b1110000101100000, 16'd41892, 16'b0001011000001110);
	test_shift(16'b1110001100011100, 16'd14945, 16'b1100011000111001);
	test_shift(16'b0000101000011001, 16'd13059, 16'b0101000011001000);
	test_shift(16'b0111001100000110, 16'd38150, 16'b1100000110011100);
	test_shift(16'b0100001110011000, 16'd21284, 16'b0011100110000100);
	test_shift(16'b0110101101110101, 16'd1529, 16'b1110101011010110);
	test_shift(16'b0100110001101101, 16'd64598, 16'b0001101101010011);
	test_shift(16'b0000011101000111, 16'd7481, 16'b1000111000001110);
	test_shift(16'b0010010001001001, 16'd24699, 16'b0100100100100010);
	test_shift(16'b1010000010110001, 16'd33702, 16'b0010110001101000);
	test_shift(16'b1011110010101001, 16'd29820, 16'b1001101111001010);
	test_shift(16'b1011110011100011, 16'd45803, 16'b0001110111100111);
	test_shift(16'b0001000111011010, 16'd7478, 16'b0111011010000100);
	test_shift(16'b1111000010011010, 16'd17779, 16'b1000010011010111);
	test_shift(16'b0000001001010010, 16'd5751, 16'b0010100100000001);
	test_shift(16'b1001001111101111, 16'd30966, 16'b1111101111100100);
	test_shift(16'b0001011100111010, 16'd25759, 16'b0000101110011101);
	test_shift(16'b1011111001110001, 16'd48092, 16'b0001101111100111);
	test_shift(16'b1110011011000000, 16'd41590, 16'b1011000000111001);
	test_shift(16'b1000110000001100, 16'd61606, 16'b0000001100100011);
	test_shift(16'b0000000111100011, 16'd41909, 16'b0011110001100000);
	test_shift(16'b1010110000111110, 16'd35743, 16'b0101011000011111);
	test_shift(16'b0000110110010101, 16'd37665, 16'b0001101100101010);
	test_shift(16'b0000100000001110, 16'd61950, 16'b1000001000000011);
	test_shift(16'b1100100010101110, 16'd32781, 16'b1101100100010101);
	test_shift(16'b0011110111011010, 16'd48978, 16'b1111011101101000);
	test_shift(16'b1011010111011011, 16'd19223, 16'b1110110111011010);
	test_shift(16'b0001000101011100, 16'd56563, 16'b1000101011100000);
	test_shift(16'b0001011000100010, 16'd33920, 16'b0001011000100010);
	test_shift(16'b1101100100011101, 16'd36888, 16'b0001110111011001);
	test_shift(16'b0101100101110001, 16'd13143, 16'b1011100010101100);
	test_shift(16'b1110100110010111, 16'd2831, 16'b1111010011001011);
	test_shift(16'b0111100101000110, 16'd60932, 16'b1001010001100111);
	test_shift(16'b1100000111111010, 16'd20144, 16'b1100000111111010);
	test_shift(16'b1001011111100111, 16'd53743, 16'b1100101111110011);
	test_shift(16'b1110101000101011, 16'd247, 16'b0001010111110101);
	test_shift(16'b0000101010001011, 16'd19768, 16'b1000101100001010);
	test_shift(16'b0010010001000000, 16'd46123, 16'b0000000100100010);
	test_shift(16'b0010111101011100, 16'd54794, 16'b0111000010111101);
	test_shift(16'b1111100001100111, 16'd32539, 16'b0011111111000011);
	test_shift(16'b1001001111110100, 16'd18807, 16'b1111101001001001);
	test_shift(16'b0000101110101011, 16'd47367, 16'b1101010110000101);
	test_shift(16'b0011100000110000, 16'd34159, 16'b0001110000011000);
	test_shift(16'b0000001101111011, 16'd45767, 16'b1011110110000001);
	test_shift(16'b1000011000100110, 16'd9411, 16'b0011000100110100);
	test_shift(16'b0001010000011000, 16'd25002, 16'b0110000001010000);
	test_shift(16'b0010100110101101, 16'd39768, 16'b1010110100101001);
	test_shift(16'b0100100100001010, 16'd62159, 16'b0010010010000101);
	test_shift(16'b0000011100000111, 16'd50899, 16'b0011100000111000);
	test_shift(16'b1110111100010100, 16'd60794, 16'b0101001110111100);
	test_shift(16'b1000000111111100, 16'd10958, 16'b0010000001111111);
	test_shift(16'b1100100101010110, 16'd7359, 16'b0110010010101011);
	test_shift(16'b0000100101111110, 16'd4800, 16'b0000100101111110);
	test_shift(16'b0001110101100111, 16'd25850, 16'b1001110001110101);
	test_shift(16'b0100110011001100, 16'd37750, 16'b0011001100010011);
	test_shift(16'b0001101110011101, 16'd17995, 16'b1110100011011100);
	test_shift(16'b1111000000000110, 16'd26188, 16'b0110111100000000);
	test_shift(16'b1000110000101101, 16'd58431, 16'b1100011000010110);
	test_shift(16'b0010111110010001, 16'd4690, 16'b1011111001000100);
	test_shift(16'b1000001011111011, 16'd58021, 16'b0101111101110000);
	test_shift(16'b1010001111110000, 16'd49888, 16'b1010001111110000);
	test_shift(16'b1011010000011101, 16'd45929, 16'b0011101101101000);
	test_shift(16'b0101000111011000, 16'd12101, 16'b0011101100001010);
	test_shift(16'b0011000000010001, 16'd35363, 16'b1000000010001001);
	test_shift(16'b1000101000110010, 16'd39806, 16'b1010001010001100);
	test_shift(16'b1000000010000111, 16'd1741, 16'b1111000000010000);
	test_shift(16'b1000101101101101, 16'd49553, 16'b0001011011011011);
	test_shift(16'b1100001101111000, 16'd1805, 16'b0001100001101111);
	test_shift(16'b1001101000011111, 16'd8543, 16'b1100110100001111);
	test_shift(16'b0010100101110111, 16'd58555, 16'b1011100101001011);
	test_shift(16'b0101100010001001, 16'd61932, 16'b1001010110001000);
	test_shift(16'b0110111010010000, 16'd36834, 16'b1011101001000001);
	test_shift(16'b0111011101011011, 16'd47656, 16'b0101101101110111);
	test_shift(16'b0101110111001010, 16'd14445, 16'b0100101110111001);
	test_shift(16'b0001011111001001, 16'd14832, 16'b0001011111001001);
	test_shift(16'b1111101001010110, 16'd57246, 16'b1011111010010101);
	test_shift(16'b0000100010110000, 16'd11488, 16'b0000100010110000);
	test_shift(16'b1101011000100010, 16'd26574, 16'b1011010110001000);
	test_shift(16'b0000010000101011, 16'd39312, 16'b0000010000101011);
	test_shift(16'b1111111100000010, 16'd10671, 16'b0111111110000001);
	test_shift(16'b0110101111110010, 16'd23703, 16'b1111100100110101);
	test_shift(16'b1110110100110111, 16'd15253, 16'b1010011011111101);
	test_shift(16'b1101000011000101, 16'd25040, 16'b1101000011000101);
	test_shift(16'b1010010110110010, 16'd32658, 16'b1001011011001010);
	test_shift(16'b0101010100111011, 16'd6253, 16'b0110101010100111);
	test_shift(16'b0011001111100010, 16'd3346, 16'b1100111110001000);
	test_shift(16'b0110111111111100, 16'd33533, 16'b1000110111111111);
	test_shift(16'b0111100011100000, 16'd49788, 16'b0000011110001110);
	test_shift(16'b0001010011111001, 16'd384, 16'b0001010011111001);
	test_shift(16'b0101001111001111, 16'd47653, 16'b0111100111101010);
	test_shift(16'b1011110000100110, 16'd10072, 16'b0010011010111100);
	test_shift(16'b1111111000100110, 16'd38060, 16'b0110111111100010);
	test_shift(16'b0101101000110101, 16'd17541, 16'b0100011010101011);
	test_shift(16'b0011110011001110, 16'd26822, 16'b0011001110001111);
	test_shift(16'b0110000101101010, 16'd58166, 16'b0101101010011000);
	test_shift(16'b1100111011001011, 16'd47732, 16'b1110110010111100);
	test_shift(16'b0001100100001110, 16'd56497, 16'b0011001000011100);
	test_shift(16'b1110101010000100, 16'd45210, 16'b0001001110101010);
	test_shift(16'b0011100010110111, 16'd15086, 16'b1100111000101101);
	test_shift(16'b1111001100010011, 16'd59885, 16'b0111111001100010);
	test_shift(16'b0110011000011001, 16'd18618, 16'b0110010110011000);
	test_shift(16'b1001111101100111, 16'd17258, 16'b1001111001111101);
	test_shift(16'b1111101110000101, 16'd45962, 16'b0001011111101110);
	test_shift(16'b1000001000110110, 16'd58843, 16'b1011010000010001);
	test_shift(16'b1101100011110110, 16'd6979, 16'b1100011110110110);
	test_shift(16'b1111001101001110, 16'd55520, 16'b1111001101001110);
	test_shift(16'b0011110101100001, 16'd34362, 16'b1000010011110101);
	test_shift(16'b1000111111011110, 16'd1789, 16'b1101000111111011);
	test_shift(16'b0011000010010101, 16'd3659, 16'b1010100110000100);
	test_shift(16'b1010001100011111, 16'd25691, 16'b1111110100011000);
	test_shift(16'b0101010101010100, 16'd15226, 16'b0101000101010101);
	test_shift(16'b0000111011101111, 16'd757, 16'b1101110111100001);
	test_shift(16'b0010000100011101, 16'd62497, 16'b0100001000111010);
	test_shift(16'b1000100111001101, 16'd63890, 16'b0010011100110110);
	test_shift(16'b0101000101100001, 16'd45498, 16'b1000010101000101);
	test_shift(16'b0101101100010001, 16'd8106, 16'b0100010101101100);
	test_shift(16'b1011000100001001, 16'd4185, 16'b0001001101100010);
	test_shift(16'b1001111110011110, 16'd58338, 16'b0111111001111010);
	test_shift(16'b0000010011110110, 16'd36148, 16'b0100111101100000);
	test_shift(16'b0000011001111001, 16'd58923, 16'b1100100000110011);
	test_shift(16'b1000100100001011, 16'd19764, 16'b1001000010111000);
	test_shift(16'b1111011100110011, 16'd19826, 16'b1101110011001111);
	test_shift(16'b0001101001100111, 16'd48164, 16'b1010011001110001);
	test_shift(16'b1011001110101000, 16'd6125, 16'b0001011001110101);
	test_shift(16'b1100001001100001, 16'd13778, 16'b0000100110000111);
	test_shift(16'b1000000110110001, 16'd15018, 16'b1100011000000110);
	test_shift(16'b0011000000010010, 16'd54506, 16'b0100100011000000);
	test_shift(16'b0111100101000100, 16'd62066, 16'b1110010100010001);
	test_shift(16'b1011011110111100, 16'd13922, 16'b1101111011110010);
	test_shift(16'b0010010001110100, 16'd47749, 16'b1000111010000100);
	test_shift(16'b0011110110001110, 16'd32729, 16'b0001110001111011);
	test_shift(16'b1010111111000100, 16'd32593, 16'b0101111110001001);
	test_shift(16'b0100010001000000, 16'd30288, 16'b0100010001000000);
	test_shift(16'b0000110000010011, 16'd59341, 16'b0110000110000010);
	test_shift(16'b0110110111100110, 16'd32120, 16'b1110011001101101);
	test_shift(16'b0111101110101010, 16'd47855, 16'b0011110111010101);
	test_shift(16'b1001011100010011, 16'd39230, 16'b1110010111000100);
	test_shift(16'b1001010100001111, 16'd65029, 16'b1010000111110010);
	test_shift(16'b1101000111010100, 16'd11200, 16'b1101000111010100);
	test_shift(16'b1001000010011101, 16'd32847, 16'b1100100001001110);
	test_shift(16'b0111001110011010, 16'd23114, 16'b0110100111001110);
	test_shift(16'b0100111001110011, 16'd1184, 16'b0100111001110011);
	test_shift(16'b1011101110010101, 16'd44600, 16'b1001010110111011);
	test_shift(16'b1110100100011000, 16'd1977, 16'b0011000111010010);
	test_shift(16'b1011100010110011, 16'd56552, 16'b1011001110111000);
	test_shift(16'b0000010100000101, 16'd9271, 16'b1000001010000010);
	test_shift(16'b1100101001111011, 16'd57586, 16'b0010100111101111);
	test_shift(16'b1001111110000000, 16'd55127, 16'b1100000001001111);
	test_shift(16'b1011001011101001, 16'd36595, 16'b1001011101001101);
	test_shift(16'b0101110111000001, 16'd46559, 16'b1010111011100000);
	test_shift(16'b1110100111000011, 16'd8550, 16'b0111000011111010);
	test_shift(16'b1101101101101101, 16'd53229, 16'b1011101101101101);
	test_shift(16'b1001101011110110, 16'd43431, 16'b0111101101001101);
	test_shift(16'b0111001101111000, 16'd1622, 16'b1101111000011100);
	test_shift(16'b1110100000100110, 16'd20864, 16'b1110100000100110);
	test_shift(16'b1100111110100011, 16'd52657, 16'b1001111101000111);
	test_shift(16'b1000110100101111, 16'd34130, 16'b0011010010111110);
	test_shift(16'b0110100001000001, 16'd15396, 16'b1000010000010110);
	test_shift(16'b1011010110011110, 16'd10740, 16'b0101100111101011);
	test_shift(16'b0101111001001000, 16'd53176, 16'b0100100001011110);
	test_shift(16'b1110011111010001, 16'd22167, 16'b1110100011110011);
	test_shift(16'b1001110111101110, 16'd41396, 16'b1101111011101001);
	test_shift(16'b1010110010101000, 16'd10045, 16'b0001010110010101);
	test_shift(16'b0000100010100011, 16'd24604, 16'b0011000010001010);
	test_shift(16'b1100011010110101, 16'd20100, 16'b0110101101011100);
	test_shift(16'b0110100001111101, 16'd49721, 16'b1111101011010000);
	test_shift(16'b0011001101101110, 16'd34323, 16'b1001101101110001);
	test_shift(16'b0001011101011001, 16'd41249, 16'b0010111010110010);
	test_shift(16'b1011111011010000, 16'd45990, 16'b1011010000101111);
	test_shift(16'b0010000100101100, 16'd61704, 16'b0010110000100001);
	test_shift(16'b1011101000111101, 16'd45830, 16'b1000111101101110);
	test_shift(16'b0110110101110001, 16'd17784, 16'b0111000101101101);
	test_shift(16'b0010011011111000, 16'd11114, 16'b1110000010011011);
	test_shift(16'b1100100001010010, 16'd60042, 16'b0100101100100001);
	test_shift(16'b0100010111001110, 16'd45856, 16'b0100010111001110);
	test_shift(16'b1110000000000001, 16'd13614, 16'b0111100000000000);
	test_shift(16'b0111000010100011, 16'd10210, 16'b1100001010001101);
	test_shift(16'b0101110100010100, 16'd8660, 16'b1101000101000101);
	test_shift(16'b1010110101100000, 16'd7325, 16'b0001010110101100);
	test_shift(16'b0000010110001000, 16'd19620, 16'b0101100010000000);
	test_shift(16'b0010111111000000, 16'd62747, 16'b0000000101111110);
	test_shift(16'b1010010100111110, 16'd57387, 16'b1111010100101001);
	test_shift(16'b0111010110101110, 16'd7066, 16'b1011100111010110);
	test_shift(16'b1110101101011010, 16'd10410, 16'b0110101110101101);
	test_shift(16'b1100000000101101, 16'd50929, 16'b1000000001011011);
	test_shift(16'b0011110010011110, 16'd25677, 16'b1100011110010011);
	test_shift(16'b0110000000010000, 16'd936, 16'b0001000001100000);
	test_shift(16'b1111000001001100, 16'd7096, 16'b0100110011110000);
	test_shift(16'b1010001100001000, 16'd54081, 16'b0100011000010001);
	test_shift(16'b0000111011101000, 16'd55794, 16'b0011101110100000);
	test_shift(16'b1110100111010011, 16'd7686, 16'b0111010011111010);
	test_shift(16'b0101110011001000, 16'd8528, 16'b0101110011001000);
	test_shift(16'b0110101110110000, 16'd6085, 16'b0111011000001101);
	test_shift(16'b0010011100110110, 16'd38602, 16'b1101100010011100);
	test_shift(16'b1101111000100011, 16'd11346, 16'b0111100010001111);
	test_shift(16'b0111011000000011, 16'd7195, 16'b0001101110110000);
	test_shift(16'b0101101111101011, 16'd63481, 16'b1101011010110111);
	test_shift(16'b1110110100010110, 16'd61254, 16'b0100010110111011);
	test_shift(16'b1011010101110110, 16'd42931, 16'b1010101110110101);
	test_shift(16'b0001001110100011, 16'd61239, 16'b1101000110001001);
	test_shift(16'b1110101011000000, 16'd34139, 16'b0000011101010110);
	test_shift(16'b1000101100100000, 16'd44645, 16'b0110010000010001);
	test_shift(16'b1110011011011000, 16'd22629, 16'b1101101100011100);
	test_shift(16'b0011010011000010, 16'd29567, 16'b0001101001100001);
	test_shift(16'b1010110000110111, 16'd5214, 16'b1110101100001101);
	test_shift(16'b0110100001000111, 16'd39169, 16'b1101000010001110);
	test_shift(16'b1101111000100010, 16'd31553, 16'b1011110001000101);
	test_shift(16'b1011010111100100, 16'd61405, 16'b1001011010111100);
	test_shift(16'b1110111100011110, 16'd42876, 16'b1110111011110001);
	test_shift(16'b1010000100001101, 16'd27704, 16'b0000110110100001);
	test_shift(16'b0110100011011110, 16'd60034, 16'b1010001101111001);
	test_shift(16'b0010001010100110, 16'd14275, 16'b0001010100110001);
	test_shift(16'b1011000000000111, 16'd1763, 16'b1000000000111101);
	test_shift(16'b1001110100111101, 16'd6909, 16'b1011001110100111);
	test_shift(16'b1001011010100011, 16'd24525, 16'b0111001011010100);
	test_shift(16'b1111000100111110, 16'd44187, 16'b1111011110001001);

    $display("SUCCESS :: FINISH CALLED FROM END OF FILE!");
    $finish;

end


endmodule

