
`timescale 1ns / 1ps
module rotl_tb;

logic clk;
logic [15:0] data, shifted, n_shifts;

rotr ROTR(
    .data_i(data),
    .n_i(n_shifts),
    .data_o(shifted)
);

task test_shift(input logic [15:0] test_data, input logic [15:0] n, input logic [15:0] correct);
    data <= test_data;
    n_shifts <= n;
    #2;

    assert(shifted == correct)
        else begin
            $error("Bad Shift: 0x%x >> 0x%x: 0x%x, Needed: 0x%x", data, n_shifts, shifted, correct);
            $finish;
        end
endtask


always begin
    clk = 1'b0;
    #1;
    clk = 1'b1;
    #1;
end


initial begin
    $fsdbDumpfile("dump.fsdb");
	$fsdbDumpvars(0, "+all");
    data = 16'b0;

    #2;

	test_shift(16'b1011101110101000, 16'd43679, 16'b0111011101010001);
	test_shift(16'b1001101010110101, 16'd12467, 16'b1011001101010110);
	test_shift(16'b1100111000101100, 16'd6557, 16'b0111000101100110);
	test_shift(16'b1100001011101000, 16'd54164, 16'b1000110000101110);
	test_shift(16'b0111101101000111, 16'd16792, 16'b0100011101111011);
	test_shift(16'b1001001010001000, 16'd4406, 16'b0010001001001010);
	test_shift(16'b0110110111001011, 16'd49260, 16'b1101110010110110);
	test_shift(16'b1010001111000001, 16'd8450, 16'b0110100011110000);
	test_shift(16'b1011100011111000, 16'd29463, 16'b1111000101110001);
	test_shift(16'b0101101110110110, 16'd11181, 16'b1101110110110010);
	test_shift(16'b0101010100100001, 16'd60731, 16'b1010010000101010);
	test_shift(16'b0001000110110010, 16'd43933, 16'b1000110110010000);
	test_shift(16'b0101011101000111, 16'd672, 16'b0101011101000111);
	test_shift(16'b1110001001001110, 16'd60671, 16'b1100010010011101);
	test_shift(16'b0110101001111111, 16'd62049, 16'b1011010100111111);
	test_shift(16'b0010011100001101, 16'd11821, 16'b0011100001101001);
	test_shift(16'b0101101110011111, 16'd11463, 16'b0011111010110111);
	test_shift(16'b0010010001101101, 16'd32673, 16'b1001001000110110);
	test_shift(16'b0010100100101111, 16'd37459, 16'b1110010100100101);
	test_shift(16'b1000010011111101, 16'd42048, 16'b1000010011111101);
	test_shift(16'b0011001010100111, 16'd23595, 16'b0101010011100110);
	test_shift(16'b0010101010001111, 16'd47398, 16'b0011110010101010);
	test_shift(16'b0110111000000100, 16'd50250, 16'b1000000100011011);
	test_shift(16'b1011110111101011, 16'd35291, 16'b1011110101110111);
	test_shift(16'b1110001100001011, 16'd60766, 16'b1000110000101111);
	test_shift(16'b0010100101010001, 16'd9719, 16'b1010001001010010);
	test_shift(16'b1000101101000101, 16'd13943, 16'b1000101100010110);
	test_shift(16'b1101110101010100, 16'd22353, 16'b0110111010101010);
	test_shift(16'b1010111001001000, 16'd29184, 16'b1010111001001000);
	test_shift(16'b1000000000101100, 16'd26027, 16'b0000010110010000);
	test_shift(16'b0101110100010101, 16'd60156, 16'b1101000101010101);
	test_shift(16'b1011111001000000, 16'd43323, 16'b1100100000010111);
	test_shift(16'b0001011110100011, 16'd11748, 16'b0011000101111010);
	test_shift(16'b0010010101000010, 16'd16602, 16'b0101000010001001);
	test_shift(16'b1100001011101110, 16'd8642, 16'b1011000010111011);
	test_shift(16'b1110110000001101, 16'd36044, 16'b1100000011011110);
	test_shift(16'b1110001010011100, 16'd27219, 16'b1001110001010011);
	test_shift(16'b1100000110100111, 16'd12265, 16'b1101001111100000);
	test_shift(16'b1001111010110000, 16'd64059, 16'b1101011000010011);
	test_shift(16'b0100111110100100, 16'd30768, 16'b0100111110100100);
	test_shift(16'b1010011011111001, 16'd14845, 16'b0011011111001101);
	test_shift(16'b0011111010001110, 16'd52134, 16'b0011100011111010);
	test_shift(16'b1001000011010101, 16'd40476, 16'b0000110101011001);
	test_shift(16'b1010010110001011, 16'd22555, 16'b1011000101110100);
	test_shift(16'b0101110101011001, 16'd9281, 16'b1010111010101100);
	test_shift(16'b0001000110111011, 16'd10626, 16'b1100010001101110);
	test_shift(16'b0111010010111111, 16'd41804, 16'b0100101111110111);
	test_shift(16'b1001101000010000, 16'd45145, 16'b0000100001001101);
	test_shift(16'b1011011111000011, 16'd34754, 16'b1110110111110000);
	test_shift(16'b0111110011100111, 16'd41229, 16'b1110011100111011);
	test_shift(16'b1000111100101011, 16'd48555, 16'b1110010101110001);
	test_shift(16'b0100101001011000, 16'd22890, 16'b1001011000010010);
	test_shift(16'b1110111111111000, 16'd7050, 16'b1111111000111011);
	test_shift(16'b1111000010110001, 16'd18561, 16'b1111100001011000);
	test_shift(16'b0101010011000011, 16'd47530, 16'b0011000011010101);
	test_shift(16'b0110101101110100, 16'd50383, 16'b1101011011101000);
	test_shift(16'b1111011101011001, 16'd26802, 16'b0111110111010110);
	test_shift(16'b1101101001101110, 16'd29575, 16'b1101110110110100);
	test_shift(16'b0001001111111011, 16'd38144, 16'b0001001111111011);
	test_shift(16'b0011111011010000, 16'd32787, 16'b0000011111011010);
	test_shift(16'b0111001010010110, 16'd50105, 16'b0100101100111001);
	test_shift(16'b0000001011011011, 16'd44591, 16'b0000010110110110);
	test_shift(16'b1111110101010111, 16'd7274, 16'b0101010111111111);
	test_shift(16'b1101100111100011, 16'd49641, 16'b1111000111101100);
	test_shift(16'b0110010011100111, 16'd9572, 16'b0111011001001110);
	test_shift(16'b0101110011010110, 16'd50077, 16'b1110011010110010);
	test_shift(16'b0100010000010101, 16'd62592, 16'b0100010000010101);
	test_shift(16'b0011110010101011, 16'd65162, 16'b0010101011001111);
	test_shift(16'b1111010010100101, 16'd52014, 16'b1101001010010111);
	test_shift(16'b1111011010110100, 16'd19149, 16'b1011010110100111);
	test_shift(16'b1110010010110001, 16'd43017, 16'b0101100011110010);
	test_shift(16'b1110000111111111, 16'd33496, 16'b1111111111100001);
	test_shift(16'b0111100110111011, 16'd38090, 16'b0110111011011110);
	test_shift(16'b0001001110010010, 16'd52374, 16'b0100100001001110);
	test_shift(16'b0000100101011101, 16'd11636, 16'b1101000010010101);
	test_shift(16'b1001111100110100, 16'd39141, 16'b1010010011111001);
	test_shift(16'b0011010101111110, 16'd63612, 16'b0101011111100011);
	test_shift(16'b1101010110011111, 16'd9838, 16'b0101011001111111);
	test_shift(16'b0100110001110101, 16'd49566, 16'b0011000111010101);
	test_shift(16'b0010110010011001, 16'd16721, 16'b1001011001001100);
	test_shift(16'b1101110010000010, 16'd14340, 16'b0010110111001000);
	test_shift(16'b0100010010010001, 16'd65478, 16'b0100010100010010);
	test_shift(16'b1001001011100110, 16'd58688, 16'b1001001011100110);
	test_shift(16'b0010100111110101, 16'd52231, 16'b1110101001010011);
	test_shift(16'b0110000011111100, 16'd23085, 16'b0000011111100011);
	test_shift(16'b1001011010100110, 16'd20231, 16'b0100110100101101);
	test_shift(16'b0100011100010101, 16'd14427, 16'b1110001010101000);
	test_shift(16'b1000100000100100, 16'd32021, 16'b0010010001000001);
	test_shift(16'b1011010100111011, 16'd12702, 16'b1101010011101110);
	test_shift(16'b1011010111001001, 16'd14399, 16'b0110101110010011);
	test_shift(16'b0001001101000011, 16'd19620, 16'b0011000100110100);
	test_shift(16'b1000010011001110, 16'd61374, 16'b0001001100111010);
	test_shift(16'b1110100010111000, 16'd242, 16'b0011101000101110);
	test_shift(16'b0000011111011010, 16'd11326, 16'b0001111101101000);
	test_shift(16'b1000111111110110, 16'd4844, 16'b1111111101101000);
	test_shift(16'b1011100000001001, 16'd15583, 16'b0111000000010011);
	test_shift(16'b1010111111000111, 16'd26797, 16'b0111111000111101);
	test_shift(16'b1011111001000111, 16'd45155, 16'b1111011111001000);
	test_shift(16'b0001011100100010, 16'd26010, 16'b1100100010000101);
	test_shift(16'b0011001011001000, 16'd6267, 16'b0101100100000110);
	test_shift(16'b0111111011111011, 16'd42924, 16'b1110111110110111);
	test_shift(16'b0100010000111011, 16'd28752, 16'b0100010000111011);
	test_shift(16'b1010000100001000, 16'd15110, 16'b0010001010000100);
	test_shift(16'b1100110100111110, 16'd60218, 16'b0100111110110011);
	test_shift(16'b1101111001011010, 16'd35660, 16'b1110010110101101);
	test_shift(16'b0111000010111101, 16'd21705, 16'b0101111010111000);
	test_shift(16'b1100110101000011, 16'd10208, 16'b1100110101000011);
	test_shift(16'b1010000000011111, 16'd64733, 16'b0000000011111101);
	test_shift(16'b0010010101110110, 16'd31036, 16'b0101011101100010);
	test_shift(16'b1000000111111111, 16'd29905, 16'b1100000011111111);
	test_shift(16'b1111010011001011, 16'd16276, 16'b1011111101001100);
	test_shift(16'b1001011001001101, 16'd12080, 16'b1001011001001101);
	test_shift(16'b0110100001001110, 16'd50952, 16'b0100111001101000);
	test_shift(16'b0111100101001101, 16'd35830, 16'b0011010111100101);
	test_shift(16'b0110010010110011, 16'd32628, 16'b0011011001001011);
	test_shift(16'b1010010101110111, 16'd6508, 16'b0101011101111010);
	test_shift(16'b1110111100011000, 16'd38361, 16'b1000110001110111);
	test_shift(16'b0101100110010011, 16'd62447, 16'b1011001100100110);
	test_shift(16'b0100010100001000, 16'd49391, 16'b1000101000010000);
	test_shift(16'b1010010111011111, 16'd10440, 16'b1101111110100101);
	test_shift(16'b1100100011011001, 16'd52158, 16'b0010001101100111);
	test_shift(16'b0100010010110100, 16'd440, 16'b1011010001000100);
	test_shift(16'b0100111001100001, 16'd45435, 16'b1100110000101001);
	test_shift(16'b0111010001010011, 16'd59887, 16'b1110100010100110);
	test_shift(16'b0101000110000101, 16'd13417, 16'b1100001010101000);
	test_shift(16'b1011011010001101, 16'd43643, 16'b1101000110110110);
	test_shift(16'b1110000011110010, 16'd47424, 16'b1110000011110010);
	test_shift(16'b0110111010011010, 16'd28721, 16'b0011011101001101);
	test_shift(16'b1010011011001100, 16'd44071, 16'b1001100101001101);
	test_shift(16'b0001001110001001, 16'd57059, 16'b0010001001110001);
	test_shift(16'b1000001000011001, 16'd41114, 16'b1000011001100000);
	test_shift(16'b1111010100111100, 16'd20171, 16'b1010011110011110);
	test_shift(16'b0010011010101010, 16'd13449, 16'b0101010100010011);
	test_shift(16'b1111001100010101, 16'd39465, 16'b1000101011111001);
	test_shift(16'b1010100011111110, 16'd25300, 16'b1110101010001111);
	test_shift(16'b0000101100011111, 16'd14540, 16'b1011000111110000);
	test_shift(16'b1010110111110101, 16'd14791, 16'b1110101101011011);
	test_shift(16'b0001000100000001, 16'd32927, 16'b0010001000000010);
	test_shift(16'b1100011111011100, 16'd45640, 16'b1101110011000111);
	test_shift(16'b0001101101111100, 16'd16445, 16'b1101101111100000);
	test_shift(16'b1100110110011000, 16'd12942, 16'b0011011001100011);
	test_shift(16'b1100101000010011, 16'd1037, 16'b0101000010011110);
	test_shift(16'b0111110010010111, 16'd33946, 16'b0010010111011111);
	test_shift(16'b0010000001011101, 16'd7440, 16'b0010000001011101);
	test_shift(16'b1101111101111011, 16'd41804, 16'b1111011110111101);
	test_shift(16'b1101010111101010, 16'd27710, 16'b0101011110101011);
	test_shift(16'b0010000110011100, 16'd6411, 16'b0011001110000100);
	test_shift(16'b0001011000111011, 16'd8896, 16'b0001011000111011);
	test_shift(16'b0100100110000010, 16'd56095, 16'b1001001100000100);
	test_shift(16'b1010101111111101, 16'd17529, 16'b1111111011010101);
	test_shift(16'b1100101000000101, 16'd65253, 16'b0010111001010000);
	test_shift(16'b1011100110001100, 16'd56148, 16'b1100101110011000);
	test_shift(16'b1111111010100100, 16'd23977, 16'b0101001001111111);
	test_shift(16'b0010011011100000, 16'd14433, 16'b0001001101110000);
	test_shift(16'b1111001010101111, 16'd23148, 16'b0010101011111111);
	test_shift(16'b0000000110101011, 16'd845, 16'b0000110101011000);
	test_shift(16'b1101000000011110, 16'd48442, 16'b0000011110110100);
	test_shift(16'b0010111110001010, 16'd48159, 16'b0101111100010100);
	test_shift(16'b1000001000011010, 16'd430, 16'b0000100001101010);
	test_shift(16'b1111000011010111, 16'd57021, 16'b1000011010111111);
	test_shift(16'b0000111111110111, 16'd63469, 16'b0111111110111000);
	test_shift(16'b0101000100010110, 16'd16952, 16'b0001011001010001);
	test_shift(16'b0101011111011111, 16'd12963, 16'b1110101011111011);
	test_shift(16'b0110011100110010, 16'd50065, 16'b0011001110011001);
	test_shift(16'b0110110100011110, 16'd51974, 16'b0111100110110100);
	test_shift(16'b0010010011100000, 16'd42855, 16'b1100000001001001);
	test_shift(16'b0010111010111000, 16'd46847, 16'b0101110101110000);
	test_shift(16'b1001010100010001, 16'd35652, 16'b0001100101010001);
	test_shift(16'b1111010000001011, 16'd22686, 16'b1101000000101111);
	test_shift(16'b0110101100111010, 16'd25614, 16'b1010110011101001);
	test_shift(16'b0011010100011011, 16'd54326, 16'b0110110011010100);
	test_shift(16'b1010101101011101, 16'd12148, 16'b1101101010110101);
	test_shift(16'b1010111110001000, 16'd47965, 16'b0111110001000101);
	test_shift(16'b1011111110000100, 16'd29844, 16'b0100101111111000);
	test_shift(16'b0001110110011010, 16'd64783, 16'b0011101100110100);
	test_shift(16'b0010111100000111, 16'd48918, 16'b0001110010111100);
	test_shift(16'b0110010000011011, 16'd27052, 16'b0100000110110110);
	test_shift(16'b0110111110011010, 16'd55256, 16'b1001101001101111);
	test_shift(16'b0000010100000111, 16'd64001, 16'b1000001010000011);
	test_shift(16'b1100011011011100, 16'd28782, 16'b0001101101110011);
	test_shift(16'b0000011101111000, 16'd52869, 16'b1100000000111011);
	test_shift(16'b0000100101000001, 16'd23791, 16'b0001001010000010);
	test_shift(16'b0000010100100011, 16'd41148, 16'b0101001000110000);
	test_shift(16'b0011010100110110, 16'd36273, 16'b0001101010011011);
	test_shift(16'b0010000110010011, 16'd45151, 16'b0100001100100110);
	test_shift(16'b0111111000010010, 16'd38784, 16'b0111111000010010);
	test_shift(16'b1000111111010010, 16'd62058, 16'b1111010010100011);
	test_shift(16'b1100100011111101, 16'd38904, 16'b1111110111001000);
	test_shift(16'b1101110001001111, 16'd4869, 16'b0111111011100010);
	test_shift(16'b1011100000110100, 16'd6224, 16'b1011100000110100);
	test_shift(16'b0010010001000010, 16'd16234, 16'b0001000010001001);
	test_shift(16'b0111001001001100, 16'd57555, 16'b1000111001001001);
	test_shift(16'b0000111101110001, 16'd38100, 16'b0001000011110111);
	test_shift(16'b1001111010010100, 16'd3173, 16'b1010010011110100);
	test_shift(16'b1000000110000011, 16'd50842, 16'b0110000011100000);
	test_shift(16'b1110010010011100, 16'd35689, 16'b0100111001110010);
	test_shift(16'b0101000001011110, 16'd8113, 16'b0010100000101111);
	test_shift(16'b1010111110110101, 16'd60024, 16'b1011010110101111);
	test_shift(16'b0011110010001110, 16'd38267, 16'b1001000111000111);
	test_shift(16'b0111010101110001, 16'd62737, 16'b1011101010111000);
	test_shift(16'b1101001101000010, 16'd48159, 16'b1010011010000101);
	test_shift(16'b0000101010010110, 16'd13255, 16'b0010110000010101);
	test_shift(16'b0100111010000100, 16'd56162, 16'b0001001110100001);
	test_shift(16'b0010111100101001, 16'd5733, 16'b0100100101111001);
	test_shift(16'b1110110110111011, 16'd63272, 16'b1011101111101101);
	test_shift(16'b0001001000001100, 16'd35876, 16'b1100000100100000);
	test_shift(16'b0001110011011110, 16'd1334, 16'b0111100001110011);
	test_shift(16'b0001101010110111, 16'd35696, 16'b0001101010110111);
	test_shift(16'b1010000110101000, 16'd2399, 16'b0100001101010001);
	test_shift(16'b1110000000110101, 16'd16023, 16'b0110101111000000);
	test_shift(16'b1110011111111101, 16'd6245, 16'b1110111100111111);
	test_shift(16'b1000111001111101, 16'd9144, 16'b0111110110001110);
	test_shift(16'b0000001100001100, 16'd29228, 16'b0011000011000000);
	test_shift(16'b0110110110011010, 16'd64858, 16'b0110011010011011);
	test_shift(16'b0111101100100001, 16'd15262, 16'b1110110010000101);
	test_shift(16'b0100010111111010, 16'd30737, 16'b0010001011111101);
	test_shift(16'b1010000100000001, 16'd14683, 16'b0010000000110100);
	test_shift(16'b1011000111111111, 16'd27420, 16'b0001111111111011);
	test_shift(16'b1001111010011111, 16'd8834, 16'b1110011110100111);
	test_shift(16'b0001101111000010, 16'd2491, 16'b0111100001000011);
	test_shift(16'b1011101011000001, 16'd62111, 16'b0111010110000011);
	test_shift(16'b1000010100011010, 16'd33115, 16'b1010001101010000);
	test_shift(16'b0010100111000101, 16'd24622, 16'b1010011100010100);
	test_shift(16'b1010011010110111, 16'd34331, 16'b1101011011110100);
	test_shift(16'b1100001111010100, 16'd49103, 16'b1000011110101001);
	test_shift(16'b1000010011100110, 16'd21834, 16'b0011100110100001);
	test_shift(16'b0011011110000000, 16'd62295, 16'b0000000001101111);
	test_shift(16'b1011110110000001, 16'd39547, 16'b1011000000110111);
	test_shift(16'b0100000110000000, 16'd3361, 16'b0010000011000000);
	test_shift(16'b0111010010110110, 16'd31428, 16'b0110011101001011);
	test_shift(16'b0101000000100011, 16'd37206, 16'b1000110101000000);
	test_shift(16'b1110110100110101, 16'd52097, 16'b1111011010011010);
	test_shift(16'b0110010011001011, 16'd2414, 16'b1001001100101101);
	test_shift(16'b0110101101010011, 16'd37236, 16'b0011011010110101);
	test_shift(16'b1111000101111011, 16'd35352, 16'b0111101111110001);
	test_shift(16'b0001001100100000, 16'd10974, 16'b0100110010000000);
	test_shift(16'b0000010111100111, 16'd37480, 16'b1110011100000101);
	test_shift(16'b1000110101010111, 16'd45394, 16'b1110001101010101);
	test_shift(16'b1111101010110101, 16'd63112, 16'b1011010111111010);
	test_shift(16'b0010100001101110, 16'd46249, 16'b0011011100010100);
	test_shift(16'b0111110001010000, 16'd52082, 16'b0001111100010100);
	test_shift(16'b1001100001101010, 16'd25744, 16'b1001100001101010);
	test_shift(16'b0101111010001011, 16'd6374, 16'b0010110101111010);
	test_shift(16'b0010011111010011, 16'd61079, 16'b1010011001001111);
	test_shift(16'b0001110111101111, 16'd42875, 16'b1011110111100011);
	test_shift(16'b1001011110111100, 16'd5471, 16'b0010111101111001);
	test_shift(16'b1100110010000001, 16'd55794, 16'b0111001100100000);
	test_shift(16'b1011110100100011, 16'd32351, 16'b0111101001000111);
	test_shift(16'b0011110000001100, 16'd42074, 16'b0000001100001111);
	test_shift(16'b0100000000110000, 16'd64412, 16'b0000001100000100);
	test_shift(16'b0001011010001001, 16'd19869, 16'b1011010001001000);
	test_shift(16'b0110101001010111, 16'd34130, 16'b1101101010010101);
	test_shift(16'b1000000010110011, 16'd6015, 16'b0000000101100111);
	test_shift(16'b0100100100001101, 16'd29938, 16'b0101001001000011);
	test_shift(16'b0110110110101101, 16'd14653, 16'b0110110101101011);
	test_shift(16'b1111111111000100, 16'd3138, 16'b0011111111110001);
	test_shift(16'b0011010100000001, 16'd43421, 16'b1010100000001001);
	test_shift(16'b1100101011100101, 16'd2205, 16'b0101011100101110);
	test_shift(16'b1001000000100000, 16'd20130, 16'b0010010000001000);
	test_shift(16'b0100100110000010, 16'd17409, 16'b0010010011000001);
	test_shift(16'b1010011000100110, 16'd26959, 16'b0100110001001101);
	test_shift(16'b0010011001101100, 16'd27012, 16'b1100001001100110);
	test_shift(16'b1000011010101101, 16'd2588, 16'b0110101011011000);
	test_shift(16'b0101011011111111, 16'd35280, 16'b0101011011111111);
	test_shift(16'b1000110101001000, 16'd7078, 16'b0010001000110101);
	test_shift(16'b1110011000101111, 16'd50485, 16'b0111111100110001);
	test_shift(16'b1011111010111000, 16'd19702, 16'b1110001011111010);
	test_shift(16'b0011111111110001, 16'd38149, 16'b1000100111111111);
	test_shift(16'b0011101101101010, 16'd14906, 16'b1101101010001110);
	test_shift(16'b1111111011001010, 16'd30838, 16'b0010101111111011);
	test_shift(16'b1111101010100000, 16'd21088, 16'b1111101010100000);
	test_shift(16'b1001110110010100, 16'd158, 16'b0111011001010010);
	test_shift(16'b1000010110001001, 16'd23542, 16'b0010011000010110);
	test_shift(16'b1111011101000010, 16'd48182, 16'b0000101111011101);
	test_shift(16'b0111101001100101, 16'd42261, 16'b0010101111010011);
	test_shift(16'b1000010100001100, 16'd51854, 16'b0001010000110010);
	test_shift(16'b1011011111100000, 16'd20279, 16'b1100000101101111);
	test_shift(16'b1100111101001101, 16'd13269, 16'b0110111001111010);
	test_shift(16'b0000001111110100, 16'd35734, 16'b1101000000001111);
	test_shift(16'b1010001010101111, 16'd8123, 16'b0101010111110100);
	test_shift(16'b0111000011110000, 16'd29285, 16'b1000001110000111);
	test_shift(16'b0111001110101010, 16'd58682, 16'b1110101010011100);
	test_shift(16'b0010101110110110, 16'd11139, 16'b1100010101110110);
	test_shift(16'b1010110010001011, 16'd8287, 16'b0101100100010111);
	test_shift(16'b1101011110011011, 16'd54250, 16'b1110011011110101);
	test_shift(16'b0010111000001110, 16'd30600, 16'b0000111000101110);
	test_shift(16'b1010001000100010, 16'd20302, 16'b1000100010001010);
	test_shift(16'b1011011010000101, 16'd62173, 16'b1011010000101101);
	test_shift(16'b0000000101110011, 16'd61728, 16'b0000000101110011);
	test_shift(16'b0101000011010000, 16'd39732, 16'b0000010100001101);
	test_shift(16'b0100111100111111, 16'd59598, 16'b0011110011111101);
	test_shift(16'b1011110100000010, 16'd49122, 16'b1010111101000000);
	test_shift(16'b1011011101100010, 16'd7963, 16'b1110110001010110);
	test_shift(16'b0010110010001001, 16'd26367, 16'b0101100100010010);
	test_shift(16'b0111001101001100, 16'd3077, 16'b0110001110011010);
	test_shift(16'b0111000010000000, 16'd3633, 16'b0011100001000000);
	test_shift(16'b1000111100110010, 16'd53127, 16'b0110010100011110);
	test_shift(16'b1110100011011110, 16'd50428, 16'b1000110111101110);
	test_shift(16'b1000111010000000, 16'd31325, 16'b0111010000000100);
	test_shift(16'b1111101100101000, 16'd35290, 16'b1100101000111110);
	test_shift(16'b0010101101101100, 16'd30107, 16'b0110110110000101);
	test_shift(16'b0101010101011000, 16'd62535, 16'b1011000010101010);
	test_shift(16'b1010010010110111, 16'd22529, 16'b1101001001011011);
	test_shift(16'b1111001111101000, 16'd19440, 16'b1111001111101000);
	test_shift(16'b0110000111010100, 16'd51493, 16'b1010001100001110);
	test_shift(16'b0001111111111110, 16'd56982, 16'b1111100001111111);
	test_shift(16'b0010010101111010, 16'd37678, 16'b1001010111101000);
	test_shift(16'b0010110110010100, 16'd64682, 16'b0110010100001011);
	test_shift(16'b0101100111000101, 16'd48871, 16'b1000101010110011);
	test_shift(16'b0010010011010011, 16'd21576, 16'b1101001100100100);
	test_shift(16'b1001111011010101, 16'd63590, 16'b0101011001111011);
	test_shift(16'b0011011000001000, 16'd64337, 16'b0001101100000100);
	test_shift(16'b1000000100111100, 16'd1484, 16'b0001001111001000);
	test_shift(16'b1000100100011000, 16'd55959, 16'b0011000100010010);
	test_shift(16'b1101011101001101, 16'd46065, 16'b1110101110100110);
	test_shift(16'b1111110111101011, 16'd23531, 16'b1011110101111111);
	test_shift(16'b0110111000000010, 16'd34540, 16'b1110000000100110);
	test_shift(16'b0010100011010000, 16'd2413, 16'b0100011010000001);
	test_shift(16'b0001001100100001, 16'd18657, 16'b1000100110010000);
	test_shift(16'b1011011100101011, 16'd38490, 16'b1100101011101101);
	test_shift(16'b0100010110010011, 16'd27591, 16'b0010011010001011);
	test_shift(16'b1111111110100000, 16'd1116, 16'b1111101000001111);
	test_shift(16'b1001000100001100, 16'd6816, 16'b1001000100001100);
	test_shift(16'b1100011011101110, 16'd332, 16'b0110111011101100);
	test_shift(16'b0100000111101000, 16'd48673, 16'b0010000011110100);
	test_shift(16'b0111110001001000, 16'd49205, 16'b0100001111100010);
	test_shift(16'b1111110111100001, 16'd51341, 16'b1110111100001111);
	test_shift(16'b1111001001000101, 16'd36012, 16'b0010010001011111);
	test_shift(16'b1101001111111111, 16'd4282, 16'b1111111111110100);
	test_shift(16'b0100011001010011, 16'd43400, 16'b0101001101000110);
	test_shift(16'b0110011100001001, 16'd14141, 16'b0011100001001011);
	test_shift(16'b0101000111010011, 16'd20087, 16'b1010011010100011);
	test_shift(16'b1011101100111100, 16'd44130, 16'b0010111011001111);
	test_shift(16'b1101011010001100, 16'd56465, 16'b0110101101000110);
	test_shift(16'b1000011101001101, 16'd10278, 16'b0011011000011101);
	test_shift(16'b0101011001000010, 16'd32843, 16'b1100100001001010);
	test_shift(16'b1001011100101000, 16'd48130, 16'b0010010111001010);
	test_shift(16'b1111100101111111, 16'd18670, 16'b1110010111111111);
	test_shift(16'b0011011111100010, 16'd39049, 16'b1111000100011011);
	test_shift(16'b1000111010111010, 16'd48170, 16'b1010111010100011);
	test_shift(16'b0110011111000111, 16'd47109, 16'b0011101100111110);
	test_shift(16'b1010011001010100, 16'd60678, 16'b0101001010011001);
	test_shift(16'b1011100001000111, 16'd27100, 16'b1000010001111011);
	test_shift(16'b1011110111110101, 16'd31822, 16'b1111011111010110);
	test_shift(16'b1011010001100001, 16'd58886, 16'b1000011011010001);
	test_shift(16'b1010000101110010, 16'd34720, 16'b1010000101110010);
	test_shift(16'b1010010011000000, 16'd28623, 16'b0100100110000001);
	test_shift(16'b0110001001000001, 16'd27868, 16'b0010010000010110);
	test_shift(16'b0100111110000101, 16'd11264, 16'b0100111110000101);
	test_shift(16'b0010011100101011, 16'd10020, 16'b1011001001110010);
	test_shift(16'b0100000000100110, 16'd37859, 16'b1100100000000100);
	test_shift(16'b0000101111000010, 16'd47027, 16'b0100000101111000);
	test_shift(16'b1101101011101111, 16'd2180, 16'b1111110110101110);
	test_shift(16'b1010011110010100, 16'd1737, 16'b1100101001010011);
	test_shift(16'b1100100011011001, 16'd46783, 16'b1001000110110011);
	test_shift(16'b1010101001000110, 16'd49881, 16'b0010001101010101);
	test_shift(16'b0100100110111001, 16'd1040, 16'b0100100110111001);
	test_shift(16'b1101111000111011, 16'd59556, 16'b1011110111100011);
	test_shift(16'b1101000111100001, 16'd64670, 16'b0100011110000111);
	test_shift(16'b0011011000110010, 16'd10434, 16'b1000110110001100);
	test_shift(16'b0100110010110001, 16'd53569, 16'b1010011001011000);
	test_shift(16'b1111001111000100, 16'd34479, 16'b1110011110001001);
	test_shift(16'b1001110101011111, 16'd59617, 16'b1100111010101111);
	test_shift(16'b0011111111101111, 16'd4786, 16'b1100111111111011);
	test_shift(16'b0010001000000001, 16'd50386, 16'b0100100010000000);
	test_shift(16'b0101101010000001, 16'd48324, 16'b0001010110101000);
	test_shift(16'b1110011110011001, 16'd16414, 16'b1001111001100111);
	test_shift(16'b0000000010100101, 16'd62662, 16'b1001010000000010);
	test_shift(16'b0010110111010110, 16'd21985, 16'b0001011011101011);
	test_shift(16'b0001110011111100, 16'd45991, 16'b1111100000111001);
	test_shift(16'b1011011110000110, 16'd30604, 16'b0111100001101011);
	test_shift(16'b1100101100000100, 16'd10497, 16'b0110010110000010);
	test_shift(16'b0110111101100001, 16'd49542, 16'b1000010110111101);
	test_shift(16'b0100101010101110, 16'd50041, 16'b0101011100100101);
	test_shift(16'b1011110011001111, 16'd23480, 16'b1100111110111100);
	test_shift(16'b0010001111000000, 16'd11462, 16'b0000000010001111);
	test_shift(16'b1101011011010000, 16'd56665, 16'b0110100001101011);
	test_shift(16'b1100001110100001, 16'd44587, 16'b0111010000111000);
	test_shift(16'b0101100110010010, 16'd59434, 16'b0110010010010110);
	test_shift(16'b0000000101011010, 16'd36069, 16'b1101000000001010);
	test_shift(16'b0111110001010100, 16'd46753, 16'b0011111000101010);
	test_shift(16'b0011110000100101, 16'd7969, 16'b1001111000010010);
	test_shift(16'b1111111110010111, 16'd10648, 16'b1001011111111111);
	test_shift(16'b1101111100101111, 16'd19569, 16'b1110111110010111);
	test_shift(16'b0100100000001010, 16'd33865, 16'b0000010100100100);
	test_shift(16'b0101011010011110, 16'd19150, 16'b0101101001111001);
	test_shift(16'b0001000001111110, 16'd63669, 16'b1111000010000011);
	test_shift(16'b1011011000111011, 16'd57222, 16'b1110111011011000);
	test_shift(16'b0101010000010110, 16'd35208, 16'b0001011001010100);
	test_shift(16'b1001001100111101, 16'd53574, 16'b1111011001001100);
	test_shift(16'b0001101110011100, 16'd30169, 16'b1100111000001101);
	test_shift(16'b1101000100001000, 16'd25463, 16'b0001000110100010);
	test_shift(16'b0100011110011100, 16'd41323, 16'b1111001110001000);
	test_shift(16'b0100011000011010, 16'd65047, 16'b0011010010001100);
	test_shift(16'b0000111001000101, 16'd60544, 16'b0000111001000101);
	test_shift(16'b0100100110000010, 16'd17078, 16'b0000100100100110);
	test_shift(16'b1101100111000100, 16'd13460, 16'b0100110110011100);
	test_shift(16'b1010111011111001, 16'd20595, 16'b0011010111011111);
	test_shift(16'b1010111111011100, 16'd33833, 16'b1110111001010111);
	test_shift(16'b0000101110101000, 16'd19598, 16'b0010111010100000);
	test_shift(16'b0110011111000110, 16'd31886, 16'b1001111100011001);
	test_shift(16'b0011010000000010, 16'd19908, 16'b0010001101000000);
	test_shift(16'b1101110011000110, 16'd41305, 16'b0110001101101110);
	test_shift(16'b1001000101101011, 16'd64845, 16'b1000101101011100);
	test_shift(16'b1100100110100010, 16'd42683, 16'b0011010001011001);
	test_shift(16'b1001000101011010, 16'd25637, 16'b1101010010001010);
	test_shift(16'b0011110110100101, 16'd64154, 16'b0110100101001111);
	test_shift(16'b0000010100111001, 16'd60020, 16'b1001000001010011);
	test_shift(16'b0010010101111000, 16'd61059, 16'b0000010010101111);
	test_shift(16'b0011010100101111, 16'd32249, 16'b1001011110011010);
	test_shift(16'b1010011101111001, 16'd26789, 16'b1100110100111011);
	test_shift(16'b1010111101000001, 16'd5945, 16'b1010000011010111);
	test_shift(16'b1010011011101110, 16'd43901, 16'b0011011101110101);
	test_shift(16'b1011011101001101, 16'd41873, 16'b1101101110100110);
	test_shift(16'b1011010010011100, 16'd40520, 16'b1001110010110100);
	test_shift(16'b1001001011001110, 16'd20595, 16'b1101001001011001);
	test_shift(16'b0001101100111011, 16'd17187, 16'b0110001101100111);
	test_shift(16'b1111111010110111, 16'd36508, 16'b1110101101111111);
	test_shift(16'b0100110001100010, 16'd48144, 16'b0100110001100010);
	test_shift(16'b1111001101101010, 16'd59712, 16'b1111001101101010);
	test_shift(16'b1110100010011011, 16'd37358, 16'b1010001001101111);
	test_shift(16'b1110110010101010, 16'd64508, 16'b1100101010101110);
	test_shift(16'b0110100001100101, 16'd14251, 16'b0000110010101101);
	test_shift(16'b1011100000101000, 16'd38826, 16'b0000101000101110);
	test_shift(16'b0110011100110010, 16'd5632, 16'b0110011100110010);
	test_shift(16'b0001000111010111, 16'd45950, 16'b0100011101011100);
	test_shift(16'b1000100010010101, 16'd14069, 16'b1010110001000100);
	test_shift(16'b1101100111000011, 16'd41001, 16'b1110000111101100);
	test_shift(16'b1001100001101001, 16'd31284, 16'b1001100110000110);
	test_shift(16'b1001101101100001, 16'd22719, 16'b0011011011000011);
	test_shift(16'b0001110111100010, 16'd21026, 16'b1000011101111000);
	test_shift(16'b0110110010000010, 16'd27377, 16'b0011011001000001);
	test_shift(16'b0000101001001111, 16'd18318, 16'b0010100100111100);
	test_shift(16'b0000111110111100, 16'd20203, 16'b1111011110000001);
	test_shift(16'b0111101001001110, 16'd2821, 16'b0111001111010010);
	test_shift(16'b1101101000110011, 16'd45045, 16'b1001111011010001);
	test_shift(16'b0000001110001100, 16'd64914, 16'b0000000011100011);
	test_shift(16'b0110100001000000, 16'd9807, 16'b1101000010000000);
	test_shift(16'b0011001011000110, 16'd4143, 16'b0110010110001100);
	test_shift(16'b0001000100110000, 16'd35457, 16'b0000100010011000);
	test_shift(16'b0100110100001101, 16'd58704, 16'b0100110100001101);
	test_shift(16'b1001011011101110, 16'd55907, 16'b1101001011011101);
	test_shift(16'b1010111011100100, 16'd799, 16'b0101110111001001);
	test_shift(16'b0001101100001100, 16'd39745, 16'b0000110110000110);
	test_shift(16'b0101010011000011, 16'd25869, 16'b1010011000011010);
	test_shift(16'b0100111101000000, 16'd3973, 16'b0000001001111010);
	test_shift(16'b0101101111110010, 16'd16261, 16'b1001001011011111);
	test_shift(16'b0000001000001111, 16'd48594, 16'b1100000010000011);
	test_shift(16'b1101001100111011, 16'd19497, 16'b1001110111101001);
	test_shift(16'b1010011010000001, 16'd22882, 16'b0110100110100000);
	test_shift(16'b1001111010110111, 16'd64873, 16'b0101101111001111);
	test_shift(16'b1010000111101001, 16'd25798, 16'b1010011010000111);
	test_shift(16'b0000010001110010, 16'd25829, 16'b1001000000100011);
	test_shift(16'b1000001111001100, 16'd44878, 16'b0000111100110010);
	test_shift(16'b1010000100010000, 16'd35976, 16'b0001000010100001);
	test_shift(16'b1000110000011000, 16'd34999, 16'b0011000100011000);
	test_shift(16'b0111100010001110, 16'd30318, 16'b1110001000111001);
	test_shift(16'b1010110111001100, 16'd4267, 16'b1011100110010101);
	test_shift(16'b1100010010110100, 16'd300, 16'b0100101101001100);
	test_shift(16'b0101000010101000, 16'd40409, 16'b0101010000101000);
	test_shift(16'b0011100110000000, 16'd4910, 16'b1110011000000000);
	test_shift(16'b0100110111010001, 16'd15826, 16'b0101001101110100);
	test_shift(16'b1111001111001110, 16'd50493, 16'b1001111001110111);
	test_shift(16'b0000111010010110, 16'd18158, 16'b0011101001011000);
	test_shift(16'b0011001110100100, 16'd23988, 16'b0100001100111010);
	test_shift(16'b0100000001100011, 16'd50116, 16'b0011010000000110);
	test_shift(16'b1000110101101100, 16'd45316, 16'b1100100011010110);
	test_shift(16'b0001000011010100, 16'd9124, 16'b0100000100001101);
	test_shift(16'b1001011101010110, 16'd54247, 16'b1010110100101110);
	test_shift(16'b0111101011010011, 16'd46398, 16'b1110101101001101);
	test_shift(16'b1011010101101000, 16'd43315, 16'b0001011010101101);
	test_shift(16'b0100110000011000, 16'd7795, 16'b0000100110000011);
	test_shift(16'b1010110101001111, 16'd9848, 16'b0100111110101101);
	test_shift(16'b1110000010111110, 16'd64228, 16'b1110111000001011);
	test_shift(16'b0000000001010011, 16'd29356, 16'b0000010100110000);
	test_shift(16'b1101111101000111, 16'd54163, 16'b1111101111101000);
	test_shift(16'b0011111100011011, 16'd20905, 16'b1000110110011111);
	test_shift(16'b1110101010000100, 16'd29225, 16'b0100001001110101);
	test_shift(16'b1100001010000111, 16'd27663, 16'b1000010100001111);
	test_shift(16'b0000011000001111, 16'd60431, 16'b0000110000011110);
	test_shift(16'b1100110000111011, 16'd8417, 16'b1110011000011101);
	test_shift(16'b0001101100001100, 16'd52754, 16'b0000011011000011);
	test_shift(16'b0011011110001011, 16'd56551, 16'b0001011001101111);
	test_shift(16'b1001111001111110, 16'd60333, 16'b1111001111110100);
	test_shift(16'b0011011111001011, 16'd55295, 16'b0110111110010110);
	test_shift(16'b1001011001101000, 16'd46459, 16'b1100110100010010);
	test_shift(16'b1100101011011001, 16'd53642, 16'b1011011001110010);
	test_shift(16'b1101101010100101, 16'd19944, 16'b1010010111011010);
	test_shift(16'b1100010001100100, 16'd48585, 16'b0011001001100010);
	test_shift(16'b0001111101100000, 16'd32164, 16'b0000000111110110);
	test_shift(16'b0110101100111011, 16'd27366, 16'b1110110110101100);
	test_shift(16'b0000001110001000, 16'd48047, 16'b0000011100010000);
	test_shift(16'b0000110111110101, 16'd46656, 16'b0000110111110101);
	test_shift(16'b0010101101110011, 16'd35630, 16'b1010110111001100);
	test_shift(16'b1001000011100000, 16'd18771, 16'b0001001000011100);
	test_shift(16'b0010110110011111, 16'd17192, 16'b1001111100101101);
	test_shift(16'b1010010010010000, 16'd11937, 16'b0101001001001000);
	test_shift(16'b0111001100110101, 16'd17771, 16'b0110011010101110);
	test_shift(16'b0110111110101011, 16'd17605, 16'b0101101101111101);
	test_shift(16'b0001101001100100, 16'd3392, 16'b0001101001100100);
	test_shift(16'b1001011011010111, 16'd30918, 16'b0101111001011011);
	test_shift(16'b1010011001101100, 16'd52308, 16'b1100101001100110);
	test_shift(16'b0010000100110101, 16'd12146, 16'b0100100001001101);
	test_shift(16'b1100010011111001, 16'd64130, 16'b0111000100111110);
	test_shift(16'b1111010011000101, 16'd14640, 16'b1111010011000101);
	test_shift(16'b1011100100000100, 16'd48116, 16'b0100101110010000);
	test_shift(16'b1101100110010101, 16'd12922, 16'b0110010101110110);
	test_shift(16'b0001110101000101, 16'd26180, 16'b0101000111010100);
	test_shift(16'b0001111101101011, 16'd26474, 16'b1101101011000111);
	test_shift(16'b0010001110000011, 16'd10055, 16'b0000011001000111);
	test_shift(16'b0110101110100101, 16'd25744, 16'b0110101110100101);
	test_shift(16'b1010101010111001, 16'd13478, 16'b1110011010101010);
	test_shift(16'b0001101101001101, 16'd64494, 16'b0110110100110100);
	test_shift(16'b0111011111010101, 16'd29590, 16'b0101010111011111);
	test_shift(16'b0100011110001001, 16'd50147, 16'b0010100011110001);
	test_shift(16'b1101010010100100, 16'd11607, 16'b0100100110101001);
	test_shift(16'b0000001001011011, 16'd10006, 16'b0110110000001001);
	test_shift(16'b0010101100000010, 16'd59683, 16'b0100010101100000);
	test_shift(16'b1001111101110001, 16'd32516, 16'b0001100111110111);
	test_shift(16'b0100101010100101, 16'd50301, 16'b0101010100101010);
	test_shift(16'b1010100111000100, 16'd17293, 16'b0100111000100101);
	test_shift(16'b1100011100100110, 16'd7512, 16'b0010011011000111);
	test_shift(16'b0110000011101001, 16'd8977, 16'b1011000001110100);
	test_shift(16'b1111100011001000, 16'd41182, 16'b1110001100100011);
	test_shift(16'b0001001011111010, 16'd7817, 16'b0111110100001001);
	test_shift(16'b1011110000011011, 16'd23067, 16'b1000001101110111);
	test_shift(16'b1101000111000110, 16'd16883, 16'b1101101000111000);
	test_shift(16'b1000101010100101, 16'd56938, 16'b1010100101100010);
	test_shift(16'b1010000011111010, 16'd42309, 16'b1101010100000111);
	test_shift(16'b1111101000000101, 16'd53722, 16'b1000000101111110);
	test_shift(16'b0111101001110000, 16'd53707, 16'b0100111000001111);
	test_shift(16'b0000101011100000, 16'd55082, 16'b1011100000000010);
	test_shift(16'b1100101010001111, 16'd31680, 16'b1100101010001111);
	test_shift(16'b0101011111101001, 16'd14502, 16'b1010010101011111);
	test_shift(16'b0101110011101101, 16'd20173, 16'b1110011101101010);
	test_shift(16'b0010001001111100, 16'd26253, 16'b0001001111100001);
	test_shift(16'b1000001010101110, 16'd41904, 16'b1000001010101110);
	test_shift(16'b1101101100001010, 16'd47510, 16'b0010101101101100);
	test_shift(16'b1011111101101111, 16'd12558, 16'b1111110110111110);
	test_shift(16'b1011011000011010, 16'd9090, 16'b1010110110000110);
	test_shift(16'b1110100111110100, 16'd29404, 16'b1001111101001110);
	test_shift(16'b1101101110010010, 16'd12845, 16'b1101110010010110);
	test_shift(16'b0000111101110111, 16'd17080, 16'b0111011100001111);
	test_shift(16'b0100100111111011, 16'd45239, 16'b1111011010010011);
	test_shift(16'b0101101000100011, 16'd17675, 16'b0100010001101011);
	test_shift(16'b1111001101010010, 16'd52899, 16'b0101111001101010);
	test_shift(16'b1001100010101000, 16'd10980, 16'b1000100110001010);
	test_shift(16'b0001111100001110, 16'd57292, 16'b1111000011100001);
	test_shift(16'b1000111111000011, 16'd14597, 16'b0001110001111110);
	test_shift(16'b0000101111010101, 16'd4097, 16'b1000010111101010);
	test_shift(16'b0000001011101011, 16'd31394, 16'b1100000010111010);
	test_shift(16'b0011000111100010, 16'd15932, 16'b0001111000100011);
	test_shift(16'b0111101001100100, 16'd20101, 16'b0010001111010011);
	test_shift(16'b1001110111011100, 16'd14221, 16'b1110111011100100);
	test_shift(16'b0111011001111100, 16'd23683, 16'b1000111011001111);
	test_shift(16'b1110010000010000, 16'd54316, 16'b0100000100001110);
	test_shift(16'b1100011111010110, 16'd48399, 16'b1000111110101101);
	test_shift(16'b1100010000010111, 16'd64590, 16'b0001000001011111);
	test_shift(16'b1000100101010100, 16'd7232, 16'b1000100101010100);
	test_shift(16'b0101100001010111, 16'd593, 16'b1010110000101011);
	test_shift(16'b0010011010011011, 16'd16165, 16'b1101100100110100);
	test_shift(16'b0000000111110000, 16'd12037, 16'b1000000000001111);
	test_shift(16'b1111111101000110, 16'd1608, 16'b0100011011111111);
	test_shift(16'b0100111111111011, 16'd11671, 16'b1111011010011111);
	test_shift(16'b1111001100111010, 16'd8355, 16'b0101111001100111);
	test_shift(16'b0101100011110110, 16'd5661, 16'b1100011110110010);
	test_shift(16'b1111010000101100, 16'd12032, 16'b1111010000101100);
	test_shift(16'b0110100111100001, 16'd8122, 16'b0111100001011010);
	test_shift(16'b0101000011000000, 16'd34864, 16'b0101000011000000);
	test_shift(16'b1101101010000111, 16'd39288, 16'b1000011111011010);
	test_shift(16'b0001110111010011, 16'd33885, 16'b1110111010011000);
	test_shift(16'b1111011101010111, 16'd32065, 16'b1111101110101011);
	test_shift(16'b1100000011010010, 16'd11357, 16'b0000011010010110);
	test_shift(16'b0101001010000101, 16'd7479, 16'b0000101010100101);
	test_shift(16'b1111010100000100, 16'd28324, 16'b0100111101010000);
	test_shift(16'b1101000101011101, 16'd41424, 16'b1101000101011101);
	test_shift(16'b1011100001100111, 16'd16840, 16'b0110011110111000);
	test_shift(16'b1000110110111110, 16'd49118, 16'b0011011011111010);
	test_shift(16'b1110001101011100, 16'd17373, 16'b0001101011100111);
	test_shift(16'b0100111110110001, 16'd58321, 16'b1010011111011000);
	test_shift(16'b1110111110001101, 16'd39874, 16'b0111101111100011);
	test_shift(16'b1001100100100110, 16'd1556, 16'b0110100110010010);
	test_shift(16'b1101111000100010, 16'd53442, 16'b1011011110001000);
	test_shift(16'b1010100011011001, 16'd58944, 16'b1010100011011001);
	test_shift(16'b1000101111000110, 16'd27450, 16'b1111000110100010);
	test_shift(16'b0011010110010100, 16'd15732, 16'b0100001101011001);
	test_shift(16'b1101011011101100, 16'd6605, 16'b1011011101100110);
	test_shift(16'b0000110111000110, 16'd18907, 16'b1011100011000001);
	test_shift(16'b0011110110011011, 16'd60219, 16'b1011001101100111);
	test_shift(16'b0100101001100000, 16'd59041, 16'b0010010100110000);
	test_shift(16'b1100110001110000, 16'd25194, 16'b0001110000110011);
	test_shift(16'b0001101010000110, 16'd27833, 16'b0100001100001101);
	test_shift(16'b0011010111100011, 16'd51805, 16'b1010111100011001);
	test_shift(16'b1111110010000000, 16'd25408, 16'b1111110010000000);
	test_shift(16'b0101001011010110, 16'd41821, 16'b1001011010110010);
	test_shift(16'b1000111011100110, 16'd60092, 16'b1110111001101000);
	test_shift(16'b1111000100110010, 16'd33519, 16'b1110001001100101);
	test_shift(16'b1001100011111000, 16'd35611, 16'b0001111100010011);
	test_shift(16'b0100011111010000, 16'd40393, 16'b1110100000100011);
	test_shift(16'b1011100010101000, 16'd28872, 16'b1010100010111000);
	test_shift(16'b0111110000000000, 16'd13324, 16'b1100000000000111);
	test_shift(16'b1101001010001000, 16'd61461, 16'b0100011010010100);
	test_shift(16'b1101111001010111, 16'd61969, 16'b1110111100101011);
	test_shift(16'b1101000011010110, 16'd37927, 16'b1010110110100001);
	test_shift(16'b0101011100101000, 16'd26719, 16'b1010111001010000);
	test_shift(16'b0111000100111000, 16'd55750, 16'b1110000111000100);
	test_shift(16'b1011010001011111, 16'd62463, 16'b0110100010111111);
	test_shift(16'b1011101110001001, 16'd45430, 16'b0010011011101110);
	test_shift(16'b0111010011011001, 16'd55473, 16'b1011101001101100);
	test_shift(16'b1111001101110100, 16'd6654, 16'b1100110111010011);
	test_shift(16'b1000111100001010, 16'd49869, 16'b0111100001010100);
	test_shift(16'b0111011100001000, 16'd50179, 16'b0000111011100001);
	test_shift(16'b1010111001001011, 16'd24432, 16'b1010111001001011);
	test_shift(16'b1001010110111101, 16'd25158, 16'b1111011001010110);
	test_shift(16'b0111111110000001, 16'd36938, 16'b1110000001011111);
	test_shift(16'b0010001111011111, 16'd48640, 16'b0010001111011111);
	test_shift(16'b1000110100010010, 16'd23464, 16'b0001001010001101);
	test_shift(16'b0010000010011110, 16'd8908, 16'b0000100111100010);
	test_shift(16'b0100101010011001, 16'd46804, 16'b1001010010101001);
	test_shift(16'b0101000011101111, 16'd8963, 16'b1110101000011101);
	test_shift(16'b1111000001011010, 16'd26410, 16'b0001011010111100);
	test_shift(16'b0000100010101001, 16'd3418, 16'b0010101001000010);
	test_shift(16'b1100000101110101, 16'd61106, 16'b0111000001011101);
	test_shift(16'b1011011101000101, 16'd30051, 16'b1011011011101000);
	test_shift(16'b0100000110100000, 16'd5046, 16'b1000000100000110);
	test_shift(16'b0111110110110101, 16'd27654, 16'b1101010111110110);
	test_shift(16'b1100110001100001, 16'd53779, 16'b0011100110001100);
	test_shift(16'b0110011100110001, 16'd31605, 16'b1000101100111001);
	test_shift(16'b1111111001101111, 16'd22960, 16'b1111111001101111);
	test_shift(16'b1111001110011011, 16'd31200, 16'b1111001110011011);
	test_shift(16'b0110111000011010, 16'd50761, 16'b0000110100110111);
	test_shift(16'b1101001100101000, 16'd28440, 16'b0010100011010011);
	test_shift(16'b1110111010100010, 16'd55415, 16'b0100010111011101);
	test_shift(16'b1000010011000000, 16'd47252, 16'b0000100001001100);
	test_shift(16'b0011000101110001, 16'd52334, 16'b1100010111000100);
	test_shift(16'b1010001011100110, 16'd17066, 16'b1011100110101000);
	test_shift(16'b0100110011101111, 16'd25350, 16'b1011110100110011);
	test_shift(16'b0111101011001011, 16'd47915, 16'b0101100101101111);
	test_shift(16'b1111011010001100, 16'd52284, 16'b0110100011001111);
	test_shift(16'b1101110011101111, 16'd64021, 16'b0111111011100111);
	test_shift(16'b0101001010011101, 16'd17295, 16'b1010010100111010);
	test_shift(16'b1010100100110100, 16'd39402, 16'b0100110100101010);
	test_shift(16'b1011101110101001, 16'd40905, 16'b1101010011011101);
	test_shift(16'b1101000110000100, 16'd37863, 16'b0000100110100011);
	test_shift(16'b0010101010110110, 16'd15991, 16'b0110110001010101);
	test_shift(16'b0101001110100110, 16'd5052, 16'b0011101001100101);
	test_shift(16'b1001101000000111, 16'd10318, 16'b0110100000011110);
	test_shift(16'b0000100000011000, 16'd34232, 16'b0001100000001000);
	test_shift(16'b1110001010100011, 16'd34700, 16'b0010101000111110);
	test_shift(16'b1001100101011001, 16'd6846, 16'b0110010101100110);
	test_shift(16'b0011000100010010, 16'd54847, 16'b0110001000100100);
	test_shift(16'b1000000011100000, 16'd6428, 16'b0000111000001000);
	test_shift(16'b1001001010101111, 16'd25563, 16'b0101010111110010);
	test_shift(16'b1101001100101110, 16'd65522, 16'b1011010011001011);
	test_shift(16'b1011001001110011, 16'd1865, 16'b0011100111011001);
	test_shift(16'b0110001010001001, 16'd1789, 16'b0001010001001011);
	test_shift(16'b1111001001100111, 16'd25035, 16'b0100110011111110);
	test_shift(16'b0101011101010011, 16'd52404, 16'b0011010101110101);
	test_shift(16'b0110001000111000, 16'd29088, 16'b0110001000111000);
	test_shift(16'b0110010011010000, 16'd16489, 16'b0110100000110010);
	test_shift(16'b1101010110100101, 16'd29851, 16'b1011010010111010);
	test_shift(16'b1010010110010101, 16'd20791, 16'b0010101101001011);
	test_shift(16'b1001011000101001, 16'd16122, 16'b1000101001100101);
	test_shift(16'b0001100000001101, 16'd10818, 16'b0100011000000011);
	test_shift(16'b1000001011000011, 16'd48761, 16'b0110000111000001);
	test_shift(16'b0000110100011011, 16'd14454, 16'b0110110000110100);
	test_shift(16'b1011011101101010, 16'd64524, 16'b0111011010101011);
	test_shift(16'b1001100101101010, 16'd8658, 16'b1010011001011010);
	test_shift(16'b1111111001110011, 16'd13779, 16'b0111111111001110);
	test_shift(16'b1011010111100001, 16'd39024, 16'b1011010111100001);
	test_shift(16'b1010100111001000, 16'd25884, 16'b1001110010001010);
	test_shift(16'b1100010110010110, 16'd53013, 16'b1011011000101100);
	test_shift(16'b1000101010110010, 16'd35570, 16'b1010001010101100);
	test_shift(16'b1100010111101111, 16'd16275, 16'b1111100010111101);
	test_shift(16'b0010111001101111, 16'd13729, 16'b1001011100110111);
	test_shift(16'b0001100001011010, 16'd49182, 16'b0110000101101000);
	test_shift(16'b0010101001111110, 16'd14747, 16'b0100111111000101);
	test_shift(16'b1001100011010001, 16'd7143, 16'b1010001100110001);
	test_shift(16'b0100000111001110, 16'd7578, 16'b0111001110010000);
	test_shift(16'b1010010101111110, 16'd7726, 16'b1001010111111010);
	test_shift(16'b1100000010111001, 16'd51652, 16'b1001110000001011);
	test_shift(16'b1000100100101000, 16'd40540, 16'b1001001010001000);
	test_shift(16'b0110100111000110, 16'd36148, 16'b0110011010011100);
	test_shift(16'b1100101010000111, 16'd63208, 16'b1000011111001010);
	test_shift(16'b1011111000101010, 16'd8045, 16'b1111000101010101);
	test_shift(16'b0100110000001111, 16'd45277, 16'b0110000001111010);
	test_shift(16'b1111111110111111, 16'd43344, 16'b1111111110111111);
	test_shift(16'b1011011010110101, 16'd39974, 16'b1101011011011010);
	test_shift(16'b1010110100000001, 16'd48430, 16'b1011010000000110);
	test_shift(16'b0011110001111000, 16'd31317, 16'b1100000111100011);
	test_shift(16'b1001000101110001, 16'd57730, 16'b0110010001011100);
	test_shift(16'b0001110100111110, 16'd38699, 16'b1010011111000011);
	test_shift(16'b0100010001110010, 16'd19666, 16'b1001000100011100);
	test_shift(16'b0000011101100011, 16'd39265, 16'b1000001110110001);
	test_shift(16'b1000000101011010, 16'd46610, 16'b1010000001010110);
	test_shift(16'b1101000010111011, 16'd15850, 16'b0010111011110100);
	test_shift(16'b0111010001110011, 16'd8311, 16'b1110011011101000);
	test_shift(16'b1000000000001111, 16'd9080, 16'b0000111110000000);
	test_shift(16'b0011110010010101, 16'd27634, 16'b0100111100100101);
	test_shift(16'b1100010101111111, 16'd50736, 16'b1100010101111111);
	test_shift(16'b0101001110010011, 16'd49568, 16'b0101001110010011);
	test_shift(16'b1100110111010101, 16'd22711, 16'b1010101110011011);
	test_shift(16'b1101011110110011, 16'd26170, 16'b1110110011110101);
	test_shift(16'b0001110111001000, 16'd51926, 16'b0010000001110111);
	test_shift(16'b0110000010010000, 16'd27851, 16'b0001001000001100);
	test_shift(16'b1100101011001001, 16'd35764, 16'b1001110010101100);
	test_shift(16'b0111011001111000, 16'd2661, 16'b1100001110110011);
	test_shift(16'b1101001001101000, 16'd25175, 16'b1101000110100100);
	test_shift(16'b1100101100011100, 16'd64918, 16'b0111001100101100);
	test_shift(16'b1101110010110000, 16'd27561, 16'b0101100001101110);
	test_shift(16'b1011100111101100, 16'd42369, 16'b0101110011110110);
	test_shift(16'b1010100010100110, 16'd18657, 16'b0101010001010011);
	test_shift(16'b0111110010011101, 16'd49185, 16'b1011111001001110);
	test_shift(16'b0000000001101010, 16'd33861, 16'b0101000000000011);
	test_shift(16'b0000100100110010, 16'd53642, 16'b0100110010000010);
	test_shift(16'b0001000110111100, 16'd51200, 16'b0001000110111100);
	test_shift(16'b0001000000010000, 16'd11174, 16'b0100000001000000);
	test_shift(16'b1010111111110101, 16'd53507, 16'b1011010111111110);
	test_shift(16'b0111001111001110, 16'd57267, 16'b1100111001111001);
	test_shift(16'b1000110010111100, 16'd13558, 16'b1111001000110010);
	test_shift(16'b1101100001101100, 16'd60880, 16'b1101100001101100);
	test_shift(16'b0100010110000010, 16'd54590, 16'b0001011000001001);
	test_shift(16'b0110110001111110, 16'd16510, 16'b1011000111111001);
	test_shift(16'b1111010100100001, 16'd35798, 16'b1000011111010100);
	test_shift(16'b1101001100001101, 16'd23917, 16'b1001100001101110);
	test_shift(16'b1110101011110000, 16'd35667, 16'b0001110101011110);
	test_shift(16'b0000001001001001, 16'd19894, 16'b0010010000001001);
	test_shift(16'b1100011100001110, 16'd54283, 16'b1110000111011000);
	test_shift(16'b1101011011111100, 16'd15218, 16'b0011010110111111);
	test_shift(16'b1111111101111101, 16'd4241, 16'b1111111110111110);
	test_shift(16'b0010101101101011, 16'd36772, 16'b1011001010110110);
	test_shift(16'b0011000000000000, 16'd46068, 16'b0000001100000000);
	test_shift(16'b0111100001100010, 16'd30235, 16'b0000110001001111);
	test_shift(16'b1100100101011010, 16'd62987, 16'b0010101101011001);
	test_shift(16'b1110100110010001, 16'd14480, 16'b1110100110010001);
	test_shift(16'b0000001010110111, 16'd12006, 16'b1101110000001010);
	test_shift(16'b1011101000110111, 16'd63559, 16'b0110111101110100);
	test_shift(16'b1110011101110011, 16'd62796, 16'b0111011100111110);
	test_shift(16'b0111110011100110, 16'd26399, 16'b1111100111001100);
	test_shift(16'b1000100110111001, 16'd24227, 16'b0011000100110111);
	test_shift(16'b1000110111010001, 16'd11388, 16'b1101110100011000);
	test_shift(16'b1110111101110011, 16'd35449, 16'b1011100111110111);
	test_shift(16'b1100101000100010, 16'd29956, 16'b0010110010100010);
	test_shift(16'b1001100100111100, 16'd58988, 16'b1001001111001001);
	test_shift(16'b1000101110011010, 16'd4168, 16'b1001101010001011);
	test_shift(16'b1001001001010100, 16'd24241, 16'b0100100100101010);
	test_shift(16'b1010010111000101, 16'd47524, 16'b0101101001011100);
	test_shift(16'b0001000010110111, 16'd16578, 16'b1100010000101101);
	test_shift(16'b1100000001110001, 16'd13307, 16'b0000111000111000);
	test_shift(16'b1010110011101000, 16'd26775, 16'b1101000101011001);
	test_shift(16'b0001010000101100, 16'd11324, 16'b0100001011000001);
	test_shift(16'b0010100000001010, 16'd54526, 16'b1010000000101000);
	test_shift(16'b1101101100000101, 16'd5350, 16'b0001011101101100);
	test_shift(16'b1111010000001110, 16'd35632, 16'b1111010000001110);
	test_shift(16'b0000111011001000, 16'd64503, 16'b1001000000011101);
	test_shift(16'b0010101000100001, 16'd41716, 16'b0001001010100010);
	test_shift(16'b0111110000000000, 16'd22952, 16'b0000000001111100);
	test_shift(16'b1111111000101100, 16'd1785, 16'b0001011001111111);
	test_shift(16'b0001111010000010, 16'd19095, 16'b0000010000111101);
	test_shift(16'b1111010110010010, 16'd5467, 16'b1011001001011110);
	test_shift(16'b1110100001111101, 16'd16964, 16'b1101111010000111);
	test_shift(16'b0001110001100001, 16'd63907, 16'b0010001110001100);
	test_shift(16'b0000100011100000, 16'd52799, 16'b0001000111000000);
	test_shift(16'b0101111101001110, 16'd9817, 16'b1010011100101111);
	test_shift(16'b1111010110000110, 16'd14920, 16'b1000011011110101);
	test_shift(16'b1010001101100000, 16'd58569, 16'b1011000001010001);
	test_shift(16'b1110100111000010, 16'd31833, 16'b1110000101110100);
	test_shift(16'b0101000011001011, 16'd14327, 16'b1001011010100001);
	test_shift(16'b0100111001010110, 16'd54834, 16'b1001001110010101);
	test_shift(16'b0011000011001101, 16'd57579, 16'b0001100110100110);
	test_shift(16'b0000010000001111, 16'd49968, 16'b0000010000001111);
	test_shift(16'b0000101100000000, 16'd33566, 16'b0010110000000000);
	test_shift(16'b0011000000110110, 16'd44209, 16'b0001100000011011);
	test_shift(16'b1100010010001001, 16'd62677, 16'b0100111000100100);
	test_shift(16'b1010111111001000, 16'd61132, 16'b1111110010001010);
	test_shift(16'b1001101001101110, 16'd65143, 16'b1101110100110100);
	test_shift(16'b1011101000000111, 16'd31336, 16'b0000011110111010);
	test_shift(16'b1000101001110000, 16'd29867, 16'b0100111000010001);
	test_shift(16'b1111010100100101, 16'd11205, 16'b0010111110101001);
	test_shift(16'b1010000101001010, 16'd41581, 16'b0000101001010101);
	test_shift(16'b1000111001010110, 16'd46281, 16'b0010101101000111);
	test_shift(16'b1100010100100001, 16'd10119, 16'b0100001110001010);
	test_shift(16'b0101100010110010, 16'd10884, 16'b0010010110001011);
	test_shift(16'b0110110000010100, 16'd25753, 16'b0000101000110110);
	test_shift(16'b1001001110110010, 16'd38391, 16'b0110010100100111);
	test_shift(16'b0111001011011010, 16'd21190, 16'b0110100111001011);
	test_shift(16'b1110011101111011, 16'd28143, 16'b1100111011110111);
	test_shift(16'b0011010100111011, 16'd43696, 16'b0011010100111011);
	test_shift(16'b1010111010001000, 16'd38967, 16'b0001000101011101);
	test_shift(16'b1100011110111101, 16'd38828, 16'b0111101111011100);
	test_shift(16'b1000100001001110, 16'd16722, 16'b1010001000010011);
	test_shift(16'b0100110111100101, 16'd9679, 16'b1001101111001010);
	test_shift(16'b0001001011000010, 16'd33202, 16'b1000010010110000);
	test_shift(16'b1000001101100111, 16'd44892, 16'b0011011001111000);
	test_shift(16'b1000111010110100, 16'd39270, 16'b1101001000111010);
	test_shift(16'b1001000100011011, 16'd5735, 16'b0011011100100010);
	test_shift(16'b1101100011001011, 16'd14562, 16'b1111011000110010);
	test_shift(16'b0110101000101011, 16'd40711, 16'b0101011011010100);
	test_shift(16'b1111111111101100, 16'd12685, 16'b1111111101100111);
	test_shift(16'b1010011010001011, 16'd15399, 16'b0001011101001101);
	test_shift(16'b0111100101100110, 16'd11129, 16'b1011001100111100);
	test_shift(16'b0000110011110011, 16'd17732, 16'b0011000011001111);
	test_shift(16'b1010100000010100, 16'd16642, 16'b0010101000000101);
	test_shift(16'b0010110111010010, 16'd1717, 16'b1001000101101110);
	test_shift(16'b0001100111101000, 16'd60046, 16'b0110011110100000);
	test_shift(16'b0110101000100110, 16'd50548, 16'b0110011010100010);
	test_shift(16'b0011100001100011, 16'd8694, 16'b1000110011100001);
	test_shift(16'b1001010101011011, 16'd37333, 16'b1101110010101010);
	test_shift(16'b1000101101000000, 16'd11633, 16'b0100010110100000);
	test_shift(16'b0101011011100000, 16'd21187, 16'b0000101011011100);
	test_shift(16'b0101100011010011, 16'd35601, 16'b1010110001101001);
	test_shift(16'b0000010110010100, 16'd41701, 16'b1010000000101100);
	test_shift(16'b0011011001100010, 16'd37231, 16'b0110110011000100);
	test_shift(16'b0011110110011100, 16'd25604, 16'b1100001111011001);
	test_shift(16'b1011010111011000, 16'd11579, 16'b1011101100010110);
	test_shift(16'b1110010010011011, 16'd42134, 16'b0110111110010010);
	test_shift(16'b1001011000010011, 16'd16561, 16'b1100101100001001);
	test_shift(16'b0001010010110001, 16'd31855, 16'b0010100101100010);
	test_shift(16'b1111010111101011, 16'd64427, 16'b1011110101111110);
	test_shift(16'b0101001011110101, 16'd41429, 16'b1010101010010111);
	test_shift(16'b1101101000101101, 16'd27028, 16'b1101110110100010);
	test_shift(16'b0000111000011011, 16'd6887, 16'b0011011000011100);
	test_shift(16'b0000001111000001, 16'd45601, 16'b1000000111100000);
	test_shift(16'b0001111100000110, 16'd34483, 16'b1100001111100000);
	test_shift(16'b1001010111001101, 16'd62094, 16'b0101011100110110);
	test_shift(16'b0110001011001110, 16'd56943, 16'b1100010110011100);
	test_shift(16'b0111111111010010, 16'd17261, 16'b1111111010010011);
	test_shift(16'b0001001110000100, 16'd32339, 16'b1000001001110000);
	test_shift(16'b0000001100001001, 16'd62917, 16'b0100100000011000);
	test_shift(16'b0000011010001000, 16'd11365, 16'b0100000000110100);
	test_shift(16'b1101111000011000, 16'd30202, 16'b1000011000110111);
	test_shift(16'b1100110011010101, 16'd45286, 16'b0101011100110011);
	test_shift(16'b1111111111010011, 16'd54188, 16'b1111110100111111);
	test_shift(16'b1110100111111101, 16'd51490, 16'b0111101001111111);
	test_shift(16'b1011011011110000, 16'd41648, 16'b1011011011110000);
	test_shift(16'b1011101001100111, 16'd38079, 16'b0111010011001111);
	test_shift(16'b0111101000000101, 16'd59954, 16'b0101111010000001);
	test_shift(16'b0011000011110110, 16'd231, 16'b1110110001100001);
	test_shift(16'b0000011000100111, 16'd23484, 16'b0110001001110000);
	test_shift(16'b1110100111101110, 16'd39754, 16'b0111101110111010);
	test_shift(16'b0000011010101011, 16'd36196, 16'b1011000001101010);
	test_shift(16'b1100001100110101, 16'd3459, 16'b1011100001100110);
	test_shift(16'b0111100111111100, 16'd39064, 16'b1111110001111001);
	test_shift(16'b1110100101100111, 16'd63273, 16'b1011001111110100);
	test_shift(16'b0000010000110001, 16'd6024, 16'b0011000100000100);
	test_shift(16'b0101001110001000, 16'd48352, 16'b0101001110001000);
	test_shift(16'b1000111111000111, 16'd9873, 16'b1100011111100011);
	test_shift(16'b0000011001011100, 16'd27799, 16'b1011100000001100);
	test_shift(16'b0110001111011010, 16'd16174, 16'b1000111101101001);
	test_shift(16'b0101111011110010, 16'd52368, 16'b0101111011110010);
	test_shift(16'b0101011100100100, 16'd49963, 16'b1110010010001010);
	test_shift(16'b0100001101100001, 16'd16688, 16'b0100001101100001);
	test_shift(16'b0101101101000010, 16'd62373, 16'b0001001011011010);
	test_shift(16'b1101110000100010, 16'd15476, 16'b0010110111000010);
	test_shift(16'b0000000011101010, 16'd51152, 16'b0000000011101010);
	test_shift(16'b1100111000001101, 16'd1809, 16'b1110011100000110);
	test_shift(16'b0100010100001110, 16'd39576, 16'b0000111001000101);
	test_shift(16'b1011110000001101, 16'd34768, 16'b1011110000001101);
	test_shift(16'b1000100010100001, 16'd36294, 16'b1000011000100010);
	test_shift(16'b0000100010111111, 16'd6603, 16'b0001011111100001);
	test_shift(16'b0010000110111100, 16'd6204, 16'b0001101111000010);
	test_shift(16'b0001010111111010, 16'd63117, 16'b1010111111010000);
	test_shift(16'b1001011001000000, 16'd23552, 16'b1001011001000000);
	test_shift(16'b1101111110010110, 16'd15362, 16'b1011011111100101);
	test_shift(16'b0010110001000000, 16'd38392, 16'b0100000000101100);
	test_shift(16'b1111010010100000, 16'd3628, 16'b0100101000001111);
	test_shift(16'b0100001010001011, 16'd42677, 16'b0101101000010100);
	test_shift(16'b1011101000110110, 16'd52451, 16'b1101011101000110);
	test_shift(16'b0000010010000001, 16'd51746, 16'b0100000100100000);
	test_shift(16'b1000100100001000, 16'd47585, 16'b0100010010000100);
	test_shift(16'b1110000011111100, 16'd56312, 16'b1111110011100000);
	test_shift(16'b0001010000011011, 16'd16324, 16'b1011000101000001);
	test_shift(16'b0100011111100100, 16'd16541, 16'b0011111100100010);
	test_shift(16'b0110111110111001, 16'd32442, 16'b1110111001011011);
	test_shift(16'b0010001111010001, 16'd18616, 16'b1101000100100011);
	test_shift(16'b0110001000001011, 16'd35849, 16'b0000010110110001);
	test_shift(16'b0001001101101001, 16'd30733, 16'b1001101101001000);
	test_shift(16'b1100001110100001, 16'd19312, 16'b1100001110100001);
	test_shift(16'b0001100110011101, 16'd37643, 16'b0011001110100011);
	test_shift(16'b1001100011111010, 16'd27608, 16'b1111101010011000);
	test_shift(16'b0110001000110101, 16'd38125, 16'b0001000110101011);
	test_shift(16'b0100101001101011, 16'd21653, 16'b0101101001010011);
	test_shift(16'b0000101010110100, 16'd7075, 16'b1000000101010110);
	test_shift(16'b1100111000011001, 16'd20852, 16'b1001110011100001);
	test_shift(16'b1100101011110100, 16'd42730, 16'b1011110100110010);
	test_shift(16'b0101010010011110, 16'd59694, 16'b0101001001111001);
	test_shift(16'b1100111001001100, 16'd14496, 16'b1100111001001100);
	test_shift(16'b1001100111101011, 16'd38136, 16'b1110101110011001);
	test_shift(16'b0111011101000011, 16'd9264, 16'b0111011101000011);
	test_shift(16'b0010100101000001, 16'd209, 16'b1001010010100000);
	test_shift(16'b0001000101111110, 16'd3830, 16'b1111100001000101);
	test_shift(16'b1101011000010000, 16'd58329, 16'b0000100001101011);
	test_shift(16'b1010111110110100, 16'd48043, 16'b1111011010010101);
	test_shift(16'b1100110010011001, 16'd30188, 16'b1100100110011100);
	test_shift(16'b1000010110111101, 16'd37289, 16'b1101111011000010);
	test_shift(16'b0000110100101011, 16'd59034, 16'b0100101011000011);
	test_shift(16'b1111011010010011, 16'd62847, 16'b1110110100100111);
	test_shift(16'b1110011011000010, 16'd44090, 16'b1011000010111001);
	test_shift(16'b0101101000111111, 16'd45534, 16'b0110100011111101);
	test_shift(16'b1101111000001101, 16'd3575, 16'b0001101110111100);
	test_shift(16'b0000001001001010, 16'd26148, 16'b1010000000100100);
	test_shift(16'b0111110101101010, 16'd13563, 16'b1010110101001111);
	test_shift(16'b0101011011011010, 16'd47389, 16'b1011011011010010);
	test_shift(16'b1011110011100111, 16'd59865, 16'b0111001111011110);
	test_shift(16'b1101000100001010, 16'd13144, 16'b0000101011010001);
	test_shift(16'b1001011011010011, 16'd52964, 16'b0011100101101101);
	test_shift(16'b0111100010010101, 16'd28468, 16'b0101011110001001);
	test_shift(16'b0001101110111111, 16'd34905, 16'b1101111110001101);
	test_shift(16'b1000010001010010, 16'd13476, 16'b0010100001000101);
	test_shift(16'b0001010001110011, 16'd2761, 16'b0011100110001010);
	test_shift(16'b0001100000110101, 16'd5906, 16'b0100011000001101);
	test_shift(16'b1100111010101000, 16'd29364, 16'b1000110011101010);
	test_shift(16'b1101001111110100, 16'd35784, 16'b1111010011010011);
	test_shift(16'b1100000101000011, 16'd16009, 16'b1010000111100000);
	test_shift(16'b0110110101111001, 16'd41408, 16'b0110110101111001);
	test_shift(16'b0000110001111000, 16'd56221, 16'b0110001111000000);
	test_shift(16'b1010000011011010, 16'd50575, 16'b0100000110110101);
	test_shift(16'b1101001111010011, 16'd47236, 16'b0011110100111101);
	test_shift(16'b0000100010000111, 16'd21614, 16'b0010001000011100);
	test_shift(16'b0001010100110000, 16'd52653, 16'b1010100110000000);
	test_shift(16'b0010000111110011, 16'd45278, 16'b1000011111001100);
	test_shift(16'b0011010010110110, 16'd28272, 16'b0011010010110110);
	test_shift(16'b1011110011000000, 16'd38104, 16'b1100000010111100);
	test_shift(16'b1010110101111111, 16'd42156, 16'b1101011111111010);
	test_shift(16'b0101111001001111, 16'd21371, 16'b1100100111101011);
	test_shift(16'b0011010101110101, 16'd60915, 16'b1010011010101110);
	test_shift(16'b0011000100101010, 16'd39434, 16'b0100101010001100);
	test_shift(16'b0100000011011001, 16'd137, 16'b0110110010100000);
	test_shift(16'b0111000101001111, 16'd23487, 16'b1110001010011110);
	test_shift(16'b1111000010110100, 16'd44645, 16'b1010011110000101);
	test_shift(16'b0110111110000101, 16'd63214, 16'b1011111000010101);
	test_shift(16'b1000001000100010, 16'd44066, 16'b1010000010001000);
	test_shift(16'b0000111101000100, 16'd51357, 16'b0111101000100000);
	test_shift(16'b1010000001011010, 16'd25060, 16'b1010101000000101);
	test_shift(16'b1100101110100001, 16'd48407, 16'b0100001110010111);
	test_shift(16'b0101010001110011, 16'd23513, 16'b0011100110101010);
	test_shift(16'b0110000010101100, 16'd37239, 16'b0101100011000001);
	test_shift(16'b1110111101000101, 16'd2554, 16'b1101000101111011);
	test_shift(16'b0001100101100000, 16'd13975, 16'b1100000000110010);
	test_shift(16'b0011011001001000, 16'd55689, 16'b0010010000011011);
	test_shift(16'b1100101110110101, 16'd21822, 16'b0010111011010111);
	test_shift(16'b1000010100100101, 16'd38223, 16'b0000101001001011);
	test_shift(16'b1010100111010101, 16'd33093, 16'b1010110101001110);
	test_shift(16'b1000010001011011, 16'd41796, 16'b1011100001000101);
	test_shift(16'b1010111100011010, 16'd41755, 16'b1110001101010101);
	test_shift(16'b0011000011100111, 16'd64798, 16'b1100001110011100);
	test_shift(16'b1001001010111010, 16'd6353, 16'b0100100101011101);
	test_shift(16'b1010100100100001, 16'd25004, 16'b1001001000011010);
	test_shift(16'b0010110100000100, 16'd58589, 16'b0110100000100001);
	test_shift(16'b0111110101100111, 16'd2699, 16'b1010110011101111);
	test_shift(16'b0100010011011001, 16'd35478, 16'b0110010100010011);
	test_shift(16'b0000011001101000, 16'd43479, 16'b1101000000001100);
	test_shift(16'b0110101000000111, 16'd1925, 16'b0011101101010000);
	test_shift(16'b1110010111110010, 16'd13108, 16'b0010111001011111);
	test_shift(16'b1110000110011010, 16'd3055, 16'b1100001100110101);
	test_shift(16'b1000011011011001, 16'd63907, 16'b0011000011011011);
	test_shift(16'b1110111011110100, 16'd21604, 16'b0100111011101111);
	test_shift(16'b1110110000010000, 16'd62539, 16'b1000001000011101);
	test_shift(16'b0000001111001111, 16'd52295, 16'b1001111000000111);
	test_shift(16'b1000011011111000, 16'd2675, 16'b0001000011011111);
	test_shift(16'b1010010010011111, 16'd17104, 16'b1010010010011111);
	test_shift(16'b0101010010110101, 16'd42071, 16'b0110101010101001);
	test_shift(16'b1110010011001110, 16'd39944, 16'b1100111011100100);
	test_shift(16'b1010100010011001, 16'd7445, 16'b1100110101000100);
	test_shift(16'b0110011111100110, 16'd36363, 16'b1111110011001100);
	test_shift(16'b0101000111111001, 16'd50374, 16'b1110010101000111);
	test_shift(16'b0101111110001101, 16'd33576, 16'b1000110101011111);
	test_shift(16'b1000011010001100, 16'd27018, 16'b1010001100100001);
	test_shift(16'b1010111111011000, 16'd56082, 16'b0010101111110110);
	test_shift(16'b0101101101101010, 16'd35422, 16'b0110110110101001);
	test_shift(16'b0100101000001011, 16'd45660, 16'b1010000010110100);
	test_shift(16'b0110011101101100, 16'd38618, 16'b1101101100011001);
	test_shift(16'b1011101110111101, 16'd18565, 16'b1110110111011101);
	test_shift(16'b1101001111101101, 16'd61630, 16'b0100111110110111);
	test_shift(16'b1001100000101100, 16'd49364, 16'b1100100110000010);
	test_shift(16'b0101110001001111, 16'd28645, 16'b0111101011100010);
	test_shift(16'b1100011101011111, 16'd54481, 16'b1110001110101111);
	test_shift(16'b0100100000100000, 16'd47625, 16'b0001000000100100);
	test_shift(16'b1011010001001000, 16'd8569, 16'b0010010001011010);
	test_shift(16'b1001001001111000, 16'd22970, 16'b1001111000100100);
	test_shift(16'b0101110001111011, 16'd33733, 16'b1101101011100011);
	test_shift(16'b0110001111101001, 16'd531, 16'b0010110001111101);
	test_shift(16'b0000011000001011, 16'd43341, 16'b0011000001011000);
	test_shift(16'b1110011010111100, 16'd13863, 16'b0111100111001101);
	test_shift(16'b1000000101010100, 16'd53053, 16'b0000101010100100);
	test_shift(16'b1001100111110100, 16'd35288, 16'b1111010010011001);
	test_shift(16'b1110001011111100, 16'd37022, 16'b1000101111110011);
	test_shift(16'b1111110110100111, 16'd15613, 16'b1110110100111111);
	test_shift(16'b1110010001101111, 16'd872, 16'b0110111111100100);
	test_shift(16'b0011001110100100, 16'd27232, 16'b0011001110100100);
	test_shift(16'b0011011110011010, 16'd13734, 16'b0110100011011110);
	test_shift(16'b1000010100001011, 16'd50584, 16'b0000101110000101);
	test_shift(16'b0000000101111011, 16'd33281, 16'b1000000010111101);
	test_shift(16'b1000101111110000, 16'd15827, 16'b0001000101111110);
	test_shift(16'b1100101100001001, 16'd65466, 16'b1100001001110010);
	test_shift(16'b1010101110000100, 16'd5390, 16'b1010111000010010);
	test_shift(16'b1010011100111111, 16'd56427, 16'b1110011111110100);
	test_shift(16'b0100100001111110, 16'd64300, 16'b1000011111100100);
	test_shift(16'b1100111010000000, 16'd31896, 16'b1000000011001110);
	test_shift(16'b0111111101110100, 16'd53318, 16'b1101000111111101);

    $display("SUCCESS :: FINISH CALLED FROM END OF FILE!");
    $finish;

end


endmodule

