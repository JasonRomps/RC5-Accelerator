`define K_size 128 // Key size (PARAMETER)
`define W_size 16 // word size (PARAMETER)
`define T 26 // 2*(number of rounds + 1)

// COMMENT THIS DEFINE OUT FOR ALL 10,000 TEST CASES!!!!
`define FULL

`timescale 1ns / 1ps
module key_tb;

logic start;
logic clk;
logic rst;
logic[`K_size-1:0] key;
logic[`W_size-1:0] sub [`T];
logic ready;

keygen Keygen(.*);

default clocking ckb @(posedge clk);
    input sub, ready;
    output rst, key, start;
endclocking

always begin
    clk = 1'b0;
    #1;
    clk = 1'b1;
    #1;
end

task reset();
    rst <= 1;
    ##1;
    rst <= 0;
    ##1;
endtask

task test_expansion(logic[`K_size-1:0] test_key, logic [`W_size-1:0] test_subkey [`T]);
    key <= test_key;
    start <= 1;
    ##1;

    start <= 0;

    while(~ready) begin
        ##1;
    end

    for(int i = 0; i < `T; i++) begin
        assert(test_subkey[i] == sub[i])
            else begin
                $error("Bad Subkey Value: 0x%x at position %0d, should be 0x%x", sub[i], i, test_subkey[i]);
                $finish;
            end
    end
endtask

initial begin
    $fsdbDumpfile("dump.fsdb");
	$fsdbDumpvars(0, "+all");
    key <= 0;
    rst <= 0;
    start <= 0;

    #2;

    reset();

	test_expansion(128'hff6437a2d84a29d2692a5848177da494, {16'd58031, 16'd55734, 16'd39026, 16'd34949, 16'd44626, 16'd26908, 16'd30331, 16'd9073, 16'd14534, 16'd8516, 16'd51677, 16'd48415, 16'd37976, 16'd10818, 16'd50175, 16'd3407, 16'd64641, 16'd50058, 16'd35322, 16'd8098, 16'd7148, 16'd39892, 16'd62986, 16'd40991, 16'd37102, 16'd15450});
	test_expansion(128'h5db04132e8875cce57b0d8d3b50d15dc, {16'd44782, 16'd1932, 16'd40049, 16'd42159, 16'd8711, 16'd60465, 16'd11744, 16'd22533, 16'd3089, 16'd32921, 16'd31501, 16'd28196, 16'd43557, 16'd53578, 16'd14750, 16'd56645, 16'd44849, 16'd56293, 16'd51715, 16'd60018, 16'd59739, 16'd36058, 16'd4932, 16'd2481, 16'd58364, 16'd64461});
	test_expansion(128'h995dad14e730c7c877076770b635e622, {16'd36021, 16'd36148, 16'd16253, 16'd38450, 16'd30131, 16'd1570, 16'd57838, 16'd51666, 16'd33874, 16'd40434, 16'd17844, 16'd5254, 16'd50710, 16'd58262, 16'd9333, 16'd48966, 16'd455, 16'd35267, 16'd14254, 16'd36809, 16'd50441, 16'd30566, 16'd54158, 16'd14507, 16'd33554, 16'd8743});
	test_expansion(128'ha474e2eb1ed2b8b4f2fb5a5e4a4470a9, {16'd48493, 16'd15361, 16'd8111, 16'd25986, 16'd44216, 16'd47784, 16'd36247, 16'd22111, 16'd29307, 16'd22810, 16'd62633, 16'd40133, 16'd42817, 16'd44493, 16'd33692, 16'd38110, 16'd5689, 16'd49855, 16'd64669, 16'd45120, 16'd7903, 16'd49993, 16'd9787, 16'd59473, 16'd13379, 16'd8491});
	test_expansion(128'h1be82cdcc3a2fd6f44520d427501e175, {16'd1868, 16'd7044, 16'd32642, 16'd3273, 16'd33246, 16'd47455, 16'd37089, 16'd47072, 16'd31832, 16'd63729, 16'd15097, 16'd44849, 16'd52354, 16'd14502, 16'd2140, 16'd8714, 16'd59841, 16'd6768, 16'd42547, 16'd4546, 16'd22258, 16'd34556, 16'd12981, 16'd19021, 16'd48073, 16'd20931});
	test_expansion(128'h283b92a0463442508e682818248de078, {16'd1388, 16'd12219, 16'd29107, 16'd38456, 16'd3758, 16'd12168, 16'd4235, 16'd61023, 16'd62475, 16'd14896, 16'd29826, 16'd25852, 16'd9928, 16'd54836, 16'd15684, 16'd42594, 16'd6835, 16'd36566, 16'd48747, 16'd36323, 16'd27660, 16'd37206, 16'd40840, 16'd14404, 16'd56395, 16'd21711});
	test_expansion(128'ha30f563cb673a3c897d91ac2bf24d217, {16'd41196, 16'd53778, 16'd22584, 16'd17684, 16'd13120, 16'd48182, 16'd46699, 16'd43805, 16'd41209, 16'd63110, 16'd27174, 16'd20484, 16'd49280, 16'd39554, 16'd10963, 16'd40749, 16'd60197, 16'd15715, 16'd59934, 16'd51105, 16'd41046, 16'd20871, 16'd42061, 16'd48338, 16'd14283, 16'd38837});
	test_expansion(128'h53607407f7790ab20c6732db12da5b99, {16'd25029, 16'd11553, 16'd47383, 16'd34348, 16'd14314, 16'd11300, 16'd6455, 16'd3950, 16'd6355, 16'd26957, 16'd32332, 16'd42299, 16'd50629, 16'd65216, 16'd36896, 16'd49325, 16'd58006, 16'd21792, 16'd55964, 16'd17916, 16'd7043, 16'd32951, 16'd2560, 16'd51863, 16'd28170, 16'd16811});
	test_expansion(128'h7005bc0bd7f3b68a2a44ea3b2896a6d1, {16'd62281, 16'd1432, 16'd25842, 16'd1778, 16'd20143, 16'd15557, 16'd39216, 16'd15198, 16'd49538, 16'd61088, 16'd27365, 16'd10159, 16'd26063, 16'd8051, 16'd6815, 16'd7326, 16'd47940, 16'd12975, 16'd6664, 16'd203, 16'd45025, 16'd27782, 16'd46589, 16'd36818, 16'd42276, 16'd32989});
	test_expansion(128'hd15df1bb1ed32c4f62ea8ee3ace8c7f0, {16'd51994, 16'd22304, 16'd17190, 16'd26788, 16'd14094, 16'd64805, 16'd7986, 16'd45294, 16'd53714, 16'd54566, 16'd15859, 16'd913, 16'd49641, 16'd10303, 16'd40974, 16'd27692, 16'd58944, 16'd38172, 16'd40233, 16'd50581, 16'd20000, 16'd42496, 16'd65051, 16'd8068, 16'd52138, 16'd29127});
	
	`ifdef FULL
	
	test_expansion(128'he4bd49bfefe240d8c699f86709673ee8, {16'd13158, 16'd12368, 16'd36588, 16'd9161, 16'd32625, 16'd29116, 16'd47353, 16'd53641, 16'd50120, 16'd40213, 16'd20206, 16'd10459, 16'd44500, 16'd61389, 16'd14298, 16'd59599, 16'd59504, 16'd58231, 16'd396, 16'd65192, 16'd40741, 16'd56378, 16'd25966, 16'd7390, 16'd24379, 16'd44075});
	test_expansion(128'hf0c92f7b53872d11a5121159ff74bf18, {16'd42101, 16'd53252, 16'd13984, 16'd58075, 16'd8420, 16'd8742, 16'd31229, 16'd18768, 16'd46368, 16'd36623, 16'd13771, 16'd36881, 16'd11443, 16'd21945, 16'd33116, 16'd29317, 16'd32417, 16'd31175, 16'd42039, 16'd15017, 16'd20377, 16'd13139, 16'd46568, 16'd39019, 16'd37443, 16'd61299});
	test_expansion(128'h931e8601faefe2492aa7a5ba7239f26e, {16'd17273, 16'd16054, 16'd21383, 16'd60797, 16'd30891, 16'd6357, 16'd55000, 16'd7670, 16'd48468, 16'd57414, 16'd62164, 16'd57438, 16'd4904, 16'd25906, 16'd716, 16'd173, 16'd11913, 16'd61588, 16'd25077, 16'd63192, 16'd51626, 16'd58812, 16'd39051, 16'd33545, 16'd28671, 16'd10065});
	test_expansion(128'hec7655ad487e5677bcd806bf16327993, {16'd42182, 16'd64214, 16'd45867, 16'd3031, 16'd58742, 16'd3746, 16'd34171, 16'd6264, 16'd55998, 16'd50014, 16'd55567, 16'd32873, 16'd42546, 16'd56711, 16'd62962, 16'd10975, 16'd13938, 16'd43885, 16'd59413, 16'd40181, 16'd61100, 16'd19543, 16'd54099, 16'd42447, 16'd57951, 16'd60533});
	test_expansion(128'h18ea18a147084b2570a4ff911bc14480, {16'd5437, 16'd47909, 16'd58120, 16'd12358, 16'd60024, 16'd26663, 16'd49033, 16'd19089, 16'd1823, 16'd59979, 16'd59966, 16'd42122, 16'd3308, 16'd8243, 16'd24629, 16'd62982, 16'd44715, 16'd9862, 16'd19798, 16'd27539, 16'd29699, 16'd30331, 16'd2649, 16'd12537, 16'd34063, 16'd42521});
	test_expansion(128'h2f19097c2d1ea767dd140b328d56efcc, {16'd41961, 16'd64341, 16'd11865, 16'd63208, 16'd34994, 16'd64377, 16'd33234, 16'd16172, 16'd14521, 16'd64549, 16'd15076, 16'd53324, 16'd33502, 16'd10611, 16'd58969, 16'd58558, 16'd36278, 16'd46582, 16'd29847, 16'd59398, 16'd46073, 16'd41490, 16'd2319, 16'd40644, 16'd50635, 16'd31361});
	test_expansion(128'h49a40f5fbaf6e9b8f51c3ce7fed67649, {16'd35010, 16'd52734, 16'd20880, 16'd54225, 16'd46885, 16'd61752, 16'd5209, 16'd24417, 16'd19821, 16'd47075, 16'd22036, 16'd32988, 16'd12573, 16'd25010, 16'd48357, 16'd56020, 16'd28678, 16'd7408, 16'd52101, 16'd29582, 16'd64419, 16'd47689, 16'd27951, 16'd4429, 16'd51394, 16'd7128});
	test_expansion(128'hfb62038d01d6f90aad536ba17e306d61, {16'd63748, 16'd42270, 16'd36455, 16'd40100, 16'd6997, 16'd54024, 16'd21146, 16'd55598, 16'd56836, 16'd21214, 16'd49170, 16'd16666, 16'd49731, 16'd29161, 16'd46943, 16'd2066, 16'd23118, 16'd17047, 16'd3508, 16'd54083, 16'd56818, 16'd13543, 16'd9632, 16'd42815, 16'd15723, 16'd58160});
	test_expansion(128'h0f5902274cd86b852c6d03a395aee561, {16'd48457, 16'd54127, 16'd61599, 16'd22749, 16'd16986, 16'd14417, 16'd6464, 16'd2234, 16'd48382, 16'd52610, 16'd43710, 16'd63690, 16'd35530, 16'd27204, 16'd38271, 16'd14940, 16'd12856, 16'd810, 16'd58502, 16'd10215, 16'd61827, 16'd42562, 16'd7052, 16'd18184, 16'd36088, 16'd34064});
	test_expansion(128'hf6b1e7546a03ede5e8d4610b09df5577, {16'd42239, 16'd37999, 16'd50967, 16'd47703, 16'd42219, 16'd963, 16'd751, 16'd38929, 16'd24286, 16'd42674, 16'd50660, 16'd12889, 16'd59154, 16'd53783, 16'd342, 16'd62704, 16'd63020, 16'd38048, 16'd54604, 16'd41658, 16'd16677, 16'd3215, 16'd55092, 16'd23216, 16'd53324, 16'd37375});
	test_expansion(128'h8ab2774758e7df79b45ee17558e51db7, {16'd38561, 16'd9068, 16'd27262, 16'd20104, 16'd52643, 16'd15381, 16'd42856, 16'd43972, 16'd40201, 16'd32978, 16'd54550, 16'd50441, 16'd13390, 16'd51838, 16'd43599, 16'd25213, 16'd10439, 16'd19968, 16'd62667, 16'd44894, 16'd55918, 16'd58112, 16'd10618, 16'd2271, 16'd34379, 16'd34795});
	test_expansion(128'hfa46d3f2b0af87fb5ec0daf5e7ee6fce, {16'd64576, 16'd17877, 16'd33235, 16'd53669, 16'd43478, 16'd1341, 16'd58747, 16'd34197, 16'd63228, 16'd11752, 16'd46700, 16'd11160, 16'd15318, 16'd13840, 16'd44203, 16'd48997, 16'd38375, 16'd28882, 16'd56576, 16'd57572, 16'd61035, 16'd33865, 16'd12728, 16'd9713, 16'd56062, 16'd25933});
	test_expansion(128'heb7983e38aa2321c4b42902e48409813, {16'd3792, 16'd12504, 16'd41309, 16'd24384, 16'd2786, 16'd45838, 16'd3588, 16'd55279, 16'd11181, 16'd64838, 16'd26212, 16'd23005, 16'd38023, 16'd6178, 16'd11050, 16'd62610, 16'd42291, 16'd43649, 16'd5214, 16'd5483, 16'd14198, 16'd223, 16'd10802, 16'd39322, 16'd25561, 16'd56249});
	test_expansion(128'hd9c26c06b5a11e65a577aee686fd3384, {16'd55340, 16'd39795, 16'd46180, 16'd37744, 16'd2252, 16'd52668, 16'd62864, 16'd21352, 16'd43461, 16'd50391, 16'd59574, 16'd22132, 16'd21942, 16'd48696, 16'd6551, 16'd5448, 16'd5524, 16'd11120, 16'd47228, 16'd37755, 16'd1177, 16'd17668, 16'd59707, 16'd47983, 16'd44259, 16'd28362});
	test_expansion(128'h33b980e4a7c0e8db7a0604ea3e681fab, {16'd7003, 16'd8739, 16'd36631, 16'd5635, 16'd54930, 16'd61378, 16'd48145, 16'd37520, 16'd40308, 16'd17956, 16'd46140, 16'd58592, 16'd33637, 16'd8571, 16'd17506, 16'd28950, 16'd7867, 16'd5987, 16'd49705, 16'd5019, 16'd39921, 16'd38386, 16'd56694, 16'd50717, 16'd31090, 16'd23428});
	test_expansion(128'hd8f1c51e1b857e1ed5bc550678107fd6, {16'd40527, 16'd34770, 16'd4332, 16'd37431, 16'd61374, 16'd8898, 16'd17295, 16'd55886, 16'd1742, 16'd853, 16'd38333, 16'd22247, 16'd49873, 16'd2500, 16'd55091, 16'd53988, 16'd19814, 16'd53010, 16'd64409, 16'd9996, 16'd54316, 16'd25923, 16'd7556, 16'd43192, 16'd61419, 16'd53683});
	test_expansion(128'h95756bc3cbe9a9b17bd67e5b6733423f, {16'd22244, 16'd12210, 16'd28970, 16'd5404, 16'd18772, 16'd30467, 16'd9334, 16'd18792, 16'd27842, 16'd54259, 16'd18504, 16'd12780, 16'd42184, 16'd43680, 16'd12888, 16'd2311, 16'd8659, 16'd30408, 16'd45572, 16'd63517, 16'd5676, 16'd16335, 16'd56975, 16'd20788, 16'd36084, 16'd30919});
	test_expansion(128'h66b0e7a3dfb571190ae283b56d20b9a9, {16'd39232, 16'd62227, 16'd49262, 16'd855, 16'd47122, 16'd49294, 16'd16242, 16'd16443, 16'd27714, 16'd18505, 16'd26056, 16'd3961, 16'd50021, 16'd57171, 16'd50390, 16'd17198, 16'd10283, 16'd30379, 16'd54065, 16'd18052, 16'd38371, 16'd10965, 16'd36234, 16'd57436, 16'd11417, 16'd15107});
	test_expansion(128'h98e5303347ddc3a62fe50c9697bdb1d7, {16'd15839, 16'd33193, 16'd9041, 16'd45976, 16'd56263, 16'd5310, 16'd36874, 16'd61224, 16'd23078, 16'd11223, 16'd34390, 16'd44316, 16'd52119, 16'd55532, 16'd45329, 16'd64468, 16'd49755, 16'd21502, 16'd53291, 16'd51745, 16'd49768, 16'd60144, 16'd46594, 16'd36641, 16'd4840, 16'd20789});
	test_expansion(128'hfb4ffb611799301f82eb6bdbe9d932cb, {16'd25927, 16'd6856, 16'd56207, 16'd45319, 16'd30306, 16'd23492, 16'd7673, 16'd3420, 16'd65081, 16'd48581, 16'd10826, 16'd7263, 16'd1973, 16'd62307, 16'd43378, 16'd23251, 16'd53126, 16'd42105, 16'd25558, 16'd5634, 16'd31659, 16'd7502, 16'd212, 16'd30336, 16'd45565, 16'd4086});
	test_expansion(128'ha355c8ad0594c3c8edd8d4b262afbcb0, {16'd63314, 16'd19033, 16'd19699, 16'd34797, 16'd15872, 16'd53221, 16'd31112, 16'd16933, 16'd10222, 16'd42665, 16'd51213, 16'd12266, 16'd4141, 16'd39153, 16'd50189, 16'd55416, 16'd12501, 16'd13881, 16'd46886, 16'd14816, 16'd21829, 16'd61354, 16'd14608, 16'd63063, 16'd53590, 16'd32740});
	test_expansion(128'h7293bcd066b8af8383bd8295c50f6090, {16'd7719, 16'd62540, 16'd6785, 16'd59519, 16'd45080, 16'd39789, 16'd44932, 16'd24711, 16'd49413, 16'd58218, 16'd60059, 16'd44277, 16'd9380, 16'd30587, 16'd26062, 16'd11097, 16'd16277, 16'd4059, 16'd33197, 16'd11339, 16'd33388, 16'd15034, 16'd19790, 16'd55389, 16'd12315, 16'd13602});
	test_expansion(128'h1678d34656f50b01e69c17d2ee1ece06, {16'd40187, 16'd11740, 16'd16844, 16'd33562, 16'd53628, 16'd29150, 16'd61247, 16'd34072, 16'd35019, 16'd3477, 16'd934, 16'd50100, 16'd39703, 16'd50636, 16'd36532, 16'd10552, 16'd5492, 16'd44240, 16'd43341, 16'd33361, 16'd23575, 16'd59357, 16'd19591, 16'd49676, 16'd17043, 16'd46665});
	test_expansion(128'hae602636bf05cc0a4fcd39fc1e3e9716, {16'd46623, 16'd65059, 16'd62026, 16'd23288, 16'd62596, 16'd1273, 16'd25113, 16'd53454, 16'd23596, 16'd24672, 16'd14124, 16'd57144, 16'd62473, 16'd727, 16'd24345, 16'd49089, 16'd31219, 16'd15226, 16'd8674, 16'd30082, 16'd19367, 16'd7965, 16'd13840, 16'd13435, 16'd23414, 16'd14119});
	test_expansion(128'hc2fb05f71369f1b122dcda46e72bbcae, {16'd56807, 16'd2857, 16'd51110, 16'd25165, 16'd4615, 16'd43205, 16'd15464, 16'd43197, 16'd54150, 16'd58622, 16'd2705, 16'd36592, 16'd48240, 16'd47166, 16'd29566, 16'd60416, 16'd11676, 16'd44005, 16'd5208, 16'd60424, 16'd58439, 16'd25888, 16'd40117, 16'd31251, 16'd37115, 16'd37046});
	test_expansion(128'h4b9729a41e5fb2d0941c7c55f87cac0c, {16'd26181, 16'd64732, 16'd2920, 16'd3692, 16'd35002, 16'd39146, 16'd30597, 16'd53263, 16'd43720, 16'd37239, 16'd3534, 16'd25382, 16'd58381, 16'd40609, 16'd38185, 16'd8332, 16'd13580, 16'd36790, 16'd59316, 16'd50192, 16'd16983, 16'd37878, 16'd6791, 16'd39682, 16'd43464, 16'd60437});
	test_expansion(128'hcfe86ca08e7c408afbee7414744a3e73, {16'd29812, 16'd35484, 16'd8266, 16'd22058, 16'd52834, 16'd30348, 16'd21545, 16'd18632, 16'd54830, 16'd37789, 16'd63316, 16'd7715, 16'd29265, 16'd19450, 16'd18215, 16'd53316, 16'd2931, 16'd5114, 16'd53942, 16'd17883, 16'd59827, 16'd1146, 16'd24839, 16'd31634, 16'd14881, 16'd17482});
	test_expansion(128'h7780bf1e4bdb113857e39ba90001f246, {16'd13594, 16'd6907, 16'd35961, 16'd53364, 16'd12765, 16'd34973, 16'd48387, 16'd27849, 16'd18851, 16'd22498, 16'd38280, 16'd62219, 16'd5364, 16'd28335, 16'd11706, 16'd28893, 16'd18006, 16'd62241, 16'd19728, 16'd1771, 16'd18165, 16'd20178, 16'd38634, 16'd11486, 16'd10864, 16'd47340});
	test_expansion(128'hb0a40fa6579c6360305f98ccc4befaa2, {16'd65122, 16'd16895, 16'd58663, 16'd2034, 16'd45616, 16'd60573, 16'd36335, 16'd55230, 16'd30247, 16'd16643, 16'd63716, 16'd21038, 16'd34041, 16'd41047, 16'd59634, 16'd14836, 16'd23320, 16'd24117, 16'd24748, 16'd4222, 16'd6788, 16'd1193, 16'd36321, 16'd35610, 16'd65200, 16'd50972});
	test_expansion(128'h164a2059d94139563ea6503401ba920f, {16'd4707, 16'd16430, 16'd51324, 16'd45682, 16'd5645, 16'd32203, 16'd49378, 16'd39972, 16'd13362, 16'd6105, 16'd62531, 16'd5492, 16'd51294, 16'd24315, 16'd31706, 16'd53956, 16'd28059, 16'd30540, 16'd32794, 16'd13340, 16'd26609, 16'd17954, 16'd49084, 16'd1112, 16'd27540, 16'd51857});
	test_expansion(128'hef00ee37993ba20827816d4aa717ef39, {16'd52488, 16'd52890, 16'd9476, 16'd20914, 16'd18415, 16'd2061, 16'd10442, 16'd21129, 16'd27335, 16'd15323, 16'd18258, 16'd9385, 16'd24319, 16'd18032, 16'd52172, 16'd12342, 16'd40235, 16'd21453, 16'd2470, 16'd6765, 16'd1440, 16'd60126, 16'd10407, 16'd31097, 16'd47466, 16'd8470});
	test_expansion(128'h59e9d323ca6da08ebf33e0e4fd9f7dd9, {16'd29933, 16'd40021, 16'd47659, 16'd39250, 16'd2358, 16'd6199, 16'd36154, 16'd29490, 16'd52733, 16'd5258, 16'd5206, 16'd7153, 16'd54607, 16'd37149, 16'd33639, 16'd24227, 16'd33966, 16'd62415, 16'd20745, 16'd23057, 16'd53796, 16'd8730, 16'd59735, 16'd59468, 16'd20831, 16'd49852});
	test_expansion(128'h9205f97bfbe9c046dda7c9ad52fefe18, {16'd50257, 16'd621, 16'd24936, 16'd48398, 16'd54682, 16'd51065, 16'd13557, 16'd26530, 16'd10, 16'd27970, 16'd14054, 16'd44816, 16'd44393, 16'd43716, 16'd29316, 16'd57279, 16'd40656, 16'd25559, 16'd35237, 16'd52872, 16'd56915, 16'd35235, 16'd32903, 16'd47357, 16'd22225, 16'd22670});
	test_expansion(128'h17af1399d38cf7491bf72f48dcff199a, {16'd60195, 16'd34479, 16'd1817, 16'd53057, 16'd52701, 16'd43177, 16'd17923, 16'd43539, 16'd30803, 16'd11540, 16'd63866, 16'd46462, 16'd38543, 16'd56486, 16'd54293, 16'd54551, 16'd57294, 16'd23070, 16'd46725, 16'd34684, 16'd17386, 16'd60962, 16'd64492, 16'd48003, 16'd43401, 16'd12200});
	test_expansion(128'h85bf8b65f2f4802a58fa7dcd2438e352, {16'd25879, 16'd57078, 16'd30576, 16'd39157, 16'd23994, 16'd6264, 16'd5862, 16'd27705, 16'd3273, 16'd28071, 16'd22235, 16'd34733, 16'd22391, 16'd47610, 16'd60740, 16'd10737, 16'd1866, 16'd6716, 16'd27922, 16'd36104, 16'd21951, 16'd6451, 16'd25095, 16'd5357, 16'd62529, 16'd1637});
	test_expansion(128'ha7f8b1af3ffff45919c1bce135e7a9b6, {16'd40191, 16'd50762, 16'd35207, 16'd42995, 16'd17324, 16'd16757, 16'd11455, 16'd555, 16'd47436, 16'd50044, 16'd61423, 16'd57595, 16'd18736, 16'd56683, 16'd36205, 16'd21846, 16'd41669, 16'd17003, 16'd13095, 16'd337, 16'd8979, 16'd10004, 16'd3852, 16'd38223, 16'd10595, 16'd58183});
	test_expansion(128'h1a8a15e2a89f6198a0ad87c0aa5755ac, {16'd16692, 16'd58393, 16'd32886, 16'd1912, 16'd15427, 16'd53445, 16'd10876, 16'd12985, 16'd16356, 16'd7730, 16'd42935, 16'd56244, 16'd25199, 16'd7819, 16'd53231, 16'd29798, 16'd63414, 16'd59578, 16'd2816, 16'd51800, 16'd4925, 16'd33078, 16'd49190, 16'd27272, 16'd25288, 16'd30169});
	test_expansion(128'hb7dd02f7393ea947bc09606b175326ce, {16'd55448, 16'd49447, 16'd47999, 16'd5516, 16'd52505, 16'd58944, 16'd38818, 16'd27495, 16'd28129, 16'd9056, 16'd22030, 16'd45380, 16'd31299, 16'd5732, 16'd93, 16'd23653, 16'd60808, 16'd41734, 16'd47538, 16'd55421, 16'd48365, 16'd56348, 16'd10991, 16'd19263, 16'd13604, 16'd39361});
	test_expansion(128'h46f19656e8e66ba619de4de6873877bf, {16'd63325, 16'd15276, 16'd62050, 16'd48629, 16'd43126, 16'd23263, 16'd1017, 16'd61657, 16'd30206, 16'd45744, 16'd53256, 16'd3904, 16'd8403, 16'd50810, 16'd2232, 16'd18790, 16'd53391, 16'd18383, 16'd10872, 16'd4517, 16'd20909, 16'd8023, 16'd32726, 16'd3977, 16'd42442, 16'd7550});
	test_expansion(128'h0abde3eba9ce23b46eaccd6ce8b9a556, {16'd60436, 16'd60529, 16'd53752, 16'd10214, 16'd54395, 16'd53156, 16'd6308, 16'd31327, 16'd27687, 16'd65151, 16'd22959, 16'd60458, 16'd8384, 16'd25840, 16'd28374, 16'd60250, 16'd29248, 16'd57905, 16'd10175, 16'd14328, 16'd25389, 16'd56513, 16'd19715, 16'd64981, 16'd50589, 16'd3237});
	test_expansion(128'h84d085767bfc338b4592282b63b3d041, {16'd44737, 16'd18082, 16'd28962, 16'd40572, 16'd17271, 16'd2334, 16'd30792, 16'd28971, 16'd25789, 16'd1243, 16'd39173, 16'd1513, 16'd27101, 16'd9336, 16'd42726, 16'd37570, 16'd47826, 16'd29691, 16'd8310, 16'd15450, 16'd9751, 16'd49944, 16'd20231, 16'd17134, 16'd30562, 16'd57240});
	test_expansion(128'h57e039d4278d3cdc693552f007c1e0fe, {16'd44738, 16'd13275, 16'd57825, 16'd46952, 16'd64726, 16'd19764, 16'd39003, 16'd1670, 16'd18399, 16'd16614, 16'd19978, 16'd45044, 16'd45491, 16'd59355, 16'd36678, 16'd5535, 16'd45305, 16'd46090, 16'd47115, 16'd2018, 16'd45934, 16'd11973, 16'd35838, 16'd10218, 16'd24185, 16'd14764});
	test_expansion(128'hf40a5568b3f89954ef203c11a85055e3, {16'd59540, 16'd8496, 16'd54207, 16'd7671, 16'd36846, 16'd7205, 16'd25050, 16'd29633, 16'd42392, 16'd6102, 16'd34292, 16'd53882, 16'd12286, 16'd4733, 16'd7738, 16'd19226, 16'd27238, 16'd14671, 16'd45852, 16'd45359, 16'd12364, 16'd37067, 16'd50704, 16'd32778, 16'd20192, 16'd24161});
	test_expansion(128'h7f923c40a9a61e961a832967f127b6fd, {16'd50690, 16'd43368, 16'd47512, 16'd3276, 16'd42416, 16'd57533, 16'd27150, 16'd7770, 16'd27139, 16'd22876, 16'd56194, 16'd5029, 16'd15060, 16'd7765, 16'd35004, 16'd36906, 16'd621, 16'd34457, 16'd39057, 16'd46967, 16'd8234, 16'd24946, 16'd4339, 16'd13290, 16'd643, 16'd52290});
	test_expansion(128'hfffd5a97ecd9c86aaf15c2f2b4464b14, {16'd22701, 16'd21392, 16'd36964, 16'd61538, 16'd44984, 16'd16166, 16'd46409, 16'd59916, 16'd59796, 16'd2414, 16'd61351, 16'd8491, 16'd64128, 16'd8426, 16'd18799, 16'd22095, 16'd36465, 16'd54598, 16'd50224, 16'd12835, 16'd65103, 16'd44265, 16'd50833, 16'd39242, 16'd27241, 16'd59342});
	test_expansion(128'h9af78b1a599f23a45131ecb6668cd364, {16'd52417, 16'd57413, 16'd4969, 16'd43702, 16'd12293, 16'd18347, 16'd6150, 16'd28266, 16'd44319, 16'd7537, 16'd36152, 16'd62161, 16'd42201, 16'd31116, 16'd15730, 16'd44232, 16'd5309, 16'd46345, 16'd9758, 16'd11079, 16'd55577, 16'd53772, 16'd25379, 16'd53594, 16'd26437, 16'd23862});
	test_expansion(128'ha0143cec8eb8c8ca5e06a1cb8bd611c2, {16'd5970, 16'd30866, 16'd35766, 16'd58590, 16'd63304, 16'd32675, 16'd28479, 16'd65354, 16'd56609, 16'd16761, 16'd31375, 16'd20005, 16'd29746, 16'd46024, 16'd8655, 16'd55299, 16'd16069, 16'd29773, 16'd56883, 16'd59575, 16'd56671, 16'd51173, 16'd25190, 16'd4473, 16'd30620, 16'd35063});
	test_expansion(128'h9835d7acaf39d09b31e712955af2e35b, {16'd7379, 16'd35936, 16'd57169, 16'd2820, 16'd13399, 16'd53360, 16'd33845, 16'd21460, 16'd18539, 16'd32657, 16'd27255, 16'd42737, 16'd21834, 16'd44674, 16'd59374, 16'd42324, 16'd49122, 16'd12038, 16'd43150, 16'd61677, 16'd19713, 16'd60992, 16'd45400, 16'd8701, 16'd59149, 16'd51848});
	test_expansion(128'h155d49bebeaa77953b49815447fc7e01, {16'd12678, 16'd2695, 16'd37651, 16'd58920, 16'd14596, 16'd19377, 16'd41970, 16'd58668, 16'd17806, 16'd14772, 16'd57796, 16'd59485, 16'd59224, 16'd197, 16'd42759, 16'd31974, 16'd58497, 16'd12493, 16'd128, 16'd15680, 16'd26940, 16'd45706, 16'd47034, 16'd37981, 16'd2071, 16'd33830});
	test_expansion(128'hb18dd44d84fcdbf9af4a4f0cd7c9f0fc, {16'd39624, 16'd48080, 16'd29467, 16'd8620, 16'd14606, 16'd25287, 16'd51693, 16'd13414, 16'd56923, 16'd3357, 16'd36621, 16'd41863, 16'd33899, 16'd8732, 16'd38832, 16'd1506, 16'd56195, 16'd40154, 16'd34694, 16'd12589, 16'd18049, 16'd17997, 16'd64884, 16'd44973, 16'd48266, 16'd9002});
	test_expansion(128'h0e73ebde53bbaf72f11312541f57f559, {16'd10495, 16'd45034, 16'd7321, 16'd3426, 16'd48773, 16'd23430, 16'd52721, 16'd15274, 16'd35101, 16'd32076, 16'd1368, 16'd23271, 16'd30206, 16'd30980, 16'd10477, 16'd32556, 16'd24123, 16'd18988, 16'd13666, 16'd9185, 16'd54088, 16'd11382, 16'd18591, 16'd9185, 16'd12483, 16'd59468});
	test_expansion(128'h2eec1e0968327a1c006b4b603492d717, {16'd15923, 16'd47225, 16'd41692, 16'd3105, 16'd34406, 16'd29719, 16'd41539, 16'd5598, 16'd42756, 16'd45997, 16'd8802, 16'd53522, 16'd63058, 16'd51082, 16'd59502, 16'd40774, 16'd10611, 16'd9311, 16'd64132, 16'd62121, 16'd32318, 16'd62060, 16'd27071, 16'd15166, 16'd48421, 16'd29565});
	test_expansion(128'hfb33773096e88d157908d56425da7515, {16'd56514, 16'd1612, 16'd40388, 16'd29056, 16'd45797, 16'd32221, 16'd22766, 16'd48872, 16'd54909, 16'd25158, 16'd21881, 16'd4490, 16'd24744, 16'd38831, 16'd60892, 16'd15261, 16'd53398, 16'd6614, 16'd47316, 16'd22798, 16'd9558, 16'd60396, 16'd36451, 16'd35425, 16'd35446, 16'd30696});
	test_expansion(128'h0fa1002718e5e019661c331a3fda357f, {16'd64665, 16'd41294, 16'd37493, 16'd39038, 16'd57763, 16'd30667, 16'd40445, 16'd41842, 16'd3254, 16'd52039, 16'd33916, 16'd12529, 16'd28531, 16'd16199, 16'd18934, 16'd64486, 16'd51947, 16'd25321, 16'd14283, 16'd32658, 16'd25713, 16'd59914, 16'd34721, 16'd49623, 16'd35098, 16'd12515});
	test_expansion(128'h5a16331b870d15f9a474db2a39dd0b85, {16'd46196, 16'd62023, 16'd41070, 16'd58666, 16'd31755, 16'd1417, 16'd9169, 16'd1090, 16'd5752, 16'd25643, 16'd29541, 16'd49988, 16'd64871, 16'd36476, 16'd16476, 16'd51791, 16'd10723, 16'd64333, 16'd61910, 16'd43328, 16'd738, 16'd41610, 16'd40934, 16'd19393, 16'd37260, 16'd54204});
	test_expansion(128'h1ca5b15f8b5fb9a3c767ecbe47b41302, {16'd64154, 16'd8625, 16'd62812, 16'd55619, 16'd59251, 16'd15769, 16'd150, 16'd36467, 16'd12422, 16'd42790, 16'd15821, 16'd28948, 16'd45187, 16'd55352, 16'd53474, 16'd39297, 16'd22611, 16'd64851, 16'd39814, 16'd22885, 16'd1040, 16'd50142, 16'd58618, 16'd285, 16'd49334, 16'd49114});
	test_expansion(128'h415d61407b94e81c653c09535d49bc37, {16'd42077, 16'd27648, 16'd1210, 16'd2549, 16'd55650, 16'd50582, 16'd26557, 16'd41186, 16'd23187, 16'd44307, 16'd53289, 16'd50857, 16'd8393, 16'd56894, 16'd43732, 16'd34689, 16'd48046, 16'd34039, 16'd49513, 16'd33485, 16'd38455, 16'd17450, 16'd50249, 16'd52545, 16'd49061, 16'd33316});
	test_expansion(128'hdf24b6750c519e08733c8c873eaa3ff4, {16'd27310, 16'd29652, 16'd55233, 16'd36125, 16'd3829, 16'd54348, 16'd9708, 16'd5672, 16'd3934, 16'd11771, 16'd7821, 16'd49830, 16'd21187, 16'd31736, 16'd34353, 16'd64040, 16'd28199, 16'd12067, 16'd36114, 16'd12758, 16'd33807, 16'd56622, 16'd50742, 16'd37059, 16'd35819, 16'd62365});
	test_expansion(128'h2f58bc6458f3e97bef7abd4ba9e4c7af, {16'd49171, 16'd62129, 16'd36994, 16'd2105, 16'd11335, 16'd24170, 16'd28092, 16'd128, 16'd267, 16'd13229, 16'd17946, 16'd41230, 16'd47609, 16'd36726, 16'd20373, 16'd27746, 16'd27047, 16'd40814, 16'd13614, 16'd3888, 16'd11607, 16'd33793, 16'd28300, 16'd2541, 16'd46047, 16'd18955});
	test_expansion(128'h004eff869b3ed343643eb1b50e8e8148, {16'd4413, 16'd41730, 16'd60850, 16'd60721, 16'd16074, 16'd32029, 16'd19505, 16'd21599, 16'd42609, 16'd40677, 16'd63730, 16'd43725, 16'd2311, 16'd9451, 16'd31734, 16'd43588, 16'd12247, 16'd59982, 16'd32622, 16'd33871, 16'd64510, 16'd49296, 16'd17994, 16'd11102, 16'd4952, 16'd48241});
	test_expansion(128'habb70fa8856baac799492cbb1ea782e7, {16'd25407, 16'd58202, 16'd3898, 16'd38646, 16'd4296, 16'd59145, 16'd53820, 16'd16028, 16'd51425, 16'd24814, 16'd61665, 16'd60938, 16'd3298, 16'd19527, 16'd1543, 16'd14644, 16'd20836, 16'd54531, 16'd14116, 16'd45905, 16'd46424, 16'd48682, 16'd5587, 16'd57780, 16'd42259, 16'd1170});
	test_expansion(128'h047d2a6fc834d631292de02adc07cf7e, {16'd7844, 16'd21721, 16'd1865, 16'd59656, 16'd37303, 16'd18265, 16'd54607, 16'd40805, 16'd12823, 16'd26332, 16'd46329, 16'd27914, 16'd5066, 16'd376, 16'd28844, 16'd5543, 16'd47345, 16'd54527, 16'd63740, 16'd17534, 16'd38027, 16'd60263, 16'd58577, 16'd27041, 16'd44361, 16'd48649});
	test_expansion(128'h3d92b29a3cee7420d28eaf7dd6491031, {16'd50058, 16'd14532, 16'd54474, 16'd31668, 16'd5233, 16'd60132, 16'd10134, 16'd51339, 16'd9839, 16'd17564, 16'd34502, 16'd59757, 16'd39122, 16'd43594, 16'd51843, 16'd26563, 16'd48259, 16'd4910, 16'd31679, 16'd20878, 16'd47763, 16'd62792, 16'd9720, 16'd3537, 16'd40467, 16'd15822});
	test_expansion(128'hebd361f57dc897d26e895b7c9e530b3b, {16'd47792, 16'd34213, 16'd56637, 16'd13768, 16'd17183, 16'd15203, 16'd50211, 16'd11862, 16'd17285, 16'd62221, 16'd61226, 16'd27430, 16'd13184, 16'd8840, 16'd42714, 16'd20343, 16'd4436, 16'd1796, 16'd13407, 16'd5507, 16'd44755, 16'd64056, 16'd50831, 16'd55801, 16'd48704, 16'd22673});
	test_expansion(128'h0cb05f758e0c1780bf4b8068450707da, {16'd18110, 16'd14513, 16'd17161, 16'd17198, 16'd54541, 16'd10188, 16'd36944, 16'd25957, 16'd52465, 16'd36222, 16'd7928, 16'd44326, 16'd28478, 16'd23412, 16'd9251, 16'd24651, 16'd24796, 16'd46875, 16'd40540, 16'd33790, 16'd35905, 16'd1401, 16'd46220, 16'd9398, 16'd20336, 16'd17085});
	test_expansion(128'haed49be178d874b8d635f96e80ced9b8, {16'd47036, 16'd2111, 16'd43726, 16'd36522, 16'd43453, 16'd20245, 16'd50692, 16'd18666, 16'd60826, 16'd16889, 16'd5212, 16'd21420, 16'd8118, 16'd55287, 16'd8168, 16'd35553, 16'd30322, 16'd24801, 16'd27790, 16'd46407, 16'd56408, 16'd10094, 16'd10412, 16'd6233, 16'd43424, 16'd56925});
	test_expansion(128'h23b4b5dd8b541fc116d3be239746ca4b, {16'd47183, 16'd54905, 16'd13160, 16'd34580, 16'd2783, 16'd18469, 16'd5817, 16'd32331, 16'd17521, 16'd51536, 16'd61296, 16'd13871, 16'd56409, 16'd33683, 16'd31378, 16'd16557, 16'd54218, 16'd27459, 16'd34769, 16'd35307, 16'd16704, 16'd31760, 16'd9779, 16'd45653, 16'd9294, 16'd15532});
	test_expansion(128'h44f08bbaa87bebbb1bc33712aed864fa, {16'd39800, 16'd3585, 16'd52957, 16'd38373, 16'd27761, 16'd5335, 16'd23127, 16'd4666, 16'd3284, 16'd22614, 16'd33635, 16'd4704, 16'd28950, 16'd53877, 16'd32015, 16'd62873, 16'd14718, 16'd47102, 16'd27687, 16'd1419, 16'd36458, 16'd19615, 16'd22018, 16'd9487, 16'd63708, 16'd62525});
	test_expansion(128'h1a0ee3a7281a4242e27d300b6f2b1613, {16'd52362, 16'd16379, 16'd37134, 16'd39599, 16'd45985, 16'd22720, 16'd39165, 16'd42735, 16'd49505, 16'd57087, 16'd23352, 16'd53888, 16'd61931, 16'd35538, 16'd52951, 16'd59480, 16'd39767, 16'd34018, 16'd29535, 16'd6774, 16'd32811, 16'd23893, 16'd48203, 16'd59677, 16'd5316, 16'd54789});
	test_expansion(128'h149828b7dee23d06c1ab9e3fbab98eec, {16'd36306, 16'd50108, 16'd23592, 16'd41621, 16'd36989, 16'd46672, 16'd5518, 16'd60675, 16'd23454, 16'd57637, 16'd13757, 16'd45127, 16'd29326, 16'd35728, 16'd25867, 16'd2474, 16'd46578, 16'd32458, 16'd43076, 16'd6251, 16'd13616, 16'd49208, 16'd16105, 16'd22098, 16'd27032, 16'd14351});
	test_expansion(128'h8a93d27741a9ef3f069f549b4e029cc6, {16'd59584, 16'd25055, 16'd53895, 16'd64927, 16'd35109, 16'd26889, 16'd27052, 16'd63195, 16'd23049, 16'd49401, 16'd55951, 16'd57825, 16'd7971, 16'd42507, 16'd39949, 16'd42933, 16'd10278, 16'd2259, 16'd18049, 16'd56287, 16'd5154, 16'd22440, 16'd13859, 16'd35011, 16'd22091, 16'd8063});
	test_expansion(128'h18829121577ed378399f76b2db211a18, {16'd6405, 16'd40056, 16'd41387, 16'd55221, 16'd40437, 16'd57815, 16'd23554, 16'd5961, 16'd60370, 16'd57791, 16'd33631, 16'd37358, 16'd2182, 16'd17956, 16'd10974, 16'd31152, 16'd11453, 16'd43494, 16'd2680, 16'd57809, 16'd37615, 16'd25067, 16'd30792, 16'd63181, 16'd195, 16'd38010});
	test_expansion(128'h1d512bc91ff69af0852d804879755607, {16'd507, 16'd2324, 16'd2944, 16'd25208, 16'd5951, 16'd48957, 16'd61335, 16'd35532, 16'd11907, 16'd54720, 16'd54574, 16'd34824, 16'd50606, 16'd39252, 16'd26408, 16'd41647, 16'd58977, 16'd53134, 16'd17606, 16'd14109, 16'd745, 16'd21104, 16'd8416, 16'd22799, 16'd21074, 16'd21064});
	test_expansion(128'h1cce6ca417b61c1b4ce117ae710f988b, {16'd59728, 16'd58661, 16'd29597, 16'd59526, 16'd31032, 16'd6682, 16'd1504, 16'd11410, 16'd52329, 16'd50455, 16'd8017, 16'd65402, 16'd39609, 16'd52658, 16'd59465, 16'd48290, 16'd50469, 16'd34098, 16'd51637, 16'd465, 16'd21151, 16'd30178, 16'd30675, 16'd48279, 16'd11614, 16'd25275});
	test_expansion(128'h3b197d93d6b0e58b6ebedfaa832d9f86, {16'd58220, 16'd6996, 16'd14862, 16'd23539, 16'd42434, 16'd57790, 16'd16297, 16'd47271, 16'd14443, 16'd15485, 16'd18919, 16'd41965, 16'd39268, 16'd49320, 16'd3418, 16'd41424, 16'd10608, 16'd7730, 16'd49069, 16'd17618, 16'd4485, 16'd19396, 16'd22751, 16'd45629, 16'd23680, 16'd29839});
	test_expansion(128'h85af780d764a4a5b080f69008d9d46c5, {16'd33564, 16'd37558, 16'd32643, 16'd47618, 16'd38270, 16'd11741, 16'd55820, 16'd9837, 16'd24475, 16'd51218, 16'd26778, 16'd18567, 16'd10217, 16'd59068, 16'd33355, 16'd45792, 16'd28712, 16'd26146, 16'd35949, 16'd33619, 16'd10628, 16'd42152, 16'd26358, 16'd332, 16'd39666, 16'd13657});
	test_expansion(128'h323e733d8a8e9ed99e7ea6607befa831, {16'd10655, 16'd49681, 16'd46012, 16'd46409, 16'd38205, 16'd50483, 16'd14781, 16'd52698, 16'd61915, 16'd58041, 16'd22242, 16'd64443, 16'd64584, 16'd44997, 16'd62461, 16'd21995, 16'd979, 16'd55163, 16'd57281, 16'd2452, 16'd4430, 16'd9755, 16'd28982, 16'd32345, 16'd27757, 16'd429});
	test_expansion(128'h725986eddc95044fd412b7339290205b, {16'd47919, 16'd29750, 16'd3562, 16'd4383, 16'd50785, 16'd1375, 16'd26822, 16'd7691, 16'd2048, 16'd15397, 16'd55882, 16'd30231, 16'd57110, 16'd48306, 16'd48237, 16'd17015, 16'd5117, 16'd40537, 16'd54948, 16'd5744, 16'd4755, 16'd31415, 16'd59329, 16'd53937, 16'd32386, 16'd44284});
	test_expansion(128'h0133ab6dc665d945eb25e3a8ebc851de, {16'd4431, 16'd4451, 16'd42056, 16'd54235, 16'd55390, 16'd38602, 16'd25831, 16'd56891, 16'd43649, 16'd44002, 16'd65144, 16'd6084, 16'd52803, 16'd57300, 16'd47386, 16'd6605, 16'd42731, 16'd22323, 16'd35980, 16'd1864, 16'd19862, 16'd40627, 16'd28100, 16'd57943, 16'd61633, 16'd640});
	test_expansion(128'h1d64550e2b626d543a267645ea8f7918, {16'd11255, 16'd13272, 16'd1231, 16'd22180, 16'd58009, 16'd11799, 16'd58690, 16'd18248, 16'd21861, 16'd7874, 16'd5016, 16'd32439, 16'd2632, 16'd29812, 16'd64375, 16'd4446, 16'd43933, 16'd62205, 16'd16251, 16'd27144, 16'd63496, 16'd57691, 16'd39069, 16'd33968, 16'd65203, 16'd41298});
	test_expansion(128'h37c47596aa729f6de88310165af9432f, {16'd32457, 16'd9199, 16'd14325, 16'd56319, 16'd40803, 16'd9359, 16'd57047, 16'd42612, 16'd48245, 16'd41245, 16'd7165, 16'd18601, 16'd60949, 16'd20074, 16'd16000, 16'd9011, 16'd36035, 16'd22910, 16'd63533, 16'd12561, 16'd29747, 16'd63832, 16'd60563, 16'd28055, 16'd55206, 16'd49232});
	test_expansion(128'h59fef812fe356cec3e89233b82a77f5f, {16'd57150, 16'd65239, 16'd9175, 16'd28254, 16'd36808, 16'd35605, 16'd51252, 16'd23839, 16'd33178, 16'd46261, 16'd49666, 16'd59593, 16'd14200, 16'd62282, 16'd62862, 16'd52235, 16'd36474, 16'd7311, 16'd8699, 16'd10334, 16'd1698, 16'd47319, 16'd7459, 16'd61312, 16'd41942, 16'd29200});
	test_expansion(128'h3660111d907e3267ca0495d1d7049614, {16'd25561, 16'd56596, 16'd6108, 16'd48226, 16'd10082, 16'd10984, 16'd26177, 16'd2520, 16'd44283, 16'd42747, 16'd26044, 16'd56494, 16'd28695, 16'd46192, 16'd37349, 16'd13753, 16'd49446, 16'd26343, 16'd49978, 16'd30397, 16'd23272, 16'd30699, 16'd39460, 16'd16199, 16'd32832, 16'd3616});
	test_expansion(128'h44be5ce8f14bcbec7b52ea7de9815f72, {16'd11592, 16'd9451, 16'd24148, 16'd54535, 16'd2501, 16'd63581, 16'd57134, 16'd9948, 16'd23214, 16'd64855, 16'd39702, 16'd5018, 16'd45708, 16'd14913, 16'd36482, 16'd51414, 16'd11871, 16'd31801, 16'd39608, 16'd18855, 16'd31795, 16'd20992, 16'd29828, 16'd30473, 16'd6997, 16'd10690});
	test_expansion(128'h525cc212e4d5bdaf2dee070ba49754e1, {16'd65282, 16'd22760, 16'd45575, 16'd25553, 16'd26073, 16'd53484, 16'd17169, 16'd26958, 16'd11908, 16'd51583, 16'd52781, 16'd49806, 16'd48375, 16'd46163, 16'd53474, 16'd36880, 16'd24490, 16'd19535, 16'd10634, 16'd9827, 16'd20732, 16'd50873, 16'd45296, 16'd51592, 16'd43989, 16'd46768});
	test_expansion(128'h5bc67eed2b00c28754d0f3e199499638, {16'd19292, 16'd28085, 16'd49558, 16'd65414, 16'd63927, 16'd33342, 16'd53574, 16'd40986, 16'd2762, 16'd56520, 16'd15975, 16'd60186, 16'd28203, 16'd20805, 16'd43036, 16'd5054, 16'd5256, 16'd44873, 16'd35298, 16'd41894, 16'd36591, 16'd38618, 16'd61840, 16'd9900, 16'd23342, 16'd55849});
	test_expansion(128'h9c0fd2148d3103a7cc823b8ba5850f3d, {16'd11345, 16'd54435, 16'd1096, 16'd7019, 16'd10948, 16'd22741, 16'd3483, 16'd48909, 16'd56999, 16'd38635, 16'd41959, 16'd64435, 16'd61103, 16'd36010, 16'd40666, 16'd36017, 16'd5901, 16'd47842, 16'd51606, 16'd55680, 16'd56815, 16'd9951, 16'd45392, 16'd2642, 16'd21422, 16'd19492});
	test_expansion(128'hf25fb356cb4c2a710882e63d981798ac, {16'd20900, 16'd31391, 16'd51441, 16'd23, 16'd47300, 16'd28778, 16'd6416, 16'd140, 16'd26971, 16'd27234, 16'd1004, 16'd57485, 16'd50513, 16'd5399, 16'd61756, 16'd34093, 16'd28729, 16'd63021, 16'd43062, 16'd8628, 16'd43647, 16'd35569, 16'd23031, 16'd44701, 16'd5261, 16'd12649});
	test_expansion(128'h9ebe2dade24be9769b5fa7c275df7a78, {16'd29897, 16'd56932, 16'd42577, 16'd41075, 16'd50621, 16'd25243, 16'd34942, 16'd16836, 16'd6235, 16'd28965, 16'd42875, 16'd42546, 16'd54267, 16'd15286, 16'd64964, 16'd61538, 16'd27381, 16'd3791, 16'd55658, 16'd52686, 16'd16346, 16'd27128, 16'd13108, 16'd5069, 16'd10652, 16'd15436});
	test_expansion(128'hfe18351734ad38909e220e23db3f80ba, {16'd3182, 16'd51031, 16'd6603, 16'd22920, 16'd2190, 16'd56196, 16'd26766, 16'd42698, 16'd37041, 16'd26640, 16'd14936, 16'd37015, 16'd22607, 16'd60233, 16'd664, 16'd34230, 16'd46083, 16'd34845, 16'd63325, 16'd19886, 16'd666, 16'd1722, 16'd62191, 16'd23495, 16'd46372, 16'd27453});
	test_expansion(128'hf9b532efa65a627cb47c0de14df019e4, {16'd60610, 16'd19033, 16'd7333, 16'd3219, 16'd24737, 16'd64193, 16'd42044, 16'd61498, 16'd33152, 16'd43413, 16'd60987, 16'd6380, 16'd48076, 16'd12441, 16'd56053, 16'd63957, 16'd37070, 16'd304, 16'd26372, 16'd30790, 16'd57267, 16'd22993, 16'd42392, 16'd56310, 16'd27868, 16'd60508});
	test_expansion(128'h001c3079287a41e7eeac6d3c0ab9c9f9, {16'd26370, 16'd9082, 16'd24244, 16'd53611, 16'd31408, 16'd55230, 16'd39473, 16'd24282, 16'd31138, 16'd1671, 16'd50781, 16'd9149, 16'd21901, 16'd3068, 16'd4967, 16'd11293, 16'd10338, 16'd12006, 16'd11209, 16'd32801, 16'd40727, 16'd36430, 16'd27453, 16'd49097, 16'd48244, 16'd12084});
	test_expansion(128'ha23b283e7e90eac084f4d005cec5ef17, {16'd59546, 16'd61689, 16'd37684, 16'd13055, 16'd14381, 16'd39724, 16'd18353, 16'd21010, 16'd35688, 16'd48855, 16'd1017, 16'd60594, 16'd49692, 16'd8576, 16'd47202, 16'd33294, 16'd62351, 16'd30117, 16'd18746, 16'd45568, 16'd53970, 16'd37855, 16'd46925, 16'd25569, 16'd12120, 16'd43073});
	test_expansion(128'h0b0f728e25d6f156f9f3f908f32c547f, {16'd39383, 16'd33431, 16'd27023, 16'd45553, 16'd54308, 16'd39711, 16'd32661, 16'd26790, 16'd44245, 16'd64295, 16'd26082, 16'd32759, 16'd48758, 16'd1184, 16'd5258, 16'd52332, 16'd7580, 16'd17577, 16'd27373, 16'd42339, 16'd50455, 16'd55430, 16'd40137, 16'd19340, 16'd58489, 16'd24357});
	test_expansion(128'h1d52701fac4fd71d0a5619d39e1cefc0, {16'd22540, 16'd26358, 16'd51668, 16'd40769, 16'd38589, 16'd7365, 16'd1414, 16'd47213, 16'd9912, 16'd39833, 16'd49029, 16'd64131, 16'd20656, 16'd64331, 16'd58736, 16'd13958, 16'd47087, 16'd51235, 16'd6687, 16'd16632, 16'd44860, 16'd35503, 16'd15345, 16'd10352, 16'd54886, 16'd4391});
	test_expansion(128'h34661aa8f504d49ea5e858f43ac918be, {16'd21235, 16'd24738, 16'd54754, 16'd20525, 16'd36860, 16'd50703, 16'd56759, 16'd39126, 16'd41406, 16'd26058, 16'd50502, 16'd23427, 16'd22094, 16'd63237, 16'd25943, 16'd5847, 16'd7618, 16'd38842, 16'd18205, 16'd28990, 16'd38593, 16'd44294, 16'd31707, 16'd30606, 16'd33317, 16'd15895});
	test_expansion(128'h499c0470130439b1e49264693fda396c, {16'd9148, 16'd57079, 16'd56428, 16'd43481, 16'd42335, 16'd5221, 16'd29829, 16'd63391, 16'd43550, 16'd8017, 16'd14821, 16'd62263, 16'd5644, 16'd332, 16'd60418, 16'd63891, 16'd60890, 16'd7706, 16'd61913, 16'd34775, 16'd46134, 16'd35797, 16'd6814, 16'd9058, 16'd34930, 16'd32216});
	test_expansion(128'h3bdb73bf2e983f296c2fcde0459a3a61, {16'd29869, 16'd9891, 16'd31596, 16'd12641, 16'd2050, 16'd9018, 16'd42106, 16'd27308, 16'd60034, 16'd56414, 16'd19407, 16'd1281, 16'd57149, 16'd13859, 16'd4905, 16'd41640, 16'd44375, 16'd41692, 16'd13105, 16'd28520, 16'd31621, 16'd25416, 16'd19681, 16'd34847, 16'd29753, 16'd50619});
	test_expansion(128'h5499f941c7395cc160ac20691501f369, {16'd27075, 16'd32527, 16'd59764, 16'd2206, 16'd7064, 16'd51096, 16'd13043, 16'd7137, 16'd6727, 16'd24158, 16'd35485, 16'd48104, 16'd53789, 16'd5220, 16'd23867, 16'd12570, 16'd11690, 16'd16549, 16'd41527, 16'd23902, 16'd13568, 16'd34794, 16'd42361, 16'd64967, 16'd14966, 16'd45262});
	test_expansion(128'h48b3d9e0f3890fad84f30ee455aaf6c8, {16'd56796, 16'd1960, 16'd57552, 16'd62705, 16'd27945, 16'd24258, 16'd8499, 16'd59012, 16'd56635, 16'd39287, 16'd23630, 16'd27885, 16'd28029, 16'd8415, 16'd62306, 16'd53049, 16'd57508, 16'd2658, 16'd40054, 16'd19615, 16'd45533, 16'd46372, 16'd10503, 16'd11361, 16'd39737, 16'd4178});
	test_expansion(128'h354a38afe7faa5f5644721b180c9a7bd, {16'd32978, 16'd56393, 16'd63574, 16'd35641, 16'd1725, 16'd15604, 16'd51894, 16'd63781, 16'd27777, 16'd13744, 16'd23832, 16'd15149, 16'd31026, 16'd30143, 16'd64551, 16'd13211, 16'd51622, 16'd26013, 16'd38876, 16'd48698, 16'd62631, 16'd10071, 16'd6925, 16'd27845, 16'd4900, 16'd343});
	test_expansion(128'h10a3517b97b2247f0b59438edb0c924c, {16'd14901, 16'd11051, 16'd55276, 16'd47844, 16'd31471, 16'd32444, 16'd58128, 16'd12585, 16'd45770, 16'd27566, 16'd9319, 16'd30451, 16'd35618, 16'd29893, 16'd51069, 16'd14063, 16'd50193, 16'd46903, 16'd30002, 16'd44899, 16'd2932, 16'd23418, 16'd60767, 16'd51029, 16'd5831, 16'd15216});
	test_expansion(128'he5740e0702cd3ca881f1dccdb33d01ec, {16'd41292, 16'd21193, 16'd1381, 16'd10049, 16'd30353, 16'd56912, 16'd36533, 16'd42430, 16'd39512, 16'd61877, 16'd7605, 16'd23739, 16'd34847, 16'd63156, 16'd32347, 16'd13710, 16'd41158, 16'd6395, 16'd64748, 16'd14466, 16'd27014, 16'd7267, 16'd63144, 16'd32870, 16'd62950, 16'd40746});
	test_expansion(128'hff06ff030483641423e15bee8b0e3954, {16'd10524, 16'd25344, 16'd48159, 16'd54343, 16'd5291, 16'd32874, 16'd30377, 16'd49180, 16'd16043, 16'd35737, 16'd27792, 16'd41567, 16'd64540, 16'd59892, 16'd15937, 16'd15980, 16'd9785, 16'd61050, 16'd22845, 16'd57518, 16'd39385, 16'd40925, 16'd19397, 16'd38345, 16'd38296, 16'd38935});
	test_expansion(128'h951af15ce671b446777b6dbc73ca61bd, {16'd43372, 16'd50607, 16'd3115, 16'd59248, 16'd31896, 16'd57530, 16'd50198, 16'd284, 16'd11405, 16'd2859, 16'd28581, 16'd19202, 16'd51484, 16'd33507, 16'd50296, 16'd18361, 16'd57122, 16'd31718, 16'd61310, 16'd16791, 16'd10139, 16'd20943, 16'd21301, 16'd62752, 16'd31292, 16'd41901});
	test_expansion(128'hd529651d37f59ecc9999c46df66d3167, {16'd34663, 16'd46212, 16'd23172, 16'd1651, 16'd53667, 16'd64647, 16'd41927, 16'd47453, 16'd15183, 16'd59669, 16'd58602, 16'd59236, 16'd57136, 16'd17209, 16'd50822, 16'd32182, 16'd20280, 16'd48369, 16'd8749, 16'd33539, 16'd58832, 16'd30074, 16'd38886, 16'd28687, 16'd36185, 16'd22094});
	test_expansion(128'hcfaddac5d8c1bef8a1994c762abf197f, {16'd2409, 16'd14569, 16'd39877, 16'd55129, 16'd59059, 16'd7040, 16'd59431, 16'd53085, 16'd52839, 16'd32743, 16'd28412, 16'd24461, 16'd48030, 16'd11622, 16'd37777, 16'd44891, 16'd34733, 16'd46363, 16'd53305, 16'd22040, 16'd40981, 16'd13624, 16'd33285, 16'd34402, 16'd45910, 16'd53139});
	test_expansion(128'h4bb2f2d5b3a89ac95ea173fe851878ff, {16'd36142, 16'd46368, 16'd30441, 16'd31068, 16'd6839, 16'd63099, 16'd25099, 16'd3115, 16'd25581, 16'd43449, 16'd61268, 16'd50703, 16'd22535, 16'd23324, 16'd44281, 16'd61001, 16'd23116, 16'd20098, 16'd54807, 16'd23213, 16'd20706, 16'd49607, 16'd61569, 16'd14847, 16'd24054, 16'd18293});
	test_expansion(128'ha0a60d0db4806c0036a477ae5e649916, {16'd8651, 16'd9568, 16'd25109, 16'd28744, 16'd47173, 16'd35913, 16'd6729, 16'd52775, 16'd8966, 16'd458, 16'd35270, 16'd32079, 16'd36190, 16'd2389, 16'd2631, 16'd32479, 16'd40976, 16'd62779, 16'd52850, 16'd65393, 16'd64008, 16'd12822, 16'd37138, 16'd54650, 16'd57992, 16'd198});
	test_expansion(128'h21543a6cd4f79dead36770432e063389, {16'd43442, 16'd40560, 16'd9571, 16'd33533, 16'd3540, 16'd62602, 16'd61872, 16'd34544, 16'd41835, 16'd58550, 16'd23175, 16'd15238, 16'd37727, 16'd47177, 16'd17168, 16'd2486, 16'd47923, 16'd38327, 16'd42024, 16'd44672, 16'd58483, 16'd3791, 16'd57758, 16'd25288, 16'd1870, 16'd57931});
	test_expansion(128'h73c24748c3e6c5ea68e44daf33e7c274, {16'd29552, 16'd38679, 16'd52761, 16'd50111, 16'd18320, 16'd7277, 16'd47712, 16'd57209, 16'd4135, 16'd11045, 16'd43484, 16'd15213, 16'd43425, 16'd2733, 16'd24164, 16'd52941, 16'd29691, 16'd37248, 16'd64420, 16'd59314, 16'd35871, 16'd50559, 16'd61876, 16'd53416, 16'd18551, 16'd36535});
	test_expansion(128'h1c21fe3eabee8c5923c9fbb31a048177, {16'd54353, 16'd13547, 16'd6872, 16'd49967, 16'd58099, 16'd46123, 16'd56326, 16'd33407, 16'd2832, 16'd54192, 16'd49403, 16'd57066, 16'd28713, 16'd60292, 16'd24599, 16'd31626, 16'd29529, 16'd7233, 16'd48730, 16'd8147, 16'd50066, 16'd4505, 16'd63428, 16'd33725, 16'd27105, 16'd45018});
	test_expansion(128'hcd3cfb219b859220ef3a33760f033718, {16'd1443, 16'd59035, 16'd46532, 16'd19081, 16'd60393, 16'd45130, 16'd23891, 16'd7691, 16'd40410, 16'd21898, 16'd41752, 16'd443, 16'd18473, 16'd35567, 16'd24520, 16'd53315, 16'd62041, 16'd46005, 16'd51114, 16'd16247, 16'd53324, 16'd64255, 16'd6485, 16'd45808, 16'd17467, 16'd14272});
	test_expansion(128'h6cf1a6e05c087710db261c1ee88590af, {16'd43363, 16'd26369, 16'd35512, 16'd53940, 16'd18426, 16'd39569, 16'd22879, 16'd12704, 16'd19598, 16'd1170, 16'd2291, 16'd22716, 16'd47792, 16'd58059, 16'd25932, 16'd16210, 16'd39075, 16'd12872, 16'd28494, 16'd5154, 16'd8212, 16'd23856, 16'd4659, 16'd44717, 16'd25955, 16'd18267});
	test_expansion(128'h74aa3badd8f2502ed134790b52afc9de, {16'd18419, 16'd18418, 16'd61114, 16'd53299, 16'd43538, 16'd35959, 16'd38395, 16'd40353, 16'd1037, 16'd45444, 16'd58209, 16'd2205, 16'd6737, 16'd27690, 16'd24086, 16'd21798, 16'd34586, 16'd62960, 16'd62677, 16'd40834, 16'd14789, 16'd57494, 16'd27193, 16'd5419, 16'd42717, 16'd20038});
	test_expansion(128'h1c461b94169fb41a6107c4bebeda3a69, {16'd32971, 16'd34919, 16'd15916, 16'd27181, 16'd25093, 16'd21236, 16'd39376, 16'd6336, 16'd54212, 16'd11785, 16'd53308, 16'd41891, 16'd52619, 16'd40515, 16'd6208, 16'd61768, 16'd20222, 16'd49855, 16'd42445, 16'd15113, 16'd2007, 16'd64516, 16'd16600, 16'd55773, 16'd55923, 16'd39230});
	test_expansion(128'hdadd87910359574a5af27433bee22497, {16'd29058, 16'd59512, 16'd38994, 16'd49310, 16'd10131, 16'd167, 16'd48879, 16'd13916, 16'd38155, 16'd43418, 16'd24876, 16'd44665, 16'd43922, 16'd13194, 16'd24742, 16'd36582, 16'd43187, 16'd55916, 16'd61161, 16'd51677, 16'd53640, 16'd17449, 16'd21101, 16'd18735, 16'd34481, 16'd18915});
	test_expansion(128'he74420209cafe555fcbdae437b54491d, {16'd4990, 16'd1469, 16'd24092, 16'd62250, 16'd48371, 16'd34316, 16'd33106, 16'd2456, 16'd41861, 16'd48287, 16'd56641, 16'd40926, 16'd24080, 16'd7705, 16'd44065, 16'd5790, 16'd24717, 16'd8707, 16'd14448, 16'd35945, 16'd52058, 16'd48980, 16'd27901, 16'd7241, 16'd46521, 16'd46853});
	test_expansion(128'he5c1a83ef6c77e2543cfd45ed6eb7614, {16'd59703, 16'd3140, 16'd27160, 16'd9946, 16'd21025, 16'd35430, 16'd16069, 16'd59675, 16'd61048, 16'd47714, 16'd56239, 16'd12238, 16'd877, 16'd26954, 16'd58877, 16'd45366, 16'd42263, 16'd37074, 16'd54106, 16'd21643, 16'd36990, 16'd881, 16'd32784, 16'd23077, 16'd38454, 16'd58290});
	test_expansion(128'h43ae15038affd697118da74546e7b6f0, {16'd27248, 16'd2626, 16'd9444, 16'd38733, 16'd25225, 16'd8046, 16'd9427, 16'd60572, 16'd48444, 16'd28933, 16'd14143, 16'd52716, 16'd20470, 16'd42023, 16'd44407, 16'd36333, 16'd41177, 16'd7057, 16'd24140, 16'd20012, 16'd25748, 16'd27048, 16'd23196, 16'd64752, 16'd9803, 16'd27082});
	test_expansion(128'h041d3751b00c27bfad79e5be40147490, {16'd14737, 16'd38194, 16'd9506, 16'd59641, 16'd10622, 16'd53313, 16'd43876, 16'd56593, 16'd35786, 16'd7851, 16'd55305, 16'd59810, 16'd43853, 16'd31091, 16'd6694, 16'd11736, 16'd35127, 16'd36952, 16'd24160, 16'd29453, 16'd32414, 16'd14305, 16'd25412, 16'd20554, 16'd26207, 16'd53743});
	test_expansion(128'h963c1588c5f1dc4d6844510b5254bf7d, {16'd30617, 16'd52716, 16'd13807, 16'd38263, 16'd31318, 16'd49975, 16'd50859, 16'd28442, 16'd63168, 16'd49899, 16'd10901, 16'd28399, 16'd61762, 16'd28246, 16'd4314, 16'd35900, 16'd35531, 16'd28016, 16'd62761, 16'd12042, 16'd11796, 16'd17481, 16'd35655, 16'd37105, 16'd18988, 16'd6596});
	test_expansion(128'h25dc62d02ac06f646fc1cb0e9bd481e9, {16'd61597, 16'd59536, 16'd9325, 16'd16750, 16'd62045, 16'd21358, 16'd38394, 16'd13945, 16'd9735, 16'd8323, 16'd3122, 16'd20690, 16'd58453, 16'd43776, 16'd61132, 16'd64379, 16'd21419, 16'd46459, 16'd24366, 16'd45838, 16'd18936, 16'd12291, 16'd13364, 16'd49257, 16'd19732, 16'd23331});
	test_expansion(128'hc65dcad92a70a033fe54beb965055a3f, {16'd8136, 16'd1853, 16'd8222, 16'd32719, 16'd48288, 16'd8545, 16'd44338, 16'd63630, 16'd5540, 16'd62849, 16'd44909, 16'd9086, 16'd17623, 16'd29248, 16'd44405, 16'd51814, 16'd26654, 16'd38858, 16'd39498, 16'd44435, 16'd58976, 16'd43699, 16'd27743, 16'd45671, 16'd3599, 16'd42890});
	test_expansion(128'hfcbc90fc9f9d86366b388ae720efda86, {16'd42130, 16'd26230, 16'd45342, 16'd61372, 16'd44078, 16'd16011, 16'd34437, 16'd63226, 16'd6147, 16'd4818, 16'd19225, 16'd30729, 16'd48165, 16'd38641, 16'd25549, 16'd58470, 16'd60489, 16'd4120, 16'd43264, 16'd28516, 16'd31412, 16'd61401, 16'd33485, 16'd53567, 16'd3790, 16'd65424});
	test_expansion(128'hdb37dcc15bd52a0eba3b0b1a17764db8, {16'd2478, 16'd38611, 16'd28218, 16'd23811, 16'd24714, 16'd9347, 16'd44832, 16'd10689, 16'd47029, 16'd21167, 16'd17420, 16'd6597, 16'd52784, 16'd23500, 16'd57588, 16'd44134, 16'd60366, 16'd51802, 16'd34780, 16'd6670, 16'd8130, 16'd12879, 16'd48340, 16'd18468, 16'd52800, 16'd11941});
	test_expansion(128'h573ba02e6dfe4359560ddc188b97ebf6, {16'd5344, 16'd54650, 16'd36913, 16'd5415, 16'd58178, 16'd46247, 16'd5698, 16'd64858, 16'd20961, 16'd63054, 16'd9579, 16'd53800, 16'd38785, 16'd3760, 16'd14833, 16'd4128, 16'd18943, 16'd61992, 16'd25372, 16'd13273, 16'd19903, 16'd5487, 16'd610, 16'd8194, 16'd11102, 16'd26391});
	test_expansion(128'h76ebd6cc97f92714b622d44f974a7c9f, {16'd20374, 16'd13795, 16'd33908, 16'd1496, 16'd40241, 16'd17988, 16'd40559, 16'd23793, 16'd19531, 16'd32704, 16'd37529, 16'd61203, 16'd12339, 16'd38239, 16'd55874, 16'd47993, 16'd53111, 16'd12699, 16'd14748, 16'd50560, 16'd15577, 16'd57098, 16'd43712, 16'd13123, 16'd7136, 16'd58917});
	test_expansion(128'h65e9e7f91c23c9fe20089f1d25035003, {16'd53996, 16'd22902, 16'd15745, 16'd32065, 16'd25988, 16'd46815, 16'd5063, 16'd2734, 16'd4803, 16'd6129, 16'd30553, 16'd49570, 16'd964, 16'd48929, 16'd57774, 16'd57569, 16'd40015, 16'd43167, 16'd28548, 16'd13225, 16'd2802, 16'd51470, 16'd32864, 16'd227, 16'd971, 16'd10397});
	test_expansion(128'hef2d2ad95c1407ef2524de3844082d93, {16'd65357, 16'd42592, 16'd25067, 16'd43007, 16'd14475, 16'd35701, 16'd56162, 16'd64229, 16'd55379, 16'd26929, 16'd13126, 16'd50211, 16'd33060, 16'd34808, 16'd5539, 16'd6923, 16'd45195, 16'd42102, 16'd60413, 16'd31482, 16'd25650, 16'd18265, 16'd4024, 16'd59230, 16'd35011, 16'd58163});
	test_expansion(128'hd080e8ab652ee55db2a608fbfc3a59c4, {16'd20183, 16'd21167, 16'd34350, 16'd65265, 16'd52414, 16'd53716, 16'd20813, 16'd30634, 16'd19951, 16'd49870, 16'd29850, 16'd54110, 16'd47195, 16'd44314, 16'd16096, 16'd61375, 16'd55165, 16'd19847, 16'd53795, 16'd18271, 16'd43519, 16'd49991, 16'd32325, 16'd3487, 16'd56559, 16'd31256});
	test_expansion(128'hdbebf8c7ee5febb2ec08c41efb63dbd7, {16'd42053, 16'd49601, 16'd49105, 16'd54017, 16'd32179, 16'd19122, 16'd55769, 16'd9821, 16'd26994, 16'd65097, 16'd39217, 16'd4137, 16'd31648, 16'd56403, 16'd32657, 16'd37691, 16'd48107, 16'd36831, 16'd48402, 16'd23957, 16'd46614, 16'd40958, 16'd24344, 16'd11358, 16'd48127, 16'd9955});
	test_expansion(128'h8765e19af9beefddbf52c03790ad3458, {16'd51364, 16'd9135, 16'd40793, 16'd40241, 16'd62826, 16'd15129, 16'd58328, 16'd19205, 16'd27759, 16'd52275, 16'd20522, 16'd20717, 16'd33959, 16'd21406, 16'd44029, 16'd34982, 16'd58502, 16'd55025, 16'd30512, 16'd23173, 16'd54716, 16'd14739, 16'd60892, 16'd60390, 16'd47718, 16'd11039});
	test_expansion(128'h74e13128e742fa4f8d97d79922f19d94, {16'd36606, 16'd58407, 16'd37883, 16'd21511, 16'd38590, 16'd20289, 16'd64787, 16'd579, 16'd14607, 16'd16077, 16'd59502, 16'd35754, 16'd11240, 16'd8292, 16'd59623, 16'd21814, 16'd37565, 16'd44933, 16'd10845, 16'd31104, 16'd59361, 16'd30367, 16'd2922, 16'd63306, 16'd7320, 16'd17300});
	test_expansion(128'ha04573cdbb1cb1b42809911235282eca, {16'd26971, 16'd49281, 16'd16473, 16'd1095, 16'd34945, 16'd53954, 16'd30006, 16'd17402, 16'd52067, 16'd64823, 16'd29079, 16'd56994, 16'd34215, 16'd49005, 16'd6261, 16'd64156, 16'd4606, 16'd29637, 16'd27754, 16'd56485, 16'd65354, 16'd59, 16'd15579, 16'd21896, 16'd42036, 16'd35466});
	test_expansion(128'hcc0bf6b5ac558d978cb64bd4aba89667, {16'd17185, 16'd63999, 16'd13664, 16'd63897, 16'd53172, 16'd504, 16'd24565, 16'd16608, 16'd51355, 16'd15953, 16'd38766, 16'd58683, 16'd15264, 16'd52131, 16'd50547, 16'd62819, 16'd63894, 16'd37715, 16'd55468, 16'd36936, 16'd48517, 16'd35274, 16'd15710, 16'd2850, 16'd399, 16'd54137});
	test_expansion(128'h46435087d8983481dec5aca1a278ca0c, {16'd49720, 16'd37482, 16'd25357, 16'd7983, 16'd37030, 16'd16845, 16'd19169, 16'd48965, 16'd17517, 16'd29220, 16'd20670, 16'd44029, 16'd54870, 16'd6540, 16'd19427, 16'd54055, 16'd55345, 16'd52811, 16'd27457, 16'd57319, 16'd63306, 16'd30523, 16'd4025, 16'd31744, 16'd57685, 16'd26617});
	test_expansion(128'hab458404157216e3b188a3ed8ea85044, {16'd15565, 16'd61968, 16'd11750, 16'd14053, 16'd36239, 16'd32123, 16'd29048, 16'd31981, 16'd4890, 16'd32922, 16'd34383, 16'd58612, 16'd30963, 16'd53595, 16'd30759, 16'd57223, 16'd27120, 16'd50187, 16'd9904, 16'd2579, 16'd10323, 16'd53533, 16'd6712, 16'd53094, 16'd40514, 16'd45374});
	test_expansion(128'h5a5f2e010a596f6eeace4d35276b2f49, {16'd22809, 16'd100, 16'd20484, 16'd41807, 16'd44438, 16'd11626, 16'd7036, 16'd11474, 16'd57618, 16'd52024, 16'd65089, 16'd64174, 16'd56426, 16'd31872, 16'd52494, 16'd45948, 16'd38148, 16'd28663, 16'd45945, 16'd38794, 16'd41043, 16'd62549, 16'd17079, 16'd1049, 16'd24495, 16'd60076});
	test_expansion(128'h4214488ed6d366a5d2c040b0340cbf7f, {16'd58779, 16'd62550, 16'd10512, 16'd56266, 16'd8943, 16'd15605, 16'd38187, 16'd2846, 16'd4538, 16'd44960, 16'd40541, 16'd56309, 16'd13628, 16'd41376, 16'd4058, 16'd49000, 16'd47508, 16'd40286, 16'd48116, 16'd64918, 16'd24666, 16'd48248, 16'd13658, 16'd52804, 16'd45207, 16'd33840});
	test_expansion(128'he59da378ddb45224c599d0a5f97b6fed, {16'd51250, 16'd7593, 16'd358, 16'd39599, 16'd34158, 16'd47836, 16'd28327, 16'd25086, 16'd21872, 16'd57632, 16'd45102, 16'd47523, 16'd48639, 16'd16643, 16'd61840, 16'd37920, 16'd3320, 16'd4738, 16'd26201, 16'd95, 16'd26393, 16'd59933, 16'd10555, 16'd63711, 16'd64293, 16'd49738});
	test_expansion(128'h7826785baeb61471ac6692ca5a860f7e, {16'd15491, 16'd60904, 16'd15826, 16'd59965, 16'd47712, 16'd41324, 16'd51810, 16'd64878, 16'd27862, 16'd31840, 16'd32981, 16'd14221, 16'd3205, 16'd58860, 16'd57448, 16'd42536, 16'd4111, 16'd28292, 16'd52645, 16'd35195, 16'd20772, 16'd64477, 16'd63983, 16'd31316, 16'd17245, 16'd13909});
	test_expansion(128'hb4bff70d9f1d1594439587066b8c81ca, {16'd16000, 16'd19857, 16'd36793, 16'd50078, 16'd17549, 16'd13352, 16'd12520, 16'd11024, 16'd45416, 16'd18649, 16'd61749, 16'd61482, 16'd5354, 16'd23681, 16'd43377, 16'd5720, 16'd33887, 16'd58916, 16'd55152, 16'd14749, 16'd29458, 16'd47932, 16'd14134, 16'd11865, 16'd41702, 16'd60578});
	test_expansion(128'h7b2b4a0307fee38cb6fd7fbb2ce37b76, {16'd26686, 16'd29248, 16'd18047, 16'd55763, 16'd36929, 16'd26710, 16'd7566, 16'd43806, 16'd2817, 16'd36993, 16'd28872, 16'd4320, 16'd56829, 16'd25112, 16'd35886, 16'd51243, 16'd16683, 16'd58276, 16'd30964, 16'd18435, 16'd30334, 16'd59745, 16'd2493, 16'd15445, 16'd39852, 16'd64087});
	test_expansion(128'h5be55eef7624e4b045ce6dd94a2cb836, {16'd48744, 16'd27353, 16'd13490, 16'd49719, 16'd44284, 16'd13017, 16'd54416, 16'd61229, 16'd10091, 16'd46490, 16'd34513, 16'd23355, 16'd58150, 16'd59954, 16'd61615, 16'd21255, 16'd33712, 16'd36886, 16'd36149, 16'd6240, 16'd25670, 16'd36332, 16'd56924, 16'd8527, 16'd24172, 16'd18323});
	test_expansion(128'h102ffc190866aa4e285e2a2ac10c8e56, {16'd12678, 16'd4565, 16'd64473, 16'd64056, 16'd4325, 16'd52700, 16'd12368, 16'd8437, 16'd41812, 16'd4761, 16'd37926, 16'd2835, 16'd9900, 16'd24036, 16'd64630, 16'd14042, 16'd12712, 16'd55025, 16'd10519, 16'd48689, 16'd3657, 16'd55051, 16'd49997, 16'd28887, 16'd59955, 16'd55986});
	test_expansion(128'h6623cb9a47cb3141d654c54fc7cd6aba, {16'd17554, 16'd37756, 16'd32160, 16'd65407, 16'd26564, 16'd7701, 16'd42917, 16'd42248, 16'd41388, 16'd36217, 16'd36722, 16'd17702, 16'd17579, 16'd7196, 16'd44704, 16'd57732, 16'd14557, 16'd13168, 16'd21266, 16'd48809, 16'd55404, 16'd32891, 16'd12918, 16'd55704, 16'd31780, 16'd39414});
	test_expansion(128'haff48ece304966ee9dbeea086aa28121, {16'd46854, 16'd14065, 16'd19612, 16'd53221, 16'd50729, 16'd32649, 16'd19465, 16'd15535, 16'd62892, 16'd3479, 16'd25340, 16'd52559, 16'd50229, 16'd51112, 16'd58854, 16'd25530, 16'd63996, 16'd25577, 16'd60687, 16'd41314, 16'd2445, 16'd61964, 16'd8606, 16'd52029, 16'd59912, 16'd23065});
	test_expansion(128'hd8f8207ec4c8795a1c30a8d494a07773, {16'd34130, 16'd41905, 16'd22987, 16'd62727, 16'd57816, 16'd49329, 16'd21232, 16'd12419, 16'd22880, 16'd16341, 16'd26223, 16'd7470, 16'd35688, 16'd27578, 16'd46443, 16'd51279, 16'd41109, 16'd41101, 16'd30782, 16'd21245, 16'd17157, 16'd61880, 16'd28913, 16'd7834, 16'd59077, 16'd952});
	test_expansion(128'h498fe5649ad345f2a644752ab49e663e, {16'd54269, 16'd30291, 16'd17508, 16'd17105, 16'd20486, 16'd22826, 16'd21263, 16'd342, 16'd17755, 16'd36745, 16'd63041, 16'd56276, 16'd19908, 16'd17446, 16'd11799, 16'd48822, 16'd10735, 16'd13996, 16'd13690, 16'd8329, 16'd24747, 16'd60831, 16'd14140, 16'd29640, 16'd47922, 16'd25164});
	test_expansion(128'hd6eb0475b44a126d9f738bd16d551eb4, {16'd6436, 16'd35497, 16'd32923, 16'd25217, 16'd64089, 16'd54672, 16'd49469, 16'd8876, 16'd15892, 16'd13774, 16'd58070, 16'd14449, 16'd28614, 16'd49104, 16'd34248, 16'd26417, 16'd29498, 16'd14003, 16'd37778, 16'd5490, 16'd36510, 16'd22535, 16'd10384, 16'd43756, 16'd19249, 16'd30150});
	test_expansion(128'hcc697d9b4e1c8b048e248dc7231e4ec9, {16'd45742, 16'd11502, 16'd50590, 16'd48731, 16'd56910, 16'd6041, 16'd46679, 16'd2157, 16'd49708, 16'd49829, 16'd56264, 16'd18061, 16'd13561, 16'd34902, 16'd17223, 16'd44923, 16'd43977, 16'd45889, 16'd16331, 16'd37149, 16'd47518, 16'd6555, 16'd13400, 16'd52975, 16'd51073, 16'd25279});
	test_expansion(128'h08ab0d7314db816c22c8c03a49c43db2, {16'd64144, 16'd19349, 16'd65323, 16'd36406, 16'd2176, 16'd24328, 16'd22185, 16'd34497, 16'd57032, 16'd64759, 16'd26223, 16'd17869, 16'd54625, 16'd6920, 16'd11963, 16'd190, 16'd41876, 16'd38748, 16'd58122, 16'd37860, 16'd57309, 16'd11618, 16'd31661, 16'd60868, 16'd53255, 16'd11718});
	test_expansion(128'hf2e712c93bf322d57436d7e1aa24efdd, {16'd18486, 16'd61650, 16'd56640, 16'd5145, 16'd25120, 16'd64890, 16'd25611, 16'd63841, 16'd49182, 16'd45400, 16'd44917, 16'd59680, 16'd28440, 16'd37673, 16'd5326, 16'd8396, 16'd13239, 16'd24753, 16'd64862, 16'd62159, 16'd19044, 16'd54600, 16'd50637, 16'd5066, 16'd2715, 16'd55462});
	test_expansion(128'h5e5a0f4f07eca99cd453452e0ba9b41a, {16'd49837, 16'd59749, 16'd18065, 16'd51853, 16'd111, 16'd59624, 16'd17304, 16'd42932, 16'd30918, 16'd30531, 16'd56922, 16'd5055, 16'd54520, 16'd44411, 16'd43460, 16'd15904, 16'd25353, 16'd41528, 16'd16767, 16'd34710, 16'd32123, 16'd18615, 16'd32471, 16'd58945, 16'd22517, 16'd60434});
	test_expansion(128'hab50fa86fa7a808460d2d66a148b611b, {16'd16879, 16'd45287, 16'd22148, 16'd2620, 16'd3280, 16'd6400, 16'd846, 16'd15025, 16'd35042, 16'd35630, 16'd36867, 16'd57262, 16'd57349, 16'd1828, 16'd14723, 16'd25831, 16'd49359, 16'd7995, 16'd16998, 16'd612, 16'd20590, 16'd6152, 16'd48671, 16'd7164, 16'd58525, 16'd23344});
	test_expansion(128'h02033ff7513353f1db9deab6bcc803f7, {16'd8735, 16'd50113, 16'd8971, 16'd39422, 16'd22872, 16'd62963, 16'd61256, 16'd4241, 16'd558, 16'd16423, 16'd42592, 16'd49116, 16'd667, 16'd13215, 16'd54218, 16'd17811, 16'd50299, 16'd57514, 16'd36635, 16'd48498, 16'd33250, 16'd24041, 16'd221, 16'd23897, 16'd33832, 16'd58987});
	test_expansion(128'hf5ceb73260c3b6c84f48189d0ed05bc5, {16'd28250, 16'd56963, 16'd51905, 16'd61136, 16'd6711, 16'd54437, 16'd40934, 16'd59830, 16'd24701, 16'd43862, 16'd1631, 16'd38225, 16'd46738, 16'd42904, 16'd19675, 16'd24721, 16'd25552, 16'd59556, 16'd65192, 16'd54119, 16'd3264, 16'd55333, 16'd13728, 16'd8859, 16'd44287, 16'd22263});
	test_expansion(128'hedc410dfb8035ecd88545021f5229be7, {16'd58112, 16'd10247, 16'd60205, 16'd7250, 16'd17898, 16'd49956, 16'd64701, 16'd65032, 16'd13771, 16'd2622, 16'd58962, 16'd41039, 16'd26062, 16'd22012, 16'd8646, 16'd6040, 16'd10849, 16'd16011, 16'd31261, 16'd2448, 16'd46721, 16'd54781, 16'd29784, 16'd53653, 16'd57648, 16'd35850});
	test_expansion(128'h16a41acadddb8c66eee168c816e506fc, {16'd41402, 16'd45673, 16'd65460, 16'd21347, 16'd23947, 16'd47769, 16'd50155, 16'd473, 16'd30463, 16'd35028, 16'd6250, 16'd38760, 16'd6485, 16'd51209, 16'd4615, 16'd43299, 16'd61650, 16'd13303, 16'd6963, 16'd36682, 16'd30925, 16'd53430, 16'd53618, 16'd49191, 16'd47927, 16'd46697});
	test_expansion(128'hc0103e2c9eb6e91b417c570d7685fd26, {16'd52385, 16'd25668, 16'd39317, 16'd50239, 16'd20762, 16'd33264, 16'd64493, 16'd15403, 16'd53698, 16'd3209, 16'd50491, 16'd30164, 16'd25488, 16'd51978, 16'd5612, 16'd17267, 16'd10810, 16'd14346, 16'd47642, 16'd28279, 16'd39827, 16'd5709, 16'd2105, 16'd46816, 16'd41472, 16'd8654});
	test_expansion(128'hb8c8bd1841f2ec2f028f0713ab7d608d, {16'd55876, 16'd56163, 16'd23930, 16'd18877, 16'd53173, 16'd7715, 16'd34877, 16'd37974, 16'd5727, 16'd24512, 16'd41473, 16'd44460, 16'd47860, 16'd60216, 16'd44845, 16'd43115, 16'd1873, 16'd40743, 16'd43443, 16'd1179, 16'd14066, 16'd41867, 16'd37981, 16'd57624, 16'd25433, 16'd48860});
	test_expansion(128'h23933a0b44ed3215f99ec9f7c2d8141c, {16'd20933, 16'd57603, 16'd46123, 16'd54756, 16'd52374, 16'd49598, 16'd7813, 16'd55319, 16'd5225, 16'd54885, 16'd17490, 16'd62757, 16'd63586, 16'd43996, 16'd26291, 16'd62061, 16'd48656, 16'd24519, 16'd28148, 16'd18971, 16'd1648, 16'd55055, 16'd52901, 16'd25604, 16'd21512, 16'd35200});
	test_expansion(128'he77b4ebe3cdc2aff197b752c8c08dc40, {16'd12631, 16'd45511, 16'd59597, 16'd13956, 16'd57657, 16'd27088, 16'd6455, 16'd58427, 16'd4238, 16'd20556, 16'd13817, 16'd41342, 16'd30129, 16'd50129, 16'd61896, 16'd4234, 16'd49345, 16'd38716, 16'd23191, 16'd58119, 16'd6790, 16'd43444, 16'd6733, 16'd14996, 16'd49103, 16'd14595});
	test_expansion(128'hd9c818338f26281caed064ef810e0f77, {16'd30986, 16'd54479, 16'd59321, 16'd17700, 16'd43290, 16'd56933, 16'd29226, 16'd57781, 16'd52918, 16'd16509, 16'd7138, 16'd8945, 16'd38182, 16'd7983, 16'd36700, 16'd21927, 16'd24565, 16'd56399, 16'd2067, 16'd37111, 16'd4929, 16'd22174, 16'd35210, 16'd39284, 16'd38412, 16'd17508});
	test_expansion(128'h29153bdeec3fe537a062953d9371063d, {16'd8731, 16'd31310, 16'd30576, 16'd25447, 16'd29333, 16'd24208, 16'd40857, 16'd8917, 16'd33672, 16'd55683, 16'd19870, 16'd43828, 16'd12773, 16'd14074, 16'd26391, 16'd39323, 16'd38407, 16'd59086, 16'd21867, 16'd61965, 16'd40721, 16'd6420, 16'd7816, 16'd19587, 16'd24360, 16'd22225});
	test_expansion(128'hb18754f6de15ccd8903f73ea5a990475, {16'd21942, 16'd71, 16'd15034, 16'd39413, 16'd65309, 16'd58833, 16'd29633, 16'd49146, 16'd40912, 16'd25448, 16'd12018, 16'd3899, 16'd61308, 16'd30632, 16'd37916, 16'd57222, 16'd21216, 16'd43816, 16'd43013, 16'd17744, 16'd24909, 16'd28537, 16'd41467, 16'd13557, 16'd42143, 16'd51131});
	test_expansion(128'h654798e8eee0ee569928f07281ae73d1, {16'd38762, 16'd11091, 16'd5584, 16'd49270, 16'd48154, 16'd29008, 16'd22291, 16'd18511, 16'd50036, 16'd26310, 16'd65193, 16'd34951, 16'd45749, 16'd32246, 16'd23682, 16'd55159, 16'd59149, 16'd50184, 16'd5136, 16'd13926, 16'd6938, 16'd47742, 16'd58818, 16'd5484, 16'd14542, 16'd26875});
	test_expansion(128'hac42af44f2fac5665fa6751162e5ff97, {16'd13681, 16'd55276, 16'd2174, 16'd57273, 16'd4456, 16'd31455, 16'd17330, 16'd32358, 16'd7278, 16'd3537, 16'd44706, 16'd61590, 16'd21760, 16'd26657, 16'd42225, 16'd42451, 16'd60548, 16'd48353, 16'd2131, 16'd62343, 16'd23494, 16'd45695, 16'd35760, 16'd30276, 16'd32018, 16'd36828});
	test_expansion(128'hd73dfc2ece0052f6a7a6cbe8ac3ae0a3, {16'd56379, 16'd34609, 16'd63651, 16'd47705, 16'd11191, 16'd24914, 16'd29132, 16'd48227, 16'd42454, 16'd18533, 16'd41403, 16'd65242, 16'd34414, 16'd61280, 16'd18755, 16'd39207, 16'd36247, 16'd31577, 16'd46060, 16'd44697, 16'd58524, 16'd20300, 16'd58288, 16'd4455, 16'd63264, 16'd40563});
	test_expansion(128'h6f8d260f3cfd2d3492be5da423f7c2e5, {16'd31060, 16'd6777, 16'd57973, 16'd48666, 16'd1526, 16'd53908, 16'd32837, 16'd61706, 16'd56847, 16'd50814, 16'd22600, 16'd36716, 16'd63411, 16'd1166, 16'd21137, 16'd34177, 16'd59522, 16'd57693, 16'd61927, 16'd21404, 16'd43143, 16'd49263, 16'd27825, 16'd39346, 16'd61692, 16'd12554});
	test_expansion(128'hd9a853e1f2ff976a3e65bf05df0bdbe0, {16'd14, 16'd20547, 16'd25509, 16'd49928, 16'd50921, 16'd44874, 16'd36541, 16'd15016, 16'd1984, 16'd49, 16'd4942, 16'd4520, 16'd40493, 16'd32568, 16'd7443, 16'd32312, 16'd60146, 16'd38664, 16'd29494, 16'd40491, 16'd21036, 16'd57435, 16'd26208, 16'd41829, 16'd64531, 16'd18398});
	test_expansion(128'hfb18b2bcf65a0dc1e7ed3fcf48ecf0a3, {16'd10790, 16'd8100, 16'd41689, 16'd3272, 16'd46270, 16'd9090, 16'd17882, 16'd3804, 16'd54632, 16'd38608, 16'd8009, 16'd64598, 16'd20142, 16'd50109, 16'd49480, 16'd24095, 16'd2167, 16'd28914, 16'd35021, 16'd7294, 16'd14515, 16'd6372, 16'd56677, 16'd47898, 16'd21193, 16'd41822});
	test_expansion(128'hb47af2419720d72eb925a24d7c4ef5ab, {16'd14318, 16'd36297, 16'd41676, 16'd15187, 16'd56696, 16'd61085, 16'd29951, 16'd27514, 16'd24732, 16'd28975, 16'd29852, 16'd32647, 16'd23380, 16'd63585, 16'd48358, 16'd15793, 16'd21007, 16'd40091, 16'd62369, 16'd5094, 16'd15189, 16'd4101, 16'd1066, 16'd22675, 16'd36381, 16'd606});
	test_expansion(128'h7f2f77daf09b3275292ce5b1f541c62f, {16'd62872, 16'd6202, 16'd62875, 16'd38358, 16'd57799, 16'd16851, 16'd49754, 16'd59751, 16'd60465, 16'd7943, 16'd5406, 16'd4052, 16'd26948, 16'd52135, 16'd22467, 16'd23338, 16'd41723, 16'd64021, 16'd22565, 16'd22778, 16'd10014, 16'd62834, 16'd39360, 16'd32044, 16'd28378, 16'd6544});
	test_expansion(128'h44b956989174bb546df1a152bfdc3fb2, {16'd52214, 16'd51310, 16'd298, 16'd46432, 16'd47058, 16'd49110, 16'd12509, 16'd35228, 16'd12899, 16'd60965, 16'd47222, 16'd26101, 16'd56534, 16'd2063, 16'd57193, 16'd8844, 16'd56727, 16'd42974, 16'd21328, 16'd42606, 16'd30293, 16'd38381, 16'd37500, 16'd30682, 16'd48427, 16'd40220});
	test_expansion(128'hc1d30e6c3a69a15b9188f01a311759b8, {16'd55930, 16'd42506, 16'd32630, 16'd2719, 16'd49603, 16'd57118, 16'd64679, 16'd55960, 16'd21442, 16'd756, 16'd29482, 16'd27278, 16'd30026, 16'd30899, 16'd1116, 16'd54682, 16'd57028, 16'd53335, 16'd32673, 16'd57583, 16'd51586, 16'd34661, 16'd65274, 16'd49187, 16'd2930, 16'd24809});
	test_expansion(128'heeab233eaebb5cccfc8fe713f4f8bf86, {16'd11013, 16'd41205, 16'd1234, 16'd12430, 16'd26931, 16'd39014, 16'd41592, 16'd23205, 16'd8801, 16'd59541, 16'd27589, 16'd52390, 16'd8949, 16'd40802, 16'd10813, 16'd20432, 16'd42603, 16'd60621, 16'd17377, 16'd20018, 16'd18299, 16'd58825, 16'd33144, 16'd4208, 16'd29875, 16'd18552});
	test_expansion(128'heda64de7ee41875dc01a0a77ebb5008b, {16'd54710, 16'd59128, 16'd29106, 16'd17270, 16'd46241, 16'd39291, 16'd62497, 16'd13451, 16'd53934, 16'd33603, 16'd59651, 16'd11907, 16'd34727, 16'd36509, 16'd26744, 16'd2385, 16'd41447, 16'd43021, 16'd53599, 16'd35744, 16'd34770, 16'd52289, 16'd55599, 16'd55017, 16'd55804, 16'd64689});
	test_expansion(128'h7c993b6a3068073f2b7da969c99a2950, {16'd18631, 16'd24790, 16'd968, 16'd27336, 16'd40138, 16'd63275, 16'd23322, 16'd63100, 16'd17312, 16'd64807, 16'd21839, 16'd22676, 16'd11111, 16'd8314, 16'd29943, 16'd28036, 16'd52064, 16'd21093, 16'd39849, 16'd35394, 16'd11935, 16'd49077, 16'd8839, 16'd2554, 16'd65326, 16'd17418});
	test_expansion(128'h3db0b690664f60fb1a55e67b2133587c, {16'd38824, 16'd36352, 16'd8525, 16'd63689, 16'd3482, 16'd39447, 16'd12508, 16'd44217, 16'd38963, 16'd61587, 16'd11803, 16'd53604, 16'd52871, 16'd26831, 16'd4895, 16'd45061, 16'd25299, 16'd28989, 16'd42304, 16'd40379, 16'd34782, 16'd44436, 16'd20579, 16'd38540, 16'd22270, 16'd46273});
	test_expansion(128'h871ca1c37244586f26780c1f5e1ee0db, {16'd25968, 16'd29597, 16'd1129, 16'd14246, 16'd44149, 16'd9209, 16'd44946, 16'd61609, 16'd10097, 16'd48893, 16'd63580, 16'd43679, 16'd24713, 16'd33049, 16'd16016, 16'd58945, 16'd29709, 16'd4707, 16'd39571, 16'd52079, 16'd15756, 16'd48917, 16'd41464, 16'd12682, 16'd58875, 16'd39327});
	test_expansion(128'hd615a565ca97b86445b602272574fc91, {16'd8132, 16'd21448, 16'd63134, 16'd57979, 16'd62997, 16'd60144, 16'd26894, 16'd65283, 16'd646, 16'd2678, 16'd16986, 16'd3379, 16'd9779, 16'd32365, 16'd24823, 16'd39855, 16'd18424, 16'd29908, 16'd30483, 16'd10731, 16'd42141, 16'd47356, 16'd28618, 16'd27670, 16'd49483, 16'd56912});
	test_expansion(128'hd1ef85762412a1a08ad7c5deb7b6c0be, {16'd53232, 16'd210, 16'd10780, 16'd35435, 16'd32977, 16'd33733, 16'd55783, 16'd42326, 16'd37342, 16'd65396, 16'd26459, 16'd16849, 16'd24487, 16'd35181, 16'd7931, 16'd5772, 16'd61243, 16'd47773, 16'd48464, 16'd47185, 16'd17676, 16'd50763, 16'd24000, 16'd29238, 16'd11322, 16'd12224});
	test_expansion(128'hf89f2696b1722b8dbe97d6cfe69aa5c2, {16'd44278, 16'd30389, 16'd29732, 16'd23353, 16'd37110, 16'd41748, 16'd42372, 16'd13480, 16'd43025, 16'd42445, 16'd13604, 16'd15391, 16'd32980, 16'd37613, 16'd21909, 16'd63142, 16'd47067, 16'd23018, 16'd31448, 16'd63540, 16'd56653, 16'd4992, 16'd8809, 16'd6207, 16'd63298, 16'd10001});
	test_expansion(128'he00eccd5d88d3f6e4ade706d19559784, {16'd9014, 16'd61770, 16'd45057, 16'd36390, 16'd27949, 16'd1157, 16'd23917, 16'd23654, 16'd33086, 16'd65287, 16'd27463, 16'd37602, 16'd58922, 16'd62945, 16'd13698, 16'd22973, 16'd52197, 16'd58219, 16'd38406, 16'd43993, 16'd18529, 16'd14827, 16'd5594, 16'd35544, 16'd47763, 16'd32151});
	test_expansion(128'hce56184aa6987f2c5f9e212f70a81574, {16'd63999, 16'd43189, 16'd48339, 16'd7140, 16'd63257, 16'd26673, 16'd33405, 16'd42684, 16'd50785, 16'd48976, 16'd57836, 16'd36584, 16'd39013, 16'd14813, 16'd20785, 16'd32188, 16'd53857, 16'd32320, 16'd9995, 16'd19452, 16'd7345, 16'd34673, 16'd53822, 16'd23400, 16'd51899, 16'd25142});
	test_expansion(128'h85b78c0e8c2ffabf1c6dea08749a43ec, {16'd3315, 16'd63022, 16'd38930, 16'd39802, 16'd53877, 16'd52214, 16'd34170, 16'd59605, 16'd33549, 16'd14530, 16'd36206, 16'd26135, 16'd49397, 16'd49049, 16'd25747, 16'd20741, 16'd47753, 16'd53606, 16'd23341, 16'd47782, 16'd18538, 16'd36449, 16'd16770, 16'd37052, 16'd10795, 16'd47876});
	test_expansion(128'h8729fde1b78f930c858795e08c14a0da, {16'd30142, 16'd26320, 16'd2189, 16'd58753, 16'd58521, 16'd33030, 16'd12982, 16'd19554, 16'd64556, 16'd34508, 16'd17316, 16'd21019, 16'd44454, 16'd64350, 16'd46259, 16'd1881, 16'd15662, 16'd22399, 16'd14435, 16'd2630, 16'd29746, 16'd25340, 16'd15823, 16'd20365, 16'd10916, 16'd44260});
	test_expansion(128'hd189817e5a80440e30da3cdb48207944, {16'd64907, 16'd33342, 16'd38603, 16'd43560, 16'd58331, 16'd59990, 16'd1383, 16'd51273, 16'd10381, 16'd6351, 16'd4062, 16'd6505, 16'd55413, 16'd29573, 16'd42627, 16'd27706, 16'd9078, 16'd20884, 16'd12229, 16'd17289, 16'd13650, 16'd43426, 16'd26295, 16'd51395, 16'd10952, 16'd47648});
	test_expansion(128'h5192a220ad94ed6d1631d986a39721a7, {16'd61823, 16'd60370, 16'd1941, 16'd52291, 16'd52269, 16'd62028, 16'd28687, 16'd3908, 16'd49110, 16'd18674, 16'd30759, 16'd38021, 16'd44435, 16'd10547, 16'd44924, 16'd14333, 16'd4319, 16'd45475, 16'd47678, 16'd39788, 16'd60389, 16'd59752, 16'd63516, 16'd17211, 16'd11142, 16'd13296});
	test_expansion(128'h86abfaad82cee8c9fef57464bb4f7cf6, {16'd63797, 16'd59533, 16'd12906, 16'd26989, 16'd922, 16'd4382, 16'd42455, 16'd37935, 16'd45578, 16'd59916, 16'd3890, 16'd20089, 16'd49737, 16'd14703, 16'd26411, 16'd51240, 16'd2513, 16'd7472, 16'd55852, 16'd36048, 16'd4569, 16'd28152, 16'd42021, 16'd3354, 16'd10658, 16'd39909});
	test_expansion(128'h23aebb4952fdc65735d0010ba9759f94, {16'd2027, 16'd53734, 16'd46000, 16'd51143, 16'd57120, 16'd25864, 16'd29937, 16'd64416, 16'd24903, 16'd48912, 16'd38559, 16'd41444, 16'd27089, 16'd59600, 16'd28477, 16'd988, 16'd232, 16'd19644, 16'd24938, 16'd13134, 16'd13533, 16'd946, 16'd46707, 16'd46692, 16'd1499, 16'd2026});
	test_expansion(128'hcd00c6c50b5985d08a7cba0bdf470ebc, {16'd29230, 16'd50862, 16'd16506, 16'd15179, 16'd5518, 16'd61367, 16'd44523, 16'd59482, 16'd1255, 16'd55738, 16'd48753, 16'd26021, 16'd3872, 16'd33617, 16'd34169, 16'd21802, 16'd65446, 16'd5339, 16'd50365, 16'd45357, 16'd17193, 16'd52725, 16'd61942, 16'd59988, 16'd14659, 16'd19451});
	test_expansion(128'hb5cd6e2d4d82c88a845ca086f4974cc0, {16'd23888, 16'd19961, 16'd55016, 16'd21167, 16'd54979, 16'd63173, 16'd36071, 16'd55515, 16'd45891, 16'd7640, 16'd51441, 16'd63149, 16'd39148, 16'd47456, 16'd27158, 16'd64447, 16'd14281, 16'd48899, 16'd12186, 16'd18756, 16'd7553, 16'd40189, 16'd61838, 16'd29951, 16'd37406, 16'd43820});
	test_expansion(128'h3531f2a3556f5b2238b2877e73b8c106, {16'd62167, 16'd12577, 16'd21537, 16'd52983, 16'd33412, 16'd9118, 16'd51224, 16'd415, 16'd44027, 16'd41611, 16'd15314, 16'd4204, 16'd64031, 16'd20836, 16'd55705, 16'd63179, 16'd47690, 16'd50375, 16'd21520, 16'd40684, 16'd21698, 16'd35472, 16'd60786, 16'd318, 16'd35492, 16'd16202});
	test_expansion(128'h615f0bf648c3679099debe22fcb22e5f, {16'd53867, 16'd37791, 16'd2000, 16'd5806, 16'd45907, 16'd34993, 16'd9682, 16'd60280, 16'd15452, 16'd30466, 16'd46137, 16'd40342, 16'd61536, 16'd65366, 16'd63089, 16'd56593, 16'd34413, 16'd33696, 16'd43179, 16'd11926, 16'd44975, 16'd41644, 16'd33019, 16'd43564, 16'd57918, 16'd53497});
	test_expansion(128'hcdde39e17df37bac7c738829d4916d7f, {16'd55568, 16'd49569, 16'd4812, 16'd19828, 16'd58664, 16'd26590, 16'd10697, 16'd17103, 16'd25050, 16'd6914, 16'd10964, 16'd44679, 16'd14326, 16'd10030, 16'd57011, 16'd61455, 16'd31637, 16'd19289, 16'd19434, 16'd31150, 16'd56975, 16'd25334, 16'd13187, 16'd22646, 16'd2275, 16'd19277});
	test_expansion(128'h60f1608992e6c2fc13c21fa8bf99c904, {16'd53817, 16'd63687, 16'd44127, 16'd29798, 16'd63339, 16'd19768, 16'd42032, 16'd31363, 16'd37939, 16'd19136, 16'd36193, 16'd44483, 16'd27859, 16'd953, 16'd52008, 16'd5952, 16'd35471, 16'd39601, 16'd59918, 16'd18672, 16'd16688, 16'd33969, 16'd32046, 16'd27525, 16'd18740, 16'd48184});
	test_expansion(128'h6efcc5372eb03186039319d9d84a90a2, {16'd21322, 16'd26880, 16'd19740, 16'd35867, 16'd18251, 16'd1370, 16'd64855, 16'd15424, 16'd32567, 16'd7195, 16'd15081, 16'd59444, 16'd8496, 16'd37977, 16'd28411, 16'd45830, 16'd30896, 16'd16219, 16'd34300, 16'd48960, 16'd27319, 16'd42321, 16'd47635, 16'd1197, 16'd61794, 16'd46221});
	test_expansion(128'h2dceab4c70a7c2ffa0c0c5705d5bda4e, {16'd22794, 16'd10903, 16'd54295, 16'd22103, 16'd5174, 16'd8706, 16'd53990, 16'd24211, 16'd57617, 16'd43147, 16'd43723, 16'd44308, 16'd45295, 16'd33328, 16'd7908, 16'd38288, 16'd60093, 16'd6209, 16'd49635, 16'd34924, 16'd47498, 16'd43602, 16'd53854, 16'd12261, 16'd43716, 16'd35498});
	test_expansion(128'h62a10951b2628b662ab70bd4502be38c, {16'd51593, 16'd4492, 16'd7310, 16'd34812, 16'd48822, 16'd59941, 16'd64773, 16'd53662, 16'd63481, 16'd46102, 16'd19054, 16'd13484, 16'd13934, 16'd28167, 16'd5922, 16'd15129, 16'd15114, 16'd32502, 16'd21671, 16'd27097, 16'd61725, 16'd64632, 16'd32175, 16'd22947, 16'd40771, 16'd16912});
	test_expansion(128'h8d823c8d4368c5b0b2cf7d0aa5a0843b, {16'd50051, 16'd14950, 16'd293, 16'd13506, 16'd3396, 16'd36069, 16'd35575, 16'd54887, 16'd18796, 16'd3228, 16'd58117, 16'd8621, 16'd64809, 16'd47622, 16'd37862, 16'd25584, 16'd22799, 16'd48448, 16'd25129, 16'd56738, 16'd32103, 16'd40499, 16'd61596, 16'd40673, 16'd39501, 16'd6268});
	test_expansion(128'h5fa6caed22ec7716f31103dbd3788dfe, {16'd46053, 16'd13423, 16'd52440, 16'd46749, 16'd58152, 16'd42954, 16'd26873, 16'd43909, 16'd18499, 16'd30267, 16'd36660, 16'd10582, 16'd54465, 16'd3403, 16'd22798, 16'd22153, 16'd61167, 16'd24953, 16'd60017, 16'd27702, 16'd45700, 16'd47297, 16'd54380, 16'd50540, 16'd61840, 16'd11823});
	test_expansion(128'hb0c8bca16d44ec4d1af9ab49204936e3, {16'd63934, 16'd20361, 16'd12595, 16'd6139, 16'd35190, 16'd59745, 16'd50852, 16'd20445, 16'd47216, 16'd59086, 16'd55388, 16'd45175, 16'd4011, 16'd62810, 16'd31234, 16'd42119, 16'd49585, 16'd25377, 16'd7302, 16'd28451, 16'd21448, 16'd43165, 16'd18732, 16'd42288, 16'd53385, 16'd45472});
	test_expansion(128'h25e1fb48ed79f0ab7cd3b15b8c1474b8, {16'd58705, 16'd15451, 16'd61901, 16'd28948, 16'd21249, 16'd44842, 16'd5999, 16'd26269, 16'd48781, 16'd63720, 16'd25916, 16'd55458, 16'd25549, 16'd51247, 16'd55680, 16'd15148, 16'd12966, 16'd435, 16'd1377, 16'd29668, 16'd49623, 16'd30457, 16'd51634, 16'd29063, 16'd57552, 16'd2587});
	test_expansion(128'hd68962d4ace0ec28a8697de635f71efd, {16'd47917, 16'd7300, 16'd50470, 16'd18425, 16'd34684, 16'd17601, 16'd32001, 16'd4885, 16'd30266, 16'd55207, 16'd59131, 16'd27088, 16'd58111, 16'd63024, 16'd49017, 16'd44963, 16'd895, 16'd40126, 16'd41995, 16'd51857, 16'd48533, 16'd16708, 16'd50083, 16'd28146, 16'd42847, 16'd51958});
	test_expansion(128'h28f3bf6b47a2cc65c30a9a05e0af50ae, {16'd7492, 16'd12694, 16'd15815, 16'd26230, 16'd50398, 16'd31455, 16'd22205, 16'd662, 16'd8030, 16'd27508, 16'd20686, 16'd26959, 16'd20416, 16'd64603, 16'd48623, 16'd31170, 16'd64605, 16'd18482, 16'd145, 16'd12671, 16'd9078, 16'd26645, 16'd3285, 16'd43208, 16'd65390, 16'd65282});
	test_expansion(128'h085f12f0e3bcc30c17892e707e8e0309, {16'd48721, 16'd42332, 16'd62718, 16'd15531, 16'd32018, 16'd48957, 16'd20299, 16'd8496, 16'd37596, 16'd61287, 16'd20728, 16'd64079, 16'd26234, 16'd51822, 16'd12453, 16'd2865, 16'd55999, 16'd21012, 16'd46631, 16'd9769, 16'd27105, 16'd49017, 16'd30159, 16'd27138, 16'd24971, 16'd8186});
	test_expansion(128'h80fd9e277b4110c63082141205e7dd04, {16'd47895, 16'd38290, 16'd61669, 16'd2017, 16'd28013, 16'd11989, 16'd39094, 16'd4521, 16'd27367, 16'd45656, 16'd4781, 16'd33667, 16'd40562, 16'd3779, 16'd39261, 16'd62259, 16'd22362, 16'd19898, 16'd31767, 16'd57813, 16'd45906, 16'd38499, 16'd64578, 16'd11430, 16'd40185, 16'd61147});
	test_expansion(128'h844e3989cafb7efde81f386eb43ff8f6, {16'd8631, 16'd41375, 16'd3294, 16'd62938, 16'd54811, 16'd14789, 16'd43061, 16'd4802, 16'd16004, 16'd8891, 16'd44734, 16'd54666, 16'd19784, 16'd10531, 16'd42259, 16'd35838, 16'd11822, 16'd14624, 16'd4191, 16'd44029, 16'd18531, 16'd55471, 16'd20854, 16'd27437, 16'd12176, 16'd57713});
	test_expansion(128'ha7284c84cd73a988cb44aaeb992b7f27, {16'd37981, 16'd52906, 16'd16928, 16'd30711, 16'd47998, 16'd13112, 16'd38952, 16'd9762, 16'd44917, 16'd42927, 16'd14248, 16'd30511, 16'd38705, 16'd41271, 16'd8592, 16'd8875, 16'd22893, 16'd52962, 16'd14240, 16'd23532, 16'd59087, 16'd11749, 16'd32117, 16'd49821, 16'd59894, 16'd63372});
	test_expansion(128'h40b824959327909365b357b81d4df80c, {16'd15241, 16'd10856, 16'd56537, 16'd44286, 16'd54948, 16'd51435, 16'd58849, 16'd17292, 16'd14014, 16'd56999, 16'd34341, 16'd50275, 16'd56627, 16'd22819, 16'd63241, 16'd14603, 16'd64774, 16'd61627, 16'd9264, 16'd49694, 16'd16219, 16'd1844, 16'd49213, 16'd10660, 16'd12123, 16'd26321});
	test_expansion(128'h972d1dfc0a9342c0a5df2a2c91e6da1b, {16'd2077, 16'd40070, 16'd11871, 16'd23258, 16'd25484, 16'd25507, 16'd43777, 16'd28872, 16'd26832, 16'd44288, 16'd24360, 16'd39427, 16'd38934, 16'd27213, 16'd42861, 16'd48580, 16'd30181, 16'd58549, 16'd42741, 16'd41100, 16'd36063, 16'd62514, 16'd23470, 16'd30534, 16'd53793, 16'd33225});
	test_expansion(128'h8d7505275f9454db769ee5067c2c3c0f, {16'd29874, 16'd27630, 16'd26998, 16'd40674, 16'd19890, 16'd29355, 16'd44106, 16'd58419, 16'd49687, 16'd12934, 16'd39150, 16'd18985, 16'd10212, 16'd36389, 16'd50683, 16'd26833, 16'd52810, 16'd9590, 16'd25102, 16'd50743, 16'd53995, 16'd42681, 16'd15025, 16'd39897, 16'd40880, 16'd8047});
	test_expansion(128'h2ca4c1151da285688d9e5bacbe41e780, {16'd40534, 16'd55940, 16'd32365, 16'd34387, 16'd39530, 16'd8619, 16'd13128, 16'd35026, 16'd46145, 16'd6610, 16'd47976, 16'd25620, 16'd26029, 16'd46178, 16'd40716, 16'd15070, 16'd20290, 16'd13913, 16'd26830, 16'd33748, 16'd59658, 16'd36516, 16'd29234, 16'd23918, 16'd27018, 16'd17355});
	test_expansion(128'hfdb2e1e856401ecfed3750434b822496, {16'd58260, 16'd23276, 16'd64676, 16'd11021, 16'd28493, 16'd30396, 16'd9530, 16'd25218, 16'd22888, 16'd43040, 16'd17913, 16'd46325, 16'd25991, 16'd61364, 16'd32628, 16'd40373, 16'd17519, 16'd60988, 16'd35965, 16'd11401, 16'd15158, 16'd37345, 16'd36164, 16'd50599, 16'd52794, 16'd44438});
	test_expansion(128'h19f4d99147ac47b8f416643bae958326, {16'd44148, 16'd54254, 16'd47924, 16'd44695, 16'd22236, 16'd12694, 16'd54351, 16'd45772, 16'd43808, 16'd22192, 16'd42431, 16'd3900, 16'd25489, 16'd60083, 16'd62504, 16'd26079, 16'd7718, 16'd9796, 16'd4674, 16'd50497, 16'd7503, 16'd54437, 16'd53359, 16'd36377, 16'd4661, 16'd47663});
	test_expansion(128'he94023485d593eb54306ba735b62fd40, {16'd24554, 16'd64535, 16'd21979, 16'd57001, 16'd23875, 16'd23662, 16'd61757, 16'd43502, 16'd20783, 16'd53506, 16'd12206, 16'd29768, 16'd31378, 16'd3300, 16'd46536, 16'd9727, 16'd14045, 16'd5630, 16'd55632, 16'd31056, 16'd1936, 16'd22019, 16'd48862, 16'd59695, 16'd54397, 16'd34998});
	test_expansion(128'h8bfb4545e346d8d41e158ebcad8bfd55, {16'd14712, 16'd38540, 16'd64683, 16'd4318, 16'd36949, 16'd14506, 16'd48313, 16'd61942, 16'd44503, 16'd41400, 16'd45084, 16'd12486, 16'd59399, 16'd5712, 16'd28890, 16'd17870, 16'd40411, 16'd21054, 16'd4096, 16'd34613, 16'd22152, 16'd5087, 16'd64912, 16'd42178, 16'd42505, 16'd39293});
	test_expansion(128'h1078a17e6a8d9c5aedd85c7f861ff334, {16'd39816, 16'd12305, 16'd3220, 16'd14878, 16'd58514, 16'd15105, 16'd48927, 16'd35082, 16'd55181, 16'd25479, 16'd19027, 16'd4544, 16'd9927, 16'd26206, 16'd11591, 16'd6200, 16'd65056, 16'd63597, 16'd3080, 16'd23842, 16'd25017, 16'd27761, 16'd65029, 16'd37085, 16'd63242, 16'd1419});
	test_expansion(128'h0b9e6c62375d554341a42c08c061ddac, {16'd56382, 16'd42226, 16'd64123, 16'd59522, 16'd59106, 16'd59091, 16'd38488, 16'd52136, 16'd39392, 16'd64812, 16'd49864, 16'd60061, 16'd53768, 16'd5685, 16'd25372, 16'd22178, 16'd3318, 16'd18998, 16'd48582, 16'd12218, 16'd63347, 16'd56060, 16'd37886, 16'd16184, 16'd30926, 16'd61876});
	test_expansion(128'h360539d1af0f9c37a2fc0d571ef5e9d9, {16'd27153, 16'd16487, 16'd52361, 16'd47213, 16'd23194, 16'd45763, 16'd18805, 16'd6094, 16'd65174, 16'd61370, 16'd55643, 16'd41785, 16'd15816, 16'd64128, 16'd59783, 16'd5246, 16'd63830, 16'd37497, 16'd40946, 16'd11959, 16'd41285, 16'd13795, 16'd893, 16'd24190, 16'd56618, 16'd8659});
	test_expansion(128'hdad260588c257185b4bdb9cfe82694a7, {16'd34791, 16'd52151, 16'd11332, 16'd35971, 16'd12536, 16'd43116, 16'd59595, 16'd17004, 16'd23898, 16'd695, 16'd27720, 16'd1448, 16'd61161, 16'd5766, 16'd26951, 16'd20022, 16'd42761, 16'd638, 16'd10763, 16'd53569, 16'd41441, 16'd58310, 16'd18427, 16'd30241, 16'd12706, 16'd9964});
	test_expansion(128'h96e1e51ee1aa0243e2fbe4aee4d042f3, {16'd38886, 16'd48350, 16'd4319, 16'd41208, 16'd50874, 16'd42163, 16'd28799, 16'd63241, 16'd43804, 16'd46511, 16'd16930, 16'd46477, 16'd10959, 16'd15095, 16'd43594, 16'd43113, 16'd58855, 16'd60467, 16'd63803, 16'd35877, 16'd9184, 16'd50734, 16'd53192, 16'd54372, 16'd33458, 16'd2572});
	test_expansion(128'h91e788506ad08d76cb74093f45e46de6, {16'd6562, 16'd7698, 16'd20212, 16'd39415, 16'd37087, 16'd41300, 16'd30618, 16'd43213, 16'd11412, 16'd35073, 16'd46698, 16'd26493, 16'd24696, 16'd33642, 16'd49773, 16'd35988, 16'd53855, 16'd49384, 16'd64914, 16'd43895, 16'd34830, 16'd50711, 16'd22943, 16'd31220, 16'd63483, 16'd19582});
	test_expansion(128'h22bcd7a172e0a45b4059e545b0446a4f, {16'd58222, 16'd18434, 16'd14519, 16'd32634, 16'd7400, 16'd36654, 16'd30420, 16'd37607, 16'd28222, 16'd11990, 16'd43653, 16'd32832, 16'd708, 16'd29965, 16'd64063, 16'd38445, 16'd62915, 16'd53111, 16'd26592, 16'd13645, 16'd13303, 16'd47489, 16'd36168, 16'd43857, 16'd41279, 16'd47676});
	test_expansion(128'h5f61d6bf851f8eaf17e7a538f31b1fc5, {16'd46304, 16'd24610, 16'd9476, 16'd9824, 16'd44070, 16'd12469, 16'd32201, 16'd14861, 16'd13756, 16'd64332, 16'd41832, 16'd47443, 16'd29177, 16'd10407, 16'd11625, 16'd34777, 16'd17931, 16'd61251, 16'd61523, 16'd45283, 16'd39498, 16'd14598, 16'd23413, 16'd11177, 16'd49633, 16'd54770});
	test_expansion(128'h693405ab6e455dc959d42766c29d239e, {16'd12326, 16'd45253, 16'd33838, 16'd7140, 16'd36423, 16'd53019, 16'd6023, 16'd28406, 16'd18920, 16'd19913, 16'd55556, 16'd14172, 16'd48568, 16'd11085, 16'd39498, 16'd7301, 16'd18103, 16'd22461, 16'd28560, 16'd1709, 16'd51868, 16'd27995, 16'd33647, 16'd39710, 16'd57000, 16'd17025});
	test_expansion(128'h4a6ebeda495af123d33f0e9adfa1a74e, {16'd59007, 16'd43556, 16'd8500, 16'd27458, 16'd50499, 16'd57089, 16'd40051, 16'd37323, 16'd43058, 16'd2648, 16'd52867, 16'd50762, 16'd28132, 16'd58224, 16'd17204, 16'd35676, 16'd36160, 16'd32293, 16'd60703, 16'd3803, 16'd46268, 16'd26737, 16'd39898, 16'd56678, 16'd37082, 16'd10820});
	test_expansion(128'h8e39898c0923d31b56b19c065e16875c, {16'd44474, 16'd32208, 16'd45893, 16'd17234, 16'd21426, 16'd3643, 16'd32068, 16'd37068, 16'd4935, 16'd59786, 16'd25095, 16'd59513, 16'd47387, 16'd21471, 16'd29234, 16'd64716, 16'd16282, 16'd62394, 16'd6217, 16'd43414, 16'd38912, 16'd1383, 16'd52732, 16'd52959, 16'd47427, 16'd30559});
	test_expansion(128'hbea3c553f97ca58c8fc588b7ca158c5f, {16'd35562, 16'd44912, 16'd45165, 16'd60053, 16'd53852, 16'd51096, 16'd63851, 16'd29562, 16'd56041, 16'd53487, 16'd59888, 16'd11340, 16'd31289, 16'd64249, 16'd18634, 16'd7486, 16'd36113, 16'd30522, 16'd45575, 16'd40309, 16'd46610, 16'd20035, 16'd9499, 16'd13719, 16'd62290, 16'd44045});
	test_expansion(128'hafc5705ab6ff3f8468133dfaccd9ec9a, {16'd6693, 16'd28433, 16'd60380, 16'd27160, 16'd58766, 16'd27348, 16'd991, 16'd53291, 16'd64426, 16'd14788, 16'd13930, 16'd9395, 16'd39217, 16'd58110, 16'd60225, 16'd47728, 16'd26827, 16'd41721, 16'd33773, 16'd60598, 16'd53728, 16'd16959, 16'd37107, 16'd13723, 16'd40238, 16'd48730});
	test_expansion(128'h2ba85b2a18a5d9c5bcc86a17ed30fda0, {16'd25207, 16'd44191, 16'd1169, 16'd63403, 16'd39260, 16'd59487, 16'd18309, 16'd2763, 16'd18554, 16'd51399, 16'd32136, 16'd32496, 16'd11766, 16'd40890, 16'd35101, 16'd52306, 16'd12526, 16'd65158, 16'd26769, 16'd53755, 16'd29893, 16'd48744, 16'd7247, 16'd32118, 16'd495, 16'd43945});
	test_expansion(128'hd5a9049cb5d284fec75763cec0e1656f, {16'd224, 16'd56926, 16'd9355, 16'd40964, 16'd13155, 16'd54345, 16'd16192, 16'd25165, 16'd18535, 16'd54637, 16'd8862, 16'd63879, 16'd12565, 16'd65460, 16'd44612, 16'd46701, 16'd10494, 16'd52289, 16'd8258, 16'd53718, 16'd38795, 16'd12458, 16'd8964, 16'd20443, 16'd53532, 16'd62654});
	test_expansion(128'h881837edd874d946086517709a75f6c4, {16'd60001, 16'd42733, 16'd11478, 16'd50436, 16'd42223, 16'd30159, 16'd4453, 16'd19435, 16'd24639, 16'd28707, 16'd6619, 16'd53958, 16'd479, 16'd31593, 16'd41970, 16'd1367, 16'd37228, 16'd2143, 16'd3148, 16'd37961, 16'd65010, 16'd50750, 16'd59228, 16'd18135, 16'd16723, 16'd30871});
	test_expansion(128'h3ebbd02b1981b8c6c5ba175698c83fa5, {16'd8496, 16'd30849, 16'd5510, 16'd7056, 16'd56497, 16'd53666, 16'd13973, 16'd15618, 16'd21038, 16'd6196, 16'd46649, 16'd59862, 16'd11368, 16'd38489, 16'd45822, 16'd28381, 16'd53295, 16'd25146, 16'd53633, 16'd35769, 16'd6368, 16'd28067, 16'd7936, 16'd14545, 16'd47787, 16'd3920});
	test_expansion(128'h1f8323795430a4013dc447e8dfca14c6, {16'd25657, 16'd21951, 16'd2353, 16'd36697, 16'd47451, 16'd5050, 16'd59052, 16'd65174, 16'd37093, 16'd8690, 16'd48819, 16'd8478, 16'd51720, 16'd24490, 16'd24202, 16'd23854, 16'd24121, 16'd51945, 16'd40145, 16'd31674, 16'd18623, 16'd52105, 16'd3229, 16'd53833, 16'd55840, 16'd32791});
	test_expansion(128'h2d4ca08cc9b58d75d6fbe096f6e03ea5, {16'd61185, 16'd2907, 16'd26385, 16'd23151, 16'd18684, 16'd16984, 16'd29090, 16'd59475, 16'd30398, 16'd17688, 16'd32577, 16'd60574, 16'd10186, 16'd16507, 16'd57301, 16'd54989, 16'd29595, 16'd15548, 16'd53849, 16'd59808, 16'd43921, 16'd61039, 16'd34137, 16'd17176, 16'd40681, 16'd13460});
	test_expansion(128'h6569f136891b9f510e5b5e4877771281, {16'd52840, 16'd38233, 16'd49222, 16'd31433, 16'd62258, 16'd25493, 16'd12958, 16'd48924, 16'd38974, 16'd35531, 16'd29910, 16'd55791, 16'd60891, 16'd31981, 16'd45728, 16'd35903, 16'd25837, 16'd15262, 16'd4175, 16'd52399, 16'd58757, 16'd63529, 16'd61112, 16'd18937, 16'd17408, 16'd4465});
	test_expansion(128'hf0b5c35fcd623a923632be203bce8829, {16'd48161, 16'd5613, 16'd41954, 16'd40422, 16'd27987, 16'd34071, 16'd32989, 16'd65473, 16'd21775, 16'd16496, 16'd27448, 16'd56347, 16'd7717, 16'd58262, 16'd62931, 16'd49818, 16'd52781, 16'd46408, 16'd7425, 16'd24651, 16'd34470, 16'd38586, 16'd16609, 16'd4812, 16'd44135, 16'd24523});
	test_expansion(128'h4ffbecf97fb28e345bd8ded7cc16e93b, {16'd25916, 16'd57336, 16'd35383, 16'd20051, 16'd1281, 16'd53883, 16'd5763, 16'd10888, 16'd46431, 16'd3272, 16'd63808, 16'd57375, 16'd18376, 16'd1789, 16'd21037, 16'd1444, 16'd49404, 16'd23482, 16'd54612, 16'd48790, 16'd21866, 16'd48078, 16'd14947, 16'd11293, 16'd23769, 16'd52717});
	test_expansion(128'h80d067948adf0dd4c135244f7d8e6d6e, {16'd65105, 16'd46485, 16'd14626, 16'd27146, 16'd46440, 16'd18809, 16'd17684, 16'd43923, 16'd40547, 16'd24666, 16'd50025, 16'd880, 16'd44477, 16'd15506, 16'd52112, 16'd44457, 16'd11417, 16'd53648, 16'd48270, 16'd2942, 16'd33774, 16'd51701, 16'd2656, 16'd64504, 16'd64917, 16'd24593});
	test_expansion(128'h0ca7d1fb9778d2885cac4ae231bbe68d, {16'd15249, 16'd13756, 16'd21783, 16'd11778, 16'd27072, 16'd6706, 16'd64785, 16'd19117, 16'd53251, 16'd20071, 16'd42046, 16'd15088, 16'd7265, 16'd41431, 16'd27959, 16'd13875, 16'd249, 16'd18248, 16'd11685, 16'd42854, 16'd42388, 16'd30338, 16'd61263, 16'd27994, 16'd21868, 16'd35477});
	test_expansion(128'h2723b648f1900ab0519d56717bebf3c8, {16'd39039, 16'd46369, 16'd6193, 16'd31307, 16'd32669, 16'd32038, 16'd38328, 16'd59743, 16'd2501, 16'd10336, 16'd52498, 16'd1389, 16'd2544, 16'd34886, 16'd39639, 16'd10622, 16'd20927, 16'd30887, 16'd10927, 16'd64704, 16'd3596, 16'd43125, 16'd44574, 16'd46601, 16'd65422, 16'd27651});
	test_expansion(128'h7502e7e9839cdbd6de3b6f3ba6ce3dc8, {16'd30724, 16'd46325, 16'd50941, 16'd48162, 16'd10750, 16'd27196, 16'd42074, 16'd53821, 16'd10285, 16'd47225, 16'd57460, 16'd5072, 16'd14361, 16'd12036, 16'd20828, 16'd39968, 16'd52964, 16'd59076, 16'd46637, 16'd50791, 16'd50234, 16'd14558, 16'd3064, 16'd41582, 16'd30418, 16'd51755});
	test_expansion(128'hf1284797f9f16fb6a6051e9f060dfd90, {16'd2131, 16'd2697, 16'd23133, 16'd1161, 16'd57623, 16'd5327, 16'd12714, 16'd21437, 16'd1514, 16'd30057, 16'd28085, 16'd50434, 16'd3357, 16'd42708, 16'd61501, 16'd43825, 16'd31641, 16'd60274, 16'd59643, 16'd25152, 16'd29822, 16'd39535, 16'd3990, 16'd43027, 16'd44755, 16'd46926});
	test_expansion(128'h5598b4a60d09a2c75cfd519cbd520b24, {16'd21763, 16'd61545, 16'd55325, 16'd27073, 16'd43138, 16'd2912, 16'd16236, 16'd38254, 16'd1657, 16'd23553, 16'd41704, 16'd64184, 16'd29354, 16'd48149, 16'd7294, 16'd811, 16'd43623, 16'd1094, 16'd2577, 16'd57053, 16'd24966, 16'd28090, 16'd6529, 16'd57013, 16'd9947, 16'd20235});
	test_expansion(128'h5f3514a859caf27fcbbd9ca6f005b811, {16'd30146, 16'd6414, 16'd19305, 16'd30916, 16'd32490, 16'd57491, 16'd22118, 16'd64127, 16'd10153, 16'd27887, 16'd59017, 16'd28185, 16'd32784, 16'd659, 16'd34740, 16'd25207, 16'd869, 16'd18722, 16'd22980, 16'd25788, 16'd22927, 16'd24529, 16'd10518, 16'd1039, 16'd51819, 16'd16758});
	test_expansion(128'hfe824f2e386478452f88f136de3dcb50, {16'd2112, 16'd5352, 16'd59450, 16'd51630, 16'd37198, 16'd62618, 16'd47893, 16'd27086, 16'd62276, 16'd41342, 16'd50849, 16'd15324, 16'd58573, 16'd58312, 16'd29971, 16'd64833, 16'd19430, 16'd24836, 16'd24179, 16'd39507, 16'd39932, 16'd31210, 16'd34762, 16'd33509, 16'd61934, 16'd26218});
	test_expansion(128'h63c1ac3eca0c492b9d299a1bb92d037b, {16'd55544, 16'd26820, 16'd34681, 16'd64254, 16'd41400, 16'd12826, 16'd50943, 16'd6566, 16'd52736, 16'd53387, 16'd60581, 16'd44223, 16'd54480, 16'd60491, 16'd64554, 16'd55057, 16'd64499, 16'd42326, 16'd10911, 16'd35722, 16'd49570, 16'd54487, 16'd41147, 16'd12464, 16'd52231, 16'd31621});
	test_expansion(128'hd6a361cdc334c9c951d59b37dfee289a, {16'd18079, 16'd12255, 16'd4768, 16'd30248, 16'd43205, 16'd41840, 16'd34216, 16'd26762, 16'd17520, 16'd58072, 16'd40845, 16'd23152, 16'd64005, 16'd57969, 16'd59474, 16'd22929, 16'd11495, 16'd60854, 16'd50839, 16'd634, 16'd38038, 16'd52093, 16'd41269, 16'd16804, 16'd48348, 16'd17857});
	test_expansion(128'h5c3cea9ad96f24ee3ce708dc2cf06f5e, {16'd4913, 16'd38845, 16'd24300, 16'd48377, 16'd11897, 16'd62821, 16'd22151, 16'd35924, 16'd17497, 16'd2641, 16'd31756, 16'd59659, 16'd62971, 16'd31613, 16'd16601, 16'd8509, 16'd22357, 16'd11222, 16'd3585, 16'd46607, 16'd10584, 16'd12466, 16'd49670, 16'd49968, 16'd28526, 16'd55297});
	test_expansion(128'h22ae0af21e1e6f2505cfbe0b7611a98c, {16'd14404, 16'd26827, 16'd34552, 16'd46975, 16'd39756, 16'd56134, 16'd43694, 16'd33987, 16'd51419, 16'd30023, 16'd46224, 16'd42136, 16'd24420, 16'd50489, 16'd34140, 16'd33967, 16'd20788, 16'd62844, 16'd718, 16'd56942, 16'd12584, 16'd47546, 16'd64656, 16'd40133, 16'd21825, 16'd65525});
	test_expansion(128'h04380a8c20b029fd68cff7ca03ed4dfb, {16'd5409, 16'd45945, 16'd59674, 16'd15749, 16'd40480, 16'd18867, 16'd5848, 16'd54882, 16'd62947, 16'd18570, 16'd6561, 16'd56993, 16'd44720, 16'd36293, 16'd21014, 16'd1256, 16'd840, 16'd3339, 16'd42331, 16'd42896, 16'd59708, 16'd1352, 16'd15358, 16'd21061, 16'd57533, 16'd23848});
	test_expansion(128'hbf06aa1624884014115974906818592f, {16'd2135, 16'd53130, 16'd58369, 16'd34195, 16'd16888, 16'd13063, 16'd34008, 16'd41322, 16'd41590, 16'd51555, 16'd29572, 16'd56053, 16'd39545, 16'd64037, 16'd32633, 16'd64263, 16'd31820, 16'd50869, 16'd6279, 16'd11731, 16'd30664, 16'd17706, 16'd35793, 16'd64568, 16'd49463, 16'd6222});
	test_expansion(128'h3750b3e2afe66790116bcbfbf35b1881, {16'd41799, 16'd8771, 16'd20277, 16'd57615, 16'd64009, 16'd18787, 16'd43510, 16'd1355, 16'd23103, 16'd35351, 16'd8767, 16'd32887, 16'd50089, 16'd34401, 16'd48030, 16'd6882, 16'd12853, 16'd64460, 16'd48864, 16'd39286, 16'd18239, 16'd1147, 16'd62599, 16'd6960, 16'd48427, 16'd38219});
	test_expansion(128'h9d22267da8e5ef0a9af3fd586acd62dd, {16'd11775, 16'd33163, 16'd22567, 16'd50636, 16'd5954, 16'd36738, 16'd7103, 16'd20946, 16'd56702, 16'd23142, 16'd37567, 16'd4429, 16'd44335, 16'd17152, 16'd58272, 16'd56458, 16'd41866, 16'd63071, 16'd61569, 16'd30261, 16'd12404, 16'd29361, 16'd27393, 16'd7231, 16'd62724, 16'd4170});
	test_expansion(128'he0514d54a21308a0ab9f145cb7ca2ec0, {16'd33781, 16'd54972, 16'd62184, 16'd60300, 16'd44097, 16'd40476, 16'd49147, 16'd48851, 16'd63455, 16'd60105, 16'd2008, 16'd32756, 16'd8361, 16'd9282, 16'd35764, 16'd57671, 16'd51341, 16'd25526, 16'd61142, 16'd41124, 16'd36157, 16'd54654, 16'd24580, 16'd18976, 16'd26271, 16'd10295});
	test_expansion(128'hc5af5dafece7498084a514024122fb19, {16'd569, 16'd24439, 16'd43578, 16'd20376, 16'd26008, 16'd57568, 16'd25465, 16'd48821, 16'd1679, 16'd8775, 16'd64376, 16'd58413, 16'd41018, 16'd38477, 16'd62784, 16'd41441, 16'd42610, 16'd45848, 16'd35131, 16'd19798, 16'd63431, 16'd48037, 16'd58099, 16'd57517, 16'd1963, 16'd35777});
	test_expansion(128'h380def9107fc15e53683871932ae3f08, {16'd32065, 16'd22112, 16'd48304, 16'd1189, 16'd1861, 16'd23184, 16'd6617, 16'd40579, 16'd48429, 16'd50136, 16'd26464, 16'd3538, 16'd1303, 16'd24893, 16'd54179, 16'd18414, 16'd39616, 16'd17091, 16'd31309, 16'd42489, 16'd19122, 16'd33071, 16'd33737, 16'd24985, 16'd33083, 16'd12036});
	test_expansion(128'h99149e194115bc1b12e533d6b66ee1fd, {16'd24016, 16'd10968, 16'd25956, 16'd25665, 16'd46249, 16'd10066, 16'd61696, 16'd24468, 16'd64054, 16'd46547, 16'd14331, 16'd31668, 16'd47508, 16'd57761, 16'd21280, 16'd40525, 16'd9262, 16'd58872, 16'd8118, 16'd57293, 16'd36638, 16'd63930, 16'd52819, 16'd47712, 16'd15717, 16'd26471});
	test_expansion(128'h2421913622506bb0ad996b82de5fc98a, {16'd29232, 16'd20487, 16'd41688, 16'd19865, 16'd11186, 16'd52827, 16'd4069, 16'd19044, 16'd64148, 16'd39703, 16'd32754, 16'd30491, 16'd24521, 16'd16762, 16'd52291, 16'd30988, 16'd48118, 16'd49975, 16'd40054, 16'd2777, 16'd11663, 16'd58195, 16'd47691, 16'd64701, 16'd58106, 16'd21819});
	test_expansion(128'hee8f588c4d5903382a656fa249261119, {16'd23874, 16'd46175, 16'd61960, 16'd23082, 16'd40517, 16'd31544, 16'd39851, 16'd15371, 16'd20326, 16'd14111, 16'd833, 16'd44247, 16'd9117, 16'd3021, 16'd44085, 16'd64876, 16'd50552, 16'd58085, 16'd13658, 16'd36283, 16'd8047, 16'd32447, 16'd1494, 16'd28170, 16'd34302, 16'd12115});
	test_expansion(128'hb614ce07565fa64e628a22b445df0d85, {16'd58364, 16'd27100, 16'd48320, 16'd19391, 16'd26426, 16'd2542, 16'd31632, 16'd35508, 16'd40367, 16'd50994, 16'd46100, 16'd26713, 16'd63281, 16'd61040, 16'd46288, 16'd37995, 16'd29465, 16'd61037, 16'd7192, 16'd49032, 16'd18538, 16'd57171, 16'd21703, 16'd39803, 16'd52949, 16'd32232});
	test_expansion(128'hf27fc121934839e379202df7b9217396, {16'd62511, 16'd25099, 16'd19589, 16'd15455, 16'd52238, 16'd10154, 16'd45382, 16'd56741, 16'd2966, 16'd49410, 16'd41334, 16'd29335, 16'd57926, 16'd57928, 16'd40589, 16'd11253, 16'd17958, 16'd52466, 16'd21004, 16'd48604, 16'd40147, 16'd43894, 16'd43912, 16'd24028, 16'd39993, 16'd21479});
	test_expansion(128'he73b3c9604e8ca864791e40eb24ba46d, {16'd33652, 16'd2579, 16'd22395, 16'd59895, 16'd16590, 16'd10913, 16'd54668, 16'd24733, 16'd50038, 16'd43955, 16'd25667, 16'd61704, 16'd8960, 16'd16232, 16'd53674, 16'd25348, 16'd7257, 16'd8774, 16'd54676, 16'd30128, 16'd12492, 16'd15695, 16'd678, 16'd27378, 16'd5535, 16'd25236});
	test_expansion(128'hb9dcfd329992af61e615a64165623fbb, {16'd33284, 16'd11427, 16'd29177, 16'd44041, 16'd5025, 16'd26375, 16'd13975, 16'd50920, 16'd14641, 16'd37447, 16'd7126, 16'd38838, 16'd17961, 16'd65124, 16'd14958, 16'd33164, 16'd677, 16'd40039, 16'd4860, 16'd25961, 16'd65471, 16'd60344, 16'd53254, 16'd40710, 16'd22328, 16'd26106});
	test_expansion(128'hde57f4e2f1eeccb27e484c98da9722b6, {16'd5468, 16'd45677, 16'd45648, 16'd59576, 16'd9653, 16'd59911, 16'd13876, 16'd38476, 16'd8416, 16'd30071, 16'd40956, 16'd63347, 16'd51373, 16'd29455, 16'd36217, 16'd41912, 16'd43433, 16'd36758, 16'd27332, 16'd60318, 16'd31706, 16'd19106, 16'd493, 16'd19722, 16'd58235, 16'd54232});
	test_expansion(128'hb77e9efdd16944febf4a7cf85d9f6810, {16'd652, 16'd56400, 16'd18445, 16'd30160, 16'd58142, 16'd8562, 16'd57738, 16'd25853, 16'd59915, 16'd37149, 16'd18807, 16'd2394, 16'd7792, 16'd13561, 16'd35106, 16'd26647, 16'd36506, 16'd43900, 16'd22184, 16'd40949, 16'd15716, 16'd6521, 16'd55891, 16'd30943, 16'd23157, 16'd55911});
	test_expansion(128'h02039eb65475631c030df2ae0bf64347, {16'd22159, 16'd59919, 16'd7593, 16'd22893, 16'd64395, 16'd45704, 16'd49223, 16'd10629, 16'd41507, 16'd51190, 16'd14980, 16'd48250, 16'd19773, 16'd37713, 16'd44295, 16'd20888, 16'd61833, 16'd22850, 16'd27567, 16'd10356, 16'd57920, 16'd33586, 16'd5612, 16'd42196, 16'd53964, 16'd16087});
	test_expansion(128'hf04c94999a7c05d6e4282ee43a591e31, {16'd61437, 16'd5027, 16'd49805, 16'd47309, 16'd52622, 16'd51616, 16'd42157, 16'd59495, 16'd44446, 16'd16083, 16'd31913, 16'd56911, 16'd33077, 16'd20370, 16'd59261, 16'd20741, 16'd56690, 16'd15363, 16'd48992, 16'd3125, 16'd48687, 16'd43232, 16'd52624, 16'd28908, 16'd8812, 16'd6912});
	test_expansion(128'h6a56fa84e0d5a0b64e78d79d28816f86, {16'd49226, 16'd50369, 16'd30725, 16'd51696, 16'd43346, 16'd55148, 16'd61169, 16'd53260, 16'd9829, 16'd21038, 16'd24764, 16'd55466, 16'd31195, 16'd27012, 16'd48408, 16'd35894, 16'd15876, 16'd64239, 16'd15198, 16'd30125, 16'd28712, 16'd24245, 16'd14299, 16'd7330, 16'd34095, 16'd7629});
	test_expansion(128'hbdbd15793ff7aabde478c9f39000cccf, {16'd17663, 16'd14809, 16'd6070, 16'd28624, 16'd25424, 16'd61492, 16'd31961, 16'd22749, 16'd24883, 16'd51328, 16'd30472, 16'd62555, 16'd469, 16'd52335, 16'd18371, 16'd9388, 16'd4484, 16'd58696, 16'd5023, 16'd44569, 16'd566, 16'd56937, 16'd5063, 16'd45441, 16'd239, 16'd9986});
	test_expansion(128'h52a3e02a88a404ac5777372245a9fe4d, {16'd64629, 16'd41906, 16'd13140, 16'd60562, 16'd46667, 16'd20499, 16'd16716, 16'd39755, 16'd61753, 16'd33092, 16'd7771, 16'd24683, 16'd26134, 16'd18643, 16'd37705, 16'd28625, 16'd43204, 16'd34509, 16'd27662, 16'd3508, 16'd62367, 16'd14608, 16'd32253, 16'd55461, 16'd59237, 16'd65454});
	test_expansion(128'h9714d0dd1797bb864aeeaaa959a7f2cd, {16'd65170, 16'd32562, 16'd18128, 16'd13499, 16'd30839, 16'd6620, 16'd51357, 16'd26530, 16'd44113, 16'd5171, 16'd45138, 16'd52367, 16'd17843, 16'd11661, 16'd4479, 16'd63863, 16'd5202, 16'd29135, 16'd56736, 16'd12209, 16'd29623, 16'd58132, 16'd60930, 16'd39276, 16'd52451, 16'd45879});
	test_expansion(128'h28d927e30fb2cb165de038494b29b636, {16'd52065, 16'd21636, 16'd64003, 16'd5752, 16'd11879, 16'd1610, 16'd26175, 16'd25726, 16'd46284, 16'd36207, 16'd45902, 16'd32208, 16'd5032, 16'd50120, 16'd10052, 16'd37326, 16'd26414, 16'd44320, 16'd17666, 16'd35825, 16'd24393, 16'd55306, 16'd31218, 16'd60020, 16'd29546, 16'd16891});
	test_expansion(128'h16b551fc7e6496acefe84f58dd7b7359, {16'd40095, 16'd26112, 16'd44656, 16'd47562, 16'd15311, 16'd41526, 16'd30783, 16'd50069, 16'd25644, 16'd28166, 16'd16688, 16'd27170, 16'd24132, 16'd45046, 16'd48180, 16'd3805, 16'd5324, 16'd585, 16'd10368, 16'd64066, 16'd29287, 16'd55817, 16'd19923, 16'd8030, 16'd43045, 16'd21068});
	test_expansion(128'hdb14b0a9f39a42b7d2e4536f1ec48b4c, {16'd45907, 16'd19245, 16'd34210, 16'd41656, 16'd9098, 16'd52400, 16'd26920, 16'd236, 16'd33741, 16'd48228, 16'd43421, 16'd47474, 16'd24540, 16'd22495, 16'd17261, 16'd35720, 16'd21908, 16'd28428, 16'd30238, 16'd3559, 16'd24891, 16'd37734, 16'd2461, 16'd21125, 16'd31253, 16'd10099});
	test_expansion(128'h04d4d76063177c0ada163975620dbc89, {16'd38868, 16'd14546, 16'd47874, 16'd32718, 16'd55069, 16'd51526, 16'd44770, 16'd33589, 16'd34143, 16'd53727, 16'd34696, 16'd19747, 16'd39225, 16'd54798, 16'd48904, 16'd23258, 16'd55553, 16'd23271, 16'd12518, 16'd51634, 16'd35979, 16'd54943, 16'd35712, 16'd9757, 16'd20583, 16'd19859});
	test_expansion(128'hcaf1d836676129a7d1c20fa91ee9db90, {16'd27640, 16'd19242, 16'd55069, 16'd62407, 16'd25330, 16'd50007, 16'd10277, 16'd38112, 16'd10082, 16'd35350, 16'd25295, 16'd34039, 16'd9322, 16'd47561, 16'd15829, 16'd59535, 16'd46898, 16'd41724, 16'd24789, 16'd14008, 16'd9743, 16'd10982, 16'd24863, 16'd51472, 16'd21319, 16'd60079});
	test_expansion(128'h9b8b0fa366e8c8f94b387fb0800d7c8e, {16'd56786, 16'd29897, 16'd34644, 16'd3149, 16'd15583, 16'd50636, 16'd42124, 16'd24750, 16'd44235, 16'd3077, 16'd47829, 16'd51201, 16'd52543, 16'd62129, 16'd51125, 16'd798, 16'd54706, 16'd10794, 16'd9649, 16'd737, 16'd30926, 16'd27753, 16'd5104, 16'd65336, 16'd18647, 16'd25174});
	test_expansion(128'habedea8c38807127960e8fbe3e015178, {16'd10684, 16'd22285, 16'd48645, 16'd27500, 16'd34887, 16'd34660, 16'd29472, 16'd62522, 16'd44897, 16'd3771, 16'd63456, 16'd24950, 16'd16538, 16'd50134, 16'd9480, 16'd27845, 16'd50594, 16'd2592, 16'd56503, 16'd57546, 16'd43280, 16'd10731, 16'd14038, 16'd58713, 16'd31554, 16'd22650});
	test_expansion(128'h438ac89339e6c91728397c5bd745077d, {16'd55547, 16'd17684, 16'd36406, 16'd38835, 16'd28294, 16'd12588, 16'd53708, 16'd53902, 16'd40308, 16'd12238, 16'd27239, 16'd47518, 16'd15357, 16'd60246, 16'd4590, 16'd2909, 16'd5704, 16'd48855, 16'd46335, 16'd19723, 16'd14231, 16'd27694, 16'd55244, 16'd26321, 16'd25807, 16'd61478});
	test_expansion(128'h8435dc148306438c17aa629d8de2abe8, {16'd39123, 16'd55183, 16'd16055, 16'd10744, 16'd7574, 16'd29737, 16'd46295, 16'd2164, 16'd3693, 16'd40732, 16'd39269, 16'd49035, 16'd59664, 16'd17421, 16'd47054, 16'd15488, 16'd57527, 16'd22584, 16'd63394, 16'd53029, 16'd46748, 16'd40910, 16'd13058, 16'd42409, 16'd39079, 16'd23819});
	test_expansion(128'ha84d5f4eee52f063416a2897117a1f5a, {16'd34252, 16'd17051, 16'd50151, 16'd4396, 16'd27157, 16'd51352, 16'd21811, 16'd46514, 16'd24061, 16'd28813, 16'd21535, 16'd4111, 16'd49862, 16'd50117, 16'd43950, 16'd45209, 16'd35279, 16'd45186, 16'd7058, 16'd57788, 16'd3295, 16'd47830, 16'd57264, 16'd33841, 16'd7346, 16'd15387});
	test_expansion(128'h7c15d842d2dbe3ac0231496de3bdee00, {16'd57105, 16'd40629, 16'd52874, 16'd49506, 16'd42362, 16'd64177, 16'd27336, 16'd49399, 16'd63314, 16'd32383, 16'd1071, 16'd48488, 16'd7020, 16'd4382, 16'd46407, 16'd21972, 16'd12994, 16'd49822, 16'd64643, 16'd39755, 16'd24437, 16'd44876, 16'd55620, 16'd30161, 16'd47217, 16'd14812});
	test_expansion(128'ha1a0b4c1ade49afb6fbddabcc32c5426, {16'd13447, 16'd50651, 16'd41788, 16'd28600, 16'd37175, 16'd21450, 16'd19239, 16'd10386, 16'd10027, 16'd20796, 16'd55552, 16'd46483, 16'd17750, 16'd35797, 16'd36130, 16'd49985, 16'd60085, 16'd37613, 16'd56661, 16'd33394, 16'd51421, 16'd44934, 16'd32185, 16'd19689, 16'd15641, 16'd33687});
	test_expansion(128'h6aa9cc449c5be61553c1661ffcb226ed, {16'd51101, 16'd1772, 16'd21333, 16'd294, 16'd9341, 16'd50605, 16'd60775, 16'd325, 16'd17835, 16'd14753, 16'd22035, 16'd40238, 16'd669, 16'd19070, 16'd62887, 16'd44733, 16'd23799, 16'd56058, 16'd45694, 16'd38863, 16'd27075, 16'd10681, 16'd7029, 16'd39720, 16'd14989, 16'd27172});
	test_expansion(128'hd269bcc7c0c7aa23b9cb7f4f4442ad99, {16'd44521, 16'd33728, 16'd3285, 16'd3946, 16'd41009, 16'd38583, 16'd4223, 16'd19752, 16'd5528, 16'd17803, 16'd41630, 16'd26560, 16'd23029, 16'd63535, 16'd39638, 16'd36743, 16'd13788, 16'd49015, 16'd46335, 16'd5593, 16'd49324, 16'd4036, 16'd3326, 16'd34421, 16'd10261, 16'd57702});
	test_expansion(128'h21bdddeb9d8fcf79e1be341bb6cf3104, {16'd39671, 16'd12168, 16'd46843, 16'd4592, 16'd16529, 16'd56172, 16'd52876, 16'd50852, 16'd45880, 16'd32220, 16'd53551, 16'd49992, 16'd19048, 16'd58415, 16'd58137, 16'd39254, 16'd44736, 16'd45722, 16'd2946, 16'd17935, 16'd39790, 16'd3964, 16'd62700, 16'd13003, 16'd5341, 16'd19214});
	test_expansion(128'h004ca4d517b99c9cd22cc6087739705f, {16'd54637, 16'd37830, 16'd7879, 16'd64074, 16'd19624, 16'd32062, 16'd30, 16'd64768, 16'd37953, 16'd29662, 16'd22406, 16'd29869, 16'd6325, 16'd18156, 16'd49763, 16'd11798, 16'd9661, 16'd20106, 16'd42907, 16'd17054, 16'd36834, 16'd44416, 16'd64048, 16'd53709, 16'd33625, 16'd55450});
	test_expansion(128'h8916e986d625870f215541274817c803, {16'd24791, 16'd59885, 16'd18970, 16'd51366, 16'd16278, 16'd45810, 16'd58701, 16'd63046, 16'd15580, 16'd49283, 16'd20341, 16'd588, 16'd47986, 16'd3479, 16'd3753, 16'd54599, 16'd57557, 16'd57748, 16'd47130, 16'd57015, 16'd49379, 16'd55803, 16'd10854, 16'd33473, 16'd568, 16'd24804});
	test_expansion(128'hc80578efcd2dceba40698e9ed8e80216, {16'd26315, 16'd23208, 16'd12631, 16'd12510, 16'd61771, 16'd27532, 16'd54561, 16'd57528, 16'd43274, 16'd24827, 16'd54946, 16'd17478, 16'd6275, 16'd44733, 16'd31242, 16'd10583, 16'd46879, 16'd8306, 16'd21672, 16'd3086, 16'd40589, 16'd45878, 16'd18581, 16'd44590, 16'd44512, 16'd41053});
	test_expansion(128'h686f88a7995afb2b7ff93e7f2398400a, {16'd40660, 16'd42460, 16'd27187, 16'd53747, 16'd22419, 16'd16917, 16'd50796, 16'd9442, 16'd54996, 16'd47532, 16'd40663, 16'd17213, 16'd56569, 16'd23686, 16'd46476, 16'd9298, 16'd31423, 16'd34359, 16'd49801, 16'd55935, 16'd19831, 16'd24531, 16'd38772, 16'd50769, 16'd28670, 16'd41351});
	test_expansion(128'h047b7dcb6d229d29ec47ad62e39da649, {16'd44004, 16'd14809, 16'd49928, 16'd51041, 16'd4854, 16'd36781, 16'd16951, 16'd39911, 16'd42698, 16'd62017, 16'd17607, 16'd12632, 16'd136, 16'd64973, 16'd13926, 16'd12969, 16'd64580, 16'd53334, 16'd47549, 16'd11460, 16'd48249, 16'd20404, 16'd36925, 16'd1585, 16'd3516, 16'd16558});
	test_expansion(128'h58e5ac621684ecd5f9cf4f0fbae0bca0, {16'd4767, 16'd7348, 16'd44713, 16'd60507, 16'd22481, 16'd42941, 16'd57743, 16'd13099, 16'd13390, 16'd20853, 16'd863, 16'd3587, 16'd54206, 16'd12100, 16'd48140, 16'd37534, 16'd47734, 16'd13759, 16'd60712, 16'd28032, 16'd11153, 16'd11398, 16'd16834, 16'd7024, 16'd8318, 16'd30734});
	test_expansion(128'h94993e9c0182531999150453144ad6e5, {16'd56490, 16'd49686, 16'd39952, 16'd57184, 16'd25866, 16'd16352, 16'd47045, 16'd15859, 16'd64351, 16'd35002, 16'd19639, 16'd12542, 16'd53244, 16'd52620, 16'd62276, 16'd38355, 16'd37186, 16'd31153, 16'd48149, 16'd56840, 16'd28427, 16'd44481, 16'd4519, 16'd57167, 16'd49331, 16'd55690});
	test_expansion(128'hac7067ef2b98289a4db53deda66aa45f, {16'd849, 16'd38813, 16'd50924, 16'd38372, 16'd52559, 16'd9858, 16'd23027, 16'd58707, 16'd56827, 16'd36388, 16'd62753, 16'd43404, 16'd8791, 16'd23671, 16'd47474, 16'd58402, 16'd8262, 16'd59943, 16'd11708, 16'd33474, 16'd18398, 16'd56377, 16'd17432, 16'd12593, 16'd46985, 16'd34777});
	test_expansion(128'had82e1e895169d623caaadc94a040ffb, {16'd53435, 16'd63311, 16'd61691, 16'd7109, 16'd397, 16'd33878, 16'd22327, 16'd31756, 16'd19065, 16'd13401, 16'd14858, 16'd20876, 16'd33002, 16'd43562, 16'd17896, 16'd58525, 16'd45543, 16'd38230, 16'd42322, 16'd5214, 16'd11918, 16'd9213, 16'd20817, 16'd19377, 16'd25725, 16'd30914});
	test_expansion(128'h8faf049d25365b1c79076ec9e18c45ba, {16'd4341, 16'd33596, 16'd4983, 16'd27787, 16'd25223, 16'd5718, 16'd14822, 16'd50646, 16'd55546, 16'd46592, 16'd2764, 16'd58425, 16'd34311, 16'd54905, 16'd61175, 16'd20027, 16'd51512, 16'd33678, 16'd38149, 16'd64643, 16'd29321, 16'd39740, 16'd5414, 16'd64019, 16'd48625, 16'd2880});
	test_expansion(128'h92d2920c8c6be3c2a553f8786c06b1d7, {16'd47310, 16'd37946, 16'd11407, 16'd36326, 16'd63796, 16'd25161, 16'd48571, 16'd41897, 16'd10622, 16'd9455, 16'd18544, 16'd49718, 16'd50908, 16'd50060, 16'd751, 16'd11959, 16'd4205, 16'd10736, 16'd61271, 16'd39988, 16'd14159, 16'd47447, 16'd31253, 16'd54323, 16'd4201, 16'd18315});
	test_expansion(128'h87713e2146c95d70c946489b1cccfada, {16'd50929, 16'd55787, 16'd59033, 16'd41235, 16'd24533, 16'd27591, 16'd59213, 16'd16366, 16'd39331, 16'd19514, 16'd64663, 16'd27685, 16'd22926, 16'd14308, 16'd42350, 16'd37910, 16'd13321, 16'd7350, 16'd63303, 16'd9183, 16'd17402, 16'd56637, 16'd38496, 16'd45478, 16'd26995, 16'd61331});
	test_expansion(128'h39db01566de86745285be619766885c9, {16'd46898, 16'd2892, 16'd9673, 16'd43981, 16'd19387, 16'd27375, 16'd11340, 16'd16368, 16'd52330, 16'd40182, 16'd38522, 16'd50093, 16'd6008, 16'd25042, 16'd58450, 16'd47654, 16'd30624, 16'd25467, 16'd21584, 16'd15871, 16'd65512, 16'd51603, 16'd7122, 16'd9754, 16'd51404, 16'd24331});
	test_expansion(128'h5585e68681ee89348439ff5e34935324, {16'd50069, 16'd53863, 16'd56683, 16'd54269, 16'd22984, 16'd16293, 16'd50700, 16'd22673, 16'd22312, 16'd35707, 16'd38980, 16'd53655, 16'd6083, 16'd47987, 16'd63314, 16'd54833, 16'd16472, 16'd2000, 16'd49772, 16'd23811, 16'd26572, 16'd33566, 16'd30924, 16'd62132, 16'd3904, 16'd24129});
	test_expansion(128'h6dc52de223d6a16c5144be3782494ac1, {16'd59135, 16'd58482, 16'd25334, 16'd31978, 16'd54165, 16'd29181, 16'd4143, 16'd28711, 16'd20401, 16'd38236, 16'd28677, 16'd7348, 16'd26435, 16'd29806, 16'd25883, 16'd13540, 16'd19160, 16'd39743, 16'd63070, 16'd41515, 16'd21874, 16'd21341, 16'd9152, 16'd56062, 16'd56035, 16'd58748});
	test_expansion(128'h6c9f24e8df45bc37b46a6505f64ea4e6, {16'd47639, 16'd7375, 16'd24864, 16'd33248, 16'd24724, 16'd54191, 16'd56681, 16'd52724, 16'd17641, 16'd29862, 16'd34598, 16'd17375, 16'd7024, 16'd48899, 16'd28416, 16'd43839, 16'd8986, 16'd54198, 16'd14400, 16'd31272, 16'd504, 16'd48948, 16'd78, 16'd58864, 16'd52775, 16'd18779});
	test_expansion(128'h6de6e130e0b722c438fbddf63a83dae3, {16'd33981, 16'd15180, 16'd9593, 16'd13289, 16'd3483, 16'd61497, 16'd61669, 16'd55320, 16'd10715, 16'd17961, 16'd48740, 16'd1459, 16'd40206, 16'd9369, 16'd16281, 16'd16048, 16'd49688, 16'd31124, 16'd39388, 16'd7134, 16'd28343, 16'd60944, 16'd29376, 16'd31735, 16'd55718, 16'd29381});
	test_expansion(128'heda2df2becf883984575eae4cd75a94b, {16'd60019, 16'd3737, 16'd58683, 16'd24352, 16'd49624, 16'd48329, 16'd33089, 16'd39105, 16'd29897, 16'd27251, 16'd19205, 16'd56924, 16'd23881, 16'd41201, 16'd12649, 16'd56893, 16'd17238, 16'd26641, 16'd16845, 16'd64434, 16'd1489, 16'd30594, 16'd48792, 16'd63789, 16'd48208, 16'd62755});
	test_expansion(128'ha80e3cbe931867ea0309670395c0aada, {16'd35355, 16'd13225, 16'd52916, 16'd16312, 16'd23181, 16'd14949, 16'd6129, 16'd5488, 16'd38920, 16'd25256, 16'd32789, 16'd5869, 16'd15950, 16'd34998, 16'd16542, 16'd52072, 16'd32438, 16'd16613, 16'd1147, 16'd41160, 16'd7824, 16'd37742, 16'd42759, 16'd34410, 16'd16503, 16'd9496});
	test_expansion(128'h0e2a6fc578938d56fdf7ab5a7f9b7c5e, {16'd55528, 16'd51569, 16'd24160, 16'd12767, 16'd53370, 16'd17589, 16'd17074, 16'd28302, 16'd21046, 16'd58308, 16'd63646, 16'd64699, 16'd9642, 16'd23638, 16'd34418, 16'd46381, 16'd26655, 16'd7715, 16'd60995, 16'd52025, 16'd51248, 16'd53091, 16'd21108, 16'd43996, 16'd55885, 16'd64948});
	test_expansion(128'h3aa3840d3cbc97b65a090d32cef1a436, {16'd18282, 16'd54706, 16'd35953, 16'd29498, 16'd33496, 16'd62382, 16'd36289, 16'd29477, 16'd61187, 16'd24313, 16'd45675, 16'd53549, 16'd17462, 16'd12521, 16'd19897, 16'd63554, 16'd57485, 16'd16193, 16'd36905, 16'd5652, 16'd41125, 16'd34400, 16'd29120, 16'd36926, 16'd37522, 16'd14456});
	test_expansion(128'h93bd5a18862594b166d07a9dccb55cfe, {16'd29441, 16'd63645, 16'd18320, 16'd58244, 16'd57233, 16'd15452, 16'd22935, 16'd23188, 16'd30972, 16'd37263, 16'd63762, 16'd5251, 16'd20222, 16'd46666, 16'd55807, 16'd30597, 16'd18833, 16'd54405, 16'd10099, 16'd10294, 16'd12211, 16'd54133, 16'd17080, 16'd63053, 16'd17356, 16'd3879});
	test_expansion(128'hdc6d6e68c14969400f31a1198a912c02, {16'd30129, 16'd35010, 16'd43183, 16'd57577, 16'd5198, 16'd51421, 16'd25930, 16'd4802, 16'd38528, 16'd55787, 16'd18608, 16'd34510, 16'd34697, 16'd20830, 16'd22405, 16'd38763, 16'd54222, 16'd40327, 16'd33049, 16'd47255, 16'd6336, 16'd5807, 16'd8489, 16'd43020, 16'd39122, 16'd56063});
	test_expansion(128'haf7b2c728a18874369f8112317f087a1, {16'd11509, 16'd26227, 16'd53547, 16'd45671, 16'd9974, 16'd50809, 16'd12631, 16'd36481, 16'd6597, 16'd42236, 16'd8012, 16'd31352, 16'd10575, 16'd3020, 16'd38340, 16'd16320, 16'd27455, 16'd44243, 16'd28757, 16'd30263, 16'd37978, 16'd22420, 16'd17608, 16'd43567, 16'd43430, 16'd509});
	test_expansion(128'h9c10ca80e4e53f0b6bd8e0db4c5ad57b, {16'd64229, 16'd10511, 16'd1942, 16'd24896, 16'd14578, 16'd47652, 16'd34632, 16'd5656, 16'd50652, 16'd26535, 16'd61985, 16'd36268, 16'd61702, 16'd7385, 16'd50266, 16'd9063, 16'd56584, 16'd30324, 16'd61980, 16'd41220, 16'd5757, 16'd27491, 16'd28535, 16'd41874, 16'd6068, 16'd45060});
	test_expansion(128'h805ea06d4d10026a2c9df85050624eb4, {16'd33633, 16'd7341, 16'd24787, 16'd52111, 16'd62461, 16'd12220, 16'd13556, 16'd54387, 16'd14014, 16'd41770, 16'd55953, 16'd51741, 16'd52544, 16'd22559, 16'd18400, 16'd21414, 16'd36953, 16'd5999, 16'd34257, 16'd289, 16'd7048, 16'd40605, 16'd2591, 16'd42222, 16'd32725, 16'd33209});
	test_expansion(128'hddb0fbfafd3c898cc1d73bc03954cd4a, {16'd57927, 16'd26382, 16'd3690, 16'd60348, 16'd5641, 16'd37255, 16'd18393, 16'd22266, 16'd45270, 16'd10600, 16'd12300, 16'd33088, 16'd31010, 16'd49718, 16'd64686, 16'd4756, 16'd42923, 16'd10140, 16'd50198, 16'd55224, 16'd48957, 16'd60163, 16'd64979, 16'd19361, 16'd15290, 16'd13751});
	test_expansion(128'h7d3ce4f9464d594ca3006d7d7cb097f2, {16'd61237, 16'd35424, 16'd4205, 16'd60632, 16'd27991, 16'd53864, 16'd40979, 16'd38879, 16'd6205, 16'd15672, 16'd29237, 16'd26499, 16'd38122, 16'd45149, 16'd57123, 16'd61198, 16'd64842, 16'd59127, 16'd29818, 16'd34734, 16'd61805, 16'd61591, 16'd46225, 16'd31130, 16'd27242, 16'd39805});
	test_expansion(128'h06e97e16c94ad4c0aa39500e3241fb81, {16'd24562, 16'd58763, 16'd28149, 16'd15422, 16'd30715, 16'd25296, 16'd47460, 16'd17635, 16'd15578, 16'd60929, 16'd62351, 16'd7171, 16'd38484, 16'd18260, 16'd28944, 16'd36631, 16'd50716, 16'd61360, 16'd59262, 16'd62719, 16'd13906, 16'd50905, 16'd45079, 16'd17610, 16'd56957, 16'd3758});
	test_expansion(128'hde4ea5e395924e8d4ff503b5ce3400ed, {16'd49578, 16'd17158, 16'd34940, 16'd26249, 16'd9205, 16'd64455, 16'd60353, 16'd12537, 16'd22009, 16'd14782, 16'd36472, 16'd53076, 16'd64554, 16'd11604, 16'd42298, 16'd22926, 16'd17925, 16'd53637, 16'd3657, 16'd43666, 16'd46707, 16'd5411, 16'd10513, 16'd24631, 16'd32743, 16'd18501});
	test_expansion(128'ha94596c87d86b151e01aa6e1f97b46f3, {16'd17274, 16'd33824, 16'd14742, 16'd29450, 16'd26498, 16'd41557, 16'd30229, 16'd44919, 16'd37825, 16'd51911, 16'd37432, 16'd18521, 16'd27891, 16'd28402, 16'd61326, 16'd32151, 16'd51198, 16'd61190, 16'd56838, 16'd14362, 16'd20944, 16'd33904, 16'd41612, 16'd50273, 16'd56532, 16'd27931});
	test_expansion(128'h69871f1484af67595002887140842e50, {16'd5362, 16'd24243, 16'd50201, 16'd38045, 16'd3831, 16'd17751, 16'd30530, 16'd49180, 16'd49623, 16'd2329, 16'd4391, 16'd48257, 16'd1245, 16'd43388, 16'd39865, 16'd38466, 16'd31414, 16'd49619, 16'd46905, 16'd55489, 16'd53704, 16'd375, 16'd61746, 16'd49839, 16'd15076, 16'd21407});
	test_expansion(128'h955970ec5862fde5155423b49a0a4d62, {16'd23798, 16'd49880, 16'd39412, 16'd63905, 16'd48663, 16'd26784, 16'd8897, 16'd34436, 16'd27344, 16'd31358, 16'd17609, 16'd52624, 16'd34189, 16'd15514, 16'd26290, 16'd11303, 16'd11530, 16'd4055, 16'd15535, 16'd41840, 16'd20128, 16'd57185, 16'd57560, 16'd44384, 16'd56241, 16'd18707});
	test_expansion(128'h9417f29af1a0a45e64053df272aaf55e, {16'd14344, 16'd25139, 16'd33870, 16'd10478, 16'd1348, 16'd18846, 16'd52601, 16'd4023, 16'd8336, 16'd49464, 16'd8028, 16'd63171, 16'd6545, 16'd58825, 16'd22478, 16'd2710, 16'd32561, 16'd13369, 16'd36820, 16'd25603, 16'd8369, 16'd39863, 16'd54843, 16'd5827, 16'd2084, 16'd55693});
	test_expansion(128'h212e7e458ffa600babe63f5024e2eb53, {16'd4538, 16'd27324, 16'd4114, 16'd62965, 16'd18157, 16'd25639, 16'd14826, 16'd10578, 16'd54596, 16'd39508, 16'd1333, 16'd38141, 16'd29388, 16'd49008, 16'd33032, 16'd46075, 16'd6444, 16'd8266, 16'd56712, 16'd17948, 16'd26989, 16'd13394, 16'd29320, 16'd58714, 16'd54490, 16'd12598});
	test_expansion(128'h7dd52f5e53363f832d3cd423899ec7bd, {16'd30172, 16'd10624, 16'd27956, 16'd34027, 16'd15661, 16'd25068, 16'd2135, 16'd6917, 16'd55602, 16'd44085, 16'd23698, 16'd42056, 16'd23613, 16'd6356, 16'd55898, 16'd64380, 16'd31321, 16'd38695, 16'd11791, 16'd31073, 16'd54408, 16'd46056, 16'd31171, 16'd2172, 16'd54706, 16'd22720});
	test_expansion(128'h566efe5e9edce6d1f7384f17feb03614, {16'd10376, 16'd7282, 16'd40053, 16'd56744, 16'd7189, 16'd9725, 16'd24897, 16'd10080, 16'd1660, 16'd2733, 16'd22136, 16'd49452, 16'd40943, 16'd42327, 16'd37066, 16'd36010, 16'd26675, 16'd39534, 16'd55499, 16'd64860, 16'd51148, 16'd45284, 16'd58504, 16'd9876, 16'd25240, 16'd41564});
	test_expansion(128'hd41ae03d51aebf3cee306a2d27c2d013, {16'd61635, 16'd15406, 16'd3713, 16'd20472, 16'd64622, 16'd23333, 16'd36313, 16'd41988, 16'd28920, 16'd65035, 16'd40984, 16'd32686, 16'd62470, 16'd60173, 16'd50986, 16'd59064, 16'd52825, 16'd30362, 16'd49017, 16'd63393, 16'd21463, 16'd62247, 16'd65181, 16'd4256, 16'd15305, 16'd40434});
	test_expansion(128'h4bf19f813473a87b989ef426d81294e1, {16'd5392, 16'd36913, 16'd55089, 16'd27252, 16'd64528, 16'd36579, 16'd19945, 16'd26017, 16'd48574, 16'd31308, 16'd15501, 16'd18084, 16'd27658, 16'd12987, 16'd31073, 16'd57577, 16'd65486, 16'd54983, 16'd48559, 16'd10806, 16'd46925, 16'd37159, 16'd3085, 16'd36552, 16'd56149, 16'd15889});
	test_expansion(128'hcb178a00847335d131b707e70807fc41, {16'd60330, 16'd17008, 16'd10484, 16'd44385, 16'd44401, 16'd8369, 16'd55206, 16'd30250, 16'd61194, 16'd9609, 16'd29293, 16'd12216, 16'd47607, 16'd13997, 16'd58074, 16'd47499, 16'd27842, 16'd49253, 16'd46738, 16'd44077, 16'd53421, 16'd32910, 16'd38423, 16'd15723, 16'd52512, 16'd64900});
	test_expansion(128'hd473759ac447fa98c20958cd7507c938, {16'd10845, 16'd51572, 16'd55484, 16'd56355, 16'd4264, 16'd55500, 16'd12966, 16'd64611, 16'd15921, 16'd41564, 16'd63669, 16'd17225, 16'd14249, 16'd7920, 16'd4476, 16'd60460, 16'd6543, 16'd36389, 16'd59420, 16'd23503, 16'd46743, 16'd243, 16'd4100, 16'd37166, 16'd32057, 16'd46903});
	test_expansion(128'he2d6dedd1f56426dec1f176493b2f1e0, {16'd46899, 16'd15821, 16'd64253, 16'd61694, 16'd51018, 16'd44547, 16'd25631, 16'd26200, 16'd44775, 16'd40512, 16'd64795, 16'd38007, 16'd3671, 16'd60179, 16'd10318, 16'd36551, 16'd41075, 16'd62672, 16'd12608, 16'd8355, 16'd28490, 16'd50759, 16'd6478, 16'd57279, 16'd36937, 16'd46085});
	test_expansion(128'h45aaefff547b79166dc9f3bc3c593ba2, {16'd64843, 16'd17325, 16'd63467, 16'd7196, 16'd51928, 16'd287, 16'd11244, 16'd40075, 16'd35082, 16'd60917, 16'd43407, 16'd38883, 16'd54347, 16'd57574, 16'd62369, 16'd30393, 16'd52146, 16'd41765, 16'd37546, 16'd24707, 16'd35752, 16'd51260, 16'd60044, 16'd498, 16'd8349, 16'd5182});
	test_expansion(128'h64e2806d6e487219556d9b66e62f52f4, {16'd50125, 16'd63728, 16'd61346, 16'd62672, 16'd40646, 16'd50660, 16'd2843, 16'd54240, 16'd34479, 16'd33279, 16'd50608, 16'd1797, 16'd35558, 16'd51021, 16'd4750, 16'd31190, 16'd13130, 16'd11474, 16'd15833, 16'd9248, 16'd30861, 16'd22085, 16'd37051, 16'd12406, 16'd27148, 16'd34683});
	test_expansion(128'h9afd6a16baa1658805786531f12b0002, {16'd58890, 16'd11353, 16'd4351, 16'd36706, 16'd1586, 16'd17897, 16'd45496, 16'd25768, 16'd60141, 16'd23233, 16'd45350, 16'd32752, 16'd6774, 16'd33777, 16'd61404, 16'd7662, 16'd49725, 16'd45802, 16'd49307, 16'd40866, 16'd21383, 16'd34881, 16'd23434, 16'd64630, 16'd217, 16'd45578});
	test_expansion(128'h2e1ecf77579d2350b97c483956998424, {16'd21750, 16'd39855, 16'd54632, 16'd31868, 16'd64593, 16'd16138, 16'd15386, 16'd21365, 16'd38576, 16'd36773, 16'd32101, 16'd31408, 16'd103, 16'd13991, 16'd12841, 16'd5868, 16'd64015, 16'd37200, 16'd42852, 16'd17614, 16'd19138, 16'd20803, 16'd10106, 16'd54922, 16'd48419, 16'd36861});
	test_expansion(128'h61d4e30ab6cbcf92a5825ec6224fc474, {16'd47421, 16'd44143, 16'd64749, 16'd4535, 16'd59267, 16'd53424, 16'd49351, 16'd18121, 16'd30549, 16'd5331, 16'd40439, 16'd4959, 16'd24321, 16'd4122, 16'd21569, 16'd39882, 16'd55518, 16'd17394, 16'd57243, 16'd6728, 16'd27371, 16'd43254, 16'd4172, 16'd49371, 16'd42335, 16'd11732});
	test_expansion(128'h101041e315781177f3ebd492e007fbf3, {16'd16752, 16'd6794, 16'd38288, 16'd47916, 16'd7508, 16'd22892, 16'd6889, 16'd63276, 16'd31117, 16'd37696, 16'd30879, 16'd42107, 16'd33645, 16'd55953, 16'd39472, 16'd1546, 16'd22000, 16'd61359, 16'd64285, 16'd46258, 16'd54977, 16'd61422, 16'd28273, 16'd20308, 16'd1770, 16'd20718});
	test_expansion(128'h9a402d9ff0db3e928dd058207da7ac32, {16'd19701, 16'd12275, 16'd49947, 16'd29683, 16'd25366, 16'd17547, 16'd53043, 16'd40367, 16'd21604, 16'd11510, 16'd25663, 16'd25793, 16'd38947, 16'd46035, 16'd58753, 16'd22938, 16'd4213, 16'd29744, 16'd42748, 16'd63189, 16'd21534, 16'd14245, 16'd5041, 16'd13046, 16'd2371, 16'd11534});
	test_expansion(128'h7a772da62a12cb9c601831559bf7ff7a, {16'd59110, 16'd18845, 16'd7474, 16'd56159, 16'd5174, 16'd22547, 16'd56567, 16'd46618, 16'd30868, 16'd53610, 16'd19913, 16'd63612, 16'd11618, 16'd63588, 16'd54446, 16'd11096, 16'd62277, 16'd21516, 16'd25995, 16'd17593, 16'd31755, 16'd4480, 16'd22501, 16'd21478, 16'd52960, 16'd12249});
	test_expansion(128'h3aef7bef59e821177b965b70fdc02999, {16'd1952, 16'd46016, 16'd15788, 16'd20109, 16'd62653, 16'd31530, 16'd50498, 16'd7049, 16'd58220, 16'd35903, 16'd43344, 16'd4270, 16'd34374, 16'd15549, 16'd54370, 16'd54028, 16'd51571, 16'd61319, 16'd17948, 16'd58264, 16'd57327, 16'd7149, 16'd42491, 16'd37418, 16'd31678, 16'd47838});
	test_expansion(128'h013eba9c652054f7dfed300fe4df6e12, {16'd43501, 16'd54155, 16'd32387, 16'd55979, 16'd53202, 16'd28241, 16'd49093, 16'd35821, 16'd38036, 16'd42980, 16'd54025, 16'd4628, 16'd20527, 16'd38690, 16'd58848, 16'd375, 16'd6341, 16'd31526, 16'd10995, 16'd18534, 16'd30628, 16'd13331, 16'd42944, 16'd2887, 16'd43707, 16'd31514});
	test_expansion(128'he24d197037444c3cf577e6640024fb91, {16'd54597, 16'd25375, 16'd22560, 16'd30537, 16'd40042, 16'd59161, 16'd26807, 16'd41727, 16'd5301, 16'd21284, 16'd50940, 16'd14929, 16'd30227, 16'd52432, 16'd2244, 16'd38396, 16'd23577, 16'd1312, 16'd18294, 16'd45046, 16'd45906, 16'd6822, 16'd10405, 16'd19483, 16'd15189, 16'd26562});
	test_expansion(128'ha38857285d8ef67851f8b89ff9920ea9, {16'd14028, 16'd7400, 16'd53115, 16'd891, 16'd11319, 16'd18733, 16'd61836, 16'd33035, 16'd33505, 16'd50048, 16'd2590, 16'd40233, 16'd61417, 16'd25978, 16'd29570, 16'd59664, 16'd49525, 16'd26557, 16'd13590, 16'd24992, 16'd14677, 16'd8634, 16'd22613, 16'd9578, 16'd51054, 16'd19984});
	test_expansion(128'h35aec4a2b14129cf535db5cdc28e26af, {16'd18050, 16'd46910, 16'd62042, 16'd18657, 16'd46033, 16'd59166, 16'd7179, 16'd51398, 16'd63137, 16'd26662, 16'd22014, 16'd6708, 16'd14023, 16'd290, 16'd44354, 16'd8829, 16'd10190, 16'd4827, 16'd32858, 16'd32882, 16'd21728, 16'd41892, 16'd57781, 16'd42887, 16'd43387, 16'd53702});
	test_expansion(128'h30b8fd4e496e14774ad1df91c3f533ac, {16'd12778, 16'd7223, 16'd35754, 16'd1497, 16'd4295, 16'd17354, 16'd52880, 16'd33878, 16'd37699, 16'd33647, 16'd20286, 16'd62016, 16'd56229, 16'd1, 16'd53103, 16'd36733, 16'd10805, 16'd33101, 16'd57707, 16'd39726, 16'd43789, 16'd23391, 16'd35357, 16'd59019, 16'd14029, 16'd64226});
	test_expansion(128'h7e7acf496f1c1a516c5fe9c94632b942, {16'd1183, 16'd50381, 16'd42423, 16'd57017, 16'd41876, 16'd65305, 16'd26123, 16'd47850, 16'd2565, 16'd24705, 16'd21174, 16'd18452, 16'd6096, 16'd6445, 16'd40835, 16'd12366, 16'd11372, 16'd39914, 16'd30588, 16'd5992, 16'd17465, 16'd7225, 16'd26349, 16'd17952, 16'd15805, 16'd1645});
	test_expansion(128'he7bdc5dfc077e44bb7fd2efb385a4342, {16'd36930, 16'd29776, 16'd53220, 16'd51255, 16'd24791, 16'd24177, 16'd2903, 16'd17955, 16'd27649, 16'd56204, 16'd40690, 16'd57545, 16'd36796, 16'd35172, 16'd20701, 16'd52785, 16'd15925, 16'd26721, 16'd16090, 16'd11727, 16'd46633, 16'd59215, 16'd34723, 16'd17426, 16'd62295, 16'd32697});
	test_expansion(128'hb61cef1c372befe63132e1fb8b926512, {16'd11707, 16'd13801, 16'd40005, 16'd19401, 16'd50675, 16'd11887, 16'd56565, 16'd23684, 16'd35960, 16'd37255, 16'd48970, 16'd54892, 16'd56687, 16'd60952, 16'd61617, 16'd54630, 16'd37270, 16'd34307, 16'd62905, 16'd36831, 16'd30300, 16'd59211, 16'd12103, 16'd13099, 16'd38931, 16'd32680});
	test_expansion(128'hf47527aecb20d6fdeb01246fae437680, {16'd34944, 16'd11109, 16'd29952, 16'd16146, 16'd22065, 16'd22402, 16'd49012, 16'd1594, 16'd6744, 16'd18624, 16'd16947, 16'd17345, 16'd54158, 16'd34089, 16'd14324, 16'd32013, 16'd60727, 16'd46008, 16'd32449, 16'd5523, 16'd21094, 16'd63761, 16'd1523, 16'd606, 16'd64018, 16'd45179});
	test_expansion(128'h72c278c6a1ac78a2c5591cf4deb97880, {16'd54096, 16'd15404, 16'd55311, 16'd52845, 16'd16155, 16'd5954, 16'd40043, 16'd22907, 16'd33275, 16'd61206, 16'd10491, 16'd23478, 16'd58588, 16'd49309, 16'd5441, 16'd48938, 16'd28425, 16'd2914, 16'd16975, 16'd31131, 16'd11737, 16'd61159, 16'd50670, 16'd42323, 16'd22715, 16'd50109});
	test_expansion(128'h4640ef261efa4f75cecb8ebdec62b17e, {16'd14473, 16'd56081, 16'd61720, 16'd32524, 16'd59186, 16'd10373, 16'd640, 16'd24472, 16'd54629, 16'd32017, 16'd18282, 16'd57783, 16'd40094, 16'd57067, 16'd14752, 16'd13891, 16'd15189, 16'd21012, 16'd60704, 16'd53296, 16'd10935, 16'd51442, 16'd1810, 16'd7314, 16'd13095, 16'd61934});
	test_expansion(128'h173dd82e79b0a3fb7b470e69e1984ee3, {16'd33867, 16'd8365, 16'd4533, 16'd63302, 16'd37275, 16'd32341, 16'd11653, 16'd42462, 16'd24304, 16'd52565, 16'd64056, 16'd64851, 16'd46450, 16'd47495, 16'd12215, 16'd44525, 16'd42605, 16'd47300, 16'd10004, 16'd39338, 16'd24367, 16'd10071, 16'd50321, 16'd24790, 16'd6996, 16'd4973});
	test_expansion(128'hc0476fed1162e88979741c972182e743, {16'd36696, 16'd561, 16'd45839, 16'd35053, 16'd19335, 16'd59894, 16'd32062, 16'd58058, 16'd33257, 16'd41225, 16'd6605, 16'd28110, 16'd17289, 16'd38446, 16'd29320, 16'd26925, 16'd33605, 16'd49424, 16'd65099, 16'd30778, 16'd48077, 16'd2510, 16'd54297, 16'd5236, 16'd33195, 16'd6507});
	test_expansion(128'h836b085ea5a2310e70e52b3c8a8f1ce2, {16'd48742, 16'd58868, 16'd5092, 16'd62293, 16'd12600, 16'd10638, 16'd19334, 16'd56792, 16'd36598, 16'd37416, 16'd41457, 16'd32083, 16'd50441, 16'd13352, 16'd35872, 16'd13254, 16'd13869, 16'd37362, 16'd49109, 16'd64613, 16'd30873, 16'd37735, 16'd44545, 16'd13916, 16'd16906, 16'd6003});
	test_expansion(128'he92e626fc6bbe452f9130c8f347c8a6d, {16'd5308, 16'd11932, 16'd42439, 16'd52247, 16'd18284, 16'd29813, 16'd65189, 16'd64506, 16'd1332, 16'd58466, 16'd42511, 16'd14808, 16'd34094, 16'd53156, 16'd65096, 16'd18543, 16'd14635, 16'd36027, 16'd12021, 16'd26263, 16'd31682, 16'd50407, 16'd3902, 16'd27595, 16'd17504, 16'd27631});
	test_expansion(128'h437f15e64f6f34a8429daae09068ef40, {16'd61599, 16'd57491, 16'd13130, 16'd9543, 16'd48625, 16'd22652, 16'd62911, 16'd14659, 16'd19481, 16'd33809, 16'd8981, 16'd61900, 16'd39483, 16'd9187, 16'd47287, 16'd7306, 16'd31837, 16'd27920, 16'd58103, 16'd60881, 16'd4856, 16'd6906, 16'd22239, 16'd28182, 16'd23151, 16'd44509});
	test_expansion(128'h101f872a82a613529bcf64073c65076b, {16'd32322, 16'd57033, 16'd33813, 16'd17488, 16'd30103, 16'd8484, 16'd63849, 16'd9229, 16'd45693, 16'd61184, 16'd23783, 16'd36960, 16'd60154, 16'd57414, 16'd51769, 16'd56252, 16'd44164, 16'd44525, 16'd11070, 16'd13413, 16'd40199, 16'd8247, 16'd37115, 16'd37025, 16'd23459, 16'd19104});
	test_expansion(128'h783b79c1108a9ec98e1ffd156bee4ef9, {16'd18577, 16'd57404, 16'd5211, 16'd54479, 16'd33449, 16'd25958, 16'd14455, 16'd21377, 16'd57104, 16'd20566, 16'd13534, 16'd6288, 16'd53918, 16'd47509, 16'd37653, 16'd62245, 16'd54762, 16'd3629, 16'd31915, 16'd24383, 16'd26968, 16'd313, 16'd4306, 16'd12992, 16'd42558, 16'd51740});
	test_expansion(128'he0e53a100a1421feddcc46a370b5058f, {16'd8091, 16'd41421, 16'd5679, 16'd21521, 16'd193, 16'd9345, 16'd38962, 16'd35747, 16'd27590, 16'd3988, 16'd53776, 16'd19436, 16'd48964, 16'd58225, 16'd36164, 16'd14085, 16'd40200, 16'd42267, 16'd12764, 16'd1076, 16'd10552, 16'd20915, 16'd3251, 16'd14764, 16'd58421, 16'd31136});
	test_expansion(128'h696f18fb4e947927a864c57b32de750a, {16'd65202, 16'd38720, 16'd8883, 16'd9136, 16'd18645, 16'd8535, 16'd55485, 16'd15616, 16'd10743, 16'd2181, 16'd6725, 16'd51221, 16'd2430, 16'd60602, 16'd29203, 16'd2468, 16'd36155, 16'd8302, 16'd33768, 16'd39695, 16'd34794, 16'd443, 16'd24954, 16'd58777, 16'd54371, 16'd5180});
	test_expansion(128'h5c9bc9c0c4d1777221f1a349a0472bca, {16'd25094, 16'd14849, 16'd1450, 16'd32149, 16'd34871, 16'd65086, 16'd23867, 16'd20345, 16'd12928, 16'd56621, 16'd7343, 16'd55517, 16'd33144, 16'd62531, 16'd24710, 16'd57199, 16'd13163, 16'd35600, 16'd60623, 16'd9141, 16'd38726, 16'd33817, 16'd48851, 16'd11654, 16'd47260, 16'd43009});
	test_expansion(128'he24a1f98173ad9c9679051d32effc37a, {16'd5035, 16'd56538, 16'd25141, 16'd11467, 16'd49246, 16'd40025, 16'd39430, 16'd57444, 16'd52756, 16'd26543, 16'd50183, 16'd65175, 16'd60131, 16'd44626, 16'd26577, 16'd51821, 16'd5241, 16'd48208, 16'd62334, 16'd40892, 16'd32107, 16'd32630, 16'd6860, 16'd7571, 16'd47368, 16'd28785});
	test_expansion(128'h90b52e819f7c97705f3b807fa1c19292, {16'd27874, 16'd55789, 16'd55103, 16'd16531, 16'd51889, 16'd61648, 16'd25344, 16'd42085, 16'd18230, 16'd42940, 16'd30992, 16'd25687, 16'd49789, 16'd23526, 16'd37355, 16'd64406, 16'd10919, 16'd16852, 16'd49514, 16'd40947, 16'd30975, 16'd11618, 16'd909, 16'd63624, 16'd18045, 16'd18468});
	test_expansion(128'hdf5570fe834096b94f2b417df7fd0c29, {16'd44599, 16'd20736, 16'd54789, 16'd8379, 16'd30045, 16'd38350, 16'd8068, 16'd59029, 16'd39873, 16'd65284, 16'd8466, 16'd30787, 16'd37753, 16'd7252, 16'd57249, 16'd23306, 16'd19203, 16'd9578, 16'd14460, 16'd15014, 16'd2457, 16'd62731, 16'd33083, 16'd42888, 16'd5867, 16'd2655});
	test_expansion(128'h87cc850ca354d4435f8366e3302df894, {16'd49821, 16'd10173, 16'd57093, 16'd61114, 16'd13638, 16'd32171, 16'd6202, 16'd24984, 16'd10646, 16'd17261, 16'd9702, 16'd24349, 16'd6275, 16'd17204, 16'd9535, 16'd38072, 16'd8392, 16'd559, 16'd34728, 16'd4332, 16'd45285, 16'd35749, 16'd50486, 16'd59596, 16'd11172, 16'd45520});
	test_expansion(128'h18f712fb6e710731f9339b2aa2e34c93, {16'd20832, 16'd62624, 16'd59763, 16'd10462, 16'd42996, 16'd44567, 16'd15288, 16'd6025, 16'd9206, 16'd14792, 16'd58789, 16'd62247, 16'd56106, 16'd1565, 16'd17537, 16'd5343, 16'd36909, 16'd51926, 16'd63868, 16'd59816, 16'd14249, 16'd12008, 16'd65261, 16'd13647, 16'd1384, 16'd36361});
	test_expansion(128'h14a979982240fa03dcfee61214f44abd, {16'd60730, 16'd11740, 16'd6189, 16'd21050, 16'd45497, 16'd7247, 16'd50252, 16'd55859, 16'd43672, 16'd46629, 16'd17205, 16'd30484, 16'd39665, 16'd25572, 16'd35105, 16'd41905, 16'd62346, 16'd17679, 16'd46198, 16'd29646, 16'd41986, 16'd41215, 16'd44154, 16'd28221, 16'd59406, 16'd62159});
	test_expansion(128'hf6b141aa985abaecbf05b0fbf51241c8, {16'd56335, 16'd34012, 16'd23018, 16'd28956, 16'd63704, 16'd61365, 16'd5469, 16'd7773, 16'd48485, 16'd28263, 16'd32552, 16'd58633, 16'd60264, 16'd46972, 16'd41526, 16'd35563, 16'd12337, 16'd21645, 16'd17409, 16'd22672, 16'd47000, 16'd27711, 16'd14622, 16'd52901, 16'd46206, 16'd1892});
	test_expansion(128'h5040a360c9c29c4d3f480da2d07d41cd, {16'd64626, 16'd63739, 16'd65444, 16'd51675, 16'd15417, 16'd38162, 16'd25142, 16'd64211, 16'd840, 16'd12868, 16'd61799, 16'd25833, 16'd7676, 16'd50340, 16'd59903, 16'd63352, 16'd6305, 16'd28224, 16'd63728, 16'd31656, 16'd64632, 16'd7938, 16'd12053, 16'd45590, 16'd45516, 16'd5688});
	test_expansion(128'hba22ed5bf83f67f6c140ff363e5b7275, {16'd13559, 16'd45921, 16'd57904, 16'd50355, 16'd52072, 16'd7313, 16'd44005, 16'd4029, 16'd55350, 16'd47387, 16'd42210, 16'd20469, 16'd64801, 16'd13516, 16'd57447, 16'd42354, 16'd48943, 16'd48798, 16'd38993, 16'd58123, 16'd32272, 16'd30824, 16'd899, 16'd61078, 16'd15161, 16'd55091});
	test_expansion(128'ha7154edc79a7a39b4c8b18faa2c6c534, {16'd57120, 16'd46007, 16'd53853, 16'd59035, 16'd34083, 16'd59159, 16'd37076, 16'd9612, 16'd25416, 16'd44446, 16'd46398, 16'd39170, 16'd26476, 16'd25663, 16'd29229, 16'd40948, 16'd30045, 16'd16868, 16'd47661, 16'd47333, 16'd17230, 16'd58735, 16'd38930, 16'd63263, 16'd24970, 16'd35577});
	test_expansion(128'h5220f26ddccf0aa522468dce5e95e86b, {16'd9685, 16'd23022, 16'd8687, 16'd41197, 16'd29720, 16'd29847, 16'd55052, 16'd22767, 16'd58223, 16'd54428, 16'd38099, 16'd48115, 16'd10070, 16'd62293, 16'd52043, 16'd65510, 16'd64531, 16'd56577, 16'd60152, 16'd8970, 16'd56477, 16'd65275, 16'd47486, 16'd32937, 16'd47213, 16'd65307});
	test_expansion(128'he85d7182d7718e3b05246c8c1fcdd77c, {16'd40532, 16'd52387, 16'd44332, 16'd43750, 16'd62074, 16'd43978, 16'd49874, 16'd40930, 16'd56222, 16'd47949, 16'd25136, 16'd3313, 16'd61772, 16'd6812, 16'd43624, 16'd6357, 16'd34166, 16'd18140, 16'd58572, 16'd14780, 16'd58384, 16'd35174, 16'd39894, 16'd57249, 16'd33880, 16'd15529});
	test_expansion(128'h3bda071263e55c6d0d44414f2f51d516, {16'd16476, 16'd27930, 16'd47112, 16'd16394, 16'd52056, 16'd12224, 16'd49688, 16'd20851, 16'd64956, 16'd479, 16'd28068, 16'd39495, 16'd15845, 16'd41043, 16'd32981, 16'd29047, 16'd37034, 16'd39431, 16'd12390, 16'd64426, 16'd56621, 16'd57379, 16'd39603, 16'd21478, 16'd37013, 16'd17983});
	test_expansion(128'h2613b7d774b62b2ee8aa125a9237c895, {16'd59617, 16'd4684, 16'd40887, 16'd50461, 16'd57551, 16'd8163, 16'd11678, 16'd8662, 16'd30202, 16'd18266, 16'd6086, 16'd25259, 16'd24638, 16'd18818, 16'd37331, 16'd39358, 16'd56935, 16'd27991, 16'd6198, 16'd10370, 16'd32262, 16'd16344, 16'd38326, 16'd54039, 16'd13805, 16'd39805});
	test_expansion(128'hb5216e8e4f2094e8b9a2dea29960d569, {16'd14514, 16'd22600, 16'd10147, 16'd24552, 16'd7768, 16'd57124, 16'd5319, 16'd53293, 16'd47304, 16'd9797, 16'd37160, 16'd1842, 16'd30186, 16'd42041, 16'd48220, 16'd48357, 16'd49106, 16'd19434, 16'd2672, 16'd9338, 16'd40518, 16'd26815, 16'd47582, 16'd43990, 16'd34113, 16'd3061});
	test_expansion(128'h368297e2f0c28d01ae8892789a5ec95d, {16'd3317, 16'd30637, 16'd62847, 16'd40709, 16'd62723, 16'd22416, 16'd46466, 16'd34030, 16'd26258, 16'd49345, 16'd6818, 16'd58309, 16'd21902, 16'd23454, 16'd22544, 16'd17727, 16'd51520, 16'd23104, 16'd13131, 16'd53032, 16'd23375, 16'd39753, 16'd26349, 16'd14786, 16'd20025, 16'd61796});
	test_expansion(128'he82c2842e4223af207d272723d292e49, {16'd2383, 16'd48359, 16'd55036, 16'd42305, 16'd40296, 16'd19242, 16'd38412, 16'd7587, 16'd59379, 16'd50186, 16'd58323, 16'd4648, 16'd56168, 16'd17033, 16'd39460, 16'd6348, 16'd27315, 16'd9767, 16'd43406, 16'd47418, 16'd8909, 16'd35028, 16'd51647, 16'd36073, 16'd37602, 16'd580});
	test_expansion(128'h22af06e458a5e2468e0f9d1f4ce150b4, {16'd50671, 16'd55667, 16'd15368, 16'd20575, 16'd62115, 16'd42074, 16'd33603, 16'd30764, 16'd50846, 16'd59800, 16'd59316, 16'd1140, 16'd45062, 16'd53502, 16'd17374, 16'd48272, 16'd63375, 16'd54817, 16'd27091, 16'd59351, 16'd56513, 16'd575, 16'd61271, 16'd64150, 16'd512, 16'd24656});
	test_expansion(128'ha4156de7ed479000e1f6ef7f7983e2e3, {16'd49565, 16'd20610, 16'd41872, 16'd57888, 16'd12945, 16'd50217, 16'd45002, 16'd6229, 16'd46110, 16'd9298, 16'd6105, 16'd64487, 16'd40498, 16'd41401, 16'd64561, 16'd56446, 16'd59673, 16'd38309, 16'd12390, 16'd19032, 16'd61735, 16'd12697, 16'd42406, 16'd19859, 16'd56465, 16'd37493});
	test_expansion(128'hb36ebe72943d5989c942e979e87fc2fb, {16'd27184, 16'd13634, 16'd30244, 16'd13497, 16'd64019, 16'd33353, 16'd15327, 16'd64083, 16'd20690, 16'd224, 16'd54475, 16'd27070, 16'd50078, 16'd58498, 16'd46722, 16'd4591, 16'd43534, 16'd19028, 16'd39031, 16'd62627, 16'd14043, 16'd18019, 16'd6472, 16'd23256, 16'd8757, 16'd46864});
	test_expansion(128'h31db280fcd6dd1033e76c6496a54c92d, {16'd36597, 16'd62554, 16'd32154, 16'd57921, 16'd30506, 16'd431, 16'd8359, 16'd5008, 16'd58965, 16'd39192, 16'd54047, 16'd54389, 16'd65522, 16'd11522, 16'd52960, 16'd16079, 16'd53069, 16'd35934, 16'd45147, 16'd7997, 16'd41888, 16'd36950, 16'd20542, 16'd16422, 16'd30927, 16'd56613});
	test_expansion(128'h270921902a335ba9b94f80449cca852f, {16'd14489, 16'd14338, 16'd39860, 16'd2677, 16'd55675, 16'd2460, 16'd31545, 16'd52285, 16'd19875, 16'd35507, 16'd16077, 16'd10432, 16'd27447, 16'd41569, 16'd33070, 16'd15080, 16'd56070, 16'd36170, 16'd51497, 16'd6666, 16'd53158, 16'd16375, 16'd49644, 16'd39387, 16'd56314, 16'd13993});
	test_expansion(128'hd97e4dae0ce3f2bef2c8133797efb882, {16'd53133, 16'd37739, 16'd59164, 16'd7138, 16'd14129, 16'd58986, 16'd21767, 16'd5943, 16'd7969, 16'd5895, 16'd17698, 16'd64585, 16'd24269, 16'd12938, 16'd1587, 16'd39306, 16'd18821, 16'd64158, 16'd59534, 16'd44678, 16'd18358, 16'd18486, 16'd44719, 16'd4693, 16'd63565, 16'd64008});
	test_expansion(128'h011c2defe371b07553f2121362e3c2b1, {16'd34566, 16'd41284, 16'd33569, 16'd60467, 16'd44388, 16'd15432, 16'd9486, 16'd19719, 16'd54247, 16'd22149, 16'd21775, 16'd14305, 16'd10341, 16'd29575, 16'd10194, 16'd10477, 16'd47747, 16'd4510, 16'd36849, 16'd28073, 16'd49899, 16'd6575, 16'd7278, 16'd8459, 16'd16375, 16'd13507});
	test_expansion(128'h199e5d4140d313e33826a3abbe31b3c1, {16'd36092, 16'd34468, 16'd53703, 16'd16044, 16'd10408, 16'd1579, 16'd58761, 16'd1978, 16'd57072, 16'd31162, 16'd13423, 16'd37119, 16'd27862, 16'd592, 16'd1357, 16'd64496, 16'd44393, 16'd20306, 16'd8587, 16'd62177, 16'd621, 16'd62369, 16'd9534, 16'd45498, 16'd65329, 16'd39522});
	test_expansion(128'h3487b80b2578b8a42e8b29e4805d7698, {16'd45001, 16'd22860, 16'd14531, 16'd2695, 16'd21470, 16'd63826, 16'd56136, 16'd2269, 16'd49343, 16'd22439, 16'd19753, 16'd5551, 16'd45953, 16'd47902, 16'd12512, 16'd43617, 16'd38082, 16'd46733, 16'd50021, 16'd42076, 16'd35475, 16'd15579, 16'd33113, 16'd18352, 16'd45859, 16'd36154});
	test_expansion(128'hd5df0818c7721ba6ca0b23256cb72aa9, {16'd15288, 16'd43865, 16'd63243, 16'd16599, 16'd40059, 16'd2895, 16'd38681, 16'd9948, 16'd26818, 16'd16075, 16'd28543, 16'd30778, 16'd47613, 16'd21679, 16'd2706, 16'd30912, 16'd53518, 16'd41343, 16'd58123, 16'd57866, 16'd55111, 16'd47718, 16'd5880, 16'd59561, 16'd59535, 16'd15564});
	test_expansion(128'hf47915b6cc36e7f4dd25c42c9b04ce69, {16'd22019, 16'd379, 16'd4077, 16'd36922, 16'd25574, 16'd53128, 16'd9947, 16'd19514, 16'd29657, 16'd16768, 16'd26792, 16'd59923, 16'd33009, 16'd41855, 16'd14080, 16'd22065, 16'd34457, 16'd35758, 16'd30035, 16'd64454, 16'd33139, 16'd55007, 16'd16684, 16'd58156, 16'd10509, 16'd37384});
	test_expansion(128'h782ea2433c59b9be040a26068ca36f9c, {16'd43168, 16'd10682, 16'd32351, 16'd17444, 16'd42377, 16'd61671, 16'd16306, 16'd21880, 16'd40910, 16'd40439, 16'd11115, 16'd920, 16'd18509, 16'd29100, 16'd3044, 16'd23618, 16'd58698, 16'd50796, 16'd38005, 16'd7210, 16'd62982, 16'd37560, 16'd26095, 16'd698, 16'd8487, 16'd14825});
	test_expansion(128'hd9104cb93ef621bb56f0a01c3e1a9581, {16'd19897, 16'd23963, 16'd40123, 16'd9196, 16'd41544, 16'd9943, 16'd37374, 16'd33377, 16'd53807, 16'd48165, 16'd28654, 16'd37454, 16'd29671, 16'd21371, 16'd62535, 16'd5587, 16'd30209, 16'd37815, 16'd1393, 16'd37548, 16'd62509, 16'd56409, 16'd50862, 16'd10149, 16'd46838, 16'd38183});
	test_expansion(128'hd7102a53eb5579a1c9df97975e333500, {16'd14232, 16'd51533, 16'd53172, 16'd61174, 16'd27098, 16'd5700, 16'd4310, 16'd51909, 16'd56583, 16'd62421, 16'd45839, 16'd48200, 16'd30428, 16'd16823, 16'd49043, 16'd23985, 16'd9218, 16'd39933, 16'd12420, 16'd28294, 16'd25700, 16'd13549, 16'd59241, 16'd6792, 16'd8554, 16'd54020});
	test_expansion(128'h05c129315b39ee784a965e4dc2669bb8, {16'd40114, 16'd40965, 16'd11298, 16'd3899, 16'd63112, 16'd7854, 16'd44611, 16'd65531, 16'd42924, 16'd48946, 16'd52956, 16'd54563, 16'd20348, 16'd27544, 16'd18330, 16'd38646, 16'd23151, 16'd40117, 16'd8944, 16'd3359, 16'd22628, 16'd62348, 16'd44681, 16'd14113, 16'd20122, 16'd60510});
	test_expansion(128'hf13e9ceab7d3349765b299b2b8ee3a3c, {16'd49692, 16'd58999, 16'd30609, 16'd34321, 16'd3165, 16'd14303, 16'd37591, 16'd40411, 16'd38335, 16'd48552, 16'd8948, 16'd4046, 16'd19326, 16'd2642, 16'd30374, 16'd31590, 16'd20195, 16'd12, 16'd30782, 16'd4092, 16'd60845, 16'd10978, 16'd56502, 16'd9932, 16'd60665, 16'd27392});
	test_expansion(128'h74831a62fcf1aaff007a55c9f92d80d2, {16'd23395, 16'd11175, 16'd26009, 16'd65401, 16'd6110, 16'd39868, 16'd10665, 16'd24613, 16'd22717, 16'd10129, 16'd31468, 16'd64004, 16'd42772, 16'd51667, 16'd22019, 16'd11655, 16'd13745, 16'd39034, 16'd29223, 16'd13388, 16'd65420, 16'd33599, 16'd54775, 16'd65166, 16'd50475, 16'd13680});
	test_expansion(128'h791fff0acef814b823ac2c6446bb2d86, {16'd59221, 16'd43607, 16'd53903, 16'd7528, 16'd54982, 16'd54334, 16'd33343, 16'd64960, 16'd25348, 16'd47579, 16'd47190, 16'd15327, 16'd22071, 16'd1912, 16'd4524, 16'd64378, 16'd56947, 16'd53263, 16'd10925, 16'd7078, 16'd56699, 16'd41994, 16'd14701, 16'd964, 16'd58259, 16'd56742});
	test_expansion(128'hdc6c1d584146a3aaf8ff06d6baa51fff, {16'd11211, 16'd41923, 16'd5230, 16'd14386, 16'd32542, 16'd50821, 16'd62846, 16'd53468, 16'd38595, 16'd63941, 16'd14196, 16'd42679, 16'd33089, 16'd26287, 16'd15187, 16'd24029, 16'd34969, 16'd22830, 16'd34623, 16'd10224, 16'd60879, 16'd21266, 16'd59140, 16'd13340, 16'd22795, 16'd4818});
	test_expansion(128'h4436f3201b2cdb792a3f041e7d054500, {16'd6638, 16'd53019, 16'd37898, 16'd20940, 16'd54994, 16'd49324, 16'd24993, 16'd3642, 16'd27702, 16'd23746, 16'd8575, 16'd61530, 16'd60544, 16'd20147, 16'd11404, 16'd38658, 16'd59627, 16'd65262, 16'd20144, 16'd65459, 16'd51697, 16'd64046, 16'd1340, 16'd47052, 16'd60147, 16'd35005});
	test_expansion(128'h14cd8f4fb7851edd35fe6138e0bf8127, {16'd25503, 16'd55061, 16'd37879, 16'd31785, 16'd32901, 16'd15563, 16'd27856, 16'd52100, 16'd12356, 16'd30323, 16'd19512, 16'd55243, 16'd2140, 16'd3170, 16'd61290, 16'd62463, 16'd15653, 16'd23166, 16'd17048, 16'd59754, 16'd1233, 16'd41811, 16'd21274, 16'd39292, 16'd24659, 16'd43553});
	test_expansion(128'haf04610d1e72727a627061058d7b448f, {16'd21874, 16'd22253, 16'd52981, 16'd55698, 16'd57179, 16'd58159, 16'd24719, 16'd61807, 16'd33512, 16'd44508, 16'd2630, 16'd2966, 16'd1584, 16'd30126, 16'd60733, 16'd45813, 16'd42919, 16'd43408, 16'd875, 16'd5939, 16'd64730, 16'd43672, 16'd27855, 16'd35888, 16'd60983, 16'd47648});
	test_expansion(128'h716683bf81f8823fe53865312ed32d28, {16'd3217, 16'd18210, 16'd58577, 16'd50510, 16'd59622, 16'd41070, 16'd25750, 16'd10131, 16'd58436, 16'd9182, 16'd11267, 16'd44914, 16'd35565, 16'd6904, 16'd23506, 16'd49420, 16'd9762, 16'd23591, 16'd60715, 16'd23523, 16'd40817, 16'd39732, 16'd63225, 16'd58809, 16'd18226, 16'd41279});
	test_expansion(128'h02b357c84a85f6ed8f55528a196d7359, {16'd15416, 16'd16929, 16'd1345, 16'd61198, 16'd17768, 16'd14302, 16'd2975, 16'd51069, 16'd34219, 16'd12860, 16'd18189, 16'd15650, 16'd16344, 16'd56293, 16'd37306, 16'd46536, 16'd65361, 16'd8154, 16'd53218, 16'd54134, 16'd62464, 16'd11349, 16'd60453, 16'd51360, 16'd45182, 16'd19808});
	test_expansion(128'h9bd040c932c8ab16576c5dba3d33d723, {16'd52588, 16'd29105, 16'd55623, 16'd31088, 16'd4402, 16'd64289, 16'd7291, 16'd27294, 16'd63572, 16'd21893, 16'd21196, 16'd46042, 16'd17957, 16'd41778, 16'd3239, 16'd21263, 16'd64454, 16'd12792, 16'd59890, 16'd3257, 16'd57412, 16'd56928, 16'd55474, 16'd17247, 16'd6043, 16'd54488});
	test_expansion(128'hd971b44fdc0d8f6e10f9e59f0b028a39, {16'd39115, 16'd15280, 16'd59698, 16'd45738, 16'd34047, 16'd5532, 16'd3807, 16'd45020, 16'd41390, 16'd50906, 16'd47776, 16'd40606, 16'd25214, 16'd2924, 16'd17695, 16'd28637, 16'd41722, 16'd10153, 16'd41904, 16'd3669, 16'd41050, 16'd64149, 16'd55260, 16'd40289, 16'd16862, 16'd13566});
	test_expansion(128'hb38ca098fc5614a838641529875f7cfe, {16'd38922, 16'd61113, 16'd30981, 16'd10116, 16'd51283, 16'd39210, 16'd61988, 16'd57959, 16'd38947, 16'd8986, 16'd42503, 16'd4906, 16'd9381, 16'd1994, 16'd30882, 16'd18172, 16'd349, 16'd16753, 16'd40585, 16'd11814, 16'd7608, 16'd19989, 16'd35953, 16'd46297, 16'd6185, 16'd62935});
	test_expansion(128'hc705665d0d97e14c91780ff3e1009224, {16'd56958, 16'd35640, 16'd30103, 16'd47598, 16'd35762, 16'd20908, 16'd30739, 16'd38894, 16'd55184, 16'd27124, 16'd27412, 16'd59272, 16'd51443, 16'd45039, 16'd55672, 16'd65118, 16'd53655, 16'd22709, 16'd399, 16'd8706, 16'd24043, 16'd65112, 16'd12471, 16'd33481, 16'd55337, 16'd50466});
	test_expansion(128'h33a9e6b84a57bb9ff59ecc142f3e69fc, {16'd12616, 16'd19275, 16'd41176, 16'd4583, 16'd62217, 16'd37725, 16'd57001, 16'd27793, 16'd32039, 16'd38251, 16'd64925, 16'd44247, 16'd3290, 16'd64448, 16'd58361, 16'd54348, 16'd25819, 16'd40949, 16'd15959, 16'd51166, 16'd52295, 16'd2386, 16'd64779, 16'd50389, 16'd42682, 16'd29332});
	test_expansion(128'h1c202df97ed3c70140da81f288036207, {16'd54017, 16'd55278, 16'd11558, 16'd45582, 16'd53923, 16'd30296, 16'd38760, 16'd46770, 16'd37100, 16'd56644, 16'd532, 16'd29150, 16'd8577, 16'd12796, 16'd30965, 16'd2365, 16'd38489, 16'd56004, 16'd32521, 16'd3615, 16'd20021, 16'd42891, 16'd3097, 16'd20105, 16'd12773, 16'd8591});
	test_expansion(128'h618d7a786952e6507fe1be6fb23d154f, {16'd59585, 16'd4735, 16'd20171, 16'd39562, 16'd10616, 16'd62318, 16'd28899, 16'd26206, 16'd32974, 16'd36716, 16'd26712, 16'd38639, 16'd28156, 16'd26463, 16'd49318, 16'd2298, 16'd616, 16'd47538, 16'd31230, 16'd23491, 16'd38276, 16'd47232, 16'd30408, 16'd47904, 16'd25859, 16'd55423});
	test_expansion(128'h5eedb4a6bebb8d9f36dbdc358f9e4dfe, {16'd13644, 16'd16927, 16'd23895, 16'd10067, 16'd55813, 16'd64456, 16'd10773, 16'd38521, 16'd56290, 16'd25245, 16'd48469, 16'd44987, 16'd23879, 16'd7097, 16'd57607, 16'd6361, 16'd22061, 16'd57250, 16'd56032, 16'd34945, 16'd25495, 16'd1002, 16'd271, 16'd62229, 16'd25244, 16'd27582});
	test_expansion(128'h2877655d906ac52932ea322c249c3bb2, {16'd27612, 16'd4741, 16'd29114, 16'd38367, 16'd45918, 16'd47978, 16'd13887, 16'd35696, 16'd14642, 16'd33044, 16'd54010, 16'd52417, 16'd19212, 16'd53074, 16'd51942, 16'd45415, 16'd8603, 16'd14447, 16'd218, 16'd5989, 16'd10306, 16'd6254, 16'd7323, 16'd5807, 16'd12051, 16'd39903});
	test_expansion(128'h081288319eaf595f6170548077acc0cb, {16'd60914, 16'd37888, 16'd48358, 16'd57125, 16'd60010, 16'd50289, 16'd45225, 16'd14884, 16'd45642, 16'd57732, 16'd30567, 16'd39634, 16'd11882, 16'd12062, 16'd27437, 16'd63730, 16'd53952, 16'd16150, 16'd15747, 16'd2361, 16'd40302, 16'd35134, 16'd14561, 16'd51972, 16'd31269, 16'd26485});
	test_expansion(128'h4980aac02043877348dda51ba05625f5, {16'd55835, 16'd14969, 16'd46556, 16'd21983, 16'd29222, 16'd35277, 16'd4466, 16'd57040, 16'd19646, 16'd42952, 16'd50016, 16'd6230, 16'd32838, 16'd5193, 16'd56787, 16'd56113, 16'd40937, 16'd6565, 16'd61469, 16'd60898, 16'd25883, 16'd55589, 16'd1287, 16'd36440, 16'd18082, 16'd35820});
	test_expansion(128'h88ec34c7216386b3675044c91dd52cbd, {16'd55453, 16'd13825, 16'd11541, 16'd28230, 16'd37110, 16'd47157, 16'd21058, 16'd53839, 16'd12869, 16'd33951, 16'd39110, 16'd7470, 16'd367, 16'd21161, 16'd32399, 16'd33642, 16'd3325, 16'd53387, 16'd4994, 16'd2851, 16'd1876, 16'd21820, 16'd33183, 16'd61473, 16'd39093, 16'd2755});
	test_expansion(128'h00f32b0c8e0b57f9fb0ffea09d633d50, {16'd26910, 16'd61329, 16'd8463, 16'd35800, 16'd46888, 16'd26986, 16'd50869, 16'd43786, 16'd64962, 16'd26421, 16'd57133, 16'd12367, 16'd9560, 16'd48214, 16'd60686, 16'd21793, 16'd28077, 16'd6713, 16'd56175, 16'd48611, 16'd30498, 16'd48180, 16'd54723, 16'd60814, 16'd37504, 16'd16533});
	test_expansion(128'h9ac558a6ff3b652b99b333c5654cc0e4, {16'd7790, 16'd53521, 16'd26863, 16'd58382, 16'd28490, 16'd39477, 16'd38074, 16'd31344, 16'd56528, 16'd55617, 16'd60815, 16'd5313, 16'd57864, 16'd20578, 16'd57489, 16'd48716, 16'd62922, 16'd47586, 16'd53808, 16'd38582, 16'd62804, 16'd4366, 16'd42302, 16'd46876, 16'd120, 16'd57499});
	test_expansion(128'he47e22baee41e1b2e6160238cd3105e6, {16'd32579, 16'd1265, 16'd20788, 16'd18655, 16'd41013, 16'd35203, 16'd31618, 16'd4539, 16'd24264, 16'd58944, 16'd42840, 16'd56167, 16'd48597, 16'd25417, 16'd64231, 16'd23362, 16'd35426, 16'd35933, 16'd56548, 16'd447, 16'd59745, 16'd13160, 16'd56753, 16'd15028, 16'd15779, 16'd16085});
	test_expansion(128'h72ebc0ee9f9929ab37108e9865666157, {16'd36786, 16'd36045, 16'd35830, 16'd14300, 16'd27391, 16'd37840, 16'd38491, 16'd23403, 16'd56119, 16'd8769, 16'd47893, 16'd6047, 16'd35189, 16'd61306, 16'd4587, 16'd36075, 16'd10806, 16'd38043, 16'd11955, 16'd54619, 16'd64951, 16'd51462, 16'd22265, 16'd34957, 16'd59826, 16'd61839});
	test_expansion(128'hdb2003fc0d8ad240770f41543c0fffe2, {16'd21622, 16'd33177, 16'd31120, 16'd12619, 16'd7359, 16'd26615, 16'd1935, 16'd30718, 16'd51394, 16'd58295, 16'd5727, 16'd32803, 16'd11710, 16'd13364, 16'd11994, 16'd6872, 16'd16434, 16'd25850, 16'd153, 16'd34660, 16'd41851, 16'd58829, 16'd35796, 16'd641, 16'd2915, 16'd31784});
	test_expansion(128'he6103b4deac7d3452f93c79340bde3b7, {16'd32432, 16'd25167, 16'd60877, 16'd47850, 16'd61028, 16'd56430, 16'd34971, 16'd48134, 16'd63061, 16'd4083, 16'd58003, 16'd36560, 16'd22995, 16'd63508, 16'd37706, 16'd57498, 16'd9767, 16'd17342, 16'd20061, 16'd43937, 16'd30649, 16'd64427, 16'd57631, 16'd19151, 16'd12668, 16'd29857});
	test_expansion(128'he9aab5b0899e43b9257eae0259c7ff9d, {16'd50224, 16'd18313, 16'd41864, 16'd79, 16'd14240, 16'd42353, 16'd36031, 16'd30593, 16'd18964, 16'd24435, 16'd3540, 16'd27816, 16'd62882, 16'd28060, 16'd2161, 16'd19795, 16'd45779, 16'd52055, 16'd38882, 16'd54730, 16'd15425, 16'd38470, 16'd33894, 16'd49459, 16'd22914, 16'd54833});
	test_expansion(128'h2008dd645d2a89537b3d5483a8f5e32b, {16'd25018, 16'd49422, 16'd65096, 16'd56619, 16'd10992, 16'd32778, 16'd40360, 16'd1867, 16'd52723, 16'd34319, 16'd36724, 16'd28179, 16'd42385, 16'd34278, 16'd50324, 16'd58885, 16'd37225, 16'd14970, 16'd30473, 16'd5148, 16'd44162, 16'd63769, 16'd49973, 16'd13285, 16'd38885, 16'd12598});
	test_expansion(128'h19c2a5c017d030c9ecee82dd227615e7, {16'd63518, 16'd17252, 16'd36298, 16'd1197, 16'd50782, 16'd32630, 16'd64797, 16'd16905, 16'd42846, 16'd61296, 16'd2295, 16'd44269, 16'd43320, 16'd41681, 16'd3101, 16'd24333, 16'd45716, 16'd386, 16'd49125, 16'd11531, 16'd42321, 16'd39036, 16'd40836, 16'd2652, 16'd48323, 16'd955});
	test_expansion(128'hb9b33c14144846cf00e0eedf59ea82f4, {16'd59684, 16'd52810, 16'd55297, 16'd62950, 16'd30527, 16'd6810, 16'd58854, 16'd50061, 16'd50492, 16'd19314, 16'd47765, 16'd26040, 16'd8884, 16'd47920, 16'd50138, 16'd51266, 16'd62566, 16'd3188, 16'd25979, 16'd43664, 16'd42838, 16'd28906, 16'd17390, 16'd50131, 16'd64570, 16'd2144});
	test_expansion(128'hf6a875122cb177044a864374c281f2a6, {16'd19577, 16'd45964, 16'd10161, 16'd43818, 16'd33579, 16'd61956, 16'd45455, 16'd59697, 16'd55851, 16'd10017, 16'd23327, 16'd3711, 16'd45874, 16'd4484, 16'd17077, 16'd43377, 16'd43259, 16'd29808, 16'd63322, 16'd46000, 16'd31665, 16'd63977, 16'd19250, 16'd31396, 16'd15502, 16'd40156});
	test_expansion(128'hbfdaebd82cadebefcd73a49b3ae64b45, {16'd39459, 16'd23664, 16'd5304, 16'd15216, 16'd25700, 16'd27073, 16'd18076, 16'd51129, 16'd34626, 16'd17023, 16'd495, 16'd39702, 16'd54680, 16'd10445, 16'd49427, 16'd9519, 16'd57744, 16'd19468, 16'd45305, 16'd43380, 16'd43638, 16'd2534, 16'd21240, 16'd51867, 16'd50464, 16'd65291});
	test_expansion(128'hca6f3ab45ea463337485c1a70bdcd2fd, {16'd30218, 16'd29115, 16'd49629, 16'd43728, 16'd57149, 16'd33702, 16'd9583, 16'd322, 16'd39634, 16'd31534, 16'd31128, 16'd13188, 16'd42032, 16'd61628, 16'd1657, 16'd1799, 16'd35848, 16'd44022, 16'd53514, 16'd55307, 16'd599, 16'd19125, 16'd27988, 16'd58785, 16'd49141, 16'd46858});
	test_expansion(128'h5bcc458f8e50b2f46093e4bac4669a17, {16'd37862, 16'd22309, 16'd53, 16'd29624, 16'd48077, 16'd1043, 16'd28400, 16'd7096, 16'd30537, 16'd8118, 16'd22913, 16'd38327, 16'd49191, 16'd30470, 16'd51056, 16'd7449, 16'd61090, 16'd2775, 16'd35568, 16'd53057, 16'd33247, 16'd64756, 16'd10337, 16'd50536, 16'd23931, 16'd34276});
	test_expansion(128'h44430ad45f413449b7267179a69093c9, {16'd45468, 16'd62376, 16'd60908, 16'd19647, 16'd11466, 16'd41157, 16'd53673, 16'd10909, 16'd9617, 16'd16998, 16'd7868, 16'd1058, 16'd15105, 16'd55752, 16'd54693, 16'd35120, 16'd10251, 16'd13188, 16'd37381, 16'd9852, 16'd46308, 16'd8932, 16'd10960, 16'd8391, 16'd5219, 16'd55561});
	test_expansion(128'h15a8c4b0b415613936158d7bb330be6a, {16'd20318, 16'd54476, 16'd13232, 16'd59746, 16'd53340, 16'd11913, 16'd11554, 16'd55057, 16'd4902, 16'd20985, 16'd62677, 16'd37667, 16'd40868, 16'd63934, 16'd45751, 16'd54465, 16'd44401, 16'd27381, 16'd41355, 16'd38968, 16'd41686, 16'd25253, 16'd27215, 16'd47596, 16'd13254, 16'd49478});
	test_expansion(128'he599e33faf3a0e6d0141caee3006cb2a, {16'd53842, 16'd4318, 16'd21357, 16'd47596, 16'd14412, 16'd52922, 16'd7930, 16'd25757, 16'd43614, 16'd24618, 16'd40850, 16'd10527, 16'd34430, 16'd57879, 16'd35057, 16'd9592, 16'd8308, 16'd47930, 16'd26983, 16'd54137, 16'd37535, 16'd63263, 16'd53963, 16'd23755, 16'd30145, 16'd47832});
	test_expansion(128'h43fd35870d7446ebe76b93112c4963ce, {16'd46552, 16'd4659, 16'd53712, 16'd55000, 16'd22043, 16'd53649, 16'd13663, 16'd14836, 16'd64394, 16'd24325, 16'd9864, 16'd105, 16'd13747, 16'd1005, 16'd63397, 16'd12034, 16'd14809, 16'd14983, 16'd63196, 16'd7833, 16'd42889, 16'd48678, 16'd45681, 16'd46735, 16'd31210, 16'd6366});
	test_expansion(128'h1c6e6c52c23c8cae960eddf7e7078db1, {16'd26311, 16'd12983, 16'd14163, 16'd917, 16'd39076, 16'd36942, 16'd24293, 16'd2313, 16'd1303, 16'd9802, 16'd44901, 16'd52618, 16'd11394, 16'd57838, 16'd34595, 16'd53273, 16'd3977, 16'd31430, 16'd44742, 16'd57897, 16'd15957, 16'd27970, 16'd38518, 16'd48712, 16'd29957, 16'd42312});
	test_expansion(128'h70eca0e1b7e3f867d5fc5d0b60b7e6bd, {16'd19960, 16'd33590, 16'd8989, 16'd48317, 16'd56740, 16'd27541, 16'd7639, 16'd44414, 16'd34375, 16'd58635, 16'd59184, 16'd19037, 16'd7595, 16'd7188, 16'd44332, 16'd52729, 16'd32905, 16'd27924, 16'd5381, 16'd53930, 16'd8699, 16'd47078, 16'd8611, 16'd44285, 16'd22351, 16'd34298});
	test_expansion(128'h3df9679ffc0436b4b0f603a9bf240163, {16'd40, 16'd37280, 16'd6634, 16'd32547, 16'd39428, 16'd7472, 16'd59034, 16'd13705, 16'd21478, 16'd6904, 16'd12032, 16'd41159, 16'd11786, 16'd59859, 16'd59411, 16'd19660, 16'd48642, 16'd29916, 16'd24268, 16'd55154, 16'd56019, 16'd3905, 16'd59111, 16'd20526, 16'd3611, 16'd11787});
	test_expansion(128'hbfac4c5a27dea2297f67056bf4e30c5b, {16'd48173, 16'd47780, 16'd54876, 16'd37337, 16'd5078, 16'd2757, 16'd57431, 16'd15831, 16'd14876, 16'd6296, 16'd3860, 16'd33700, 16'd40196, 16'd40853, 16'd47502, 16'd41298, 16'd64725, 16'd36941, 16'd28007, 16'd56374, 16'd2282, 16'd10795, 16'd43934, 16'd43036, 16'd26462, 16'd12712});
	test_expansion(128'hbbb2862652f299a13de5208b1776dfe5, {16'd34820, 16'd27345, 16'd43406, 16'd57096, 16'd8711, 16'd41319, 16'd13992, 16'd57709, 16'd56685, 16'd56667, 16'd47757, 16'd19355, 16'd39235, 16'd4291, 16'd51429, 16'd45101, 16'd19616, 16'd42087, 16'd46615, 16'd41672, 16'd4350, 16'd10240, 16'd24924, 16'd21937, 16'd14981, 16'd56936});
	test_expansion(128'h0b19554458872b2a80e7b153503b2a19, {16'd29269, 16'd19035, 16'd45447, 16'd58023, 16'd65087, 16'd52214, 16'd11958, 16'd59063, 16'd36227, 16'd4053, 16'd923, 16'd36084, 16'd7450, 16'd15628, 16'd28362, 16'd12988, 16'd10000, 16'd52211, 16'd31782, 16'd58010, 16'd15225, 16'd13817, 16'd17028, 16'd43342, 16'd38033, 16'd16685});
	test_expansion(128'h42d6cca7480bc1ef1af37e416a17d3eb, {16'd37856, 16'd32717, 16'd44909, 16'd51136, 16'd24870, 16'd5677, 16'd32845, 16'd9836, 16'd28345, 16'd16581, 16'd43837, 16'd38438, 16'd26694, 16'd53234, 16'd6238, 16'd9098, 16'd34578, 16'd2163, 16'd48542, 16'd15060, 16'd58062, 16'd31187, 16'd12030, 16'd64032, 16'd40323, 16'd37023});
	test_expansion(128'h17460906b29335910a91ffa325468265, {16'd182, 16'd34979, 16'd45587, 16'd60516, 16'd16006, 16'd57532, 16'd54560, 16'd39532, 16'd34785, 16'd32683, 16'd12985, 16'd64473, 16'd24474, 16'd1621, 16'd9504, 16'd4309, 16'd28024, 16'd3948, 16'd35894, 16'd56953, 16'd52247, 16'd36171, 16'd5907, 16'd50759, 16'd3231, 16'd42863});
	test_expansion(128'h5254fe5f08add42d47e88fefd25d52c9, {16'd25730, 16'd64348, 16'd47486, 16'd39908, 16'd22339, 16'd63990, 16'd56931, 16'd36762, 16'd24357, 16'd14592, 16'd63551, 16'd59869, 16'd14565, 16'd3174, 16'd58788, 16'd27339, 16'd28664, 16'd47777, 16'd49247, 16'd64795, 16'd49372, 16'd58592, 16'd52508, 16'd40190, 16'd34261, 16'd33075});
	test_expansion(128'h4a5d7b1f8a34a527a8dc79b1126f768f, {16'd63628, 16'd53972, 16'd4250, 16'd14728, 16'd61407, 16'd61567, 16'd58526, 16'd13162, 16'd21688, 16'd19132, 16'd41020, 16'd19421, 16'd31296, 16'd4406, 16'd55924, 16'd53592, 16'd11514, 16'd34686, 16'd39680, 16'd49281, 16'd62104, 16'd55659, 16'd20141, 16'd56660, 16'd18840, 16'd59761});
	test_expansion(128'hb39a2ddb00865ce10713f6115bc3471b, {16'd53343, 16'd57292, 16'd1116, 16'd2697, 16'd28837, 16'd12644, 16'd18601, 16'd55085, 16'd28568, 16'd11814, 16'd11196, 16'd64916, 16'd26949, 16'd14199, 16'd34581, 16'd17777, 16'd59925, 16'd1220, 16'd20317, 16'd15479, 16'd17307, 16'd21908, 16'd39330, 16'd36746, 16'd28009, 16'd4739});
	test_expansion(128'h5fd2d092fa9f684a392bbace002e3af7, {16'd50069, 16'd5042, 16'd38328, 16'd53562, 16'd25225, 16'd12533, 16'd36140, 16'd64208, 16'd27980, 16'd51467, 16'd56177, 16'd11622, 16'd36230, 16'd41053, 16'd29614, 16'd22241, 16'd35466, 16'd40716, 16'd36577, 16'd9420, 16'd19540, 16'd31959, 16'd65386, 16'd62693, 16'd54691, 16'd39358});
	test_expansion(128'h636fbb46302a663dfa7100d7b62ca3c5, {16'd10398, 16'd57258, 16'd63208, 16'd20186, 16'd12524, 16'd20179, 16'd32946, 16'd13362, 16'd65021, 16'd64625, 16'd38633, 16'd42618, 16'd13400, 16'd56337, 16'd64097, 16'd26817, 16'd4179, 16'd35202, 16'd59790, 16'd22499, 16'd22482, 16'd46647, 16'd50699, 16'd51251, 16'd12564, 16'd7008});
	test_expansion(128'h988e7a8f214ea24433bfdbcb582a50da, {16'd43381, 16'd4838, 16'd36507, 16'd7106, 16'd15633, 16'd65128, 16'd40699, 16'd64472, 16'd2626, 16'd1601, 16'd4898, 16'd12787, 16'd34853, 16'd10073, 16'd46034, 16'd36234, 16'd136, 16'd59011, 16'd61152, 16'd13065, 16'd11192, 16'd42759, 16'd28225, 16'd4466, 16'd61107, 16'd148});
	test_expansion(128'hf5f48c5209cf2891abebe854c362cb7c, {16'd40599, 16'd51718, 16'd37850, 16'd10752, 16'd6027, 16'd62863, 16'd20732, 16'd7636, 16'd44395, 16'd34293, 16'd19218, 16'd59662, 16'd69, 16'd36178, 16'd17104, 16'd16074, 16'd49741, 16'd44259, 16'd41645, 16'd8848, 16'd14726, 16'd56046, 16'd33944, 16'd55808, 16'd55965, 16'd12018});
	test_expansion(128'h04ff8b18e06b7be64a45048d534cb52b, {16'd37259, 16'd3310, 16'd54234, 16'd17055, 16'd58864, 16'd26986, 16'd22723, 16'd44556, 16'd50342, 16'd56906, 16'd59658, 16'd50975, 16'd25377, 16'd51459, 16'd1374, 16'd41819, 16'd19422, 16'd31988, 16'd9816, 16'd2002, 16'd1946, 16'd41305, 16'd59595, 16'd11571, 16'd33829, 16'd43236});
	test_expansion(128'h65d4886a0c99d31adaee64356e3e264a, {16'd5024, 16'd18236, 16'd36467, 16'd44033, 16'd58978, 16'd61867, 16'd14913, 16'd28829, 16'd48744, 16'd53386, 16'd28796, 16'd46892, 16'd44299, 16'd53713, 16'd44537, 16'd22946, 16'd45646, 16'd49215, 16'd65319, 16'd1484, 16'd8464, 16'd5880, 16'd57486, 16'd41940, 16'd21994, 16'd20925});
	test_expansion(128'h4ca866e3099552711af2a328ade443d7, {16'd40759, 16'd41225, 16'd61431, 16'd48308, 16'd61718, 16'd61386, 16'd41302, 16'd14545, 16'd64845, 16'd37878, 16'd27522, 16'd11381, 16'd21538, 16'd19464, 16'd51969, 16'd8564, 16'd21450, 16'd19555, 16'd41528, 16'd14635, 16'd42163, 16'd41022, 16'd59923, 16'd832, 16'd34517, 16'd42338});
	test_expansion(128'h418ee831410711f79b555116cc65dfb7, {16'd23569, 16'd62448, 16'd51723, 16'd18491, 16'd62692, 16'd33494, 16'd26480, 16'd41309, 16'd58923, 16'd2834, 16'd50094, 16'd17921, 16'd15037, 16'd37594, 16'd39781, 16'd59234, 16'd62297, 16'd49209, 16'd60959, 16'd27155, 16'd25808, 16'd42352, 16'd26653, 16'd50259, 16'd40846, 16'd51723});
	test_expansion(128'h72c6a99bed25cbda7cb3346ed417ddbd, {16'd8951, 16'd39464, 16'd59126, 16'd54629, 16'd17037, 16'd58971, 16'd59471, 16'd36604, 16'd45190, 16'd45542, 16'd8916, 16'd17909, 16'd28147, 16'd32934, 16'd31668, 16'd40698, 16'd86, 16'd20827, 16'd975, 16'd64404, 16'd4925, 16'd58511, 16'd49956, 16'd8150, 16'd11793, 16'd59226});
	test_expansion(128'hf7c60338affc2ff6b9c1a3790fe4ef36, {16'd16529, 16'd2026, 16'd27428, 16'd2186, 16'd43877, 16'd1410, 16'd60948, 16'd17288, 16'd12127, 16'd28664, 16'd11773, 16'd29491, 16'd37081, 16'd12021, 16'd23267, 16'd3626, 16'd19476, 16'd54344, 16'd32523, 16'd13636, 16'd11628, 16'd64400, 16'd52666, 16'd26303, 16'd26091, 16'd29903});
	test_expansion(128'hfa791bbd5653ead4189490d80679181d, {16'd56391, 16'd55499, 16'd28354, 16'd54092, 16'd418, 16'd55573, 16'd39321, 16'd56545, 16'd3745, 16'd6708, 16'd37920, 16'd54012, 16'd34837, 16'd40218, 16'd46672, 16'd8973, 16'd11218, 16'd29142, 16'd37405, 16'd4730, 16'd50994, 16'd45614, 16'd16393, 16'd34827, 16'd23309, 16'd53445});
	test_expansion(128'hcaad24022765fed924abef34f1451b31, {16'd23560, 16'd2245, 16'd20040, 16'd2005, 16'd38202, 16'd6366, 16'd17339, 16'd19714, 16'd54788, 16'd65309, 16'd53636, 16'd44347, 16'd17247, 16'd29437, 16'd15636, 16'd37823, 16'd17336, 16'd2386, 16'd14642, 16'd55138, 16'd56082, 16'd21383, 16'd30777, 16'd14119, 16'd42618, 16'd43449});
	test_expansion(128'hb85f30528a417914c7bcbcbe2869f4c5, {16'd21527, 16'd48050, 16'd28833, 16'd59883, 16'd60044, 16'd59113, 16'd39696, 16'd44499, 16'd51868, 16'd47571, 16'd60373, 16'd40654, 16'd30307, 16'd23154, 16'd22457, 16'd51409, 16'd26628, 16'd58771, 16'd53165, 16'd6918, 16'd47299, 16'd9155, 16'd31224, 16'd4565, 16'd59912, 16'd49184});
	test_expansion(128'h8c92075ff3c61b5c4a3d38dd8f044dbc, {16'd15783, 16'd15507, 16'd45169, 16'd53187, 16'd54256, 16'd41512, 16'd51486, 16'd31131, 16'd2036, 16'd15553, 16'd10339, 16'd63725, 16'd48248, 16'd49067, 16'd58827, 16'd15303, 16'd286, 16'd47462, 16'd15181, 16'd43611, 16'd15994, 16'd47385, 16'd24788, 16'd29735, 16'd18756, 16'd195});
	test_expansion(128'h5d116011ea4dbd4ea99db06745057a8d, {16'd33519, 16'd19683, 16'd28622, 16'd36340, 16'd45517, 16'd25685, 16'd51666, 16'd7846, 16'd681, 16'd59657, 16'd3797, 16'd40452, 16'd54576, 16'd17675, 16'd15569, 16'd51071, 16'd8077, 16'd46837, 16'd11275, 16'd62944, 16'd50805, 16'd51685, 16'd21582, 16'd13056, 16'd30014, 16'd11745});
	test_expansion(128'h1ab14e2aa8074489b596f78afd2eb04f, {16'd44846, 16'd16328, 16'd155, 16'd22946, 16'd36989, 16'd40109, 16'd24442, 16'd52091, 16'd21581, 16'd50990, 16'd35352, 16'd56314, 16'd35134, 16'd1795, 16'd28301, 16'd52626, 16'd9568, 16'd58237, 16'd32418, 16'd50355, 16'd57194, 16'd31324, 16'd61372, 16'd12746, 16'd19949, 16'd12029});
	test_expansion(128'h4cfcfc45e4ea6d46acd156df2061331d, {16'd2394, 16'd31842, 16'd63791, 16'd1470, 16'd2176, 16'd47767, 16'd484, 16'd10965, 16'd32525, 16'd43190, 16'd17165, 16'd52448, 16'd48052, 16'd54692, 16'd15828, 16'd8069, 16'd40933, 16'd56516, 16'd33896, 16'd40067, 16'd18886, 16'd30327, 16'd38059, 16'd18646, 16'd17552, 16'd48923});
	test_expansion(128'hb75ed3d4e68c8c2bccec148454a19257, {16'd1204, 16'd35505, 16'd27666, 16'd57917, 16'd47178, 16'd43999, 16'd54085, 16'd39460, 16'd63175, 16'd55712, 16'd6874, 16'd16577, 16'd59470, 16'd4003, 16'd60976, 16'd18579, 16'd19952, 16'd8805, 16'd18948, 16'd56729, 16'd20108, 16'd769, 16'd41840, 16'd32094, 16'd21132, 16'd2559});
	test_expansion(128'h5628e249134ec745bee9748a8fbac1fd, {16'd5231, 16'd61182, 16'd39671, 16'd56526, 16'd1914, 16'd2748, 16'd11071, 16'd28172, 16'd55534, 16'd2678, 16'd42082, 16'd11234, 16'd38691, 16'd40755, 16'd28320, 16'd45592, 16'd35123, 16'd21211, 16'd15438, 16'd50691, 16'd62129, 16'd61105, 16'd55482, 16'd43609, 16'd58906, 16'd57827});
	test_expansion(128'ha13e0d71e3daefcc754d3921292342ac, {16'd63570, 16'd57303, 16'd26958, 16'd14357, 16'd35124, 16'd6115, 16'd56156, 16'd322, 16'd28120, 16'd44335, 16'd1844, 16'd23579, 16'd7863, 16'd16358, 16'd37258, 16'd41050, 16'd25365, 16'd34188, 16'd13872, 16'd11546, 16'd716, 16'd64044, 16'd64453, 16'd31523, 16'd17289, 16'd22452});
	test_expansion(128'h6a5171c96288e44ed56cbd0b77ae87a7, {16'd1885, 16'd54696, 16'd55227, 16'd22197, 16'd19487, 16'd18558, 16'd52686, 16'd27936, 16'd27587, 16'd27195, 16'd42342, 16'd63517, 16'd48341, 16'd12966, 16'd51548, 16'd60633, 16'd30304, 16'd28744, 16'd21786, 16'd29818, 16'd30730, 16'd48760, 16'd15451, 16'd52050, 16'd49094, 16'd26890});
	test_expansion(128'h10b69797312aa0871f648cd0ea651a0f, {16'd12264, 16'd438, 16'd58901, 16'd35543, 16'd11680, 16'd58440, 16'd28287, 16'd25629, 16'd525, 16'd64081, 16'd60052, 16'd16382, 16'd60820, 16'd50554, 16'd10246, 16'd915, 16'd13150, 16'd65247, 16'd41084, 16'd36561, 16'd15881, 16'd41508, 16'd6535, 16'd22728, 16'd31753, 16'd47104});
	test_expansion(128'h51e90947ae824a02a5b910ff7746ca39, {16'd18910, 16'd55867, 16'd15082, 16'd10491, 16'd13846, 16'd47254, 16'd22707, 16'd28663, 16'd8833, 16'd6982, 16'd16762, 16'd26653, 16'd35723, 16'd15661, 16'd60856, 16'd12242, 16'd37932, 16'd58310, 16'd6130, 16'd37741, 16'd25059, 16'd21840, 16'd8664, 16'd18198, 16'd61027, 16'd40201});
	test_expansion(128'ha1d9cdc0319495682a4c30054115f6ea, {16'd8405, 16'd4488, 16'd37007, 16'd5099, 16'd62110, 16'd28617, 16'd37078, 16'd19370, 16'd56402, 16'd55678, 16'd34674, 16'd31527, 16'd9478, 16'd62255, 16'd4047, 16'd15618, 16'd9907, 16'd42136, 16'd41711, 16'd45782, 16'd3623, 16'd13814, 16'd45807, 16'd44857, 16'd11485, 16'd12653});
	test_expansion(128'h005e5bc7fd21b389ae8fe8a1750b058f, {16'd63485, 16'd51998, 16'd39776, 16'd45936, 16'd55889, 16'd51109, 16'd5730, 16'd47586, 16'd5449, 16'd33987, 16'd29345, 16'd17647, 16'd35755, 16'd46244, 16'd37628, 16'd45531, 16'd32435, 16'd34801, 16'd15879, 16'd33145, 16'd31484, 16'd63462, 16'd31082, 16'd10518, 16'd19229, 16'd32384});
	test_expansion(128'h29aac2ca67aad3a59748c4841f31516c, {16'd14982, 16'd24422, 16'd40106, 16'd14019, 16'd5099, 16'd39799, 16'd12351, 16'd35967, 16'd60793, 16'd27065, 16'd10827, 16'd52086, 16'd2896, 16'd44708, 16'd11121, 16'd30196, 16'd1075, 16'd55475, 16'd13863, 16'd29486, 16'd55426, 16'd21823, 16'd44064, 16'd50667, 16'd61344, 16'd11477});
	test_expansion(128'he92e188f8a983b38a176e09fab42ac43, {16'd23184, 16'd34993, 16'd64726, 16'd23723, 16'd26267, 16'd11447, 16'd37718, 16'd13472, 16'd33152, 16'd40467, 16'd40177, 16'd41274, 16'd30288, 16'd21344, 16'd63915, 16'd53633, 16'd43506, 16'd23299, 16'd55663, 16'd13140, 16'd35423, 16'd27589, 16'd53890, 16'd12440, 16'd62681, 16'd28626});
	test_expansion(128'hdbf30fe20507641485dc4d633c9ccc09, {16'd42584, 16'd44167, 16'd31565, 16'd50348, 16'd24745, 16'd48131, 16'd12488, 16'd63688, 16'd51925, 16'd63349, 16'd32102, 16'd30695, 16'd37454, 16'd10920, 16'd55392, 16'd46133, 16'd46371, 16'd45426, 16'd64059, 16'd5472, 16'd32932, 16'd15027, 16'd14599, 16'd34933, 16'd60432, 16'd7113});
	test_expansion(128'hc72f1bbec9a867b422daddc3f282b629, {16'd16818, 16'd23149, 16'd40015, 16'd43743, 16'd57053, 16'd4834, 16'd36184, 16'd58326, 16'd33655, 16'd41160, 16'd49982, 16'd44284, 16'd52149, 16'd31799, 16'd61719, 16'd54127, 16'd52933, 16'd2098, 16'd49854, 16'd26958, 16'd36606, 16'd17993, 16'd40068, 16'd53259, 16'd61451, 16'd1836});
	test_expansion(128'h30439c23c82b3cd21ee815ca251cfc58, {16'd38785, 16'd33700, 16'd25402, 16'd49430, 16'd1980, 16'd10244, 16'd55665, 16'd17603, 16'd52977, 16'd44175, 16'd21639, 16'd25629, 16'd44126, 16'd3970, 16'd55264, 16'd8472, 16'd45533, 16'd62297, 16'd31718, 16'd62821, 16'd57392, 16'd51066, 16'd24633, 16'd32415, 16'd54391, 16'd37920});
	test_expansion(128'h36dd8ec7d3734fa1e27cca6b9a8070ba, {16'd49970, 16'd21625, 16'd55466, 16'd47092, 16'd47396, 16'd48696, 16'd16516, 16'd49498, 16'd47967, 16'd20342, 16'd48387, 16'd10945, 16'd41178, 16'd58015, 16'd62592, 16'd3934, 16'd16626, 16'd59913, 16'd56174, 16'd29200, 16'd57553, 16'd16371, 16'd16734, 16'd25707, 16'd27327, 16'd56818});
	test_expansion(128'h0645c8325fd0efe2ca677a35a26127de, {16'd42178, 16'd57488, 16'd57191, 16'd36602, 16'd37475, 16'd24159, 16'd46416, 16'd25653, 16'd27761, 16'd25308, 16'd9137, 16'd12575, 16'd2668, 16'd44143, 16'd23209, 16'd57348, 16'd57651, 16'd220, 16'd60074, 16'd5960, 16'd64149, 16'd9110, 16'd55797, 16'd27626, 16'd21744, 16'd10033});
	test_expansion(128'h7f9288f7ae9639f54d396ae565bd3d3d, {16'd47704, 16'd41541, 16'd42935, 16'd23193, 16'd3392, 16'd38816, 16'd57632, 16'd5677, 16'd53146, 16'd40038, 16'd63493, 16'd21372, 16'd10109, 16'd41017, 16'd34098, 16'd24761, 16'd36556, 16'd23160, 16'd6464, 16'd31241, 16'd12305, 16'd16787, 16'd39076, 16'd49417, 16'd8671, 16'd49709});
	test_expansion(128'h607d588d9f2e63a3c4b74a63126dbaac, {16'd55764, 16'd33701, 16'd56138, 16'd3056, 16'd2318, 16'd12509, 16'd6530, 16'd10866, 16'd47665, 16'd50866, 16'd63342, 16'd54286, 16'd45712, 16'd4555, 16'd59786, 16'd55006, 16'd41629, 16'd32368, 16'd5385, 16'd42001, 16'd23792, 16'd42152, 16'd42984, 16'd42077, 16'd27786, 16'd32981});
	test_expansion(128'h7d2d39333e30ecbeb4fb60c0ca36daab, {16'd34931, 16'd57710, 16'd38005, 16'd62059, 16'd54267, 16'd3274, 16'd47043, 16'd29552, 16'd37142, 16'd47266, 16'd42399, 16'd46772, 16'd47647, 16'd37762, 16'd56920, 16'd58328, 16'd46342, 16'd26772, 16'd25918, 16'd24118, 16'd33217, 16'd52109, 16'd56107, 16'd19136, 16'd16455, 16'd47962});
	test_expansion(128'hdc956f1be6d0289e3000a823da93465e, {16'd52444, 16'd8418, 16'd6558, 16'd52625, 16'd8101, 16'd1869, 16'd46773, 16'd10729, 16'd57260, 16'd53262, 16'd12381, 16'd64889, 16'd26273, 16'd19410, 16'd11191, 16'd12364, 16'd713, 16'd8436, 16'd24944, 16'd38525, 16'd58473, 16'd48372, 16'd46571, 16'd15459, 16'd1717, 16'd21399});
	test_expansion(128'hc2dbf00b57f9d1c7de33486109d827db, {16'd16699, 16'd20304, 16'd43977, 16'd52042, 16'd32768, 16'd51619, 16'd29072, 16'd27461, 16'd9726, 16'd19154, 16'd47355, 16'd47973, 16'd5163, 16'd28786, 16'd31363, 16'd49661, 16'd62805, 16'd27264, 16'd9987, 16'd51509, 16'd4354, 16'd41990, 16'd27172, 16'd9514, 16'd60806, 16'd20046});
	test_expansion(128'h11aedb720df6af00cd4d0309f9d07289, {16'd35208, 16'd30060, 16'd2853, 16'd46473, 16'd30468, 16'd36344, 16'd11146, 16'd22994, 16'd63838, 16'd33772, 16'd5170, 16'd40214, 16'd16291, 16'd24614, 16'd4319, 16'd23005, 16'd50829, 16'd39729, 16'd39746, 16'd16764, 16'd47392, 16'd52999, 16'd52092, 16'd14431, 16'd35390, 16'd43326});
	test_expansion(128'hc5298c5197f148304d4d401c000ea7f7, {16'd35609, 16'd36978, 16'd14346, 16'd62964, 16'd3781, 16'd52851, 16'd14275, 16'd13958, 16'd1712, 16'd50683, 16'd12886, 16'd12455, 16'd62314, 16'd38651, 16'd55834, 16'd28493, 16'd44051, 16'd35403, 16'd30044, 16'd54950, 16'd41948, 16'd24851, 16'd44148, 16'd38489, 16'd21128, 16'd9215});
	test_expansion(128'h830df0391ce3d6d195aac307e95e7a46, {16'd32891, 16'd31778, 16'd58066, 16'd19299, 16'd40910, 16'd22142, 16'd11580, 16'd6901, 16'd65203, 16'd28675, 16'd44637, 16'd28009, 16'd58502, 16'd10379, 16'd38007, 16'd60496, 16'd48533, 16'd43173, 16'd24568, 16'd23469, 16'd40632, 16'd25935, 16'd9136, 16'd31793, 16'd25354, 16'd404});
	test_expansion(128'ha2e6e62e6bcf4f4add6b06e935dd3135, {16'd37078, 16'd13374, 16'd27442, 16'd60138, 16'd43619, 16'd47706, 16'd10337, 16'd14478, 16'd15463, 16'd8437, 16'd57513, 16'd54558, 16'd46428, 16'd14293, 16'd31928, 16'd50307, 16'd26151, 16'd20692, 16'd59499, 16'd47064, 16'd62744, 16'd50531, 16'd5059, 16'd1058, 16'd34075, 16'd22232});
	test_expansion(128'h184b4263fe0c592edc25a42f66f59648, {16'd64010, 16'd40697, 16'd54926, 16'd35622, 16'd11858, 16'd11965, 16'd5269, 16'd28432, 16'd36797, 16'd19171, 16'd26455, 16'd65348, 16'd38446, 16'd58816, 16'd18982, 16'd16749, 16'd1238, 16'd46873, 16'd65181, 16'd38270, 16'd26079, 16'd58225, 16'd6042, 16'd55986, 16'd55794, 16'd29721});
	test_expansion(128'h186c83b2e074ea77ce6e53caa937b668, {16'd59244, 16'd51600, 16'd52943, 16'd34884, 16'd28558, 16'd64101, 16'd60345, 16'd56428, 16'd15726, 16'd1988, 16'd30243, 16'd31131, 16'd46753, 16'd60491, 16'd56622, 16'd63782, 16'd20719, 16'd55867, 16'd59230, 16'd61522, 16'd37551, 16'd14315, 16'd25884, 16'd55079, 16'd59532, 16'd34886});
	test_expansion(128'hde2afa66b1851b0834de342c0921eb56, {16'd65480, 16'd33070, 16'd3261, 16'd12247, 16'd14038, 16'd34553, 16'd48445, 16'd47800, 16'd62504, 16'd6879, 16'd1204, 16'd11577, 16'd57361, 16'd17057, 16'd64177, 16'd3648, 16'd7097, 16'd36729, 16'd36855, 16'd57308, 16'd41267, 16'd55052, 16'd40749, 16'd8450, 16'd1707, 16'd49475});
	test_expansion(128'he8c670b2a45b5ed3839cfc5a8b20379b, {16'd27435, 16'd49157, 16'd445, 16'd28388, 16'd16315, 16'd62644, 16'd41805, 16'd19607, 16'd43212, 16'd4549, 16'd32896, 16'd58201, 16'd46710, 16'd5937, 16'd60034, 16'd54835, 16'd11888, 16'd47695, 16'd42221, 16'd56707, 16'd59271, 16'd42698, 16'd17333, 16'd55116, 16'd63015, 16'd12736});
	test_expansion(128'h1159ffe5c1dbf136d4d4103074a6c633, {16'd62397, 16'd55002, 16'd60586, 16'd63157, 16'd2824, 16'd52901, 16'd19818, 16'd13366, 16'd10062, 16'd749, 16'd10014, 16'd64641, 16'd50120, 16'd1628, 16'd53753, 16'd752, 16'd47475, 16'd64603, 16'd53157, 16'd13652, 16'd54742, 16'd34605, 16'd9446, 16'd54943, 16'd45570, 16'd54859});
	test_expansion(128'h1ccfd4fe3b8d6a2a50109ed6b77001c3, {16'd44748, 16'd60648, 16'd42542, 16'd29856, 16'd64198, 16'd7045, 16'd29258, 16'd35036, 16'd35795, 16'd39668, 16'd60745, 16'd19146, 16'd57532, 16'd37127, 16'd40455, 16'd59512, 16'd42041, 16'd60634, 16'd27102, 16'd8576, 16'd54567, 16'd25882, 16'd50980, 16'd47246, 16'd32084, 16'd20896});
	test_expansion(128'hb62de4254e35b81f2da1f75fd3dea50f, {16'd64061, 16'd4187, 16'd27151, 16'd29300, 16'd44857, 16'd20172, 16'd5785, 16'd35664, 16'd42891, 16'd12467, 16'd49466, 16'd12541, 16'd61422, 16'd40603, 16'd13780, 16'd58157, 16'd30016, 16'd14699, 16'd60838, 16'd20044, 16'd36781, 16'd13520, 16'd17749, 16'd41760, 16'd23394, 16'd27413});
	test_expansion(128'ha88c56d93015b4faa393893e0a0c4a9c, {16'd17196, 16'd8716, 16'd57303, 16'd11779, 16'd29386, 16'd62398, 16'd10318, 16'd28378, 16'd44408, 16'd47388, 16'd29558, 16'd49330, 16'd51849, 16'd37483, 16'd44251, 16'd53718, 16'd53244, 16'd24227, 16'd47621, 16'd4322, 16'd30360, 16'd48953, 16'd16021, 16'd63431, 16'd23985, 16'd29322});
	test_expansion(128'h5a45077247bccc84b05620c3023d4669, {16'd19569, 16'd50659, 16'd54211, 16'd44897, 16'd60653, 16'd61178, 16'd57879, 16'd53561, 16'd6586, 16'd13567, 16'd13996, 16'd1368, 16'd15812, 16'd43647, 16'd20704, 16'd60413, 16'd21209, 16'd16839, 16'd8038, 16'd8654, 16'd29907, 16'd25591, 16'd24582, 16'd22420, 16'd25574, 16'd46466});
	test_expansion(128'ha243cdb6663ce7b00f2f2d4e2486342f, {16'd25209, 16'd44995, 16'd27898, 16'd33282, 16'd885, 16'd51140, 16'd51962, 16'd37669, 16'd11140, 16'd53487, 16'd41457, 16'd15672, 16'd22504, 16'd34222, 16'd1294, 16'd63490, 16'd59651, 16'd61745, 16'd36814, 16'd39323, 16'd41915, 16'd22341, 16'd13450, 16'd38396, 16'd29354, 16'd45317});
	test_expansion(128'h3bed3cb4f753127c1468a6d6938b1622, {16'd28099, 16'd31718, 16'd20085, 16'd36016, 16'd26771, 16'd24614, 16'd54430, 16'd22970, 16'd24890, 16'd54321, 16'd29064, 16'd52490, 16'd46788, 16'd16523, 16'd47223, 16'd23931, 16'd39701, 16'd26488, 16'd53864, 16'd49130, 16'd52920, 16'd6566, 16'd10881, 16'd36170, 16'd5135, 16'd50193});
	test_expansion(128'h292161bf93fdfcedd7294b9a974c3afd, {16'd45686, 16'd55119, 16'd30155, 16'd27257, 16'd59964, 16'd3485, 16'd13841, 16'd44862, 16'd49997, 16'd58642, 16'd31040, 16'd16731, 16'd40840, 16'd13849, 16'd55543, 16'd49791, 16'd37522, 16'd9813, 16'd30271, 16'd1734, 16'd11790, 16'd30814, 16'd7084, 16'd36508, 16'd52648, 16'd8926});
	test_expansion(128'h0f6d38b7dcdc7a8210ea2856b733c933, {16'd13446, 16'd46025, 16'd1681, 16'd18230, 16'd45908, 16'd46300, 16'd57819, 16'd4698, 16'd52256, 16'd48731, 16'd43622, 16'd58206, 16'd51036, 16'd33542, 16'd49448, 16'd14274, 16'd8922, 16'd3331, 16'd13298, 16'd21649, 16'd9952, 16'd29446, 16'd65381, 16'd13099, 16'd46880, 16'd34166});
	test_expansion(128'hd753f16534268366247ae13f84e39c6a, {16'd32683, 16'd60612, 16'd42199, 16'd41320, 16'd55639, 16'd8647, 16'd24666, 16'd26080, 16'd24542, 16'd38388, 16'd38610, 16'd44644, 16'd16675, 16'd18981, 16'd23297, 16'd11401, 16'd48410, 16'd37368, 16'd16350, 16'd5826, 16'd5135, 16'd8503, 16'd61559, 16'd22623, 16'd12566, 16'd22642});
	test_expansion(128'hd5ef4ad8eb62a1fb00f1cfa69187edcd, {16'd29260, 16'd14886, 16'd37569, 16'd27421, 16'd5292, 16'd16081, 16'd6638, 16'd27575, 16'd54966, 16'd55612, 16'd5831, 16'd23791, 16'd29071, 16'd19680, 16'd14521, 16'd43708, 16'd13985, 16'd50153, 16'd16843, 16'd20784, 16'd21956, 16'd54401, 16'd56895, 16'd14080, 16'd60025, 16'd3952});
	test_expansion(128'h4397eeac188d118a5a225aa134ab635a, {16'd55879, 16'd42001, 16'd56859, 16'd46588, 16'd50192, 16'd9198, 16'd36198, 16'd21971, 16'd27518, 16'd28006, 16'd22826, 16'd9462, 16'd48585, 16'd8896, 16'd27547, 16'd5825, 16'd35126, 16'd33004, 16'd41571, 16'd37890, 16'd64642, 16'd13704, 16'd47488, 16'd63169, 16'd63002, 16'd17709});
	test_expansion(128'h820bf92812599e61fc57a758fd12b896, {16'd5676, 16'd7510, 16'd57905, 16'd58779, 16'd47255, 16'd24305, 16'd61300, 16'd26467, 16'd51593, 16'd25938, 16'd47843, 16'd51742, 16'd25256, 16'd64036, 16'd31618, 16'd37077, 16'd53510, 16'd37472, 16'd29998, 16'd26961, 16'd47888, 16'd31802, 16'd40226, 16'd45344, 16'd8109, 16'd16925});
	test_expansion(128'h08cac6effd1e8a6fd9148c5bac2ff677, {16'd54215, 16'd1845, 16'd46238, 16'd60477, 16'd54248, 16'd44662, 16'd34010, 16'd5575, 16'd48879, 16'd24387, 16'd16681, 16'd46905, 16'd56306, 16'd28885, 16'd61590, 16'd48241, 16'd41327, 16'd13109, 16'd34580, 16'd26000, 16'd51497, 16'd10133, 16'd3901, 16'd62369, 16'd19882, 16'd20773});
	test_expansion(128'h4d7bff135b93a29619d868c7f4f0e4a2, {16'd44222, 16'd56632, 16'd64160, 16'd51376, 16'd2699, 16'd49131, 16'd62221, 16'd57690, 16'd8383, 16'd8434, 16'd64910, 16'd40354, 16'd59105, 16'd25611, 16'd10234, 16'd12984, 16'd2621, 16'd50233, 16'd27685, 16'd4126, 16'd21907, 16'd61078, 16'd61169, 16'd50263, 16'd26689, 16'd52617});
	test_expansion(128'h897dbe9f2d03583d4f378fd93d59abe1, {16'd58663, 16'd11527, 16'd1295, 16'd27352, 16'd36363, 16'd20290, 16'd54225, 16'd56852, 16'd60783, 16'd61601, 16'd63026, 16'd38264, 16'd32756, 16'd45656, 16'd18838, 16'd14625, 16'd8036, 16'd64395, 16'd55302, 16'd61673, 16'd57546, 16'd6181, 16'd44577, 16'd51757, 16'd41473, 16'd31340});
	test_expansion(128'h34511566e5bc3744ca88697665876f44, {16'd18863, 16'd6024, 16'd40640, 16'd55337, 16'd3471, 16'd36977, 16'd48175, 16'd34150, 16'd2733, 16'd47216, 16'd4581, 16'd30351, 16'd46548, 16'd1168, 16'd50319, 16'd32697, 16'd23053, 16'd58856, 16'd37110, 16'd65179, 16'd24711, 16'd37051, 16'd3172, 16'd55462, 16'd37358, 16'd59857});
	test_expansion(128'he2adab98382094567214134a87a563fc, {16'd29722, 16'd11809, 16'd44350, 16'd44062, 16'd19184, 16'd45718, 16'd55382, 16'd7280, 16'd38433, 16'd39682, 16'd39137, 16'd59439, 16'd8434, 16'd1430, 16'd29518, 16'd38289, 16'd51252, 16'd2369, 16'd55582, 16'd29794, 16'd10397, 16'd31212, 16'd60555, 16'd48053, 16'd62227, 16'd45206});
	test_expansion(128'h56700b5ad3525ca39ccca8d2d55392a9, {16'd37695, 16'd50909, 16'd39077, 16'd59916, 16'd29295, 16'd31393, 16'd37684, 16'd45599, 16'd52959, 16'd23262, 16'd49350, 16'd62926, 16'd18137, 16'd3484, 16'd37561, 16'd7486, 16'd25403, 16'd54746, 16'd34459, 16'd64290, 16'd37963, 16'd32526, 16'd49581, 16'd40305, 16'd53277, 16'd61874});
	test_expansion(128'h5f35284aee871f60efdfb4f2634900f3, {16'd11084, 16'd41958, 16'd23784, 16'd18336, 16'd3419, 16'd20774, 16'd45116, 16'd55251, 16'd54796, 16'd15804, 16'd62697, 16'd45964, 16'd60263, 16'd19738, 16'd30491, 16'd547, 16'd58875, 16'd36273, 16'd62141, 16'd32320, 16'd54375, 16'd37467, 16'd658, 16'd60765, 16'd42685, 16'd27764});
	test_expansion(128'h697ea3e5966f30fbf3ec59128c15dadf, {16'd24050, 16'd30545, 16'd39155, 16'd19615, 16'd43823, 16'd46116, 16'd10007, 16'd46237, 16'd102, 16'd40787, 16'd62634, 16'd30057, 16'd46266, 16'd42176, 16'd50976, 16'd53617, 16'd26404, 16'd26560, 16'd40168, 16'd51644, 16'd21523, 16'd40051, 16'd32466, 16'd51833, 16'd30890, 16'd29523});
	test_expansion(128'ha92d761a155d1fb995c16eb049bd98ae, {16'd48632, 16'd48109, 16'd12388, 16'd41829, 16'd28914, 16'd60520, 16'd37097, 16'd54436, 16'd46691, 16'd22060, 16'd59140, 16'd4869, 16'd14623, 16'd43652, 16'd28274, 16'd59982, 16'd55669, 16'd52351, 16'd64984, 16'd18802, 16'd47592, 16'd45844, 16'd62622, 16'd25438, 16'd51775, 16'd12285});
	test_expansion(128'hebd32255f75fa0d7bb674ca8cd34acda, {16'd28879, 16'd25226, 16'd63322, 16'd53896, 16'd39360, 16'd39140, 16'd28447, 16'd40706, 16'd17280, 16'd56347, 16'd30347, 16'd54731, 16'd11178, 16'd60464, 16'd3987, 16'd34202, 16'd54074, 16'd57999, 16'd36364, 16'd55470, 16'd40597, 16'd61646, 16'd33527, 16'd42279, 16'd1427, 16'd7883});
	test_expansion(128'h19f5971a2bd4af9e89e95ff9f27c8cd7, {16'd28224, 16'd19257, 16'd63666, 16'd35278, 16'd36123, 16'd46375, 16'd35101, 16'd62351, 16'd11456, 16'd8660, 16'd45455, 16'd47670, 16'd6058, 16'd25017, 16'd9840, 16'd33104, 16'd23276, 16'd64358, 16'd27813, 16'd9803, 16'd45680, 16'd38357, 16'd6769, 16'd26757, 16'd51080, 16'd55239});
	test_expansion(128'h23609cb9ce564498bc02f831e098c38d, {16'd46369, 16'd55458, 16'd58192, 16'd5987, 16'd61652, 16'd63835, 16'd24258, 16'd53142, 16'd19408, 16'd28139, 16'd16900, 16'd55045, 16'd37117, 16'd42198, 16'd33446, 16'd58073, 16'd11397, 16'd1872, 16'd50441, 16'd17635, 16'd35234, 16'd59233, 16'd38093, 16'd47152, 16'd23350, 16'd60442});
	test_expansion(128'h57c38906f90b2e151105b8b27eeaf066, {16'd12475, 16'd62147, 16'd45305, 16'd12550, 16'd41615, 16'd19472, 16'd12320, 16'd45335, 16'd10419, 16'd54827, 16'd38945, 16'd56027, 16'd13096, 16'd19770, 16'd45151, 16'd15367, 16'd7522, 16'd21605, 16'd37871, 16'd36568, 16'd8634, 16'd28232, 16'd20596, 16'd10970, 16'd44201, 16'd52255});
	test_expansion(128'h93ebed0e9ba2f4fbec75da59ee04c311, {16'd42648, 16'd496, 16'd39468, 16'd46432, 16'd7541, 16'd45901, 16'd51750, 16'd59834, 16'd65408, 16'd30488, 16'd49724, 16'd50206, 16'd20597, 16'd36403, 16'd24651, 16'd49522, 16'd63129, 16'd15569, 16'd37256, 16'd65289, 16'd29792, 16'd18081, 16'd12186, 16'd58784, 16'd36956, 16'd9285});
	test_expansion(128'h518f116d1b5cf43c6a60c4f4054f1197, {16'd28780, 16'd49856, 16'd21671, 16'd56759, 16'd61785, 16'd37596, 16'd48725, 16'd18621, 16'd12857, 16'd52323, 16'd53849, 16'd50458, 16'd43004, 16'd11785, 16'd37326, 16'd37636, 16'd49002, 16'd6600, 16'd10770, 16'd18154, 16'd52474, 16'd26031, 16'd31574, 16'd48641, 16'd45636, 16'd5040});
	test_expansion(128'hac5da3364ed5fe0eccfea078868c4fe5, {16'd35306, 16'd58695, 16'd64581, 16'd7297, 16'd61130, 16'd10124, 16'd55586, 16'd28400, 16'd51982, 16'd7149, 16'd15813, 16'd3428, 16'd53952, 16'd56440, 16'd48866, 16'd43020, 16'd52059, 16'd2047, 16'd7902, 16'd594, 16'd55141, 16'd30676, 16'd33099, 16'd37152, 16'd35657, 16'd8263});
	test_expansion(128'h318b11065c183f6440cbed74e48dea26, {16'd26757, 16'd41069, 16'd7920, 16'd36201, 16'd8958, 16'd26663, 16'd61982, 16'd5431, 16'd15915, 16'd13977, 16'd9186, 16'd59581, 16'd15006, 16'd46818, 16'd19273, 16'd22615, 16'd40076, 16'd43968, 16'd56831, 16'd43072, 16'd31240, 16'd2277, 16'd50351, 16'd64954, 16'd47273, 16'd10790});
	test_expansion(128'h1bf9351aa83cd4fc2b041c2cecc2de38, {16'd33983, 16'd44610, 16'd47131, 16'd421, 16'd2185, 16'd52544, 16'd10118, 16'd38145, 16'd27283, 16'd18542, 16'd18137, 16'd24950, 16'd10088, 16'd31338, 16'd15651, 16'd36426, 16'd61275, 16'd11344, 16'd23585, 16'd14987, 16'd29755, 16'd8674, 16'd28090, 16'd49452, 16'd13618, 16'd49144});
	test_expansion(128'h70a16a2841abb4bad891751d330d2fa1, {16'd57542, 16'd26090, 16'd16262, 16'd59719, 16'd14618, 16'd36723, 16'd61160, 16'd18384, 16'd60037, 16'd42193, 16'd26502, 16'd27855, 16'd9228, 16'd1930, 16'd420, 16'd51346, 16'd57457, 16'd61446, 16'd6407, 16'd29604, 16'd22319, 16'd33829, 16'd48963, 16'd41911, 16'd2375, 16'd28069});
	test_expansion(128'hb66f78ec4dafd890e081cc765a517bff, {16'd44731, 16'd3984, 16'd55809, 16'd59145, 16'd62380, 16'd16729, 16'd48183, 16'd26887, 16'd30698, 16'd40683, 16'd3594, 16'd10274, 16'd26178, 16'd53811, 16'd9115, 16'd35309, 16'd63996, 16'd28774, 16'd46548, 16'd44096, 16'd10987, 16'd56275, 16'd18471, 16'd64942, 16'd42334, 16'd62115});
	test_expansion(128'h4f795c5e368b145e8002035b78f1f4f8, {16'd45023, 16'd58569, 16'd50362, 16'd62028, 16'd53728, 16'd8370, 16'd55281, 16'd29801, 16'd28997, 16'd2596, 16'd42436, 16'd18720, 16'd42552, 16'd39987, 16'd33942, 16'd18988, 16'd35298, 16'd39888, 16'd32922, 16'd27565, 16'd52948, 16'd9782, 16'd23474, 16'd7960, 16'd7631, 16'd3505});
	test_expansion(128'h9f2f3f100e78aa230f419f4bbe3b4898, {16'd60068, 16'd25341, 16'd37433, 16'd19693, 16'd63704, 16'd16357, 16'd39267, 16'd30629, 16'd55022, 16'd23569, 16'd5686, 16'd56419, 16'd57283, 16'd64701, 16'd39557, 16'd31649, 16'd22147, 16'd8524, 16'd51511, 16'd30571, 16'd43427, 16'd62149, 16'd43787, 16'd21111, 16'd47321, 16'd38802});
	test_expansion(128'h6cbaa6ad8374e21625bbed1dba767a5c, {16'd32442, 16'd3355, 16'd40050, 16'd49172, 16'd9570, 16'd21416, 16'd46866, 16'd5573, 16'd42983, 16'd21920, 16'd57120, 16'd55538, 16'd54542, 16'd23767, 16'd13143, 16'd25852, 16'd64197, 16'd47492, 16'd7077, 16'd61038, 16'd5619, 16'd24142, 16'd60894, 16'd26983, 16'd29753, 16'd14524});
	test_expansion(128'ha444f75cc2858b63d4d4d5a210136b9b, {16'd43387, 16'd17695, 16'd21160, 16'd1726, 16'd59764, 16'd14694, 16'd7726, 16'd23160, 16'd12101, 16'd33659, 16'd49342, 16'd17145, 16'd49680, 16'd63465, 16'd54812, 16'd24697, 16'd49927, 16'd19733, 16'd43338, 16'd29786, 16'd20107, 16'd42536, 16'd36009, 16'd24459, 16'd5027, 16'd20151});
	test_expansion(128'hf371fcf90ebbe8bafa96678eac6d5358, {16'd10687, 16'd22302, 16'd35527, 16'd61472, 16'd8549, 16'd34219, 16'd48190, 16'd9064, 16'd21888, 16'd14059, 16'd15818, 16'd22786, 16'd50538, 16'd7732, 16'd49727, 16'd48876, 16'd58360, 16'd7459, 16'd23854, 16'd61523, 16'd11589, 16'd49806, 16'd28932, 16'd44534, 16'd63305, 16'd61642});
	test_expansion(128'h7309cb0311c192eda881f8306df25719, {16'd18741, 16'd29983, 16'd54980, 16'd57048, 16'd7720, 16'd31845, 16'd55973, 16'd3667, 16'd42060, 16'd48314, 16'd44294, 16'd56651, 16'd2974, 16'd52193, 16'd19751, 16'd37260, 16'd31776, 16'd41841, 16'd6588, 16'd59667, 16'd11111, 16'd41828, 16'd20713, 16'd17860, 16'd16061, 16'd573});
	test_expansion(128'h05e19baaca26d9ad12bd4961783dc6c0, {16'd13155, 16'd15948, 16'd44167, 16'd15406, 16'd31031, 16'd30718, 16'd9362, 16'd17731, 16'd46796, 16'd28937, 16'd37457, 16'd47372, 16'd32850, 16'd26129, 16'd56107, 16'd56608, 16'd57340, 16'd56549, 16'd33005, 16'd20094, 16'd40516, 16'd50568, 16'd40487, 16'd38483, 16'd649, 16'd14470});
	test_expansion(128'hfea5a83879072fc49d3cfbbcbbe09377, {16'd53047, 16'd50097, 16'd3251, 16'd21770, 16'd59115, 16'd44006, 16'd14407, 16'd63388, 16'd57965, 16'd53297, 16'd45547, 16'd34993, 16'd44143, 16'd56164, 16'd48478, 16'd44190, 16'd1426, 16'd49497, 16'd34886, 16'd18044, 16'd41801, 16'd10803, 16'd39502, 16'd29261, 16'd45459, 16'd3954});
	test_expansion(128'h8f04e3974dc70bf56aa2fa0e62b21ce3, {16'd55469, 16'd60984, 16'd55588, 16'd48710, 16'd11581, 16'd19336, 16'd26304, 16'd38451, 16'd22852, 16'd57209, 16'd54328, 16'd53691, 16'd19038, 16'd46900, 16'd1492, 16'd52495, 16'd47067, 16'd15419, 16'd15682, 16'd55356, 16'd46127, 16'd45058, 16'd2022, 16'd48285, 16'd43764, 16'd37003});
	test_expansion(128'h754f2991629ad5c6d9d9e62596235e78, {16'd16183, 16'd12832, 16'd59867, 16'd65225, 16'd43669, 16'd16092, 16'd64769, 16'd3648, 16'd52987, 16'd64207, 16'd14238, 16'd37009, 16'd19777, 16'd51409, 16'd2577, 16'd6689, 16'd40103, 16'd5439, 16'd17862, 16'd29690, 16'd63131, 16'd57287, 16'd49282, 16'd15215, 16'd17313, 16'd24292});
	test_expansion(128'hc9791f82eee9d42eec028b49d3abc09e, {16'd14899, 16'd8768, 16'd37991, 16'd19262, 16'd42145, 16'd60972, 16'd32565, 16'd5586, 16'd17106, 16'd32222, 16'd10317, 16'd47282, 16'd51124, 16'd23411, 16'd55669, 16'd29420, 16'd58058, 16'd623, 16'd35419, 16'd17744, 16'd39931, 16'd35370, 16'd28692, 16'd37679, 16'd39496, 16'd49195});
	test_expansion(128'hb5263791907221b89d09389bb5c21778, {16'd55987, 16'd12150, 16'd14852, 16'd9136, 16'd48266, 16'd11163, 16'd52063, 16'd62861, 16'd61744, 16'd15866, 16'd3617, 16'd42403, 16'd10754, 16'd45712, 16'd5910, 16'd38213, 16'd271, 16'd58311, 16'd15716, 16'd27697, 16'd54705, 16'd45772, 16'd7019, 16'd6111, 16'd28092, 16'd6512});
	test_expansion(128'h2d98577e3ce0e6f64a6239ad43a4e494, {16'd20737, 16'd33526, 16'd4673, 16'd30126, 16'd18936, 16'd21490, 16'd30907, 16'd28359, 16'd44466, 16'd22085, 16'd36003, 16'd3493, 16'd24359, 16'd64870, 16'd10945, 16'd37117, 16'd4303, 16'd44039, 16'd12774, 16'd54719, 16'd41944, 16'd14872, 16'd106, 16'd28753, 16'd13039, 16'd15246});
	test_expansion(128'h129c4f2af41a85a58b025fc446fca592, {16'd55342, 16'd62540, 16'd40466, 16'd35192, 16'd41374, 16'd12642, 16'd54189, 16'd7883, 16'd27240, 16'd23842, 16'd62816, 16'd3294, 16'd54286, 16'd17831, 16'd5739, 16'd26899, 16'd23839, 16'd62737, 16'd4767, 16'd49813, 16'd53057, 16'd4488, 16'd8136, 16'd33861, 16'd50038, 16'd24402});
	test_expansion(128'h207cd69c040417997bb1a76ac0659edf, {16'd10464, 16'd61770, 16'd29032, 16'd18292, 16'd11168, 16'd43405, 16'd9913, 16'd57858, 16'd45791, 16'd13916, 16'd31274, 16'd22001, 16'd13232, 16'd51123, 16'd32039, 16'd18563, 16'd7718, 16'd55806, 16'd42111, 16'd43927, 16'd27446, 16'd49550, 16'd24672, 16'd3891, 16'd15383, 16'd31319});
	test_expansion(128'h647f2db80db414683884a41d26036d4f, {16'd64429, 16'd5358, 16'd18598, 16'd32479, 16'd560, 16'd22650, 16'd49151, 16'd37734, 16'd60766, 16'd10905, 16'd52350, 16'd16435, 16'd33184, 16'd46522, 16'd3537, 16'd56976, 16'd30148, 16'd59755, 16'd60987, 16'd880, 16'd19601, 16'd41814, 16'd60569, 16'd15441, 16'd12086, 16'd45228});
	test_expansion(128'had6552ee86b85e03139fb87d330510e1, {16'd36299, 16'd12662, 16'd28917, 16'd38413, 16'd56327, 16'd25983, 16'd51936, 16'd56445, 16'd17342, 16'd49149, 16'd51528, 16'd62467, 16'd9848, 16'd16877, 16'd46392, 16'd41313, 16'd65533, 16'd33147, 16'd57419, 16'd4867, 16'd23793, 16'd64181, 16'd62115, 16'd61896, 16'd34684, 16'd25194});
	test_expansion(128'h05270adc0f8390013a1422628c179c32, {16'd34391, 16'd64036, 16'd24842, 16'd1394, 16'd57944, 16'd42216, 16'd57223, 16'd28064, 16'd8001, 16'd6711, 16'd48731, 16'd13449, 16'd32136, 16'd40032, 16'd27102, 16'd22105, 16'd364, 16'd13260, 16'd22628, 16'd50611, 16'd13513, 16'd17792, 16'd26337, 16'd23140, 16'd41023, 16'd61464});
	test_expansion(128'hb6ab535e8bce0024e8eb58770a03ad59, {16'd5383, 16'd34699, 16'd37889, 16'd15636, 16'd23011, 16'd44268, 16'd13548, 16'd23985, 16'd51494, 16'd41527, 16'd32782, 16'd21656, 16'd7195, 16'd33002, 16'd7396, 16'd60383, 16'd5432, 16'd46015, 16'd35228, 16'd46512, 16'd2475, 16'd54533, 16'd52652, 16'd30789, 16'd12604, 16'd4886});
	test_expansion(128'hb7e267359c049f991f4a68c418c54fa4, {16'd58284, 16'd36983, 16'd20451, 16'd28259, 16'd29573, 16'd19317, 16'd57101, 16'd65514, 16'd11342, 16'd38416, 16'd46548, 16'd56087, 16'd13335, 16'd30823, 16'd20832, 16'd60407, 16'd58314, 16'd22392, 16'd21337, 16'd4167, 16'd42727, 16'd38973, 16'd42405, 16'd51478, 16'd64671, 16'd44865});
	test_expansion(128'h6b527e3d131af2d2a50dac7fe497e2fa, {16'd11816, 16'd23146, 16'd10956, 16'd38958, 16'd2155, 16'd29852, 16'd26752, 16'd59193, 16'd54161, 16'd8390, 16'd11898, 16'd48132, 16'd61770, 16'd49371, 16'd44622, 16'd1491, 16'd51076, 16'd21141, 16'd31320, 16'd15584, 16'd23467, 16'd47826, 16'd39707, 16'd3212, 16'd33407, 16'd31137});
	test_expansion(128'h582c8b730a7a17217d5dcfe4e54bbe0b, {16'd35711, 16'd34343, 16'd24782, 16'd46822, 16'd62279, 16'd59183, 16'd54803, 16'd8924, 16'd53801, 16'd63584, 16'd20742, 16'd20439, 16'd20289, 16'd47700, 16'd56918, 16'd30916, 16'd38859, 16'd50295, 16'd52385, 16'd55000, 16'd49547, 16'd52233, 16'd36086, 16'd7771, 16'd3380, 16'd10546});
	test_expansion(128'hd8702fc37661f38d797ecfc274634928, {16'd9118, 16'd33187, 16'd23067, 16'd64135, 16'd2631, 16'd9183, 16'd15894, 16'd48162, 16'd40958, 16'd29233, 16'd63026, 16'd56736, 16'd10636, 16'd2803, 16'd17525, 16'd3844, 16'd17608, 16'd9082, 16'd56899, 16'd47643, 16'd43608, 16'd40972, 16'd52330, 16'd28401, 16'd57206, 16'd48937});
	test_expansion(128'h39482075ca27ccb85ece1929310765ee, {16'd51543, 16'd967, 16'd28467, 16'd710, 16'd29149, 16'd35681, 16'd22974, 16'd2910, 16'd1393, 16'd30789, 16'd25246, 16'd12570, 16'd58555, 16'd62183, 16'd4409, 16'd63294, 16'd9630, 16'd6825, 16'd50801, 16'd10969, 16'd3636, 16'd6111, 16'd53640, 16'd50498, 16'd21114, 16'd28258});
	test_expansion(128'hb16e24bc6e439dfb99b90f3af23a94b0, {16'd50442, 16'd28648, 16'd6444, 16'd38107, 16'd35284, 16'd58908, 16'd19697, 16'd65199, 16'd7592, 16'd61156, 16'd28557, 16'd56388, 16'd31600, 16'd56337, 16'd7308, 16'd27826, 16'd34611, 16'd64577, 16'd611, 16'd44438, 16'd58407, 16'd53075, 16'd61704, 16'd56230, 16'd18858, 16'd17873});
	test_expansion(128'h0fae991bfb7915d5729143335b5af564, {16'd14067, 16'd18910, 16'd29170, 16'd49531, 16'd38098, 16'd61548, 16'd4658, 16'd42872, 16'd49253, 16'd33991, 16'd32695, 16'd722, 16'd7697, 16'd47652, 16'd488, 16'd9176, 16'd27258, 16'd39179, 16'd41624, 16'd40216, 16'd37925, 16'd60062, 16'd1631, 16'd34533, 16'd8428, 16'd14232});
	test_expansion(128'h81da7761df2203765e696b9d3633a2bc, {16'd32577, 16'd10610, 16'd45287, 16'd56396, 16'd24656, 16'd17588, 16'd20280, 16'd61158, 16'd57529, 16'd46994, 16'd45430, 16'd8000, 16'd31747, 16'd5836, 16'd13323, 16'd24928, 16'd18729, 16'd62473, 16'd48613, 16'd24058, 16'd61435, 16'd36618, 16'd3276, 16'd2580, 16'd33024, 16'd55693});
	test_expansion(128'h7e81a78a2b4b4bd34d1157e37284c36d, {16'd49388, 16'd9105, 16'd39844, 16'd9891, 16'd60818, 16'd1471, 16'd46689, 16'd43914, 16'd8920, 16'd21873, 16'd17021, 16'd43632, 16'd59955, 16'd40894, 16'd52627, 16'd47975, 16'd57648, 16'd23695, 16'd8209, 16'd8452, 16'd17548, 16'd4281, 16'd61938, 16'd57672, 16'd59512, 16'd62123});
	test_expansion(128'h286c19de4abaac2bcb05708487ec5428, {16'd10070, 16'd36602, 16'd21036, 16'd22132, 16'd48731, 16'd64104, 16'd40777, 16'd25586, 16'd840, 16'd58025, 16'd12835, 16'd13221, 16'd46350, 16'd836, 16'd41999, 16'd25261, 16'd43087, 16'd45762, 16'd40487, 16'd30449, 16'd57741, 16'd8422, 16'd16325, 16'd1196, 16'd63707, 16'd52544});
	test_expansion(128'hc70f9a9078d0a340f2102ba7ab29e57b, {16'd41152, 16'd8561, 16'd20580, 16'd37013, 16'd48492, 16'd631, 16'd25399, 16'd25955, 16'd63181, 16'd18508, 16'd25865, 16'd52537, 16'd27272, 16'd26458, 16'd31117, 16'd62725, 16'd49625, 16'd41381, 16'd51877, 16'd13664, 16'd15563, 16'd33823, 16'd12190, 16'd8697, 16'd17097, 16'd49164});
	test_expansion(128'hc92ff2a2010619c649e81463986675f5, {16'd57638, 16'd35422, 16'd64536, 16'd32826, 16'd49974, 16'd13924, 16'd26724, 16'd16887, 16'd59722, 16'd12268, 16'd24302, 16'd18526, 16'd17316, 16'd10649, 16'd715, 16'd2018, 16'd1476, 16'd5934, 16'd65467, 16'd23862, 16'd58433, 16'd30927, 16'd25560, 16'd9059, 16'd19271, 16'd44903});
	test_expansion(128'h639c2c94e8a0e7019e1c26e7b5595e9d, {16'd19847, 16'd5482, 16'd28215, 16'd19125, 16'd12945, 16'd31923, 16'd61972, 16'd40389, 16'd49291, 16'd42535, 16'd33032, 16'd1732, 16'd20633, 16'd52934, 16'd25611, 16'd30781, 16'd56038, 16'd17807, 16'd35915, 16'd4319, 16'd15473, 16'd24042, 16'd11401, 16'd50866, 16'd41539, 16'd51027});
	test_expansion(128'h260e4fb8a77ff1082570ef24f986bdcd, {16'd44263, 16'd41640, 16'd18870, 16'd19542, 16'd37416, 16'd49399, 16'd5559, 16'd36220, 16'd43283, 16'd38775, 16'd58504, 16'd54493, 16'd49266, 16'd50214, 16'd33223, 16'd52799, 16'd56801, 16'd5834, 16'd28553, 16'd6140, 16'd12959, 16'd6516, 16'd9375, 16'd28451, 16'd5601, 16'd1726});
	test_expansion(128'h6484632714171f53bad3e57e425dc9ed, {16'd61487, 16'd14785, 16'd2878, 16'd49117, 16'd48617, 16'd12516, 16'd7355, 16'd63103, 16'd51751, 16'd64397, 16'd63769, 16'd48421, 16'd40866, 16'd63003, 16'd25029, 16'd56635, 16'd19070, 16'd65139, 16'd43973, 16'd18794, 16'd17297, 16'd38693, 16'd12798, 16'd14473, 16'd30919, 16'd62196});
	test_expansion(128'he6f5150e63ffee2d746327defbc87a5f, {16'd3928, 16'd52203, 16'd43530, 16'd5984, 16'd28877, 16'd35609, 16'd55202, 16'd63425, 16'd53584, 16'd33825, 16'd1949, 16'd9331, 16'd45684, 16'd1758, 16'd56388, 16'd261, 16'd30712, 16'd52032, 16'd21062, 16'd45334, 16'd22680, 16'd62357, 16'd20148, 16'd54586, 16'd44200, 16'd30081});
	test_expansion(128'h96566ea86a75cbb0e48c17332747d3d8, {16'd52806, 16'd39454, 16'd65364, 16'd11406, 16'd48009, 16'd19580, 16'd16628, 16'd43470, 16'd53833, 16'd18827, 16'd26114, 16'd50944, 16'd12893, 16'd30110, 16'd58492, 16'd16874, 16'd28635, 16'd28907, 16'd25191, 16'd61805, 16'd65014, 16'd45128, 16'd47148, 16'd47011, 16'd50180, 16'd16004});
	test_expansion(128'he46a5d416fdf7a1864705827a2ac7a79, {16'd57091, 16'd20605, 16'd13122, 16'd64924, 16'd64009, 16'd8403, 16'd2632, 16'd10732, 16'd29951, 16'd1237, 16'd909, 16'd32498, 16'd46833, 16'd45502, 16'd25957, 16'd16002, 16'd17161, 16'd33212, 16'd40628, 16'd45129, 16'd46108, 16'd5498, 16'd12610, 16'd29078, 16'd19915, 16'd20664});
	test_expansion(128'h9ca78e0ee1e8c015451c896c7128c625, {16'd12214, 16'd13541, 16'd33743, 16'd2048, 16'd15011, 16'd15275, 16'd52245, 16'd39155, 16'd3147, 16'd54892, 16'd25893, 16'd17830, 16'd14110, 16'd41706, 16'd4424, 16'd44816, 16'd7405, 16'd6439, 16'd28996, 16'd50255, 16'd47592, 16'd2486, 16'd38958, 16'd15084, 16'd12590, 16'd37725});
	test_expansion(128'h57cfab073202bfc1cca849a930257a7b, {16'd33179, 16'd59114, 16'd18101, 16'd43205, 16'd55559, 16'd6818, 16'd45201, 16'd51642, 16'd10453, 16'd51739, 16'd48713, 16'd23750, 16'd50031, 16'd37667, 16'd36660, 16'd65144, 16'd50667, 16'd3396, 16'd5601, 16'd3782, 16'd42378, 16'd5433, 16'd59463, 16'd18665, 16'd32555, 16'd6533});
	test_expansion(128'h472001831c05321236e6f160b0a767bf, {16'd62317, 16'd6524, 16'd39371, 16'd13320, 16'd62932, 16'd19799, 16'd19881, 16'd2922, 16'd18033, 16'd1700, 16'd51162, 16'd46558, 16'd35411, 16'd38008, 16'd57901, 16'd48970, 16'd48760, 16'd51280, 16'd43961, 16'd43, 16'd57150, 16'd10885, 16'd41930, 16'd13208, 16'd48115, 16'd13672});
	test_expansion(128'h397fe2afab0f06aeab28b9038539c968, {16'd59, 16'd24894, 16'd51626, 16'd22412, 16'd7372, 16'd51939, 16'd6137, 16'd29193, 16'd49220, 16'd53119, 16'd4591, 16'd20402, 16'd2644, 16'd41281, 16'd44673, 16'd50652, 16'd832, 16'd23892, 16'd19664, 16'd26384, 16'd37517, 16'd65397, 16'd43731, 16'd61747, 16'd9338, 16'd38573});
	test_expansion(128'h2093f1806f6ec715a96c572d9b85a4ed, {16'd42898, 16'd26632, 16'd41363, 16'd16071, 16'd57130, 16'd22446, 16'd30748, 16'd55320, 16'd25875, 16'd15669, 16'd53062, 16'd10555, 16'd55889, 16'd57078, 16'd33921, 16'd15798, 16'd44995, 16'd34644, 16'd18178, 16'd56045, 16'd17434, 16'd62325, 16'd6249, 16'd59785, 16'd6539, 16'd51510});
	test_expansion(128'h30e077514284f6f6002fc91d05c161ba, {16'd37734, 16'd22885, 16'd64354, 16'd51141, 16'd33975, 16'd52824, 16'd45706, 16'd17790, 16'd19732, 16'd10498, 16'd35141, 16'd13944, 16'd19169, 16'd1603, 16'd63431, 16'd50176, 16'd8679, 16'd49049, 16'd52999, 16'd38937, 16'd44500, 16'd11849, 16'd29123, 16'd6498, 16'd44735, 16'd14101});
	test_expansion(128'hf69ab666bba6403908fd42861743d3d2, {16'd44090, 16'd57726, 16'd55464, 16'd63531, 16'd39255, 16'd12500, 16'd52814, 16'd54242, 16'd27436, 16'd46599, 16'd43120, 16'd58927, 16'd13597, 16'd42866, 16'd12708, 16'd1319, 16'd28043, 16'd6507, 16'd25626, 16'd16105, 16'd44706, 16'd32826, 16'd42775, 16'd7601, 16'd55875, 16'd35094});
	test_expansion(128'hdc400e100c49a1924f5130550a6c2318, {16'd49020, 16'd44650, 16'd19051, 16'd971, 16'd20638, 16'd37607, 16'd55811, 16'd31641, 16'd34823, 16'd11449, 16'd8009, 16'd12212, 16'd11859, 16'd134, 16'd59264, 16'd55850, 16'd6747, 16'd43842, 16'd13470, 16'd6869, 16'd57465, 16'd9955, 16'd7857, 16'd62003, 16'd62337, 16'd61221});
	test_expansion(128'h1b98a2ef96453ab0c9ae46857e7de815, {16'd40204, 16'd47821, 16'd63867, 16'd46938, 16'd63244, 16'd12298, 16'd36928, 16'd62200, 16'd38399, 16'd12999, 16'd61950, 16'd44160, 16'd65311, 16'd48105, 16'd716, 16'd53846, 16'd33814, 16'd16487, 16'd48138, 16'd3421, 16'd37730, 16'd24393, 16'd29579, 16'd1920, 16'd28494, 16'd12741});
	test_expansion(128'h5e91c4f5b4d043b095ad272c82f541a6, {16'd56912, 16'd14231, 16'd57536, 16'd27779, 16'd37361, 16'd17180, 16'd16764, 16'd41317, 16'd25021, 16'd58613, 16'd52127, 16'd21982, 16'd60220, 16'd42693, 16'd63119, 16'd19505, 16'd2606, 16'd37692, 16'd51277, 16'd38003, 16'd11666, 16'd61559, 16'd48953, 16'd11157, 16'd36239, 16'd32896});
	test_expansion(128'h2c3edbc948c454ccc0d2367f427f7d32, {16'd51656, 16'd47758, 16'd54769, 16'd61777, 16'd5288, 16'd21133, 16'd20530, 16'd50796, 16'd33019, 16'd63128, 16'd31265, 16'd58598, 16'd35708, 16'd30696, 16'd23811, 16'd3806, 16'd42321, 16'd60890, 16'd1847, 16'd40357, 16'd58061, 16'd5067, 16'd51944, 16'd25142, 16'd876, 16'd54131});
	test_expansion(128'he8e4dad71a54b26bc50013f24e28fce2, {16'd54676, 16'd22565, 16'd36939, 16'd47475, 16'd18437, 16'd45309, 16'd40756, 16'd15120, 16'd2409, 16'd42938, 16'd24901, 16'd5147, 16'd54311, 16'd27742, 16'd5293, 16'd5783, 16'd59789, 16'd7187, 16'd44167, 16'd60051, 16'd404, 16'd45925, 16'd52055, 16'd51547, 16'd31588, 16'd11844});
	test_expansion(128'h26d12c607cff4e4eaab792f40eb987db, {16'd32936, 16'd19811, 16'd63661, 16'd32737, 16'd11764, 16'd56346, 16'd47710, 16'd2418, 16'd13259, 16'd8893, 16'd2170, 16'd13601, 16'd50237, 16'd29085, 16'd580, 16'd7814, 16'd22677, 16'd57334, 16'd38922, 16'd23952, 16'd40059, 16'd42107, 16'd24671, 16'd65515, 16'd49239, 16'd57082});
	test_expansion(128'h822c7bed583e8d75bc956ad3a1d57a05, {16'd29491, 16'd35746, 16'd52427, 16'd61614, 16'd5241, 16'd41703, 16'd26797, 16'd33831, 16'd15308, 16'd2765, 16'd13403, 16'd11238, 16'd4904, 16'd28114, 16'd65366, 16'd28640, 16'd4438, 16'd58424, 16'd4483, 16'd44853, 16'd56618, 16'd25839, 16'd45565, 16'd43689, 16'd27590, 16'd44507});
	test_expansion(128'hbfd5537fd194b5e3aba09b9280bdca13, {16'd36832, 16'd21409, 16'd61417, 16'd44462, 16'd35342, 16'd33016, 16'd54649, 16'd52719, 16'd28506, 16'd45248, 16'd16743, 16'd9454, 16'd42018, 16'd16882, 16'd2581, 16'd43116, 16'd55801, 16'd18889, 16'd11587, 16'd62759, 16'd43248, 16'd11007, 16'd3367, 16'd60366, 16'd3773, 16'd58233});
	test_expansion(128'hff70567aa801c06bc3f8ef04637c0406, {16'd11030, 16'd37160, 16'd36197, 16'd21970, 16'd33587, 16'd1571, 16'd6650, 16'd4904, 16'd5633, 16'd12785, 16'd5526, 16'd17372, 16'd12541, 16'd21210, 16'd31797, 16'd62937, 16'd50925, 16'd39954, 16'd57474, 16'd46647, 16'd18989, 16'd32873, 16'd14734, 16'd38289, 16'd37764, 16'd31449});
	test_expansion(128'hb4f01e43b98a5f391b533b2f2fb2499e, {16'd55740, 16'd40472, 16'd53145, 16'd5111, 16'd857, 16'd23823, 16'd33722, 16'd5385, 16'd13568, 16'd20088, 16'd49724, 16'd7913, 16'd49391, 16'd42982, 16'd55916, 16'd60499, 16'd21043, 16'd21360, 16'd1894, 16'd51150, 16'd11493, 16'd22640, 16'd55642, 16'd27885, 16'd5677, 16'd970});
	test_expansion(128'hc327692d71576d6159002501bda23ddf, {16'd21518, 16'd31025, 16'd48800, 16'd64369, 16'd53196, 16'd51865, 16'd44389, 16'd6703, 16'd15142, 16'd22898, 16'd28762, 16'd39900, 16'd40796, 16'd50453, 16'd17313, 16'd61752, 16'd9328, 16'd60816, 16'd37155, 16'd28287, 16'd32392, 16'd18758, 16'd31525, 16'd54370, 16'd19378, 16'd40474});
	test_expansion(128'h95f15e326c847b723dd54756aaf3e2db, {16'd6158, 16'd2022, 16'd30304, 16'd23694, 16'd50061, 16'd34088, 16'd34554, 16'd40558, 16'd23950, 16'd18934, 16'd19720, 16'd3529, 16'd57052, 16'd23546, 16'd32177, 16'd63062, 16'd36592, 16'd17519, 16'd6413, 16'd22968, 16'd20509, 16'd38549, 16'd56268, 16'd46119, 16'd20745, 16'd57900});
	test_expansion(128'h7068d7fd8d1efe24be617178b1a1320c, {16'd35991, 16'd26527, 16'd50580, 16'd39001, 16'd62713, 16'd48693, 16'd29368, 16'd28387, 16'd46723, 16'd64590, 16'd23850, 16'd14863, 16'd24315, 16'd30464, 16'd61100, 16'd45935, 16'd64557, 16'd34691, 16'd9847, 16'd35609, 16'd62038, 16'd38692, 16'd15025, 16'd50838, 16'd25339, 16'd25368});
	test_expansion(128'hcb809b10ee81ccadf13a5cfcf21269bf, {16'd1298, 16'd59688, 16'd28003, 16'd55347, 16'd26232, 16'd51155, 16'd10592, 16'd58256, 16'd52058, 16'd18062, 16'd28667, 16'd26988, 16'd57154, 16'd37542, 16'd9419, 16'd26354, 16'd33750, 16'd14446, 16'd63250, 16'd55380, 16'd21186, 16'd51304, 16'd576, 16'd12875, 16'd60218, 16'd56726});
	test_expansion(128'he318c367aa3a36d6652b79d8e98076af, {16'd45416, 16'd27635, 16'd26027, 16'd45145, 16'd33186, 16'd29702, 16'd36378, 16'd59589, 16'd15179, 16'd54947, 16'd37466, 16'd28362, 16'd140, 16'd338, 16'd45357, 16'd47118, 16'd35062, 16'd1302, 16'd38074, 16'd41886, 16'd42103, 16'd55649, 16'd13529, 16'd52841, 16'd7957, 16'd54893});
	test_expansion(128'he82f1db76a2bd65f169cd3c94f849fec, {16'd24606, 16'd51908, 16'd37479, 16'd9, 16'd37954, 16'd55677, 16'd15008, 16'd32847, 16'd36618, 16'd24573, 16'd39060, 16'd9562, 16'd2096, 16'd18258, 16'd26287, 16'd3043, 16'd31427, 16'd13719, 16'd25384, 16'd45264, 16'd61191, 16'd981, 16'd28684, 16'd24469, 16'd20671, 16'd61504});
	test_expansion(128'h72744e520f466e1ab481ffcaccad90ca, {16'd51538, 16'd52349, 16'd50327, 16'd48146, 16'd44246, 16'd18869, 16'd42426, 16'd16585, 16'd25253, 16'd7113, 16'd38935, 16'd40245, 16'd46949, 16'd59998, 16'd15430, 16'd6780, 16'd53337, 16'd15158, 16'd12151, 16'd27061, 16'd14601, 16'd6125, 16'd26372, 16'd44730, 16'd22128, 16'd27342});
	test_expansion(128'h3f54ba5933f1382bb43a4a78c762cb86, {16'd8343, 16'd11534, 16'd8521, 16'd24617, 16'd15522, 16'd14217, 16'd65479, 16'd12122, 16'd37207, 16'd3373, 16'd62830, 16'd48060, 16'd22171, 16'd60153, 16'd56706, 16'd62422, 16'd36056, 16'd35796, 16'd38416, 16'd37583, 16'd58284, 16'd10386, 16'd2277, 16'd60331, 16'd47208, 16'd37533});
	test_expansion(128'h5425e83dbf7adca0506c07c32d575fda, {16'd12249, 16'd4018, 16'd57416, 16'd17484, 16'd28538, 16'd57835, 16'd23726, 16'd5191, 16'd7992, 16'd20269, 16'd19122, 16'd5592, 16'd59124, 16'd20009, 16'd61148, 16'd32710, 16'd34249, 16'd58873, 16'd151, 16'd24114, 16'd11913, 16'd38022, 16'd32663, 16'd56664, 16'd22437, 16'd45464});
	test_expansion(128'h98b4d223c4490ae6c1a5c589e570d068, {16'd42060, 16'd54733, 16'd46799, 16'd36431, 16'd36178, 16'd54038, 16'd44776, 16'd22856, 16'd48989, 16'd53637, 16'd58274, 16'd23459, 16'd8691, 16'd58927, 16'd30048, 16'd1411, 16'd5274, 16'd51101, 16'd9763, 16'd26571, 16'd45074, 16'd6460, 16'd6558, 16'd40372, 16'd8147, 16'd60123});
	test_expansion(128'h6080abc9c89f78335f3bc310378f1f3b, {16'd57056, 16'd61502, 16'd25899, 16'd62325, 16'd53199, 16'd59740, 16'd64397, 16'd16793, 16'd37334, 16'd42714, 16'd62317, 16'd46616, 16'd39418, 16'd24733, 16'd46398, 16'd37250, 16'd54107, 16'd24489, 16'd6096, 16'd25714, 16'd28571, 16'd4348, 16'd64825, 16'd42442, 16'd30812, 16'd6932});
	test_expansion(128'h1bc6b5f2046235cfdd88caebaec30b3d, {16'd15032, 16'd56568, 16'd48521, 16'd62118, 16'd34556, 16'd9124, 16'd24539, 16'd3948, 16'd22084, 16'd11371, 16'd4918, 16'd60489, 16'd25598, 16'd58616, 16'd17756, 16'd20171, 16'd33933, 16'd35581, 16'd36799, 16'd24609, 16'd41395, 16'd7469, 16'd55780, 16'd3911, 16'd3375, 16'd53250});
	test_expansion(128'h1d5632756daa2a0837a4de9020198924, {16'd42847, 16'd7276, 16'd43030, 16'd3384, 16'd2193, 16'd40306, 16'd33922, 16'd40944, 16'd9096, 16'd474, 16'd55833, 16'd45953, 16'd42575, 16'd47098, 16'd17290, 16'd51144, 16'd57499, 16'd48855, 16'd9251, 16'd5680, 16'd12342, 16'd55601, 16'd53304, 16'd6205, 16'd21075, 16'd6213});
	test_expansion(128'h4d5504477ac46025ee665d9c5be2e530, {16'd50920, 16'd17039, 16'd31469, 16'd14468, 16'd46331, 16'd62274, 16'd9073, 16'd19173, 16'd35262, 16'd31035, 16'd57376, 16'd36721, 16'd30004, 16'd31632, 16'd12856, 16'd1129, 16'd27498, 16'd2554, 16'd56701, 16'd44816, 16'd31956, 16'd13331, 16'd29249, 16'd27645, 16'd21268, 16'd35166});
	test_expansion(128'h857ef23a09cb9735ea5c4b53cfc75f8c, {16'd30163, 16'd23665, 16'd44098, 16'd60438, 16'd61607, 16'd16440, 16'd9410, 16'd48894, 16'd43723, 16'd3749, 16'd56015, 16'd22421, 16'd60306, 16'd8035, 16'd53320, 16'd42833, 16'd14048, 16'd190, 16'd50611, 16'd8112, 16'd57555, 16'd4005, 16'd39025, 16'd64636, 16'd5981, 16'd50483});
	test_expansion(128'h843d67f87c21283d16fe650bc6844bdd, {16'd48092, 16'd8173, 16'd57484, 16'd27467, 16'd40553, 16'd29293, 16'd25057, 16'd24262, 16'd3773, 16'd48159, 16'd90, 16'd45299, 16'd9513, 16'd36920, 16'd3444, 16'd1489, 16'd21044, 16'd57277, 16'd29817, 16'd53232, 16'd59282, 16'd29754, 16'd23607, 16'd24331, 16'd19592, 16'd60939});
	test_expansion(128'h5eafbe1661f6fb706bb710dd649ff2f5, {16'd27875, 16'd53315, 16'd44877, 16'd7186, 16'd18013, 16'd38632, 16'd55265, 16'd49847, 16'd49984, 16'd18111, 16'd21136, 16'd25316, 16'd33874, 16'd18565, 16'd16604, 16'd17424, 16'd22793, 16'd33500, 16'd43300, 16'd16078, 16'd20309, 16'd51705, 16'd6779, 16'd11807, 16'd6907, 16'd25129});
	test_expansion(128'h8e17d8e28f0e0000c95433030a9bf4b6, {16'd54713, 16'd45369, 16'd64908, 16'd17203, 16'd47724, 16'd45712, 16'd63096, 16'd39925, 16'd48877, 16'd55727, 16'd31971, 16'd39845, 16'd10722, 16'd23188, 16'd48507, 16'd29417, 16'd16758, 16'd15965, 16'd43225, 16'd49377, 16'd23085, 16'd53531, 16'd11738, 16'd22801, 16'd40464, 16'd48604});
	test_expansion(128'h6ffb00cf6708533d14d218f139c0e2df, {16'd24453, 16'd63123, 16'd63976, 16'd61612, 16'd18821, 16'd12833, 16'd3184, 16'd54822, 16'd2660, 16'd15242, 16'd9231, 16'd22812, 16'd54280, 16'd43512, 16'd37941, 16'd45926, 16'd20418, 16'd52581, 16'd58397, 16'd30614, 16'd13270, 16'd14475, 16'd46601, 16'd45840, 16'd43029, 16'd38895});
	test_expansion(128'h4b3c835c19168cc140504cb79b007e7a, {16'd32865, 16'd49911, 16'd55791, 16'd48181, 16'd46110, 16'd881, 16'd29544, 16'd20863, 16'd3220, 16'd20732, 16'd44819, 16'd47831, 16'd52260, 16'd34521, 16'd11106, 16'd36236, 16'd43236, 16'd48576, 16'd45769, 16'd16409, 16'd5354, 16'd62872, 16'd18059, 16'd60907, 16'd53867, 16'd63023});
	test_expansion(128'h6f0ccc913b3088ba7029265781dbff36, {16'd50022, 16'd21035, 16'd48750, 16'd10403, 16'd56462, 16'd12208, 16'd17062, 16'd41408, 16'd43535, 16'd38794, 16'd43870, 16'd15251, 16'd23324, 16'd2038, 16'd12402, 16'd54548, 16'd1216, 16'd47413, 16'd11154, 16'd42325, 16'd32345, 16'd7264, 16'd15471, 16'd48948, 16'd32476, 16'd42565});
	test_expansion(128'h62349a64e3f5e954b091ec1ddb7ef7d5, {16'd38146, 16'd30740, 16'd32234, 16'd26081, 16'd16771, 16'd35960, 16'd14463, 16'd23101, 16'd12723, 16'd42049, 16'd62550, 16'd30375, 16'd3943, 16'd33271, 16'd34069, 16'd25266, 16'd51040, 16'd27858, 16'd49009, 16'd27091, 16'd63202, 16'd2329, 16'd34336, 16'd58105, 16'd65271, 16'd48906});
	test_expansion(128'hdef99b63af47d3aa55317cf12060c647, {16'd53898, 16'd18806, 16'd28242, 16'd36722, 16'd60990, 16'd5853, 16'd3923, 16'd44897, 16'd46214, 16'd23345, 16'd22141, 16'd18277, 16'd34806, 16'd26220, 16'd21770, 16'd42093, 16'd5806, 16'd53780, 16'd38964, 16'd12434, 16'd57535, 16'd57980, 16'd24092, 16'd61858, 16'd61255, 16'd30136});
	test_expansion(128'h9d33fd0881e9d0f330baa504b9b21350, {16'd34057, 16'd24298, 16'd16566, 16'd47674, 16'd24293, 16'd21992, 16'd46062, 16'd51356, 16'd29675, 16'd31446, 16'd42469, 16'd6235, 16'd8446, 16'd64932, 16'd57538, 16'd60167, 16'd27258, 16'd16018, 16'd46813, 16'd40368, 16'd44410, 16'd26227, 16'd28728, 16'd52442, 16'd56357, 16'd8180});
	test_expansion(128'h1550e80f9d9295e9e64f08e622e7acd7, {16'd41027, 16'd31987, 16'd49684, 16'd36790, 16'd12144, 16'd31040, 16'd15870, 16'd6654, 16'd58839, 16'd48877, 16'd15930, 16'd17864, 16'd20433, 16'd37983, 16'd13389, 16'd40376, 16'd64479, 16'd39814, 16'd59272, 16'd10572, 16'd54188, 16'd48224, 16'd2068, 16'd14356, 16'd17834, 16'd60114});
	test_expansion(128'h9213aac8c5b3abecdbf7c46d135612f9, {16'd52467, 16'd23626, 16'd27869, 16'd13874, 16'd1402, 16'd12827, 16'd11358, 16'd17202, 16'd43768, 16'd5165, 16'd3259, 16'd13973, 16'd50423, 16'd60003, 16'd4409, 16'd21278, 16'd14610, 16'd48670, 16'd29409, 16'd27902, 16'd21511, 16'd17449, 16'd6505, 16'd31334, 16'd29678, 16'd20405});
	test_expansion(128'hf5bd84626f9077229a8e6fe8c5b2e704, {16'd65472, 16'd23001, 16'd43633, 16'd56936, 16'd34308, 16'd51330, 16'd48593, 16'd52725, 16'd13010, 16'd29679, 16'd65373, 16'd1367, 16'd9388, 16'd8617, 16'd4236, 16'd39467, 16'd26494, 16'd47755, 16'd59071, 16'd60907, 16'd3997, 16'd47210, 16'd40857, 16'd50993, 16'd20456, 16'd62203});
	test_expansion(128'h431fa7da63138c961340fc44907249f2, {16'd62628, 16'd57136, 16'd11207, 16'd59078, 16'd15363, 16'd22876, 16'd32774, 16'd35230, 16'd53365, 16'd27670, 16'd40683, 16'd40778, 16'd31981, 16'd61078, 16'd15346, 16'd30899, 16'd20397, 16'd5071, 16'd38298, 16'd9692, 16'd140, 16'd1590, 16'd15462, 16'd13032, 16'd8975, 16'd38083});
	test_expansion(128'h5b869d435e01ce93ee6933fc759f0e32, {16'd26619, 16'd60744, 16'd30222, 16'd50460, 16'd34405, 16'd27334, 16'd24587, 16'd45456, 16'd26687, 16'd38529, 16'd19339, 16'd32009, 16'd35982, 16'd52028, 16'd35950, 16'd10309, 16'd21396, 16'd28264, 16'd15716, 16'd64937, 16'd40697, 16'd49759, 16'd34231, 16'd47996, 16'd53784, 16'd26686});
	test_expansion(128'h31c4c196b2e54042e2c69f52c6bb54e0, {16'd25168, 16'd57262, 16'd22475, 16'd24977, 16'd12375, 16'd23624, 16'd13564, 16'd28312, 16'd15333, 16'd49483, 16'd30240, 16'd52994, 16'd19082, 16'd4860, 16'd12057, 16'd40343, 16'd780, 16'd42237, 16'd47632, 16'd16173, 16'd58741, 16'd64725, 16'd7187, 16'd50064, 16'd491, 16'd44409});
	test_expansion(128'hdd426dfb0e6d482cf4a80adc05594798, {16'd6103, 16'd62248, 16'd4040, 16'd54250, 16'd44642, 16'd10252, 16'd11535, 16'd20066, 16'd24203, 16'd24823, 16'd18012, 16'd19574, 16'd64474, 16'd30998, 16'd24750, 16'd21055, 16'd6488, 16'd56708, 16'd46129, 16'd34908, 16'd55674, 16'd54427, 16'd56329, 16'd56066, 16'd45589, 16'd46481});
	test_expansion(128'ha4793a5c98bc494a3b5044fe55a44fcb, {16'd23164, 16'd62235, 16'd6027, 16'd15939, 16'd60498, 16'd46442, 16'd44803, 16'd40597, 16'd10218, 16'd17645, 16'd64117, 16'd10981, 16'd61298, 16'd43708, 16'd40697, 16'd9400, 16'd8041, 16'd50624, 16'd9988, 16'd35670, 16'd34013, 16'd5508, 16'd6425, 16'd46135, 16'd16222, 16'd26993});
	test_expansion(128'h04b4569ffea62ed023f734ba64962c44, {16'd14797, 16'd13200, 16'd34865, 16'd53090, 16'd5397, 16'd16006, 16'd33710, 16'd46546, 16'd21830, 16'd12307, 16'd4992, 16'd14326, 16'd43719, 16'd17816, 16'd26395, 16'd33692, 16'd11919, 16'd29456, 16'd65357, 16'd50203, 16'd34816, 16'd47719, 16'd2946, 16'd27932, 16'd48154, 16'd33660});
	test_expansion(128'ha0c3f370e569b19bf2bd7e09dccd2dcb, {16'd63187, 16'd5721, 16'd21144, 16'd24441, 16'd36944, 16'd25017, 16'd48557, 16'd24797, 16'd58805, 16'd40121, 16'd43427, 16'd33370, 16'd48584, 16'd59806, 16'd28063, 16'd45577, 16'd51859, 16'd30045, 16'd1791, 16'd28065, 16'd10137, 16'd15202, 16'd44262, 16'd5215, 16'd31168, 16'd57119});
	test_expansion(128'h5d45f3884807ee24d0069227368d3a05, {16'd59116, 16'd17235, 16'd25330, 16'd31746, 16'd3762, 16'd31645, 16'd15564, 16'd52569, 16'd58301, 16'd22096, 16'd10627, 16'd24077, 16'd46256, 16'd23803, 16'd56721, 16'd32330, 16'd52078, 16'd31737, 16'd63267, 16'd64090, 16'd32360, 16'd14777, 16'd20948, 16'd6259, 16'd12184, 16'd18957});
	test_expansion(128'h4247d2d51637245d36ce32d23a2f8be3, {16'd33505, 16'd56105, 16'd23963, 16'd53152, 16'd52684, 16'd46202, 16'd42412, 16'd91, 16'd17750, 16'd3033, 16'd181, 16'd44653, 16'd33639, 16'd21572, 16'd12517, 16'd3792, 16'd1578, 16'd59206, 16'd41038, 16'd63903, 16'd1208, 16'd4625, 16'd37345, 16'd35628, 16'd13116, 16'd63127});
	test_expansion(128'h11e54b934edf82149edc89ab872b76b2, {16'd31185, 16'd34281, 16'd34117, 16'd58540, 16'd6244, 16'd17632, 16'd9326, 16'd28264, 16'd28909, 16'd49097, 16'd51146, 16'd41938, 16'd27152, 16'd58142, 16'd18199, 16'd40233, 16'd2972, 16'd21119, 16'd48277, 16'd48003, 16'd19571, 16'd29052, 16'd61434, 16'd65283, 16'd40416, 16'd52805});
	test_expansion(128'h0e57c5394c1e06009c76c02cf47bbe31, {16'd50374, 16'd63372, 16'd47188, 16'd16093, 16'd55031, 16'd5443, 16'd39223, 16'd34175, 16'd16250, 16'd4841, 16'd49230, 16'd54900, 16'd24670, 16'd5428, 16'd5628, 16'd19021, 16'd34396, 16'd19185, 16'd3821, 16'd59461, 16'd54868, 16'd38948, 16'd18102, 16'd46337, 16'd47937, 16'd48242});
	test_expansion(128'h3286d7b73ae53d7bff8762e5e782bfcb, {16'd35958, 16'd43768, 16'd21147, 16'd11668, 16'd16049, 16'd39980, 16'd60019, 16'd39168, 16'd44565, 16'd3601, 16'd9470, 16'd11089, 16'd28715, 16'd59574, 16'd17858, 16'd15467, 16'd28329, 16'd54999, 16'd6285, 16'd42475, 16'd32777, 16'd54544, 16'd14319, 16'd9109, 16'd64679, 16'd12318});
	test_expansion(128'hdceb70eae4f3455f64c9e3c4ec42889f, {16'd13517, 16'd29936, 16'd11809, 16'd11694, 16'd43791, 16'd42006, 16'd11826, 16'd57489, 16'd43774, 16'd57787, 16'd1531, 16'd44490, 16'd14596, 16'd63464, 16'd5458, 16'd5658, 16'd5662, 16'd46486, 16'd8199, 16'd55143, 16'd32579, 16'd34445, 16'd61696, 16'd58927, 16'd41259, 16'd55334});
	test_expansion(128'h6aaa35a80eb24243dbce4067ae76423f, {16'd22039, 16'd22918, 16'd3221, 16'd34474, 16'd3593, 16'd61335, 16'd5415, 16'd13260, 16'd65423, 16'd61507, 16'd26175, 16'd23773, 16'd27250, 16'd2548, 16'd39564, 16'd61827, 16'd61473, 16'd41257, 16'd41332, 16'd31048, 16'd596, 16'd27701, 16'd16216, 16'd57865, 16'd57390, 16'd32661});
	test_expansion(128'ha89cdf5f43a2b74e8f2c92222975b6c4, {16'd3349, 16'd33182, 16'd63438, 16'd55521, 16'd49483, 16'd52621, 16'd6203, 16'd6058, 16'd49815, 16'd37086, 16'd62196, 16'd37413, 16'd43886, 16'd30116, 16'd18564, 16'd4179, 16'd15555, 16'd61989, 16'd50709, 16'd28132, 16'd51283, 16'd53915, 16'd49510, 16'd24993, 16'd58731, 16'd56518});
	test_expansion(128'h82ddea2646bf6bee8f13b1e1943decb9, {16'd21565, 16'd5375, 16'd11081, 16'd18807, 16'd35440, 16'd62656, 16'd52950, 16'd28820, 16'd45097, 16'd9962, 16'd5294, 16'd38705, 16'd61875, 16'd8544, 16'd13547, 16'd13048, 16'd1325, 16'd14933, 16'd38412, 16'd54731, 16'd12144, 16'd17175, 16'd22772, 16'd32720, 16'd16022, 16'd10408});
	test_expansion(128'h159a215e1a9c41903285752f2b369d7c, {16'd6141, 16'd21244, 16'd40515, 16'd56988, 16'd60359, 16'd4521, 16'd4365, 16'd22093, 16'd13457, 16'd54709, 16'd24186, 16'd6412, 16'd44442, 16'd36384, 16'd21996, 16'd18218, 16'd61787, 16'd61784, 16'd39313, 16'd18043, 16'd36130, 16'd8059, 16'd56081, 16'd50885, 16'd14353, 16'd9807});
	test_expansion(128'hd2a2bc560b93991ac1cf14fe4f22d258, {16'd22730, 16'd11909, 16'd23392, 16'd62791, 16'd49456, 16'd61107, 16'd44153, 16'd40295, 16'd23054, 16'd3970, 16'd56159, 16'd22015, 16'd61392, 16'd44519, 16'd17466, 16'd4673, 16'd41048, 16'd14963, 16'd44614, 16'd15542, 16'd64956, 16'd51432, 16'd34453, 16'd7028, 16'd4744, 16'd43589});
	test_expansion(128'hb5a2355aca5380a3e840fb9844c16711, {16'd28762, 16'd49439, 16'd49295, 16'd44730, 16'd38936, 16'd23592, 16'd62442, 16'd42330, 16'd36264, 16'd17871, 16'd58635, 16'd14640, 16'd50993, 16'd16469, 16'd3547, 16'd48117, 16'd49217, 16'd21185, 16'd65177, 16'd3957, 16'd53695, 16'd57889, 16'd59594, 16'd14942, 16'd54881, 16'd42442});
	test_expansion(128'h4c1ab856a8aaac5356548d7023b57300, {16'd3047, 16'd28120, 16'd42801, 16'd41603, 16'd14987, 16'd47777, 16'd41626, 16'd30362, 16'd35036, 16'd64446, 16'd47013, 16'd4367, 16'd45062, 16'd30379, 16'd62521, 16'd52865, 16'd58923, 16'd34133, 16'd8185, 16'd49127, 16'd41623, 16'd30818, 16'd64786, 16'd57257, 16'd9967, 16'd27742});
	test_expansion(128'hda4ac2ac3043e33b8ac640c90efb69a2, {16'd17120, 16'd22899, 16'd30339, 16'd22348, 16'd64589, 16'd40144, 16'd34091, 16'd60780, 16'd22533, 16'd63057, 16'd20439, 16'd39251, 16'd47930, 16'd34754, 16'd55397, 16'd42540, 16'd21716, 16'd10076, 16'd32128, 16'd59032, 16'd26978, 16'd45642, 16'd3923, 16'd6579, 16'd22717, 16'd50266});
	test_expansion(128'h0e12b3b2d455641fcc986c8ed48717f3, {16'd55156, 16'd883, 16'd56405, 16'd55582, 16'd6159, 16'd23876, 16'd896, 16'd28345, 16'd31774, 16'd21867, 16'd40599, 16'd48775, 16'd2258, 16'd33620, 16'd10496, 16'd26833, 16'd14800, 16'd55487, 16'd14, 16'd42509, 16'd27655, 16'd21618, 16'd62291, 16'd47463, 16'd17007, 16'd6020});
	test_expansion(128'h10effb38ce5bbd955f13af81d8f627d7, {16'd31063, 16'd8241, 16'd55567, 16'd52277, 16'd9535, 16'd59057, 16'd59886, 16'd9226, 16'd55076, 16'd39555, 16'd33762, 16'd49246, 16'd21817, 16'd4607, 16'd60899, 16'd54715, 16'd9403, 16'd63172, 16'd5162, 16'd4743, 16'd21765, 16'd131, 16'd7690, 16'd14887, 16'd22037, 16'd40473});
	test_expansion(128'h9d18c437a8bfcdde9df14a4799fcaa6f, {16'd15132, 16'd18576, 16'd5510, 16'd62380, 16'd742, 16'd25610, 16'd58608, 16'd6769, 16'd11425, 16'd29629, 16'd62067, 16'd41465, 16'd7105, 16'd23792, 16'd7842, 16'd28020, 16'd65087, 16'd60495, 16'd56479, 16'd22935, 16'd64385, 16'd64615, 16'd4137, 16'd28740, 16'd2278, 16'd32311});
	test_expansion(128'h472e19664b35d2f384dd540b6c64959e, {16'd53804, 16'd11903, 16'd1014, 16'd21339, 16'd7129, 16'd44655, 16'd6537, 16'd29847, 16'd1130, 16'd40757, 16'd48958, 16'd2692, 16'd23506, 16'd45299, 16'd2632, 16'd31145, 16'd5573, 16'd36095, 16'd54502, 16'd45241, 16'd44026, 16'd38869, 16'd18210, 16'd28461, 16'd20741, 16'd51543});
	test_expansion(128'h7190efb241c88ee7b333c4bc92e654a9, {16'd25890, 16'd147, 16'd18248, 16'd28522, 16'd59966, 16'd27320, 16'd27966, 16'd39361, 16'd16815, 16'd16953, 16'd58736, 16'd28873, 16'd7877, 16'd31847, 16'd38987, 16'd34527, 16'd23282, 16'd5362, 16'd11264, 16'd3004, 16'd36879, 16'd22533, 16'd53386, 16'd30423, 16'd3747, 16'd40976});
	test_expansion(128'h18935f6eb1927c6e04137ef6161bbd82, {16'd35406, 16'd33336, 16'd16599, 16'd36802, 16'd12592, 16'd9880, 16'd978, 16'd41824, 16'd18378, 16'd63014, 16'd549, 16'd6289, 16'd28854, 16'd10441, 16'd12325, 16'd53673, 16'd20844, 16'd63042, 16'd39316, 16'd50079, 16'd24086, 16'd65186, 16'd26170, 16'd60906, 16'd10978, 16'd37093});
	test_expansion(128'h32232418b74fc6f6886cf9548bc0149a, {16'd32595, 16'd29256, 16'd21658, 16'd25185, 16'd18999, 16'd31050, 16'd3884, 16'd46157, 16'd19996, 16'd64735, 16'd31122, 16'd25701, 16'd59494, 16'd51465, 16'd6355, 16'd13681, 16'd800, 16'd52819, 16'd12534, 16'd41309, 16'd15462, 16'd7448, 16'd51869, 16'd30403, 16'd1485, 16'd58962});
	test_expansion(128'hb71545d16032356174aee97e11abd26f, {16'd55140, 16'd7631, 16'd44578, 16'd29582, 16'd23009, 16'd50820, 16'd14218, 16'd54250, 16'd3588, 16'd31453, 16'd33992, 16'd54543, 16'd64475, 16'd63855, 16'd35865, 16'd57358, 16'd63853, 16'd2743, 16'd4957, 16'd22502, 16'd51950, 16'd31409, 16'd14413, 16'd33433, 16'd43436, 16'd52607});
	test_expansion(128'h0025a4caca15d03883cfb6a4d32f1c52, {16'd15630, 16'd25978, 16'd23878, 16'd36017, 16'd10280, 16'd32268, 16'd6287, 16'd63753, 16'd32147, 16'd28169, 16'd50849, 16'd36081, 16'd62576, 16'd28513, 16'd55917, 16'd64371, 16'd59282, 16'd16297, 16'd33009, 16'd12972, 16'd41064, 16'd54947, 16'd19931, 16'd30972, 16'd39856, 16'd24303});
	test_expansion(128'h5631e0e089e2b35907d01b785b5db855, {16'd14333, 16'd37545, 16'd50681, 16'd36589, 16'd35596, 16'd18858, 16'd40682, 16'd2801, 16'd44940, 16'd33408, 16'd906, 16'd41232, 16'd45849, 16'd7832, 16'd17387, 16'd31136, 16'd21550, 16'd1617, 16'd27141, 16'd56049, 16'd23889, 16'd213, 16'd36526, 16'd18462, 16'd21288, 16'd21051});
	test_expansion(128'hf3ca5b0aa518116f36f635af00918932, {16'd41227, 16'd59287, 16'd62967, 16'd58871, 16'd64641, 16'd17540, 16'd11191, 16'd7781, 16'd48676, 16'd8885, 16'd30804, 16'd59785, 16'd10075, 16'd35854, 16'd32429, 16'd37271, 16'd26864, 16'd5131, 16'd61444, 16'd31829, 16'd45244, 16'd39294, 16'd45320, 16'd39941, 16'd38727, 16'd61862});
	test_expansion(128'h8a4a3c3c1d2ee513899a1a6614316cdc, {16'd18974, 16'd33523, 16'd60453, 16'd1198, 16'd46032, 16'd47008, 16'd44927, 16'd52580, 16'd30779, 16'd32351, 16'd8067, 16'd61003, 16'd34898, 16'd24787, 16'd38525, 16'd33992, 16'd46603, 16'd23201, 16'd46032, 16'd4966, 16'd48997, 16'd31338, 16'd28017, 16'd5120, 16'd44269, 16'd27918});
	test_expansion(128'h62eb7b9c88cd44c339b59d4f578cff85, {16'd52550, 16'd16406, 16'd23654, 16'd16789, 16'd53344, 16'd57862, 16'd48717, 16'd18089, 16'd42008, 16'd10283, 16'd21118, 16'd2265, 16'd3758, 16'd63730, 16'd27841, 16'd41663, 16'd8801, 16'd32346, 16'd17256, 16'd56751, 16'd57622, 16'd28366, 16'd46963, 16'd20712, 16'd48499, 16'd23996});
	test_expansion(128'hb464e08793c6805049734e1a53fba009, {16'd18182, 16'd17219, 16'd53137, 16'd49188, 16'd20239, 16'd47117, 16'd9414, 16'd14899, 16'd45454, 16'd43863, 16'd33054, 16'd26911, 16'd31167, 16'd19606, 16'd5843, 16'd56858, 16'd17688, 16'd31213, 16'd50781, 16'd52591, 16'd43080, 16'd45448, 16'd31362, 16'd36223, 16'd22909, 16'd28561});
	test_expansion(128'h1cbe761515c70e9774683f755e577467, {16'd22798, 16'd51881, 16'd56469, 16'd50016, 16'd47811, 16'd17098, 16'd39552, 16'd45908, 16'd51041, 16'd56864, 16'd64892, 16'd13358, 16'd55050, 16'd63509, 16'd23990, 16'd10090, 16'd51280, 16'd23086, 16'd27679, 16'd9555, 16'd59834, 16'd39475, 16'd43167, 16'd22884, 16'd48833, 16'd22294});
	test_expansion(128'h2d7ff7c0b387ec9f8163bbd73c962192, {16'd48154, 16'd13379, 16'd2606, 16'd51395, 16'd51781, 16'd2732, 16'd30444, 16'd61946, 16'd16360, 16'd65069, 16'd6835, 16'd52395, 16'd29017, 16'd37843, 16'd10199, 16'd35307, 16'd22262, 16'd28005, 16'd22126, 16'd7268, 16'd47905, 16'd235, 16'd25720, 16'd58040, 16'd5000, 16'd31946});
	test_expansion(128'h453af873db46f9cf442d859c702261ea, {16'd41913, 16'd51485, 16'd60638, 16'd11850, 16'd42092, 16'd8649, 16'd6929, 16'd56652, 16'd48309, 16'd7592, 16'd42802, 16'd53136, 16'd41719, 16'd4406, 16'd22863, 16'd65376, 16'd44794, 16'd17736, 16'd44522, 16'd16513, 16'd15474, 16'd34993, 16'd64211, 16'd60026, 16'd39060, 16'd37283});
	test_expansion(128'haa6531719000abb4a2f2980008aef992, {16'd26459, 16'd57622, 16'd40841, 16'd59035, 16'd6092, 16'd6720, 16'd47250, 16'd23726, 16'd12319, 16'd33237, 16'd52642, 16'd29718, 16'd20565, 16'd14782, 16'd7930, 16'd12266, 16'd43827, 16'd58595, 16'd7833, 16'd12746, 16'd29421, 16'd53672, 16'd42855, 16'd2215, 16'd8307, 16'd42691});
	test_expansion(128'hd7ad2f5e8970df3fd38c1e02b62349e2, {16'd41637, 16'd404, 16'd63978, 16'd44982, 16'd32508, 16'd11649, 16'd27064, 16'd61211, 16'd11647, 16'd55268, 16'd13127, 16'd14256, 16'd12654, 16'd28121, 16'd46439, 16'd27892, 16'd9672, 16'd38089, 16'd28683, 16'd44649, 16'd1881, 16'd51142, 16'd43492, 16'd15487, 16'd3682, 16'd56297});
	test_expansion(128'h8739629d3a966fad109a57ab8b308ee0, {16'd27859, 16'd28590, 16'd53308, 16'd63125, 16'd46322, 16'd26281, 16'd65323, 16'd22467, 16'd32006, 16'd62199, 16'd58502, 16'd36738, 16'd45067, 16'd25462, 16'd45999, 16'd41297, 16'd60595, 16'd44519, 16'd26939, 16'd4172, 16'd37154, 16'd7698, 16'd44912, 16'd58598, 16'd58214, 16'd52796});
	test_expansion(128'he3a429acfc667bd2dbc24586312a1af9, {16'd50567, 16'd20719, 16'd44840, 16'd9591, 16'd11808, 16'd8174, 16'd12323, 16'd41842, 16'd1008, 16'd50934, 16'd16315, 16'd57938, 16'd22365, 16'd44351, 16'd43490, 16'd48522, 16'd64101, 16'd1934, 16'd1656, 16'd63220, 16'd57137, 16'd59731, 16'd59929, 16'd18737, 16'd26521, 16'd48647});
	test_expansion(128'h50c8056fca87cbdcff4f16b51c14b946, {16'd280, 16'd27797, 16'd910, 16'd52348, 16'd42752, 16'd22795, 16'd52370, 16'd54351, 16'd50855, 16'd28614, 16'd3279, 16'd27880, 16'd49484, 16'd50058, 16'd34722, 16'd47892, 16'd37132, 16'd14905, 16'd49901, 16'd22007, 16'd24792, 16'd14803, 16'd18723, 16'd2129, 16'd45500, 16'd12996});
	test_expansion(128'h8525344a1cfb40499708ed198e9136b9, {16'd2778, 16'd65121, 16'd11961, 16'd17021, 16'd4382, 16'd22207, 16'd14195, 16'd27783, 16'd18809, 16'd24417, 16'd30445, 16'd13908, 16'd55878, 16'd16950, 16'd21316, 16'd11072, 16'd15244, 16'd55542, 16'd11577, 16'd5029, 16'd28429, 16'd27, 16'd29152, 16'd21975, 16'd48041, 16'd365});
	test_expansion(128'ha7187ac8850a25782d0c39732d54e2e7, {16'd38376, 16'd48121, 16'd61693, 16'd31151, 16'd16748, 16'd39615, 16'd28393, 16'd7384, 16'd17526, 16'd5709, 16'd41619, 16'd14817, 16'd37554, 16'd17998, 16'd42589, 16'd3893, 16'd14560, 16'd12795, 16'd1458, 16'd53868, 16'd33440, 16'd4305, 16'd41195, 16'd43628, 16'd43133, 16'd25396});
	test_expansion(128'hc831dcd28d48ca3e2bea13baf82e9fdf, {16'd24724, 16'd14764, 16'd1247, 16'd38729, 16'd14809, 16'd1082, 16'd43838, 16'd46279, 16'd29995, 16'd9797, 16'd54424, 16'd25167, 16'd37144, 16'd60193, 16'd64942, 16'd45490, 16'd57677, 16'd44907, 16'd65406, 16'd63306, 16'd22665, 16'd2600, 16'd17848, 16'd46392, 16'd20009, 16'd2319});
	test_expansion(128'h3edf383abc3dbcd447ea369ee6401aec, {16'd65505, 16'd1239, 16'd44602, 16'd35367, 16'd21482, 16'd52905, 16'd50306, 16'd58014, 16'd28387, 16'd57324, 16'd39607, 16'd1435, 16'd61739, 16'd58647, 16'd45325, 16'd21791, 16'd2285, 16'd40466, 16'd7680, 16'd57537, 16'd3802, 16'd33652, 16'd37143, 16'd22969, 16'd37833, 16'd23529});
	test_expansion(128'he95ef705b5f8efc70408504f9687d6c9, {16'd979, 16'd35648, 16'd29496, 16'd2975, 16'd30316, 16'd25895, 16'd27738, 16'd38892, 16'd13501, 16'd37873, 16'd15124, 16'd27649, 16'd53512, 16'd46555, 16'd28492, 16'd9583, 16'd43061, 16'd29178, 16'd12305, 16'd18890, 16'd28868, 16'd37184, 16'd10283, 16'd15631, 16'd57321, 16'd21775});
	test_expansion(128'h828011c17174d3adcda79da4f5368687, {16'd49101, 16'd11025, 16'd40232, 16'd43570, 16'd16873, 16'd31587, 16'd41999, 16'd49056, 16'd52981, 16'd19972, 16'd3694, 16'd6665, 16'd2535, 16'd46114, 16'd1518, 16'd42645, 16'd46902, 16'd63746, 16'd50024, 16'd30394, 16'd27973, 16'd57097, 16'd61188, 16'd32862, 16'd54647, 16'd23756});
	test_expansion(128'hbfe30a7d2f196d3ab161174ea261fbc2, {16'd50437, 16'd53857, 16'd57958, 16'd35329, 16'd50039, 16'd46932, 16'd20676, 16'd4174, 16'd24431, 16'd64346, 16'd38005, 16'd14046, 16'd19257, 16'd37977, 16'd38446, 16'd12109, 16'd18096, 16'd2863, 16'd8148, 16'd51970, 16'd48760, 16'd20932, 16'd35150, 16'd51328, 16'd54870, 16'd46756});
	test_expansion(128'h65ec946994f39983a536ea35e0973622, {16'd54037, 16'd9587, 16'd62211, 16'd18548, 16'd43729, 16'd10144, 16'd38058, 16'd25003, 16'd47785, 16'd54868, 16'd51293, 16'd46439, 16'd34458, 16'd44566, 16'd25764, 16'd45882, 16'd31515, 16'd10085, 16'd34677, 16'd64124, 16'd55167, 16'd45290, 16'd5687, 16'd20684, 16'd33866, 16'd41233});
	test_expansion(128'h805970dca4bf7fded9a42a9219f7795c, {16'd58924, 16'd26504, 16'd56933, 16'd39183, 16'd342, 16'd63526, 16'd29679, 16'd7953, 16'd8161, 16'd20953, 16'd4397, 16'd50074, 16'd51766, 16'd62649, 16'd25204, 16'd325, 16'd8498, 16'd19611, 16'd31574, 16'd55371, 16'd17853, 16'd45154, 16'd34167, 16'd6059, 16'd33699, 16'd6025});
	test_expansion(128'h3d7471fb16f7ddf49fcc2c71ad4690a4, {16'd630, 16'd61396, 16'd61313, 16'd53934, 16'd49042, 16'd49469, 16'd45715, 16'd7330, 16'd49294, 16'd9513, 16'd50932, 16'd61276, 16'd46380, 16'd20646, 16'd21025, 16'd29015, 16'd44940, 16'd24392, 16'd50794, 16'd44619, 16'd20961, 16'd22925, 16'd56857, 16'd57984, 16'd60557, 16'd49459});
	test_expansion(128'h03c149a0cc2e5515668e1ddcae42bf58, {16'd63908, 16'd61169, 16'd43593, 16'd3663, 16'd28135, 16'd44255, 16'd30069, 16'd41752, 16'd33723, 16'd41955, 16'd53162, 16'd14178, 16'd29300, 16'd14755, 16'd48590, 16'd22852, 16'd4245, 16'd26755, 16'd60973, 16'd26972, 16'd29663, 16'd62347, 16'd9173, 16'd58608, 16'd21751, 16'd17496});
	test_expansion(128'hde2327e0e6b050415b88f0a54cb6529b, {16'd42666, 16'd4909, 16'd51738, 16'd40449, 16'd42329, 16'd39028, 16'd13813, 16'd17853, 16'd6000, 16'd621, 16'd40106, 16'd28063, 16'd3617, 16'd41662, 16'd26424, 16'd40049, 16'd8920, 16'd1282, 16'd41004, 16'd6744, 16'd23627, 16'd24590, 16'd61042, 16'd1548, 16'd43120, 16'd19712});
	test_expansion(128'h1d1d0cbacc6ec7044ff4a143d0f37b83, {16'd47704, 16'd65210, 16'd43806, 16'd44019, 16'd62541, 16'd45800, 16'd2544, 16'd8110, 16'd4805, 16'd62132, 16'd23794, 16'd29880, 16'd7640, 16'd37286, 16'd24080, 16'd9437, 16'd27535, 16'd35332, 16'd47190, 16'd21129, 16'd40097, 16'd18706, 16'd56956, 16'd30827, 16'd6522, 16'd11857});
	test_expansion(128'hd12c018770f74337921345e1cc0e1a7e, {16'd62876, 16'd32558, 16'd34605, 16'd11310, 16'd59012, 16'd46124, 16'd8878, 16'd14294, 16'd13062, 16'd20731, 16'd16717, 16'd61634, 16'd42513, 16'd61714, 16'd649, 16'd26861, 16'd19705, 16'd1275, 16'd1223, 16'd18960, 16'd62173, 16'd33687, 16'd56233, 16'd50598, 16'd25785, 16'd61737});
	test_expansion(128'hb0404d89bd0aba235b6acc0976a71e35, {16'd48950, 16'd44745, 16'd30072, 16'd24662, 16'd4922, 16'd57527, 16'd2788, 16'd12172, 16'd63079, 16'd65479, 16'd28402, 16'd48321, 16'd61617, 16'd52073, 16'd52866, 16'd2555, 16'd41499, 16'd15347, 16'd32765, 16'd34449, 16'd50533, 16'd23738, 16'd63635, 16'd33158, 16'd30714, 16'd44523});
	test_expansion(128'h155a7fad0cca4bcdff9796ed4ca41be2, {16'd41198, 16'd60514, 16'd33653, 16'd21610, 16'd5569, 16'd44287, 16'd5467, 16'd61217, 16'd25735, 16'd976, 16'd44265, 16'd7396, 16'd34895, 16'd2521, 16'd63269, 16'd63949, 16'd1740, 16'd20738, 16'd30563, 16'd25061, 16'd27321, 16'd56682, 16'd49729, 16'd24514, 16'd20256, 16'd8818});
	test_expansion(128'he93ad8cafb0aede52563376f1b7f4040, {16'd57540, 16'd62948, 16'd31655, 16'd62529, 16'd43705, 16'd62333, 16'd57091, 16'd25181, 16'd2932, 16'd1160, 16'd53355, 16'd14879, 16'd54344, 16'd62537, 16'd3604, 16'd56933, 16'd61989, 16'd10266, 16'd29950, 16'd32440, 16'd48056, 16'd173, 16'd46789, 16'd15490, 16'd31229, 16'd26999});
	test_expansion(128'he8ccc158e21efbbbbf5802ff257b92d6, {16'd12579, 16'd63995, 16'd5134, 16'd19108, 16'd16172, 16'd36748, 16'd63109, 16'd10182, 16'd13908, 16'd37287, 16'd620, 16'd41050, 16'd20159, 16'd15499, 16'd63949, 16'd14297, 16'd48519, 16'd48092, 16'd7790, 16'd45315, 16'd61340, 16'd46865, 16'd58919, 16'd32364, 16'd58755, 16'd8395});
	test_expansion(128'h6fcd3408294ba4aee6fe492f11ecc93f, {16'd58565, 16'd15008, 16'd57122, 16'd60047, 16'd33908, 16'd60564, 16'd37901, 16'd13815, 16'd33971, 16'd10501, 16'd45074, 16'd58778, 16'd15289, 16'd38709, 16'd3364, 16'd7717, 16'd63284, 16'd14957, 16'd47496, 16'd53867, 16'd37486, 16'd4106, 16'd13312, 16'd23180, 16'd5798, 16'd44887});
	test_expansion(128'hc7e97c1987ac190fdf256e59a74343d5, {16'd50267, 16'd54786, 16'd4136, 16'd212, 16'd306, 16'd49003, 16'd6831, 16'd14566, 16'd25188, 16'd14241, 16'd29779, 16'd30968, 16'd18320, 16'd62314, 16'd2555, 16'd37860, 16'd53281, 16'd49749, 16'd119, 16'd39295, 16'd6778, 16'd57829, 16'd30686, 16'd62828, 16'd29896, 16'd3654});
	test_expansion(128'h6a9e289a6ec435f07de2172ad9cadbf1, {16'd29590, 16'd28080, 16'd59045, 16'd64330, 16'd50698, 16'd10440, 16'd58047, 16'd9427, 16'd14336, 16'd60127, 16'd26416, 16'd30696, 16'd7546, 16'd12555, 16'd15666, 16'd11037, 16'd21753, 16'd56559, 16'd31197, 16'd44555, 16'd28319, 16'd41857, 16'd47925, 16'd28429, 16'd17972, 16'd25921});
	test_expansion(128'hf2dd31569f679f7453b57491a101f2f2, {16'd21515, 16'd11511, 16'd27265, 16'd32744, 16'd23372, 16'd21784, 16'd62564, 16'd35708, 16'd18533, 16'd28047, 16'd38763, 16'd37467, 16'd25075, 16'd55493, 16'd19879, 16'd8815, 16'd17570, 16'd58022, 16'd9464, 16'd56679, 16'd47963, 16'd16434, 16'd35777, 16'd6281, 16'd54956, 16'd51050});
	test_expansion(128'hecf4994098dec1523def29e624ba6d94, {16'd6701, 16'd53298, 16'd3954, 16'd26517, 16'd30082, 16'd27172, 16'd45425, 16'd34298, 16'd33062, 16'd39489, 16'd6413, 16'd57837, 16'd32231, 16'd22152, 16'd45428, 16'd38288, 16'd7431, 16'd29403, 16'd24598, 16'd23668, 16'd34817, 16'd16754, 16'd19182, 16'd38083, 16'd7105, 16'd21685});
	test_expansion(128'h2619964672fa31c732f712689a41b09a, {16'd14791, 16'd30619, 16'd981, 16'd12947, 16'd32926, 16'd23416, 16'd13843, 16'd27698, 16'd14446, 16'd4789, 16'd2347, 16'd7018, 16'd30382, 16'd61826, 16'd31824, 16'd51233, 16'd25030, 16'd23051, 16'd28036, 16'd13095, 16'd29648, 16'd7831, 16'd15562, 16'd53446, 16'd27862, 16'd48721});
	test_expansion(128'h284d3a4cc21439264703121b69f5f22f, {16'd1141, 16'd4573, 16'd36732, 16'd3466, 16'd51356, 16'd4436, 16'd3956, 16'd19006, 16'd20213, 16'd32709, 16'd2937, 16'd22701, 16'd13672, 16'd36790, 16'd25293, 16'd42212, 16'd21301, 16'd5994, 16'd27847, 16'd59346, 16'd3714, 16'd19197, 16'd59048, 16'd29634, 16'd6534, 16'd11599});
	test_expansion(128'h8c0aee4f15a288ba93de396fc33a832e, {16'd8521, 16'd47583, 16'd55035, 16'd28830, 16'd44521, 16'd3980, 16'd46766, 16'd58173, 16'd40679, 16'd43868, 16'd40595, 16'd49136, 16'd61431, 16'd7577, 16'd5200, 16'd61565, 16'd8303, 16'd17988, 16'd21589, 16'd56890, 16'd6477, 16'd7420, 16'd29015, 16'd760, 16'd23084, 16'd46658});
	test_expansion(128'hff136d934d2fe6a4577d72a29fbdecf1, {16'd43271, 16'd12679, 16'd32976, 16'd7160, 16'd60932, 16'd35780, 16'd1222, 16'd9954, 16'd42189, 16'd11411, 16'd16298, 16'd34004, 16'd58211, 16'd55265, 16'd52378, 16'd51312, 16'd61281, 16'd26167, 16'd15769, 16'd43236, 16'd11307, 16'd63992, 16'd8472, 16'd25075, 16'd23346, 16'd49496});
	test_expansion(128'h32408ce733a10479b32e767012a23141, {16'd26833, 16'd9623, 16'd50037, 16'd27893, 16'd45695, 16'd25994, 16'd51834, 16'd63287, 16'd45946, 16'd27343, 16'd13065, 16'd42191, 16'd18685, 16'd54168, 16'd30808, 16'd43166, 16'd20710, 16'd42423, 16'd28813, 16'd40765, 16'd9696, 16'd11010, 16'd35248, 16'd21097, 16'd20346, 16'd5479});
	test_expansion(128'h2f6ec862aeb55656c816794c828844a8, {16'd21854, 16'd40832, 16'd26780, 16'd37789, 16'd54625, 16'd44509, 16'd41147, 16'd8666, 16'd47109, 16'd61972, 16'd63039, 16'd1341, 16'd8007, 16'd31601, 16'd17430, 16'd3403, 16'd29485, 16'd18500, 16'd2351, 16'd45479, 16'd1860, 16'd38225, 16'd37208, 16'd37104, 16'd26075, 16'd53925});
	test_expansion(128'h91c091e1929f6c2b79afbf15bb2899fc, {16'd27835, 16'd16912, 16'd19812, 16'd2285, 16'd38064, 16'd24022, 16'd10302, 16'd8030, 16'd17191, 16'd26314, 16'd15933, 16'd5685, 16'd12970, 16'd31703, 16'd28094, 16'd32767, 16'd2793, 16'd35842, 16'd2722, 16'd20805, 16'd34695, 16'd62142, 16'd17337, 16'd32386, 16'd50056, 16'd60302});
	test_expansion(128'h011beb2fb4d8e4d2f633af2baf0b6714, {16'd23505, 16'd58967, 16'd37335, 16'd25926, 16'd63001, 16'd63072, 16'd24369, 16'd41938, 16'd56308, 16'd62405, 16'd32715, 16'd27869, 16'd41457, 16'd10057, 16'd48390, 16'd64439, 16'd52164, 16'd24983, 16'd3435, 16'd36313, 16'd47465, 16'd60449, 16'd28715, 16'd34158, 16'd31337, 16'd61865});
	test_expansion(128'h397ba7ecc1a21fef11219105d47dea87, {16'd12734, 16'd26050, 16'd33219, 16'd2766, 16'd22765, 16'd18247, 16'd19130, 16'd32068, 16'd34376, 16'd35426, 16'd58312, 16'd60562, 16'd21317, 16'd13697, 16'd36074, 16'd57197, 16'd38955, 16'd35094, 16'd17117, 16'd60320, 16'd31202, 16'd4980, 16'd23390, 16'd62612, 16'd26970, 16'd12363});
	test_expansion(128'hbf852863c9148f2ad384b742ae4d3630, {16'd49257, 16'd974, 16'd16030, 16'd14969, 16'd26541, 16'd55970, 16'd7073, 16'd13486, 16'd8594, 16'd55956, 16'd3313, 16'd20183, 16'd57811, 16'd61910, 16'd65044, 16'd62, 16'd24757, 16'd62019, 16'd2677, 16'd1382, 16'd32894, 16'd65080, 16'd33634, 16'd45599, 16'd36099, 16'd51598});
	test_expansion(128'h843bba45858e792828856271410b45a6, {16'd22320, 16'd62988, 16'd8579, 16'd17955, 16'd7128, 16'd25237, 16'd57878, 16'd39651, 16'd39630, 16'd16010, 16'd29822, 16'd21398, 16'd3583, 16'd50258, 16'd32441, 16'd23618, 16'd36973, 16'd10888, 16'd34640, 16'd27204, 16'd12970, 16'd25445, 16'd63493, 16'd11285, 16'd1363, 16'd28524});
	test_expansion(128'h9a4c09c9f20401b45bc3e51b9deb0e07, {16'd59893, 16'd6407, 16'd8569, 16'd25318, 16'd30402, 16'd31150, 16'd33222, 16'd24404, 16'd31665, 16'd55973, 16'd36375, 16'd52419, 16'd48416, 16'd49974, 16'd3744, 16'd15708, 16'd57478, 16'd12281, 16'd56043, 16'd15970, 16'd37509, 16'd65182, 16'd33638, 16'd5370, 16'd16364, 16'd48411});
	test_expansion(128'heb324f01c55af14c1abb7abd2c1cb2f2, {16'd19107, 16'd16906, 16'd38192, 16'd56604, 16'd46517, 16'd3271, 16'd42981, 16'd28203, 16'd7560, 16'd34094, 16'd24275, 16'd17200, 16'd37673, 16'd45931, 16'd49345, 16'd26530, 16'd60120, 16'd34417, 16'd30172, 16'd40866, 16'd27332, 16'd26796, 16'd9931, 16'd45195, 16'd16099, 16'd62008});
	test_expansion(128'hc4b3f46d5833e200e37f9f68451d35e4, {16'd44126, 16'd38918, 16'd47086, 16'd64961, 16'd4461, 16'd41444, 16'd4984, 16'd12652, 16'd1867, 16'd63013, 16'd39961, 16'd55179, 16'd35779, 16'd19133, 16'd22775, 16'd50010, 16'd14153, 16'd39326, 16'd1931, 16'd25132, 16'd21232, 16'd42129, 16'd5040, 16'd38890, 16'd29719, 16'd22468});
	test_expansion(128'hcd99e744875acdfb0abaf52ce09d349f, {16'd13267, 16'd37134, 16'd55655, 16'd61898, 16'd22568, 16'd64302, 16'd22750, 16'd30834, 16'd58383, 16'd12299, 16'd63446, 16'd38042, 16'd60243, 16'd57302, 16'd5787, 16'd20131, 16'd25298, 16'd62022, 16'd18053, 16'd34132, 16'd43512, 16'd56908, 16'd32684, 16'd13200, 16'd59369, 16'd14495});
	test_expansion(128'h44772d4b72ee6000e6c9041aff8e9111, {16'd9776, 16'd34419, 16'd4905, 16'd56194, 16'd5092, 16'd11915, 16'd56901, 16'd53997, 16'd58261, 16'd10094, 16'd65360, 16'd34195, 16'd4509, 16'd31063, 16'd30610, 16'd14661, 16'd22398, 16'd3088, 16'd9288, 16'd31078, 16'd34429, 16'd53908, 16'd5597, 16'd37521, 16'd26879, 16'd2115});
	test_expansion(128'h532099c91764f4f6b6a8425c6919b20e, {16'd29729, 16'd59719, 16'd34238, 16'd253, 16'd62638, 16'd22027, 16'd16718, 16'd9078, 16'd24236, 16'd12338, 16'd24688, 16'd50368, 16'd62166, 16'd52395, 16'd31477, 16'd46157, 16'd31879, 16'd47175, 16'd8757, 16'd37486, 16'd27534, 16'd49744, 16'd34267, 16'd8260, 16'd50033, 16'd2050});
	test_expansion(128'h518540d417365525bbee9de591ff9d71, {16'd4113, 16'd22498, 16'd26824, 16'd24638, 16'd3327, 16'd25976, 16'd47059, 16'd14419, 16'd38653, 16'd58748, 16'd47555, 16'd27771, 16'd5565, 16'd5390, 16'd25872, 16'd59091, 16'd5194, 16'd46628, 16'd56596, 16'd33877, 16'd44774, 16'd64697, 16'd3422, 16'd36962, 16'd53516, 16'd2309});
	test_expansion(128'h830e37efa9b11b4d8197cbc6bd31b55a, {16'd50801, 16'd62853, 16'd21782, 16'd54598, 16'd24310, 16'd24442, 16'd48065, 16'd7482, 16'd9432, 16'd49159, 16'd4682, 16'd25175, 16'd1334, 16'd49218, 16'd53012, 16'd31650, 16'd31717, 16'd61238, 16'd20800, 16'd30250, 16'd9487, 16'd28930, 16'd55109, 16'd22517, 16'd26258, 16'd17414});
	test_expansion(128'h20be6a443c1bcaa55903a4b94d2f5bcd, {16'd34062, 16'd45054, 16'd24070, 16'd45815, 16'd59960, 16'd50304, 16'd38805, 16'd25226, 16'd28479, 16'd36427, 16'd20276, 16'd15579, 16'd37583, 16'd34499, 16'd51975, 16'd31927, 16'd43439, 16'd19306, 16'd24941, 16'd60880, 16'd31363, 16'd2561, 16'd783, 16'd15700, 16'd28764, 16'd49916});
	test_expansion(128'hd1e3a812e0b0fb437b3c77bcda220691, {16'd52239, 16'd54766, 16'd20417, 16'd39942, 16'd44726, 16'd43563, 16'd942, 16'd8896, 16'd17738, 16'd26279, 16'd32265, 16'd23492, 16'd2703, 16'd56076, 16'd14253, 16'd18793, 16'd26624, 16'd20917, 16'd49023, 16'd57368, 16'd50225, 16'd64455, 16'd26528, 16'd11929, 16'd46921, 16'd34122});
	test_expansion(128'hd6e2451c11e1543bd1b85e425d2533cd, {16'd21288, 16'd39681, 16'd31386, 16'd26588, 16'd2674, 16'd52269, 16'd13760, 16'd26999, 16'd46102, 16'd1102, 16'd63569, 16'd15543, 16'd25656, 16'd28848, 16'd9256, 16'd4757, 16'd44967, 16'd6220, 16'd51814, 16'd12521, 16'd59669, 16'd2331, 16'd42943, 16'd59158, 16'd54434, 16'd53750});
	test_expansion(128'h63905d25855f5bbc294aa0de41f2377e, {16'd24907, 16'd46247, 16'd62693, 16'd63161, 16'd36630, 16'd18189, 16'd20281, 16'd53617, 16'd55879, 16'd29555, 16'd6878, 16'd57798, 16'd6670, 16'd30261, 16'd7225, 16'd28921, 16'd37993, 16'd62764, 16'd14858, 16'd6937, 16'd44269, 16'd26456, 16'd18715, 16'd29716, 16'd39210, 16'd46665});
	test_expansion(128'h3c941304b4484ef4b11fb44350e4e489, {16'd36973, 16'd17854, 16'd55484, 16'd18366, 16'd31765, 16'd32720, 16'd16724, 16'd18929, 16'd30980, 16'd1777, 16'd19042, 16'd28931, 16'd11036, 16'd25488, 16'd35543, 16'd46084, 16'd42656, 16'd1565, 16'd42863, 16'd64637, 16'd12642, 16'd6572, 16'd23290, 16'd23610, 16'd42917, 16'd6935});
	test_expansion(128'h169f8a5058e3f6ab5829a9377ea38b07, {16'd21034, 16'd55440, 16'd37404, 16'd44912, 16'd61790, 16'd5300, 16'd43812, 16'd49651, 16'd51649, 16'd37648, 16'd28528, 16'd56661, 16'd54847, 16'd65346, 16'd55617, 16'd29665, 16'd23686, 16'd22393, 16'd19334, 16'd12585, 16'd32419, 16'd24513, 16'd12914, 16'd48893, 16'd25285, 16'd8877});
	test_expansion(128'h7ad4d7964ec4d08e8607cafd20eab60c, {16'd19065, 16'd19652, 16'd17488, 16'd42487, 16'd9424, 16'd62011, 16'd38518, 16'd33923, 16'd16124, 16'd10697, 16'd36110, 16'd39132, 16'd14670, 16'd63128, 16'd46641, 16'd14252, 16'd38934, 16'd58343, 16'd9156, 16'd44232, 16'd51078, 16'd32641, 16'd53430, 16'd39376, 16'd13277, 16'd13620});
	test_expansion(128'h65a58f0a9f012cd7f3ce9b02ae26f9ea, {16'd52809, 16'd55876, 16'd53084, 16'd37508, 16'd48134, 16'd45131, 16'd55237, 16'd9764, 16'd15077, 16'd54024, 16'd40212, 16'd604, 16'd61562, 16'd53292, 16'd16606, 16'd54909, 16'd14956, 16'd11779, 16'd15230, 16'd35664, 16'd25212, 16'd32330, 16'd25449, 16'd41683, 16'd35639, 16'd48644});
	test_expansion(128'h2576002cdf962b6b86d0b1221e8b11df, {16'd29216, 16'd13817, 16'd50031, 16'd15721, 16'd27914, 16'd33657, 16'd4618, 16'd13184, 16'd4819, 16'd17352, 16'd40590, 16'd4389, 16'd32110, 16'd45451, 16'd44304, 16'd46412, 16'd62906, 16'd42503, 16'd31469, 16'd21130, 16'd20273, 16'd799, 16'd7432, 16'd38939, 16'd4609, 16'd63855});
	test_expansion(128'h5d1bae89f43baa91d300b6bf383c695f, {16'd39680, 16'd8508, 16'd55315, 16'd11886, 16'd35479, 16'd54628, 16'd60038, 16'd28456, 16'd19280, 16'd20884, 16'd29279, 16'd21083, 16'd32316, 16'd53204, 16'd59737, 16'd26735, 16'd2817, 16'd46964, 16'd28310, 16'd40716, 16'd44300, 16'd34308, 16'd44383, 16'd24887, 16'd14344, 16'd19007});
	test_expansion(128'h6e095af7b72bf7d844c8757c3e824203, {16'd57642, 16'd35217, 16'd42689, 16'd44175, 16'd59351, 16'd125, 16'd50567, 16'd909, 16'd57898, 16'd64819, 16'd38542, 16'd62350, 16'd34154, 16'd25027, 16'd16521, 16'd26256, 16'd57753, 16'd17769, 16'd26840, 16'd59807, 16'd951, 16'd52045, 16'd7927, 16'd3757, 16'd48199, 16'd26891});
	test_expansion(128'h88559c0f4fb5e5e139026eaf35041263, {16'd11270, 16'd27169, 16'd31436, 16'd53426, 16'd16647, 16'd62754, 16'd6687, 16'd18588, 16'd45552, 16'd35600, 16'd47502, 16'd12706, 16'd11347, 16'd24550, 16'd4606, 16'd54766, 16'd52921, 16'd47725, 16'd12124, 16'd47296, 16'd38631, 16'd25318, 16'd40350, 16'd7889, 16'd46345, 16'd44885});
	test_expansion(128'h008f2ec6e59ac8cad511a343e215d769, {16'd31205, 16'd4938, 16'd45616, 16'd47263, 16'd27334, 16'd64159, 16'd62516, 16'd6826, 16'd34145, 16'd43326, 16'd42124, 16'd35551, 16'd24950, 16'd5292, 16'd43131, 16'd50056, 16'd32567, 16'd14365, 16'd9391, 16'd11516, 16'd49122, 16'd38211, 16'd9460, 16'd8812, 16'd15951, 16'd16500});
	test_expansion(128'h86a555fe884b022902a9bc58d767ba1f, {16'd1164, 16'd549, 16'd25482, 16'd13377, 16'd50648, 16'd43121, 16'd56403, 16'd65480, 16'd19304, 16'd61721, 16'd30963, 16'd38841, 16'd56846, 16'd47828, 16'd5742, 16'd32582, 16'd62563, 16'd64968, 16'd18879, 16'd31613, 16'd32986, 16'd11809, 16'd15355, 16'd5034, 16'd13577, 16'd51574});
	test_expansion(128'he42271803a04471b1ff51caf7976514c, {16'd18560, 16'd28691, 16'd57081, 16'd9839, 16'd11588, 16'd22332, 16'd1985, 16'd47860, 16'd50042, 16'd31498, 16'd63419, 16'd59009, 16'd10778, 16'd59541, 16'd10133, 16'd45877, 16'd4467, 16'd5831, 16'd7072, 16'd51118, 16'd31645, 16'd20505, 16'd64624, 16'd22750, 16'd27470, 16'd19306});
	test_expansion(128'h33f83111ad26125d50adcb895387e549, {16'd54595, 16'd58758, 16'd48466, 16'd3677, 16'd19958, 16'd6315, 16'd64657, 16'd54033, 16'd10331, 16'd6809, 16'd6575, 16'd1315, 16'd24463, 16'd24995, 16'd36785, 16'd26635, 16'd19919, 16'd33461, 16'd31628, 16'd59142, 16'd34587, 16'd60622, 16'd10542, 16'd24524, 16'd21024, 16'd36664});
	test_expansion(128'hc26f638b356bd7b6528745ce329092b3, {16'd1935, 16'd87, 16'd18499, 16'd25207, 16'd52478, 16'd51547, 16'd60542, 16'd52688, 16'd1059, 16'd39562, 16'd9054, 16'd5297, 16'd60692, 16'd48268, 16'd59316, 16'd26679, 16'd29062, 16'd14077, 16'd41434, 16'd64899, 16'd48338, 16'd47214, 16'd8299, 16'd30418, 16'd14813, 16'd56656});
	test_expansion(128'hab3682c84a9d3d16cb2c9209e1e7f71b, {16'd36632, 16'd31827, 16'd40779, 16'd31068, 16'd59089, 16'd14258, 16'd3152, 16'd58310, 16'd22336, 16'd5639, 16'd20570, 16'd45470, 16'd6344, 16'd49463, 16'd64486, 16'd52978, 16'd35827, 16'd32516, 16'd22989, 16'd58187, 16'd51331, 16'd59576, 16'd6091, 16'd45203, 16'd61550, 16'd55027});
	test_expansion(128'h4c4875e5040784d4a02b0330c04f3c92, {16'd20555, 16'd9789, 16'd62778, 16'd9792, 16'd49756, 16'd34567, 16'd4286, 16'd12703, 16'd49940, 16'd27499, 16'd15263, 16'd20591, 16'd43045, 16'd57469, 16'd58249, 16'd53206, 16'd10081, 16'd29692, 16'd53369, 16'd19361, 16'd47699, 16'd25366, 16'd5871, 16'd9240, 16'd15795, 16'd36756});
	test_expansion(128'hf40eb3355f0da86e4a3ee0917d3e99ca, {16'd40613, 16'd31383, 16'd63505, 16'd58885, 16'd14498, 16'd42178, 16'd38774, 16'd43660, 16'd51220, 16'd20931, 16'd43484, 16'd25159, 16'd15245, 16'd42192, 16'd21492, 16'd62994, 16'd20185, 16'd6689, 16'd47500, 16'd63095, 16'd49298, 16'd40989, 16'd20342, 16'd36706, 16'd8007, 16'd31384});
	test_expansion(128'hc339b34917e8f044f69e4a5928d9fc6a, {16'd44988, 16'd30125, 16'd44074, 16'd47366, 16'd13543, 16'd26219, 16'd17433, 16'd45632, 16'd45501, 16'd49912, 16'd41225, 16'd6860, 16'd49513, 16'd22458, 16'd43671, 16'd5990, 16'd39497, 16'd29220, 16'd42641, 16'd5359, 16'd37284, 16'd27159, 16'd30637, 16'd47170, 16'd35521, 16'd5343});
	test_expansion(128'h0cdbb95cf442169ca8dfd6599b2fb891, {16'd58298, 16'd3998, 16'd58845, 16'd37044, 16'd54105, 16'd4002, 16'd42335, 16'd48066, 16'd55904, 16'd62062, 16'd45793, 16'd9069, 16'd26318, 16'd29142, 16'd21489, 16'd63621, 16'd51639, 16'd9251, 16'd34172, 16'd47995, 16'd37573, 16'd44843, 16'd55235, 16'd5605, 16'd6456, 16'd41639});
	test_expansion(128'h00625aef4fa9e9cd0463b4f79dcd667b, {16'd21777, 16'd7233, 16'd41243, 16'd56428, 16'd59356, 16'd15729, 16'd50021, 16'd41646, 16'd51150, 16'd11512, 16'd40875, 16'd11196, 16'd50105, 16'd2336, 16'd3043, 16'd46691, 16'd9303, 16'd202, 16'd3627, 16'd57839, 16'd6617, 16'd26530, 16'd56705, 16'd22392, 16'd8927, 16'd36781});
	test_expansion(128'h9430a88c78154d14e151dbce1c938cb3, {16'd9198, 16'd51475, 16'd49987, 16'd52392, 16'd21435, 16'd32127, 16'd27109, 16'd15815, 16'd29356, 16'd21516, 16'd26722, 16'd59203, 16'd40642, 16'd8985, 16'd59361, 16'd11919, 16'd65453, 16'd37396, 16'd56494, 16'd42038, 16'd45539, 16'd55056, 16'd39299, 16'd64450, 16'd3443, 16'd28814});
	test_expansion(128'h31a0c3f436eec9148a0bf9cf9c2e6a1c, {16'd48451, 16'd45851, 16'd9115, 16'd4619, 16'd12787, 16'd29873, 16'd63405, 16'd40585, 16'd50673, 16'd57307, 16'd4223, 16'd54987, 16'd9110, 16'd15582, 16'd34053, 16'd8059, 16'd34607, 16'd52108, 16'd38063, 16'd9601, 16'd24680, 16'd7775, 16'd22636, 16'd13571, 16'd10589, 16'd8249});
	test_expansion(128'he6886c8cfe05dc3e5f7df1180213796f, {16'd51153, 16'd15377, 16'd54654, 16'd65080, 16'd4179, 16'd28937, 16'd156, 16'd27609, 16'd36820, 16'd62277, 16'd51152, 16'd59264, 16'd25276, 16'd25697, 16'd8913, 16'd36863, 16'd11845, 16'd7964, 16'd48488, 16'd13709, 16'd33049, 16'd17685, 16'd11380, 16'd40173, 16'd8129, 16'd25628});
	test_expansion(128'h7ff2b2af8aa60a309e3e1d51ea0e1fab, {16'd63151, 16'd38945, 16'd42359, 16'd51264, 16'd55147, 16'd28170, 16'd11649, 16'd32502, 16'd14194, 16'd26035, 16'd29805, 16'd22719, 16'd59897, 16'd20039, 16'd37468, 16'd26247, 16'd25656, 16'd41366, 16'd27972, 16'd37610, 16'd57915, 16'd37686, 16'd49750, 16'd3220, 16'd48112, 16'd12190});
	test_expansion(128'hed127d2bfd7812674bc5ad4e2295c455, {16'd27657, 16'd55184, 16'd28698, 16'd22350, 16'd123, 16'd59187, 16'd5202, 16'd31817, 16'd44104, 16'd25858, 16'd56230, 16'd45277, 16'd44788, 16'd28661, 16'd65374, 16'd65107, 16'd31490, 16'd597, 16'd57129, 16'd14424, 16'd40390, 16'd38764, 16'd23985, 16'd18102, 16'd61722, 16'd24226});
	test_expansion(128'ha24941b94273f32f7f64d6b91e327ee0, {16'd49227, 16'd28093, 16'd36936, 16'd27437, 16'd48977, 16'd47204, 16'd6801, 16'd13781, 16'd45978, 16'd45560, 16'd62750, 16'd65374, 16'd25148, 16'd47411, 16'd63863, 16'd25181, 16'd21679, 16'd10786, 16'd25538, 16'd23114, 16'd24848, 16'd19697, 16'd8366, 16'd6751, 16'd42724, 16'd49986});
	test_expansion(128'h81df45bf743db97c4f16c9d79c6a1154, {16'd28166, 16'd59726, 16'd26736, 16'd55412, 16'd19358, 16'd46174, 16'd44750, 16'd10087, 16'd22216, 16'd16888, 16'd25147, 16'd31894, 16'd6067, 16'd43600, 16'd2429, 16'd15449, 16'd57429, 16'd14660, 16'd48865, 16'd41067, 16'd36323, 16'd63985, 16'd53672, 16'd543, 16'd5201, 16'd2156});
	test_expansion(128'h83eb7f02323317a82a08ecfbd1562635, {16'd10768, 16'd23247, 16'd36706, 16'd62189, 16'd1776, 16'd7334, 16'd668, 16'd7710, 16'd55594, 16'd62254, 16'd896, 16'd32198, 16'd24017, 16'd27507, 16'd5171, 16'd54966, 16'd50066, 16'd36019, 16'd60184, 16'd48250, 16'd7620, 16'd41599, 16'd59829, 16'd24749, 16'd12549, 16'd9204});
	test_expansion(128'hf9e882d5621ab00895bf3f1fb77508d3, {16'd61198, 16'd13032, 16'd59035, 16'd6181, 16'd43710, 16'd3518, 16'd64176, 16'd14082, 16'd43746, 16'd24145, 16'd2262, 16'd31712, 16'd45302, 16'd56641, 16'd59993, 16'd63147, 16'd18489, 16'd42320, 16'd63426, 16'd50155, 16'd43465, 16'd20876, 16'd55978, 16'd53859, 16'd28254, 16'd22081});
	test_expansion(128'h9e24123753ab93e0a8c20f45c63356c7, {16'd25650, 16'd52332, 16'd31337, 16'd12505, 16'd41775, 16'd51522, 16'd49459, 16'd56279, 16'd57855, 16'd62047, 16'd30176, 16'd9869, 16'd26841, 16'd55434, 16'd60215, 16'd40246, 16'd6187, 16'd22289, 16'd22128, 16'd61761, 16'd5828, 16'd138, 16'd62482, 16'd15544, 16'd26082, 16'd12624});
	test_expansion(128'h4a9e804ef4a4e7b68a180078464524de, {16'd42795, 16'd7404, 16'd8911, 16'd8971, 16'd12278, 16'd5793, 16'd24081, 16'd37639, 16'd21465, 16'd27468, 16'd64593, 16'd29562, 16'd35271, 16'd8837, 16'd18206, 16'd7479, 16'd54441, 16'd48547, 16'd24012, 16'd23776, 16'd4004, 16'd4564, 16'd25236, 16'd53439, 16'd54229, 16'd4597});
	test_expansion(128'h4f3b1004363ab4442f5e26b74e4b149e, {16'd290, 16'd43094, 16'd28807, 16'd9328, 16'd19410, 16'd36574, 16'd22998, 16'd61645, 16'd65179, 16'd51256, 16'd33891, 16'd38378, 16'd50355, 16'd27041, 16'd64203, 16'd5432, 16'd30888, 16'd65060, 16'd5949, 16'd26408, 16'd46801, 16'd38689, 16'd48244, 16'd1966, 16'd54551, 16'd64348});
	test_expansion(128'hd56c987d1a30c74fd068183f3f235393, {16'd40712, 16'd51448, 16'd55392, 16'd9600, 16'd48436, 16'd23463, 16'd37798, 16'd27810, 16'd4515, 16'd60249, 16'd37086, 16'd42761, 16'd48703, 16'd10927, 16'd43047, 16'd29134, 16'd45548, 16'd11272, 16'd45828, 16'd60903, 16'd45581, 16'd59024, 16'd65163, 16'd47258, 16'd15885, 16'd25471});
	test_expansion(128'h930e9f0b9c0a7c0cbcc0d0e28c8ef084, {16'd9241, 16'd60379, 16'd29332, 16'd20748, 16'd45125, 16'd26514, 16'd20661, 16'd24882, 16'd24029, 16'd23959, 16'd1501, 16'd18752, 16'd41596, 16'd33316, 16'd52201, 16'd18900, 16'd6685, 16'd52964, 16'd11504, 16'd22005, 16'd58488, 16'd47884, 16'd44212, 16'd25119, 16'd48360, 16'd62145});
	test_expansion(128'h52322776444c2202123b37ec4661d367, {16'd38947, 16'd57253, 16'd46848, 16'd60579, 16'd19955, 16'd46696, 16'd63922, 16'd31847, 16'd52928, 16'd33572, 16'd40041, 16'd171, 16'd33843, 16'd6400, 16'd25913, 16'd4278, 16'd22542, 16'd5817, 16'd3271, 16'd56509, 16'd27536, 16'd40242, 16'd51053, 16'd13268, 16'd27297, 16'd32112});
	test_expansion(128'h860a1f0f7cb26f45e3ef242a41ec147f, {16'd60555, 16'd4090, 16'd51816, 16'd32331, 16'd23191, 16'd48026, 16'd12377, 16'd48075, 16'd50855, 16'd8911, 16'd27221, 16'd52717, 16'd41454, 16'd47609, 16'd37179, 16'd5227, 16'd53364, 16'd18159, 16'd36212, 16'd7861, 16'd23447, 16'd6722, 16'd31980, 16'd16791, 16'd49068, 16'd15957});
	test_expansion(128'hcc11840c9b10fc181934ad21845d653d, {16'd8538, 16'd41784, 16'd20362, 16'd54870, 16'd40024, 16'd23346, 16'd57325, 16'd13238, 16'd21857, 16'd21387, 16'd47805, 16'd34369, 16'd21332, 16'd3838, 16'd52343, 16'd42277, 16'd20413, 16'd22322, 16'd1626, 16'd57327, 16'd44514, 16'd25709, 16'd34465, 16'd61945, 16'd20843, 16'd5439});
	test_expansion(128'h137c178af7fc6b7b1532e7e0b1f46918, {16'd50624, 16'd63294, 16'd20743, 16'd43100, 16'd62575, 16'd38882, 16'd10942, 16'd51627, 16'd15217, 16'd34137, 16'd16570, 16'd64718, 16'd15912, 16'd34351, 16'd35849, 16'd4508, 16'd23892, 16'd13933, 16'd9966, 16'd54356, 16'd33106, 16'd57299, 16'd13238, 16'd27250, 16'd47095, 16'd16860});
	test_expansion(128'h39aa7cfb44ef918576ce9d4b2505cd34, {16'd2320, 16'd62028, 16'd39325, 16'd14910, 16'd60499, 16'd48639, 16'd63757, 16'd35439, 16'd12539, 16'd45816, 16'd20999, 16'd39904, 16'd45141, 16'd39608, 16'd10573, 16'd45746, 16'd16235, 16'd39275, 16'd51644, 16'd20073, 16'd6011, 16'd24693, 16'd54372, 16'd8593, 16'd1500, 16'd33589});
	test_expansion(128'h73778535bf2019f6a1b594a96261e136, {16'd9372, 16'd11755, 16'd46003, 16'd8118, 16'd30379, 16'd50212, 16'd57742, 16'd33795, 16'd24709, 16'd61906, 16'd28137, 16'd22909, 16'd58788, 16'd58208, 16'd53721, 16'd13761, 16'd5658, 16'd11835, 16'd32564, 16'd65132, 16'd1891, 16'd36476, 16'd27373, 16'd13863, 16'd54416, 16'd17338});
	test_expansion(128'hc4fb44396bcb06073111c76e5005a1cc, {16'd32869, 16'd12704, 16'd36393, 16'd40123, 16'd44624, 16'd19872, 16'd48538, 16'd4867, 16'd53539, 16'd23742, 16'd41788, 16'd7659, 16'd35759, 16'd51941, 16'd57679, 16'd2296, 16'd22341, 16'd60070, 16'd13277, 16'd11379, 16'd43152, 16'd13395, 16'd18975, 16'd40917, 16'd27092, 16'd64466});
	test_expansion(128'h239fbfe3633d9a4ea312fd854204e0f6, {16'd3292, 16'd15782, 16'd56633, 16'd39628, 16'd29894, 16'd27076, 16'd9151, 16'd48271, 16'd31013, 16'd60795, 16'd9709, 16'd14127, 16'd6050, 16'd23020, 16'd59084, 16'd35566, 16'd5286, 16'd56252, 16'd39513, 16'd34413, 16'd40138, 16'd31054, 16'd5030, 16'd9566, 16'd43160, 16'd15923});
	test_expansion(128'h16ca6269bc2ef6907e67acdefd0107fd, {16'd61369, 16'd24280, 16'd22873, 16'd10734, 16'd13954, 16'd49862, 16'd56256, 16'd39031, 16'd29991, 16'd42530, 16'd64070, 16'd53943, 16'd40696, 16'd13008, 16'd33194, 16'd8654, 16'd12649, 16'd32378, 16'd4505, 16'd48830, 16'd62412, 16'd65187, 16'd55313, 16'd40987, 16'd11755, 16'd45263});
	test_expansion(128'h1f7c0835359190c1e1812f985731b1c9, {16'd30832, 16'd52880, 16'd16460, 16'd18952, 16'd35898, 16'd13757, 16'd40763, 16'd58016, 16'd3542, 16'd46257, 16'd44783, 16'd7457, 16'd29290, 16'd26699, 16'd22025, 16'd47167, 16'd13406, 16'd2765, 16'd3046, 16'd14470, 16'd27279, 16'd40739, 16'd58489, 16'd6442, 16'd8921, 16'd14763});
	test_expansion(128'h69a24235db40523a767f2016ed550cd9, {16'd64566, 16'd37408, 16'd8147, 16'd33368, 16'd55681, 16'd36096, 16'd25431, 16'd64323, 16'd1988, 16'd60168, 16'd62956, 16'd13905, 16'd46604, 16'd3113, 16'd60527, 16'd62999, 16'd47438, 16'd24592, 16'd45270, 16'd32122, 16'd7629, 16'd52175, 16'd11139, 16'd56372, 16'd13624, 16'd17890});
	test_expansion(128'h679d6d3712bbd58693712ccc352298b6, {16'd59140, 16'd19299, 16'd34296, 16'd25113, 16'd47655, 16'd48325, 16'd37660, 16'd51272, 16'd7964, 16'd30934, 16'd56715, 16'd41988, 16'd64055, 16'd52284, 16'd16320, 16'd18795, 16'd63585, 16'd6680, 16'd54961, 16'd2025, 16'd5037, 16'd23242, 16'd61021, 16'd50150, 16'd13746, 16'd22968});
	test_expansion(128'hb282dc29c0be68520e1217dbebc63ac4, {16'd61440, 16'd3066, 16'd52438, 16'd23583, 16'd40143, 16'd43194, 16'd6945, 16'd48806, 16'd14419, 16'd25223, 16'd8530, 16'd4588, 16'd31075, 16'd2201, 16'd1165, 16'd19053, 16'd43151, 16'd39165, 16'd60724, 16'd15516, 16'd58533, 16'd2853, 16'd15367, 16'd60092, 16'd33270, 16'd6015});
	test_expansion(128'hd38a410fc92e5575232d9eabba7e2871, {16'd23359, 16'd31339, 16'd49522, 16'd7849, 16'd25439, 16'd11968, 16'd55623, 16'd14914, 16'd5065, 16'd60663, 16'd55399, 16'd18182, 16'd28219, 16'd22650, 16'd9026, 16'd3900, 16'd46031, 16'd40807, 16'd24054, 16'd3003, 16'd37695, 16'd19097, 16'd52761, 16'd29656, 16'd64507, 16'd474});
	test_expansion(128'hbaadea6b5ea09cf1e534e5ea74132d35, {16'd29605, 16'd46918, 16'd15268, 16'd6649, 16'd53895, 16'd28199, 16'd56198, 16'd58923, 16'd61002, 16'd10064, 16'd9790, 16'd43252, 16'd19529, 16'd51842, 16'd44711, 16'd57810, 16'd1940, 16'd60348, 16'd53207, 16'd52070, 16'd31447, 16'd42968, 16'd1303, 16'd26200, 16'd50443, 16'd584});
	test_expansion(128'h13ce2dbe0cd599576eca8b7fa05088ac, {16'd25019, 16'd59080, 16'd7301, 16'd51815, 16'd42032, 16'd25188, 16'd2870, 16'd36523, 16'd44192, 16'd12507, 16'd8513, 16'd42538, 16'd50672, 16'd39228, 16'd15847, 16'd45892, 16'd58751, 16'd9348, 16'd50728, 16'd21666, 16'd55264, 16'd19974, 16'd18238, 16'd42784, 16'd24980, 16'd47713});
	test_expansion(128'hb51c13bc1aab905fda3728a394ccc656, {16'd2066, 16'd14695, 16'd60288, 16'd6275, 16'd51987, 16'd5921, 16'd56171, 16'd41497, 16'd23797, 16'd40709, 16'd14616, 16'd46079, 16'd2039, 16'd4790, 16'd50936, 16'd62400, 16'd11895, 16'd32757, 16'd12049, 16'd2269, 16'd12625, 16'd16088, 16'd45665, 16'd37478, 16'd29985, 16'd47315});
	test_expansion(128'h08647b00748feed67642e4622945764f, {16'd55637, 16'd19376, 16'd6913, 16'd27423, 16'd29689, 16'd39135, 16'd31652, 16'd13927, 16'd30584, 16'd4954, 16'd56984, 16'd43988, 16'd33275, 16'd57038, 16'd36294, 16'd45391, 16'd51395, 16'd36320, 16'd21342, 16'd59458, 16'd43837, 16'd46880, 16'd48865, 16'd33045, 16'd1606, 16'd13838});
	test_expansion(128'h8d75c87dad9dbbf4b7052df1282309b0, {16'd19561, 16'd12833, 16'd18190, 16'd41019, 16'd59321, 16'd63927, 16'd46880, 16'd60302, 16'd19089, 16'd23929, 16'd17535, 16'd9058, 16'd6775, 16'd27756, 16'd25708, 16'd62439, 16'd59562, 16'd54608, 16'd42956, 16'd16174, 16'd31692, 16'd37428, 16'd60087, 16'd25176, 16'd24448, 16'd48807});
	test_expansion(128'h5484abd8d8be21527b24047700db4836, {16'd47691, 16'd62815, 16'd16315, 16'd57274, 16'd10147, 16'd19111, 16'd48548, 16'd47285, 16'd28988, 16'd27623, 16'd36234, 16'd36845, 16'd47074, 16'd10770, 16'd20865, 16'd45122, 16'd7374, 16'd50535, 16'd33139, 16'd37834, 16'd54098, 16'd37947, 16'd26525, 16'd14944, 16'd7310, 16'd9779});
	test_expansion(128'h4067ff700b13dfcb8c927f5390a21f95, {16'd54197, 16'd30242, 16'd16500, 16'd47681, 16'd376, 16'd17752, 16'd25843, 16'd18287, 16'd44759, 16'd28951, 16'd52380, 16'd8852, 16'd61421, 16'd33594, 16'd37349, 16'd53261, 16'd7068, 16'd46694, 16'd29106, 16'd48541, 16'd60097, 16'd2845, 16'd6567, 16'd22631, 16'd9989, 16'd1818});
	test_expansion(128'hb4a53539f8c5c79a7ae3fa1c4d178a17, {16'd28336, 16'd1049, 16'd7625, 16'd54287, 16'd2017, 16'd22434, 16'd23306, 16'd30262, 16'd17884, 16'd39940, 16'd57292, 16'd4736, 16'd59165, 16'd23952, 16'd28045, 16'd57885, 16'd20136, 16'd60932, 16'd11813, 16'd36297, 16'd60963, 16'd3869, 16'd25484, 16'd23080, 16'd57651, 16'd4322});
	test_expansion(128'h42a0f49aa8d92381cd4f5f3c76deac68, {16'd53481, 16'd23479, 16'd27409, 16'd46133, 16'd26659, 16'd29878, 16'd50547, 16'd7732, 16'd60032, 16'd30941, 16'd3277, 16'd5397, 16'd25071, 16'd24357, 16'd25045, 16'd26705, 16'd60668, 16'd57712, 16'd43731, 16'd3337, 16'd15808, 16'd52324, 16'd16460, 16'd11846, 16'd29980, 16'd61758});
	test_expansion(128'hc80489b88c05095c573ca97a0b3eaa4f, {16'd38234, 16'd19584, 16'd34475, 16'd44570, 16'd36402, 16'd39009, 16'd10878, 16'd35928, 16'd6365, 16'd1184, 16'd15418, 16'd51028, 16'd45899, 16'd7265, 16'd35909, 16'd3849, 16'd57616, 16'd39551, 16'd51250, 16'd30141, 16'd29608, 16'd26017, 16'd61950, 16'd36718, 16'd19276, 16'd42029});
	test_expansion(128'ha500caf43a85043d4b062417818562a9, {16'd48878, 16'd27788, 16'd35402, 16'd17499, 16'd30001, 16'd46877, 16'd40911, 16'd40850, 16'd50934, 16'd13075, 16'd43967, 16'd61551, 16'd58747, 16'd44430, 16'd690, 16'd31155, 16'd4040, 16'd54650, 16'd10711, 16'd7708, 16'd14697, 16'd27301, 16'd25912, 16'd8297, 16'd48141, 16'd3022});
	test_expansion(128'heb2acd6b4a4dabe4c97ff57180a98302, {16'd23653, 16'd42613, 16'd37139, 16'd61528, 16'd9318, 16'd20124, 16'd16410, 16'd5058, 16'd43111, 16'd15163, 16'd33867, 16'd62389, 16'd61849, 16'd16817, 16'd40019, 16'd49220, 16'd7304, 16'd38539, 16'd9791, 16'd26991, 16'd23860, 16'd55755, 16'd1898, 16'd59425, 16'd61692, 16'd17477});
	test_expansion(128'h8b556641e3184c871a02de305986765b, {16'd6433, 16'd46501, 16'd25855, 16'd60549, 16'd33215, 16'd41152, 16'd33786, 16'd6728, 16'd59341, 16'd61504, 16'd22749, 16'd44274, 16'd48007, 16'd3320, 16'd57340, 16'd6470, 16'd23860, 16'd37847, 16'd35940, 16'd6027, 16'd64296, 16'd26304, 16'd5680, 16'd5496, 16'd36536, 16'd34959});
	test_expansion(128'hbf97629f2f6ed940d65dfc0c79532a8c, {16'd38890, 16'd37809, 16'd19878, 16'd33608, 16'd25120, 16'd10982, 16'd45855, 16'd55277, 16'd23530, 16'd63380, 16'd48057, 16'd37760, 16'd26381, 16'd3839, 16'd47714, 16'd2621, 16'd22187, 16'd46534, 16'd46811, 16'd12308, 16'd64454, 16'd6766, 16'd27378, 16'd32300, 16'd48617, 16'd60215});
	test_expansion(128'hd0c2881be1a257811432882296e32870, {16'd1171, 16'd32198, 16'd55542, 16'd60475, 16'd59540, 16'd34096, 16'd65008, 16'd30420, 16'd58315, 16'd27762, 16'd41833, 16'd29418, 16'd61995, 16'd17845, 16'd6950, 16'd63358, 16'd44801, 16'd21481, 16'd4556, 16'd40380, 16'd57289, 16'd52850, 16'd28965, 16'd15811, 16'd33935, 16'd35031});
	test_expansion(128'h1222263cb0b71ed95d4e07285cd4fe84, {16'd43392, 16'd36614, 16'd59314, 16'd683, 16'd6971, 16'd59480, 16'd33382, 16'd58792, 16'd2336, 16'd23327, 16'd26217, 16'd37024, 16'd42785, 16'd1676, 16'd24396, 16'd29756, 16'd25155, 16'd43120, 16'd54221, 16'd11849, 16'd55121, 16'd62287, 16'd9687, 16'd45128, 16'd19579, 16'd59098});
	test_expansion(128'h9bf90cbae3877d444a7c39142bec0a40, {16'd62465, 16'd33807, 16'd49651, 16'd63918, 16'd26810, 16'd47702, 16'd14652, 16'd36022, 16'd36289, 16'd15, 16'd64332, 16'd18716, 16'd63298, 16'd26175, 16'd42582, 16'd39199, 16'd15227, 16'd51290, 16'd26513, 16'd1876, 16'd56685, 16'd37384, 16'd33270, 16'd48054, 16'd39465, 16'd44282});
	test_expansion(128'h8d1703a704c916075b99ed083323298a, {16'd49723, 16'd57325, 16'd23777, 16'd2549, 16'd53031, 16'd47729, 16'd59265, 16'd53970, 16'd25344, 16'd26903, 16'd50027, 16'd12801, 16'd1853, 16'd30155, 16'd27788, 16'd17398, 16'd19493, 16'd44634, 16'd22526, 16'd24450, 16'd32918, 16'd61561, 16'd14306, 16'd19560, 16'd40869, 16'd2810});
	test_expansion(128'heb11df8444d0bf925c1a05839d6c0563, {16'd41553, 16'd13805, 16'd20367, 16'd38791, 16'd7273, 16'd3995, 16'd35005, 16'd3160, 16'd45947, 16'd55053, 16'd51151, 16'd42504, 16'd5792, 16'd53622, 16'd60938, 16'd32144, 16'd49685, 16'd59048, 16'd43075, 16'd4861, 16'd33898, 16'd5415, 16'd39590, 16'd19119, 16'd44220, 16'd45470});
	test_expansion(128'h647b13ce64ba32add8ae54471a841e9b, {16'd16394, 16'd32177, 16'd49662, 16'd59491, 16'd58290, 16'd61999, 16'd31267, 16'd64176, 16'd1631, 16'd13651, 16'd51363, 16'd53716, 16'd12874, 16'd30389, 16'd40899, 16'd11044, 16'd6791, 16'd65390, 16'd27943, 16'd18984, 16'd31590, 16'd53955, 16'd59190, 16'd6480, 16'd39574, 16'd13357});
	test_expansion(128'hd85cbb35ed60be56533aee62f3823b17, {16'd33041, 16'd61178, 16'd45463, 16'd28411, 16'd28999, 16'd20349, 16'd31732, 16'd27315, 16'd29546, 16'd46560, 16'd34864, 16'd64914, 16'd26102, 16'd31908, 16'd32144, 16'd34461, 16'd12164, 16'd27425, 16'd59438, 16'd24438, 16'd497, 16'd15759, 16'd37321, 16'd2104, 16'd6516, 16'd63644});
	test_expansion(128'h38e88f5d474bbe3f0ebc337a7031b33e, {16'd24837, 16'd26374, 16'd57579, 16'd19316, 16'd5420, 16'd12227, 16'd42672, 16'd4203, 16'd61863, 16'd61906, 16'd65160, 16'd49803, 16'd62933, 16'd61723, 16'd53245, 16'd13348, 16'd13464, 16'd29663, 16'd58435, 16'd24906, 16'd17858, 16'd28570, 16'd6341, 16'd26299, 16'd53800, 16'd31451});
	test_expansion(128'h20f83fb91e01cfff91a05b95fab7ae1d, {16'd37922, 16'd6269, 16'd37333, 16'd9658, 16'd6979, 16'd35634, 16'd50563, 16'd19094, 16'd51026, 16'd21822, 16'd61222, 16'd49379, 16'd20909, 16'd62122, 16'd5222, 16'd4961, 16'd22969, 16'd6857, 16'd30921, 16'd21394, 16'd13799, 16'd6702, 16'd11711, 16'd58489, 16'd27338, 16'd64351});
	test_expansion(128'h293fefa9ec311b2dce57a52b4388ed58, {16'd30370, 16'd47845, 16'd25960, 16'd761, 16'd20231, 16'd41568, 16'd48988, 16'd50216, 16'd49495, 16'd23324, 16'd55546, 16'd7144, 16'd40083, 16'd64196, 16'd51173, 16'd52811, 16'd48187, 16'd54709, 16'd17318, 16'd35459, 16'd4106, 16'd50880, 16'd41758, 16'd8632, 16'd57885, 16'd5472});
	test_expansion(128'h07fa44da9b82c32981d36fdb6380eaf2, {16'd45519, 16'd41799, 16'd54705, 16'd29344, 16'd56793, 16'd54850, 16'd24257, 16'd61779, 16'd22966, 16'd31276, 16'd6123, 16'd4922, 16'd59282, 16'd1103, 16'd15348, 16'd25370, 16'd56265, 16'd8183, 16'd52842, 16'd63224, 16'd62518, 16'd29721, 16'd56121, 16'd47308, 16'd53125, 16'd22115});
	test_expansion(128'h492ce1c0f9b97fdbf67e5d1792855126, {16'd58325, 16'd65309, 16'd3083, 16'd23022, 16'd63536, 16'd29302, 16'd48302, 16'd398, 16'd38064, 16'd53500, 16'd30617, 16'd36633, 16'd63978, 16'd36304, 16'd17244, 16'd45215, 16'd28399, 16'd48559, 16'd7194, 16'd43119, 16'd58332, 16'd13898, 16'd61345, 16'd31484, 16'd40780, 16'd29534});
	test_expansion(128'h76d1edf1bbdd823fe4ac02c025d30d29, {16'd9505, 16'd18671, 16'd14981, 16'd38588, 16'd25916, 16'd13313, 16'd36129, 16'd60989, 16'd49256, 16'd12193, 16'd53480, 16'd33531, 16'd56181, 16'd33988, 16'd14899, 16'd45983, 16'd8076, 16'd27813, 16'd53604, 16'd9995, 16'd40848, 16'd11820, 16'd60440, 16'd42117, 16'd32305, 16'd29073});
	test_expansion(128'h70bd7017874ea132ed86992e626a5fc5, {16'd30416, 16'd29256, 16'd32504, 16'd44505, 16'd57488, 16'd16636, 16'd2329, 16'd37948, 16'd51960, 16'd43768, 16'd44908, 16'd14524, 16'd21207, 16'd56901, 16'd53268, 16'd6756, 16'd47552, 16'd61340, 16'd846, 16'd63303, 16'd43211, 16'd62041, 16'd17639, 16'd43360, 16'd59884, 16'd22954});
	test_expansion(128'h92850cc4df872b4898fb102c79769df6, {16'd45929, 16'd39472, 16'd63496, 16'd57769, 16'd36935, 16'd38449, 16'd50684, 16'd46238, 16'd59212, 16'd29507, 16'd47667, 16'd55533, 16'd24855, 16'd30301, 16'd8554, 16'd19353, 16'd18449, 16'd11525, 16'd39149, 16'd39058, 16'd44770, 16'd53575, 16'd27223, 16'd7837, 16'd48478, 16'd34981});
	test_expansion(128'h1fb4d977df80268f752746ee90e70a88, {16'd51469, 16'd64612, 16'd4401, 16'd47147, 16'd37326, 16'd20007, 16'd25429, 16'd37745, 16'd47224, 16'd34233, 16'd20381, 16'd37800, 16'd23029, 16'd61896, 16'd21701, 16'd60980, 16'd17900, 16'd2667, 16'd40416, 16'd5350, 16'd548, 16'd59524, 16'd54198, 16'd27179, 16'd7503, 16'd29834});
	test_expansion(128'h16799901c549caf55c055d211ea8d510, {16'd33458, 16'd15924, 16'd17983, 16'd48178, 16'd48630, 16'd47921, 16'd35191, 16'd1564, 16'd32957, 16'd9471, 16'd27379, 16'd6314, 16'd31133, 16'd4762, 16'd21822, 16'd23026, 16'd39619, 16'd61107, 16'd6258, 16'd63385, 16'd43372, 16'd4316, 16'd40706, 16'd29280, 16'd13624, 16'd8534});
	test_expansion(128'hc68f6a053d7d6935b26eb5d0df8b7b3e, {16'd34804, 16'd39443, 16'd29875, 16'd33565, 16'd30544, 16'd47208, 16'd47029, 16'd43424, 16'd44743, 16'd26212, 16'd28276, 16'd55485, 16'd57233, 16'd53131, 16'd9293, 16'd46088, 16'd52357, 16'd44576, 16'd40703, 16'd50138, 16'd39185, 16'd62621, 16'd35720, 16'd24621, 16'd41862, 16'd52640});
	test_expansion(128'h2c9e469812df7c734417f2987753a163, {16'd60914, 16'd28502, 16'd62103, 16'd49031, 16'd27712, 16'd18852, 16'd52823, 16'd54616, 16'd330, 16'd15128, 16'd40159, 16'd24459, 16'd17862, 16'd51524, 16'd63640, 16'd17314, 16'd3573, 16'd21198, 16'd4235, 16'd33737, 16'd14275, 16'd45315, 16'd46615, 16'd19329, 16'd48457, 16'd14761});
	test_expansion(128'hcccd80dae91889194a21cf126f0ac892, {16'd46336, 16'd29730, 16'd30227, 16'd10819, 16'd30488, 16'd20482, 16'd49280, 16'd54274, 16'd8247, 16'd14040, 16'd43389, 16'd20379, 16'd14847, 16'd29368, 16'd65143, 16'd5776, 16'd49736, 16'd45348, 16'd53515, 16'd12483, 16'd36725, 16'd23005, 16'd4419, 16'd33729, 16'd42221, 16'd2969});
	test_expansion(128'h26e1736437fceace7de2728a0f6725b6, {16'd36489, 16'd64222, 16'd44559, 16'd25746, 16'd6557, 16'd5087, 16'd35599, 16'd33190, 16'd50940, 16'd24847, 16'd7291, 16'd62529, 16'd36841, 16'd27039, 16'd17929, 16'd8789, 16'd18275, 16'd61706, 16'd1619, 16'd14482, 16'd40030, 16'd65148, 16'd38013, 16'd1589, 16'd44797, 16'd44487});
	test_expansion(128'h2b6fada194f028e49b23880085d78749, {16'd38368, 16'd15549, 16'd58686, 16'd60873, 16'd8143, 16'd65490, 16'd10733, 16'd23920, 16'd49979, 16'd11483, 16'd50263, 16'd25262, 16'd51365, 16'd5059, 16'd26448, 16'd31993, 16'd4217, 16'd36186, 16'd15176, 16'd25065, 16'd6082, 16'd54635, 16'd34244, 16'd64801, 16'd59139, 16'd14806});
	test_expansion(128'h9630a946fbd6b4624fe72cd6c07de6e6, {16'd32484, 16'd54805, 16'd19130, 16'd56424, 16'd51566, 16'd32161, 16'd55851, 16'd52650, 16'd9845, 16'd15577, 16'd25969, 16'd26107, 16'd61945, 16'd23565, 16'd41138, 16'd45618, 16'd40999, 16'd9196, 16'd33383, 16'd44496, 16'd10965, 16'd9143, 16'd20875, 16'd43992, 16'd27946, 16'd31723});
	test_expansion(128'h4a9924e8c1deb8dd5a20e17f9b656a5e, {16'd45856, 16'd49391, 16'd19713, 16'd42100, 16'd47966, 16'd58368, 16'd47247, 16'd5487, 16'd9166, 16'd24961, 16'd60201, 16'd38452, 16'd38320, 16'd36503, 16'd41438, 16'd36944, 16'd45413, 16'd60405, 16'd18458, 16'd28664, 16'd6875, 16'd5742, 16'd46588, 16'd53546, 16'd9529, 16'd20212});
	test_expansion(128'hc46ad693abe6d1fdef2f6791fbc9266f, {16'd26038, 16'd38493, 16'd20380, 16'd38883, 16'd19036, 16'd33053, 16'd64786, 16'd4574, 16'd31529, 16'd38916, 16'd51439, 16'd3152, 16'd37616, 16'd33014, 16'd38356, 16'd26140, 16'd65480, 16'd31148, 16'd18913, 16'd61493, 16'd41057, 16'd12181, 16'd52255, 16'd20501, 16'd22677, 16'd20205});
	test_expansion(128'hbe1ed46530d652986af599b27db065f9, {16'd1960, 16'd27406, 16'd59340, 16'd10513, 16'd13563, 16'd57602, 16'd6258, 16'd59440, 16'd4496, 16'd15691, 16'd29852, 16'd56622, 16'd47199, 16'd28933, 16'd60107, 16'd16592, 16'd2788, 16'd3955, 16'd26827, 16'd15317, 16'd1358, 16'd33088, 16'd33907, 16'd33865, 16'd51495, 16'd32918});
	test_expansion(128'h9344ce956fbb32f7dd04601e0896a69d, {16'd41981, 16'd45324, 16'd33542, 16'd13602, 16'd48497, 16'd536, 16'd25876, 16'd58497, 16'd45920, 16'd63914, 16'd28484, 16'd34809, 16'd31209, 16'd8734, 16'd37304, 16'd584, 16'd19928, 16'd36955, 16'd30046, 16'd39602, 16'd63895, 16'd15204, 16'd20744, 16'd24988, 16'd60669, 16'd46189});
	test_expansion(128'h7f13448b31d3cd6a3149c2a40a3172a0, {16'd45171, 16'd26619, 16'd33882, 16'd35225, 16'd13646, 16'd42973, 16'd9989, 16'd28381, 16'd34772, 16'd43254, 16'd28954, 16'd25083, 16'd46037, 16'd11642, 16'd53058, 16'd8668, 16'd10711, 16'd45991, 16'd7688, 16'd9678, 16'd12779, 16'd24192, 16'd16070, 16'd20006, 16'd60101, 16'd57670});
	test_expansion(128'h975d75d187bd2f2f8dd183c72294f30a, {16'd63874, 16'd1643, 16'd61666, 16'd28640, 16'd56321, 16'd10009, 16'd64704, 16'd17268, 16'd35842, 16'd17855, 16'd11632, 16'd45836, 16'd19214, 16'd29527, 16'd55772, 16'd12324, 16'd18550, 16'd63280, 16'd8117, 16'd28460, 16'd12087, 16'd17956, 16'd42755, 16'd50138, 16'd29602, 16'd31802});
	test_expansion(128'h2e0e9d312e6aeb2e58fead36de84c560, {16'd22269, 16'd45329, 16'd50326, 16'd47818, 16'd26510, 16'd27838, 16'd60041, 16'd18239, 16'd49361, 16'd59893, 16'd59926, 16'd25022, 16'd62731, 16'd53832, 16'd49286, 16'd2864, 16'd54954, 16'd56526, 16'd45331, 16'd20881, 16'd3422, 16'd57628, 16'd42672, 16'd61180, 16'd21823, 16'd6392});
	test_expansion(128'h6d73522714ab167a5bc1a7a1c43d3390, {16'd5347, 16'd709, 16'd4607, 16'd33955, 16'd2410, 16'd39799, 16'd11241, 16'd13035, 16'd14159, 16'd20988, 16'd32848, 16'd47008, 16'd59654, 16'd18634, 16'd14806, 16'd23628, 16'd1429, 16'd4730, 16'd39071, 16'd58158, 16'd50089, 16'd59537, 16'd28012, 16'd3773, 16'd13133, 16'd61089});
	test_expansion(128'hf31b4902e02d419a5a0e2432c2dbed57, {16'd53245, 16'd65013, 16'd19396, 16'd30414, 16'd36455, 16'd26257, 16'd33274, 16'd7995, 16'd63771, 16'd42214, 16'd52788, 16'd43633, 16'd40729, 16'd28099, 16'd42830, 16'd7235, 16'd6050, 16'd44949, 16'd26664, 16'd16998, 16'd62360, 16'd59020, 16'd23140, 16'd15503, 16'd41815, 16'd42203});
	test_expansion(128'hadb553ed2a59c5fecf61e06a4f2a008e, {16'd9523, 16'd52111, 16'd30176, 16'd17634, 16'd17055, 16'd21239, 16'd55902, 16'd60131, 16'd28532, 16'd64170, 16'd24082, 16'd2114, 16'd31793, 16'd30081, 16'd10810, 16'd16629, 16'd16802, 16'd61035, 16'd39343, 16'd21240, 16'd18035, 16'd5320, 16'd32165, 16'd18815, 16'd5927, 16'd54656});
	test_expansion(128'hfdcef2ef384894a9b5f287b114a060d2, {16'd62282, 16'd37724, 16'd54877, 16'd36813, 16'd39238, 16'd39290, 16'd19105, 16'd33194, 16'd12063, 16'd63333, 16'd47537, 16'd41400, 16'd10405, 16'd1227, 16'd54025, 16'd16793, 16'd686, 16'd24247, 16'd37557, 16'd42023, 16'd13223, 16'd18186, 16'd61096, 16'd42408, 16'd1893, 16'd18178});
	test_expansion(128'hdcace69f1c868b4bf33a3081a9162dc9, {16'd65023, 16'd41748, 16'd63173, 16'd18987, 16'd53582, 16'd23710, 16'd64321, 16'd13704, 16'd16485, 16'd59486, 16'd12819, 16'd8389, 16'd27375, 16'd65016, 16'd18019, 16'd21119, 16'd58307, 16'd5248, 16'd31074, 16'd41378, 16'd621, 16'd64725, 16'd15002, 16'd358, 16'd17144, 16'd35494});
	test_expansion(128'hbbb30ffb396d7c526477f6029af91187, {16'd55321, 16'd52211, 16'd2020, 16'd14542, 16'd62448, 16'd5294, 16'd19690, 16'd60310, 16'd46719, 16'd30153, 16'd5418, 16'd5792, 16'd51147, 16'd64804, 16'd13332, 16'd14616, 16'd2839, 16'd12397, 16'd43800, 16'd8184, 16'd46628, 16'd63012, 16'd15585, 16'd52325, 16'd7550, 16'd45325});
	test_expansion(128'hfc6e3ea011733575f1547fc1e128fa31, {16'd52667, 16'd48510, 16'd55829, 16'd28364, 16'd42721, 16'd22099, 16'd2200, 16'd27092, 16'd9761, 16'd51369, 16'd52224, 16'd44895, 16'd31846, 16'd62057, 16'd59351, 16'd46109, 16'd24988, 16'd61464, 16'd12009, 16'd4361, 16'd28167, 16'd54672, 16'd1752, 16'd35467, 16'd61358, 16'd3341});
	test_expansion(128'he0a7514ed639c1357c53eba375e393a9, {16'd23209, 16'd31707, 16'd59427, 16'd48178, 16'd33967, 16'd53322, 16'd3013, 16'd30165, 16'd62020, 16'd8665, 16'd53248, 16'd26907, 16'd51925, 16'd7004, 16'd11018, 16'd27222, 16'd5814, 16'd42733, 16'd16566, 16'd39206, 16'd14442, 16'd36403, 16'd31971, 16'd5724, 16'd43524, 16'd10552});
	test_expansion(128'hd1bbd920cafbc27c10c4be44df83c7c4, {16'd62365, 16'd25429, 16'd53768, 16'd8623, 16'd64837, 16'd12272, 16'd8438, 16'd58812, 16'd27376, 16'd44467, 16'd45906, 16'd45740, 16'd45305, 16'd28196, 16'd20655, 16'd54448, 16'd23370, 16'd1583, 16'd3529, 16'd17471, 16'd39268, 16'd22176, 16'd29841, 16'd51096, 16'd3710, 16'd56365});
	test_expansion(128'hd699fae3f51197e87187966eed06d22e, {16'd57550, 16'd20170, 16'd29139, 16'd34444, 16'd45972, 16'd60367, 16'd21195, 16'd50950, 16'd57200, 16'd60667, 16'd16878, 16'd3133, 16'd21968, 16'd49652, 16'd59414, 16'd28638, 16'd11082, 16'd32344, 16'd41413, 16'd33238, 16'd43223, 16'd55329, 16'd48069, 16'd14161, 16'd24888, 16'd35713});
	test_expansion(128'h9da7ec436ef435587b1da8583165b997, {16'd62549, 16'd26186, 16'd51486, 16'd61925, 16'd55308, 16'd24566, 16'd60673, 16'd36633, 16'd2782, 16'd59314, 16'd3181, 16'd55698, 16'd4440, 16'd46522, 16'd35815, 16'd49192, 16'd25009, 16'd61305, 16'd46748, 16'd22420, 16'd54142, 16'd26513, 16'd42681, 16'd29190, 16'd18533, 16'd58477});
	test_expansion(128'h2799e1f4e1d58f4504e438a0ebbdf0fa, {16'd6756, 16'd65503, 16'd42406, 16'd40223, 16'd51263, 16'd63327, 16'd6401, 16'd28049, 16'd32501, 16'd48012, 16'd55201, 16'd41316, 16'd37569, 16'd17284, 16'd63815, 16'd27504, 16'd36213, 16'd42793, 16'd52826, 16'd26476, 16'd56274, 16'd6152, 16'd44826, 16'd27912, 16'd63441, 16'd27444});
	test_expansion(128'h8491e86873d36962b659a56e64f38f1c, {16'd55272, 16'd54558, 16'd35598, 16'd29318, 16'd64266, 16'd27807, 16'd49602, 16'd50295, 16'd9139, 16'd32354, 16'd25126, 16'd59392, 16'd10553, 16'd30528, 16'd23893, 16'd30731, 16'd37692, 16'd43190, 16'd31485, 16'd30453, 16'd43962, 16'd9462, 16'd44874, 16'd62993, 16'd30499, 16'd52463});
	test_expansion(128'h736bbbdf9a56ffe6e8cd53b2f61645b8, {16'd60850, 16'd38657, 16'd39833, 16'd62126, 16'd4471, 16'd46448, 16'd46147, 16'd60656, 16'd51272, 16'd24655, 16'd50541, 16'd40097, 16'd1168, 16'd12742, 16'd34399, 16'd51665, 16'd31346, 16'd7840, 16'd59187, 16'd58117, 16'd20565, 16'd33009, 16'd55685, 16'd58477, 16'd21040, 16'd10486});
	test_expansion(128'hf3d261ebd3ea551ab812010a88f7c68a, {16'd1409, 16'd38332, 16'd55817, 16'd36495, 16'd64881, 16'd38466, 16'd2009, 16'd21063, 16'd43192, 16'd33792, 16'd63478, 16'd27365, 16'd4052, 16'd8318, 16'd52010, 16'd24040, 16'd61219, 16'd55139, 16'd58288, 16'd25080, 16'd25462, 16'd52196, 16'd6277, 16'd19930, 16'd45801, 16'd4565});
	test_expansion(128'h414cd05223927d13b6d163191f8139c6, {16'd5144, 16'd42196, 16'd48353, 16'd21652, 16'd5940, 16'd47585, 16'd48179, 16'd9288, 16'd49494, 16'd22647, 16'd49348, 16'd19825, 16'd28761, 16'd20487, 16'd58496, 16'd43849, 16'd42254, 16'd39702, 16'd43417, 16'd53154, 16'd57299, 16'd16432, 16'd12068, 16'd63014, 16'd18360, 16'd11786});
	test_expansion(128'h45ef58c2358ecd851b173bbec04b829e, {16'd33241, 16'd56457, 16'd37718, 16'd33917, 16'd33216, 16'd2105, 16'd42426, 16'd4751, 16'd4857, 16'd3223, 16'd20595, 16'd57211, 16'd45171, 16'd62356, 16'd52110, 16'd53376, 16'd64299, 16'd13233, 16'd54833, 16'd63707, 16'd17097, 16'd10570, 16'd64177, 16'd55127, 16'd22152, 16'd35974});
	test_expansion(128'hf8e236a861f51f2f14f3bafb127eb7eb, {16'd33475, 16'd43886, 16'd28031, 16'd43940, 16'd39727, 16'd31934, 16'd49016, 16'd60064, 16'd61500, 16'd29953, 16'd11734, 16'd12609, 16'd17663, 16'd55734, 16'd32893, 16'd5039, 16'd23785, 16'd60906, 16'd6903, 16'd47485, 16'd23885, 16'd62030, 16'd42639, 16'd55257, 16'd20778, 16'd53702});
	test_expansion(128'haee7aa86a6028cf1a00b30ceb909612a, {16'd3761, 16'd19671, 16'd29803, 16'd45758, 16'd50216, 16'd29378, 16'd34031, 16'd8205, 16'd34412, 16'd11283, 16'd496, 16'd45452, 16'd39190, 16'd10607, 16'd17600, 16'd63231, 16'd14196, 16'd184, 16'd45609, 16'd32967, 16'd61602, 16'd54565, 16'd40404, 16'd36999, 16'd12885, 16'd62672});
	test_expansion(128'h6cec08e6ed238be29a5f3eba269cd88c, {16'd11468, 16'd8448, 16'd36918, 16'd43205, 16'd61523, 16'd58400, 16'd41751, 16'd2074, 16'd49846, 16'd46568, 16'd64402, 16'd61121, 16'd47349, 16'd4487, 16'd10400, 16'd27498, 16'd49368, 16'd41884, 16'd45375, 16'd56698, 16'd9957, 16'd5531, 16'd64324, 16'd27012, 16'd40856, 16'd35493});
	test_expansion(128'hec7555bf5280170f2915f38603597df8, {16'd4942, 16'd65215, 16'd37924, 16'd49109, 16'd55311, 16'd3793, 16'd21232, 16'd35897, 16'd60147, 16'd59500, 16'd21575, 16'd65147, 16'd16667, 16'd51582, 16'd38291, 16'd62270, 16'd29441, 16'd65045, 16'd29612, 16'd8907, 16'd18340, 16'd4494, 16'd28943, 16'd9834, 16'd3760, 16'd45011});
	test_expansion(128'hf91970c9cc92e61511cc2cdc711802d7, {16'd20889, 16'd31171, 16'd29381, 16'd26351, 16'd32793, 16'd52568, 16'd3291, 16'd6933, 16'd37406, 16'd28447, 16'd2973, 16'd10899, 16'd51915, 16'd29502, 16'd8526, 16'd44112, 16'd26, 16'd45692, 16'd19574, 16'd37987, 16'd29212, 16'd27426, 16'd47477, 16'd63523, 16'd16146, 16'd285});
	test_expansion(128'h0ea56610dca828f28c755b79beec4485, {16'd63006, 16'd54707, 16'd33538, 16'd25986, 16'd23608, 16'd31953, 16'd26768, 16'd11499, 16'd31163, 16'd62534, 16'd39399, 16'd50925, 16'd31128, 16'd21978, 16'd57158, 16'd54741, 16'd39802, 16'd30138, 16'd1260, 16'd473, 16'd27944, 16'd945, 16'd22730, 16'd15325, 16'd60903, 16'd47663});
	test_expansion(128'h336ae68c4eb11d31bf1d7ad132631aa7, {16'd25207, 16'd20444, 16'd2957, 16'd63050, 16'd57362, 16'd57057, 16'd36512, 16'd5123, 16'd56371, 16'd40177, 16'd39712, 16'd3229, 16'd27378, 16'd47662, 16'd49928, 16'd5331, 16'd14380, 16'd5543, 16'd56147, 16'd45407, 16'd23588, 16'd40671, 16'd8620, 16'd53959, 16'd55515, 16'd17463});
	test_expansion(128'h31fdb86a7345126c20ebc9026d207338, {16'd55975, 16'd32807, 16'd64054, 16'd23655, 16'd46222, 16'd25973, 16'd6992, 16'd37925, 16'd42955, 16'd64637, 16'd27154, 16'd3065, 16'd3933, 16'd31596, 16'd1530, 16'd1895, 16'd62504, 16'd29920, 16'd13521, 16'd28909, 16'd65122, 16'd40209, 16'd56470, 16'd61232, 16'd59400, 16'd17838});
	test_expansion(128'h400e3d37968028e120cede19fe3d5763, {16'd11826, 16'd39016, 16'd51183, 16'd3311, 16'd28300, 16'd13581, 16'd10640, 16'd21149, 16'd51327, 16'd35968, 16'd45090, 16'd10386, 16'd27803, 16'd15696, 16'd29560, 16'd25973, 16'd45700, 16'd34039, 16'd33552, 16'd59063, 16'd1540, 16'd5653, 16'd56695, 16'd3873, 16'd30415, 16'd7846});
	test_expansion(128'hcd6c67815034fff2b7b415400dbfdd17, {16'd32500, 16'd3826, 16'd25690, 16'd6716, 16'd53756, 16'd10912, 16'd31409, 16'd10975, 16'd60265, 16'd20813, 16'd12459, 16'd54738, 16'd56318, 16'd760, 16'd42590, 16'd54683, 16'd12786, 16'd24470, 16'd7125, 16'd11845, 16'd43984, 16'd32973, 16'd35344, 16'd55580, 16'd56255, 16'd28205});
	test_expansion(128'h2d46978d2cfcc392f9f7bce888dd92f4, {16'd18446, 16'd22896, 16'd59799, 16'd57844, 16'd53041, 16'd1040, 16'd8405, 16'd14544, 16'd41151, 16'd19608, 16'd52829, 16'd8848, 16'd32336, 16'd65233, 16'd22429, 16'd44510, 16'd45862, 16'd1609, 16'd15763, 16'd60445, 16'd13203, 16'd46702, 16'd38497, 16'd30022, 16'd64301, 16'd57092});
	test_expansion(128'h7c68f6123a9ae8daedd395b7dcdfbab5, {16'd26536, 16'd56433, 16'd45852, 16'd57903, 16'd8174, 16'd23531, 16'd32630, 16'd54634, 16'd35603, 16'd12831, 16'd59535, 16'd36894, 16'd44780, 16'd58207, 16'd33004, 16'd5940, 16'd55783, 16'd62322, 16'd51728, 16'd34548, 16'd3408, 16'd65002, 16'd25865, 16'd32933, 16'd42402, 16'd697});
	test_expansion(128'hb81d2e6db07e99cf1eefae3707531741, {16'd33850, 16'd54447, 16'd36663, 16'd30836, 16'd4366, 16'd5077, 16'd14142, 16'd56850, 16'd2886, 16'd40332, 16'd2620, 16'd65010, 16'd19255, 16'd29413, 16'd39429, 16'd31273, 16'd42092, 16'd63593, 16'd52691, 16'd19940, 16'd23968, 16'd55029, 16'd40164, 16'd36597, 16'd9860, 16'd14239});
	test_expansion(128'h42a4306701b34d9d47878a7b8c6e4564, {16'd36624, 16'd50658, 16'd57305, 16'd33472, 16'd48170, 16'd20079, 16'd65123, 16'd55211, 16'd10012, 16'd46274, 16'd28187, 16'd62113, 16'd10731, 16'd6022, 16'd13024, 16'd15694, 16'd39221, 16'd43038, 16'd57550, 16'd38663, 16'd2380, 16'd62760, 16'd19754, 16'd12211, 16'd29952, 16'd44567});
	test_expansion(128'h2458625decdb69177126fca7b1f65d8b, {16'd31667, 16'd59038, 16'd61909, 16'd10172, 16'd2344, 16'd56656, 16'd29655, 16'd33732, 16'd3527, 16'd1129, 16'd56115, 16'd49644, 16'd28913, 16'd46704, 16'd44258, 16'd55321, 16'd31196, 16'd9388, 16'd19445, 16'd38829, 16'd44700, 16'd28327, 16'd33916, 16'd39996, 16'd30140, 16'd62319});
	test_expansion(128'h267aa18fee3e5f8606b6beb095b753ab, {16'd26766, 16'd28596, 16'd34881, 16'd20487, 16'd30828, 16'd49079, 16'd12108, 16'd16565, 16'd8883, 16'd9098, 16'd2981, 16'd15674, 16'd6269, 16'd12293, 16'd57966, 16'd30987, 16'd9413, 16'd60741, 16'd48402, 16'd38227, 16'd13606, 16'd18788, 16'd57610, 16'd50736, 16'd38022, 16'd50064});
	test_expansion(128'he069ac7a51a178943d10d018565d35f6, {16'd5069, 16'd57097, 16'd20060, 16'd39081, 16'd35499, 16'd7986, 16'd43980, 16'd12687, 16'd22170, 16'd24200, 16'd53275, 16'd49260, 16'd58578, 16'd35444, 16'd53817, 16'd34193, 16'd22496, 16'd53653, 16'd5662, 16'd32938, 16'd34649, 16'd24528, 16'd62679, 16'd29946, 16'd24681, 16'd35058});
	test_expansion(128'h4edf45d70ee70f1e6bc23cfa32f7ffa0, {16'd6009, 16'd27825, 16'd29105, 16'd35648, 16'd695, 16'd39910, 16'd49807, 16'd64264, 16'd29740, 16'd50135, 16'd50626, 16'd12878, 16'd59515, 16'd15102, 16'd10334, 16'd23747, 16'd50807, 16'd26656, 16'd59853, 16'd11495, 16'd47000, 16'd44610, 16'd25314, 16'd63743, 16'd16865, 16'd19933});
	test_expansion(128'hd4d8b7e55ab96fa569e156f27b93478c, {16'd42528, 16'd1723, 16'd39227, 16'd24580, 16'd45629, 16'd15190, 16'd58768, 16'd49563, 16'd9563, 16'd27662, 16'd25887, 16'd57893, 16'd17368, 16'd44837, 16'd51652, 16'd34508, 16'd57399, 16'd609, 16'd15151, 16'd60588, 16'd25576, 16'd33807, 16'd23325, 16'd35751, 16'd16913, 16'd59441});
	test_expansion(128'heaecb50dc360516fce62c9d0156a4f5f, {16'd48975, 16'd42056, 16'd40234, 16'd53453, 16'd64492, 16'd41544, 16'd57153, 16'd29798, 16'd50720, 16'd39946, 16'd43433, 16'd3433, 16'd58599, 16'd23704, 16'd27050, 16'd29434, 16'd36040, 16'd10083, 16'd63980, 16'd49369, 16'd36171, 16'd57149, 16'd3190, 16'd60313, 16'd60508, 16'd43418});
	test_expansion(128'he8e2af477cd15deeb66ff8dbcb11a56a, {16'd2827, 16'd29079, 16'd41912, 16'd41854, 16'd12196, 16'd18477, 16'd33587, 16'd15499, 16'd20585, 16'd53988, 16'd26424, 16'd10923, 16'd56038, 16'd40259, 16'd8544, 16'd1864, 16'd18805, 16'd4799, 16'd44908, 16'd20753, 16'd59148, 16'd7582, 16'd22507, 16'd54859, 16'd38425, 16'd48125});
	test_expansion(128'hee83effcbd8db688123059e22a795057, {16'd8526, 16'd46250, 16'd46709, 16'd64502, 16'd6212, 16'd7700, 16'd23453, 16'd35015, 16'd1526, 16'd24416, 16'd46559, 16'd2835, 16'd52293, 16'd5172, 16'd54835, 16'd63903, 16'd19990, 16'd60148, 16'd33616, 16'd42874, 16'd13621, 16'd5392, 16'd23274, 16'd56133, 16'd64073, 16'd29777});
	test_expansion(128'hd37799c3c0810dea58497a849df7439c, {16'd15156, 16'd6330, 16'd14967, 16'd33349, 16'd685, 16'd8988, 16'd22423, 16'd26811, 16'd53969, 16'd59015, 16'd45365, 16'd4046, 16'd7471, 16'd63865, 16'd1610, 16'd26674, 16'd24265, 16'd46648, 16'd60081, 16'd35630, 16'd46078, 16'd23959, 16'd17639, 16'd45427, 16'd40777, 16'd3586});
	test_expansion(128'hfe90bd7f07f9e0386415338ed51c171e, {16'd8009, 16'd27433, 16'd20742, 16'd39884, 16'd33180, 16'd35926, 16'd18579, 16'd63806, 16'd10965, 16'd9784, 16'd33239, 16'd26722, 16'd39876, 16'd31770, 16'd21931, 16'd37889, 16'd27583, 16'd27555, 16'd40209, 16'd23235, 16'd5491, 16'd65182, 16'd59157, 16'd30814, 16'd53361, 16'd39401});
	test_expansion(128'hd7b41334c4cc0ac1b822da46561b0416, {16'd63799, 16'd55252, 16'd62269, 16'd1229, 16'd55839, 16'd60001, 16'd1870, 16'd60520, 16'd27727, 16'd5814, 16'd57209, 16'd23702, 16'd65414, 16'd4585, 16'd18936, 16'd11098, 16'd48263, 16'd18974, 16'd47185, 16'd33234, 16'd43275, 16'd34628, 16'd11622, 16'd43819, 16'd32082, 16'd11197});
	test_expansion(128'h78c86d0185e3bc9deb89f15fdbb16fd1, {16'd59226, 16'd8243, 16'd50945, 16'd15719, 16'd44900, 16'd32840, 16'd52596, 16'd15791, 16'd49924, 16'd17595, 16'd44920, 16'd53946, 16'd19807, 16'd52108, 16'd4908, 16'd3111, 16'd345, 16'd24973, 16'd4077, 16'd10792, 16'd7471, 16'd27893, 16'd3836, 16'd54193, 16'd19974, 16'd15716});
	test_expansion(128'h844e94ff8337d74d1efbae437a306e03, {16'd20551, 16'd54463, 16'd25357, 16'd24021, 16'd56504, 16'd20453, 16'd43006, 16'd49959, 16'd6772, 16'd37999, 16'd23664, 16'd54681, 16'd45465, 16'd54934, 16'd51967, 16'd38621, 16'd36723, 16'd32018, 16'd53911, 16'd50809, 16'd6379, 16'd2421, 16'd49297, 16'd58211, 16'd21674, 16'd35269});
	test_expansion(128'h6a9b5f4d0c34f131eaf7c9e6046b8f70, {16'd9321, 16'd57995, 16'd62881, 16'd5548, 16'd58646, 16'd55179, 16'd7017, 16'd26708, 16'd13166, 16'd14729, 16'd6741, 16'd43571, 16'd26624, 16'd5366, 16'd32538, 16'd51499, 16'd25473, 16'd36558, 16'd63058, 16'd42252, 16'd592, 16'd14448, 16'd1888, 16'd53899, 16'd31652, 16'd49951});
	test_expansion(128'h8d84e8c8659fe063e48b772b1bdc39c2, {16'd1358, 16'd58579, 16'd21334, 16'd10842, 16'd39748, 16'd965, 16'd50303, 16'd63014, 16'd35505, 16'd26431, 16'd50161, 16'd48020, 16'd43898, 16'd39277, 16'd50073, 16'd39200, 16'd32708, 16'd17202, 16'd12209, 16'd36225, 16'd2086, 16'd64740, 16'd29607, 16'd13435, 16'd20849, 16'd49070});
	test_expansion(128'h42cb5182acd51c5dcd045239d7d9fade, {16'd19849, 16'd62145, 16'd57787, 16'd61972, 16'd6451, 16'd47828, 16'd22328, 16'd48327, 16'd50390, 16'd16727, 16'd55713, 16'd61671, 16'd61631, 16'd35878, 16'd26666, 16'd50036, 16'd52194, 16'd6347, 16'd45437, 16'd28886, 16'd63183, 16'd44170, 16'd36996, 16'd40612, 16'd49900, 16'd48188});
	test_expansion(128'h65ef8ebb0bf305fb76e892ee9bdd2a79, {16'd2732, 16'd37787, 16'd14101, 16'd13549, 16'd27693, 16'd31702, 16'd38512, 16'd19347, 16'd2946, 16'd29657, 16'd19334, 16'd29367, 16'd25770, 16'd53024, 16'd23280, 16'd57472, 16'd4785, 16'd48070, 16'd52265, 16'd21496, 16'd51851, 16'd55344, 16'd49244, 16'd11483, 16'd15655, 16'd11806});
	test_expansion(128'h7ed817fb578b4f63f3863692e0b5fb82, {16'd17772, 16'd28462, 16'd1570, 16'd58841, 16'd28258, 16'd26394, 16'd23445, 16'd50911, 16'd26887, 16'd30432, 16'd23181, 16'd6698, 16'd25099, 16'd153, 16'd49027, 16'd40416, 16'd38909, 16'd32722, 16'd16724, 16'd62114, 16'd60030, 16'd45459, 16'd3416, 16'd38933, 16'd2177, 16'd7550});
	test_expansion(128'h22aa0872c776769ced4124b7357aa4b9, {16'd14390, 16'd10371, 16'd2963, 16'd28284, 16'd51839, 16'd14388, 16'd8928, 16'd34921, 16'd62219, 16'd4015, 16'd49328, 16'd45586, 16'd1460, 16'd27993, 16'd9397, 16'd4449, 16'd36989, 16'd36795, 16'd13454, 16'd42601, 16'd42821, 16'd54156, 16'd24123, 16'd769, 16'd21702, 16'd57877});
	test_expansion(128'h2aa20aa9ddd1aadb7045f0daa3c8576a, {16'd23877, 16'd59900, 16'd4331, 16'd1579, 16'd8905, 16'd41166, 16'd23226, 16'd37058, 16'd25402, 16'd31094, 16'd58096, 16'd21918, 16'd9473, 16'd28571, 16'd39731, 16'd27301, 16'd43957, 16'd39494, 16'd51624, 16'd41813, 16'd33468, 16'd43885, 16'd48853, 16'd61312, 16'd18670, 16'd35538});
	test_expansion(128'he006da7d84370d5f69d67d52f3594a50, {16'd13014, 16'd36585, 16'd37981, 16'd6599, 16'd32457, 16'd9917, 16'd54697, 16'd10034, 16'd44187, 16'd49899, 16'd19187, 16'd34510, 16'd28130, 16'd53596, 16'd59938, 16'd49793, 16'd46974, 16'd45673, 16'd9062, 16'd8607, 16'd19144, 16'd49796, 16'd25688, 16'd50316, 16'd39602, 16'd42456});
	test_expansion(128'hea4a6880765da2570b2ada583d00bd00, {16'd38806, 16'd47155, 16'd53874, 16'd12789, 16'd50142, 16'd19847, 16'd17829, 16'd30000, 16'd20880, 16'd24017, 16'd59206, 16'd59127, 16'd60061, 16'd53892, 16'd14769, 16'd37245, 16'd47064, 16'd47837, 16'd7637, 16'd54441, 16'd11274, 16'd15090, 16'd63419, 16'd34293, 16'd18010, 16'd22843});
	test_expansion(128'h347749eae5e45eb74683a5bad509dcd6, {16'd53610, 16'd63670, 16'd34357, 16'd50197, 16'd26451, 16'd28785, 16'd26162, 16'd19587, 16'd1801, 16'd7992, 16'd41573, 16'd33703, 16'd23027, 16'd48043, 16'd47027, 16'd27020, 16'd34126, 16'd24988, 16'd52431, 16'd24786, 16'd18046, 16'd28320, 16'd45682, 16'd61441, 16'd62999, 16'd10382});
	test_expansion(128'h0f7db6801e2ac6098d41a5fd22754cf4, {16'd44565, 16'd33698, 16'd17896, 16'd34172, 16'd44591, 16'd7049, 16'd21289, 16'd22173, 16'd11192, 16'd15283, 16'd29959, 16'd36245, 16'd17947, 16'd5103, 16'd20194, 16'd65255, 16'd45794, 16'd38047, 16'd21464, 16'd8279, 16'd57141, 16'd15752, 16'd44525, 16'd11667, 16'd45642, 16'd4032});
	test_expansion(128'h8588b47e2b223aba7ecfd5842ec54574, {16'd4178, 16'd47413, 16'd31366, 16'd11725, 16'd32572, 16'd53923, 16'd50572, 16'd54536, 16'd54175, 16'd6250, 16'd42178, 16'd8782, 16'd56713, 16'd55081, 16'd12851, 16'd30028, 16'd31995, 16'd65371, 16'd44777, 16'd31147, 16'd13840, 16'd63667, 16'd32999, 16'd24859, 16'd4848, 16'd25734});
	test_expansion(128'h6489002780350f88f767dc15bc1f5e1e, {16'd27243, 16'd42956, 16'd1675, 16'd21312, 16'd35456, 16'd53189, 16'd1398, 16'd12651, 16'd17140, 16'd47055, 16'd51008, 16'd23571, 16'd885, 16'd13179, 16'd3125, 16'd49043, 16'd53187, 16'd50995, 16'd54736, 16'd47050, 16'd6792, 16'd42812, 16'd21422, 16'd16772, 16'd32556, 16'd49286});
	test_expansion(128'ha5cec442a8d050e3dc97d1e784e3a032, {16'd29203, 16'd45653, 16'd10825, 16'd20558, 16'd34830, 16'd18739, 16'd5810, 16'd64841, 16'd1745, 16'd53067, 16'd24151, 16'd35289, 16'd64431, 16'd28299, 16'd50431, 16'd54449, 16'd53562, 16'd43687, 16'd14948, 16'd3940, 16'd61922, 16'd49763, 16'd48566, 16'd32486, 16'd26845, 16'd59458});
	test_expansion(128'h3c3b752238e7e1d3d35fe0ad6b391c33, {16'd52787, 16'd26408, 16'd62613, 16'd44155, 16'd34531, 16'd40530, 16'd43466, 16'd36728, 16'd55055, 16'd20439, 16'd6412, 16'd60223, 16'd34558, 16'd52491, 16'd48632, 16'd37051, 16'd31128, 16'd1420, 16'd12285, 16'd12868, 16'd53485, 16'd27526, 16'd62780, 16'd3763, 16'd19715, 16'd9476});
	test_expansion(128'hb0a2fefd8ee67ef2868bc3b68d1f21f6, {16'd56067, 16'd49318, 16'd26284, 16'd20451, 16'd16552, 16'd16797, 16'd6352, 16'd44391, 16'd12196, 16'd6694, 16'd3145, 16'd39428, 16'd32847, 16'd54613, 16'd62004, 16'd2008, 16'd39930, 16'd49232, 16'd19714, 16'd54527, 16'd3859, 16'd907, 16'd7556, 16'd16994, 16'd35254, 16'd4180});
	test_expansion(128'hdff06ca0301e50c1ad5155c86a232b90, {16'd59410, 16'd24479, 16'd19543, 16'd51307, 16'd59302, 16'd19424, 16'd18383, 16'd5668, 16'd23940, 16'd54650, 16'd530, 16'd15610, 16'd20868, 16'd32532, 16'd5335, 16'd59987, 16'd39764, 16'd51551, 16'd12460, 16'd44494, 16'd7246, 16'd38326, 16'd9377, 16'd60608, 16'd2931, 16'd55177});
	test_expansion(128'hde06f5a954cec523705b2722a50dedfe, {16'd8900, 16'd25018, 16'd27199, 16'd14661, 16'd45750, 16'd15512, 16'd826, 16'd21891, 16'd62536, 16'd41063, 16'd44041, 16'd3227, 16'd29288, 16'd24602, 16'd1190, 16'd48010, 16'd9620, 16'd27681, 16'd55197, 16'd59253, 16'd29312, 16'd42829, 16'd4186, 16'd41803, 16'd8238, 16'd8778});
	test_expansion(128'h95785bf02b2da49e71f815213406ae68, {16'd44635, 16'd57760, 16'd1233, 16'd54569, 16'd39105, 16'd52177, 16'd20192, 16'd21498, 16'd35676, 16'd7909, 16'd16999, 16'd51272, 16'd37483, 16'd27731, 16'd39623, 16'd1172, 16'd18240, 16'd7852, 16'd22474, 16'd37768, 16'd26130, 16'd59964, 16'd63630, 16'd6832, 16'd13419, 16'd19747});
	test_expansion(128'h6c522cbafeaf6f1b614e90cfc09e0d33, {16'd34883, 16'd17270, 16'd43108, 16'd5115, 16'd41747, 16'd24755, 16'd25027, 16'd9765, 16'd61838, 16'd906, 16'd31758, 16'd1919, 16'd30340, 16'd45561, 16'd59046, 16'd25502, 16'd41696, 16'd11986, 16'd47260, 16'd43527, 16'd36230, 16'd10398, 16'd56461, 16'd40186, 16'd42868, 16'd7876});
	test_expansion(128'hbbc7ab08df770a65de0f831ae767a403, {16'd44157, 16'd38072, 16'd20509, 16'd22051, 16'd59369, 16'd52383, 16'd47190, 16'd43290, 16'd43714, 16'd42274, 16'd31889, 16'd40105, 16'd58585, 16'd7418, 16'd1027, 16'd30990, 16'd6934, 16'd27161, 16'd50128, 16'd4084, 16'd6467, 16'd22616, 16'd34956, 16'd2780, 16'd63057, 16'd21728});
	test_expansion(128'h45eee0e6afb0f09d33828ccc67179fde, {16'd44934, 16'd16423, 16'd60008, 16'd18505, 16'd64214, 16'd33659, 16'd35385, 16'd40432, 16'd6188, 16'd22490, 16'd49866, 16'd57143, 16'd34096, 16'd40931, 16'd11146, 16'd42402, 16'd15528, 16'd31559, 16'd4671, 16'd36182, 16'd63150, 16'd34299, 16'd3947, 16'd61658, 16'd58080, 16'd61061});
	test_expansion(128'h215a0758b36d6dae4ef0a16ae1c13753, {16'd49471, 16'd1123, 16'd54584, 16'd17200, 16'd44964, 16'd37398, 16'd48509, 16'd24058, 16'd2468, 16'd33900, 16'd22008, 16'd19761, 16'd356, 16'd63209, 16'd30129, 16'd50680, 16'd4902, 16'd34187, 16'd55217, 16'd42836, 16'd35914, 16'd54529, 16'd53112, 16'd27263, 16'd59636, 16'd25575});
	test_expansion(128'h78ad1a8d39f92b5a8cddb1c42bd4fe3f, {16'd44518, 16'd26329, 16'd30153, 16'd34640, 16'd10477, 16'd33745, 16'd13805, 16'd61835, 16'd12022, 16'd5508, 16'd34124, 16'd20616, 16'd35071, 16'd19095, 16'd17946, 16'd22634, 16'd63394, 16'd18036, 16'd33676, 16'd48223, 16'd44555, 16'd56927, 16'd48738, 16'd6462, 16'd32062, 16'd50878});
	test_expansion(128'h774718649b1bd348da5e9c1b51238594, {16'd50171, 16'd5579, 16'd10251, 16'd4384, 16'd62169, 16'd1774, 16'd33357, 16'd59410, 16'd16209, 16'd28120, 16'd20876, 16'd8876, 16'd8745, 16'd3263, 16'd27499, 16'd43927, 16'd25446, 16'd61206, 16'd4519, 16'd45587, 16'd21857, 16'd4806, 16'd54177, 16'd19584, 16'd65095, 16'd33068});
	test_expansion(128'hbc200fcbc0d8a796b0171d77d5783af9, {16'd24575, 16'd20851, 16'd56180, 16'd22532, 16'd18229, 16'd50053, 16'd45447, 16'd25388, 16'd33695, 16'd50939, 16'd13300, 16'd63728, 16'd21689, 16'd58995, 16'd2280, 16'd60179, 16'd41125, 16'd38932, 16'd27002, 16'd15594, 16'd41233, 16'd15991, 16'd24839, 16'd25067, 16'd39063, 16'd7320});
	test_expansion(128'hab59ef193014cb0de1e0d813d6dd47e2, {16'd58072, 16'd28575, 16'd63880, 16'd36090, 16'd31761, 16'd29037, 16'd12672, 16'd25985, 16'd44655, 16'd19200, 16'd62403, 16'd32597, 16'd34980, 16'd17607, 16'd60051, 16'd39013, 16'd11482, 16'd27622, 16'd2480, 16'd27487, 16'd54635, 16'd505, 16'd30412, 16'd7163, 16'd2432, 16'd13867});
	test_expansion(128'h19f35eb2914b1a0f4f9cb05a8f7467a7, {16'd44679, 16'd24007, 16'd54605, 16'd12342, 16'd29423, 16'd39640, 16'd28216, 16'd55917, 16'd7599, 16'd44922, 16'd39185, 16'd22004, 16'd8380, 16'd8008, 16'd63836, 16'd19472, 16'd10480, 16'd5714, 16'd24680, 16'd2899, 16'd58196, 16'd24204, 16'd57680, 16'd21310, 16'd27228, 16'd51981});
	test_expansion(128'ha20e38e23964b231ce03e3507390e4f1, {16'd62303, 16'd53861, 16'd39515, 16'd30369, 16'd6421, 16'd43402, 16'd41310, 16'd37817, 16'd61563, 16'd43858, 16'd22998, 16'd60359, 16'd12184, 16'd38698, 16'd40704, 16'd42165, 16'd49208, 16'd35989, 16'd64929, 16'd19759, 16'd56731, 16'd36917, 16'd41780, 16'd39262, 16'd44799, 16'd50060});
	test_expansion(128'h2f2172827cacc5cedf58f716737726bd, {16'd12663, 16'd63291, 16'd31335, 16'd2853, 16'd60704, 16'd55579, 16'd52323, 16'd60396, 16'd4868, 16'd42439, 16'd19892, 16'd2487, 16'd14306, 16'd60614, 16'd55438, 16'd15044, 16'd16755, 16'd30827, 16'd26685, 16'd29245, 16'd58973, 16'd13751, 16'd32480, 16'd53331, 16'd44363, 16'd27440});
	test_expansion(128'hab63b79071a6084dcd3c6b3d37b9a399, {16'd41118, 16'd34456, 16'd35099, 16'd41766, 16'd41110, 16'd18180, 16'd35888, 16'd22237, 16'd19862, 16'd26061, 16'd64882, 16'd42738, 16'd56907, 16'd46417, 16'd19443, 16'd40760, 16'd30707, 16'd44024, 16'd64302, 16'd52800, 16'd65130, 16'd64096, 16'd22668, 16'd63261, 16'd913, 16'd63852});
	test_expansion(128'he4d8d5b0fbb3299aadfcb61d3f14abbe, {16'd52187, 16'd41306, 16'd48693, 16'd40769, 16'd31128, 16'd24737, 16'd18519, 16'd3475, 16'd15243, 16'd848, 16'd52723, 16'd15030, 16'd26764, 16'd9595, 16'd39104, 16'd53860, 16'd7785, 16'd8721, 16'd38275, 16'd9915, 16'd52124, 16'd17290, 16'd48938, 16'd41441, 16'd3679, 16'd37593});
	test_expansion(128'hb11eea7bee2be24f608915043d52a64f, {16'd12073, 16'd39718, 16'd41095, 16'd63930, 16'd11594, 16'd63835, 16'd20943, 16'd46602, 16'd24597, 16'd45488, 16'd34043, 16'd18485, 16'd7859, 16'd37827, 16'd28217, 16'd9857, 16'd41034, 16'd28862, 16'd12346, 16'd52899, 16'd48988, 16'd35043, 16'd5037, 16'd21481, 16'd35638, 16'd37232});
	test_expansion(128'hdbb29304271c30c3d6cfbcb98039d32a, {16'd3278, 16'd29019, 16'd6949, 16'd17189, 16'd44119, 16'd43510, 16'd35256, 16'd50200, 16'd12623, 16'd31203, 16'd9248, 16'd59519, 16'd58765, 16'd2361, 16'd46568, 16'd25108, 16'd39285, 16'd2611, 16'd13819, 16'd30597, 16'd19438, 16'd8480, 16'd11021, 16'd27794, 16'd25274, 16'd2717});
	test_expansion(128'h6bf311ea869da6d0d68aca1f9aa76e91, {16'd49645, 16'd62426, 16'd38092, 16'd12920, 16'd13795, 16'd54944, 16'd48860, 16'd36380, 16'd6034, 16'd64244, 16'd63853, 16'd33936, 16'd11575, 16'd41383, 16'd17817, 16'd12136, 16'd38292, 16'd33967, 16'd6629, 16'd14155, 16'd59761, 16'd52363, 16'd45939, 16'd31464, 16'd13334, 16'd45194});
	test_expansion(128'hdc5fa2d831a77c662c10f91b53d518a1, {16'd35511, 16'd19467, 16'd13071, 16'd1188, 16'd24683, 16'd18348, 16'd13257, 16'd2816, 16'd22750, 16'd1134, 16'd15279, 16'd41299, 16'd27007, 16'd31820, 16'd40488, 16'd8695, 16'd62947, 16'd703, 16'd64528, 16'd46315, 16'd59084, 16'd38561, 16'd5123, 16'd53885, 16'd15503, 16'd36060});
	test_expansion(128'h6d12ca882b68be396bddb127e9d1e2b7, {16'd50433, 16'd57196, 16'd33187, 16'd12856, 16'd7192, 16'd38991, 16'd32651, 16'd32257, 16'd49925, 16'd22031, 16'd35719, 16'd12534, 16'd22628, 16'd42617, 16'd18206, 16'd63039, 16'd57136, 16'd19478, 16'd39937, 16'd28108, 16'd50736, 16'd49893, 16'd11406, 16'd37142, 16'd62248, 16'd27499});
	test_expansion(128'hb118e0a75431b68063d7ce33541cd168, {16'd10862, 16'd33029, 16'd14135, 16'd64552, 16'd50241, 16'd51327, 16'd22113, 16'd9475, 16'd2503, 16'd20667, 16'd53239, 16'd13980, 16'd27801, 16'd41740, 16'd45520, 16'd53083, 16'd54963, 16'd16480, 16'd33618, 16'd35450, 16'd56336, 16'd11265, 16'd59210, 16'd30190, 16'd22941, 16'd60070});
	test_expansion(128'h14fba124e0d2944763ade196f8dca6c9, {16'd46242, 16'd49256, 16'd49061, 16'd740, 16'd25558, 16'd29836, 16'd20637, 16'd37833, 16'd19393, 16'd39876, 16'd32968, 16'd42030, 16'd56570, 16'd37946, 16'd62716, 16'd1457, 16'd30779, 16'd33582, 16'd28778, 16'd26718, 16'd9068, 16'd31901, 16'd18490, 16'd17226, 16'd64576, 16'd41045});
	test_expansion(128'hd3428c6a610d4a578a85e91a422fc103, {16'd59743, 16'd11661, 16'd32838, 16'd41063, 16'd16118, 16'd64853, 16'd42540, 16'd48235, 16'd22126, 16'd673, 16'd28554, 16'd32540, 16'd51241, 16'd26798, 16'd31814, 16'd1110, 16'd13601, 16'd40861, 16'd5119, 16'd33402, 16'd64876, 16'd56250, 16'd59360, 16'd47846, 16'd57707, 16'd47832});
	test_expansion(128'h53ec9d452d4ac1a05ed7d99e2e9677b0, {16'd18565, 16'd381, 16'd62791, 16'd4537, 16'd26143, 16'd16406, 16'd18798, 16'd34060, 16'd36052, 16'd55467, 16'd9957, 16'd24218, 16'd13225, 16'd64168, 16'd30397, 16'd2788, 16'd41478, 16'd58848, 16'd32004, 16'd22961, 16'd7733, 16'd5521, 16'd46280, 16'd25617, 16'd40536, 16'd10538});
	test_expansion(128'hcaa0b870eca65044453cf4b1365375f3, {16'd63259, 16'd29962, 16'd41643, 16'd22734, 16'd39620, 16'd34410, 16'd7204, 16'd1487, 16'd2417, 16'd22529, 16'd30589, 16'd8190, 16'd41213, 16'd29510, 16'd59408, 16'd36437, 16'd22816, 16'd17717, 16'd38303, 16'd5637, 16'd12115, 16'd26335, 16'd35946, 16'd14889, 16'd24732, 16'd27557});
	test_expansion(128'h0b43d2c7a1a58785ac38749f317eec45, {16'd30788, 16'd34756, 16'd41453, 16'd54077, 16'd58516, 16'd6481, 16'd22994, 16'd26910, 16'd4449, 16'd9940, 16'd815, 16'd26644, 16'd25484, 16'd34275, 16'd52346, 16'd29046, 16'd23361, 16'd4534, 16'd43659, 16'd40239, 16'd61833, 16'd52988, 16'd59611, 16'd61836, 16'd44512, 16'd53354});
	test_expansion(128'h7e13f8540b89cc97f3bf42bcac976056, {16'd32175, 16'd28755, 16'd53087, 16'd16574, 16'd27576, 16'd51869, 16'd46790, 16'd38886, 16'd55501, 16'd27456, 16'd62625, 16'd8782, 16'd22791, 16'd35487, 16'd51643, 16'd4646, 16'd52755, 16'd57323, 16'd56593, 16'd39429, 16'd17948, 16'd23694, 16'd36756, 16'd13479, 16'd12697, 16'd48617});
	test_expansion(128'hc7c360a85c1f352cc26000185069240d, {16'd26327, 16'd37581, 16'd20676, 16'd34230, 16'd54715, 16'd6262, 16'd60031, 16'd6460, 16'd2846, 16'd60836, 16'd62133, 16'd57797, 16'd61825, 16'd4948, 16'd10262, 16'd12661, 16'd33571, 16'd39036, 16'd41064, 16'd14472, 16'd28232, 16'd43721, 16'd42912, 16'd39317, 16'd64576, 16'd1551});
	test_expansion(128'h36b0dd271d6aed7d1e032629e0664f48, {16'd58549, 16'd43560, 16'd17643, 16'd7760, 16'd26438, 16'd65343, 16'd28354, 16'd16328, 16'd20099, 16'd2898, 16'd29646, 16'd14543, 16'd20, 16'd33461, 16'd9537, 16'd39747, 16'd897, 16'd17597, 16'd53214, 16'd47265, 16'd737, 16'd60914, 16'd52594, 16'd4923, 16'd1333, 16'd34899});
	test_expansion(128'h87143f4f337bf2c11466fd2b635dc64f, {16'd31156, 16'd12386, 16'd49126, 16'd4915, 16'd61783, 16'd20003, 16'd24271, 16'd11761, 16'd51436, 16'd29052, 16'd60853, 16'd16300, 16'd44889, 16'd60553, 16'd60406, 16'd53587, 16'd48882, 16'd26805, 16'd50445, 16'd56667, 16'd11945, 16'd14307, 16'd37687, 16'd62183, 16'd55410, 16'd24261});
	test_expansion(128'he46267b81d96255a3563570bbe01263a, {16'd18973, 16'd35188, 16'd1491, 16'd27429, 16'd55215, 16'd59165, 16'd22991, 16'd8004, 16'd6312, 16'd17210, 16'd59339, 16'd19147, 16'd46386, 16'd63289, 16'd35043, 16'd14723, 16'd32339, 16'd43742, 16'd27117, 16'd47367, 16'd53658, 16'd913, 16'd31818, 16'd345, 16'd3033, 16'd56796});
	test_expansion(128'ha03052f24b16e0c27b4a734e9e069078, {16'd54104, 16'd33997, 16'd56162, 16'd55857, 16'd23340, 16'd563, 16'd63665, 16'd62415, 16'd599, 16'd310, 16'd23614, 16'd16409, 16'd29034, 16'd26505, 16'd31349, 16'd22414, 16'd14614, 16'd53245, 16'd9260, 16'd36910, 16'd47254, 16'd53567, 16'd57316, 16'd1922, 16'd5783, 16'd5775});
	test_expansion(128'he15a81454c889a23ad118c9fe24e41ad, {16'd50959, 16'd31776, 16'd13962, 16'd57441, 16'd45028, 16'd54530, 16'd37773, 16'd5585, 16'd59467, 16'd22242, 16'd46339, 16'd53125, 16'd43090, 16'd50903, 16'd63623, 16'd31920, 16'd60137, 16'd1020, 16'd16763, 16'd28301, 16'd28085, 16'd2189, 16'd44597, 16'd53236, 16'd63923, 16'd58437});
	test_expansion(128'h7a1134d04d0e5d8f236f89c9f0363b5f, {16'd58597, 16'd30497, 16'd34162, 16'd51936, 16'd34771, 16'd63442, 16'd47046, 16'd17878, 16'd37774, 16'd36904, 16'd8177, 16'd46917, 16'd54752, 16'd20097, 16'd25847, 16'd65007, 16'd32823, 16'd22430, 16'd1310, 16'd5680, 16'd45480, 16'd7181, 16'd24307, 16'd4401, 16'd42330, 16'd14402});
	test_expansion(128'ha40f8aaad9eca21b23510e3cf4c01464, {16'd13866, 16'd40132, 16'd24482, 16'd54963, 16'd5532, 16'd36793, 16'd34183, 16'd6648, 16'd33755, 16'd55478, 16'd49701, 16'd4716, 16'd57030, 16'd9540, 16'd58921, 16'd24710, 16'd43649, 16'd59427, 16'd2459, 16'd40952, 16'd40433, 16'd40731, 16'd32299, 16'd50729, 16'd64881, 16'd21002});
	test_expansion(128'hca79d142603497f70572fd6d09b9407a, {16'd47202, 16'd40993, 16'd27685, 16'd64434, 16'd59799, 16'd2926, 16'd22117, 16'd64454, 16'd700, 16'd65451, 16'd63110, 16'd46999, 16'd34819, 16'd4137, 16'd63912, 16'd7645, 16'd61854, 16'd12832, 16'd49562, 16'd2969, 16'd4500, 16'd24020, 16'd28835, 16'd43646, 16'd56680, 16'd33639});
	test_expansion(128'h09eb00ba154916b5254f893be61b9d86, {16'd39818, 16'd6624, 16'd26802, 16'd19905, 16'd44636, 16'd13494, 16'd40233, 16'd53474, 16'd35024, 16'd63128, 16'd36885, 16'd47487, 16'd50983, 16'd26961, 16'd4651, 16'd33034, 16'd31581, 16'd58976, 16'd26235, 16'd10912, 16'd32659, 16'd53204, 16'd38605, 16'd19416, 16'd42988, 16'd969});
	test_expansion(128'hdc4911a4b2a39021bc428da7b5282ba2, {16'd52520, 16'd41551, 16'd57747, 16'd38929, 16'd31861, 16'd4431, 16'd61522, 16'd59711, 16'd19806, 16'd61463, 16'd59844, 16'd11136, 16'd62256, 16'd31278, 16'd27150, 16'd5890, 16'd2615, 16'd30638, 16'd23547, 16'd3958, 16'd31040, 16'd20643, 16'd39663, 16'd36435, 16'd61857, 16'd50874});
	test_expansion(128'he030c3e756631a95c482a5519d04a59f, {16'd63603, 16'd9316, 16'd12432, 16'd2607, 16'd49847, 16'd3736, 16'd38668, 16'd49009, 16'd33203, 16'd26382, 16'd64079, 16'd53934, 16'd31582, 16'd56029, 16'd45690, 16'd379, 16'd6072, 16'd31809, 16'd11808, 16'd58745, 16'd55920, 16'd7681, 16'd32091, 16'd59314, 16'd58873, 16'd41192});
	test_expansion(128'hc1d43ec2d9dac44fbbfbece1e00f6c83, {16'd47127, 16'd11057, 16'd40212, 16'd21460, 16'd6075, 16'd35525, 16'd48502, 16'd36987, 16'd3037, 16'd23388, 16'd45930, 16'd3735, 16'd60143, 16'd5975, 16'd51496, 16'd45222, 16'd47369, 16'd21014, 16'd40489, 16'd1637, 16'd42955, 16'd41274, 16'd27951, 16'd28568, 16'd36642, 16'd36988});
	test_expansion(128'h26a74d884375e4e688ddaa34a0cfa955, {16'd53757, 16'd60104, 16'd13292, 16'd23629, 16'd14583, 16'd13491, 16'd2647, 16'd7318, 16'd60186, 16'd36265, 16'd23824, 16'd9930, 16'd57177, 16'd14875, 16'd51195, 16'd57919, 16'd9147, 16'd40198, 16'd13711, 16'd56658, 16'd53850, 16'd33752, 16'd58797, 16'd23816, 16'd55646, 16'd846});
	test_expansion(128'hda940b06dbbfccd86bac536c339ff601, {16'd9395, 16'd40444, 16'd20378, 16'd30921, 16'd32698, 16'd64602, 16'd14365, 16'd64885, 16'd28671, 16'd39025, 16'd51925, 16'd22366, 16'd12834, 16'd2620, 16'd54270, 16'd3502, 16'd42932, 16'd30440, 16'd10126, 16'd56388, 16'd39690, 16'd23315, 16'd20607, 16'd15020, 16'd31967, 16'd45324});
	test_expansion(128'hac0de5a4addf2027c3a1e48fedff23bf, {16'd25009, 16'd40283, 16'd59321, 16'd12612, 16'd41775, 16'd49871, 16'd7671, 16'd61507, 16'd15796, 16'd32228, 16'd36198, 16'd47607, 16'd24668, 16'd30150, 16'd19015, 16'd47021, 16'd56224, 16'd44815, 16'd6480, 16'd20578, 16'd2181, 16'd18496, 16'd20800, 16'd21889, 16'd31863, 16'd55199});
	test_expansion(128'h6c29836ecf857d40b4eb7e572dff685f, {16'd24899, 16'd47350, 16'd36721, 16'd9218, 16'd51636, 16'd44703, 16'd57376, 16'd19966, 16'd30627, 16'd49468, 16'd48782, 16'd26798, 16'd19770, 16'd12654, 16'd15745, 16'd3583, 16'd5264, 16'd150, 16'd16322, 16'd38690, 16'd60330, 16'd25859, 16'd25588, 16'd64782, 16'd23315, 16'd55677});
	test_expansion(128'h7452e01841c40623d401de3f290cd8e1, {16'd22951, 16'd43350, 16'd56658, 16'd9549, 16'd17285, 16'd48066, 16'd27588, 16'd59783, 16'd15681, 16'd65121, 16'd60660, 16'd22123, 16'd60427, 16'd33906, 16'd28268, 16'd25421, 16'd63220, 16'd24073, 16'd62931, 16'd44363, 16'd14711, 16'd52413, 16'd2855, 16'd63641, 16'd60548, 16'd50103});
	test_expansion(128'h79bd0fac428f614a55252f3abc6c0252, {16'd35352, 16'd41181, 16'd25266, 16'd19981, 16'd48443, 16'd45556, 16'd334, 16'd37757, 16'd26567, 16'd50649, 16'd51391, 16'd43345, 16'd10196, 16'd46553, 16'd22523, 16'd38885, 16'd32238, 16'd51797, 16'd45955, 16'd42745, 16'd36926, 16'd2947, 16'd4714, 16'd19256, 16'd52985, 16'd23488});
	test_expansion(128'hd5931601a87ef4395a909dc6a1c3064b, {16'd9772, 16'd1634, 16'd46159, 16'd46510, 16'd43158, 16'd47150, 16'd63396, 16'd60840, 16'd43578, 16'd41531, 16'd3491, 16'd59529, 16'd37842, 16'd54169, 16'd22120, 16'd15961, 16'd50618, 16'd57032, 16'd997, 16'd33207, 16'd22213, 16'd40861, 16'd36844, 16'd50314, 16'd32380, 16'd16567});
	test_expansion(128'h3687d907d930cf7a42281a889952b93b, {16'd44417, 16'd38636, 16'd6029, 16'd59118, 16'd65400, 16'd485, 16'd14144, 16'd33609, 16'd24931, 16'd32231, 16'd16549, 16'd10595, 16'd19615, 16'd37559, 16'd2082, 16'd29001, 16'd39595, 16'd31794, 16'd18294, 16'd20030, 16'd1838, 16'd47352, 16'd38566, 16'd979, 16'd59551, 16'd58606});
	test_expansion(128'h0a387b6fe3aafe7e18558a96aa7d2e50, {16'd30139, 16'd48276, 16'd21454, 16'd7351, 16'd61406, 16'd51311, 16'd12422, 16'd10365, 16'd43292, 16'd18674, 16'd43589, 16'd9071, 16'd14023, 16'd64779, 16'd53235, 16'd44698, 16'd46001, 16'd15395, 16'd49875, 16'd24522, 16'd25981, 16'd47813, 16'd9987, 16'd21339, 16'd32745, 16'd37573});
	test_expansion(128'hf5d263a7374674ca57e061698330843d, {16'd41089, 16'd26385, 16'd45644, 16'd50428, 16'd51494, 16'd60573, 16'd49889, 16'd7298, 16'd4955, 16'd45414, 16'd11453, 16'd22933, 16'd7625, 16'd31561, 16'd7833, 16'd16541, 16'd39007, 16'd43320, 16'd16943, 16'd23284, 16'd20836, 16'd62868, 16'd37432, 16'd36495, 16'd24276, 16'd32689});
	test_expansion(128'h63c036e6b31333955f3f67f17eeafcb3, {16'd25814, 16'd24828, 16'd16918, 16'd31506, 16'd3205, 16'd55094, 16'd15671, 16'd15804, 16'd20525, 16'd38931, 16'd27006, 16'd52468, 16'd50703, 16'd21968, 16'd38224, 16'd61584, 16'd47503, 16'd6575, 16'd24818, 16'd50143, 16'd16645, 16'd43397, 16'd35550, 16'd40091, 16'd2009, 16'd11806});
	test_expansion(128'h19dc5d9f826101ff2f7e10350d3345c6, {16'd26590, 16'd27451, 16'd3315, 16'd2737, 16'd17863, 16'd18741, 16'd19380, 16'd23154, 16'd60774, 16'd50989, 16'd15469, 16'd40601, 16'd22834, 16'd42968, 16'd30690, 16'd62729, 16'd5254, 16'd50173, 16'd41908, 16'd41323, 16'd26507, 16'd58152, 16'd35296, 16'd12919, 16'd11332, 16'd44642});
	test_expansion(128'h7b1d7f7c06a418134dd473f50534e7d0, {16'd6340, 16'd21691, 16'd22935, 16'd22350, 16'd9253, 16'd16868, 16'd28172, 16'd14151, 16'd13918, 16'd27603, 16'd52780, 16'd28966, 16'd62429, 16'd54130, 16'd24983, 16'd6316, 16'd59033, 16'd28963, 16'd31598, 16'd64660, 16'd64370, 16'd2267, 16'd48864, 16'd45273, 16'd26474, 16'd60263});
	test_expansion(128'h53c6aac2093f44b1a031fec9d52ed369, {16'd43802, 16'd21382, 16'd63539, 16'd7103, 16'd33118, 16'd23371, 16'd489, 16'd39739, 16'd38835, 16'd12577, 16'd61428, 16'd9237, 16'd46023, 16'd12897, 16'd30782, 16'd43514, 16'd3664, 16'd19908, 16'd39747, 16'd8666, 16'd54362, 16'd7929, 16'd53435, 16'd44114, 16'd26561, 16'd36116});
	test_expansion(128'h64fa07a09559809844d05a8dc5eee5a4, {16'd11137, 16'd1291, 16'd21314, 16'd12256, 16'd27432, 16'd9875, 16'd57147, 16'd51687, 16'd9558, 16'd29563, 16'd50789, 16'd63889, 16'd51543, 16'd27870, 16'd40239, 16'd51188, 16'd65379, 16'd10839, 16'd46393, 16'd57140, 16'd58340, 16'd52068, 16'd42186, 16'd57225, 16'd2014, 16'd6381});
	test_expansion(128'h03145b61201e37a67c87a596f1188e5d, {16'd27201, 16'd20197, 16'd64240, 16'd8425, 16'd263, 16'd3995, 16'd42114, 16'd9624, 16'd18713, 16'd54071, 16'd39745, 16'd31871, 16'd6783, 16'd36654, 16'd50420, 16'd54611, 16'd37517, 16'd62646, 16'd23538, 16'd20722, 16'd35257, 16'd46113, 16'd18684, 16'd25451, 16'd44298, 16'd65211});
	test_expansion(128'habc5aee82f35a8375a85833d3be9bc55, {16'd29291, 16'd52099, 16'd30228, 16'd4851, 16'd50797, 16'd53159, 16'd42999, 16'd32265, 16'd42509, 16'd17017, 16'd7299, 16'd19837, 16'd22640, 16'd44584, 16'd19029, 16'd31433, 16'd33778, 16'd16192, 16'd32219, 16'd63178, 16'd24341, 16'd26408, 16'd55162, 16'd62201, 16'd40662, 16'd58604});
	test_expansion(128'h09628f3540076e01b11d5f7940498c1a, {16'd14123, 16'd31921, 16'd41437, 16'd19993, 16'd64533, 16'd13550, 16'd21769, 16'd1041, 16'd9189, 16'd25514, 16'd9557, 16'd49984, 16'd33143, 16'd56195, 16'd60916, 16'd19067, 16'd3057, 16'd16021, 16'd43157, 16'd50194, 16'd22289, 16'd54309, 16'd14507, 16'd46459, 16'd14593, 16'd56547});
	test_expansion(128'hc2fc47511c12c24c593058cb648d766d, {16'd50060, 16'd21401, 16'd23553, 16'd61140, 16'd23555, 16'd40547, 16'd61387, 16'd30162, 16'd9947, 16'd6800, 16'd60855, 16'd37914, 16'd21109, 16'd15702, 16'd6320, 16'd41101, 16'd49584, 16'd18095, 16'd51346, 16'd50860, 16'd56083, 16'd21845, 16'd55123, 16'd46695, 16'd5704, 16'd8160});
	test_expansion(128'h8138aca0a2fc09526f01eb684e9cb7b1, {16'd23584, 16'd27978, 16'd43907, 16'd28538, 16'd55064, 16'd57308, 16'd26677, 16'd2365, 16'd40815, 16'd19584, 16'd43928, 16'd51490, 16'd54058, 16'd60875, 16'd50906, 16'd28622, 16'd1499, 16'd37531, 16'd16412, 16'd34040, 16'd5148, 16'd35349, 16'd39425, 16'd53064, 16'd27419, 16'd25353});
	test_expansion(128'he9dea8ae87d18f032485ba5a4b07c367, {16'd25815, 16'd32039, 16'd61270, 16'd64717, 16'd15848, 16'd29466, 16'd15980, 16'd6756, 16'd52667, 16'd21093, 16'd64253, 16'd13865, 16'd34300, 16'd1828, 16'd48702, 16'd18747, 16'd20737, 16'd41689, 16'd63284, 16'd58773, 16'd6421, 16'd37555, 16'd43442, 16'd52929, 16'd62680, 16'd7387});
	test_expansion(128'h6ced26c60058f26622588cdd09b176b7, {16'd20306, 16'd17377, 16'd23223, 16'd5424, 16'd48301, 16'd56571, 16'd38260, 16'd125, 16'd33131, 16'd4013, 16'd28833, 16'd40395, 16'd56689, 16'd17065, 16'd37809, 16'd56133, 16'd56403, 16'd39572, 16'd30791, 16'd62248, 16'd46397, 16'd53543, 16'd58747, 16'd64052, 16'd32202, 16'd42298});
	test_expansion(128'h296f82a38f7642682dae1ed88689b8ee, {16'd12524, 16'd15206, 16'd62338, 16'd43693, 16'd16508, 16'd44815, 16'd23120, 16'd26726, 16'd45871, 16'd48595, 16'd60497, 16'd63803, 16'd22313, 16'd17167, 16'd22676, 16'd914, 16'd33686, 16'd13688, 16'd49712, 16'd39574, 16'd28029, 16'd16127, 16'd28698, 16'd17811, 16'd41270, 16'd42320});
	test_expansion(128'h842544362ac5aa68826b76cd93e55fa6, {16'd4495, 16'd63850, 16'd7089, 16'd47146, 16'd15464, 16'd27965, 16'd37905, 16'd54952, 16'd53466, 16'd11890, 16'd1755, 16'd47795, 16'd27509, 16'd62902, 16'd12994, 16'd21672, 16'd43842, 16'd27454, 16'd30839, 16'd16132, 16'd46343, 16'd63754, 16'd51164, 16'd21938, 16'd2840, 16'd17211});
	test_expansion(128'h482e10bb512545f4fe7d8f6aeef08989, {16'd34446, 16'd19741, 16'd25691, 16'd27181, 16'd53125, 16'd60466, 16'd28093, 16'd17608, 16'd9032, 16'd47594, 16'd62585, 16'd41561, 16'd26520, 16'd55615, 16'd1402, 16'd38897, 16'd50566, 16'd28685, 16'd29417, 16'd35644, 16'd30136, 16'd43133, 16'd43765, 16'd26097, 16'd63657, 16'd52668});
	test_expansion(128'h059728064005a6d6f7993d6fbf3ca3a1, {16'd33093, 16'd9167, 16'd32546, 16'd18835, 16'd117, 16'd12946, 16'd15807, 16'd53801, 16'd27276, 16'd4912, 16'd22603, 16'd47448, 16'd64165, 16'd13522, 16'd34998, 16'd64269, 16'd21450, 16'd26157, 16'd8469, 16'd5597, 16'd35202, 16'd1876, 16'd63809, 16'd59850, 16'd60590, 16'd23835});
	test_expansion(128'hd493b2620a0e8505eaed472ba08c718e, {16'd39360, 16'd48397, 16'd18751, 16'd5545, 16'd61094, 16'd4319, 16'd31284, 16'd48732, 16'd47644, 16'd47725, 16'd36974, 16'd47500, 16'd64749, 16'd14819, 16'd33894, 16'd28539, 16'd54958, 16'd27855, 16'd2461, 16'd43073, 16'd25928, 16'd65526, 16'd23418, 16'd28871, 16'd62500, 16'd18054});
	test_expansion(128'hf2dee907f61f45a42421bb7802391c5d, {16'd35452, 16'd21703, 16'd19001, 16'd24169, 16'd38410, 16'd3923, 16'd41324, 16'd44171, 16'd45381, 16'd23693, 16'd30314, 16'd38724, 16'd48686, 16'd10632, 16'd40698, 16'd34695, 16'd16179, 16'd4695, 16'd57293, 16'd55337, 16'd46656, 16'd36185, 16'd36802, 16'd58780, 16'd56539, 16'd19399});
	test_expansion(128'he1608655546ec1ad13b7ad0b05414431, {16'd64150, 16'd5604, 16'd39735, 16'd59951, 16'd57724, 16'd22201, 16'd10252, 16'd26319, 16'd36573, 16'd7589, 16'd53412, 16'd60697, 16'd58268, 16'd45484, 16'd51053, 16'd51435, 16'd64067, 16'd21812, 16'd48440, 16'd54250, 16'd11559, 16'd51310, 16'd26129, 16'd32301, 16'd34050, 16'd16903});
	test_expansion(128'h5f267c95457085acaef1f18653df4829, {16'd5866, 16'd4093, 16'd59523, 16'd19137, 16'd26329, 16'd15351, 16'd48418, 16'd16481, 16'd49452, 16'd45669, 16'd36504, 16'd35893, 16'd14722, 16'd12927, 16'd50657, 16'd21272, 16'd24596, 16'd40639, 16'd24641, 16'd8964, 16'd56619, 16'd49366, 16'd5354, 16'd3949, 16'd13934, 16'd21270});
	test_expansion(128'h633ec5e796e10aae8ed69a50f2b2b783, {16'd65097, 16'd35469, 16'd53711, 16'd47795, 16'd4687, 16'd51821, 16'd31927, 16'd24780, 16'd27986, 16'd58962, 16'd29108, 16'd26176, 16'd11495, 16'd43586, 16'd55275, 16'd24215, 16'd58172, 16'd26585, 16'd1650, 16'd13691, 16'd26580, 16'd21366, 16'd54733, 16'd1264, 16'd9083, 16'd17865});
	test_expansion(128'h2e491f11603acbad667a8311e299dc41, {16'd9137, 16'd60786, 16'd39529, 16'd30300, 16'd26810, 16'd59189, 16'd12821, 16'd13992, 16'd28290, 16'd34578, 16'd33238, 16'd38348, 16'd31628, 16'd47748, 16'd42364, 16'd11246, 16'd5558, 16'd19050, 16'd36963, 16'd64527, 16'd40976, 16'd33044, 16'd49500, 16'd24670, 16'd55147, 16'd37458});
	test_expansion(128'h2645de920f7e1a0f3a72715c9d136f34, {16'd6620, 16'd33391, 16'd33813, 16'd38759, 16'd54288, 16'd16741, 16'd61711, 16'd42656, 16'd25241, 16'd46901, 16'd1505, 16'd18148, 16'd31071, 16'd48236, 16'd44198, 16'd58140, 16'd32977, 16'd61821, 16'd54088, 16'd15764, 16'd22551, 16'd20858, 16'd3575, 16'd41832, 16'd62252, 16'd29807});
	test_expansion(128'hd8b99d8be39d3ff4dfe8ed9ba95ccb29, {16'd55299, 16'd46143, 16'd47837, 16'd131, 16'd58101, 16'd40142, 16'd46227, 16'd43727, 16'd32402, 16'd3446, 16'd5832, 16'd17266, 16'd57949, 16'd61776, 16'd17104, 16'd17937, 16'd33445, 16'd55502, 16'd58212, 16'd10474, 16'd13822, 16'd1951, 16'd22362, 16'd58110, 16'd63387, 16'd9662});
	test_expansion(128'h53f076808479ae772524f0ed31d3dce4, {16'd38412, 16'd58160, 16'd43369, 16'd10477, 16'd3085, 16'd22247, 16'd19322, 16'd11316, 16'd54736, 16'd31170, 16'd50921, 16'd50282, 16'd54751, 16'd19645, 16'd38832, 16'd18643, 16'd29367, 16'd53161, 16'd14251, 16'd59495, 16'd64916, 16'd53359, 16'd15449, 16'd45399, 16'd7576, 16'd61189});
	test_expansion(128'h453dd3a6e0e791a22e609e7c9d847f83, {16'd18414, 16'd6209, 16'd58804, 16'd22224, 16'd43361, 16'd54988, 16'd31223, 16'd60201, 16'd26970, 16'd48451, 16'd11467, 16'd17813, 16'd18274, 16'd8106, 16'd31114, 16'd61945, 16'd28442, 16'd54085, 16'd21822, 16'd42992, 16'd25579, 16'd25822, 16'd40537, 16'd7018, 16'd60953, 16'd29764});
	test_expansion(128'h4993eb2eed77470f7920d9d0225007d6, {16'd19179, 16'd27954, 16'd46725, 16'd11839, 16'd42375, 16'd57472, 16'd3582, 16'd56554, 16'd20614, 16'd52532, 16'd47650, 16'd22578, 16'd32538, 16'd41929, 16'd59326, 16'd19465, 16'd9842, 16'd61034, 16'd9377, 16'd42196, 16'd2068, 16'd6973, 16'd64119, 16'd56543, 16'd38709, 16'd65206});
	test_expansion(128'hc6d962078ffd3f42f565f06a3bfd325e, {16'd30128, 16'd32522, 16'd38270, 16'd19399, 16'd399, 16'd9356, 16'd50343, 16'd31654, 16'd56826, 16'd61087, 16'd3387, 16'd1691, 16'd38821, 16'd43044, 16'd20840, 16'd63627, 16'd43229, 16'd17519, 16'd36755, 16'd57216, 16'd7338, 16'd28924, 16'd24336, 16'd49484, 16'd40962, 16'd23077});
	test_expansion(128'h082ca00bc6314e887b654d113616d3b0, {16'd42409, 16'd11179, 16'd10602, 16'd12984, 16'd7097, 16'd39712, 16'd25839, 16'd4414, 16'd20741, 16'd13738, 16'd64371, 16'd12377, 16'd46525, 16'd58169, 16'd64528, 16'd52692, 16'd49828, 16'd17782, 16'd40506, 16'd63698, 16'd35133, 16'd16588, 16'd34505, 16'd28496, 16'd61844, 16'd48650});
	test_expansion(128'h986988b0c7c32c04ae7dd38b0b919daf, {16'd49795, 16'd54931, 16'd6332, 16'd64534, 16'd5253, 16'd31886, 16'd8477, 16'd13849, 16'd26191, 16'd59808, 16'd59014, 16'd43856, 16'd12304, 16'd2924, 16'd53736, 16'd5919, 16'd3567, 16'd8589, 16'd14676, 16'd12652, 16'd42245, 16'd63603, 16'd37553, 16'd9083, 16'd38416, 16'd34793});
	test_expansion(128'h33f0d664e719dacda63bf40fdb04335a, {16'd31166, 16'd42843, 16'd43019, 16'd24274, 16'd39593, 16'd5472, 16'd58933, 16'd26425, 16'd4500, 16'd25988, 16'd43923, 16'd18928, 16'd22821, 16'd45472, 16'd6085, 16'd28646, 16'd52703, 16'd48404, 16'd20223, 16'd6671, 16'd7585, 16'd53204, 16'd6709, 16'd32034, 16'd50084, 16'd38715});
	test_expansion(128'h9e2daa042e8f9030303d4d5d8105562c, {16'd8471, 16'd59211, 16'd57305, 16'd40314, 16'd39197, 16'd35704, 16'd63928, 16'd40271, 16'd14897, 16'd824, 16'd39522, 16'd34248, 16'd22908, 16'd18548, 16'd26422, 16'd20145, 16'd2308, 16'd3058, 16'd34982, 16'd3866, 16'd5216, 16'd36141, 16'd20756, 16'd26884, 16'd52943, 16'd3668});
	test_expansion(128'h7f2dbb0ec91e42ca9ed46956ee63127a, {16'd23389, 16'd46707, 16'd23506, 16'd2181, 16'd45655, 16'd49401, 16'd15772, 16'd15007, 16'd3599, 16'd65172, 16'd25514, 16'd6928, 16'd60830, 16'd8185, 16'd52778, 16'd2445, 16'd7262, 16'd4010, 16'd13501, 16'd48433, 16'd8482, 16'd51330, 16'd51613, 16'd5706, 16'd41145, 16'd55164});
	test_expansion(128'h795910dee7b9c0aa547174ccc4681246, {16'd17723, 16'd39454, 16'd3596, 16'd47412, 16'd2844, 16'd54036, 16'd20832, 16'd44480, 16'd32108, 16'd46035, 16'd58471, 16'd19968, 16'd34952, 16'd14039, 16'd23691, 16'd42980, 16'd48658, 16'd39099, 16'd60068, 16'd47536, 16'd13105, 16'd26986, 16'd53560, 16'd56857, 16'd32541, 16'd25674});
	test_expansion(128'hcb308e080510ac127cc2d886892b15ea, {16'd31272, 16'd7218, 16'd43441, 16'd35003, 16'd15501, 16'd47071, 16'd22733, 16'd62387, 16'd28270, 16'd47912, 16'd11532, 16'd18367, 16'd62985, 16'd46673, 16'd29473, 16'd18698, 16'd10852, 16'd30864, 16'd1223, 16'd17337, 16'd63479, 16'd22926, 16'd37200, 16'd48134, 16'd21071, 16'd46195});
	test_expansion(128'he96ac6a0b6b589ae48fb55dac1af0a70, {16'd14977, 16'd18702, 16'd52835, 16'd40161, 16'd4681, 16'd65529, 16'd53276, 16'd51844, 16'd11192, 16'd61675, 16'd45055, 16'd42716, 16'd36414, 16'd9690, 16'd51749, 16'd55789, 16'd32315, 16'd1203, 16'd9831, 16'd58067, 16'd47719, 16'd20268, 16'd52219, 16'd3580, 16'd45762, 16'd17315});
	test_expansion(128'he738e275452fde89ad8a70a18dc8bffa, {16'd61253, 16'd8237, 16'd4496, 16'd55783, 16'd44441, 16'd28037, 16'd58446, 16'd32507, 16'd18069, 16'd16624, 16'd46305, 16'd20519, 16'd60405, 16'd49565, 16'd441, 16'd33124, 16'd59019, 16'd37038, 16'd22509, 16'd42555, 16'd6162, 16'd29418, 16'd33019, 16'd615, 16'd9847, 16'd32870});
	test_expansion(128'hbf7b514b70960fa9e6463276fadfd862, {16'd22779, 16'd30752, 16'd59528, 16'd36745, 16'd34763, 16'd22356, 16'd51833, 16'd39392, 16'd494, 16'd8593, 16'd1889, 16'd62268, 16'd43499, 16'd31258, 16'd36474, 16'd53695, 16'd15726, 16'd27923, 16'd5762, 16'd5604, 16'd30794, 16'd52374, 16'd16788, 16'd51343, 16'd45705, 16'd27216});
	test_expansion(128'hac56e084239603ac4cc5dbceeb949a00, {16'd13535, 16'd13931, 16'd19048, 16'd46232, 16'd18038, 16'd58816, 16'd19554, 16'd18383, 16'd62351, 16'd59752, 16'd2661, 16'd30472, 16'd3546, 16'd37718, 16'd15954, 16'd45076, 16'd36053, 16'd16888, 16'd15727, 16'd5564, 16'd50276, 16'd88, 16'd58248, 16'd23083, 16'd16942, 16'd26196});
	test_expansion(128'h03739f3c049d3e6c57e8ced715a50bc3, {16'd40027, 16'd28125, 16'd39839, 16'd18705, 16'd59742, 16'd42273, 16'd55421, 16'd30824, 16'd36433, 16'd63367, 16'd18480, 16'd4162, 16'd9260, 16'd5080, 16'd24064, 16'd43670, 16'd27643, 16'd17281, 16'd18550, 16'd6313, 16'd485, 16'd28960, 16'd51742, 16'd21506, 16'd24690, 16'd14110});
	test_expansion(128'h8c1cd2c974e1f89cddfa5eea0ac42bfc, {16'd42324, 16'd1141, 16'd27118, 16'd36644, 16'd31074, 16'd20115, 16'd13045, 16'd1539, 16'd55665, 16'd42241, 16'd12151, 16'd29546, 16'd22456, 16'd1736, 16'd57497, 16'd21498, 16'd26250, 16'd36599, 16'd42365, 16'd39156, 16'd8661, 16'd63210, 16'd40077, 16'd17438, 16'd28973, 16'd3575});
	test_expansion(128'hc11c1b8a11b749430257d3e0dc3e6b2b, {16'd29519, 16'd15578, 16'd39837, 16'd56692, 16'd43271, 16'd15243, 16'd39522, 16'd1427, 16'd15811, 16'd53866, 16'd12310, 16'd62113, 16'd9572, 16'd45547, 16'd30885, 16'd53669, 16'd51255, 16'd63813, 16'd19570, 16'd18242, 16'd60468, 16'd25307, 16'd51747, 16'd24833, 16'd65432, 16'd41069});
	test_expansion(128'habc9d91951f08e2d374dd0d328fd3057, {16'd34638, 16'd18170, 16'd35024, 16'd53605, 16'd56040, 16'd53733, 16'd54509, 16'd42016, 16'd46991, 16'd57713, 16'd47822, 16'd10955, 16'd31601, 16'd25624, 16'd54310, 16'd7452, 16'd64287, 16'd42487, 16'd39996, 16'd55762, 16'd13108, 16'd4741, 16'd43096, 16'd30692, 16'd30713, 16'd22979});
	test_expansion(128'hca8fd39363f2220a0a9f64da5b62939d, {16'd55282, 16'd24227, 16'd26521, 16'd56173, 16'd43001, 16'd51070, 16'd6604, 16'd19474, 16'd37091, 16'd20675, 16'd16865, 16'd49119, 16'd6321, 16'd59264, 16'd12144, 16'd53524, 16'd16363, 16'd28998, 16'd19131, 16'd40789, 16'd25034, 16'd64279, 16'd20359, 16'd4146, 16'd17577, 16'd30693});
	test_expansion(128'ha1e60bd83bcbe02ba3247056e51f47b2, {16'd39491, 16'd7808, 16'd50706, 16'd51563, 16'd31281, 16'd29358, 16'd45194, 16'd27995, 16'd11156, 16'd2928, 16'd63571, 16'd46452, 16'd37463, 16'd30197, 16'd30777, 16'd9914, 16'd60211, 16'd44954, 16'd31683, 16'd59701, 16'd6212, 16'd26611, 16'd9121, 16'd62126, 16'd3236, 16'd5877});
	test_expansion(128'h9909571ff7306453bc2fbee920aa7804, {16'd52318, 16'd44918, 16'd15170, 16'd9089, 16'd8005, 16'd58550, 16'd7883, 16'd59019, 16'd6324, 16'd41171, 16'd4986, 16'd37987, 16'd52353, 16'd36638, 16'd8598, 16'd44440, 16'd55262, 16'd25469, 16'd42182, 16'd11026, 16'd6715, 16'd64879, 16'd37482, 16'd34975, 16'd3010, 16'd50562});
	test_expansion(128'h73cd94d261b3003c381b1ad2964cf488, {16'd52528, 16'd33635, 16'd58442, 16'd34533, 16'd14154, 16'd12223, 16'd61648, 16'd5454, 16'd45958, 16'd51094, 16'd52003, 16'd38256, 16'd29792, 16'd19612, 16'd57465, 16'd47782, 16'd64599, 16'd53151, 16'd56146, 16'd51912, 16'd9725, 16'd36902, 16'd51451, 16'd8394, 16'd12597, 16'd46748});
	test_expansion(128'hac30276f8ce9978728aef0805caa9ef0, {16'd25535, 16'd58923, 16'd4896, 16'd62698, 16'd21438, 16'd13256, 16'd58982, 16'd22625, 16'd57560, 16'd16734, 16'd47677, 16'd49705, 16'd40369, 16'd23265, 16'd48750, 16'd25874, 16'd28420, 16'd62439, 16'd3, 16'd40147, 16'd54307, 16'd43851, 16'd17203, 16'd23109, 16'd23529, 16'd34077});
	test_expansion(128'hfe19b61e4812c29fb119e4e4fbf2c242, {16'd59325, 16'd5472, 16'd62250, 16'd46651, 16'd12912, 16'd25356, 16'd4467, 16'd63123, 16'd53788, 16'd24607, 16'd56765, 16'd29436, 16'd34995, 16'd46240, 16'd65115, 16'd1784, 16'd33691, 16'd64196, 16'd5800, 16'd20410, 16'd43171, 16'd23281, 16'd33721, 16'd24396, 16'd46754, 16'd16337});
	test_expansion(128'he6f08734ee00915fd242c5cd23008b60, {16'd12981, 16'd33231, 16'd50463, 16'd24559, 16'd1608, 16'd15130, 16'd21796, 16'd8843, 16'd24975, 16'd42671, 16'd11395, 16'd45956, 16'd59964, 16'd45696, 16'd22764, 16'd15103, 16'd15913, 16'd64047, 16'd9195, 16'd58408, 16'd16247, 16'd54345, 16'd15327, 16'd39714, 16'd31663, 16'd14677});
	test_expansion(128'h6c5b7f51746162597e394dacbadc6d39, {16'd53778, 16'd16499, 16'd59894, 16'd3817, 16'd36054, 16'd37898, 16'd2544, 16'd37407, 16'd6639, 16'd13384, 16'd19150, 16'd10629, 16'd27593, 16'd21551, 16'd25722, 16'd52669, 16'd8036, 16'd31719, 16'd20589, 16'd40638, 16'd2882, 16'd5042, 16'd46930, 16'd13093, 16'd59942, 16'd23721});
	test_expansion(128'hc9a6838863fe59ebb4cb43062f2dbbc4, {16'd55938, 16'd51511, 16'd4791, 16'd50015, 16'd51982, 16'd50263, 16'd15889, 16'd33821, 16'd15851, 16'd10148, 16'd25513, 16'd28987, 16'd9937, 16'd37528, 16'd21019, 16'd64046, 16'd15124, 16'd53526, 16'd60316, 16'd12295, 16'd11622, 16'd43975, 16'd46331, 16'd18052, 16'd7807, 16'd25428});
	test_expansion(128'h7ae36f58ae5c6c7896563fd04fc8df2b, {16'd55812, 16'd29211, 16'd4304, 16'd33504, 16'd34775, 16'd20989, 16'd14969, 16'd2775, 16'd43647, 16'd11614, 16'd43679, 16'd50202, 16'd10043, 16'd22118, 16'd54000, 16'd23591, 16'd63022, 16'd24164, 16'd36286, 16'd62601, 16'd18988, 16'd41291, 16'd24182, 16'd23641, 16'd6188, 16'd35682});
	test_expansion(128'had7a1bd43622e9a245851dea9cee17c3, {16'd43306, 16'd3997, 16'd63324, 16'd44390, 16'd12382, 16'd32781, 16'd48609, 16'd42423, 16'd14890, 16'd33571, 16'd60194, 16'd49229, 16'd39517, 16'd23511, 16'd15046, 16'd25494, 16'd29206, 16'd21932, 16'd23480, 16'd32687, 16'd61067, 16'd46070, 16'd41424, 16'd5259, 16'd3823, 16'd60205});
	test_expansion(128'h93f0b9f1468dc5be07aa06447a2c7fa9, {16'd19455, 16'd20708, 16'd34201, 16'd8647, 16'd33781, 16'd27204, 16'd41070, 16'd13128, 16'd56049, 16'd45933, 16'd48433, 16'd30596, 16'd17375, 16'd49335, 16'd4415, 16'd28213, 16'd6146, 16'd55228, 16'd57727, 16'd47325, 16'd50929, 16'd7128, 16'd43082, 16'd18189, 16'd26542, 16'd59971});
	test_expansion(128'h5ed8ca9b89bb1309e0c91d938c98978b, {16'd63404, 16'd6674, 16'd30747, 16'd34617, 16'd41803, 16'd38846, 16'd6275, 16'd5478, 16'd35474, 16'd972, 16'd26585, 16'd28064, 16'd61373, 16'd2014, 16'd11950, 16'd1671, 16'd36228, 16'd39321, 16'd5965, 16'd26566, 16'd43770, 16'd63642, 16'd18442, 16'd10817, 16'd1814, 16'd20783});
	test_expansion(128'hc518fd85f503633650842f3d1d7a1071, {16'd32260, 16'd50397, 16'd42673, 16'd4991, 16'd6397, 16'd56661, 16'd32739, 16'd57322, 16'd63376, 16'd65349, 16'd37026, 16'd40191, 16'd28872, 16'd32922, 16'd51017, 16'd32149, 16'd3509, 16'd62975, 16'd62769, 16'd30621, 16'd24777, 16'd19315, 16'd19598, 16'd44783, 16'd13913, 16'd64397});
	test_expansion(128'h98b35c63819d9cad4c5ed7778f02dec6, {16'd27222, 16'd25588, 16'd6034, 16'd47736, 16'd52310, 16'd60547, 16'd46545, 16'd15275, 16'd3808, 16'd26480, 16'd57354, 16'd32731, 16'd44920, 16'd1951, 16'd54278, 16'd45820, 16'd6905, 16'd57833, 16'd15074, 16'd32951, 16'd65239, 16'd23669, 16'd6617, 16'd12059, 16'd21567, 16'd12561});
	test_expansion(128'hf1b82e147c2ab438f9659abd89f34841, {16'd47357, 16'd10848, 16'd36005, 16'd32087, 16'd44177, 16'd20784, 16'd6537, 16'd53161, 16'd15247, 16'd64185, 16'd3112, 16'd8205, 16'd28485, 16'd27258, 16'd59937, 16'd17840, 16'd15377, 16'd64180, 16'd61757, 16'd60823, 16'd38608, 16'd33400, 16'd57729, 16'd28031, 16'd25391, 16'd14619});
	test_expansion(128'h1b2ef93d916a53446c3f49b00079972d, {16'd38829, 16'd5799, 16'd18628, 16'd45589, 16'd44240, 16'd11109, 16'd11587, 16'd53224, 16'd24576, 16'd64231, 16'd2685, 16'd7743, 16'd41282, 16'd39626, 16'd49019, 16'd8059, 16'd45446, 16'd32316, 16'd30308, 16'd35839, 16'd14356, 16'd4836, 16'd33737, 16'd29847, 16'd51429, 16'd52155});
	test_expansion(128'h4f106801fb0bb3e9153844127293ac04, {16'd48635, 16'd5146, 16'd9939, 16'd25355, 16'd53192, 16'd65037, 16'd59431, 16'd56822, 16'd47933, 16'd40414, 16'd37461, 16'd41709, 16'd3411, 16'd37261, 16'd41896, 16'd6825, 16'd18699, 16'd43238, 16'd65275, 16'd17184, 16'd359, 16'd690, 16'd55333, 16'd63687, 16'd17794, 16'd29495});
	test_expansion(128'he28db7c7f4a823ecafdd5053ff9c215f, {16'd51499, 16'd35402, 16'd61738, 16'd51185, 16'd55340, 16'd61146, 16'd52670, 16'd55958, 16'd43485, 16'd49578, 16'd51473, 16'd47879, 16'd23559, 16'd33342, 16'd6706, 16'd64989, 16'd32322, 16'd63481, 16'd44989, 16'd2555, 16'd1909, 16'd50967, 16'd38089, 16'd18820, 16'd24789, 16'd7589});
	test_expansion(128'h4bb64d4bb9a09d7ed3e64662b074279d, {16'd37837, 16'd47717, 16'd29691, 16'd57834, 16'd59008, 16'd20829, 16'd6825, 16'd32037, 16'd55028, 16'd37631, 16'd10132, 16'd1508, 16'd8047, 16'd43671, 16'd33135, 16'd39458, 16'd58664, 16'd58014, 16'd64057, 16'd49784, 16'd10653, 16'd18456, 16'd6556, 16'd38762, 16'd62527, 16'd38282});
	test_expansion(128'h4ee84954eefeba16fb046346a4ca116a, {16'd21636, 16'd26091, 16'd54188, 16'd25024, 16'd37185, 16'd55124, 16'd23564, 16'd59217, 16'd54578, 16'd63859, 16'd32294, 16'd33136, 16'd62129, 16'd31717, 16'd15189, 16'd29346, 16'd5548, 16'd59683, 16'd25724, 16'd38811, 16'd50550, 16'd58684, 16'd40460, 16'd40581, 16'd21158, 16'd404});
	test_expansion(128'h58a0c841df4efebc6604458eb738911c, {16'd9580, 16'd18077, 16'd30943, 16'd64419, 16'd55215, 16'd53087, 16'd23183, 16'd46317, 16'd355, 16'd33864, 16'd13728, 16'd4753, 16'd25370, 16'd11413, 16'd43146, 16'd17184, 16'd18688, 16'd47183, 16'd29812, 16'd23843, 16'd8175, 16'd17600, 16'd53596, 16'd37633, 16'd10475, 16'd9854});
	test_expansion(128'he541f4b19e878d50bd54bdae87415391, {16'd9091, 16'd43853, 16'd27175, 16'd48352, 16'd47158, 16'd50421, 16'd13410, 16'd18798, 16'd19654, 16'd51933, 16'd11639, 16'd19438, 16'd19708, 16'd43359, 16'd29923, 16'd11382, 16'd17294, 16'd14214, 16'd6101, 16'd17118, 16'd50419, 16'd50231, 16'd1780, 16'd37448, 16'd1530, 16'd63385});
	test_expansion(128'h43e11ff4d661e254dadfd0072a706bd5, {16'd14555, 16'd18485, 16'd3383, 16'd46769, 16'd22483, 16'd21123, 16'd54994, 16'd39402, 16'd35889, 16'd2255, 16'd42433, 16'd5564, 16'd47096, 16'd33527, 16'd32357, 16'd54170, 16'd60601, 16'd30775, 16'd13837, 16'd2459, 16'd33710, 16'd10259, 16'd41785, 16'd4493, 16'd59837, 16'd41235});
	test_expansion(128'h86a7836244d23311e90e62d4794e8546, {16'd19668, 16'd60348, 16'd8797, 16'd53685, 16'd7547, 16'd24985, 16'd51362, 16'd19810, 16'd10002, 16'd61451, 16'd17556, 16'd23547, 16'd36124, 16'd33296, 16'd5005, 16'd32101, 16'd43026, 16'd18444, 16'd17928, 16'd40556, 16'd34771, 16'd25630, 16'd33802, 16'd8737, 16'd22196, 16'd12973});
	test_expansion(128'h60d1acb608785f975cfff09c03ea547f, {16'd42571, 16'd6678, 16'd15882, 16'd1374, 16'd3466, 16'd53980, 16'd37525, 16'd22198, 16'd7078, 16'd13213, 16'd27945, 16'd6084, 16'd10699, 16'd16467, 16'd49788, 16'd38525, 16'd17159, 16'd63745, 16'd56198, 16'd12819, 16'd60326, 16'd18759, 16'd48411, 16'd25263, 16'd51350, 16'd56131});
	test_expansion(128'h0a431ba27e8b215b4ca3a426b9ad8319, {16'd65156, 16'd51272, 16'd36245, 16'd14917, 16'd22516, 16'd51503, 16'd14740, 16'd41577, 16'd10912, 16'd40508, 16'd11108, 16'd2490, 16'd1653, 16'd53071, 16'd49720, 16'd7592, 16'd30674, 16'd23340, 16'd37824, 16'd8134, 16'd59058, 16'd37345, 16'd9696, 16'd15833, 16'd14318, 16'd11355});
	test_expansion(128'he993ff67bbbf380c6c083152feb7b335, {16'd60169, 16'd60559, 16'd43263, 16'd25478, 16'd51953, 16'd64264, 16'd31273, 16'd60149, 16'd61347, 16'd2311, 16'd24946, 16'd20965, 16'd65097, 16'd25122, 16'd42491, 16'd6986, 16'd26295, 16'd18845, 16'd5156, 16'd3444, 16'd49494, 16'd16944, 16'd17784, 16'd44540, 16'd38908, 16'd62528});
	test_expansion(128'h5f473a754efc43f8e861577a16829f33, {16'd12405, 16'd48642, 16'd47024, 16'd45097, 16'd24910, 16'd38514, 16'd2207, 16'd56544, 16'd17073, 16'd51778, 16'd15426, 16'd30553, 16'd35590, 16'd43141, 16'd56465, 16'd28859, 16'd21612, 16'd19076, 16'd41996, 16'd47281, 16'd32604, 16'd2348, 16'd54049, 16'd48028, 16'd34606, 16'd32427});
	test_expansion(128'h85128ae8e0cef6285c6485639bd4a75a, {16'd16905, 16'd46631, 16'd60445, 16'd27789, 16'd19010, 16'd63044, 16'd13610, 16'd1246, 16'd396, 16'd596, 16'd9037, 16'd55286, 16'd6384, 16'd41059, 16'd49969, 16'd38571, 16'd28829, 16'd6880, 16'd29820, 16'd60411, 16'd33842, 16'd33064, 16'd49849, 16'd30288, 16'd48618, 16'd52646});
	test_expansion(128'hd7c9c69dd0298150b8e8f5723f828d3a, {16'd10620, 16'd26016, 16'd20873, 16'd5191, 16'd57668, 16'd50242, 16'd47361, 16'd18870, 16'd43075, 16'd11455, 16'd31610, 16'd10467, 16'd51490, 16'd57757, 16'd43645, 16'd45452, 16'd37488, 16'd26823, 16'd62580, 16'd49673, 16'd12171, 16'd45547, 16'd29158, 16'd62665, 16'd46673, 16'd24928});
	test_expansion(128'h60cc68cd108c43ac6bc9b6d0f4097a07, {16'd12820, 16'd58577, 16'd10509, 16'd26083, 16'd7288, 16'd29694, 16'd54310, 16'd62024, 16'd63448, 16'd21626, 16'd929, 16'd51200, 16'd4801, 16'd18823, 16'd47541, 16'd38268, 16'd31509, 16'd33559, 16'd53068, 16'd30423, 16'd9667, 16'd36259, 16'd31770, 16'd5061, 16'd53382, 16'd6261});
	test_expansion(128'h5b191086d5b4f86cd297b92eeb57da23, {16'd35244, 16'd40399, 16'd26733, 16'd62145, 16'd40576, 16'd54714, 16'd34468, 16'd33092, 16'd53739, 16'd8153, 16'd4061, 16'd15187, 16'd37086, 16'd34416, 16'd50701, 16'd23497, 16'd41245, 16'd39948, 16'd62433, 16'd34383, 16'd52683, 16'd22648, 16'd54238, 16'd37517, 16'd28968, 16'd38449});
	test_expansion(128'h2050b5819ab6a38a8adb4d20796181dc, {16'd61307, 16'd9632, 16'd32943, 16'd33383, 16'd50421, 16'd30658, 16'd7180, 16'd51821, 16'd19349, 16'd22225, 16'd52577, 16'd64320, 16'd1151, 16'd35436, 16'd25562, 16'd1458, 16'd14052, 16'd18671, 16'd6905, 16'd10043, 16'd38868, 16'd63559, 16'd4032, 16'd15584, 16'd59966, 16'd10046});
	test_expansion(128'hb933df5b662f940ab3acb91388883f06, {16'd59412, 16'd55165, 16'd8174, 16'd54627, 16'd17617, 16'd31940, 16'd32227, 16'd25629, 16'd20692, 16'd3939, 16'd3841, 16'd6693, 16'd45859, 16'd56866, 16'd5305, 16'd40937, 16'd47466, 16'd7595, 16'd37477, 16'd2998, 16'd25076, 16'd34256, 16'd9982, 16'd55324, 16'd30762, 16'd32426});
	test_expansion(128'h5c336d255871b04bf4820706560e8349, {16'd48698, 16'd60387, 16'd4028, 16'd6042, 16'd33693, 16'd61476, 16'd34205, 16'd18173, 16'd57131, 16'd15864, 16'd32183, 16'd4757, 16'd3608, 16'd27667, 16'd40526, 16'd23235, 16'd52908, 16'd2052, 16'd4409, 16'd50875, 16'd12011, 16'd17485, 16'd8435, 16'd19834, 16'd30515, 16'd55676});
	test_expansion(128'hae4b0b352d470a99fc69b4f332c9e026, {16'd20720, 16'd27991, 16'd30959, 16'd37047, 16'd22804, 16'd27389, 16'd14204, 16'd45269, 16'd21056, 16'd65519, 16'd11753, 16'd54677, 16'd48168, 16'd7265, 16'd43390, 16'd60668, 16'd39324, 16'd54761, 16'd27461, 16'd9105, 16'd42316, 16'd1804, 16'd28689, 16'd32449, 16'd9838, 16'd62538});
	test_expansion(128'hb83d1963431d89a1df51cc1b805be423, {16'd26451, 16'd52553, 16'd36052, 16'd30975, 16'd61158, 16'd58933, 16'd26569, 16'd51649, 16'd64395, 16'd43112, 16'd23881, 16'd42576, 16'd43840, 16'd61626, 16'd64392, 16'd64820, 16'd45641, 16'd51910, 16'd11202, 16'd64314, 16'd2381, 16'd30627, 16'd37603, 16'd60825, 16'd20410, 16'd40765});
	test_expansion(128'hb2f831071a29445beb2af6ff648cfeef, {16'd61379, 16'd53842, 16'd49865, 16'd41395, 16'd24277, 16'd33961, 16'd28402, 16'd25869, 16'd12190, 16'd4193, 16'd7309, 16'd35604, 16'd50787, 16'd53438, 16'd20932, 16'd36139, 16'd37373, 16'd42507, 16'd24827, 16'd51757, 16'd51377, 16'd45260, 16'd18685, 16'd64147, 16'd13612, 16'd35310});
	test_expansion(128'h4970dbb76114446590b684c4b4b672f5, {16'd50452, 16'd266, 16'd8996, 16'd14972, 16'd50064, 16'd23092, 16'd4567, 16'd64970, 16'd8827, 16'd47881, 16'd63964, 16'd22989, 16'd30685, 16'd18826, 16'd62277, 16'd12861, 16'd62003, 16'd51, 16'd55159, 16'd38489, 16'd25340, 16'd32587, 16'd57873, 16'd27192, 16'd13960, 16'd63259});
	test_expansion(128'h0e94649277824543fd96f8946926f813, {16'd13684, 16'd62801, 16'd22069, 16'd56663, 16'd50651, 16'd61557, 16'd43571, 16'd14484, 16'd31217, 16'd52802, 16'd49916, 16'd15364, 16'd48530, 16'd21494, 16'd44490, 16'd56676, 16'd13715, 16'd61808, 16'd23465, 16'd51207, 16'd35023, 16'd17522, 16'd3833, 16'd37789, 16'd25227, 16'd47423});
	test_expansion(128'h2d549fa7333db860c6513d6685c6184f, {16'd27079, 16'd4981, 16'd64797, 16'd80, 16'd56883, 16'd20934, 16'd53216, 16'd1595, 16'd41595, 16'd37584, 16'd5835, 16'd52749, 16'd15194, 16'd43020, 16'd19996, 16'd1588, 16'd21716, 16'd1760, 16'd46835, 16'd5026, 16'd42748, 16'd25873, 16'd8290, 16'd26476, 16'd61856, 16'd53528});
	test_expansion(128'h0e40ce19d99d9712e23b06c636efa68b, {16'd2970, 16'd3635, 16'd33866, 16'd21500, 16'd10120, 16'd54391, 16'd23998, 16'd57794, 16'd44309, 16'd55554, 16'd53016, 16'd28597, 16'd44530, 16'd41666, 16'd18293, 16'd22964, 16'd57812, 16'd28840, 16'd38773, 16'd19640, 16'd41227, 16'd38175, 16'd46662, 16'd45494, 16'd22642, 16'd2283});
	test_expansion(128'hd9e527c8125f1d6e887596662b13ccbd, {16'd17656, 16'd62158, 16'd7778, 16'd13825, 16'd24932, 16'd61178, 16'd38418, 16'd7996, 16'd20045, 16'd44533, 16'd44050, 16'd3535, 16'd12394, 16'd10295, 16'd60651, 16'd4352, 16'd7558, 16'd5831, 16'd11963, 16'd60651, 16'd22191, 16'd36128, 16'd13670, 16'd53476, 16'd39366, 16'd35213});
	test_expansion(128'h4996722383d28477eb2b968698c10243, {16'd41521, 16'd42837, 16'd12308, 16'd12996, 16'd45230, 16'd57521, 16'd10711, 16'd49364, 16'd7201, 16'd64439, 16'd3297, 16'd22862, 16'd27640, 16'd53439, 16'd10794, 16'd7134, 16'd2377, 16'd25483, 16'd58349, 16'd10809, 16'd15845, 16'd43406, 16'd46185, 16'd9658, 16'd23158, 16'd38760});
	test_expansion(128'h1b9d83f55952aad9e371ffcccb327142, {16'd29416, 16'd50610, 16'd2124, 16'd57471, 16'd53652, 16'd23701, 16'd37930, 16'd3123, 16'd43485, 16'd10770, 16'd33285, 16'd45821, 16'd16014, 16'd11616, 16'd54436, 16'd35911, 16'd7229, 16'd8097, 16'd42127, 16'd45845, 16'd23379, 16'd11210, 16'd29237, 16'd56179, 16'd38244, 16'd63632});
	test_expansion(128'h11e4e68e15c29156ff080ae6fad993e5, {16'd52060, 16'd61387, 16'd10524, 16'd25384, 16'd21269, 16'd54911, 16'd34067, 16'd40721, 16'd54071, 16'd7268, 16'd52708, 16'd25193, 16'd33082, 16'd16350, 16'd11435, 16'd11396, 16'd25100, 16'd43806, 16'd61904, 16'd32344, 16'd48830, 16'd50381, 16'd10716, 16'd38502, 16'd61831, 16'd7781});
	test_expansion(128'h771a7d60788f4969a06322d76c51e89b, {16'd2609, 16'd55710, 16'd63180, 16'd54500, 16'd37700, 16'd49637, 16'd54294, 16'd43813, 16'd59333, 16'd58713, 16'd5897, 16'd21345, 16'd11318, 16'd18129, 16'd14325, 16'd21915, 16'd29721, 16'd46951, 16'd47144, 16'd15755, 16'd36790, 16'd32403, 16'd17260, 16'd45166, 16'd64833, 16'd9717});
	test_expansion(128'hc217a02ec11a0262b5dba91144124168, {16'd30793, 16'd32200, 16'd43669, 16'd1887, 16'd22836, 16'd41421, 16'd44721, 16'd50480, 16'd11469, 16'd63772, 16'd29261, 16'd56245, 16'd10915, 16'd49879, 16'd18461, 16'd46175, 16'd1380, 16'd46641, 16'd46006, 16'd52816, 16'd62088, 16'd56313, 16'd35250, 16'd40473, 16'd19034, 16'd18514});
	test_expansion(128'h3277ec7b1d66c994f766fdfa63f0b9c5, {16'd53751, 16'd13443, 16'd64113, 16'd15896, 16'd40360, 16'd62074, 16'd10611, 16'd54852, 16'd8686, 16'd21641, 16'd33288, 16'd57182, 16'd11732, 16'd35652, 16'd18476, 16'd28179, 16'd63263, 16'd61568, 16'd9175, 16'd21521, 16'd25075, 16'd55422, 16'd33641, 16'd57738, 16'd46402, 16'd1245});
	test_expansion(128'hbee37cc037b776f02c19dc1ac0a74881, {16'd63820, 16'd48373, 16'd42358, 16'd32076, 16'd11791, 16'd5270, 16'd57828, 16'd9093, 16'd58624, 16'd40942, 16'd31338, 16'd979, 16'd15704, 16'd61509, 16'd46666, 16'd26393, 16'd10419, 16'd17478, 16'd38801, 16'd15868, 16'd56986, 16'd64356, 16'd18001, 16'd33823, 16'd45399, 16'd40519});
	test_expansion(128'hf4d2b4a265410ec79470a8b9e4d801bb, {16'd37824, 16'd64339, 16'd64836, 16'd57182, 16'd61197, 16'd25259, 16'd62232, 16'd19830, 16'd30540, 16'd15204, 16'd58262, 16'd27698, 16'd10019, 16'd24143, 16'd57892, 16'd61088, 16'd12250, 16'd16473, 16'd34491, 16'd45748, 16'd32524, 16'd17758, 16'd23658, 16'd11273, 16'd10700, 16'd1593});
	test_expansion(128'h44450d3c69e532e07bf5ec61f7a12c36, {16'd4786, 16'd15090, 16'd37633, 16'd25891, 16'd42176, 16'd34527, 16'd14632, 16'd27567, 16'd44639, 16'd54590, 16'd54132, 16'd20229, 16'd15219, 16'd28667, 16'd8156, 16'd23098, 16'd10766, 16'd64272, 16'd57184, 16'd28173, 16'd7782, 16'd48331, 16'd42243, 16'd4286, 16'd34892, 16'd1842});
	test_expansion(128'he77f8a19dcaecda64842b4602bb6d870, {16'd54164, 16'd37101, 16'd19318, 16'd50198, 16'd4886, 16'd21734, 16'd103, 16'd24393, 16'd27096, 16'd56351, 16'd13225, 16'd59377, 16'd43355, 16'd24367, 16'd55771, 16'd34177, 16'd15570, 16'd65254, 16'd447, 16'd65056, 16'd28478, 16'd40987, 16'd6503, 16'd11295, 16'd50504, 16'd58943});
	test_expansion(128'h46bc13b247ea4ae29e2c25f180a1d034, {16'd14877, 16'd37244, 16'd52250, 16'd13039, 16'd62678, 16'd25652, 16'd50728, 16'd51315, 16'd37175, 16'd48162, 16'd2429, 16'd51447, 16'd21080, 16'd52504, 16'd12871, 16'd37642, 16'd2487, 16'd61479, 16'd23058, 16'd15754, 16'd49472, 16'd6833, 16'd3734, 16'd42420, 16'd51846, 16'd36721});
	test_expansion(128'h1e9d080843e16fa18fcbd28509c9e297, {16'd32723, 16'd48886, 16'd9066, 16'd52819, 16'd62563, 16'd7419, 16'd9504, 16'd34734, 16'd46930, 16'd39419, 16'd4316, 16'd4803, 16'd31158, 16'd56722, 16'd50415, 16'd10031, 16'd14826, 16'd21935, 16'd1852, 16'd10281, 16'd6763, 16'd52143, 16'd1029, 16'd21201, 16'd19444, 16'd24550});
	test_expansion(128'hd99290ac7e11be0b510b01e0fa3e8d8b, {16'd53171, 16'd63996, 16'd29552, 16'd8216, 16'd35535, 16'd43097, 16'd22567, 16'd4930, 16'd60530, 16'd10824, 16'd5023, 16'd9441, 16'd45270, 16'd8376, 16'd52753, 16'd57640, 16'd5437, 16'd39904, 16'd18550, 16'd32680, 16'd35414, 16'd54342, 16'd32774, 16'd4627, 16'd44401, 16'd47551});
	test_expansion(128'h255782436b0772befc5defc11b2ef56f, {16'd7957, 16'd43457, 16'd22415, 16'd44231, 16'd27018, 16'd3952, 16'd34172, 16'd22341, 16'd6083, 16'd26240, 16'd59586, 16'd57479, 16'd53323, 16'd52339, 16'd36684, 16'd9448, 16'd4798, 16'd44590, 16'd52842, 16'd43522, 16'd50550, 16'd26477, 16'd61416, 16'd25660, 16'd15746, 16'd49292});
	test_expansion(128'h9201171d8504c8bf02e872a83d24c951, {16'd14146, 16'd54785, 16'd55773, 16'd35357, 16'd57810, 16'd27149, 16'd301, 16'd42806, 16'd15552, 16'd24870, 16'd64373, 16'd10818, 16'd46582, 16'd61507, 16'd8946, 16'd39540, 16'd35262, 16'd42241, 16'd23078, 16'd18666, 16'd60611, 16'd13837, 16'd63149, 16'd12679, 16'd17189, 16'd31987});
	test_expansion(128'h02d3fff2afcbbf049985d2a87ccfda11, {16'd16355, 16'd45061, 16'd18593, 16'd23196, 16'd16365, 16'd38320, 16'd25031, 16'd49162, 16'd11330, 16'd33117, 16'd56325, 16'd42365, 16'd20340, 16'd8269, 16'd33004, 16'd25965, 16'd58452, 16'd60776, 16'd37686, 16'd28301, 16'd44716, 16'd21966, 16'd11104, 16'd59244, 16'd28765, 16'd60129});
	test_expansion(128'h73f1a3a1e2941ed293de646cfd937e33, {16'd36163, 16'd61429, 16'd17174, 16'd40414, 16'd42703, 16'd16343, 16'd37530, 16'd22700, 16'd41759, 16'd14276, 16'd51019, 16'd21427, 16'd16771, 16'd38349, 16'd42108, 16'd11796, 16'd11899, 16'd31451, 16'd11686, 16'd23921, 16'd20639, 16'd25466, 16'd63997, 16'd15285, 16'd5971, 16'd52320});
	test_expansion(128'h830cb3aa50fd76ef009f30114a65bfe5, {16'd47336, 16'd28938, 16'd65368, 16'd1051, 16'd41621, 16'd28439, 16'd47775, 16'd43931, 16'd43482, 16'd15796, 16'd40747, 16'd21424, 16'd56372, 16'd4520, 16'd13978, 16'd56394, 16'd2518, 16'd18038, 16'd36835, 16'd54408, 16'd29191, 16'd64233, 16'd61359, 16'd10692, 16'd29935, 16'd36186});
	test_expansion(128'ha2e267d3a9d264be855ffd013808b566, {16'd50118, 16'd48085, 16'd52072, 16'd58707, 16'd9397, 16'd19705, 16'd45840, 16'd41458, 16'd23360, 16'd23819, 16'd27355, 16'd21514, 16'd57850, 16'd25014, 16'd9835, 16'd24446, 16'd28735, 16'd50975, 16'd23773, 16'd41685, 16'd47521, 16'd57277, 16'd50360, 16'd34943, 16'd4653, 16'd12857});
	test_expansion(128'h1758930ec19a997b96dec75f2300afe6, {16'd33555, 16'd38789, 16'd534, 16'd7011, 16'd40589, 16'd30333, 16'd38343, 16'd16086, 16'd21865, 16'd37994, 16'd50074, 16'd40870, 16'd23936, 16'd16884, 16'd17704, 16'd25537, 16'd2090, 16'd43076, 16'd51614, 16'd12388, 16'd30793, 16'd2919, 16'd36858, 16'd35090, 16'd14555, 16'd16430});
	test_expansion(128'hbc08e475dcfbf72c86468556906c47da, {16'd46937, 16'd51257, 16'd12743, 16'd25350, 16'd53001, 16'd5036, 16'd4157, 16'd59849, 16'd47722, 16'd37227, 16'd14658, 16'd56842, 16'd20486, 16'd45024, 16'd13383, 16'd63929, 16'd6398, 16'd10781, 16'd50564, 16'd36878, 16'd27064, 16'd28049, 16'd24374, 16'd40471, 16'd12162, 16'd43770});
	test_expansion(128'h2793d0625e558073fc1292163641afa0, {16'd39333, 16'd14717, 16'd40862, 16'd22577, 16'd44709, 16'd43821, 16'd52153, 16'd44812, 16'd39798, 16'd45382, 16'd55658, 16'd21254, 16'd28120, 16'd21979, 16'd56009, 16'd56753, 16'd14390, 16'd58580, 16'd64106, 16'd12660, 16'd36352, 16'd36926, 16'd32184, 16'd42898, 16'd33410, 16'd22959});
	test_expansion(128'h800c78f6f09014be68668346a759006e, {16'd38138, 16'd38825, 16'd12805, 16'd50039, 16'd45259, 16'd64028, 16'd15043, 16'd29570, 16'd45728, 16'd18041, 16'd44033, 16'd39452, 16'd27227, 16'd25077, 16'd26803, 16'd16253, 16'd36157, 16'd8479, 16'd48876, 16'd22700, 16'd23492, 16'd23627, 16'd3616, 16'd31833, 16'd25939, 16'd4692});
	test_expansion(128'h9bdc357f386298cbcffe75467dfa1919, {16'd58020, 16'd50932, 16'd26054, 16'd19249, 16'd55087, 16'd9123, 16'd27184, 16'd23938, 16'd20476, 16'd34385, 16'd51297, 16'd19662, 16'd16069, 16'd17333, 16'd19156, 16'd46486, 16'd33447, 16'd57083, 16'd14256, 16'd25047, 16'd58472, 16'd17141, 16'd20792, 16'd16751, 16'd33775, 16'd56377});
	test_expansion(128'hbb461d8933793bbc19f505effab045b3, {16'd21384, 16'd2539, 16'd47887, 16'd44213, 16'd53915, 16'd44324, 16'd45747, 16'd61067, 16'd59731, 16'd25244, 16'd17327, 16'd58484, 16'd36090, 16'd42095, 16'd58946, 16'd14087, 16'd12087, 16'd22829, 16'd18089, 16'd41585, 16'd1109, 16'd28618, 16'd65499, 16'd31374, 16'd1133, 16'd16437});
	test_expansion(128'h85c243cbca37a54438e837d530376af7, {16'd5443, 16'd55170, 16'd41255, 16'd57006, 16'd32172, 16'd27651, 16'd13984, 16'd4042, 16'd41469, 16'd50667, 16'd23665, 16'd64399, 16'd13676, 16'd3173, 16'd35424, 16'd38460, 16'd37275, 16'd64749, 16'd40119, 16'd24018, 16'd35188, 16'd30801, 16'd14345, 16'd14396, 16'd19959, 16'd14435});
	test_expansion(128'h20742e528d12dc313ee8d96c3fa77f1b, {16'd29736, 16'd4047, 16'd48128, 16'd65279, 16'd46174, 16'd34583, 16'd34611, 16'd52176, 16'd25437, 16'd16598, 16'd27360, 16'd60023, 16'd51567, 16'd3865, 16'd61082, 16'd44649, 16'd8991, 16'd26282, 16'd4479, 16'd23039, 16'd46271, 16'd50509, 16'd47817, 16'd46565, 16'd28294, 16'd45393});
	test_expansion(128'hec986cff81df35be8f8eba7c4dcd1927, {16'd19758, 16'd33621, 16'd34971, 16'd39138, 16'd40610, 16'd44210, 16'd41729, 16'd38813, 16'd43368, 16'd44692, 16'd8255, 16'd28670, 16'd47880, 16'd18651, 16'd52666, 16'd17763, 16'd7484, 16'd10353, 16'd50799, 16'd17758, 16'd5220, 16'd45497, 16'd51652, 16'd57495, 16'd11862, 16'd16845});
	test_expansion(128'h6827b6c00aaf970bec6dc9390f26574b, {16'd51268, 16'd62718, 16'd38371, 16'd60000, 16'd46486, 16'd27519, 16'd8766, 16'd15959, 16'd28684, 16'd48546, 16'd32761, 16'd61308, 16'd35591, 16'd39250, 16'd34467, 16'd2288, 16'd34029, 16'd17536, 16'd4296, 16'd18641, 16'd59988, 16'd18714, 16'd45105, 16'd48439, 16'd50611, 16'd22410});
	test_expansion(128'hb6e1d6b3765d36bdc56ebdf94f558525, {16'd30361, 16'd23497, 16'd21459, 16'd60650, 16'd19984, 16'd65039, 16'd14114, 16'd42462, 16'd29643, 16'd18542, 16'd12065, 16'd23332, 16'd4092, 16'd45829, 16'd3063, 16'd27727, 16'd30512, 16'd37991, 16'd19820, 16'd31220, 16'd7805, 16'd41687, 16'd812, 16'd37863, 16'd43809, 16'd7392});
	test_expansion(128'h80d84e8fd46b603ff0c3f78a0fd96d68, {16'd17824, 16'd63249, 16'd64347, 16'd37441, 16'd53692, 16'd52656, 16'd51882, 16'd24486, 16'd48976, 16'd62850, 16'd34275, 16'd56324, 16'd60968, 16'd17388, 16'd60670, 16'd31332, 16'd21186, 16'd28109, 16'd44422, 16'd8386, 16'd2738, 16'd16547, 16'd44674, 16'd31760, 16'd61004, 16'd12390});
	test_expansion(128'h509b2d7c6d73d6f94efbdf58c3102c9e, {16'd18040, 16'd10006, 16'd30829, 16'd22917, 16'd45022, 16'd55612, 16'd64423, 16'd2741, 16'd19165, 16'd20885, 16'd38218, 16'd16765, 16'd56373, 16'd19124, 16'd23283, 16'd17488, 16'd56948, 16'd43246, 16'd16149, 16'd25859, 16'd57781, 16'd57825, 16'd19142, 16'd28261, 16'd19003, 16'd4226});
	test_expansion(128'h127d828b6d60f8feb320fcfcb62c1a39, {16'd58479, 16'd36536, 16'd52450, 16'd26141, 16'd53656, 16'd26034, 16'd14740, 16'd59710, 16'd47850, 16'd54865, 16'd11643, 16'd41128, 16'd35513, 16'd271, 16'd36119, 16'd38203, 16'd46922, 16'd24828, 16'd1312, 16'd23663, 16'd512, 16'd30609, 16'd30333, 16'd32787, 16'd65356, 16'd16768});
	test_expansion(128'hf5efe7afb13ec8ce7138135e8b9a6c4f, {16'd5279, 16'd6457, 16'd18422, 16'd11467, 16'd137, 16'd36566, 16'd61339, 16'd50138, 16'd42154, 16'd35248, 16'd21092, 16'd10838, 16'd7667, 16'd59005, 16'd1187, 16'd12527, 16'd33510, 16'd59906, 16'd7948, 16'd41572, 16'd3157, 16'd3684, 16'd36463, 16'd9089, 16'd33001, 16'd48469});
	test_expansion(128'h12e63492eacb11d9c31cecad1281ccc7, {16'd22368, 16'd26863, 16'd37684, 16'd16290, 16'd60594, 16'd41271, 16'd58140, 16'd28700, 16'd21706, 16'd5792, 16'd53757, 16'd48980, 16'd27566, 16'd38290, 16'd37422, 16'd42860, 16'd16864, 16'd33754, 16'd3303, 16'd5054, 16'd8936, 16'd10016, 16'd7549, 16'd39137, 16'd40901, 16'd58650});
	test_expansion(128'h5fc4a471e4f793ab5f2b0fd6cb918126, {16'd14492, 16'd31906, 16'd45039, 16'd41569, 16'd38506, 16'd33483, 16'd14624, 16'd18946, 16'd27447, 16'd57966, 16'd5822, 16'd31769, 16'd33831, 16'd28655, 16'd64737, 16'd48341, 16'd22390, 16'd7690, 16'd29955, 16'd8141, 16'd46502, 16'd50468, 16'd59553, 16'd59636, 16'd47438, 16'd51063});
	test_expansion(128'hace608637d2feafa1a890c6754efcfb5, {16'd57032, 16'd17471, 16'd57669, 16'd20493, 16'd64262, 16'd30940, 16'd21109, 16'd44091, 16'd795, 16'd895, 16'd31938, 16'd6633, 16'd32997, 16'd31214, 16'd39714, 16'd30964, 16'd61139, 16'd46106, 16'd31580, 16'd2515, 16'd40474, 16'd42678, 16'd7483, 16'd53259, 16'd4744, 16'd50837});
	test_expansion(128'h429ea6b722ecab8a20fdc8bdda88fee1, {16'd36233, 16'd3466, 16'd24920, 16'd26915, 16'd55537, 16'd15634, 16'd54723, 16'd26990, 16'd33355, 16'd60256, 16'd5935, 16'd37556, 16'd36046, 16'd4849, 16'd20860, 16'd30486, 16'd23822, 16'd10174, 16'd17600, 16'd3098, 16'd60270, 16'd52015, 16'd56301, 16'd47481, 16'd64486, 16'd29677});
	test_expansion(128'he02cfc2acec54892292437fd4c56b444, {16'd8604, 16'd31467, 16'd51125, 16'd27099, 16'd51183, 16'd46687, 16'd20306, 16'd16668, 16'd47831, 16'd38619, 16'd9461, 16'd51796, 16'd28717, 16'd23968, 16'd65304, 16'd12787, 16'd28379, 16'd15368, 16'd61958, 16'd47663, 16'd40700, 16'd20027, 16'd30384, 16'd42024, 16'd20605, 16'd18823});
	test_expansion(128'h2d49e35dc2fab50744dadf6acadef0c0, {16'd18227, 16'd62140, 16'd54582, 16'd57511, 16'd11459, 16'd64289, 16'd3593, 16'd40105, 16'd60458, 16'd3023, 16'd52827, 16'd36447, 16'd7931, 16'd20421, 16'd43605, 16'd8255, 16'd62857, 16'd29463, 16'd55319, 16'd61370, 16'd14295, 16'd55673, 16'd29369, 16'd24601, 16'd16558, 16'd65052});
	test_expansion(128'h9f7f714feebcac628683bb663cd771fc, {16'd21739, 16'd3183, 16'd56464, 16'd13631, 16'd38275, 16'd37183, 16'd3172, 16'd3794, 16'd29951, 16'd31678, 16'd44553, 16'd48961, 16'd41347, 16'd54231, 16'd36386, 16'd10804, 16'd3385, 16'd34207, 16'd33760, 16'd1900, 16'd65070, 16'd6428, 16'd52155, 16'd42776, 16'd58965, 16'd1844});
	test_expansion(128'h0f3fb7ab7ddbc62556e489dcec880576, {16'd55501, 16'd34292, 16'd5360, 16'd28362, 16'd57306, 16'd29435, 16'd8314, 16'd55220, 16'd18886, 16'd46219, 16'd60226, 16'd2796, 16'd58062, 16'd12642, 16'd13599, 16'd65460, 16'd57258, 16'd15381, 16'd7159, 16'd58673, 16'd56717, 16'd61796, 16'd28194, 16'd4790, 16'd7241, 16'd63658});
	test_expansion(128'h5320780b651d94af078b7e3922456d5c, {16'd62303, 16'd43275, 16'd21299, 16'd47060, 16'd38274, 16'd57291, 16'd30524, 16'd38583, 16'd33209, 16'd57475, 16'd45040, 16'd64778, 16'd13661, 16'd48599, 16'd18011, 16'd19269, 16'd59514, 16'd25170, 16'd5263, 16'd48981, 16'd13740, 16'd62022, 16'd2497, 16'd11851, 16'd11933, 16'd934});
	test_expansion(128'h5cca362576c7d28b5ca9c7b5e7fee188, {16'd25473, 16'd57380, 16'd113, 16'd15675, 16'd28442, 16'd11193, 16'd37634, 16'd37645, 16'd55971, 16'd24050, 16'd54328, 16'd33237, 16'd3163, 16'd60511, 16'd26572, 16'd55810, 16'd25981, 16'd15856, 16'd45645, 16'd4170, 16'd11035, 16'd39114, 16'd44562, 16'd44206, 16'd37134, 16'd64725});
	test_expansion(128'h250c0e1a5e090945c24500501ad5ae81, {16'd12163, 16'd12722, 16'd29076, 16'd40369, 16'd39470, 16'd20977, 16'd10430, 16'd17099, 16'd6148, 16'd42956, 16'd18923, 16'd51048, 16'd29957, 16'd65427, 16'd30597, 16'd18942, 16'd32261, 16'd21619, 16'd35237, 16'd31542, 16'd16081, 16'd52641, 16'd18731, 16'd31853, 16'd15328, 16'd57370});
	test_expansion(128'hbc1666205c1189f4b60bbb5f0b75fb35, {16'd34787, 16'd48029, 16'd31296, 16'd3169, 16'd46163, 16'd45268, 16'd24200, 16'd6217, 16'd36246, 16'd42860, 16'd28713, 16'd54593, 16'd43945, 16'd2494, 16'd11026, 16'd62233, 16'd56188, 16'd34834, 16'd5490, 16'd43459, 16'd8439, 16'd62704, 16'd7896, 16'd47532, 16'd46693, 16'd45939});
	test_expansion(128'h1d6f6ccc102c97f16adab97a2885dc12, {16'd28234, 16'd28262, 16'd697, 16'd18280, 16'd35127, 16'd29744, 16'd44422, 16'd20382, 16'd57263, 16'd33377, 16'd21060, 16'd19989, 16'd37416, 16'd42581, 16'd53852, 16'd42238, 16'd62088, 16'd2785, 16'd29194, 16'd31568, 16'd3523, 16'd38394, 16'd54229, 16'd40077, 16'd14883, 16'd39553});
	test_expansion(128'h2cf2fec1c75e43b43ecc4eed59d07535, {16'd37566, 16'd49107, 16'd40794, 16'd59525, 16'd11107, 16'd8901, 16'd40832, 16'd59727, 16'd44319, 16'd17456, 16'd13488, 16'd62338, 16'd42159, 16'd9358, 16'd25078, 16'd34432, 16'd56874, 16'd23466, 16'd27864, 16'd53985, 16'd44592, 16'd54444, 16'd3806, 16'd4236, 16'd10107, 16'd48263});
	test_expansion(128'haf03e07788a5bfc6abe9d9fbdaac931e, {16'd34348, 16'd27134, 16'd25298, 16'd33401, 16'd27664, 16'd38562, 16'd44517, 16'd3606, 16'd55408, 16'd65357, 16'd58142, 16'd2660, 16'd17674, 16'd60868, 16'd58627, 16'd7496, 16'd32266, 16'd54063, 16'd48682, 16'd47569, 16'd48766, 16'd22971, 16'd14521, 16'd16045, 16'd29664, 16'd57213});
	test_expansion(128'h1a0dd51bd1a43d652b1bcce2d10e5085, {16'd45499, 16'd23694, 16'd35539, 16'd53903, 16'd31142, 16'd15960, 16'd12370, 16'd65048, 16'd7107, 16'd17011, 16'd56121, 16'd29558, 16'd17639, 16'd28058, 16'd60430, 16'd59353, 16'd39526, 16'd39981, 16'd56271, 16'd43891, 16'd46335, 16'd3794, 16'd57023, 16'd1808, 16'd48713, 16'd57458});
	test_expansion(128'h43c278e9cf493db4a9a31f05e195ef9c, {16'd18756, 16'd50483, 16'd26139, 16'd26449, 16'd1872, 16'd15203, 16'd2981, 16'd22963, 16'd21687, 16'd23965, 16'd60472, 16'd22124, 16'd19020, 16'd35578, 16'd21740, 16'd48361, 16'd44747, 16'd53373, 16'd43888, 16'd22267, 16'd40461, 16'd8395, 16'd30928, 16'd19530, 16'd17995, 16'd64649});
	test_expansion(128'h73984002d45e256657ac81102e654630, {16'd12470, 16'd36108, 16'd52007, 16'd6730, 16'd45252, 16'd51037, 16'd2281, 16'd26325, 16'd20186, 16'd53120, 16'd57123, 16'd60337, 16'd50024, 16'd47267, 16'd46740, 16'd8862, 16'd34094, 16'd59944, 16'd48957, 16'd61109, 16'd14845, 16'd31880, 16'd28232, 16'd21919, 16'd8930, 16'd38643});
	test_expansion(128'h35968749e090ed62b0f04de9c23e61cc, {16'd44439, 16'd15975, 16'd47670, 16'd47638, 16'd24264, 16'd7318, 16'd60601, 16'd40704, 16'd37999, 16'd30300, 16'd42440, 16'd5187, 16'd46294, 16'd40881, 16'd26904, 16'd8541, 16'd50463, 16'd35767, 16'd20711, 16'd46090, 16'd8247, 16'd21010, 16'd43493, 16'd59070, 16'd25445, 16'd35442});
	test_expansion(128'h36d673129708ed6289cd13919c97d4b9, {16'd6497, 16'd19467, 16'd59344, 16'd46004, 16'd56161, 16'd53046, 16'd41518, 16'd4798, 16'd62879, 16'd20433, 16'd18055, 16'd5282, 16'd47321, 16'd17084, 16'd65431, 16'd45081, 16'd15343, 16'd62667, 16'd45877, 16'd21928, 16'd19848, 16'd60898, 16'd1459, 16'd8908, 16'd34964, 16'd9871});
	test_expansion(128'h9abb807e86ffe961b46226fa4620ebf4, {16'd35184, 16'd8105, 16'd39606, 16'd26958, 16'd25597, 16'd49308, 16'd8315, 16'd33705, 16'd5809, 16'd40804, 16'd37612, 16'd37596, 16'd38173, 16'd42158, 16'd19029, 16'd5914, 16'd14451, 16'd60098, 16'd13516, 16'd52606, 16'd33977, 16'd14091, 16'd4971, 16'd17421, 16'd45798, 16'd31558});
	test_expansion(128'h4a19106a659075f849f22d72b0a2b199, {16'd5924, 16'd41349, 16'd21792, 16'd24984, 16'd9169, 16'd32115, 16'd13313, 16'd52301, 16'd65241, 16'd16731, 16'd36855, 16'd45670, 16'd36458, 16'd60883, 16'd29881, 16'd65521, 16'd45799, 16'd46876, 16'd28699, 16'd42215, 16'd58411, 16'd35835, 16'd49324, 16'd33582, 16'd33873, 16'd44280});
	test_expansion(128'h4a3987a63870ac71b12589b917e40190, {16'd4415, 16'd9283, 16'd25647, 16'd20390, 16'd10988, 16'd53034, 16'd41178, 16'd44113, 16'd62806, 16'd22270, 16'd19731, 16'd4147, 16'd50144, 16'd48685, 16'd61198, 16'd56293, 16'd2897, 16'd12340, 16'd6119, 16'd19033, 16'd63738, 16'd57111, 16'd4616, 16'd46464, 16'd47272, 16'd55663});
	test_expansion(128'h22472957a43286c3330efbbf3ebebf70, {16'd44918, 16'd22997, 16'd10258, 16'd18646, 16'd57746, 16'd35748, 16'd38813, 16'd25797, 16'd16018, 16'd54443, 16'd15284, 16'd33964, 16'd56786, 16'd37625, 16'd63902, 16'd14957, 16'd24397, 16'd50946, 16'd2763, 16'd51944, 16'd44612, 16'd53932, 16'd61533, 16'd35458, 16'd23094, 16'd3139});
	test_expansion(128'h94d94b968238e5d82696938f7928d4fc, {16'd41620, 16'd62020, 16'd62719, 16'd64166, 16'd276, 16'd50167, 16'd26295, 16'd1337, 16'd48790, 16'd14840, 16'd43709, 16'd38438, 16'd41814, 16'd38624, 16'd34976, 16'd46234, 16'd47643, 16'd14519, 16'd27484, 16'd43713, 16'd50764, 16'd35112, 16'd3667, 16'd22803, 16'd19928, 16'd4513});
	test_expansion(128'ha7c68448bdcb11469ea43e22fd26739f, {16'd25036, 16'd26902, 16'd30021, 16'd45779, 16'd38817, 16'd26491, 16'd53417, 16'd13063, 16'd7917, 16'd48945, 16'd43930, 16'd11745, 16'd15403, 16'd38245, 16'd52153, 16'd59724, 16'd3037, 16'd14204, 16'd14814, 16'd49764, 16'd49642, 16'd1060, 16'd35440, 16'd27900, 16'd44491, 16'd35064});
	test_expansion(128'h1854b7733b57673ae4106dc53f14f832, {16'd21070, 16'd27367, 16'd42648, 16'd63489, 16'd9075, 16'd51534, 16'd9020, 16'd22471, 16'd43468, 16'd42768, 16'd3136, 16'd6665, 16'd43079, 16'd28480, 16'd23316, 16'd50334, 16'd54402, 16'd27886, 16'd34949, 16'd43192, 16'd437, 16'd35350, 16'd30184, 16'd17318, 16'd14339, 16'd47684});
	test_expansion(128'hc6299ce61f6e6b307ad5493f56af2481, {16'd50690, 16'd1151, 16'd32901, 16'd59453, 16'd22909, 16'd20449, 16'd49222, 16'd40856, 16'd41698, 16'd19836, 16'd41015, 16'd38900, 16'd34056, 16'd59636, 16'd49366, 16'd8082, 16'd8336, 16'd59847, 16'd8309, 16'd46610, 16'd26404, 16'd49920, 16'd14330, 16'd3157, 16'd64174, 16'd25008});
	test_expansion(128'h173ad9e52eef37267eb91d3dccecd1f2, {16'd61702, 16'd18915, 16'd46622, 16'd53505, 16'd21164, 16'd32741, 16'd42801, 16'd7277, 16'd17562, 16'd53346, 16'd57608, 16'd8714, 16'd51324, 16'd59691, 16'd13059, 16'd7339, 16'd38773, 16'd53150, 16'd2949, 16'd18914, 16'd22232, 16'd64863, 16'd10247, 16'd44829, 16'd23826, 16'd46444});
	test_expansion(128'h1c1f5130ada12e878ed4d6e85af8c9f7, {16'd11896, 16'd12799, 16'd33495, 16'd58465, 16'd5858, 16'd4700, 16'd2072, 16'd29327, 16'd48920, 16'd21977, 16'd58991, 16'd55335, 16'd37996, 16'd22861, 16'd34085, 16'd15825, 16'd4, 16'd38643, 16'd33071, 16'd45200, 16'd56165, 16'd38750, 16'd31261, 16'd31392, 16'd30015, 16'd238});
	test_expansion(128'h37986b4b393c5322692be40835526dc8, {16'd29896, 16'd24625, 16'd37501, 16'd57457, 16'd21657, 16'd1099, 16'd13448, 16'd58066, 16'd53014, 16'd57701, 16'd53512, 16'd63214, 16'd11256, 16'd325, 16'd56689, 16'd54843, 16'd34065, 16'd57336, 16'd28794, 16'd18103, 16'd27659, 16'd57746, 16'd15769, 16'd45378, 16'd16058, 16'd32106});
	test_expansion(128'h4951de01ce98e20be8475d1ccc2f77df, {16'd18415, 16'd4533, 16'd6346, 16'd9151, 16'd50713, 16'd59623, 16'd39206, 16'd2793, 16'd61596, 16'd4718, 16'd6041, 16'd4687, 16'd21531, 16'd34430, 16'd50047, 16'd43724, 16'd47200, 16'd8958, 16'd10139, 16'd40204, 16'd38491, 16'd49414, 16'd34272, 16'd53358, 16'd25673, 16'd41124});
	test_expansion(128'h4bbfc6cc24a03e90740a249eb64b48ea, {16'd58715, 16'd61356, 16'd4806, 16'd23125, 16'd17099, 16'd63958, 16'd7602, 16'd37341, 16'd50724, 16'd47995, 16'd61872, 16'd40831, 16'd4947, 16'd54565, 16'd48977, 16'd48767, 16'd14943, 16'd40277, 16'd57285, 16'd3907, 16'd9088, 16'd34089, 16'd49488, 16'd48669, 16'd45571, 16'd38836});
	test_expansion(128'h8a26211d7895a4938c1d99c946175812, {16'd19218, 16'd26770, 16'd37544, 16'd37497, 16'd6302, 16'd12637, 16'd65439, 16'd16851, 16'd9940, 16'd3651, 16'd25781, 16'd63663, 16'd39201, 16'd41312, 16'd50362, 16'd34235, 16'd35980, 16'd51577, 16'd9993, 16'd4272, 16'd12710, 16'd63283, 16'd65277, 16'd11563, 16'd50596, 16'd43438});
	test_expansion(128'hea481ac297c89c6938b5bd1d30118c72, {16'd16599, 16'd39472, 16'd33964, 16'd57323, 16'd14599, 16'd50899, 16'd15898, 16'd24308, 16'd1443, 16'd31498, 16'd60625, 16'd23744, 16'd10670, 16'd42565, 16'd33157, 16'd8056, 16'd61044, 16'd62555, 16'd27489, 16'd31474, 16'd57971, 16'd56052, 16'd58703, 16'd29676, 16'd39439, 16'd30109});
	test_expansion(128'h71cf51052f79739b86c765909dbea900, {16'd39785, 16'd49493, 16'd1322, 16'd59821, 16'd28365, 16'd52035, 16'd16055, 16'd39434, 16'd28803, 16'd30418, 16'd20633, 16'd49039, 16'd8744, 16'd40122, 16'd51516, 16'd32224, 16'd9859, 16'd54117, 16'd40054, 16'd58074, 16'd34230, 16'd997, 16'd28319, 16'd40152, 16'd57358, 16'd45150});
	test_expansion(128'h6e9d6749329b432cf28d54b5068cb1f7, {16'd9227, 16'd33815, 16'd26944, 16'd42932, 16'd21627, 16'd15038, 16'd40992, 16'd17945, 16'd32137, 16'd4836, 16'd7165, 16'd57561, 16'd59246, 16'd38527, 16'd1603, 16'd1554, 16'd49200, 16'd49092, 16'd45451, 16'd33180, 16'd13586, 16'd38959, 16'd31096, 16'd58137, 16'd51792, 16'd45619});
	test_expansion(128'h7ff19acc96074517f5af8f2e5fe0ad70, {16'd28130, 16'd1707, 16'd3444, 16'd60611, 16'd41205, 16'd57176, 16'd56986, 16'd28085, 16'd54283, 16'd23877, 16'd62580, 16'd54695, 16'd62936, 16'd8892, 16'd6439, 16'd11620, 16'd27256, 16'd55445, 16'd37097, 16'd51702, 16'd43456, 16'd56889, 16'd45640, 16'd36702, 16'd44673, 16'd26931});
	test_expansion(128'h274cb15542654f19fccebfdf69e2bb27, {16'd51186, 16'd20758, 16'd52529, 16'd51587, 16'd46715, 16'd22733, 16'd5832, 16'd21718, 16'd17121, 16'd46124, 16'd24688, 16'd10596, 16'd1831, 16'd16139, 16'd3848, 16'd54498, 16'd8683, 16'd8772, 16'd10680, 16'd64443, 16'd59360, 16'd28319, 16'd43133, 16'd448, 16'd64351, 16'd32425});
	test_expansion(128'hc5f4cbe724dbce6e88540945575c4757, {16'd33901, 16'd60578, 16'd3632, 16'd48466, 16'd57059, 16'd62108, 16'd23716, 16'd18083, 16'd42756, 16'd3522, 16'd49023, 16'd56763, 16'd4895, 16'd13801, 16'd177, 16'd6584, 16'd24182, 16'd20335, 16'd19629, 16'd62977, 16'd51535, 16'd5887, 16'd19165, 16'd22798, 16'd40113, 16'd37542});
	test_expansion(128'h91fddaf3d23fe293274cf73655a1bb7c, {16'd58451, 16'd25402, 16'd3084, 16'd3051, 16'd34135, 16'd47772, 16'd40805, 16'd19865, 16'd745, 16'd25388, 16'd12292, 16'd22268, 16'd46889, 16'd42594, 16'd49691, 16'd48989, 16'd399, 16'd10777, 16'd63136, 16'd1241, 16'd36717, 16'd7317, 16'd30160, 16'd37947, 16'd62667, 16'd49405});
	test_expansion(128'h4bb4dc88481f4320a214035d601a7759, {16'd54789, 16'd54324, 16'd21998, 16'd8545, 16'd16257, 16'd19362, 16'd11947, 16'd31059, 16'd2021, 16'd16905, 16'd30425, 16'd18781, 16'd37999, 16'd59678, 16'd21100, 16'd56600, 16'd4924, 16'd20810, 16'd12017, 16'd17688, 16'd5840, 16'd1246, 16'd45186, 16'd44275, 16'd8091, 16'd36555});
	test_expansion(128'h11aff0c4769235c6e04f9ee2e88afe8c, {16'd52509, 16'd35692, 16'd45977, 16'd20156, 16'd50559, 16'd35552, 16'd11871, 16'd34504, 16'd34073, 16'd5841, 16'd19308, 16'd28329, 16'd15469, 16'd3413, 16'd38516, 16'd46466, 16'd63387, 16'd12109, 16'd5785, 16'd61691, 16'd44537, 16'd44257, 16'd64778, 16'd2158, 16'd41863, 16'd39191});
	test_expansion(128'h0cd3aea7ac63f196e6f3eae5d7671412, {16'd57559, 16'd57816, 16'd22432, 16'd15911, 16'd64416, 16'd5139, 16'd6800, 16'd38414, 16'd10689, 16'd36414, 16'd50871, 16'd33454, 16'd3946, 16'd62303, 16'd26406, 16'd33513, 16'd28568, 16'd54270, 16'd34223, 16'd53716, 16'd28889, 16'd37831, 16'd17554, 16'd28053, 16'd50756, 16'd7673});
	test_expansion(128'h25ca04de23c1928371344af2af9d8ad5, {16'd6323, 16'd34551, 16'd898, 16'd41777, 16'd18433, 16'd28459, 16'd38148, 16'd18191, 16'd1527, 16'd4729, 16'd42728, 16'd47363, 16'd47738, 16'd4564, 16'd20681, 16'd14469, 16'd38882, 16'd7994, 16'd64572, 16'd51662, 16'd13599, 16'd43551, 16'd31239, 16'd30098, 16'd61134, 16'd62715});
	test_expansion(128'h7a9bbc22ce9b7890c2e1a4112bfe3e1a, {16'd32358, 16'd3690, 16'd29527, 16'd52871, 16'd13426, 16'd6392, 16'd54520, 16'd18433, 16'd25733, 16'd18464, 16'd29530, 16'd33927, 16'd1827, 16'd50903, 16'd49516, 16'd27213, 16'd61413, 16'd53271, 16'd59513, 16'd42176, 16'd61223, 16'd14878, 16'd56883, 16'd61473, 16'd35602, 16'd1202});
	test_expansion(128'h3e23011e71d7169553f25a59bdaacf7b, {16'd56476, 16'd20679, 16'd49222, 16'd42955, 16'd58585, 16'd51971, 16'd1123, 16'd30923, 16'd58902, 16'd2052, 16'd19813, 16'd28761, 16'd20811, 16'd19711, 16'd16029, 16'd60254, 16'd11219, 16'd17819, 16'd6877, 16'd12356, 16'd50094, 16'd8427, 16'd7412, 16'd33137, 16'd38218, 16'd19352});
	test_expansion(128'h1902640b6380063c1ee11806e90f2b97, {16'd35821, 16'd48159, 16'd45564, 16'd45936, 16'd37572, 16'd57201, 16'd5989, 16'd28857, 16'd39623, 16'd27399, 16'd41057, 16'd24902, 16'd1718, 16'd33744, 16'd16547, 16'd19615, 16'd17241, 16'd59449, 16'd48283, 16'd8427, 16'd62507, 16'd61938, 16'd13413, 16'd56301, 16'd42009, 16'd46196});
	test_expansion(128'h1f95630ca8ee7ffd33ba9d9463540525, {16'd46610, 16'd23468, 16'd15936, 16'd36271, 16'd14200, 16'd2822, 16'd16247, 16'd60662, 16'd16269, 16'd64689, 16'd65056, 16'd44900, 16'd57218, 16'd46525, 16'd46551, 16'd48192, 16'd41008, 16'd42314, 16'd59706, 16'd13837, 16'd61162, 16'd4349, 16'd18040, 16'd50447, 16'd41157, 16'd37236});
	test_expansion(128'h6e3c698592276b85b5d1715b381bfdd7, {16'd22252, 16'd42700, 16'd9805, 16'd1403, 16'd33530, 16'd56087, 16'd40161, 16'd50057, 16'd7682, 16'd1526, 16'd20717, 16'd29186, 16'd21663, 16'd25993, 16'd32564, 16'd13765, 16'd7520, 16'd42055, 16'd3381, 16'd7586, 16'd47780, 16'd38713, 16'd10142, 16'd63738, 16'd61060, 16'd39241});
	test_expansion(128'h41e3926064ec310fdc67115f547cfc8b, {16'd48138, 16'd39992, 16'd61795, 16'd45377, 16'd36885, 16'd28210, 16'd60676, 16'd7165, 16'd52583, 16'd39005, 16'd58591, 16'd57685, 16'd45065, 16'd32680, 16'd5760, 16'd14371, 16'd55744, 16'd5426, 16'd44528, 16'd32421, 16'd62580, 16'd17088, 16'd58234, 16'd13803, 16'd5767, 16'd22079});
	test_expansion(128'h0adf149017dd952ec51642870d45ca32, {16'd1692, 16'd41670, 16'd41912, 16'd23741, 16'd59311, 16'd46483, 16'd27097, 16'd18768, 16'd4188, 16'd9200, 16'd31673, 16'd31287, 16'd11389, 16'd62842, 16'd5650, 16'd20676, 16'd23991, 16'd26339, 16'd54003, 16'd61072, 16'd12622, 16'd51989, 16'd40287, 16'd55840, 16'd41284, 16'd10301});
	test_expansion(128'h5d5f440a77846e1fdc16de0d328ddca2, {16'd17180, 16'd60865, 16'd43944, 16'd28163, 16'd11674, 16'd2564, 16'd59485, 16'd65276, 16'd23928, 16'd41595, 16'd37706, 16'd32782, 16'd36283, 16'd9970, 16'd32144, 16'd49433, 16'd51789, 16'd37110, 16'd12033, 16'd51315, 16'd10167, 16'd13949, 16'd29924, 16'd44488, 16'd34500, 16'd28392});
	test_expansion(128'h3e872f82b80c50101fe36910289f1df5, {16'd59980, 16'd29013, 16'd20384, 16'd55368, 16'd17176, 16'd39196, 16'd12282, 16'd32007, 16'd32391, 16'd39690, 16'd15844, 16'd62063, 16'd53840, 16'd11376, 16'd47710, 16'd51870, 16'd44002, 16'd41910, 16'd10281, 16'd5873, 16'd50591, 16'd17954, 16'd34301, 16'd13580, 16'd55470, 16'd15770});
	test_expansion(128'h2a64d09623b749090c6cd3ba26e21c53, {16'd5267, 16'd58954, 16'd25761, 16'd62893, 16'd24891, 16'd45659, 16'd8426, 16'd39275, 16'd29292, 16'd15451, 16'd48320, 16'd55385, 16'd34192, 16'd1997, 16'd60217, 16'd56500, 16'd55716, 16'd52693, 16'd26780, 16'd50016, 16'd42670, 16'd64850, 16'd34440, 16'd7013, 16'd20153, 16'd43009});
	test_expansion(128'hf895c50e49497b2abad9de4bda919333, {16'd44544, 16'd12673, 16'd53705, 16'd1402, 16'd47118, 16'd14304, 16'd1551, 16'd46115, 16'd53806, 16'd46487, 16'd32964, 16'd5397, 16'd44045, 16'd33306, 16'd13924, 16'd13274, 16'd38790, 16'd52865, 16'd7047, 16'd28794, 16'd5230, 16'd34365, 16'd4429, 16'd57137, 16'd47413, 16'd45203});
	test_expansion(128'he0b426f7707794dc1f1c01ad49e4c3cf, {16'd3269, 16'd39177, 16'd60351, 16'd27518, 16'd19735, 16'd20416, 16'd14253, 16'd38159, 16'd51381, 16'd43827, 16'd51116, 16'd5640, 16'd63361, 16'd34401, 16'd59607, 16'd2417, 16'd17152, 16'd37958, 16'd4562, 16'd18150, 16'd56164, 16'd27225, 16'd26823, 16'd16183, 16'd22455, 16'd15276});
	test_expansion(128'h6c9c8078902e5d6efea1b17c218dd904, {16'd33592, 16'd10640, 16'd59521, 16'd21455, 16'd44350, 16'd6690, 16'd39551, 16'd21951, 16'd19676, 16'd29177, 16'd49464, 16'd53152, 16'd24643, 16'd44460, 16'd56150, 16'd25529, 16'd48763, 16'd16230, 16'd48893, 16'd54750, 16'd59636, 16'd16464, 16'd58022, 16'd38793, 16'd19047, 16'd65277});
	test_expansion(128'hcfff512c733a7bb0c88dbca0fba8fe12, {16'd22519, 16'd63274, 16'd36018, 16'd58152, 16'd45487, 16'd22529, 16'd5557, 16'd17613, 16'd63932, 16'd25949, 16'd65503, 16'd16611, 16'd53029, 16'd58135, 16'd42924, 16'd33339, 16'd11973, 16'd61163, 16'd16539, 16'd23764, 16'd4276, 16'd520, 16'd877, 16'd8838, 16'd46488, 16'd14324});
	test_expansion(128'he0c41f7279a53773ea80519dc3df8dac, {16'd29893, 16'd2263, 16'd52280, 16'd9982, 16'd7661, 16'd49126, 16'd13774, 16'd38344, 16'd46557, 16'd7591, 16'd26082, 16'd34494, 16'd32963, 16'd22153, 16'd5817, 16'd23743, 16'd47600, 16'd59608, 16'd4572, 16'd4840, 16'd2116, 16'd24326, 16'd62442, 16'd8822, 16'd13729, 16'd63622});
	test_expansion(128'h40030760f1fc17888720dacc5a48b39d, {16'd6116, 16'd44865, 16'd19548, 16'd18400, 16'd5362, 16'd43354, 16'd41333, 16'd7169, 16'd17522, 16'd61213, 16'd18872, 16'd27966, 16'd43099, 16'd11502, 16'd39390, 16'd9228, 16'd10288, 16'd47494, 16'd33482, 16'd59472, 16'd53000, 16'd43794, 16'd56565, 16'd18278, 16'd15701, 16'd32538});
	test_expansion(128'he8377c79436db57b58435570cb922d05, {16'd15884, 16'd31387, 16'd56924, 16'd59719, 16'd41669, 16'd52300, 16'd3462, 16'd12872, 16'd50172, 16'd253, 16'd22548, 16'd17058, 16'd28939, 16'd31579, 16'd4206, 16'd41298, 16'd28059, 16'd40108, 16'd13845, 16'd33634, 16'd53654, 16'd39225, 16'd42448, 16'd56018, 16'd32436, 16'd40123});
	test_expansion(128'hfb1aacbb0d603b706a64ec2d38d4d256, {16'd29804, 16'd42028, 16'd34145, 16'd62972, 16'd1181, 16'd11721, 16'd30737, 16'd46191, 16'd27120, 16'd18431, 16'd53753, 16'd7455, 16'd59048, 16'd27545, 16'd49948, 16'd20401, 16'd37872, 16'd10162, 16'd37168, 16'd56892, 16'd21514, 16'd20682, 16'd45900, 16'd64535, 16'd60136, 16'd42246});
	test_expansion(128'hb49f0ae259b8f53aadd1d3c39b741b14, {16'd61188, 16'd17180, 16'd14854, 16'd37525, 16'd58924, 16'd10700, 16'd12971, 16'd49520, 16'd39787, 16'd36958, 16'd25289, 16'd22000, 16'd64879, 16'd31463, 16'd47732, 16'd32310, 16'd29554, 16'd56887, 16'd64932, 16'd24044, 16'd58248, 16'd45496, 16'd10775, 16'd15637, 16'd42374, 16'd53620});
	test_expansion(128'hd47e2130562bda83e451738f4a2b9a8f, {16'd48699, 16'd1846, 16'd1384, 16'd61308, 16'd63980, 16'd34210, 16'd34627, 16'd45911, 16'd55051, 16'd23945, 16'd44410, 16'd12284, 16'd28264, 16'd12605, 16'd20149, 16'd52814, 16'd56968, 16'd48754, 16'd28289, 16'd23103, 16'd58616, 16'd12847, 16'd17871, 16'd39647, 16'd38937, 16'd8973});
	test_expansion(128'hf8b65b2e0f9cd41144ca3d7ca6d91dc1, {16'd44330, 16'd10858, 16'd54517, 16'd3165, 16'd5751, 16'd63018, 16'd23894, 16'd47367, 16'd59258, 16'd18482, 16'd11826, 16'd11961, 16'd41158, 16'd63192, 16'd61277, 16'd10750, 16'd36337, 16'd47495, 16'd53153, 16'd49661, 16'd10683, 16'd9066, 16'd34783, 16'd30283, 16'd11581, 16'd36263});
	test_expansion(128'h32223ad236aa64b05e6d603db188d9c9, {16'd38666, 16'd4599, 16'd40766, 16'd13532, 16'd15523, 16'd45309, 16'd44017, 16'd15909, 16'd41187, 16'd52926, 16'd8802, 16'd11273, 16'd58875, 16'd59728, 16'd47235, 16'd25610, 16'd6552, 16'd22669, 16'd61768, 16'd41528, 16'd5723, 16'd47095, 16'd43169, 16'd5053, 16'd45556, 16'd33507});
	test_expansion(128'h3238f8ee223b5157edad20f48ec3d425, {16'd59081, 16'd1171, 16'd6920, 16'd7699, 16'd30940, 16'd25758, 16'd48581, 16'd48904, 16'd7753, 16'd4734, 16'd36263, 16'd30193, 16'd36477, 16'd26474, 16'd42005, 16'd43319, 16'd43892, 16'd58508, 16'd62722, 16'd31297, 16'd10621, 16'd38996, 16'd32959, 16'd1474, 16'd34872, 16'd13455});
	test_expansion(128'h848ef4fe09e7c33cc1731c6c12372702, {16'd20232, 16'd7205, 16'd50769, 16'd10278, 16'd28379, 16'd18438, 16'd55353, 16'd53594, 16'd47222, 16'd64627, 16'd2836, 16'd26212, 16'd11279, 16'd55700, 16'd50699, 16'd21808, 16'd60407, 16'd1460, 16'd45218, 16'd12873, 16'd37558, 16'd45963, 16'd46744, 16'd42628, 16'd4175, 16'd18247});
	test_expansion(128'h71c9733276d18efa154b7a3731dfa1e0, {16'd48363, 16'd38769, 16'd10437, 16'd63541, 16'd10243, 16'd43749, 16'd9011, 16'd28461, 16'd49403, 16'd33248, 16'd19675, 16'd8622, 16'd3059, 16'd26248, 16'd63797, 16'd33488, 16'd37346, 16'd64647, 16'd57711, 16'd21932, 16'd10106, 16'd29072, 16'd47608, 16'd63405, 16'd59918, 16'd4042});
	test_expansion(128'hff136c22734edb5034893fbe17a5cfdf, {16'd60922, 16'd22753, 16'd21338, 16'd4014, 16'd33924, 16'd29589, 16'd63437, 16'd24355, 16'd54504, 16'd18653, 16'd64869, 16'd60513, 16'd28447, 16'd5896, 16'd11127, 16'd33619, 16'd4530, 16'd33427, 16'd58836, 16'd19330, 16'd20198, 16'd24804, 16'd63959, 16'd47250, 16'd62457, 16'd37022});
	test_expansion(128'h0fb9bd663e5c241e3c7a7cd549bf3095, {16'd39639, 16'd23776, 16'd55329, 16'd28274, 16'd22745, 16'd13976, 16'd54824, 16'd5743, 16'd9102, 16'd61001, 16'd1707, 16'd34248, 16'd48844, 16'd38171, 16'd35935, 16'd53542, 16'd24640, 16'd50186, 16'd48231, 16'd18746, 16'd32560, 16'd21692, 16'd40985, 16'd39600, 16'd43899, 16'd10504});
	test_expansion(128'h4bd5607cce3ffb568b0f8c0bebf42dd8, {16'd36076, 16'd25768, 16'd9271, 16'd34338, 16'd40248, 16'd54325, 16'd40446, 16'd34820, 16'd4845, 16'd14545, 16'd59362, 16'd14656, 16'd35105, 16'd32697, 16'd20344, 16'd62848, 16'd5884, 16'd28880, 16'd24792, 16'd14175, 16'd26324, 16'd11919, 16'd440, 16'd12928, 16'd52422, 16'd45290});
	test_expansion(128'hc5f2295137032144481cd4f72f629db6, {16'd62209, 16'd47875, 16'd6435, 16'd53728, 16'd41309, 16'd12340, 16'd54242, 16'd11674, 16'd24959, 16'd16760, 16'd56733, 16'd63833, 16'd13676, 16'd44800, 16'd2567, 16'd64283, 16'd27173, 16'd44197, 16'd36941, 16'd27986, 16'd39544, 16'd38829, 16'd43888, 16'd55261, 16'd4928, 16'd38586});
	test_expansion(128'h64f6b3033609aede89abe734a4eda19f, {16'd30696, 16'd23397, 16'd23622, 16'd58409, 16'd6838, 16'd11365, 16'd44174, 16'd13808, 16'd35432, 16'd14792, 16'd60543, 16'd15845, 16'd43542, 16'd49371, 16'd33825, 16'd19069, 16'd53518, 16'd61437, 16'd2800, 16'd34076, 16'd11281, 16'd48325, 16'd8449, 16'd16604, 16'd48410, 16'd36813});
	test_expansion(128'hd415679f2ae02cf88391165f7ee10e50, {16'd25083, 16'd45704, 16'd17570, 16'd60, 16'd30997, 16'd24819, 16'd21901, 16'd37282, 16'd39319, 16'd63944, 16'd55171, 16'd31732, 16'd34293, 16'd39565, 16'd16720, 16'd714, 16'd47254, 16'd57437, 16'd54508, 16'd48328, 16'd50186, 16'd23515, 16'd4958, 16'd50752, 16'd59177, 16'd2917});
	test_expansion(128'h8e07642ba4b22e044f10d2843fd0c125, {16'd44137, 16'd40305, 16'd12716, 16'd59091, 16'd29726, 16'd37896, 16'd14777, 16'd39152, 16'd61061, 16'd34360, 16'd46911, 16'd31508, 16'd17379, 16'd32565, 16'd2562, 16'd3671, 16'd58002, 16'd30128, 16'd45899, 16'd30655, 16'd11417, 16'd8154, 16'd59150, 16'd10612, 16'd8236, 16'd45646});
	test_expansion(128'hd00f219961c9df745789b458a9fa5de9, {16'd32440, 16'd48173, 16'd24046, 16'd42483, 16'd27276, 16'd20623, 16'd42182, 16'd52850, 16'd32915, 16'd41157, 16'd43139, 16'd54529, 16'd31960, 16'd60761, 16'd33654, 16'd57455, 16'd60427, 16'd46337, 16'd48066, 16'd33814, 16'd51717, 16'd59754, 16'd45503, 16'd11275, 16'd57463, 16'd63458});
	test_expansion(128'h0aa10c1f6f2783f518f1309dfeaa917d, {16'd47898, 16'd48923, 16'd45915, 16'd39706, 16'd29309, 16'd47306, 16'd11512, 16'd4504, 16'd26217, 16'd39048, 16'd42144, 16'd18985, 16'd23846, 16'd51160, 16'd6916, 16'd48967, 16'd39092, 16'd61888, 16'd14744, 16'd64611, 16'd15452, 16'd5959, 16'd60447, 16'd15739, 16'd11074, 16'd44725});
	test_expansion(128'h3dd2a1e724c5d43db6edd4dd61bd54b3, {16'd41311, 16'd29722, 16'd40212, 16'd54821, 16'd15057, 16'd6996, 16'd31164, 16'd51573, 16'd4969, 16'd54275, 16'd1801, 16'd14807, 16'd47095, 16'd1758, 16'd13612, 16'd17281, 16'd31198, 16'd38086, 16'd26856, 16'd1311, 16'd30412, 16'd48411, 16'd64568, 16'd39917, 16'd64742, 16'd44063});
	test_expansion(128'hb5c162c958f71682783b3f50bf03dfa4, {16'd51079, 16'd64142, 16'd35092, 16'd25225, 16'd20045, 16'd6372, 16'd43147, 16'd45453, 16'd20403, 16'd30553, 16'd6458, 16'd19398, 16'd47620, 16'd55696, 16'd31266, 16'd2057, 16'd31246, 16'd33111, 16'd53271, 16'd3723, 16'd250, 16'd44319, 16'd49573, 16'd46348, 16'd59710, 16'd25397});
	test_expansion(128'h4bba6eb793da8d69f49f3d54fde71440, {16'd4848, 16'd701, 16'd49107, 16'd55423, 16'd55815, 16'd31950, 16'd50775, 16'd40293, 16'd8534, 16'd37927, 16'd33599, 16'd9531, 16'd38715, 16'd34224, 16'd11313, 16'd6580, 16'd8072, 16'd17456, 16'd35385, 16'd49362, 16'd36525, 16'd65018, 16'd13065, 16'd59593, 16'd5190, 16'd63156});
	test_expansion(128'h6c353e07ceb20adf470e11e7cebd8c6a, {16'd13455, 16'd12337, 16'd29607, 16'd17435, 16'd6571, 16'd37781, 16'd55229, 16'd52498, 16'd62934, 16'd31658, 16'd53306, 16'd3491, 16'd15744, 16'd15177, 16'd3504, 16'd42560, 16'd16566, 16'd23784, 16'd13182, 16'd40527, 16'd61207, 16'd26612, 16'd54976, 16'd9955, 16'd32058, 16'd8092});
	test_expansion(128'hc976ce3f76117b335f00b3733a24942c, {16'd57991, 16'd34887, 16'd17072, 16'd37436, 16'd46029, 16'd32108, 16'd33078, 16'd44722, 16'd21730, 16'd19481, 16'd17619, 16'd43803, 16'd42989, 16'd36656, 16'd13820, 16'd39833, 16'd61074, 16'd56603, 16'd37234, 16'd38558, 16'd42504, 16'd33109, 16'd41783, 16'd813, 16'd26282, 16'd13066});
	test_expansion(128'h57c10a526aa6743d4cf107793c25db79, {16'd56270, 16'd62845, 16'd52172, 16'd22823, 16'd39065, 16'd7090, 16'd40261, 16'd21282, 16'd38766, 16'd8940, 16'd35519, 16'd51870, 16'd19047, 16'd10972, 16'd5723, 16'd22460, 16'd34264, 16'd6805, 16'd61594, 16'd16403, 16'd20158, 16'd22352, 16'd15133, 16'd53930, 16'd46482, 16'd38183});
	test_expansion(128'hfa437c017da9f9abaaf2c53101c30a34, {16'd59778, 16'd9400, 16'd16392, 16'd50037, 16'd23588, 16'd38589, 16'd50987, 16'd50678, 16'd27889, 16'd59989, 16'd49236, 16'd60826, 16'd59304, 16'd12259, 16'd39114, 16'd65315, 16'd13578, 16'd45135, 16'd33366, 16'd29009, 16'd59825, 16'd37033, 16'd29493, 16'd15580, 16'd2503, 16'd35465});
	test_expansion(128'h36d21d1d4a1d97b5240f1cbb18b7e0da, {16'd34823, 16'd65262, 16'd61081, 16'd56274, 16'd32054, 16'd7120, 16'd40089, 16'd17774, 16'd31473, 16'd62903, 16'd49693, 16'd31337, 16'd27210, 16'd32457, 16'd56123, 16'd10939, 16'd64601, 16'd47843, 16'd9159, 16'd38473, 16'd20399, 16'd17591, 16'd12262, 16'd7148, 16'd13808, 16'd40726});
	test_expansion(128'h065ffd0b0539680b68e5cd2357e9c9cb, {16'd36218, 16'd59435, 16'd19170, 16'd56969, 16'd61286, 16'd29580, 16'd17272, 16'd48619, 16'd16043, 16'd1866, 16'd38193, 16'd11162, 16'd3289, 16'd40199, 16'd2795, 16'd18545, 16'd13552, 16'd2368, 16'd8820, 16'd8368, 16'd52618, 16'd31663, 16'd63959, 16'd30273, 16'd1417, 16'd40147});
	test_expansion(128'h68dc1f2a9ffcda8e6af01cf0e5f55155, {16'd16460, 16'd32491, 16'd53223, 16'd5256, 16'd49589, 16'd9568, 16'd21288, 16'd39739, 16'd56071, 16'd12811, 16'd10304, 16'd17496, 16'd52965, 16'd6621, 16'd39561, 16'd21005, 16'd33456, 16'd24212, 16'd5124, 16'd26715, 16'd47686, 16'd850, 16'd2621, 16'd43505, 16'd60042, 16'd58835});
	test_expansion(128'h27b712ef52da3f4be53a46fcd6ed93e2, {16'd17756, 16'd56495, 16'd13774, 16'd58343, 16'd33022, 16'd61204, 16'd33869, 16'd63488, 16'd4151, 16'd37300, 16'd43964, 16'd59230, 16'd64681, 16'd60029, 16'd36186, 16'd61424, 16'd7610, 16'd25923, 16'd35857, 16'd60747, 16'd6867, 16'd44123, 16'd6103, 16'd11630, 16'd25236, 16'd62152});
	test_expansion(128'hdf8b6cf97026ff2542820fc5e3c4e877, {16'd3212, 16'd45221, 16'd49753, 16'd48022, 16'd19263, 16'd31440, 16'd57942, 16'd30532, 16'd15861, 16'd9551, 16'd26688, 16'd1524, 16'd15235, 16'd5511, 16'd40360, 16'd35747, 16'd42515, 16'd32470, 16'd4704, 16'd42032, 16'd33849, 16'd9169, 16'd35253, 16'd32824, 16'd16708, 16'd6731});
	test_expansion(128'h7797672b2b5ecd878f95a134f4f0b07d, {16'd45329, 16'd38773, 16'd50385, 16'd32310, 16'd25929, 16'd43552, 16'd45410, 16'd42394, 16'd34718, 16'd29579, 16'd55947, 16'd37062, 16'd36069, 16'd15596, 16'd46964, 16'd9976, 16'd47672, 16'd39561, 16'd38777, 16'd14146, 16'd26201, 16'd44386, 16'd16321, 16'd18385, 16'd2285, 16'd63324});
	test_expansion(128'haf5f5f30e4b29d4275a5a51db271a7b5, {16'd26573, 16'd48036, 16'd52248, 16'd16270, 16'd52420, 16'd25856, 16'd25301, 16'd25932, 16'd37242, 16'd49716, 16'd32335, 16'd10840, 16'd10294, 16'd28794, 16'd65195, 16'd54884, 16'd15775, 16'd46234, 16'd14217, 16'd55882, 16'd17767, 16'd42297, 16'd34054, 16'd45310, 16'd55142, 16'd3259});
	test_expansion(128'h5a20d5283b2145dad4f2b6b4bd7f86d1, {16'd17391, 16'd50173, 16'd38341, 16'd23543, 16'd52604, 16'd33566, 16'd24141, 16'd49662, 16'd45723, 16'd8087, 16'd43304, 16'd4562, 16'd24360, 16'd21030, 16'd62156, 16'd42202, 16'd59270, 16'd50531, 16'd42168, 16'd61220, 16'd25793, 16'd49592, 16'd55496, 16'd52208, 16'd26555, 16'd37363});
	test_expansion(128'ha902ff7be78cf4240e488dd90285dbf0, {16'd44295, 16'd46173, 16'd37645, 16'd56587, 16'd37794, 16'd49227, 16'd11449, 16'd57786, 16'd515, 16'd16889, 16'd24965, 16'd33231, 16'd55804, 16'd56721, 16'd54418, 16'd31916, 16'd22273, 16'd8385, 16'd21432, 16'd17470, 16'd64756, 16'd10660, 16'd18517, 16'd20309, 16'd65305, 16'd20509});
	test_expansion(128'hecb66576784bc16afa1d85d449eca472, {16'd50615, 16'd61520, 16'd33848, 16'd45884, 16'd22616, 16'd36273, 16'd53061, 16'd50660, 16'd64433, 16'd53761, 16'd59715, 16'd39322, 16'd30151, 16'd17491, 16'd54128, 16'd14150, 16'd33362, 16'd10665, 16'd50250, 16'd5737, 16'd38426, 16'd43824, 16'd22389, 16'd12700, 16'd57072, 16'd23026});
	test_expansion(128'h4efabca001d9bbb56f2dd4772c7667ee, {16'd43719, 16'd60865, 16'd52953, 16'd19973, 16'd62521, 16'd50128, 16'd43569, 16'd29498, 16'd4720, 16'd1005, 16'd27217, 16'd15403, 16'd5181, 16'd1804, 16'd46337, 16'd19202, 16'd35857, 16'd53523, 16'd49486, 16'd2339, 16'd37618, 16'd2222, 16'd33054, 16'd13032, 16'd27786, 16'd53363});
	test_expansion(128'h12d932498b2441e10d6d7e7375c4f3d7, {16'd22088, 16'd42567, 16'd64079, 16'd58826, 16'd41466, 16'd12203, 16'd54114, 16'd56706, 16'd39374, 16'd20817, 16'd63679, 16'd20567, 16'd4235, 16'd27458, 16'd41322, 16'd52983, 16'd21484, 16'd1665, 16'd10744, 16'd11184, 16'd31832, 16'd20505, 16'd12960, 16'd19376, 16'd1136, 16'd11665});
	test_expansion(128'h5c1ee7239de355a53d8235d75b9cfef8, {16'd49094, 16'd37736, 16'd33188, 16'd52879, 16'd128, 16'd62875, 16'd58223, 16'd13471, 16'd13891, 16'd60042, 16'd35704, 16'd31904, 16'd44428, 16'd3973, 16'd9973, 16'd32991, 16'd22583, 16'd32752, 16'd38384, 16'd5283, 16'd30249, 16'd18148, 16'd31367, 16'd17803, 16'd3606, 16'd3298});
	test_expansion(128'ha065d068ed7bd28e0e1d80bd8650d532, {16'd11959, 16'd10857, 16'd13678, 16'd31192, 16'd26169, 16'd6491, 16'd19115, 16'd26057, 16'd7755, 16'd38236, 16'd62802, 16'd25623, 16'd5404, 16'd14264, 16'd38225, 16'd25733, 16'd17009, 16'd27045, 16'd53435, 16'd44573, 16'd17551, 16'd58485, 16'd37646, 16'd54415, 16'd34399, 16'd31440});
	test_expansion(128'he8245220ff61351190b95ae84152217c, {16'd63187, 16'd5051, 16'd10600, 16'd34672, 16'd10766, 16'd16505, 16'd17826, 16'd51241, 16'd38871, 16'd48443, 16'd22115, 16'd708, 16'd9155, 16'd13168, 16'd19171, 16'd17953, 16'd13399, 16'd7240, 16'd58771, 16'd11075, 16'd17045, 16'd57454, 16'd32219, 16'd35099, 16'd17615, 16'd50961});
	test_expansion(128'hf9cd5e364b7eaca93b7c288c495cc19a, {16'd48125, 16'd35962, 16'd7749, 16'd41584, 16'd35776, 16'd30624, 16'd20989, 16'd20224, 16'd41487, 16'd52408, 16'd47577, 16'd41855, 16'd7655, 16'd5338, 16'd14260, 16'd60049, 16'd27568, 16'd742, 16'd19347, 16'd40015, 16'd56853, 16'd41423, 16'd2063, 16'd40558, 16'd33671, 16'd41932});
	test_expansion(128'h6fdcde684bf7bc8e9cb81596a8f37e96, {16'd38889, 16'd21018, 16'd481, 16'd13837, 16'd61485, 16'd4899, 16'd56722, 16'd4953, 16'd7097, 16'd30476, 16'd23491, 16'd29165, 16'd6994, 16'd23991, 16'd61838, 16'd62749, 16'd21924, 16'd64954, 16'd6494, 16'd20237, 16'd19762, 16'd39540, 16'd12861, 16'd26438, 16'd51623, 16'd15416});
	test_expansion(128'hefb41bdcaac901677a4257f230d920b1, {16'd50835, 16'd12791, 16'd10343, 16'd50314, 16'd42016, 16'd44694, 16'd47157, 16'd13756, 16'd29044, 16'd50312, 16'd59591, 16'd12821, 16'd33629, 16'd35489, 16'd61317, 16'd50671, 16'd3217, 16'd23048, 16'd47062, 16'd31437, 16'd58449, 16'd54564, 16'd59738, 16'd14234, 16'd25004, 16'd143});
	test_expansion(128'h9c46e0ec49c8dd2a4d4b4badf3fff24d, {16'd53511, 16'd58195, 16'd40426, 16'd40452, 16'd32121, 16'd1884, 16'd51189, 16'd44486, 16'd391, 16'd47606, 16'd21295, 16'd13432, 16'd7137, 16'd30544, 16'd30798, 16'd46058, 16'd16641, 16'd24185, 16'd6959, 16'd53888, 16'd24323, 16'd55892, 16'd6381, 16'd2777, 16'd8899, 16'd6189});
	test_expansion(128'h2196411798d8b77073d2ddd78587c62c, {16'd19268, 16'd38700, 16'd44804, 16'd26277, 16'd45554, 16'd28476, 16'd35507, 16'd48547, 16'd37078, 16'd40992, 16'd33464, 16'd46563, 16'd16367, 16'd1700, 16'd58032, 16'd25305, 16'd56299, 16'd21782, 16'd8828, 16'd55672, 16'd60065, 16'd2468, 16'd30542, 16'd42792, 16'd17981, 16'd15463});
	test_expansion(128'hbc37b544bdd3feb989ec5b1080a47569, {16'd56708, 16'd35609, 16'd42779, 16'd16968, 16'd28517, 16'd53574, 16'd61808, 16'd5253, 16'd51647, 16'd15497, 16'd28164, 16'd4681, 16'd61370, 16'd30602, 16'd60061, 16'd25610, 16'd24515, 16'd63117, 16'd15155, 16'd43060, 16'd26945, 16'd30494, 16'd60334, 16'd38835, 16'd45676, 16'd49211});
	test_expansion(128'h1c2faf02fd0c46b9b5aa64c23ed1fca4, {16'd9651, 16'd50727, 16'd14780, 16'd60369, 16'd37398, 16'd16720, 16'd30784, 16'd7644, 16'd23283, 16'd59478, 16'd51464, 16'd28604, 16'd6424, 16'd44217, 16'd13823, 16'd1130, 16'd63470, 16'd51336, 16'd44540, 16'd38868, 16'd61347, 16'd43328, 16'd34582, 16'd64168, 16'd5765, 16'd1142});
	test_expansion(128'h8331f18845f40996afbd7a542156cff2, {16'd34934, 16'd13568, 16'd19625, 16'd30339, 16'd20148, 16'd1312, 16'd7738, 16'd62273, 16'd23417, 16'd29068, 16'd37791, 16'd13651, 16'd24021, 16'd9650, 16'd17798, 16'd32092, 16'd16450, 16'd41304, 16'd60662, 16'd26571, 16'd16635, 16'd61165, 16'd47636, 16'd25275, 16'd22646, 16'd47576});
	test_expansion(128'h541c87c45859b8a62a7c20f065a9da71, {16'd7227, 16'd35129, 16'd15722, 16'd20785, 16'd57438, 16'd53166, 16'd63136, 16'd28177, 16'd16644, 16'd31668, 16'd57504, 16'd3021, 16'd47449, 16'd29584, 16'd49445, 16'd28852, 16'd36996, 16'd29285, 16'd22066, 16'd6487, 16'd60817, 16'd58430, 16'd302, 16'd32570, 16'd2351, 16'd4643});
	test_expansion(128'h40788e7f7a527f4d4282ef67603af9d5, {16'd22314, 16'd26939, 16'd64402, 16'd48833, 16'd30073, 16'd22035, 16'd825, 16'd10397, 16'd26529, 16'd41944, 16'd3624, 16'd58760, 16'd16166, 16'd29234, 16'd4765, 16'd15757, 16'd15471, 16'd11493, 16'd57453, 16'd45985, 16'd19061, 16'd18869, 16'd25867, 16'd51724, 16'd48622, 16'd42780});
	test_expansion(128'h78a789946032a82528edcf61b8fb21cc, {16'd41259, 16'd42322, 16'd14488, 16'd63180, 16'd51108, 16'd6120, 16'd28399, 16'd28913, 16'd18559, 16'd50251, 16'd58171, 16'd41650, 16'd6721, 16'd61174, 16'd33986, 16'd43234, 16'd798, 16'd30889, 16'd2943, 16'd29382, 16'd42980, 16'd27466, 16'd53989, 16'd35915, 16'd47123, 16'd3852});
	test_expansion(128'he6f7ecf7c883f305da2f360d1500c249, {16'd11052, 16'd43937, 16'd52960, 16'd33499, 16'd47436, 16'd7387, 16'd1767, 16'd56201, 16'd25164, 16'd41274, 16'd12452, 16'd48196, 16'd32503, 16'd28724, 16'd55522, 16'd40664, 16'd15504, 16'd58528, 16'd32389, 16'd26799, 16'd10150, 16'd43348, 16'd33588, 16'd15777, 16'd11339, 16'd34909});
	test_expansion(128'hc4ec243dd0c24070fb21a9a5d9de8bb3, {16'd418, 16'd12035, 16'd62173, 16'd32131, 16'd863, 16'd21820, 16'd28813, 16'd64040, 16'd14331, 16'd49049, 16'd19441, 16'd9301, 16'd28477, 16'd6258, 16'd10862, 16'd6534, 16'd48170, 16'd3097, 16'd43261, 16'd13120, 16'd36257, 16'd31791, 16'd52889, 16'd45068, 16'd52934, 16'd6209});
	test_expansion(128'h2e735dc1eed0b50612e2cc0a50e18206, {16'd26656, 16'd4116, 16'd46830, 16'd60791, 16'd42744, 16'd36782, 16'd40309, 16'd27736, 16'd2871, 16'd6270, 16'd58159, 16'd43951, 16'd773, 16'd100, 16'd59575, 16'd25378, 16'd53893, 16'd59319, 16'd55667, 16'd27297, 16'd5785, 16'd52873, 16'd46295, 16'd56070, 16'd65041, 16'd61270});
	test_expansion(128'h2f281cccc96c92d87cd4ab16424e5764, {16'd17318, 16'd30904, 16'd5894, 16'd22550, 16'd65052, 16'd3630, 16'd5829, 16'd35021, 16'd17559, 16'd49024, 16'd53990, 16'd44321, 16'd29609, 16'd60940, 16'd33458, 16'd41561, 16'd42186, 16'd56703, 16'd9149, 16'd44619, 16'd58663, 16'd55900, 16'd61428, 16'd38814, 16'd20748, 16'd19866});
	test_expansion(128'h9aafc3a07696f36f20a1a6e0a868c5de, {16'd37773, 16'd3053, 16'd64897, 16'd55197, 16'd583, 16'd49488, 16'd11824, 16'd15914, 16'd53214, 16'd23031, 16'd30669, 16'd14843, 16'd24549, 16'd8139, 16'd51258, 16'd8034, 16'd20306, 16'd7879, 16'd41733, 16'd29457, 16'd62029, 16'd20800, 16'd15653, 16'd10430, 16'd60778, 16'd60190});
	test_expansion(128'h902401e30c6febba354a5205fc7c9f6c, {16'd18396, 16'd61651, 16'd13548, 16'd51991, 16'd13245, 16'd32164, 16'd16319, 16'd59459, 16'd35313, 16'd34865, 16'd47685, 16'd39126, 16'd8613, 16'd19776, 16'd43374, 16'd64112, 16'd19842, 16'd15984, 16'd24106, 16'd49717, 16'd48526, 16'd19414, 16'd59863, 16'd30339, 16'd33539, 16'd55611});
	test_expansion(128'h5b6cc6678a794cb53b38742ca247ecd4, {16'd21434, 16'd39762, 16'd7417, 16'd7929, 16'd25767, 16'd45678, 16'd31018, 16'd26436, 16'd43340, 16'd4551, 16'd4363, 16'd48759, 16'd10663, 16'd42526, 16'd39484, 16'd27231, 16'd11783, 16'd23447, 16'd12259, 16'd4228, 16'd17651, 16'd28947, 16'd19380, 16'd10055, 16'd9269, 16'd52237});
	test_expansion(128'h130cc31a0afa8c5877deeb572130222c, {16'd32947, 16'd52985, 16'd37234, 16'd61950, 16'd52488, 16'd17420, 16'd50992, 16'd52499, 16'd8095, 16'd51930, 16'd59496, 16'd54566, 16'd45261, 16'd3651, 16'd33510, 16'd5369, 16'd45818, 16'd51289, 16'd10713, 16'd40805, 16'd52732, 16'd7484, 16'd39403, 16'd53058, 16'd52008, 16'd33483});
	test_expansion(128'h14bbe38e755683881ea8aa8f1bc55917, {16'd52180, 16'd1848, 16'd57598, 16'd13211, 16'd11900, 16'd20713, 16'd23366, 16'd3178, 16'd36793, 16'd42927, 16'd26029, 16'd41711, 16'd62096, 16'd41226, 16'd51770, 16'd2898, 16'd53841, 16'd48009, 16'd42722, 16'd50857, 16'd38899, 16'd24829, 16'd52752, 16'd4990, 16'd46175, 16'd3487});
	test_expansion(128'h92ce5d7585c150dd905021978672fef7, {16'd17075, 16'd29431, 16'd3976, 16'd34277, 16'd44911, 16'd11417, 16'd20715, 16'd60108, 16'd21314, 16'd43595, 16'd2109, 16'd39214, 16'd39553, 16'd62651, 16'd19412, 16'd44031, 16'd62565, 16'd10078, 16'd11557, 16'd2362, 16'd8832, 16'd18002, 16'd15741, 16'd29083, 16'd26722, 16'd59494});
	test_expansion(128'ha23371166cb920c4b989f3b5366827e1, {16'd40265, 16'd8917, 16'd14419, 16'd52305, 16'd15058, 16'd54848, 16'd47515, 16'd33348, 16'd31295, 16'd65312, 16'd16913, 16'd15268, 16'd29679, 16'd1758, 16'd42874, 16'd50229, 16'd2572, 16'd54955, 16'd59079, 16'd47886, 16'd30962, 16'd13855, 16'd48231, 16'd58223, 16'd28720, 16'd61419});
	test_expansion(128'hb661571cfe26f671b011738361b65fb8, {16'd7332, 16'd10895, 16'd24690, 16'd47912, 16'd35687, 16'd59229, 16'd314, 16'd50211, 16'd18363, 16'd34362, 16'd18916, 16'd62435, 16'd22571, 16'd39245, 16'd54503, 16'd54089, 16'd5478, 16'd44459, 16'd907, 16'd49431, 16'd2729, 16'd47063, 16'd31917, 16'd22147, 16'd18732, 16'd57811});
	test_expansion(128'h7aa8678ef082eae68fe2cc1e65631c6d, {16'd24724, 16'd15247, 16'd36152, 16'd58294, 16'd42661, 16'd38303, 16'd2238, 16'd1463, 16'd47882, 16'd57253, 16'd30032, 16'd1671, 16'd24454, 16'd2411, 16'd12119, 16'd8719, 16'd64182, 16'd13624, 16'd27640, 16'd29975, 16'd37495, 16'd46924, 16'd47098, 16'd27797, 16'd43586, 16'd40535});
	test_expansion(128'h568d6d2d52572e50e408bcc0737375e8, {16'd55489, 16'd64462, 16'd19597, 16'd2143, 16'd5355, 16'd33621, 16'd40981, 16'd47996, 16'd51717, 16'd36550, 16'd20995, 16'd13291, 16'd37877, 16'd37074, 16'd4127, 16'd8510, 16'd41108, 16'd58007, 16'd18270, 16'd62925, 16'd7149, 16'd35731, 16'd38119, 16'd22850, 16'd21032, 16'd6932});
	test_expansion(128'hae103f2e866e9336128ac73969b055ef, {16'd1414, 16'd10882, 16'd59135, 16'd57820, 16'd12592, 16'd37846, 16'd25026, 16'd44492, 16'd52208, 16'd25170, 16'd26017, 16'd41994, 16'd35557, 16'd22131, 16'd58932, 16'd587, 16'd10294, 16'd63992, 16'd57730, 16'd52439, 16'd11697, 16'd32816, 16'd47699, 16'd22289, 16'd30246, 16'd6328});
	test_expansion(128'hdc6eabae8b7c9ac39926973dec72cead, {16'd55725, 16'd40710, 16'd11110, 16'd38690, 16'd22378, 16'd49928, 16'd29993, 16'd28402, 16'd22631, 16'd52790, 16'd7024, 16'd62089, 16'd57854, 16'd4825, 16'd38839, 16'd57810, 16'd56800, 16'd15179, 16'd53063, 16'd31999, 16'd35427, 16'd51538, 16'd49719, 16'd5572, 16'd40447, 16'd64396});
	test_expansion(128'h1d9a1c3f1191fb753f471d4d5ecdec9d, {16'd53870, 16'd10027, 16'd2193, 16'd23820, 16'd39999, 16'd43421, 16'd7734, 16'd55255, 16'd17535, 16'd41790, 16'd52205, 16'd8791, 16'd28111, 16'd37232, 16'd48779, 16'd31949, 16'd43404, 16'd52156, 16'd17068, 16'd64674, 16'd33978, 16'd35272, 16'd5482, 16'd19665, 16'd50478, 16'd49312});
	test_expansion(128'hac7b7236bd86ec20cbc0e19eadf09013, {16'd36193, 16'd52480, 16'd28382, 16'd55291, 16'd4014, 16'd19877, 16'd18917, 16'd14237, 16'd47617, 16'd42151, 16'd8125, 16'd52467, 16'd50849, 16'd18955, 16'd29131, 16'd64192, 16'd43119, 16'd4315, 16'd65308, 16'd40075, 16'd57596, 16'd43133, 16'd471, 16'd35037, 16'd11909, 16'd42844});
	test_expansion(128'hb46aefd900b91b1ff2024fc0fe488862, {16'd14491, 16'd47754, 16'd49247, 16'd44320, 16'd63882, 16'd38362, 16'd25611, 16'd58497, 16'd62138, 16'd21880, 16'd54610, 16'd31183, 16'd64396, 16'd7082, 16'd51323, 16'd21808, 16'd53060, 16'd32036, 16'd5995, 16'd34294, 16'd26620, 16'd42365, 16'd23619, 16'd11079, 16'd16319, 16'd30099});
	test_expansion(128'h23afc5b2fa056c50cd452d8c94170ccb, {16'd53595, 16'd41511, 16'd24671, 16'd41841, 16'd26886, 16'd63781, 16'd44980, 16'd21379, 16'd59090, 16'd32211, 16'd2025, 16'd33742, 16'd12848, 16'd1733, 16'd2215, 16'd1107, 16'd8737, 16'd35167, 16'd61367, 16'd8249, 16'd16337, 16'd33570, 16'd207, 16'd18414, 16'd41180, 16'd24846});
	test_expansion(128'ha2280b5868827d8bca66f276e6ba9785, {16'd25475, 16'd38839, 16'd36867, 16'd16370, 16'd47745, 16'd30526, 16'd48931, 16'd63307, 16'd8843, 16'd61056, 16'd24913, 16'd5667, 16'd23606, 16'd42967, 16'd57223, 16'd40381, 16'd24901, 16'd10715, 16'd44214, 16'd55269, 16'd56353, 16'd3420, 16'd196, 16'd18280, 16'd37557, 16'd1912});
	test_expansion(128'hb83dfdf504becfc11c343417172f522c, {16'd45405, 16'd30880, 16'd33547, 16'd28599, 16'd55853, 16'd2298, 16'd19151, 16'd50161, 16'd29712, 16'd1076, 16'd1352, 16'd8674, 16'd31545, 16'd57008, 16'd43661, 16'd35165, 16'd54851, 16'd18322, 16'd57683, 16'd21527, 16'd18768, 16'd52881, 16'd8748, 16'd32817, 16'd48439, 16'd40358});
	test_expansion(128'h8aee973cddb2ad9a8517d480382dfc33, {16'd27841, 16'd3135, 16'd27026, 16'd56407, 16'd45566, 16'd55659, 16'd14551, 16'd55850, 16'd44589, 16'd56027, 16'd45440, 16'd9274, 16'd39617, 16'd62641, 16'd61205, 16'd64113, 16'd42346, 16'd26624, 16'd41719, 16'd37042, 16'd38005, 16'd12388, 16'd32187, 16'd44171, 16'd9806, 16'd49321});
	test_expansion(128'h65be21d214d61d50640e6b07a11e51f5, {16'd15979, 16'd36042, 16'd29690, 16'd39654, 16'd11336, 16'd61076, 16'd51505, 16'd61238, 16'd36561, 16'd49257, 16'd12208, 16'd33564, 16'd54638, 16'd44043, 16'd16618, 16'd62112, 16'd3971, 16'd14288, 16'd5514, 16'd41017, 16'd26396, 16'd35801, 16'd11926, 16'd24663, 16'd15697, 16'd44726});
	test_expansion(128'hff424f5d442b66e00b1fe4f0152f01bc, {16'd28528, 16'd41172, 16'd9292, 16'd12777, 16'd47666, 16'd42676, 16'd7706, 16'd25630, 16'd51203, 16'd20367, 16'd29282, 16'd47695, 16'd48401, 16'd33936, 16'd23883, 16'd54369, 16'd20569, 16'd20898, 16'd58492, 16'd38376, 16'd25416, 16'd37275, 16'd14724, 16'd61744, 16'd464, 16'd34986});
	test_expansion(128'h56359754a97423900102b7a75236bf78, {16'd21625, 16'd45848, 16'd49602, 16'd19595, 16'd578, 16'd25329, 16'd49050, 16'd54577, 16'd22173, 16'd31692, 16'd32481, 16'd9236, 16'd50157, 16'd34858, 16'd49307, 16'd12655, 16'd43607, 16'd63711, 16'd44491, 16'd49719, 16'd53758, 16'd11926, 16'd23492, 16'd32927, 16'd9002, 16'd42854});
	test_expansion(128'h84f2013ed331373536c629324f4b600e, {16'd33613, 16'd46300, 16'd37959, 16'd11524, 16'd14643, 16'd12429, 16'd32467, 16'd53997, 16'd42873, 16'd37631, 16'd7071, 16'd33644, 16'd11782, 16'd62537, 16'd45105, 16'd35074, 16'd20317, 16'd7861, 16'd37185, 16'd1971, 16'd42381, 16'd25251, 16'd44956, 16'd48685, 16'd2543, 16'd49722});
	test_expansion(128'hc9c166e00353920a4a9d7b973ca0c11e, {16'd13160, 16'd4465, 16'd6861, 16'd43560, 16'd61285, 16'd37579, 16'd63381, 16'd54214, 16'd10742, 16'd15166, 16'd509, 16'd62001, 16'd8138, 16'd53358, 16'd18026, 16'd42720, 16'd35543, 16'd45310, 16'd19886, 16'd21993, 16'd38285, 16'd29256, 16'd8830, 16'd64314, 16'd344, 16'd54016});
	test_expansion(128'h5084ceb1c5372ae50765fa1c12fdd908, {16'd14709, 16'd43638, 16'd5292, 16'd5435, 16'd13546, 16'd24932, 16'd1734, 16'd42404, 16'd21982, 16'd11756, 16'd10109, 16'd42049, 16'd14303, 16'd51596, 16'd35527, 16'd42130, 16'd37505, 16'd11318, 16'd21166, 16'd10132, 16'd37662, 16'd41399, 16'd15494, 16'd620, 16'd21851, 16'd40484});
	test_expansion(128'h43d098eb836af25aae9b89558e30c20b, {16'd45286, 16'd10338, 16'd1164, 16'd13825, 16'd46647, 16'd23832, 16'd53989, 16'd25932, 16'd46595, 16'd56787, 16'd20179, 16'd7906, 16'd1131, 16'd63488, 16'd55336, 16'd7476, 16'd43913, 16'd34160, 16'd38385, 16'd55523, 16'd39750, 16'd43638, 16'd39172, 16'd48769, 16'd22042, 16'd11223});
	test_expansion(128'hd039cc18a4b46f12b3627d8ae21341ef, {16'd48154, 16'd60283, 16'd63509, 16'd2385, 16'd13818, 16'd18288, 16'd24031, 16'd51913, 16'd20807, 16'd4089, 16'd56231, 16'd50479, 16'd33710, 16'd35006, 16'd24780, 16'd12974, 16'd8347, 16'd14267, 16'd11551, 16'd54931, 16'd29207, 16'd30647, 16'd5219, 16'd29410, 16'd56663, 16'd37598});
	test_expansion(128'h3c48c4aa35c45216723a5c43447f8bbd, {16'd23812, 16'd31389, 16'd42256, 16'd29374, 16'd7344, 16'd30852, 16'd59236, 16'd61352, 16'd34955, 16'd55306, 16'd46387, 16'd45089, 16'd48151, 16'd25120, 16'd42758, 16'd21213, 16'd64643, 16'd41825, 16'd18751, 16'd43860, 16'd2781, 16'd51439, 16'd53884, 16'd65162, 16'd29143, 16'd31738});
	test_expansion(128'hc16fc21c2f4aed758b46ce7aba730dd9, {16'd59131, 16'd25643, 16'd24315, 16'd41275, 16'd6486, 16'd41066, 16'd7932, 16'd21201, 16'd17905, 16'd44379, 16'd20336, 16'd29695, 16'd54784, 16'd49045, 16'd37643, 16'd34928, 16'd19310, 16'd61355, 16'd60543, 16'd18869, 16'd23911, 16'd36456, 16'd22471, 16'd29655, 16'd52436, 16'd20050});
	test_expansion(128'he6bf3cf9843d59f4ea191cab7e9fbc61, {16'd10009, 16'd3719, 16'd28123, 16'd26084, 16'd62023, 16'd9834, 16'd51850, 16'd7650, 16'd52713, 16'd1707, 16'd57679, 16'd45164, 16'd2365, 16'd12341, 16'd39406, 16'd7616, 16'd21081, 16'd44721, 16'd29755, 16'd56520, 16'd11527, 16'd49626, 16'd48333, 16'd48691, 16'd6707, 16'd17604});
	test_expansion(128'h1a21ab5a457cdfdb0edf28d72a83fdfb, {16'd47273, 16'd49569, 16'd60110, 16'd39136, 16'd23550, 16'd38456, 16'd53141, 16'd21127, 16'd27583, 16'd24464, 16'd7125, 16'd1488, 16'd61626, 16'd11303, 16'd62931, 16'd59054, 16'd31100, 16'd65483, 16'd7214, 16'd36079, 16'd61967, 16'd52435, 16'd26922, 16'd65239, 16'd42481, 16'd19843});
	test_expansion(128'h346950c8c53abf79569272e6a8902a85, {16'd29040, 16'd23035, 16'd57664, 16'd48965, 16'd26186, 16'd43534, 16'd46599, 16'd7533, 16'd29592, 16'd15664, 16'd32185, 16'd37872, 16'd23583, 16'd18200, 16'd33595, 16'd64127, 16'd404, 16'd1953, 16'd44716, 16'd38929, 16'd49608, 16'd61352, 16'd64965, 16'd28168, 16'd54924, 16'd15879});
	test_expansion(128'hb76ebedc7fb5bc44dd1727dbb3ed77df, {16'd21045, 16'd33389, 16'd18423, 16'd23854, 16'd47853, 16'd2703, 16'd1688, 16'd34417, 16'd30894, 16'd22016, 16'd16663, 16'd44089, 16'd21249, 16'd42500, 16'd8106, 16'd46705, 16'd39647, 16'd5165, 16'd14077, 16'd36402, 16'd55435, 16'd7974, 16'd30417, 16'd8238, 16'd35677, 16'd44618});
	test_expansion(128'hb67ce888d2bc2537c878420b2be7eeaa, {16'd7344, 16'd36136, 16'd29289, 16'd26515, 16'd37709, 16'd44002, 16'd40878, 16'd34321, 16'd1603, 16'd36030, 16'd60857, 16'd21465, 16'd12850, 16'd15061, 16'd56199, 16'd27347, 16'd50814, 16'd42973, 16'd3549, 16'd38306, 16'd9689, 16'd14735, 16'd42123, 16'd39471, 16'd8829, 16'd45699});
	test_expansion(128'h9c73222ba222b6932a896ee27ae7d7cc, {16'd18767, 16'd62228, 16'd51184, 16'd2886, 16'd34889, 16'd55966, 16'd37480, 16'd23060, 16'd26203, 16'd16322, 16'd7431, 16'd7289, 16'd39492, 16'd53612, 16'd13231, 16'd59035, 16'd34798, 16'd1358, 16'd7992, 16'd45846, 16'd57892, 16'd4841, 16'd32768, 16'd58859, 16'd37746, 16'd44185});
	test_expansion(128'h7e2cc13c3cfe62cfd0d75b9bd598e9e8, {16'd56837, 16'd63876, 16'd61501, 16'd13518, 16'd21033, 16'd52515, 16'd7436, 16'd47975, 16'd5630, 16'd48788, 16'd55538, 16'd48651, 16'd38735, 16'd57089, 16'd10830, 16'd38377, 16'd3412, 16'd45921, 16'd12505, 16'd9440, 16'd19864, 16'd878, 16'd27882, 16'd1673, 16'd54714, 16'd16532});
	test_expansion(128'h2c2210e71de043c5173f8770fe05ebe4, {16'd57446, 16'd12731, 16'd59613, 16'd18326, 16'd36446, 16'd63965, 16'd33480, 16'd35404, 16'd36533, 16'd54929, 16'd38757, 16'd41695, 16'd55432, 16'd24004, 16'd59909, 16'd11517, 16'd31346, 16'd48447, 16'd33571, 16'd34639, 16'd65415, 16'd36668, 16'd23504, 16'd50687, 16'd52972, 16'd61074});
	test_expansion(128'hf3b63dd3214666f7bd582f39798e2312, {16'd956, 16'd4795, 16'd24448, 16'd28396, 16'd27724, 16'd62120, 16'd32743, 16'd8721, 16'd54558, 16'd13285, 16'd57004, 16'd27806, 16'd63792, 16'd32512, 16'd26265, 16'd64925, 16'd12934, 16'd30162, 16'd31684, 16'd28456, 16'd58160, 16'd5955, 16'd19752, 16'd37434, 16'd59794, 16'd48591});
	test_expansion(128'hf0bd7079832ebc79dfbb8137897a31f8, {16'd35087, 16'd38482, 16'd39715, 16'd17879, 16'd9084, 16'd11861, 16'd5114, 16'd15701, 16'd45280, 16'd15022, 16'd39396, 16'd37557, 16'd19399, 16'd47233, 16'd19799, 16'd13045, 16'd11320, 16'd21552, 16'd33124, 16'd36447, 16'd17313, 16'd20572, 16'd23920, 16'd27491, 16'd31054, 16'd61522});
	test_expansion(128'hda49b6522743098dc0b4d6cbda2b278f, {16'd48174, 16'd31415, 16'd49097, 16'd21676, 16'd28742, 16'd10396, 16'd43718, 16'd22823, 16'd15816, 16'd61195, 16'd52780, 16'd29411, 16'd7934, 16'd55900, 16'd19347, 16'd59792, 16'd19173, 16'd56410, 16'd60241, 16'd29763, 16'd41571, 16'd25159, 16'd31498, 16'd37418, 16'd1063, 16'd47682});
	test_expansion(128'hcdbe71ce0e80b50ebc252ab1bdcd4821, {16'd56947, 16'd23016, 16'd33273, 16'd30034, 16'd57293, 16'd63650, 16'd52761, 16'd19087, 16'd30429, 16'd45775, 16'd11087, 16'd28432, 16'd47963, 16'd5234, 16'd27010, 16'd20529, 16'd52612, 16'd21037, 16'd64345, 16'd41369, 16'd56984, 16'd58574, 16'd59061, 16'd34802, 16'd42006, 16'd31521});
	test_expansion(128'h073ce1849a163a9b93a0dba20557ae71, {16'd40910, 16'd22307, 16'd7146, 16'd65067, 16'd56116, 16'd51302, 16'd17478, 16'd47261, 16'd60069, 16'd33381, 16'd51618, 16'd16614, 16'd36353, 16'd31229, 16'd47073, 16'd35570, 16'd61777, 16'd55599, 16'd19979, 16'd19076, 16'd33270, 16'd54024, 16'd14232, 16'd46640, 16'd24336, 16'd13615});
	test_expansion(128'hd06bb7f1df57f9acceac87b5dc398a81, {16'd7145, 16'd60998, 16'd56812, 16'd52070, 16'd46486, 16'd56097, 16'd62380, 16'd62318, 16'd34100, 16'd30903, 16'd63671, 16'd24504, 16'd57920, 16'd58935, 16'd7783, 16'd46906, 16'd288, 16'd7015, 16'd44440, 16'd45066, 16'd44730, 16'd41279, 16'd47077, 16'd1121, 16'd58902, 16'd21397});
	test_expansion(128'hbd34fb85892a6872eb8cda3a18a1d941, {16'd31103, 16'd52058, 16'd65470, 16'd4815, 16'd28853, 16'd64699, 16'd33413, 16'd54634, 16'd48457, 16'd32893, 16'd363, 16'd25904, 16'd34080, 16'd42561, 16'd16543, 16'd33945, 16'd34877, 16'd31324, 16'd29311, 16'd29817, 16'd1588, 16'd48762, 16'd16677, 16'd44260, 16'd29317, 16'd8627});
	test_expansion(128'hdd4745e117ebe88f561b16e6d3b14dcd, {16'd24091, 16'd24806, 16'd10765, 16'd2177, 16'd17721, 16'd52834, 16'd35267, 16'd51340, 16'd1866, 16'd52919, 16'd55473, 16'd62135, 16'd7516, 16'd46738, 16'd33524, 16'd50882, 16'd56692, 16'd55903, 16'd2965, 16'd15399, 16'd38583, 16'd32754, 16'd365, 16'd62430, 16'd9491, 16'd61743});
	test_expansion(128'h49f05db258a39add2cfc201a9e642110, {16'd57416, 16'd60577, 16'd60399, 16'd60760, 16'd8153, 16'd44392, 16'd14219, 16'd37097, 16'd3520, 16'd20833, 16'd56933, 16'd27466, 16'd47674, 16'd51609, 16'd55337, 16'd40964, 16'd36812, 16'd18910, 16'd59649, 16'd51598, 16'd32423, 16'd4914, 16'd685, 16'd55869, 16'd51102, 16'd4251});
	test_expansion(128'h2797d7135e8b44b5ae9f93c25fa5616a, {16'd10397, 16'd27870, 16'd17754, 16'd61183, 16'd16849, 16'd22119, 16'd37287, 16'd33756, 16'd10732, 16'd7048, 16'd1421, 16'd53124, 16'd39923, 16'd3911, 16'd51322, 16'd28014, 16'd9394, 16'd20573, 16'd61241, 16'd47282, 16'd39023, 16'd24903, 16'd32908, 16'd40258, 16'd18779, 16'd15836});
	test_expansion(128'h0bdbe119d45ae54779693ef20bea0122, {16'd26539, 16'd59581, 16'd29129, 16'd44798, 16'd640, 16'd6673, 16'd47074, 16'd22803, 16'd10804, 16'd44236, 16'd58214, 16'd9543, 16'd33119, 16'd45704, 16'd31928, 16'd18752, 16'd16139, 16'd57353, 16'd15892, 16'd47079, 16'd63490, 16'd7853, 16'd8636, 16'd38529, 16'd52937, 16'd38267});
	test_expansion(128'h681a0af715ac6503287d563d01b3b9eb, {16'd40909, 16'd38074, 16'd48774, 16'd50165, 16'd30849, 16'd19833, 16'd4824, 16'd28615, 16'd34881, 16'd20242, 16'd63716, 16'd63018, 16'd57601, 16'd24654, 16'd29461, 16'd12491, 16'd2168, 16'd46547, 16'd46988, 16'd54942, 16'd6739, 16'd18184, 16'd5186, 16'd46700, 16'd40945, 16'd47180});
	test_expansion(128'hbda8cade70c94ab96311bd9b4fdb6f89, {16'd6918, 16'd13829, 16'd26495, 16'd16752, 16'd62812, 16'd36012, 16'd46345, 16'd25303, 16'd5282, 16'd44289, 16'd26569, 16'd63597, 16'd58391, 16'd27681, 16'd20052, 16'd26172, 16'd47805, 16'd50950, 16'd52670, 16'd36581, 16'd51892, 16'd54891, 16'd39938, 16'd36392, 16'd53318, 16'd51478});
	test_expansion(128'h997eb1af174a42b2a52c0a29babcefa6, {16'd26125, 16'd17083, 16'd6306, 16'd24437, 16'd54404, 16'd2328, 16'd63465, 16'd31943, 16'd38403, 16'd24493, 16'd2436, 16'd11064, 16'd65086, 16'd15247, 16'd7513, 16'd42769, 16'd16916, 16'd19487, 16'd14479, 16'd4964, 16'd30939, 16'd5490, 16'd37968, 16'd43640, 16'd38639, 16'd15387});
	test_expansion(128'hb9cdebc2cde11ab6b510a3c7527565aa, {16'd29460, 16'd63637, 16'd28656, 16'd60412, 16'd42034, 16'd37257, 16'd22046, 16'd58533, 16'd3703, 16'd8995, 16'd46635, 16'd27006, 16'd7479, 16'd44515, 16'd52280, 16'd17390, 16'd43043, 16'd18685, 16'd13093, 16'd32930, 16'd39440, 16'd27158, 16'd57813, 16'd62368, 16'd37830, 16'd64475});
	test_expansion(128'h03303c6cf4a4e5bd80029e0dfdf7f035, {16'd9013, 16'd27222, 16'd64028, 16'd42700, 16'd48643, 16'd41407, 16'd22667, 16'd36441, 16'd60780, 16'd19358, 16'd8082, 16'd52098, 16'd8524, 16'd39039, 16'd2697, 16'd61902, 16'd35029, 16'd27324, 16'd9624, 16'd22490, 16'd20154, 16'd37292, 16'd57366, 16'd60254, 16'd7763, 16'd34821});
	test_expansion(128'h76521ae215409bdb564e868dc39865e6, {16'd44579, 16'd157, 16'd9760, 16'd39541, 16'd54342, 16'd57339, 16'd1479, 16'd8245, 16'd47963, 16'd7560, 16'd19443, 16'd30883, 16'd55348, 16'd8091, 16'd64402, 16'd59945, 16'd59018, 16'd28896, 16'd39495, 16'd40141, 16'd57513, 16'd10669, 16'd41457, 16'd37327, 16'd25308, 16'd41147});
	test_expansion(128'hec8db12fd30e37e2a63fdabcc6295fac, {16'd63532, 16'd12224, 16'd10981, 16'd59645, 16'd52644, 16'd42859, 16'd6138, 16'd3507, 16'd60104, 16'd21401, 16'd52046, 16'd52257, 16'd46105, 16'd17166, 16'd53630, 16'd35536, 16'd18529, 16'd33727, 16'd41436, 16'd5892, 16'd36263, 16'd13691, 16'd7332, 16'd57946, 16'd17307, 16'd32894});
	test_expansion(128'hd0631ff8662a318fb737281b94963f87, {16'd3638, 16'd25515, 16'd28200, 16'd25090, 16'd50312, 16'd8353, 16'd13365, 16'd27301, 16'd15879, 16'd22303, 16'd43620, 16'd53016, 16'd45087, 16'd41674, 16'd59634, 16'd1090, 16'd51569, 16'd39871, 16'd43763, 16'd50325, 16'd15101, 16'd63721, 16'd60726, 16'd36721, 16'd16761, 16'd23262});
	test_expansion(128'h3cf862d4383f255b85bfe451621bfa58, {16'd23975, 16'd35301, 16'd64535, 16'd7999, 16'd37542, 16'd57562, 16'd28977, 16'd29832, 16'd27801, 16'd49814, 16'd54469, 16'd4558, 16'd4605, 16'd60173, 16'd24378, 16'd19082, 16'd54474, 16'd42524, 16'd27211, 16'd10845, 16'd34191, 16'd56297, 16'd31895, 16'd8419, 16'd53624, 16'd36118});
	test_expansion(128'hdfc7e9228b041d0048cb86b622b7d017, {16'd63340, 16'd63932, 16'd1539, 16'd36849, 16'd19090, 16'd57263, 16'd24115, 16'd39866, 16'd30162, 16'd11576, 16'd45521, 16'd28871, 16'd61668, 16'd13745, 16'd28083, 16'd65045, 16'd64056, 16'd35273, 16'd33630, 16'd11182, 16'd45784, 16'd47614, 16'd51042, 16'd61607, 16'd63504, 16'd48671});
	test_expansion(128'h44978263f91687ea20636d6f06d0477d, {16'd41703, 16'd15467, 16'd32392, 16'd37942, 16'd31740, 16'd17332, 16'd60911, 16'd40975, 16'd55912, 16'd50079, 16'd12569, 16'd53015, 16'd27759, 16'd35869, 16'd42834, 16'd17949, 16'd59118, 16'd41459, 16'd39335, 16'd21686, 16'd41600, 16'd7938, 16'd58457, 16'd9744, 16'd19639, 16'd27495});
	test_expansion(128'hc54a12213ce827e0de5491117dc38c10, {16'd57576, 16'd32365, 16'd37560, 16'd34063, 16'd34108, 16'd14635, 16'd56017, 16'd60832, 16'd64580, 16'd53490, 16'd41306, 16'd49201, 16'd43789, 16'd50808, 16'd1779, 16'd22665, 16'd4295, 16'd39457, 16'd9618, 16'd40495, 16'd17740, 16'd1627, 16'd53698, 16'd26087, 16'd21159, 16'd59455});
	test_expansion(128'hc8beb8300ea1612a06cd9a7f3369bb7b, {16'd55116, 16'd30341, 16'd11703, 16'd4569, 16'd8645, 16'd21029, 16'd50338, 16'd5689, 16'd12921, 16'd53191, 16'd27002, 16'd46683, 16'd15263, 16'd45962, 16'd27963, 16'd19808, 16'd48771, 16'd7071, 16'd60232, 16'd24612, 16'd21434, 16'd23744, 16'd63305, 16'd10566, 16'd13360, 16'd56723});
	test_expansion(128'h02b1756c9a953bcf432e0bf5839beb6c, {16'd39266, 16'd25402, 16'd24144, 16'd17542, 16'd39117, 16'd20872, 16'd62447, 16'd44858, 16'd19273, 16'd12352, 16'd12972, 16'd60929, 16'd34358, 16'd42223, 16'd49289, 16'd49178, 16'd39577, 16'd32415, 16'd64255, 16'd13213, 16'd35762, 16'd56433, 16'd17455, 16'd10996, 16'd11386, 16'd26587});
	test_expansion(128'hbe164cf9d3ca72b4a375ced7e308932f, {16'd3487, 16'd62029, 16'd57986, 16'd53563, 16'd1780, 16'd9555, 16'd18034, 16'd38472, 16'd38549, 16'd40732, 16'd58350, 16'd19554, 16'd32909, 16'd37431, 16'd49339, 16'd9472, 16'd12017, 16'd11671, 16'd6777, 16'd43886, 16'd46589, 16'd52158, 16'd34697, 16'd1651, 16'd11823, 16'd51168});
	test_expansion(128'h628febef830541c1fdc1fa9957cd9019, {16'd21692, 16'd45628, 16'd35113, 16'd31708, 16'd17134, 16'd16056, 16'd53762, 16'd32226, 16'd57185, 16'd42497, 16'd36967, 16'd64385, 16'd30382, 16'd57068, 16'd50546, 16'd62102, 16'd43138, 16'd58448, 16'd53463, 16'd10878, 16'd13317, 16'd7213, 16'd55602, 16'd30705, 16'd47347, 16'd42806});
	test_expansion(128'h7c380f86a6edcdf06c69c616d79f5f29, {16'd12264, 16'd25149, 16'd22213, 16'd22399, 16'd62373, 16'd47086, 16'd894, 16'd44281, 16'd61466, 16'd1240, 16'd24943, 16'd44253, 16'd18238, 16'd40489, 16'd52876, 16'd30837, 16'd37053, 16'd57507, 16'd9491, 16'd4993, 16'd2649, 16'd36439, 16'd38082, 16'd24604, 16'd12774, 16'd2446});
	test_expansion(128'hda1b497984d8c331f6f9866107beb863, {16'd38321, 16'd52963, 16'd48207, 16'd17326, 16'd48294, 16'd10883, 16'd8260, 16'd62160, 16'd22714, 16'd21700, 16'd43296, 16'd48200, 16'd30162, 16'd33065, 16'd19300, 16'd15440, 16'd55565, 16'd40342, 16'd5330, 16'd28992, 16'd47089, 16'd51982, 16'd21917, 16'd63099, 16'd23071, 16'd51705});
	test_expansion(128'hcb6fb71ede445255a719d3251961c91a, {16'd45586, 16'd6673, 16'd31825, 16'd33768, 16'd9603, 16'd5127, 16'd26343, 16'd38717, 16'd44320, 16'd24741, 16'd1931, 16'd9283, 16'd55748, 16'd3654, 16'd54345, 16'd34037, 16'd23765, 16'd55984, 16'd44743, 16'd40901, 16'd34277, 16'd7070, 16'd40494, 16'd19341, 16'd9436, 16'd64987});
	test_expansion(128'h3173546897c5d5e09c1eb30089caf7cc, {16'd27162, 16'd44307, 16'd40929, 16'd25203, 16'd61225, 16'd6847, 16'd9520, 16'd29394, 16'd31142, 16'd43900, 16'd43553, 16'd59386, 16'd3262, 16'd36544, 16'd50274, 16'd4929, 16'd45814, 16'd61885, 16'd46829, 16'd10754, 16'd16916, 16'd57712, 16'd12711, 16'd36397, 16'd3798, 16'd61302});
	test_expansion(128'hba8998afee46405a241a2e25589fb075, {16'd6720, 16'd16392, 16'd224, 16'd39542, 16'd2402, 16'd5754, 16'd2262, 16'd13821, 16'd25706, 16'd23456, 16'd39834, 16'd20522, 16'd5903, 16'd35559, 16'd585, 16'd32277, 16'd39884, 16'd21603, 16'd14269, 16'd50815, 16'd7640, 16'd65304, 16'd57885, 16'd25525, 16'd57404, 16'd36517});
	test_expansion(128'hdc0349cb2b64a07f6257b2a0513c7b74, {16'd5242, 16'd62674, 16'd49221, 16'd35113, 16'd11494, 16'd20244, 16'd26935, 16'd56168, 16'd63391, 16'd8570, 16'd28648, 16'd5629, 16'd48564, 16'd45780, 16'd31408, 16'd53174, 16'd63488, 16'd38558, 16'd40484, 16'd3372, 16'd48965, 16'd22793, 16'd22358, 16'd8486, 16'd59085, 16'd40853});
	test_expansion(128'h4eab269aa3863c911217c0b54a9765b7, {16'd64196, 16'd55202, 16'd28664, 16'd48456, 16'd64832, 16'd40487, 16'd18453, 16'd18642, 16'd52055, 16'd8151, 16'd59376, 16'd36946, 16'd53549, 16'd9623, 16'd23633, 16'd45222, 16'd44254, 16'd58918, 16'd22347, 16'd47175, 16'd24432, 16'd27664, 16'd44736, 16'd27919, 16'd11742, 16'd37044});
	test_expansion(128'h5bb4332b7ab344a43dedfbf2dbb6b628, {16'd10898, 16'd42355, 16'd41354, 16'd48556, 16'd53562, 16'd32640, 16'd27044, 16'd34985, 16'd64721, 16'd32617, 16'd12961, 16'd46795, 16'd48645, 16'd41806, 16'd36759, 16'd53828, 16'd23876, 16'd27686, 16'd60404, 16'd6141, 16'd60192, 16'd51503, 16'd49857, 16'd25983, 16'd28931, 16'd9958});
	test_expansion(128'h22e3f7bfdd027c484bce92227ca67904, {16'd46372, 16'd40331, 16'd26428, 16'd59511, 16'd7812, 16'd53387, 16'd53173, 16'd14105, 16'd56606, 16'd4367, 16'd10769, 16'd12773, 16'd24368, 16'd34616, 16'd12791, 16'd20619, 16'd15715, 16'd14288, 16'd62107, 16'd14215, 16'd17041, 16'd62897, 16'd6702, 16'd41272, 16'd30000, 16'd53584});
	test_expansion(128'h8331322ace7dc1cd9f377b94f195f663, {16'd63457, 16'd22059, 16'd29473, 16'd45333, 16'd64338, 16'd36457, 16'd59312, 16'd63263, 16'd48032, 16'd6953, 16'd52828, 16'd45241, 16'd25674, 16'd29717, 16'd65177, 16'd214, 16'd61211, 16'd43896, 16'd12812, 16'd16033, 16'd38136, 16'd22556, 16'd4045, 16'd39369, 16'd33303, 16'd45819});
	test_expansion(128'h0f4f55ac5c0606834dae7807df77966e, {16'd43527, 16'd30457, 16'd4329, 16'd64659, 16'd28472, 16'd43367, 16'd15346, 16'd5623, 16'd38286, 16'd3519, 16'd41061, 16'd19201, 16'd45945, 16'd35847, 16'd54787, 16'd42084, 16'd23105, 16'd18896, 16'd59839, 16'd31145, 16'd37510, 16'd40753, 16'd54219, 16'd53104, 16'd49631, 16'd27053});
	test_expansion(128'hec30e4aaf9de9458c65ce02122c0fe0b, {16'd25220, 16'd14325, 16'd35630, 16'd63354, 16'd52969, 16'd34240, 16'd12453, 16'd61432, 16'd43037, 16'd34850, 16'd14693, 16'd54041, 16'd54596, 16'd56499, 16'd8277, 16'd27914, 16'd14304, 16'd42581, 16'd4550, 16'd11577, 16'd39638, 16'd27241, 16'd14261, 16'd25749, 16'd56400, 16'd31396});
	test_expansion(128'hbb99815f51981d2bff286746d4da643b, {16'd25577, 16'd58865, 16'd15077, 16'd6025, 16'd55594, 16'd65173, 16'd20000, 16'd28809, 16'd59236, 16'd27872, 16'd44702, 16'd20068, 16'd49343, 16'd36035, 16'd22441, 16'd19540, 16'd4462, 16'd58445, 16'd39906, 16'd44417, 16'd12342, 16'd55675, 16'd60288, 16'd3687, 16'd51110, 16'd34044});
	test_expansion(128'h7e8ea340fe2a34b7612115c325696090, {16'd31983, 16'd48541, 16'd36538, 16'd56384, 16'd63914, 16'd36401, 16'd23866, 16'd8621, 16'd11423, 16'd59545, 16'd58329, 16'd36139, 16'd58281, 16'd33598, 16'd46248, 16'd53943, 16'd21977, 16'd28410, 16'd25248, 16'd48369, 16'd62039, 16'd2258, 16'd30318, 16'd52541, 16'd60771, 16'd36114});
	test_expansion(128'h251669a819e8f2bc245d170575672dc0, {16'd59896, 16'd6986, 16'd63779, 16'd46533, 16'd2058, 16'd1984, 16'd57180, 16'd45623, 16'd10564, 16'd21222, 16'd33845, 16'd58793, 16'd61817, 16'd1916, 16'd19899, 16'd27028, 16'd18814, 16'd36535, 16'd53002, 16'd58139, 16'd26530, 16'd28887, 16'd54105, 16'd59436, 16'd49151, 16'd611});
	test_expansion(128'h6887ca8db65793f1fb7e7fba77e0c9a8, {16'd24005, 16'd46800, 16'd1703, 16'd2421, 16'd39166, 16'd25674, 16'd56853, 16'd7218, 16'd53061, 16'd49996, 16'd18689, 16'd27999, 16'd25290, 16'd12391, 16'd58555, 16'd41064, 16'd58254, 16'd56342, 16'd46212, 16'd18904, 16'd47325, 16'd19787, 16'd59274, 16'd27799, 16'd7605, 16'd27040});
	test_expansion(128'h25e2906440289d66517b5efed251cf3f, {16'd44287, 16'd19520, 16'd36733, 16'd54268, 16'd25721, 16'd18090, 16'd64918, 16'd46634, 16'd36032, 16'd17136, 16'd64928, 16'd45105, 16'd37577, 16'd7747, 16'd45708, 16'd15109, 16'd35629, 16'd45776, 16'd45874, 16'd44411, 16'd44309, 16'd23062, 16'd44308, 16'd53984, 16'd348, 16'd26687});
	test_expansion(128'h73465017ef4bec8d4ffd71d684481004, {16'd56501, 16'd31220, 16'd7843, 16'd23152, 16'd40675, 16'd28366, 16'd29282, 16'd58885, 16'd57847, 16'd18469, 16'd41076, 16'd3423, 16'd45830, 16'd54150, 16'd40576, 16'd13460, 16'd20642, 16'd30591, 16'd557, 16'd12456, 16'd42714, 16'd25876, 16'd27210, 16'd41282, 16'd8076, 16'd44246});
	test_expansion(128'h74dd76fccd48c98ac7fc36441ff34ba3, {16'd59349, 16'd53520, 16'd28817, 16'd20028, 16'd11244, 16'd36293, 16'd59772, 16'd11438, 16'd64185, 16'd2230, 16'd6826, 16'd7042, 16'd42082, 16'd23157, 16'd39166, 16'd56203, 16'd45985, 16'd47285, 16'd15969, 16'd16800, 16'd22889, 16'd5462, 16'd26239, 16'd5292, 16'd28406, 16'd54986});
	test_expansion(128'he3f76fe221bf1f1b57bb1afa6b632459, {16'd50634, 16'd39308, 16'd33121, 16'd64058, 16'd64469, 16'd13755, 16'd36952, 16'd47943, 16'd38354, 16'd38567, 16'd17638, 16'd55502, 16'd30343, 16'd64482, 16'd33111, 16'd18547, 16'd37962, 16'd32486, 16'd33533, 16'd28848, 16'd941, 16'd19169, 16'd56815, 16'd64254, 16'd27600, 16'd6035});
	test_expansion(128'h98d74529bf1c980961208535df68b76f, {16'd36779, 16'd9211, 16'd56988, 16'd42907, 16'd60771, 16'd10229, 16'd58420, 16'd27986, 16'd48726, 16'd52076, 16'd9081, 16'd29163, 16'd46727, 16'd50852, 16'd838, 16'd61900, 16'd22961, 16'd29388, 16'd54282, 16'd62090, 16'd53775, 16'd63632, 16'd22247, 16'd50833, 16'd63561, 16'd32972});
	test_expansion(128'hc16d4099c87475f100b5d0e1b59eb656, {16'd14771, 16'd28834, 16'd40820, 16'd27059, 16'd21789, 16'd55603, 16'd45951, 16'd22482, 16'd5653, 16'd12513, 16'd54216, 16'd15244, 16'd40023, 16'd34608, 16'd14685, 16'd14923, 16'd39481, 16'd64855, 16'd16058, 16'd4656, 16'd18065, 16'd27677, 16'd58042, 16'd32770, 16'd20611, 16'd16921});
	test_expansion(128'h414c5d306825e7e7a32af84a42d5475b, {16'd19138, 16'd12918, 16'd33347, 16'd35311, 16'd17490, 16'd35728, 16'd39862, 16'd12300, 16'd54818, 16'd22908, 16'd18100, 16'd16551, 16'd12260, 16'd64118, 16'd48074, 16'd14074, 16'd26313, 16'd20193, 16'd50168, 16'd42139, 16'd59683, 16'd23280, 16'd32773, 16'd51477, 16'd37243, 16'd18286});
	test_expansion(128'h0636248af75a92d7c7bdfb171ef6c9ce, {16'd26549, 16'd14152, 16'd47373, 16'd6061, 16'd49833, 16'd34082, 16'd14414, 16'd47994, 16'd59656, 16'd30519, 16'd47335, 16'd41592, 16'd31495, 16'd38063, 16'd35741, 16'd48675, 16'd58014, 16'd36367, 16'd32141, 16'd57353, 16'd34164, 16'd42659, 16'd13856, 16'd2296, 16'd38751, 16'd28748});
	test_expansion(128'he2d345b1714e96352c1846e3c1416adb, {16'd44897, 16'd55204, 16'd12913, 16'd62601, 16'd8424, 16'd44084, 16'd58553, 16'd34947, 16'd42260, 16'd5472, 16'd46831, 16'd3936, 16'd40340, 16'd25178, 16'd3211, 16'd3752, 16'd47581, 16'd21719, 16'd2412, 16'd59146, 16'd52170, 16'd34775, 16'd57869, 16'd13668, 16'd21302, 16'd42729});
	test_expansion(128'h600af497a958f72ae82f965bca8ae927, {16'd48441, 16'd59141, 16'd59459, 16'd49134, 16'd33188, 16'd30032, 16'd21043, 16'd8035, 16'd31273, 16'd63513, 16'd57453, 16'd3350, 16'd13368, 16'd44442, 16'd53406, 16'd16699, 16'd22066, 16'd5715, 16'd29148, 16'd35758, 16'd17812, 16'd10277, 16'd7605, 16'd42846, 16'd19159, 16'd5141});
	test_expansion(128'h6f0ce19ca3d4219ce86b9f1b66e2d585, {16'd51988, 16'd35876, 16'd31473, 16'd21208, 16'd23785, 16'd38360, 16'd16373, 16'd31538, 16'd9881, 16'd27817, 16'd34243, 16'd14313, 16'd38986, 16'd28381, 16'd12717, 16'd53744, 16'd4392, 16'd6772, 16'd34595, 16'd2937, 16'd11647, 16'd58486, 16'd60355, 16'd14993, 16'd57310, 16'd39217});
	test_expansion(128'ha90fedc6405c61010c873db59802a550, {16'd41345, 16'd19233, 16'd34281, 16'd55331, 16'd52899, 16'd48470, 16'd50774, 16'd59529, 16'd43898, 16'd61192, 16'd30726, 16'd61221, 16'd58489, 16'd37810, 16'd29022, 16'd45838, 16'd65357, 16'd20033, 16'd63517, 16'd30851, 16'd53805, 16'd40811, 16'd37840, 16'd30046, 16'd1879, 16'd12323});
	test_expansion(128'h3e54ced177fc14f5f5ed47ef00241fbf, {16'd44112, 16'd48634, 16'd7255, 16'd31325, 16'd53561, 16'd55394, 16'd26968, 16'd53251, 16'd2908, 16'd49408, 16'd53785, 16'd25770, 16'd51781, 16'd49837, 16'd12736, 16'd61190, 16'd22229, 16'd38342, 16'd60556, 16'd60055, 16'd42614, 16'd46379, 16'd33414, 16'd29802, 16'd30220, 16'd23629});
	test_expansion(128'h8b565bb162f2970310f671dd43a1cc5a, {16'd32243, 16'd30357, 16'd54329, 16'd42877, 16'd31409, 16'd51113, 16'd57843, 16'd55173, 16'd4015, 16'd57057, 16'd36501, 16'd44827, 16'd13644, 16'd64586, 16'd46275, 16'd7371, 16'd18569, 16'd61056, 16'd51619, 16'd9977, 16'd49937, 16'd30317, 16'd26439, 16'd17830, 16'd17154, 16'd1118});
	test_expansion(128'h9919d3f4970bf198974d90c1517c8316, {16'd50761, 16'd28037, 16'd33679, 16'd3793, 16'd20259, 16'd35405, 16'd18027, 16'd2520, 16'd30718, 16'd41683, 16'd24243, 16'd21455, 16'd1191, 16'd45625, 16'd4236, 16'd12412, 16'd7592, 16'd65017, 16'd32970, 16'd37615, 16'd41425, 16'd19594, 16'd58869, 16'd48492, 16'd6152, 16'd11033});
	test_expansion(128'h9fcb646495b0d8e9b3d44b4b38ecc80e, {16'd62303, 16'd12491, 16'd32209, 16'd4971, 16'd23555, 16'd30438, 16'd51162, 16'd37425, 16'd19805, 16'd7932, 16'd19969, 16'd62824, 16'd55351, 16'd3421, 16'd26720, 16'd52049, 16'd63509, 16'd35279, 16'd55308, 16'd46103, 16'd58514, 16'd5676, 16'd13865, 16'd24378, 16'd35192, 16'd54806});
	test_expansion(128'h73b8384bcfdfa295fb80a615e0d650c5, {16'd2571, 16'd1722, 16'd60256, 16'd8263, 16'd8629, 16'd41067, 16'd46156, 16'd56868, 16'd33546, 16'd8792, 16'd58988, 16'd55601, 16'd40122, 16'd13775, 16'd58099, 16'd25138, 16'd56487, 16'd53888, 16'd12708, 16'd54830, 16'd6690, 16'd35616, 16'd16469, 16'd41451, 16'd61439, 16'd55263});
	test_expansion(128'h97e852500edae737521daa79e58abcda, {16'd40773, 16'd63175, 16'd397, 16'd58255, 16'd24995, 16'd1975, 16'd51088, 16'd24700, 16'd19564, 16'd25021, 16'd12311, 16'd63238, 16'd22765, 16'd26716, 16'd49290, 16'd46297, 16'd12223, 16'd36183, 16'd32439, 16'd62996, 16'd56526, 16'd46615, 16'd23940, 16'd7732, 16'd8202, 16'd34162});
	test_expansion(128'h21ace3032c655b06276f23470358cbe4, {16'd4699, 16'd39480, 16'd17995, 16'd53717, 16'd917, 16'd47144, 16'd30720, 16'd17453, 16'd25592, 16'd49288, 16'd36632, 16'd23066, 16'd34731, 16'd28958, 16'd40424, 16'd59985, 16'd14345, 16'd62773, 16'd15519, 16'd40351, 16'd12700, 16'd43731, 16'd2980, 16'd37494, 16'd8562, 16'd39003});
	test_expansion(128'h0cac5ab00d50172acfab4bda3a5bea0b, {16'd30427, 16'd36243, 16'd47120, 16'd9710, 16'd43172, 16'd7039, 16'd19788, 16'd26696, 16'd24343, 16'd12986, 16'd37168, 16'd33071, 16'd59966, 16'd19036, 16'd29227, 16'd63217, 16'd46753, 16'd46669, 16'd12000, 16'd2784, 16'd22865, 16'd18604, 16'd57520, 16'd44769, 16'd55365, 16'd20102});
	test_expansion(128'hfa3a6cfcfef9b6188af01e4246280881, {16'd25024, 16'd61462, 16'd33986, 16'd32549, 16'd35236, 16'd36596, 16'd15120, 16'd49677, 16'd1522, 16'd32354, 16'd29741, 16'd26263, 16'd41732, 16'd36718, 16'd47616, 16'd19367, 16'd58397, 16'd18573, 16'd6820, 16'd14427, 16'd2080, 16'd5554, 16'd45906, 16'd26437, 16'd62868, 16'd15689});
	test_expansion(128'hf628a9fe4db554318707759a9c24548f, {16'd43875, 16'd2022, 16'd42910, 16'd19756, 16'd15783, 16'd53393, 16'd19637, 16'd57282, 16'd5268, 16'd17400, 16'd57860, 16'd26407, 16'd8269, 16'd9680, 16'd43213, 16'd611, 16'd31414, 16'd56186, 16'd51321, 16'd61971, 16'd34732, 16'd7556, 16'd62128, 16'd63767, 16'd4936, 16'd31101});
	test_expansion(128'hbe46794bf4c2ec744b5960b61db739e8, {16'd29236, 16'd31998, 16'd30706, 16'd7055, 16'd11002, 16'd30601, 16'd47741, 16'd8493, 16'd47635, 16'd16270, 16'd40937, 16'd6217, 16'd62698, 16'd153, 16'd15830, 16'd9094, 16'd34603, 16'd60513, 16'd49580, 16'd15311, 16'd57565, 16'd57276, 16'd14988, 16'd13382, 16'd21175, 16'd44296});
	test_expansion(128'h3643374bfc9b0483fce40ebf310203a0, {16'd59772, 16'd18213, 16'd6380, 16'd53041, 16'd17215, 16'd33122, 16'd63960, 16'd7973, 16'd59498, 16'd16734, 16'd57831, 16'd9573, 16'd60141, 16'd57957, 16'd40365, 16'd9142, 16'd40689, 16'd58112, 16'd42744, 16'd63718, 16'd34910, 16'd44857, 16'd64636, 16'd862, 16'd54721, 16'd16042});
	test_expansion(128'h5d4acafbaf2a982aa4c6a2813c490f6b, {16'd51378, 16'd39345, 16'd10331, 16'd25056, 16'd26470, 16'd62627, 16'd23937, 16'd32481, 16'd42306, 16'd46580, 16'd28619, 16'd3206, 16'd39163, 16'd48434, 16'd5238, 16'd18388, 16'd57, 16'd8960, 16'd34326, 16'd40863, 16'd18586, 16'd46733, 16'd45246, 16'd24654, 16'd64159, 16'd31794});
	test_expansion(128'h9ac81e9466473fbbed600e6b2d858ba5, {16'd27576, 16'd42792, 16'd38305, 16'd31127, 16'd57715, 16'd49162, 16'd36663, 16'd52847, 16'd61217, 16'd61185, 16'd56025, 16'd45282, 16'd64639, 16'd36997, 16'd36059, 16'd17953, 16'd14478, 16'd36861, 16'd31486, 16'd16143, 16'd64647, 16'd24731, 16'd31023, 16'd21298, 16'd65358, 16'd14859});
	test_expansion(128'h11f6ddaf4ce2f1acd4e5f8d9992b9d93, {16'd23498, 16'd17390, 16'd54039, 16'd36568, 16'd7602, 16'd21852, 16'd61912, 16'd7408, 16'd50465, 16'd36282, 16'd26351, 16'd65026, 16'd11691, 16'd10011, 16'd59584, 16'd20843, 16'd58707, 16'd34431, 16'd21140, 16'd5192, 16'd18301, 16'd61591, 16'd57969, 16'd29966, 16'd48539, 16'd8596});
	test_expansion(128'hfce6764f2f7df0566bf6a4b77b8978a7, {16'd55048, 16'd30032, 16'd57057, 16'd59484, 16'd30886, 16'd7860, 16'd14236, 16'd52701, 16'd18690, 16'd43059, 16'd59559, 16'd14423, 16'd62849, 16'd38546, 16'd21272, 16'd8517, 16'd41886, 16'd50411, 16'd22008, 16'd22331, 16'd37945, 16'd7891, 16'd65075, 16'd38327, 16'd6355, 16'd24605});
	test_expansion(128'h50abd361247615bd03bab96235ecd8e9, {16'd17019, 16'd19840, 16'd41020, 16'd17888, 16'd52558, 16'd54204, 16'd50427, 16'd14836, 16'd42241, 16'd6121, 16'd44124, 16'd38790, 16'd38037, 16'd7517, 16'd46159, 16'd46263, 16'd22597, 16'd40242, 16'd44403, 16'd20150, 16'd9100, 16'd46545, 16'd34693, 16'd31910, 16'd14063, 16'd35980});
	test_expansion(128'h098d60663a7097e31d0147aa2138282f, {16'd26980, 16'd20720, 16'd36989, 16'd30726, 16'd15809, 16'd1035, 16'd23593, 16'd35712, 16'd34252, 16'd25054, 16'd2184, 16'd20882, 16'd58018, 16'd29377, 16'd20799, 16'd27325, 16'd23074, 16'd1639, 16'd6533, 16'd15193, 16'd18773, 16'd36427, 16'd35011, 16'd31638, 16'd10944, 16'd51389});
	test_expansion(128'h11c751ba3287ad44899156e6c2917856, {16'd43430, 16'd8832, 16'd36044, 16'd52385, 16'd35152, 16'd16808, 16'd741, 16'd26739, 16'd63419, 16'd33119, 16'd13430, 16'd58272, 16'd1691, 16'd37705, 16'd57970, 16'd30245, 16'd59574, 16'd34419, 16'd17538, 16'd46241, 16'd27296, 16'd52152, 16'd17641, 16'd129, 16'd35917, 16'd55644});
	test_expansion(128'h78a4610c9139625a803186a3170a9609, {16'd49782, 16'd41790, 16'd20486, 16'd12925, 16'd34908, 16'd27232, 16'd7066, 16'd43471, 16'd29833, 16'd18843, 16'd51745, 16'd63119, 16'd40834, 16'd55329, 16'd12203, 16'd27540, 16'd37477, 16'd59897, 16'd59595, 16'd24135, 16'd34118, 16'd14990, 16'd49526, 16'd8373, 16'd55404, 16'd56074});
	test_expansion(128'h2d8f9b1d741ce8cd703ee3ab28146285, {16'd22181, 16'd38873, 16'd38174, 16'd22690, 16'd58652, 16'd4419, 16'd64212, 16'd8157, 16'd59422, 16'd4596, 16'd58944, 16'd42299, 16'd30254, 16'd4817, 16'd9023, 16'd64140, 16'd53524, 16'd55780, 16'd63487, 16'd43934, 16'd61148, 16'd62742, 16'd63433, 16'd34296, 16'd5672, 16'd37417});
	test_expansion(128'hacd33f4955bad200e830bbf191f4c345, {16'd32489, 16'd27057, 16'd40339, 16'd27369, 16'd5176, 16'd63654, 16'd27620, 16'd6044, 16'd42480, 16'd15253, 16'd20489, 16'd53269, 16'd63735, 16'd51089, 16'd46748, 16'd46939, 16'd16345, 16'd19223, 16'd25224, 16'd49412, 16'd49261, 16'd4274, 16'd47944, 16'd1477, 16'd53186, 16'd58536});
	test_expansion(128'hdff4075370dc633cfd35ea2fa3ab37d4, {16'd45788, 16'd12679, 16'd58354, 16'd48262, 16'd60594, 16'd2202, 16'd50022, 16'd37422, 16'd23332, 16'd27995, 16'd29388, 16'd15230, 16'd15930, 16'd13010, 16'd55969, 16'd8337, 16'd13882, 16'd10425, 16'd55765, 16'd53285, 16'd7175, 16'd21775, 16'd32554, 16'd388, 16'd26672, 16'd40052});
	test_expansion(128'hdb37e2e7cd6274914f146fdc369beabd, {16'd52918, 16'd43292, 16'd22605, 16'd42958, 16'd13821, 16'd19514, 16'd16380, 16'd63964, 16'd2645, 16'd47479, 16'd14887, 16'd45815, 16'd44443, 16'd57491, 16'd39289, 16'd61665, 16'd4693, 16'd52667, 16'd12460, 16'd48483, 16'd22024, 16'd27799, 16'd30239, 16'd28608, 16'd2983, 16'd8328});
	test_expansion(128'ha83d7472cf5978ab8a51d871273c79ee, {16'd53043, 16'd58520, 16'd64186, 16'd32328, 16'd51673, 16'd59434, 16'd51812, 16'd44568, 16'd10908, 16'd22714, 16'd26047, 16'd35707, 16'd35194, 16'd2243, 16'd24248, 16'd15961, 16'd59498, 16'd6370, 16'd11204, 16'd20069, 16'd58738, 16'd20131, 16'd17320, 16'd6334, 16'd10432, 16'd5641});
	test_expansion(128'hac6da7883957844b5473020592aec66b, {16'd35617, 16'd38583, 16'd51466, 16'd20037, 16'd23082, 16'd43025, 16'd12683, 16'd5703, 16'd15897, 16'd11798, 16'd36154, 16'd36351, 16'd45124, 16'd40806, 16'd39585, 16'd44784, 16'd56586, 16'd46802, 16'd6791, 16'd16894, 16'd39507, 16'd18127, 16'd59723, 16'd51159, 16'd6730, 16'd29386});
	test_expansion(128'h60b9d6520216a57b642629c20f97c910, {16'd5723, 16'd65506, 16'd20950, 16'd20666, 16'd2523, 16'd39752, 16'd47465, 16'd31122, 16'd50279, 16'd414, 16'd65161, 16'd25468, 16'd56025, 16'd5699, 16'd53383, 16'd23728, 16'd61168, 16'd25588, 16'd37299, 16'd19652, 16'd48508, 16'd52340, 16'd55366, 16'd64692, 16'd19772, 16'd52903});
	test_expansion(128'hab83cf39841e4108c033fe4f2aea3243, {16'd43942, 16'd52686, 16'd2931, 16'd13370, 16'd50039, 16'd24321, 16'd14642, 16'd30425, 16'd62482, 16'd1328, 16'd59787, 16'd47995, 16'd30335, 16'd23433, 16'd59396, 16'd21481, 16'd38565, 16'd60682, 16'd58973, 16'd13383, 16'd12861, 16'd24909, 16'd4882, 16'd53609, 16'd48424, 16'd53607});
	test_expansion(128'h2c949f692a890ee2dcc0b5969c61b6d4, {16'd59174, 16'd12771, 16'd21445, 16'd39730, 16'd1407, 16'd43285, 16'd47469, 16'd63796, 16'd12872, 16'd11272, 16'd12886, 16'd27611, 16'd56729, 16'd34539, 16'd51471, 16'd21318, 16'd46649, 16'd11066, 16'd22782, 16'd59792, 16'd32690, 16'd12685, 16'd32342, 16'd6943, 16'd9088, 16'd54034});
	test_expansion(128'h555f5849cf5054074ee269312cfbd3f9, {16'd8637, 16'd56225, 16'd48021, 16'd7141, 16'd11458, 16'd60269, 16'd15499, 16'd47331, 16'd13670, 16'd45064, 16'd59638, 16'd34081, 16'd62977, 16'd11830, 16'd17865, 16'd12578, 16'd61344, 16'd19600, 16'd14670, 16'd23252, 16'd40669, 16'd13446, 16'd19966, 16'd5043, 16'd19068, 16'd396});
	test_expansion(128'he5e513cf4e3a2712a0469ace5011a130, {16'd7091, 16'd8670, 16'd7579, 16'd55541, 16'd696, 16'd8763, 16'd63236, 16'd40332, 16'd54269, 16'd56231, 16'd35164, 16'd16786, 16'd46940, 16'd18486, 16'd55839, 16'd41667, 16'd18733, 16'd24042, 16'd19246, 16'd22924, 16'd35480, 16'd1476, 16'd47219, 16'd59947, 16'd3038, 16'd36053});
	test_expansion(128'hfac55ff094e10174434bb103aa27d4a0, {16'd45929, 16'd63079, 16'd53822, 16'd22542, 16'd7237, 16'd17045, 16'd6894, 16'd26421, 16'd25132, 16'd48146, 16'd9130, 16'd34519, 16'd18587, 16'd1112, 16'd43678, 16'd7242, 16'd7437, 16'd21968, 16'd3166, 16'd15813, 16'd63419, 16'd28140, 16'd226, 16'd47366, 16'd660, 16'd14440});
	test_expansion(128'hc24bcc1076a7457a092ff9cc78802cd9, {16'd45026, 16'd40886, 16'd42268, 16'd56991, 16'd40662, 16'd10370, 16'd53772, 16'd50238, 16'd17666, 16'd6727, 16'd27276, 16'd21576, 16'd62180, 16'd22088, 16'd53339, 16'd19539, 16'd52360, 16'd7593, 16'd17439, 16'd31018, 16'd33252, 16'd6952, 16'd60231, 16'd24295, 16'd36585, 16'd61931});
	test_expansion(128'h1c4faa5b3ece023b8115d9d12d1b39f1, {16'd35095, 16'd33219, 16'd62516, 16'd30304, 16'd25526, 16'd3717, 16'd59508, 16'd48830, 16'd39998, 16'd53171, 16'd62153, 16'd19518, 16'd62047, 16'd46039, 16'd24972, 16'd63233, 16'd17810, 16'd58079, 16'd43491, 16'd23507, 16'd22183, 16'd51738, 16'd50997, 16'd8553, 16'd42368, 16'd3085});
	test_expansion(128'hfe55a8317d8dfcd6a5fa3f977d1a0f0e, {16'd27885, 16'd53138, 16'd41652, 16'd52995, 16'd16324, 16'd33733, 16'd40768, 16'd5995, 16'd26966, 16'd36119, 16'd5717, 16'd30722, 16'd19638, 16'd40693, 16'd35251, 16'd12006, 16'd39073, 16'd54597, 16'd3492, 16'd17724, 16'd2808, 16'd24989, 16'd27254, 16'd30460, 16'd4343, 16'd58020});
	test_expansion(128'hd524e472efb2b83b56049702af2a4477, {16'd23493, 16'd26656, 16'd16565, 16'd48499, 16'd24340, 16'd9483, 16'd7201, 16'd11401, 16'd46136, 16'd956, 16'd45140, 16'd24676, 16'd48348, 16'd4436, 16'd53828, 16'd23398, 16'd6210, 16'd52808, 16'd4300, 16'd64640, 16'd36861, 16'd12439, 16'd1297, 16'd28210, 16'd43650, 16'd36950});
	test_expansion(128'hf02632b27d1f7e2d91a3b4d5f206d325, {16'd54563, 16'd61411, 16'd53250, 16'd486, 16'd26037, 16'd41957, 16'd32108, 16'd45032, 16'd58435, 16'd4527, 16'd49373, 16'd49658, 16'd48245, 16'd39551, 16'd39215, 16'd58665, 16'd47760, 16'd45263, 16'd57808, 16'd36291, 16'd33264, 16'd25798, 16'd57694, 16'd32069, 16'd49505, 16'd42031});
	test_expansion(128'h966aacb31fa49630731c2d968b9d8557, {16'd21742, 16'd65112, 16'd23882, 16'd19009, 16'd24434, 16'd49347, 16'd56135, 16'd62480, 16'd8401, 16'd9546, 16'd41759, 16'd65127, 16'd8609, 16'd43163, 16'd25650, 16'd41887, 16'd59358, 16'd5, 16'd6072, 16'd14756, 16'd60837, 16'd19216, 16'd13928, 16'd30156, 16'd21658, 16'd56958});
	test_expansion(128'h73709d3ebd70e79565c2f419f93fc7e8, {16'd47379, 16'd52081, 16'd38854, 16'd34625, 16'd47890, 16'd268, 16'd22480, 16'd30247, 16'd22975, 16'd10018, 16'd39629, 16'd35535, 16'd17719, 16'd45032, 16'd11171, 16'd24747, 16'd14959, 16'd4741, 16'd6325, 16'd8257, 16'd28776, 16'd40591, 16'd5928, 16'd60872, 16'd56994, 16'd38416});
	test_expansion(128'h7e61fa43531136f3567d9de33ff4deae, {16'd18184, 16'd21117, 16'd60715, 16'd30466, 16'd50472, 16'd33829, 16'd27630, 16'd36119, 16'd45265, 16'd4860, 16'd37451, 16'd31005, 16'd535, 16'd6742, 16'd48505, 16'd27820, 16'd1456, 16'd27512, 16'd35792, 16'd46457, 16'd42569, 16'd42394, 16'd48459, 16'd15150, 16'd54146, 16'd37597});
	test_expansion(128'h2d55fc56f61b3bd2150f780b3b4c9fab, {16'd13193, 16'd10238, 16'd61307, 16'd27672, 16'd48100, 16'd11227, 16'd25093, 16'd17813, 16'd32850, 16'd34164, 16'd23785, 16'd30552, 16'd15714, 16'd13994, 16'd60574, 16'd25895, 16'd37070, 16'd64690, 16'd27747, 16'd32560, 16'd32066, 16'd57423, 16'd10565, 16'd58542, 16'd7848, 16'd10581});
	test_expansion(128'h5d94593a0c4da672dfa731b4ce132177, {16'd14251, 16'd15033, 16'd40244, 16'd8503, 16'd25208, 16'd41869, 16'd28362, 16'd15179, 16'd65241, 16'd64719, 16'd38767, 16'd32212, 16'd62950, 16'd2826, 16'd41621, 16'd10756, 16'd878, 16'd17067, 16'd35028, 16'd21901, 16'd16378, 16'd14705, 16'd65465, 16'd16570, 16'd36877, 16'd47660});
	test_expansion(128'h28facf962fcc8f8e3112940d15fdc507, {16'd50305, 16'd29304, 16'd1460, 16'd13197, 16'd32634, 16'd34006, 16'd35417, 16'd48068, 16'd15127, 16'd5295, 16'd55710, 16'd27127, 16'd32794, 16'd63511, 16'd57946, 16'd45873, 16'd62904, 16'd11831, 16'd23250, 16'd3318, 16'd62425, 16'd4118, 16'd48685, 16'd50787, 16'd50897, 16'd63788});
	test_expansion(128'ha3cfc03b3e0b762dbd36383add7b0273, {16'd14599, 16'd4654, 16'd6176, 16'd42378, 16'd35216, 16'd20704, 16'd27659, 16'd18956, 16'd369, 16'd53411, 16'd3962, 16'd59871, 16'd1955, 16'd21208, 16'd21283, 16'd7989, 16'd26596, 16'd3399, 16'd3086, 16'd65131, 16'd57573, 16'd47816, 16'd24307, 16'd6712, 16'd39940, 16'd8543});
	test_expansion(128'h97cd69851e9af9a477bdb481926a190e, {16'd6930, 16'd15645, 16'd27786, 16'd63707, 16'd45971, 16'd14580, 16'd18271, 16'd40669, 16'd15152, 16'd42204, 16'd8552, 16'd14727, 16'd50171, 16'd55635, 16'd25183, 16'd1559, 16'd37897, 16'd13640, 16'd43327, 16'd24129, 16'd46203, 16'd40215, 16'd58292, 16'd6540, 16'd17002, 16'd9269});
	test_expansion(128'h3875ef8a94a39c0a9bf8ebe8d03f8a12, {16'd32809, 16'd11386, 16'd43652, 16'd56989, 16'd17055, 16'd1642, 16'd45072, 16'd15512, 16'd20893, 16'd2234, 16'd5227, 16'd42765, 16'd32611, 16'd997, 16'd16744, 16'd35579, 16'd50086, 16'd27847, 16'd29347, 16'd29784, 16'd43579, 16'd45737, 16'd53931, 16'd2269, 16'd38195, 16'd45142});
	test_expansion(128'hbdec2a747a1027e1cc8701afaab0b180, {16'd14120, 16'd28598, 16'd21987, 16'd2295, 16'd5963, 16'd18765, 16'd40228, 16'd28607, 16'd18609, 16'd4809, 16'd30008, 16'd6886, 16'd16993, 16'd11237, 16'd57875, 16'd37073, 16'd36420, 16'd35638, 16'd31222, 16'd56796, 16'd14786, 16'd4990, 16'd59347, 16'd27490, 16'd7564, 16'd44251});
	test_expansion(128'hc58b637f823624a892c226df9f39172d, {16'd29403, 16'd44951, 16'd12222, 16'd15770, 16'd16776, 16'd3597, 16'd58329, 16'd19579, 16'd1432, 16'd10420, 16'd59182, 16'd3686, 16'd31939, 16'd35914, 16'd11519, 16'd58420, 16'd21167, 16'd7777, 16'd56553, 16'd38109, 16'd52384, 16'd3615, 16'd18043, 16'd34621, 16'd22045, 16'd9011});
	test_expansion(128'h596834cad232b2860628217f1c6eff77, {16'd5151, 16'd52519, 16'd12509, 16'd33082, 16'd20691, 16'd24907, 16'd44935, 16'd42016, 16'd47746, 16'd32255, 16'd48992, 16'd54168, 16'd42693, 16'd52347, 16'd27651, 16'd39692, 16'd57350, 16'd16999, 16'd21618, 16'd100, 16'd55339, 16'd18685, 16'd56628, 16'd44988, 16'd4986, 16'd48675});
	test_expansion(128'h04d1c527f2f4b4c4452713bdecb7bdcc, {16'd19985, 16'd57860, 16'd24496, 16'd47303, 16'd36093, 16'd21022, 16'd63882, 16'd18226, 16'd56888, 16'd27572, 16'd14594, 16'd18110, 16'd30088, 16'd52878, 16'd48816, 16'd10028, 16'd21925, 16'd24107, 16'd41733, 16'd65530, 16'd16343, 16'd3600, 16'd16757, 16'd2677, 16'd18402, 16'd37554});
	test_expansion(128'hf20ff40d2b2b9554e695378d8ae55aa6, {16'd47899, 16'd41161, 16'd35256, 16'd39079, 16'd47654, 16'd48584, 16'd57047, 16'd45882, 16'd54191, 16'd38591, 16'd2258, 16'd60247, 16'd62016, 16'd44746, 16'd48983, 16'd33229, 16'd21611, 16'd64372, 16'd16730, 16'd34388, 16'd12898, 16'd12939, 16'd5090, 16'd9050, 16'd59302, 16'd65309});
	test_expansion(128'ha2aaef8f6fcda26f232aeeca838810fd, {16'd43299, 16'd47356, 16'd13532, 16'd31259, 16'd11457, 16'd29579, 16'd17375, 16'd33966, 16'd55537, 16'd56058, 16'd32240, 16'd43420, 16'd52672, 16'd63829, 16'd2585, 16'd29206, 16'd52522, 16'd42504, 16'd30169, 16'd41463, 16'd42357, 16'd40271, 16'd21496, 16'd55074, 16'd15582, 16'd61386});
	test_expansion(128'h0626783a151c57ed77c384644f3bc773, {16'd21787, 16'd18872, 16'd36286, 16'd47595, 16'd12958, 16'd25490, 16'd55669, 16'd1146, 16'd39416, 16'd53331, 16'd20637, 16'd10299, 16'd53327, 16'd48332, 16'd28831, 16'd31165, 16'd16099, 16'd39642, 16'd50421, 16'd64533, 16'd22106, 16'd12163, 16'd44806, 16'd33835, 16'd26793, 16'd21113});
	test_expansion(128'hf18b564e87626ead8c1e10dde4efbadf, {16'd11917, 16'd42313, 16'd15380, 16'd294, 16'd40384, 16'd58835, 16'd44989, 16'd52855, 16'd246, 16'd21762, 16'd9308, 16'd20074, 16'd49703, 16'd53529, 16'd9715, 16'd6710, 16'd904, 16'd61985, 16'd58907, 16'd20657, 16'd14076, 16'd24906, 16'd59830, 16'd21947, 16'd41945, 16'd36068});
	test_expansion(128'h6592f96071cbe55dd6735a8b71ca6fba, {16'd31473, 16'd40763, 16'd240, 16'd26822, 16'd5645, 16'd53097, 16'd53564, 16'd27942, 16'd56408, 16'd18239, 16'd2061, 16'd44078, 16'd38367, 16'd54584, 16'd19332, 16'd16002, 16'd25870, 16'd31424, 16'd8546, 16'd9645, 16'd5916, 16'd54755, 16'd9631, 16'd42491, 16'd46263, 16'd1694});
	test_expansion(128'h38682635a6357bacd00eb3071ed9e601, {16'd44232, 16'd45391, 16'd32619, 16'd43073, 16'd5831, 16'd24146, 16'd5120, 16'd65139, 16'd21178, 16'd16310, 16'd2906, 16'd55753, 16'd5164, 16'd41131, 16'd12597, 16'd49287, 16'd62283, 16'd10502, 16'd62220, 16'd14687, 16'd42077, 16'd9500, 16'd59750, 16'd13706, 16'd17999, 16'd32350});
	test_expansion(128'h4690271a4cfa91dc32d56df911bff1e8, {16'd11258, 16'd5802, 16'd26201, 16'd11575, 16'd47542, 16'd26592, 16'd32161, 16'd35949, 16'd64560, 16'd17846, 16'd48253, 16'd61692, 16'd45985, 16'd46445, 16'd20615, 16'd27690, 16'd45996, 16'd42944, 16'd31740, 16'd32383, 16'd65425, 16'd62437, 16'd8253, 16'd48953, 16'd22694, 16'd19576});
	test_expansion(128'h22f39de64b962eede03f33e0d7e4f6ed, {16'd25569, 16'd29610, 16'd28288, 16'd17343, 16'd13975, 16'd37329, 16'd43816, 16'd2378, 16'd33226, 16'd803, 16'd46445, 16'd60006, 16'd25309, 16'd13152, 16'd55853, 16'd20004, 16'd5251, 16'd30509, 16'd26141, 16'd16071, 16'd5719, 16'd47621, 16'd41405, 16'd50616, 16'd10941, 16'd57428});
	test_expansion(128'h2ba26c7f941ac20d2425e5d3ac4f57a9, {16'd17447, 16'd64606, 16'd53457, 16'd25732, 16'd59724, 16'd40529, 16'd60500, 16'd31852, 16'd38770, 16'd16395, 16'd62525, 16'd65453, 16'd16399, 16'd29023, 16'd34894, 16'd44562, 16'd6172, 16'd39227, 16'd40483, 16'd1758, 16'd11936, 16'd23532, 16'd21849, 16'd3212, 16'd7629, 16'd40287});
	test_expansion(128'h0af4616d054d674191e23adc3f0e5946, {16'd12483, 16'd57648, 16'd31358, 16'd3740, 16'd47012, 16'd25087, 16'd40658, 16'd18527, 16'd47759, 16'd55722, 16'd18614, 16'd29200, 16'd16483, 16'd39452, 16'd25426, 16'd10787, 16'd28879, 16'd28319, 16'd7306, 16'd3691, 16'd60247, 16'd63205, 16'd6905, 16'd6290, 16'd1046, 16'd24390});
	test_expansion(128'h9ed7d76adc0190870971256b3177224f, {16'd19140, 16'd43558, 16'd14673, 16'd1338, 16'd55759, 16'd55790, 16'd42460, 16'd26088, 16'd18426, 16'd43848, 16'd46069, 16'd12127, 16'd17731, 16'd21595, 16'd43932, 16'd18058, 16'd18875, 16'd11712, 16'd38534, 16'd58562, 16'd35636, 16'd57956, 16'd38771, 16'd39266, 16'd19939, 16'd21314});
	test_expansion(128'h23a9b303e62aadcb8a16b1e9b5530a6e, {16'd14205, 16'd46939, 16'd62210, 16'd44534, 16'd46870, 16'd37507, 16'd9012, 16'd24999, 16'd3002, 16'd8259, 16'd23928, 16'd51008, 16'd7047, 16'd14264, 16'd22346, 16'd23332, 16'd6303, 16'd50061, 16'd30920, 16'd20718, 16'd55089, 16'd63448, 16'd43703, 16'd56172, 16'd49305, 16'd2147});
	test_expansion(128'h544cf4c705febe6535f76702fcc65988, {16'd46275, 16'd38942, 16'd3222, 16'd6137, 16'd18264, 16'd31077, 16'd42626, 16'd4254, 16'd5392, 16'd44139, 16'd35848, 16'd12800, 16'd5091, 16'd37999, 16'd14868, 16'd63992, 16'd17944, 16'd44848, 16'd22492, 16'd30770, 16'd59933, 16'd19203, 16'd46397, 16'd1193, 16'd4642, 16'd14295});
	test_expansion(128'h16f74c45bf341419af744bb3c70ae614, {16'd23547, 16'd22469, 16'd34493, 16'd19230, 16'd53989, 16'd56770, 16'd14460, 16'd32163, 16'd7895, 16'd53729, 16'd60906, 16'd36917, 16'd5894, 16'd42172, 16'd15994, 16'd32361, 16'd25040, 16'd26932, 16'd46222, 16'd24587, 16'd31430, 16'd61236, 16'd49257, 16'd56268, 16'd5418, 16'd46998});
	test_expansion(128'h9e15aa9e6a34a4a314d2c6f033c25f96, {16'd12687, 16'd52929, 16'd53634, 16'd46351, 16'd20202, 16'd55201, 16'd28839, 16'd22911, 16'd5066, 16'd38887, 16'd36370, 16'd46800, 16'd17782, 16'd32015, 16'd22446, 16'd45482, 16'd16846, 16'd18642, 16'd48029, 16'd12557, 16'd63073, 16'd9867, 16'd51561, 16'd1372, 16'd63928, 16'd2195});
	test_expansion(128'hbc57637b98f625cff1d161afe2a5cb3f, {16'd18465, 16'd34701, 16'd49334, 16'd43316, 16'd53124, 16'd44428, 16'd31681, 16'd37384, 16'd17238, 16'd15894, 16'd47307, 16'd37668, 16'd57897, 16'd45479, 16'd62863, 16'd36460, 16'd30867, 16'd64065, 16'd56683, 16'd48456, 16'd49725, 16'd6630, 16'd40947, 16'd63396, 16'd37279, 16'd16677});
	test_expansion(128'h46d7d667b9aead2194eeba722a71a2ab, {16'd17193, 16'd58783, 16'd5532, 16'd3203, 16'd56419, 16'd10316, 16'd31184, 16'd4804, 16'd51108, 16'd44575, 16'd38681, 16'd64173, 16'd50058, 16'd55456, 16'd46117, 16'd51786, 16'd62936, 16'd19552, 16'd32107, 16'd21432, 16'd39197, 16'd57094, 16'd14087, 16'd27688, 16'd3432, 16'd11678});
	test_expansion(128'h400e575449d8ed6d074d7ad70de96bee, {16'd22559, 16'd64085, 16'd12210, 16'd1938, 16'd29610, 16'd40932, 16'd33540, 16'd22835, 16'd58292, 16'd54578, 16'd1375, 16'd60965, 16'd11423, 16'd37551, 16'd62752, 16'd26940, 16'd34319, 16'd1719, 16'd8955, 16'd57252, 16'd34010, 16'd27977, 16'd791, 16'd2490, 16'd56291, 16'd19720});
	test_expansion(128'h79e460836c5aa8f358d75e4a068b0fc7, {16'd62868, 16'd7889, 16'd10764, 16'd57077, 16'd40769, 16'd2906, 16'd49647, 16'd45644, 16'd16436, 16'd22515, 16'd40881, 16'd48063, 16'd763, 16'd41447, 16'd28016, 16'd24880, 16'd40764, 16'd56078, 16'd8883, 16'd20181, 16'd64485, 16'd40421, 16'd25293, 16'd46089, 16'd46819, 16'd14598});
	test_expansion(128'h4859ed6728f5c9401420310e6892bcac, {16'd49651, 16'd9757, 16'd34216, 16'd38409, 16'd50086, 16'd11756, 16'd13539, 16'd34187, 16'd17283, 16'd16058, 16'd15773, 16'd12569, 16'd62185, 16'd33642, 16'd62903, 16'd2006, 16'd14441, 16'd6782, 16'd9250, 16'd4404, 16'd37961, 16'd17747, 16'd63353, 16'd62414, 16'd53582, 16'd5570});
	test_expansion(128'h759f786110362bfa1de814d2c4935a4a, {16'd2351, 16'd24509, 16'd17084, 16'd13957, 16'd32230, 16'd65353, 16'd15841, 16'd26008, 16'd45989, 16'd20599, 16'd61545, 16'd11780, 16'd10991, 16'd20464, 16'd57766, 16'd8430, 16'd35982, 16'd17111, 16'd57148, 16'd47715, 16'd43055, 16'd21449, 16'd40420, 16'd34451, 16'd42015, 16'd12826});
	test_expansion(128'h7517ce865fe63b83c28ef5299ebc3deb, {16'd23803, 16'd18335, 16'd50482, 16'd38169, 16'd13541, 16'd4925, 16'd39354, 16'd59607, 16'd51970, 16'd61456, 16'd3016, 16'd24444, 16'd54353, 16'd26839, 16'd61762, 16'd44627, 16'd24464, 16'd26612, 16'd36593, 16'd340, 16'd40808, 16'd22373, 16'd9018, 16'd63786, 16'd30046, 16'd41569});
	test_expansion(128'h14a48d26a0d2b99a761a2ff791a404b5, {16'd18204, 16'd34295, 16'd39172, 16'd44411, 16'd8342, 16'd42054, 16'd14681, 16'd60582, 16'd4259, 16'd38254, 16'd4879, 16'd13760, 16'd10736, 16'd25807, 16'd17822, 16'd43930, 16'd17135, 16'd37996, 16'd58009, 16'd45943, 16'd21250, 16'd36773, 16'd63848, 16'd28482, 16'd59940, 16'd55999});
	test_expansion(128'hf71fa2163d0dff74050e2ffe4b47286d, {16'd5475, 16'd41756, 16'd25996, 16'd34146, 16'd33819, 16'd35261, 16'd51469, 16'd58009, 16'd24036, 16'd40659, 16'd56276, 16'd48088, 16'd15999, 16'd61870, 16'd30034, 16'd5254, 16'd35881, 16'd40712, 16'd55357, 16'd31989, 16'd34645, 16'd412, 16'd34873, 16'd20373, 16'd56932, 16'd50327});
	test_expansion(128'h50c5635ce305b6c994182f0a806e74b3, {16'd60797, 16'd15852, 16'd28257, 16'd16177, 16'd45720, 16'd22786, 16'd30918, 16'd15072, 16'd39022, 16'd29451, 16'd46214, 16'd41708, 16'd37863, 16'd11529, 16'd38203, 16'd31473, 16'd55642, 16'd21056, 16'd24178, 16'd21954, 16'd23098, 16'd52990, 16'd10342, 16'd18665, 16'd7311, 16'd4389});
	test_expansion(128'h693d196fa32228326205310dc86086bb, {16'd21016, 16'd36897, 16'd59554, 16'd39231, 16'd19876, 16'd11693, 16'd42438, 16'd39632, 16'd63880, 16'd5718, 16'd25254, 16'd44368, 16'd31236, 16'd1388, 16'd52168, 16'd10563, 16'd33338, 16'd23237, 16'd43683, 16'd59215, 16'd56964, 16'd33344, 16'd14525, 16'd44700, 16'd44585, 16'd3598});
	test_expansion(128'he306d15a9ce69f13d7a0414f2a64588f, {16'd21631, 16'd15106, 16'd37528, 16'd48604, 16'd58394, 16'd26499, 16'd50712, 16'd24683, 16'd51387, 16'd38408, 16'd45629, 16'd56474, 16'd42785, 16'd50411, 16'd45267, 16'd58797, 16'd46959, 16'd23029, 16'd26738, 16'd16811, 16'd29582, 16'd65113, 16'd57235, 16'd777, 16'd55477, 16'd64460});
	test_expansion(128'h7a37fd1e2e3af8f962a332d44c7f647b, {16'd64071, 16'd35925, 16'd41614, 16'd39866, 16'd4065, 16'd14325, 16'd30305, 16'd11116, 16'd45823, 16'd31070, 16'd44502, 16'd59898, 16'd20904, 16'd46664, 16'd38695, 16'd63100, 16'd43790, 16'd55697, 16'd56328, 16'd27656, 16'd8398, 16'd51780, 16'd58529, 16'd14798, 16'd48144, 16'd49363});
	test_expansion(128'h2ca55c837aa5edc4e88bd54e18e4f527, {16'd4059, 16'd43330, 16'd15274, 16'd62453, 16'd2775, 16'd60109, 16'd62337, 16'd31514, 16'd26570, 16'd15924, 16'd21583, 16'd9916, 16'd61730, 16'd47348, 16'd22971, 16'd38905, 16'd58316, 16'd5267, 16'd8396, 16'd4083, 16'd45940, 16'd61667, 16'd222, 16'd10549, 16'd48857, 16'd43184});
	test_expansion(128'h2e8ba8f7ad2ae7c4407afe7690b0ac09, {16'd54375, 16'd60123, 16'd10861, 16'd28971, 16'd13508, 16'd41285, 16'd45432, 16'd25550, 16'd50563, 16'd27649, 16'd29324, 16'd54267, 16'd64723, 16'd55764, 16'd47241, 16'd22325, 16'd46127, 16'd37009, 16'd10584, 16'd3594, 16'd33894, 16'd9122, 16'd15948, 16'd65531, 16'd13011, 16'd63957});
	test_expansion(128'h608da01fd99e356b022effec5cbe0e8e, {16'd25932, 16'd2321, 16'd45612, 16'd51625, 16'd448, 16'd22481, 16'd57699, 16'd59499, 16'd11866, 16'd5262, 16'd60226, 16'd27411, 16'd7531, 16'd29977, 16'd59375, 16'd20676, 16'd49667, 16'd34463, 16'd4222, 16'd57986, 16'd46317, 16'd23413, 16'd40338, 16'd63630, 16'd37418, 16'd58767});
	test_expansion(128'h389057e66e6bc5cfaee8d82e46f9ced8, {16'd38941, 16'd36471, 16'd52248, 16'd27375, 16'd17487, 16'd33696, 16'd20804, 16'd49698, 16'd18674, 16'd2151, 16'd18478, 16'd31635, 16'd6241, 16'd30464, 16'd32967, 16'd42849, 16'd37689, 16'd38653, 16'd52596, 16'd6860, 16'd30479, 16'd26112, 16'd6504, 16'd51827, 16'd56434, 16'd48309});
	test_expansion(128'hf81ba1606a11a8f21f8bf0923d09f5cd, {16'd9772, 16'd52457, 16'd56073, 16'd48756, 16'd37894, 16'd1915, 16'd24443, 16'd56549, 16'd48833, 16'd54673, 16'd34263, 16'd394, 16'd24862, 16'd30931, 16'd31222, 16'd8566, 16'd21392, 16'd10898, 16'd47998, 16'd34918, 16'd39664, 16'd56208, 16'd8101, 16'd60082, 16'd54436, 16'd25392});
	test_expansion(128'hc3b4227987af79541da9430220e64060, {16'd388, 16'd60287, 16'd31829, 16'd23628, 16'd20140, 16'd10863, 16'd36691, 16'd16259, 16'd6015, 16'd28976, 16'd10766, 16'd39590, 16'd51113, 16'd50116, 16'd60143, 16'd59677, 16'd46505, 16'd2522, 16'd8671, 16'd60683, 16'd57469, 16'd44971, 16'd27819, 16'd24359, 16'd36461, 16'd65514});
	test_expansion(128'ha17a2881a9935788a4a4ce6023e822c7, {16'd40072, 16'd16965, 16'd14225, 16'd10874, 16'd8663, 16'd9992, 16'd8437, 16'd53961, 16'd56215, 16'd17658, 16'd49107, 16'd37119, 16'd48661, 16'd5827, 16'd48955, 16'd59553, 16'd19005, 16'd51359, 16'd28672, 16'd6597, 16'd1912, 16'd41544, 16'd48019, 16'd50659, 16'd21990, 16'd42958});
	test_expansion(128'h8c05732209dc751f5f4a31b556e4dcef, {16'd64476, 16'd64888, 16'd5007, 16'd18793, 16'd55646, 16'd51481, 16'd10649, 16'd8691, 16'd31452, 16'd35166, 16'd64237, 16'd21233, 16'd11983, 16'd65049, 16'd24528, 16'd8397, 16'd34299, 16'd40670, 16'd48599, 16'd51238, 16'd60382, 16'd20175, 16'd357, 16'd58491, 16'd13745, 16'd47721});
	test_expansion(128'h7f636b3fd6161b3ea8ff8063ee50235e, {16'd22036, 16'd20339, 16'd43054, 16'd7566, 16'd56174, 16'd9928, 16'd18017, 16'd59634, 16'd13783, 16'd29656, 16'd5770, 16'd52859, 16'd7822, 16'd42932, 16'd53661, 16'd25843, 16'd20264, 16'd21344, 16'd15398, 16'd20956, 16'd19734, 16'd44494, 16'd51831, 16'd41930, 16'd23203, 16'd13076});
	test_expansion(128'h9e50ae08aec824c1f46433ee2999d2c1, {16'd32580, 16'd23013, 16'd57299, 16'd48881, 16'd17923, 16'd7869, 16'd29715, 16'd55797, 16'd1411, 16'd35598, 16'd54098, 16'd42734, 16'd24962, 16'd54827, 16'd16604, 16'd3007, 16'd4910, 16'd21630, 16'd30943, 16'd12693, 16'd28824, 16'd29431, 16'd62896, 16'd64548, 16'd55420, 16'd51474});
	test_expansion(128'he54f25a6461603a5281db59418edb3d9, {16'd27760, 16'd14187, 16'd35877, 16'd33188, 16'd58495, 16'd60779, 16'd20151, 16'd62599, 16'd59098, 16'd36005, 16'd35414, 16'd23088, 16'd59060, 16'd61137, 16'd53707, 16'd7131, 16'd18011, 16'd46924, 16'd43777, 16'd4928, 16'd30467, 16'd35111, 16'd52686, 16'd59142, 16'd15382, 16'd23868});
	test_expansion(128'hf426fe49ecde846f8e77df565927e9b3, {16'd63138, 16'd17805, 16'd11484, 16'd63123, 16'd34515, 16'd21469, 16'd55849, 16'd23913, 16'd58339, 16'd47472, 16'd51321, 16'd58187, 16'd15730, 16'd11361, 16'd57043, 16'd57590, 16'd44525, 16'd44628, 16'd55772, 16'd28371, 16'd18135, 16'd9734, 16'd42121, 16'd41856, 16'd42667, 16'd30414});
	test_expansion(128'he6606ccf4893e7bc239ceb81d7a2ee84, {16'd33665, 16'd23724, 16'd32432, 16'd3564, 16'd57991, 16'd46514, 16'd20027, 16'd46383, 16'd18150, 16'd9541, 16'd2715, 16'd29207, 16'd26348, 16'd25494, 16'd52508, 16'd2834, 16'd34151, 16'd63518, 16'd61772, 16'd23856, 16'd13411, 16'd34396, 16'd2878, 16'd30132, 16'd60010, 16'd9807});
	test_expansion(128'h0ae58c881652bf25af8e07793621a18d, {16'd46097, 16'd53272, 16'd48070, 16'd31649, 16'd13350, 16'd50137, 16'd63852, 16'd26759, 16'd51085, 16'd51156, 16'd46548, 16'd30161, 16'd7311, 16'd16568, 16'd38384, 16'd22403, 16'd23021, 16'd35208, 16'd26699, 16'd54989, 16'd3933, 16'd45229, 16'd16825, 16'd22707, 16'd43034, 16'd58515});
	test_expansion(128'hc93895a76dc499beb9d961b464d1085f, {16'd48654, 16'd34918, 16'd52380, 16'd38852, 16'd39809, 16'd18282, 16'd58041, 16'd3407, 16'd14654, 16'd56899, 16'd48960, 16'd14755, 16'd32893, 16'd54452, 16'd57393, 16'd6646, 16'd34914, 16'd41674, 16'd55485, 16'd65005, 16'd62701, 16'd17161, 16'd2128, 16'd3447, 16'd55141, 16'd43236});
	test_expansion(128'ha3a0cc6b6d3bf8ba3e9fa5fa2cc66899, {16'd11891, 16'd48116, 16'd31295, 16'd58114, 16'd2707, 16'd61179, 16'd15578, 16'd19347, 16'd32354, 16'd2650, 16'd33917, 16'd61663, 16'd43972, 16'd49533, 16'd36468, 16'd57433, 16'd6804, 16'd10776, 16'd4348, 16'd60177, 16'd49553, 16'd37883, 16'd45761, 16'd25115, 16'd37583, 16'd65383});
	test_expansion(128'h7917ff16a235b080a51113313af2b047, {16'd7663, 16'd63000, 16'd55758, 16'd48992, 16'd37464, 16'd35487, 16'd61727, 16'd24881, 16'd34962, 16'd50253, 16'd17044, 16'd57521, 16'd3957, 16'd4153, 16'd25595, 16'd56287, 16'd19849, 16'd45949, 16'd30962, 16'd30979, 16'd44930, 16'd18554, 16'd35064, 16'd44194, 16'd17965, 16'd22271});
	test_expansion(128'h3baa465c806d87dec13dbdbaf772d39d, {16'd39783, 16'd56503, 16'd61301, 16'd5350, 16'd55653, 16'd22838, 16'd34745, 16'd61006, 16'd48045, 16'd28047, 16'd57308, 16'd43001, 16'd32536, 16'd4065, 16'd50697, 16'd32715, 16'd59985, 16'd59521, 16'd23444, 16'd38243, 16'd41594, 16'd29317, 16'd22408, 16'd49882, 16'd15316, 16'd56596});
	test_expansion(128'hb5e7839900bd322814a78b7783de59fd, {16'd41549, 16'd21274, 16'd4804, 16'd46127, 16'd57746, 16'd46401, 16'd21447, 16'd47068, 16'd62395, 16'd52921, 16'd64203, 16'd13051, 16'd61247, 16'd55638, 16'd62990, 16'd55254, 16'd14, 16'd16378, 16'd64348, 16'd32730, 16'd25811, 16'd28204, 16'd7905, 16'd433, 16'd28985, 16'd23094});
	test_expansion(128'hbf7e2d8a8976f95e328d36a2286b63ba, {16'd61070, 16'd49756, 16'd42953, 16'd24960, 16'd41931, 16'd56883, 16'd23064, 16'd8452, 16'd24290, 16'd54866, 16'd3961, 16'd34228, 16'd53029, 16'd11324, 16'd36760, 16'd13052, 16'd59479, 16'd12842, 16'd43307, 16'd11668, 16'd44059, 16'd47256, 16'd23690, 16'd35566, 16'd4153, 16'd61812});
	test_expansion(128'h3045fa95b2deccab4d07df6d6857c15b, {16'd22026, 16'd34799, 16'd51223, 16'd14513, 16'd17012, 16'd8336, 16'd34581, 16'd10309, 16'd46509, 16'd37250, 16'd47836, 16'd5149, 16'd25321, 16'd352, 16'd56007, 16'd20460, 16'd18193, 16'd61816, 16'd15123, 16'd33634, 16'd62204, 16'd57076, 16'd33124, 16'd2381, 16'd18098, 16'd11651});
	test_expansion(128'h6f8ee1163bbeceb70ffe27a9a12e363d, {16'd29495, 16'd10675, 16'd55689, 16'd41548, 16'd48642, 16'd56037, 16'd52581, 16'd16383, 16'd32082, 16'd15016, 16'd13776, 16'd2753, 16'd40867, 16'd55135, 16'd19904, 16'd23442, 16'd2052, 16'd44396, 16'd48529, 16'd64375, 16'd37353, 16'd61552, 16'd55091, 16'd39905, 16'd50073, 16'd38});
	test_expansion(128'h687177af1c0d8efe0e8bcde84ebd048e, {16'd25537, 16'd16753, 16'd18496, 16'd41545, 16'd34788, 16'd2036, 16'd3182, 16'd43669, 16'd48786, 16'd32446, 16'd55889, 16'd64579, 16'd3123, 16'd16495, 16'd21563, 16'd42456, 16'd11342, 16'd2253, 16'd40888, 16'd59970, 16'd1534, 16'd48131, 16'd19658, 16'd2869, 16'd19317, 16'd41431});
	test_expansion(128'h038a448cf36c78392d53e243979c86c0, {16'd36270, 16'd45904, 16'd64941, 16'd20467, 16'd11296, 16'd14378, 16'd51185, 16'd37799, 16'd13142, 16'd9873, 16'd28197, 16'd11108, 16'd13582, 16'd5639, 16'd3033, 16'd41998, 16'd43318, 16'd3841, 16'd30730, 16'd43207, 16'd14104, 16'd27524, 16'd12738, 16'd7467, 16'd12372, 16'd23681});
	test_expansion(128'h0d7feff1ab77a0842a90856fb37aca5f, {16'd61629, 16'd51896, 16'd34649, 16'd58352, 16'd31578, 16'd64743, 16'd6456, 16'd8459, 16'd61470, 16'd65435, 16'd7639, 16'd58861, 16'd39224, 16'd8079, 16'd62006, 16'd55121, 16'd54373, 16'd53306, 16'd29423, 16'd65355, 16'd63497, 16'd23721, 16'd36427, 16'd53767, 16'd43515, 16'd60296});
	test_expansion(128'hce7816d0870bebd58a8a3e34c06dc7c1, {16'd51443, 16'd31436, 16'd62312, 16'd25678, 16'd4403, 16'd27830, 16'd26990, 16'd47961, 16'd59221, 16'd58399, 16'd59333, 16'd5345, 16'd2331, 16'd21494, 16'd30167, 16'd58616, 16'd42373, 16'd18504, 16'd50421, 16'd62829, 16'd50669, 16'd64134, 16'd22249, 16'd29393, 16'd7450, 16'd39351});
	test_expansion(128'h1735cd430828eedc22ce18af9119c926, {16'd62255, 16'd4055, 16'd6954, 16'd17760, 16'd58959, 16'd13866, 16'd36777, 16'd20407, 16'd13850, 16'd44040, 16'd51818, 16'd58059, 16'd19186, 16'd42984, 16'd19314, 16'd64991, 16'd55492, 16'd21835, 16'd58550, 16'd43492, 16'd54120, 16'd56314, 16'd3315, 16'd45216, 16'd5954, 16'd50739});
	test_expansion(128'h3071378a6de278bb500a9f16fdd1ddc4, {16'd21193, 16'd64695, 16'd28617, 16'd50391, 16'd64786, 16'd4114, 16'd58672, 16'd64303, 16'd10457, 16'd17379, 16'd19257, 16'd45486, 16'd55575, 16'd3493, 16'd24620, 16'd38927, 16'd25207, 16'd51521, 16'd56770, 16'd49732, 16'd27103, 16'd34246, 16'd45398, 16'd49915, 16'd31619, 16'd17351});
	test_expansion(128'h99dcd5930842019a349734d31a89b405, {16'd56159, 16'd232, 16'd52829, 16'd30375, 16'd49249, 16'd60128, 16'd65266, 16'd43190, 16'd57716, 16'd4820, 16'd22308, 16'd16715, 16'd60114, 16'd4606, 16'd13454, 16'd46383, 16'd40135, 16'd58982, 16'd55794, 16'd35015, 16'd26400, 16'd2249, 16'd31841, 16'd19826, 16'd49181, 16'd48067});
	test_expansion(128'h81341b42ef3490ca73369742cffa65af, {16'd24678, 16'd44634, 16'd53529, 16'd46439, 16'd34944, 16'd47839, 16'd19558, 16'd54775, 16'd23900, 16'd11783, 16'd51996, 16'd12621, 16'd61708, 16'd28120, 16'd31414, 16'd12029, 16'd41199, 16'd30157, 16'd8288, 16'd54201, 16'd48483, 16'd35729, 16'd35057, 16'd36285, 16'd44729, 16'd42556});
	test_expansion(128'hac7ed1039037b1328c1bc8d3cde27652, {16'd6549, 16'd47531, 16'd9015, 16'd12504, 16'd29843, 16'd23083, 16'd10956, 16'd53963, 16'd30406, 16'd5490, 16'd39299, 16'd16652, 16'd24313, 16'd17701, 16'd28150, 16'd4776, 16'd34179, 16'd16688, 16'd2072, 16'd20918, 16'd59787, 16'd16611, 16'd21480, 16'd28704, 16'd59847, 16'd4646});
	test_expansion(128'hd0d8012f192cc03fbc6cb3a569b83dd8, {16'd13428, 16'd50741, 16'd47652, 16'd63181, 16'd10566, 16'd60901, 16'd40906, 16'd44691, 16'd62778, 16'd12905, 16'd12743, 16'd55306, 16'd3024, 16'd32590, 16'd15036, 16'd62340, 16'd60503, 16'd14588, 16'd29552, 16'd24458, 16'd39687, 16'd18777, 16'd7684, 16'd19038, 16'd4695, 16'd5834});
	test_expansion(128'haaf0601e9e33b9f4ff1fdce3393c3a35, {16'd61864, 16'd56755, 16'd39447, 16'd5134, 16'd38885, 16'd56567, 16'd12537, 16'd7754, 16'd49823, 16'd38760, 16'd52798, 16'd49302, 16'd40013, 16'd47622, 16'd8274, 16'd44573, 16'd55295, 16'd54751, 16'd20959, 16'd18221, 16'd11101, 16'd47047, 16'd59351, 16'd14562, 16'd62789, 16'd47782});
	test_expansion(128'h4c74f892bb097edf8b9df2e354013705, {16'd20142, 16'd54645, 16'd21541, 16'd9607, 16'd36460, 16'd22402, 16'd33323, 16'd57647, 16'd35037, 16'd65094, 16'd15785, 16'd23454, 16'd51284, 16'd3926, 16'd1271, 16'd13497, 16'd41793, 16'd31975, 16'd33473, 16'd53238, 16'd58431, 16'd57829, 16'd13715, 16'd3104, 16'd52853, 16'd30183});
	test_expansion(128'hdc3ec853b403017b055fea46249efc19, {16'd14546, 16'd52989, 16'd3500, 16'd35473, 16'd38448, 16'd9834, 16'd11019, 16'd13363, 16'd27081, 16'd9799, 16'd45794, 16'd52118, 16'd23634, 16'd37586, 16'd64049, 16'd52617, 16'd20972, 16'd18543, 16'd52189, 16'd59886, 16'd64841, 16'd46266, 16'd9677, 16'd35778, 16'd5917, 16'd49785});
	test_expansion(128'hafa6ba60e471f0b1d3b6dc4d772ffa5e, {16'd31071, 16'd44659, 16'd15506, 16'd43739, 16'd58994, 16'd38457, 16'd39170, 16'd18309, 16'd57073, 16'd35129, 16'd8779, 16'd48149, 16'd39045, 16'd25840, 16'd6283, 16'd64585, 16'd8168, 16'd33404, 16'd46354, 16'd55153, 16'd28250, 16'd57940, 16'd13281, 16'd62797, 16'd59197, 16'd6888});
	test_expansion(128'h68b29d7fddd0162b61e92fe7ac497a3a, {16'd24940, 16'd38230, 16'd13475, 16'd1376, 16'd23258, 16'd2225, 16'd35013, 16'd17473, 16'd30993, 16'd24107, 16'd23222, 16'd3421, 16'd41085, 16'd32380, 16'd9711, 16'd17181, 16'd34297, 16'd45970, 16'd23411, 16'd43521, 16'd4616, 16'd49608, 16'd39881, 16'd59992, 16'd26606, 16'd8203});
	test_expansion(128'hdb7add035a4ec0c55fbea046ecaa4b42, {16'd63241, 16'd6864, 16'd22601, 16'd6235, 16'd29929, 16'd19554, 16'd21766, 16'd54446, 16'd59687, 16'd40647, 16'd44920, 16'd19897, 16'd32922, 16'd46794, 16'd14839, 16'd33731, 16'd26495, 16'd7030, 16'd22770, 16'd28107, 16'd54113, 16'd21285, 16'd54002, 16'd58672, 16'd54361, 16'd60383});
	test_expansion(128'h053d19c618462e03cf4db9070e48b756, {16'd2361, 16'd36740, 16'd29308, 16'd64660, 16'd38461, 16'd53540, 16'd38217, 16'd11342, 16'd56197, 16'd60921, 16'd7705, 16'd5080, 16'd38037, 16'd8830, 16'd50879, 16'd45645, 16'd26350, 16'd36085, 16'd40978, 16'd6428, 16'd43440, 16'd53210, 16'd6624, 16'd42578, 16'd53164, 16'd11296});
	test_expansion(128'h7bf8da0b7c5b3701578cf4e469708d44, {16'd53568, 16'd30993, 16'd30957, 16'd38977, 16'd15522, 16'd49490, 16'd56211, 16'd38498, 16'd40332, 16'd14109, 16'd17200, 16'd42288, 16'd3927, 16'd62559, 16'd51237, 16'd38612, 16'd10816, 16'd45006, 16'd41398, 16'd61477, 16'd43854, 16'd39062, 16'd14420, 16'd5286, 16'd16243, 16'd37075});
	test_expansion(128'hc31bae56fe7a8db3cc605ec29afe91bf, {16'd30674, 16'd47138, 16'd20094, 16'd14786, 16'd28330, 16'd51542, 16'd29362, 16'd859, 16'd17470, 16'd45235, 16'd3826, 16'd44884, 16'd6125, 16'd27453, 16'd19483, 16'd56624, 16'd7604, 16'd58388, 16'd51387, 16'd46821, 16'd29180, 16'd42739, 16'd45611, 16'd57483, 16'd27312, 16'd52263});
	test_expansion(128'hd00c23601a4969048bbef129fa616c3c, {16'd2885, 16'd4624, 16'd63083, 16'd38777, 16'd12112, 16'd53278, 16'd25100, 16'd58925, 16'd3201, 16'd12857, 16'd19647, 16'd61970, 16'd22207, 16'd53212, 16'd36550, 16'd30464, 16'd39166, 16'd22128, 16'd2519, 16'd48331, 16'd26809, 16'd55479, 16'd5257, 16'd62572, 16'd8122, 16'd37455});
	test_expansion(128'hbbbe7f42183f296c84d70e12a5e49f89, {16'd45769, 16'd64045, 16'd55726, 16'd6685, 16'd16844, 16'd12074, 16'd25146, 16'd36081, 16'd24597, 16'd9259, 16'd8844, 16'd749, 16'd60107, 16'd396, 16'd19755, 16'd23724, 16'd39184, 16'd2992, 16'd39982, 16'd14671, 16'd29314, 16'd21639, 16'd52510, 16'd49388, 16'd32753, 16'd34332});
	test_expansion(128'hc93418577f7ef51554b521935e2d7450, {16'd12624, 16'd17676, 16'd2455, 16'd218, 16'd50597, 16'd63863, 16'd35961, 16'd14236, 16'd29039, 16'd6174, 16'd54055, 16'd17678, 16'd4932, 16'd15511, 16'd38961, 16'd2976, 16'd65206, 16'd3280, 16'd57254, 16'd59658, 16'd8391, 16'd44975, 16'd60830, 16'd44147, 16'd38286, 16'd43772});
	test_expansion(128'h963c557e022f3a89f5ba31292dbc174d, {16'd31100, 16'd41581, 16'd59342, 16'd41232, 16'd46846, 16'd60817, 16'd49054, 16'd60435, 16'd56282, 16'd895, 16'd18724, 16'd55552, 16'd61989, 16'd29145, 16'd61296, 16'd36895, 16'd51523, 16'd60333, 16'd51429, 16'd24622, 16'd42429, 16'd21579, 16'd59823, 16'd33171, 16'd39349, 16'd29783});
	test_expansion(128'h0607a11fd9d0eaf3a195008e4de324b3, {16'd27541, 16'd21232, 16'd26196, 16'd4068, 16'd47506, 16'd18406, 16'd6388, 16'd12890, 16'd42150, 16'd34678, 16'd53303, 16'd6825, 16'd53383, 16'd34377, 16'd25890, 16'd3620, 16'd59589, 16'd24479, 16'd16815, 16'd6766, 16'd49704, 16'd61257, 16'd32011, 16'd7398, 16'd7749, 16'd983});
	test_expansion(128'h5b5a5054e8f81720039096ac1e3e66a5, {16'd38637, 16'd30132, 16'd30510, 16'd47020, 16'd3002, 16'd26817, 16'd32433, 16'd51480, 16'd36855, 16'd31076, 16'd33086, 16'd56084, 16'd48923, 16'd38800, 16'd55062, 16'd51624, 16'd58756, 16'd4433, 16'd45257, 16'd49940, 16'd55212, 16'd3094, 16'd52253, 16'd33354, 16'd59846, 16'd48912});
	test_expansion(128'hb06f728f99320eee1f4a42d7a4a7c84f, {16'd56040, 16'd61887, 16'd2641, 16'd32069, 16'd56765, 16'd53915, 16'd20786, 16'd3721, 16'd12519, 16'd54967, 16'd28523, 16'd60659, 16'd58506, 16'd53737, 16'd52295, 16'd43617, 16'd41412, 16'd25370, 16'd47604, 16'd12940, 16'd6472, 16'd42990, 16'd22368, 16'd30331, 16'd37341, 16'd45945});
	test_expansion(128'h3f5dafea199ebce89308289561ddb4d1, {16'd20756, 16'd27153, 16'd16574, 16'd65206, 16'd50288, 16'd1825, 16'd25730, 16'd20621, 16'd65255, 16'd45734, 16'd38945, 16'd44588, 16'd48530, 16'd10707, 16'd2507, 16'd57637, 16'd20224, 16'd54998, 16'd33421, 16'd51820, 16'd25515, 16'd46833, 16'd25146, 16'd61974, 16'd47192, 16'd62567});
	test_expansion(128'hdd7f90f076b2a912c12942789c0d0ad7, {16'd59946, 16'd9075, 16'd61434, 16'd2307, 16'd25624, 16'd33759, 16'd53988, 16'd7482, 16'd10980, 16'd49717, 16'd38214, 16'd57810, 16'd43702, 16'd47784, 16'd15415, 16'd28813, 16'd24292, 16'd8433, 16'd55530, 16'd25257, 16'd46053, 16'd19777, 16'd49373, 16'd15421, 16'd54596, 16'd57563});
	test_expansion(128'h0679929109dc3aa60b6e8556ca49b797, {16'd1827, 16'd23012, 16'd56028, 16'd9901, 16'd13955, 16'd34132, 16'd24226, 16'd47957, 16'd2991, 16'd26251, 16'd48445, 16'd9542, 16'd5257, 16'd33311, 16'd2022, 16'd21113, 16'd48630, 16'd52651, 16'd64691, 16'd61452, 16'd50461, 16'd48812, 16'd45045, 16'd59499, 16'd56513, 16'd38304});
	test_expansion(128'hcbe0b14c7ab3d9abaebd55c47a8e5884, {16'd31812, 16'd63194, 16'd62191, 16'd41626, 16'd53853, 16'd1194, 16'd53492, 16'd45552, 16'd10325, 16'd37552, 16'd26252, 16'd18755, 16'd11750, 16'd28535, 16'd54622, 16'd47136, 16'd16369, 16'd52653, 16'd36198, 16'd22991, 16'd19839, 16'd57176, 16'd44799, 16'd24938, 16'd36929, 16'd29224});
	test_expansion(128'h547dc44eb0beb8335c2d74a9fbb79655, {16'd30702, 16'd21279, 16'd2706, 16'd33056, 16'd24488, 16'd28077, 16'd54766, 16'd21905, 16'd56942, 16'd48795, 16'd14995, 16'd3243, 16'd11981, 16'd64996, 16'd31164, 16'd60759, 16'd3035, 16'd54782, 16'd34468, 16'd44287, 16'd104, 16'd42966, 16'd46294, 16'd93, 16'd38746, 16'd48424});
	test_expansion(128'ha2dc4a836b78928b793e6833f1cd795f, {16'd13115, 16'd9307, 16'd32302, 16'd40427, 16'd61, 16'd24638, 16'd47718, 16'd41937, 16'd48495, 16'd49273, 16'd24520, 16'd33800, 16'd37164, 16'd39965, 16'd45660, 16'd49083, 16'd170, 16'd13950, 16'd62883, 16'd7348, 16'd38723, 16'd40351, 16'd10388, 16'd2965, 16'd10860, 16'd56305});
	test_expansion(128'h6c31140caaaf30e3e48b789f5560da48, {16'd44020, 16'd6382, 16'd25105, 16'd11910, 16'd44717, 16'd39211, 16'd56002, 16'd10652, 16'd5842, 16'd8988, 16'd7428, 16'd21815, 16'd18919, 16'd55764, 16'd54242, 16'd42333, 16'd31019, 16'd15020, 16'd243, 16'd55405, 16'd27602, 16'd9523, 16'd23624, 16'd15064, 16'd48841, 16'd35424});
	test_expansion(128'hddfa9cffb373cc594e3fb8d96a2749cf, {16'd54679, 16'd64452, 16'd15147, 16'd49849, 16'd49856, 16'd57987, 16'd44751, 16'd43184, 16'd51399, 16'd37229, 16'd29852, 16'd33944, 16'd52134, 16'd45958, 16'd31780, 16'd37563, 16'd9583, 16'd35384, 16'd4398, 16'd25426, 16'd25678, 16'd10857, 16'd47210, 16'd15424, 16'd31204, 16'd58285});
	test_expansion(128'h4dff9921f360e4d9747f272dfff45b65, {16'd52593, 16'd50565, 16'd27499, 16'd52983, 16'd31703, 16'd15545, 16'd18440, 16'd36090, 16'd8779, 16'd56529, 16'd50466, 16'd31775, 16'd30079, 16'd50573, 16'd62590, 16'd4804, 16'd51417, 16'd26009, 16'd46008, 16'd57481, 16'd13916, 16'd33572, 16'd62251, 16'd44789, 16'd11268, 16'd64747});
	test_expansion(128'h27e83032674fbed8bbe292822bafd153, {16'd5328, 16'd17845, 16'd30810, 16'd28847, 16'd26138, 16'd52996, 16'd24917, 16'd31834, 16'd37031, 16'd14910, 16'd36611, 16'd23274, 16'd18533, 16'd11730, 16'd21924, 16'd64754, 16'd45396, 16'd50823, 16'd16615, 16'd61537, 16'd33038, 16'd29949, 16'd40278, 16'd5408, 16'd19930, 16'd37917});
	test_expansion(128'he3b48668edef873a8b1bff4222e98312, {16'd8047, 16'd45667, 16'd57001, 16'd28698, 16'd36970, 16'd35644, 16'd54612, 16'd30743, 16'd41412, 16'd23498, 16'd49932, 16'd63514, 16'd63588, 16'd47431, 16'd64106, 16'd13247, 16'd47477, 16'd58882, 16'd27298, 16'd18204, 16'd27294, 16'd40828, 16'd31826, 16'd60774, 16'd46065, 16'd48338});
	test_expansion(128'h41fc2c906ccce8a8b395ff794f472c6a, {16'd47587, 16'd4292, 16'd14947, 16'd44560, 16'd24071, 16'd8282, 16'd7982, 16'd30765, 16'd26658, 16'd23338, 16'd40278, 16'd45885, 16'd26562, 16'd6231, 16'd46983, 16'd35343, 16'd42803, 16'd16299, 16'd56488, 16'd27024, 16'd13111, 16'd32854, 16'd65316, 16'd13679, 16'd26534, 16'd62876});
	test_expansion(128'h0acdaf7b07be22192b9b20f06ca1ace8, {16'd15996, 16'd56258, 16'd53769, 16'd40375, 16'd45095, 16'd51262, 16'd12053, 16'd9254, 16'd6117, 16'd44397, 16'd39114, 16'd58513, 16'd25731, 16'd25992, 16'd42171, 16'd2656, 16'd63221, 16'd9391, 16'd51570, 16'd63322, 16'd24289, 16'd5476, 16'd1356, 16'd47005, 16'd28088, 16'd10408});
	test_expansion(128'h640086654baf363e6d3f9c2c761c87f1, {16'd36128, 16'd6699, 16'd57204, 16'd35048, 16'd36602, 16'd28723, 16'd14203, 16'd49070, 16'd27097, 16'd1886, 16'd35780, 16'd11038, 16'd30405, 16'd8627, 16'd20938, 16'd65335, 16'd38700, 16'd17885, 16'd60590, 16'd63532, 16'd61382, 16'd46950, 16'd7677, 16'd2970, 16'd15724, 16'd3684});
	test_expansion(128'h13cd48034a2b644ca0ae0cfb07184ada, {16'd59290, 16'd52314, 16'd24951, 16'd9634, 16'd2391, 16'd33550, 16'd6271, 16'd55544, 16'd34590, 16'd54128, 16'd18142, 16'd9225, 16'd52760, 16'd36706, 16'd64036, 16'd18024, 16'd33, 16'd37319, 16'd38879, 16'd50662, 16'd62795, 16'd54966, 16'd22995, 16'd30564, 16'd13508, 16'd5202});
	test_expansion(128'h955faff2fbb0e2c91df7336f993ba7e5, {16'd33619, 16'd5973, 16'd18341, 16'd58718, 16'd58690, 16'd61601, 16'd35373, 16'd62073, 16'd23861, 16'd22875, 16'd42148, 16'd209, 16'd37714, 16'd7511, 16'd15445, 16'd13828, 16'd27177, 16'd61468, 16'd60390, 16'd22186, 16'd53925, 16'd56848, 16'd20811, 16'd31813, 16'd59108, 16'd23719});
	test_expansion(128'he04eff37559d7d3ae6985ecf7af3c60a, {16'd61459, 16'd53312, 16'd62755, 16'd31024, 16'd62134, 16'd29278, 16'd52501, 16'd14010, 16'd46206, 16'd16178, 16'd7290, 16'd20763, 16'd12497, 16'd3526, 16'd62526, 16'd41989, 16'd55866, 16'd35925, 16'd47024, 16'd8797, 16'd53170, 16'd12524, 16'd12004, 16'd14468, 16'd13819, 16'd32186});
	test_expansion(128'hde66916e0b0ea26dc44d4b0a93eb289d, {16'd41853, 16'd22195, 16'd38041, 16'd11104, 16'd53384, 16'd19729, 16'd65272, 16'd59062, 16'd38235, 16'd45634, 16'd17272, 16'd63523, 16'd8487, 16'd23613, 16'd56724, 16'd59183, 16'd63215, 16'd7277, 16'd32542, 16'd63214, 16'd25959, 16'd8541, 16'd23622, 16'd55931, 16'd13345, 16'd58786});
	test_expansion(128'h92cb896a8c6122337d290a64e20abe34, {16'd36046, 16'd48571, 16'd14730, 16'd57974, 16'd16164, 16'd21627, 16'd37287, 16'd64619, 16'd37964, 16'd12661, 16'd52348, 16'd36399, 16'd9349, 16'd48933, 16'd49176, 16'd15673, 16'd23365, 16'd56473, 16'd61935, 16'd55749, 16'd27814, 16'd27913, 16'd2474, 16'd38620, 16'd3138, 16'd18048});
	test_expansion(128'h7e515f5ba194782df513ae1bee938485, {16'd48536, 16'd43260, 16'd64231, 16'd38315, 16'd16664, 16'd18665, 16'd31388, 16'd55304, 16'd20483, 16'd35371, 16'd7014, 16'd5710, 16'd23591, 16'd17672, 16'd58672, 16'd56292, 16'd60059, 16'd50983, 16'd30702, 16'd35622, 16'd24843, 16'd19114, 16'd1261, 16'd15297, 16'd34253, 16'd51930});
	test_expansion(128'h5c643b5974067c79170089a800521aee, {16'd34601, 16'd38848, 16'd40849, 16'd60023, 16'd31015, 16'd13395, 16'd16628, 16'd38847, 16'd3922, 16'd6979, 16'd62983, 16'd27851, 16'd27372, 16'd49029, 16'd60073, 16'd27449, 16'd57158, 16'd6260, 16'd22287, 16'd49817, 16'd24506, 16'd54794, 16'd63164, 16'd51223, 16'd51814, 16'd26332});
	test_expansion(128'hd5e462b1d3047a68702285b00216df90, {16'd19370, 16'd47210, 16'd25950, 16'd37263, 16'd19452, 16'd43021, 16'd63009, 16'd15671, 16'd47137, 16'd20300, 16'd47149, 16'd38653, 16'd6960, 16'd30803, 16'd64223, 16'd47199, 16'd36351, 16'd32313, 16'd20812, 16'd7152, 16'd25898, 16'd4811, 16'd19190, 16'd12403, 16'd35844, 16'd60284});
	test_expansion(128'h286c6fbb4cb2ef7b1442aa101636db7f, {16'd40052, 16'd38797, 16'd37085, 16'd16631, 16'd49361, 16'd34469, 16'd40373, 16'd18530, 16'd65477, 16'd65514, 16'd22447, 16'd42408, 16'd46685, 16'd31135, 16'd62033, 16'd18500, 16'd57442, 16'd54631, 16'd5265, 16'd23805, 16'd36656, 16'd17610, 16'd15715, 16'd26046, 16'd42827, 16'd36940});
	test_expansion(128'h337e3063f937d493a08a49622524757e, {16'd20891, 16'd5353, 16'd52454, 16'd32523, 16'd25304, 16'd58636, 16'd55904, 16'd53840, 16'd30556, 16'd51972, 16'd7255, 16'd36251, 16'd24519, 16'd27114, 16'd25890, 16'd63667, 16'd26772, 16'd26288, 16'd7409, 16'd21397, 16'd7884, 16'd49366, 16'd1416, 16'd23591, 16'd46970, 16'd64722});
	test_expansion(128'he0299c16ebcc5d6854901bc65c45fcbe, {16'd38890, 16'd56454, 16'd2862, 16'd20167, 16'd34105, 16'd16723, 16'd5160, 16'd25777, 16'd30370, 16'd41511, 16'd26346, 16'd31119, 16'd10860, 16'd41227, 16'd23531, 16'd53164, 16'd1774, 16'd12352, 16'd6819, 16'd59278, 16'd39593, 16'd905, 16'd6361, 16'd55727, 16'd20682, 16'd46122});
	test_expansion(128'h6c71aa74457b794ef8c48c17f452f505, {16'd20391, 16'd50949, 16'd15538, 16'd38363, 16'd7220, 16'd18676, 16'd59692, 16'd43579, 16'd2287, 16'd2540, 16'd36181, 16'd58814, 16'd49764, 16'd15241, 16'd16972, 16'd608, 16'd63318, 16'd23874, 16'd36026, 16'd6439, 16'd55177, 16'd9903, 16'd36339, 16'd18930, 16'd21385, 16'd54635});
	test_expansion(128'h0e0ebdcfaaac487f99c2d86b78b9ca1f, {16'd458, 16'd29910, 16'd56552, 16'd45851, 16'd19088, 16'd15019, 16'd39302, 16'd36086, 16'd5421, 16'd13643, 16'd52879, 16'd47637, 16'd21907, 16'd58610, 16'd11866, 16'd20058, 16'd20475, 16'd62666, 16'd37572, 16'd34239, 16'd36697, 16'd16162, 16'd1347, 16'd64571, 16'd55828, 16'd24899});
	test_expansion(128'hbb406c67c45e7da24a94942d18e05eb4, {16'd39635, 16'd38438, 16'd19322, 16'd33188, 16'd37100, 16'd52399, 16'd15794, 16'd19137, 16'd37957, 16'd25000, 16'd62175, 16'd9328, 16'd27961, 16'd13974, 16'd3422, 16'd21427, 16'd27462, 16'd55409, 16'd58877, 16'd13858, 16'd46829, 16'd56862, 16'd20389, 16'd5167, 16'd61589, 16'd51421});
	test_expansion(128'hc65205090b465941647baba8f4a66536, {16'd55995, 16'd28, 16'd32885, 16'd1797, 16'd6235, 16'd26999, 16'd6585, 16'd8698, 16'd12087, 16'd18813, 16'd17711, 16'd63560, 16'd58601, 16'd3163, 16'd54195, 16'd61500, 16'd35816, 16'd50402, 16'd1307, 16'd53903, 16'd41186, 16'd43439, 16'd36656, 16'd60771, 16'd1972, 16'd13359});
	test_expansion(128'h9cf5abe180fe8046b146316a89317486, {16'd49487, 16'd27749, 16'd17540, 16'd46411, 16'd42903, 16'd33452, 16'd16666, 16'd62929, 16'd35842, 16'd25283, 16'd8147, 16'd62674, 16'd278, 16'd17625, 16'd10861, 16'd58840, 16'd50583, 16'd38961, 16'd48174, 16'd48614, 16'd60823, 16'd52546, 16'd14307, 16'd41779, 16'd32326, 16'd20531});
	test_expansion(128'h2f5dca0c3cdc2968e6e4ad1145083b73, {16'd37964, 16'd49005, 16'd46077, 16'd57322, 16'd37696, 16'd10487, 16'd41943, 16'd64654, 16'd1842, 16'd10092, 16'd63990, 16'd44543, 16'd17864, 16'd8940, 16'd15395, 16'd5263, 16'd6536, 16'd7238, 16'd20807, 16'd21505, 16'd55791, 16'd29646, 16'd21022, 16'd41095, 16'd56771, 16'd41477});
	test_expansion(128'h98a69d5cb3e3be1c98cae6bc89f2a8e3, {16'd2201, 16'd1731, 16'd55438, 16'd2713, 16'd41537, 16'd17310, 16'd42365, 16'd57868, 16'd23445, 16'd48018, 16'd291, 16'd50995, 16'd38588, 16'd45532, 16'd47955, 16'd494, 16'd61810, 16'd37947, 16'd59626, 16'd17787, 16'd26908, 16'd9498, 16'd33521, 16'd41405, 16'd20886, 16'd49341});
	test_expansion(128'h330a6fd2e3efdedcce01e80067443a23, {16'd37369, 16'd33266, 16'd38950, 16'd36949, 16'd50025, 16'd5551, 16'd56845, 16'd27160, 16'd30749, 16'd15187, 16'd7145, 16'd16916, 16'd34242, 16'd16478, 16'd58723, 16'd2118, 16'd37620, 16'd14735, 16'd19401, 16'd42079, 16'd23894, 16'd62450, 16'd16679, 16'd40380, 16'd50393, 16'd768});
	test_expansion(128'h20f4f3f2ef14d31db431a313433624da, {16'd36265, 16'd17773, 16'd50849, 16'd63030, 16'd46344, 16'd25815, 16'd59431, 16'd56286, 16'd27227, 16'd65532, 16'd61203, 16'd32791, 16'd2857, 16'd46925, 16'd59043, 16'd64889, 16'd12010, 16'd63982, 16'd2225, 16'd34213, 16'd44923, 16'd24398, 16'd18310, 16'd56161, 16'd56212, 16'd28464});
	test_expansion(128'h9a54ec9056842997b09745c7d4b58232, {16'd32804, 16'd33602, 16'd22835, 16'd41681, 16'd41877, 16'd26504, 16'd19661, 16'd23402, 16'd20365, 16'd47549, 16'd37440, 16'd12132, 16'd41266, 16'd55430, 16'd33338, 16'd31621, 16'd51008, 16'd45909, 16'd47135, 16'd22474, 16'd18723, 16'd41046, 16'd24265, 16'd18754, 16'd10841, 16'd4784});
	test_expansion(128'h7f9c44d36180525f576198bf831d3799, {16'd734, 16'd301, 16'd58153, 16'd6846, 16'd60562, 16'd43962, 16'd46649, 16'd35641, 16'd37531, 16'd65464, 16'd62503, 16'd350, 16'd49402, 16'd44859, 16'd45785, 16'd24260, 16'd1276, 16'd11333, 16'd58292, 16'd20789, 16'd23090, 16'd55072, 16'd8469, 16'd5199, 16'd15571, 16'd64848});
	test_expansion(128'h55738250c05c90f66c16198d453c4741, {16'd35004, 16'd55112, 16'd31580, 16'd59368, 16'd33740, 16'd4460, 16'd36350, 16'd13298, 16'd26024, 16'd64949, 16'd7752, 16'd15264, 16'd20972, 16'd37086, 16'd47938, 16'd18430, 16'd10324, 16'd48640, 16'd58374, 16'd45871, 16'd60792, 16'd5203, 16'd890, 16'd30381, 16'd11450, 16'd28386});
	test_expansion(128'h3f1dd6978942c713a528d3619688fe39, {16'd57019, 16'd31469, 16'd34486, 16'd27112, 16'd21678, 16'd25750, 16'd34555, 16'd16216, 16'd43273, 16'd59958, 16'd60363, 16'd56551, 16'd26320, 16'd10309, 16'd45755, 16'd65006, 16'd32437, 16'd12532, 16'd30766, 16'd15566, 16'd32238, 16'd24704, 16'd33229, 16'd45854, 16'd56420, 16'd52525});
	test_expansion(128'h712d937850ce51d6c1251492bf2686f4, {16'd63846, 16'd16869, 16'd45785, 16'd8305, 16'd42462, 16'd23265, 16'd17991, 16'd284, 16'd41001, 16'd39366, 16'd10862, 16'd17198, 16'd3270, 16'd34774, 16'd62989, 16'd19329, 16'd11766, 16'd61726, 16'd24530, 16'd56707, 16'd60437, 16'd35330, 16'd27060, 16'd17357, 16'd50425, 16'd19184});
	test_expansion(128'h1a05a82feb47fe15b61451df4db73f02, {16'd32119, 16'd59199, 16'd52846, 16'd29865, 16'd21985, 16'd50014, 16'd26920, 16'd50177, 16'd37362, 16'd19554, 16'd40150, 16'd7546, 16'd29647, 16'd18811, 16'd31392, 16'd18139, 16'd54816, 16'd58160, 16'd37973, 16'd54735, 16'd6410, 16'd24738, 16'd32189, 16'd15621, 16'd17504, 16'd32917});
	test_expansion(128'h311061ef516f1c447d7dda62ae866053, {16'd25131, 16'd13795, 16'd24611, 16'd6218, 16'd60586, 16'd25299, 16'd61721, 16'd63049, 16'd47576, 16'd37166, 16'd57013, 16'd50859, 16'd24010, 16'd37066, 16'd36132, 16'd32503, 16'd27407, 16'd8459, 16'd3846, 16'd46895, 16'd43885, 16'd42516, 16'd25334, 16'd55936, 16'd2158, 16'd11477});
	test_expansion(128'hbb2f610650f6ac01b639c55be52c5b92, {16'd12779, 16'd6104, 16'd23231, 16'd26916, 16'd53794, 16'd59689, 16'd51129, 16'd50869, 16'd8233, 16'd49997, 16'd21855, 16'd1215, 16'd38140, 16'd41391, 16'd61962, 16'd12451, 16'd36901, 16'd17286, 16'd893, 16'd35489, 16'd49075, 16'd40303, 16'd43975, 16'd25309, 16'd61654, 16'd27248});
	test_expansion(128'h4b949333b5429ec2d17da4f4e9593090, {16'd17481, 16'd29017, 16'd14532, 16'd23600, 16'd19531, 16'd37695, 16'd33915, 16'd39940, 16'd30331, 16'd62147, 16'd14812, 16'd51263, 16'd25521, 16'd37079, 16'd11004, 16'd51747, 16'd33513, 16'd57452, 16'd6460, 16'd61193, 16'd10036, 16'd24337, 16'd5197, 16'd18925, 16'd29843, 16'd25413});
	test_expansion(128'hdc07b0f138eff16dd056d15841eb7667, {16'd42298, 16'd14863, 16'd17483, 16'd32866, 16'd32880, 16'd4051, 16'd14731, 16'd55551, 16'd54070, 16'd49872, 16'd26605, 16'd36158, 16'd34893, 16'd32786, 16'd14486, 16'd8159, 16'd44822, 16'd10172, 16'd63750, 16'd7777, 16'd54964, 16'd39177, 16'd46894, 16'd22556, 16'd18209, 16'd24134});
	test_expansion(128'h6d864cdf5fd98ee06283e78fa4ec4439, {16'd49410, 16'd64750, 16'd24324, 16'd18725, 16'd50284, 16'd57277, 16'd17804, 16'd38102, 16'd57726, 16'd7302, 16'd30821, 16'd61457, 16'd39209, 16'd38143, 16'd54646, 16'd2123, 16'd37669, 16'd12246, 16'd24369, 16'd27949, 16'd18134, 16'd6255, 16'd21167, 16'd2659, 16'd18102, 16'd11931});
	test_expansion(128'hf8d25f437d96774ccce9fca8e64d4eef, {16'd64617, 16'd35011, 16'd6612, 16'd44928, 16'd26529, 16'd35223, 16'd37754, 16'd8070, 16'd61320, 16'd19654, 16'd11362, 16'd37675, 16'd39015, 16'd38394, 16'd5505, 16'd36303, 16'd50573, 16'd59629, 16'd43293, 16'd8562, 16'd62530, 16'd57357, 16'd7714, 16'd18696, 16'd40052, 16'd13376});
	test_expansion(128'h1ca3f2a38fa848e64d2723db44416851, {16'd34700, 16'd2548, 16'd35648, 16'd38207, 16'd25797, 16'd12017, 16'd34096, 16'd30071, 16'd60655, 16'd32364, 16'd1003, 16'd46329, 16'd1520, 16'd21877, 16'd39543, 16'd48442, 16'd36922, 16'd53824, 16'd58992, 16'd15934, 16'd45370, 16'd46783, 16'd50129, 16'd54705, 16'd29949, 16'd14316});
	test_expansion(128'h64c7f1a384845b45537e883b651c162a, {16'd18169, 16'd51981, 16'd20661, 16'd54954, 16'd7150, 16'd38017, 16'd31587, 16'd62067, 16'd34809, 16'd26318, 16'd5404, 16'd57747, 16'd3778, 16'd55127, 16'd60335, 16'd43398, 16'd59003, 16'd34149, 16'd25316, 16'd7218, 16'd31241, 16'd14601, 16'd40383, 16'd57433, 16'd3719, 16'd48944});
	test_expansion(128'hd791dd06d2c71b5c351f216ffb4743e0, {16'd57320, 16'd51874, 16'd53121, 16'd10655, 16'd13929, 16'd28413, 16'd13664, 16'd19024, 16'd47808, 16'd33770, 16'd8984, 16'd50300, 16'd33218, 16'd35999, 16'd3414, 16'd53458, 16'd44045, 16'd26658, 16'd846, 16'd58486, 16'd62828, 16'd16741, 16'd45151, 16'd12315, 16'd27137, 16'd24391});
	test_expansion(128'hc99f914597c7adcbdb93deea3cb742f7, {16'd45716, 16'd4839, 16'd36924, 16'd11334, 16'd4727, 16'd32699, 16'd28244, 16'd53627, 16'd49751, 16'd18132, 16'd32896, 16'd24334, 16'd895, 16'd2702, 16'd64812, 16'd51935, 16'd31650, 16'd54902, 16'd18202, 16'd22977, 16'd46126, 16'd20373, 16'd51240, 16'd58789, 16'd61871, 16'd36910});
	test_expansion(128'h5f259521e42cedfbd2380d587e8e5784, {16'd35898, 16'd5340, 16'd63431, 16'd26281, 16'd30297, 16'd10960, 16'd60094, 16'd8024, 16'd41344, 16'd46278, 16'd55870, 16'd14572, 16'd34003, 16'd47111, 16'd62, 16'd29897, 16'd13027, 16'd27729, 16'd4429, 16'd16565, 16'd38463, 16'd53474, 16'd20008, 16'd11087, 16'd17235, 16'd9579});
	test_expansion(128'h442e5d7fc71339f0d743cf950d62a58f, {16'd34492, 16'd925, 16'd5678, 16'd58851, 16'd3730, 16'd19859, 16'd49182, 16'd50508, 16'd14928, 16'd54669, 16'd22425, 16'd49442, 16'd23332, 16'd17447, 16'd469, 16'd59794, 16'd33384, 16'd18335, 16'd16580, 16'd59574, 16'd7185, 16'd49088, 16'd65404, 16'd847, 16'd12232, 16'd29410});
	test_expansion(128'heb1b42885cfa0b144e029e1e6a4fb1c1, {16'd28889, 16'd5928, 16'd59599, 16'd39009, 16'd31233, 16'd6081, 16'd1944, 16'd1416, 16'd21602, 16'd49916, 16'd7558, 16'd55826, 16'd41721, 16'd48323, 16'd26933, 16'd9165, 16'd3303, 16'd22680, 16'd43461, 16'd53723, 16'd26342, 16'd31308, 16'd11737, 16'd29474, 16'd18861, 16'd13949});
	test_expansion(128'h15d7ee289f1727c240ce5cac1d673806, {16'd45872, 16'd40222, 16'd51274, 16'd31506, 16'd62040, 16'd14122, 16'd11989, 16'd60627, 16'd5452, 16'd58545, 16'd36448, 16'd43689, 16'd61642, 16'd41415, 16'd48515, 16'd13714, 16'd30628, 16'd15818, 16'd36950, 16'd61052, 16'd39638, 16'd37630, 16'd11880, 16'd40031, 16'd792, 16'd15527});
	test_expansion(128'h725a05585699b8edaf07c2a9b1b4ae8b, {16'd62558, 16'd1905, 16'd31424, 16'd24430, 16'd21236, 16'd63598, 16'd8810, 16'd44613, 16'd12794, 16'd39353, 16'd30172, 16'd56484, 16'd19270, 16'd2715, 16'd50805, 16'd37311, 16'd40968, 16'd21942, 16'd25975, 16'd44898, 16'd12580, 16'd3933, 16'd16860, 16'd11751, 16'd17167, 16'd13808});
	test_expansion(128'hc7e5750fe40f06ab41dd0279b1a4b78d, {16'd34052, 16'd62506, 16'd42756, 16'd30709, 16'd1395, 16'd60936, 16'd29576, 16'd2635, 16'd48588, 16'd18445, 16'd1153, 16'd12003, 16'd54755, 16'd59685, 16'd41866, 16'd53725, 16'd15357, 16'd27652, 16'd42464, 16'd48821, 16'd3732, 16'd20631, 16'd26423, 16'd351, 16'd15467, 16'd2684});
	test_expansion(128'h33946f1fad17ceec527d6b2406174b65, {16'd65326, 16'd61810, 16'd38371, 16'd5665, 16'd56355, 16'd27041, 16'd55777, 16'd30965, 16'd54684, 16'd45057, 16'd8472, 16'd4311, 16'd1795, 16'd4391, 16'd44381, 16'd60823, 16'd61322, 16'd42872, 16'd7662, 16'd36915, 16'd35708, 16'd12613, 16'd34346, 16'd63529, 16'd21415, 16'd16609});
	test_expansion(128'h730c97d0d9fe1487621058332c1f6114, {16'd8427, 16'd17129, 16'd48852, 16'd34281, 16'd15516, 16'd21453, 16'd3290, 16'd34042, 16'd51428, 16'd45900, 16'd27236, 16'd50823, 16'd48076, 16'd45256, 16'd60251, 16'd60589, 16'd56555, 16'd63802, 16'd11351, 16'd47273, 16'd58524, 16'd3466, 16'd65126, 16'd4424, 16'd29625, 16'd64813});
	test_expansion(128'hf134077ede97ac1e296758278ca987c7, {16'd21207, 16'd18166, 16'd41309, 16'd53105, 16'd24083, 16'd55119, 16'd57664, 16'd55133, 16'd24996, 16'd48324, 16'd31922, 16'd42500, 16'd17989, 16'd11880, 16'd16510, 16'd28362, 16'd53541, 16'd60674, 16'd12731, 16'd8899, 16'd17509, 16'd51240, 16'd57501, 16'd16201, 16'd16314, 16'd38759});
	test_expansion(128'h671d0d3f0d1142ae9747ad4bc4926657, {16'd7413, 16'd11305, 16'd9638, 16'd40771, 16'd13007, 16'd35034, 16'd10573, 16'd37567, 16'd222, 16'd26662, 16'd10536, 16'd5278, 16'd58173, 16'd20099, 16'd32748, 16'd3051, 16'd59399, 16'd34458, 16'd6197, 16'd9554, 16'd14659, 16'd25374, 16'd42401, 16'd52237, 16'd30530, 16'd46049});
	test_expansion(128'h8020fef896a7fd6c37f64ef93e42e3b8, {16'd28408, 16'd43083, 16'd14268, 16'd20735, 16'd23980, 16'd54125, 16'd26143, 16'd54481, 16'd18643, 16'd62828, 16'd55901, 16'd38245, 16'd9204, 16'd64561, 16'd29863, 16'd3114, 16'd2136, 16'd51160, 16'd42395, 16'd56367, 16'd52006, 16'd46610, 16'd22379, 16'd41739, 16'd12336, 16'd14897});
	test_expansion(128'h15fb55280f5839424515df5a73159a3a, {16'd17610, 16'd6331, 16'd58845, 16'd50103, 16'd2831, 16'd31459, 16'd55512, 16'd34985, 16'd2427, 16'd41647, 16'd62212, 16'd32446, 16'd16873, 16'd43006, 16'd7938, 16'd7574, 16'd5435, 16'd51662, 16'd27438, 16'd9632, 16'd64624, 16'd7123, 16'd22986, 16'd31156, 16'd50404, 16'd297});
	test_expansion(128'h1e760f0290db5a7d5851f9e911a90ecd, {16'd1856, 16'd8606, 16'd46314, 16'd11909, 16'd13568, 16'd8493, 16'd31516, 16'd19653, 16'd51554, 16'd33301, 16'd59701, 16'd29483, 16'd19173, 16'd61709, 16'd36771, 16'd63064, 16'd58780, 16'd1258, 16'd46776, 16'd38055, 16'd60178, 16'd60933, 16'd34000, 16'd63130, 16'd55361, 16'd49539});
	test_expansion(128'h61b103ec333776447557cc3b9d586faa, {16'd47503, 16'd48367, 16'd62367, 16'd45115, 16'd55890, 16'd39389, 16'd29295, 16'd975, 16'd30336, 16'd9840, 16'd53952, 16'd62539, 16'd5135, 16'd14648, 16'd18143, 16'd39533, 16'd21770, 16'd58961, 16'd62130, 16'd2702, 16'd5182, 16'd9926, 16'd10120, 16'd51163, 16'd65488, 16'd6051});
	test_expansion(128'h07e63203773d5206480a76653469ac35, {16'd25464, 16'd33574, 16'd52582, 16'd206, 16'd2039, 16'd64215, 16'd22568, 16'd15785, 16'd26957, 16'd53322, 16'd31161, 16'd31455, 16'd7332, 16'd13255, 16'd8258, 16'd20327, 16'd40924, 16'd37149, 16'd35009, 16'd45011, 16'd24835, 16'd13326, 16'd5788, 16'd40600, 16'd37616, 16'd18421});
	test_expansion(128'h7b45c9a70d42ca08fa7aa1c6399c0e5e, {16'd34215, 16'd58580, 16'd49497, 16'd3449, 16'd41209, 16'd1418, 16'd17818, 16'd42275, 16'd18762, 16'd29631, 16'd61744, 16'd28697, 16'd48771, 16'd8591, 16'd33227, 16'd41834, 16'd35705, 16'd57143, 16'd1743, 16'd41700, 16'd10315, 16'd43699, 16'd64759, 16'd1139, 16'd35292, 16'd6163});
	test_expansion(128'hebe7accea64cb24393f08e90397c15a9, {16'd32898, 16'd24266, 16'd49076, 16'd966, 16'd34642, 16'd62456, 16'd63596, 16'd3028, 16'd46480, 16'd22926, 16'd38704, 16'd51377, 16'd7906, 16'd64963, 16'd49243, 16'd12858, 16'd4266, 16'd1563, 16'd12797, 16'd59015, 16'd49110, 16'd31124, 16'd38708, 16'd64607, 16'd53306, 16'd50621});
	test_expansion(128'h2c8ed00113d86bc8d517b3574b991829, {16'd60587, 16'd5164, 16'd23786, 16'd21474, 16'd47571, 16'd56034, 16'd42979, 16'd13481, 16'd9393, 16'd65084, 16'd43436, 16'd11263, 16'd25271, 16'd62453, 16'd29187, 16'd22456, 16'd51042, 16'd6060, 16'd60384, 16'd1916, 16'd47943, 16'd54021, 16'd50211, 16'd14363, 16'd19361, 16'd27203});
	test_expansion(128'h32e0f792a49425ea981fbfb175a2e2f0, {16'd33035, 16'd36421, 16'd63340, 16'd38420, 16'd32389, 16'd26644, 16'd65336, 16'd15380, 16'd23923, 16'd36759, 16'd30287, 16'd24933, 16'd5743, 16'd30825, 16'd8719, 16'd43384, 16'd65031, 16'd4273, 16'd21127, 16'd46183, 16'd62415, 16'd24168, 16'd53691, 16'd23536, 16'd36987, 16'd24353});
	test_expansion(128'h163547397b3fc12d554096606e648459, {16'd56880, 16'd64800, 16'd46355, 16'd35180, 16'd22370, 16'd44495, 16'd42540, 16'd19051, 16'd30496, 16'd61194, 16'd50465, 16'd47298, 16'd16282, 16'd46193, 16'd57584, 16'd63558, 16'd16635, 16'd32375, 16'd7783, 16'd60052, 16'd2333, 16'd32877, 16'd22172, 16'd50965, 16'd36200, 16'd62370});
	test_expansion(128'hdd80622c68730e21a17bf35f428e34dd, {16'd21253, 16'd59796, 16'd44847, 16'd54717, 16'd7742, 16'd28390, 16'd62499, 16'd12852, 16'd56168, 16'd20777, 16'd6846, 16'd61077, 16'd60960, 16'd45618, 16'd10595, 16'd40799, 16'd14643, 16'd55915, 16'd18167, 16'd16175, 16'd37387, 16'd39020, 16'd12021, 16'd26848, 16'd9930, 16'd61593});
	test_expansion(128'h6e779c6f1cd8871c978d4700ab3be029, {16'd49963, 16'd45328, 16'd12608, 16'd42222, 16'd43568, 16'd41024, 16'd24027, 16'd11258, 16'd53937, 16'd63226, 16'd10464, 16'd61538, 16'd4879, 16'd7849, 16'd55159, 16'd60620, 16'd33503, 16'd13077, 16'd49322, 16'd10994, 16'd60581, 16'd41821, 16'd2027, 16'd6127, 16'd19673, 16'd34367});
	test_expansion(128'hbc6eb1324bd08a4cf55e26cdb9f8dfb8, {16'd61810, 16'd21553, 16'd36548, 16'd17214, 16'd57577, 16'd4152, 16'd33267, 16'd9353, 16'd56489, 16'd36773, 16'd11381, 16'd59289, 16'd8410, 16'd313, 16'd26977, 16'd32255, 16'd39551, 16'd55714, 16'd35962, 16'd26389, 16'd61131, 16'd6102, 16'd57212, 16'd35059, 16'd50872, 16'd2445});
	test_expansion(128'h8506f56091aac79e544d852b18f32687, {16'd31882, 16'd11609, 16'd19650, 16'd25698, 16'd41897, 16'd832, 16'd27577, 16'd8035, 16'd57085, 16'd10177, 16'd52291, 16'd38151, 16'd24171, 16'd41228, 16'd28324, 16'd9884, 16'd40291, 16'd12871, 16'd832, 16'd53115, 16'd27945, 16'd34008, 16'd6307, 16'd41104, 16'd58120, 16'd20177});
	test_expansion(128'h6847fdc7b77c3b23163e73abf611bc02, {16'd29304, 16'd43046, 16'd52739, 16'd52673, 16'd52293, 16'd52428, 16'd109, 16'd10905, 16'd4355, 16'd57444, 16'd54516, 16'd30497, 16'd28250, 16'd57721, 16'd57415, 16'd14352, 16'd54519, 16'd45093, 16'd12791, 16'd22018, 16'd23118, 16'd17394, 16'd9306, 16'd38029, 16'd51256, 16'd28207});
	test_expansion(128'h7c6d501b714735a98da14666f1f130c2, {16'd52702, 16'd48133, 16'd57753, 16'd16261, 16'd48285, 16'd27452, 16'd28697, 16'd51386, 16'd36174, 16'd25655, 16'd31293, 16'd10984, 16'd28310, 16'd53453, 16'd55280, 16'd41076, 16'd11587, 16'd16342, 16'd23754, 16'd26506, 16'd13892, 16'd16399, 16'd4399, 16'd49894, 16'd54133, 16'd59165});
	test_expansion(128'h8d63c455e0b3ff3e3e70a817c4f2af2e, {16'd51139, 16'd63569, 16'd13673, 16'd11805, 16'd30088, 16'd19479, 16'd25901, 16'd32327, 16'd58592, 16'd6388, 16'd40725, 16'd8746, 16'd31911, 16'd1966, 16'd10203, 16'd60145, 16'd38598, 16'd54509, 16'd47576, 16'd39522, 16'd65258, 16'd23454, 16'd3155, 16'd25996, 16'd7249, 16'd43480});
	test_expansion(128'hcdaa295586d4798fe8e8d8770f0871cc, {16'd535, 16'd53167, 16'd3716, 16'd26548, 16'd14741, 16'd38157, 16'd7090, 16'd7346, 16'd3086, 16'd48031, 16'd56175, 16'd5007, 16'd15234, 16'd23680, 16'd330, 16'd21614, 16'd55911, 16'd23133, 16'd37415, 16'd8731, 16'd29193, 16'd56164, 16'd47836, 16'd45447, 16'd32360, 16'd21540});
	test_expansion(128'hc8d47e691d545db99c192cb536cf55f7, {16'd1004, 16'd42708, 16'd27564, 16'd64138, 16'd3865, 16'd19888, 16'd1527, 16'd49360, 16'd38392, 16'd1051, 16'd35174, 16'd33248, 16'd21815, 16'd43209, 16'd25852, 16'd57771, 16'd39891, 16'd2441, 16'd9252, 16'd12066, 16'd53221, 16'd59146, 16'd50923, 16'd42746, 16'd46252, 16'd8886});
	test_expansion(128'h0a48625ba6cbcd671becb32540633d2a, {16'd46777, 16'd16076, 16'd14105, 16'd45188, 16'd13460, 16'd61257, 16'd21605, 16'd55617, 16'd3079, 16'd25223, 16'd35201, 16'd41485, 16'd41825, 16'd63475, 16'd34440, 16'd14239, 16'd40989, 16'd50846, 16'd35651, 16'd26987, 16'd1692, 16'd21849, 16'd64124, 16'd5522, 16'd33720, 16'd56780});
	test_expansion(128'h71fba84fa601be6739305475c6f221de, {16'd21871, 16'd60830, 16'd64413, 16'd9099, 16'd18268, 16'd50640, 16'd52452, 16'd59141, 16'd33585, 16'd16613, 16'd10576, 16'd15556, 16'd56051, 16'd7591, 16'd7689, 16'd19888, 16'd44863, 16'd33121, 16'd35718, 16'd13188, 16'd20759, 16'd14221, 16'd10315, 16'd25629, 16'd24309, 16'd30068});
	test_expansion(128'hc3e754bd497e8f2f8b442ae77b29f9af, {16'd26855, 16'd12997, 16'd37580, 16'd26364, 16'd26692, 16'd3969, 16'd2328, 16'd47151, 16'd26221, 16'd26846, 16'd15326, 16'd21489, 16'd11714, 16'd47014, 16'd64469, 16'd39520, 16'd42147, 16'd11192, 16'd59594, 16'd40224, 16'd22481, 16'd10624, 16'd24799, 16'd53480, 16'd36156, 16'd55966});
	test_expansion(128'hb2789c3f48fd53831233a38df3ef14ec, {16'd33621, 16'd52962, 16'd49638, 16'd3574, 16'd39224, 16'd59170, 16'd24645, 16'd34163, 16'd54505, 16'd36044, 16'd20399, 16'd25263, 16'd52333, 16'd7185, 16'd22745, 16'd54409, 16'd36392, 16'd58167, 16'd22582, 16'd29912, 16'd40836, 16'd4064, 16'd33323, 16'd64938, 16'd48382, 16'd57938});
	test_expansion(128'h499761f4291a7af381ea58ea7e79ec8d, {16'd37080, 16'd28956, 16'd3344, 16'd56283, 16'd60980, 16'd849, 16'd52047, 16'd12958, 16'd16724, 16'd24985, 16'd26793, 16'd46053, 16'd19059, 16'd7350, 16'd64570, 16'd50696, 16'd33486, 16'd4740, 16'd60148, 16'd49834, 16'd20234, 16'd2375, 16'd3209, 16'd9182, 16'd38832, 16'd51227});
	test_expansion(128'h0dc31d76f85d7e729fcf3c1314661ea3, {16'd52270, 16'd52931, 16'd41540, 16'd59297, 16'd64161, 16'd62488, 16'd59345, 16'd17013, 16'd23910, 16'd63422, 16'd48025, 16'd20040, 16'd63010, 16'd28350, 16'd1720, 16'd24778, 16'd56598, 16'd31559, 16'd51594, 16'd37864, 16'd60242, 16'd61982, 16'd37615, 16'd32561, 16'd40572, 16'd64756});
	test_expansion(128'h3c7af9986cefc0dcc53f788a7ec3e734, {16'd1615, 16'd3016, 16'd63511, 16'd55818, 16'd25079, 16'd8486, 16'd25801, 16'd39535, 16'd62322, 16'd21068, 16'd63101, 16'd39836, 16'd4948, 16'd49581, 16'd23162, 16'd22579, 16'd44132, 16'd55188, 16'd56190, 16'd56349, 16'd32305, 16'd53180, 16'd34589, 16'd48869, 16'd7139, 16'd41211});
	test_expansion(128'h0405e373183ce9bbc6bc8fcfdc1f821a, {16'd55716, 16'd21084, 16'd4700, 16'd34620, 16'd24981, 16'd39674, 16'd5200, 16'd55573, 16'd37457, 16'd26100, 16'd12331, 16'd60956, 16'd30556, 16'd16344, 16'd24106, 16'd4875, 16'd65070, 16'd40060, 16'd25843, 16'd32827, 16'd57481, 16'd20990, 16'd40566, 16'd39827, 16'd57541, 16'd25318});
	test_expansion(128'hd5fb2cb332b055a8e06c221503ece592, {16'd21649, 16'd55813, 16'd257, 16'd62769, 16'd30339, 16'd12061, 16'd31481, 16'd4784, 16'd17019, 16'd57654, 16'd46080, 16'd49761, 16'd63994, 16'd20419, 16'd1940, 16'd5514, 16'd1739, 16'd1906, 16'd38052, 16'd54896, 16'd39235, 16'd23479, 16'd23371, 16'd44008, 16'd19345, 16'd1306});
	test_expansion(128'hc804ff20e977cff1b97e9556c0cddd8a, {16'd21726, 16'd10295, 16'd59617, 16'd48326, 16'd59721, 16'd25780, 16'd18060, 16'd51771, 16'd21649, 16'd63174, 16'd13889, 16'd45366, 16'd40272, 16'd53543, 16'd981, 16'd267, 16'd7884, 16'd26957, 16'd43611, 16'd24319, 16'd4970, 16'd51440, 16'd36735, 16'd15654, 16'd10355, 16'd40590});
	test_expansion(128'h7075451d3ca4d23fe0e5470e9d75bc5a, {16'd38886, 16'd25556, 16'd13704, 16'd15224, 16'd45565, 16'd29376, 16'd47227, 16'd20610, 16'd43182, 16'd6389, 16'd50361, 16'd29684, 16'd20141, 16'd16576, 16'd46992, 16'd14254, 16'd53149, 16'd40425, 16'd50078, 16'd31341, 16'd39613, 16'd624, 16'd24742, 16'd7679, 16'd3433, 16'd8030});
	test_expansion(128'h98de9d5885e0c1e12825ed94fde330bc, {16'd13763, 16'd15152, 16'd27399, 16'd6789, 16'd20373, 16'd30650, 16'd29590, 16'd37773, 16'd36036, 16'd27814, 16'd59264, 16'd42959, 16'd23182, 16'd65298, 16'd61351, 16'd2771, 16'd1928, 16'd5343, 16'd34688, 16'd23910, 16'd53102, 16'd13405, 16'd14639, 16'd9839, 16'd33013, 16'd40613});
	test_expansion(128'ha48f8175c7028676c07ef7e9e5cb22b4, {16'd35244, 16'd35093, 16'd50589, 16'd6515, 16'd63729, 16'd3004, 16'd8669, 16'd38239, 16'd19393, 16'd10519, 16'd4423, 16'd52099, 16'd48023, 16'd54505, 16'd60199, 16'd36442, 16'd916, 16'd12258, 16'd56285, 16'd9165, 16'd26051, 16'd42282, 16'd56256, 16'd29263, 16'd35742, 16'd38581});
	test_expansion(128'h6a3e110e21e6f28f5ac10cd7098d2b63, {16'd46397, 16'd63957, 16'd28322, 16'd58431, 16'd5460, 16'd40860, 16'd7450, 16'd64441, 16'd36490, 16'd36572, 16'd45129, 16'd30781, 16'd50052, 16'd18146, 16'd7399, 16'd6095, 16'd26138, 16'd47942, 16'd11541, 16'd34885, 16'd33081, 16'd35531, 16'd7561, 16'd28733, 16'd34207, 16'd54569});
	test_expansion(128'h4b653246f26a68a74389aa8a997ae138, {16'd45804, 16'd42882, 16'd57543, 16'd45577, 16'd52645, 16'd40795, 16'd14098, 16'd11752, 16'd31695, 16'd55264, 16'd23563, 16'd4712, 16'd48801, 16'd31113, 16'd43410, 16'd8509, 16'd45680, 16'd45075, 16'd64561, 16'd51784, 16'd32141, 16'd42881, 16'd33499, 16'd54669, 16'd57687, 16'd17901});
	test_expansion(128'h19b96e8a2ce8d423d08902325041dacd, {16'd35412, 16'd44787, 16'd56093, 16'd4932, 16'd24426, 16'd62625, 16'd32424, 16'd35038, 16'd15260, 16'd15818, 16'd11689, 16'd21201, 16'd26786, 16'd57535, 16'd55168, 16'd25246, 16'd48970, 16'd49815, 16'd9220, 16'd45355, 16'd7301, 16'd44432, 16'd61043, 16'd19113, 16'd39162, 16'd55536});
	test_expansion(128'hddbcc5451272e38cab20ea28c4179df5, {16'd47291, 16'd32183, 16'd372, 16'd5235, 16'd52192, 16'd35452, 16'd23016, 16'd10230, 16'd44304, 16'd43965, 16'd61230, 16'd19614, 16'd33373, 16'd37535, 16'd51056, 16'd11246, 16'd11665, 16'd13870, 16'd50977, 16'd43515, 16'd64519, 16'd58166, 16'd6032, 16'd24326, 16'd51069, 16'd54222});
	test_expansion(128'h173a2fc5ec74964d886a6f3933693fa3, {16'd36046, 16'd37944, 16'd7978, 16'd37475, 16'd26309, 16'd36884, 16'd5263, 16'd51898, 16'd15297, 16'd24777, 16'd20562, 16'd49508, 16'd86, 16'd44528, 16'd13512, 16'd15805, 16'd38114, 16'd22542, 16'd34946, 16'd13394, 16'd49902, 16'd26858, 16'd43468, 16'd27648, 16'd22250, 16'd52292});
	test_expansion(128'h339ce73bcd464197794101a62cbcbe9d, {16'd57978, 16'd48123, 16'd45802, 16'd43262, 16'd30399, 16'd18119, 16'd27332, 16'd8085, 16'd53336, 16'd33106, 16'd64721, 16'd1744, 16'd14625, 16'd30511, 16'd12201, 16'd39387, 16'd21980, 16'd48053, 16'd22945, 16'd35931, 16'd43145, 16'd2157, 16'd60, 16'd42353, 16'd64052, 16'd4085});
	test_expansion(128'hc2c852890b946b2c9dc5be9ffb879afe, {16'd45623, 16'd44998, 16'd13199, 16'd22595, 16'd2454, 16'd42979, 16'd57435, 16'd42795, 16'd1940, 16'd54351, 16'd52035, 16'd8646, 16'd27391, 16'd7640, 16'd7635, 16'd11251, 16'd57483, 16'd27594, 16'd41156, 16'd8499, 16'd2853, 16'd48083, 16'd49733, 16'd1858, 16'd37432, 16'd16515});
	test_expansion(128'h0489f8234931a17c092821b22b4aa8ea, {16'd60616, 16'd38665, 16'd4453, 16'd56078, 16'd9220, 16'd4600, 16'd20436, 16'd49728, 16'd31716, 16'd32876, 16'd58746, 16'd440, 16'd7559, 16'd12380, 16'd42948, 16'd13546, 16'd50971, 16'd46263, 16'd41575, 16'd4298, 16'd25346, 16'd48575, 16'd34655, 16'd45161, 16'd59739, 16'd17490});
	test_expansion(128'h20d03f7d7666e3223edc57c15a97c4fd, {16'd16410, 16'd25243, 16'd15411, 16'd60773, 16'd63048, 16'd65464, 16'd3257, 16'd3598, 16'd50239, 16'd6205, 16'd33392, 16'd60868, 16'd30897, 16'd32592, 16'd25184, 16'd14617, 16'd12560, 16'd7045, 16'd45281, 16'd40029, 16'd27510, 16'd60627, 16'd48363, 16'd33500, 16'd62797, 16'd16745});
	test_expansion(128'hecd0c7c87f765e01495c5c28530dbef9, {16'd52046, 16'd50184, 16'd42125, 16'd48781, 16'd3789, 16'd14003, 16'd33085, 16'd3809, 16'd4379, 16'd15567, 16'd49568, 16'd62057, 16'd41321, 16'd107, 16'd42196, 16'd8922, 16'd12003, 16'd54361, 16'd40117, 16'd31433, 16'd64260, 16'd17370, 16'd43238, 16'd16617, 16'd50100, 16'd15345});
	test_expansion(128'h30934b8d6bfd7699c649e08028ada4a0, {16'd21134, 16'd15548, 16'd62263, 16'd41633, 16'd15807, 16'd57151, 16'd23313, 16'd44669, 16'd17422, 16'd65298, 16'd20142, 16'd44873, 16'd712, 16'd664, 16'd50291, 16'd59995, 16'd21441, 16'd14832, 16'd9292, 16'd53574, 16'd58309, 16'd51030, 16'd29565, 16'd62419, 16'd32095, 16'd37461});
	test_expansion(128'hca170c4d0e7771ef1426c280f379bb11, {16'd9592, 16'd19439, 16'd43561, 16'd1930, 16'd37915, 16'd32583, 16'd28620, 16'd64847, 16'd28397, 16'd5888, 16'd34905, 16'd15958, 16'd17570, 16'd38307, 16'd53352, 16'd31873, 16'd34741, 16'd6899, 16'd59580, 16'd29388, 16'd40040, 16'd14660, 16'd34981, 16'd33016, 16'd7284, 16'd40819});
	test_expansion(128'hf8f34ef7ae848f6dfa6520bc610899f8, {16'd10573, 16'd24991, 16'd54007, 16'd50167, 16'd20470, 16'd10734, 16'd14938, 16'd3698, 16'd43217, 16'd11993, 16'd20035, 16'd40604, 16'd15184, 16'd27801, 16'd38877, 16'd53650, 16'd13221, 16'd58173, 16'd2859, 16'd64187, 16'd15818, 16'd59081, 16'd54170, 16'd60334, 16'd65232, 16'd17074});
	test_expansion(128'hebe0e05e6ddbd6fcf41394e72556c21a, {16'd25285, 16'd56452, 16'd1687, 16'd32983, 16'd46538, 16'd644, 16'd12428, 16'd10463, 16'd12846, 16'd33611, 16'd30161, 16'd48010, 16'd43883, 16'd34574, 16'd14501, 16'd3158, 16'd39230, 16'd4915, 16'd33793, 16'd42746, 16'd8768, 16'd45305, 16'd48799, 16'd3081, 16'd22253, 16'd21080});
	test_expansion(128'h045e943a384083b50cdcc699a796be75, {16'd18854, 16'd5349, 16'd62712, 16'd4178, 16'd391, 16'd19447, 16'd52677, 16'd55810, 16'd47770, 16'd5124, 16'd62525, 16'd60535, 16'd16767, 16'd11018, 16'd52322, 16'd13276, 16'd33702, 16'd3285, 16'd46948, 16'd57113, 16'd10919, 16'd34187, 16'd43341, 16'd9411, 16'd5598, 16'd51141});
	test_expansion(128'h30d0c1078df55d210b03b46502554758, {16'd18790, 16'd64218, 16'd64967, 16'd34776, 16'd34631, 16'd52205, 16'd61790, 16'd49160, 16'd24580, 16'd29013, 16'd50046, 16'd10574, 16'd56004, 16'd14773, 16'd35781, 16'd47919, 16'd18796, 16'd8102, 16'd26586, 16'd50696, 16'd33835, 16'd31695, 16'd20175, 16'd2909, 16'd30995, 16'd34333});
	test_expansion(128'heb9358a92ea81fa19fa595b92e5876dd, {16'd22437, 16'd51298, 16'd5487, 16'd64179, 16'd52632, 16'd11871, 16'd44622, 16'd27814, 16'd60749, 16'd51111, 16'd6113, 16'd21164, 16'd35326, 16'd37172, 16'd35066, 16'd46828, 16'd58872, 16'd30950, 16'd9705, 16'd42969, 16'd8718, 16'd2897, 16'd1778, 16'd42307, 16'd50478, 16'd22206});
	test_expansion(128'h2a6318aaf51a1db100fb4ccab6abb4f4, {16'd34534, 16'd20716, 16'd63502, 16'd2074, 16'd50713, 16'd42633, 16'd58296, 16'd48622, 16'd22267, 16'd64715, 16'd62756, 16'd64072, 16'd52875, 16'd14932, 16'd36988, 16'd10968, 16'd14520, 16'd14442, 16'd4715, 16'd23178, 16'd54931, 16'd7215, 16'd21452, 16'd47964, 16'd30564, 16'd58401});
	test_expansion(128'h18fb3e54f66c09db4e5c831568d582e8, {16'd7938, 16'd16093, 16'd26151, 16'd27004, 16'd26206, 16'd61732, 16'd45803, 16'd44073, 16'd13807, 16'd5973, 16'd12168, 16'd21515, 16'd45461, 16'd29910, 16'd48283, 16'd9989, 16'd6137, 16'd47923, 16'd17846, 16'd46822, 16'd52412, 16'd58858, 16'd55535, 16'd1097, 16'd62418, 16'd51082});
	test_expansion(128'h9a2268eeb8e72fdb99850237afa1d5ee, {16'd62002, 16'd43403, 16'd48919, 16'd33747, 16'd1042, 16'd21012, 16'd45571, 16'd50407, 16'd19481, 16'd17382, 16'd63935, 16'd41326, 16'd55943, 16'd58925, 16'd60593, 16'd51669, 16'd12102, 16'd261, 16'd14272, 16'd60528, 16'd10497, 16'd55899, 16'd10515, 16'd27164, 16'd57086, 16'd58770});
	test_expansion(128'h6778b64543ded25a8b8631669b6995ee, {16'd43833, 16'd32317, 16'd24736, 16'd50446, 16'd44731, 16'd50720, 16'd15271, 16'd26743, 16'd1669, 16'd41230, 16'd55934, 16'd52116, 16'd47589, 16'd7882, 16'd24360, 16'd15799, 16'd62937, 16'd6505, 16'd61015, 16'd56341, 16'd40146, 16'd32832, 16'd31036, 16'd18519, 16'd6587, 16'd26196});
	test_expansion(128'hc0f620fd5d8c33aaedb3880de71e5987, {16'd13408, 16'd1653, 16'd44993, 16'd9570, 16'd18173, 16'd56940, 16'd62820, 16'd43978, 16'd8519, 16'd63765, 16'd40618, 16'd58847, 16'd14455, 16'd65348, 16'd42329, 16'd49908, 16'd18861, 16'd18979, 16'd37877, 16'd35676, 16'd64338, 16'd55776, 16'd47840, 16'd57148, 16'd731, 16'd26753});
	test_expansion(128'h09bad3ac0cca5f11380e98b5083dadac, {16'd49322, 16'd35726, 16'd51243, 16'd24588, 16'd42078, 16'd10031, 16'd65029, 16'd34914, 16'd44027, 16'd37340, 16'd56592, 16'd6946, 16'd55400, 16'd59067, 16'd1922, 16'd33062, 16'd17161, 16'd25366, 16'd33884, 16'd24185, 16'd58038, 16'd7364, 16'd25049, 16'd7021, 16'd44607, 16'd42130});
	test_expansion(128'h457a6d6e3ebf8e5a79ced9c97020c623, {16'd50778, 16'd23289, 16'd16795, 16'd17553, 16'd39578, 16'd62076, 16'd8303, 16'd992, 16'd48433, 16'd10500, 16'd62072, 16'd6089, 16'd27431, 16'd30905, 16'd65512, 16'd21505, 16'd24764, 16'd20113, 16'd34918, 16'd64825, 16'd8872, 16'd55809, 16'd44693, 16'd46286, 16'd45010, 16'd64077});
	test_expansion(128'hb25e5222235ba84c40b64880cbc9cd33, {16'd38707, 16'd28016, 16'd36073, 16'd59403, 16'd38507, 16'd61057, 16'd11839, 16'd7061, 16'd26339, 16'd36416, 16'd33334, 16'd16643, 16'd10239, 16'd45119, 16'd45026, 16'd4825, 16'd60711, 16'd13366, 16'd14611, 16'd4685, 16'd42059, 16'd55789, 16'd18930, 16'd9612, 16'd2222, 16'd43591});
	test_expansion(128'h98568b6e208ae9759db48e6b42a2ca68, {16'd28806, 16'd36656, 16'd9798, 16'd55634, 16'd20804, 16'd49719, 16'd43261, 16'd47842, 16'd50867, 16'd61380, 16'd9247, 16'd38519, 16'd43427, 16'd45942, 16'd57090, 16'd518, 16'd60836, 16'd54607, 16'd28681, 16'd7134, 16'd51237, 16'd27321, 16'd35608, 16'd63267, 16'd29849, 16'd381});
	test_expansion(128'h0f7cd4c3fa58525c90a76c4227453f78, {16'd6759, 16'd32685, 16'd21782, 16'd43285, 16'd13982, 16'd57204, 16'd30229, 16'd12603, 16'd109, 16'd14870, 16'd36535, 16'd45400, 16'd12673, 16'd37489, 16'd19652, 16'd26615, 16'd35506, 16'd33958, 16'd35071, 16'd46445, 16'd34673, 16'd4769, 16'd25653, 16'd16493, 16'd12605, 16'd846});
	test_expansion(128'hd650cf7da65c82a156c0cb5c9734285a, {16'd3275, 16'd1363, 16'd2823, 16'd64634, 16'd25400, 16'd58870, 16'd7742, 16'd53718, 16'd51693, 16'd23682, 16'd54365, 16'd2587, 16'd30999, 16'd14522, 16'd19306, 16'd18021, 16'd54337, 16'd31344, 16'd47408, 16'd32368, 16'd43469, 16'd48581, 16'd4405, 16'd869, 16'd35870, 16'd17147});
	test_expansion(128'h19e4f9e5000b575571f5249e77236b66, {16'd55796, 16'd15019, 16'd64520, 16'd6131, 16'd61619, 16'd21039, 16'd5598, 16'd54497, 16'd16573, 16'd18626, 16'd60286, 16'd34678, 16'd39622, 16'd2560, 16'd58043, 16'd21686, 16'd15855, 16'd51768, 16'd809, 16'd56108, 16'd18355, 16'd42455, 16'd29288, 16'd58474, 16'd62980, 16'd31524});
	test_expansion(128'h472586a3ecea9f3684d44ff72be208aa, {16'd55134, 16'd12464, 16'd23021, 16'd64352, 16'd20089, 16'd58899, 16'd39200, 16'd5756, 16'd41841, 16'd49774, 16'd41565, 16'd39792, 16'd26131, 16'd56334, 16'd62238, 16'd33783, 16'd37704, 16'd59533, 16'd31955, 16'd44586, 16'd63621, 16'd18686, 16'd35940, 16'd10589, 16'd32825, 16'd30755});
	test_expansion(128'hdea68fc14494a64149695fca6fe79ea8, {16'd40408, 16'd21979, 16'd28352, 16'd59903, 16'd15062, 16'd8353, 16'd57588, 16'd47062, 16'd62355, 16'd36591, 16'd47141, 16'd54496, 16'd1164, 16'd65090, 16'd46616, 16'd36508, 16'd8697, 16'd8522, 16'd64776, 16'd50120, 16'd48921, 16'd19020, 16'd63921, 16'd51824, 16'd20984, 16'd45493});
	test_expansion(128'ha352c84ac98922b6edf0e52ac05bfb23, {16'd61764, 16'd52509, 16'd7107, 16'd27128, 16'd29954, 16'd11041, 16'd50677, 16'd49545, 16'd34661, 16'd46978, 16'd13048, 16'd1057, 16'd46440, 16'd38043, 16'd5070, 16'd53169, 16'd53524, 16'd21402, 16'd18352, 16'd15388, 16'd27418, 16'd63111, 16'd10820, 16'd30309, 16'd38878, 16'd4617});
	test_expansion(128'h470a2fa744857bd2707404c1b6547c04, {16'd37101, 16'd42274, 16'd18804, 16'd34756, 16'd3687, 16'd19343, 16'd54482, 16'd48680, 16'd2143, 16'd33753, 16'd2134, 16'd38632, 16'd20171, 16'd17356, 16'd13361, 16'd6748, 16'd62728, 16'd22846, 16'd39828, 16'd64675, 16'd31933, 16'd56499, 16'd39829, 16'd31086, 16'd30494, 16'd40309});
	test_expansion(128'hfe8d352cb00368f928c63afb17cccf76, {16'd33258, 16'd31422, 16'd38262, 16'd34962, 16'd13974, 16'd59409, 16'd35192, 16'd60222, 16'd26653, 16'd15088, 16'd53922, 16'd45499, 16'd15759, 16'd12355, 16'd50603, 16'd30386, 16'd21494, 16'd50671, 16'd26124, 16'd24038, 16'd57957, 16'd1910, 16'd14065, 16'd64760, 16'd12049, 16'd20613});
	test_expansion(128'h12c7cef313aa45b1b450efedde4dedd2, {16'd25982, 16'd19925, 16'd5713, 16'd64923, 16'd38754, 16'd7608, 16'd26652, 16'd11818, 16'd3754, 16'd967, 16'd86, 16'd3456, 16'd65055, 16'd46900, 16'd29065, 16'd4846, 16'd18896, 16'd16847, 16'd62940, 16'd52145, 16'd11613, 16'd5562, 16'd38926, 16'd60364, 16'd50711, 16'd47235});
	test_expansion(128'h6460c237746a1ce1e2329f614b07d386, {16'd28753, 16'd40587, 16'd18682, 16'd31336, 16'd8884, 16'd55182, 16'd59244, 16'd26769, 16'd38501, 16'd27102, 16'd59161, 16'd9594, 16'd29231, 16'd58023, 16'd39926, 16'd39868, 16'd64507, 16'd56366, 16'd60816, 16'd1076, 16'd61112, 16'd18380, 16'd52751, 16'd1088, 16'd15373, 16'd13411});
	test_expansion(128'h3c872257ca2310f520191b0350fafd4f, {16'd58736, 16'd5871, 16'd4887, 16'd62840, 16'd21237, 16'd53550, 16'd38231, 16'd12718, 16'd40339, 16'd15587, 16'd40267, 16'd27418, 16'd9435, 16'd64003, 16'd29062, 16'd57569, 16'd38371, 16'd19095, 16'd9362, 16'd11805, 16'd18599, 16'd36917, 16'd39875, 16'd6943, 16'd47611, 16'd669});
	test_expansion(128'h8d6382d12f5eb540c4a1e56d95bb34b1, {16'd15635, 16'd12601, 16'd26266, 16'd36049, 16'd21578, 16'd58054, 16'd46637, 16'd56266, 16'd42972, 16'd6452, 16'd36194, 16'd54378, 16'd38813, 16'd34896, 16'd2653, 16'd4151, 16'd28249, 16'd49200, 16'd37630, 16'd5154, 16'd43289, 16'd2997, 16'd32941, 16'd59676, 16'd8794, 16'd27755});
	test_expansion(128'h38cb92572a11078f4ed0cd8ca09e15dd, {16'd32683, 16'd43368, 16'd57513, 16'd63964, 16'd26846, 16'd49379, 16'd26904, 16'd64257, 16'd61102, 16'd1477, 16'd42281, 16'd5510, 16'd33426, 16'd43893, 16'd10228, 16'd23540, 16'd57879, 16'd44169, 16'd36369, 16'd49089, 16'd13832, 16'd43475, 16'd58251, 16'd46687, 16'd5176, 16'd34618});
	test_expansion(128'h44361f58e945f4c553a286b001b2fc0c, {16'd37778, 16'd24398, 16'd36029, 16'd572, 16'd27234, 16'd34547, 16'd5338, 16'd54793, 16'd18691, 16'd15854, 16'd53038, 16'd531, 16'd47756, 16'd63737, 16'd29711, 16'd27004, 16'd46262, 16'd3875, 16'd36233, 16'd52502, 16'd55855, 16'd2093, 16'd55596, 16'd31227, 16'd45435, 16'd52125});
	test_expansion(128'hcc49692dfd2559cdd1aa0fcccc6ecb2f, {16'd38674, 16'd47381, 16'd18901, 16'd42343, 16'd17553, 16'd26269, 16'd48543, 16'd63239, 16'd12401, 16'd50381, 16'd44045, 16'd62121, 16'd25499, 16'd14358, 16'd38588, 16'd52328, 16'd5937, 16'd44943, 16'd12483, 16'd62128, 16'd41924, 16'd13354, 16'd192, 16'd62862, 16'd8766, 16'd5762});
	test_expansion(128'hc39817c964c0a66dc2f441fdb27f5ff1, {16'd27839, 16'd2635, 16'd19779, 16'd40743, 16'd30083, 16'd47216, 16'd65533, 16'd56996, 16'd58417, 16'd10217, 16'd56615, 16'd52663, 16'd8723, 16'd7210, 16'd21218, 16'd32958, 16'd28490, 16'd60610, 16'd52955, 16'd45970, 16'd52231, 16'd31215, 16'd61952, 16'd43569, 16'd43509, 16'd11177});
	test_expansion(128'h2ab10e116b0da941e78c8d76b21e9c47, {16'd11942, 16'd17340, 16'd12476, 16'd13784, 16'd18028, 16'd12589, 16'd5285, 16'd54969, 16'd60540, 16'd24578, 16'd9097, 16'd57968, 16'd18143, 16'd36502, 16'd6831, 16'd14104, 16'd22062, 16'd29464, 16'd61704, 16'd52617, 16'd42083, 16'd44778, 16'd53014, 16'd16593, 16'd48756, 16'd15670});
	test_expansion(128'he445186962b517c424ad8382547283f4, {16'd18508, 16'd21596, 16'd42586, 16'd26186, 16'd44108, 16'd48085, 16'd48567, 16'd11283, 16'd43103, 16'd23122, 16'd45597, 16'd6259, 16'd51540, 16'd4481, 16'd40351, 16'd30056, 16'd41980, 16'd50299, 16'd21334, 16'd39111, 16'd39467, 16'd34531, 16'd20434, 16'd54986, 16'd1815, 16'd6179});
	test_expansion(128'h61c687b4e5bb3cd7388de7c03a7dc063, {16'd30847, 16'd17374, 16'd22263, 16'd36777, 16'd55527, 16'd3630, 16'd1723, 16'd62874, 16'd39774, 16'd42634, 16'd17604, 16'd809, 16'd13095, 16'd49092, 16'd29231, 16'd30384, 16'd25235, 16'd55017, 16'd23792, 16'd43892, 16'd63610, 16'd58486, 16'd10895, 16'd4071, 16'd29512, 16'd7543});
	test_expansion(128'hb05cd12d4b6a08efb93ec232d849339b, {16'd19549, 16'd31473, 16'd29037, 16'd45467, 16'd28878, 16'd49329, 16'd64356, 16'd49451, 16'd12654, 16'd59337, 16'd47208, 16'd25379, 16'd55197, 16'd61841, 16'd43278, 16'd11981, 16'd40507, 16'd3126, 16'd13945, 16'd7265, 16'd25549, 16'd54554, 16'd30106, 16'd29811, 16'd49593, 16'd8676});
	test_expansion(128'h26647b38f4c4c3b518954d439356b094, {16'd39120, 16'd44140, 16'd3328, 16'd299, 16'd64937, 16'd43542, 16'd1535, 16'd8167, 16'd39810, 16'd43630, 16'd55639, 16'd49987, 16'd42002, 16'd23353, 16'd15358, 16'd1034, 16'd61656, 16'd38898, 16'd27528, 16'd15038, 16'd38411, 16'd35236, 16'd18013, 16'd36080, 16'd52888, 16'd54319});
	test_expansion(128'h52e396d470e9680eed8d9ee0e58cb768, {16'd63898, 16'd16028, 16'd47555, 16'd11410, 16'd63189, 16'd51991, 16'd39611, 16'd14560, 16'd36381, 16'd9020, 16'd28921, 16'd25990, 16'd22617, 16'd8537, 16'd20471, 16'd26008, 16'd58252, 16'd35927, 16'd19728, 16'd38063, 16'd54816, 16'd36485, 16'd29583, 16'd17754, 16'd38157, 16'd8219});
	test_expansion(128'he27de93beaa6f09a7a8157c781171cec, {16'd7182, 16'd35505, 16'd59241, 16'd13182, 16'd20383, 16'd38345, 16'd53599, 16'd35012, 16'd24900, 16'd65203, 16'd37633, 16'd25328, 16'd7961, 16'd31340, 16'd53847, 16'd50710, 16'd1045, 16'd24822, 16'd48552, 16'd24951, 16'd4942, 16'd38179, 16'd10395, 16'd51698, 16'd48613, 16'd56313});
	test_expansion(128'h0ad393ad721620bb607dc20cdaf09b34, {16'd54598, 16'd33334, 16'd36743, 16'd58567, 16'd28637, 16'd22313, 16'd48091, 16'd25636, 16'd47186, 16'd14769, 16'd55853, 16'd32594, 16'd15091, 16'd13065, 16'd53835, 16'd17695, 16'd1487, 16'd48499, 16'd43713, 16'd38282, 16'd32972, 16'd10332, 16'd30287, 16'd27273, 16'd33925, 16'd44509});
	test_expansion(128'hb90794bffb825bbfb6b99258d5e87c6b, {16'd55504, 16'd28517, 16'd56012, 16'd21645, 16'd52703, 16'd4595, 16'd59472, 16'd42384, 16'd16997, 16'd48739, 16'd37132, 16'd49669, 16'd51636, 16'd1520, 16'd58423, 16'd13443, 16'd24635, 16'd58463, 16'd11445, 16'd26785, 16'd47929, 16'd11608, 16'd40470, 16'd11592, 16'd43210, 16'd19706});
	test_expansion(128'h202e37e378b4df5b3f7aaf72f0fef8a6, {16'd8159, 16'd39822, 16'd8846, 16'd17215, 16'd644, 16'd46798, 16'd25966, 16'd64010, 16'd56690, 16'd12990, 16'd41189, 16'd28192, 16'd19331, 16'd13727, 16'd27003, 16'd34125, 16'd10392, 16'd29127, 16'd26736, 16'd30452, 16'd51964, 16'd41735, 16'd58687, 16'd20491, 16'd33025, 16'd10991});
	test_expansion(128'h0def16456052d300f77edb9bfdb984a4, {16'd55688, 16'd34869, 16'd11166, 16'd9186, 16'd22061, 16'd381, 16'd5512, 16'd9224, 16'd37782, 16'd45272, 16'd1140, 16'd30253, 16'd17044, 16'd56742, 16'd53210, 16'd17463, 16'd12356, 16'd62935, 16'd45423, 16'd30598, 16'd18699, 16'd35507, 16'd62764, 16'd23162, 16'd64042, 16'd63808});
	test_expansion(128'h3d1f61adba191a2a97e6cfdfaba66f3d, {16'd32096, 16'd26066, 16'd7060, 16'd13829, 16'd43835, 16'd11649, 16'd46768, 16'd50000, 16'd42162, 16'd52928, 16'd49288, 16'd22734, 16'd65124, 16'd18979, 16'd19867, 16'd19219, 16'd60220, 16'd57376, 16'd54024, 16'd60136, 16'd6153, 16'd2264, 16'd50596, 16'd52183, 16'd62332, 16'd29543});
	test_expansion(128'h32a522cf4aac0a0cd34ff479414a5b9f, {16'd48433, 16'd2240, 16'd28402, 16'd20652, 16'd16100, 16'd62039, 16'd6810, 16'd63638, 16'd24419, 16'd15634, 16'd36228, 16'd62018, 16'd8356, 16'd49951, 16'd50284, 16'd1270, 16'd38132, 16'd20032, 16'd59210, 16'd474, 16'd17171, 16'd5646, 16'd27946, 16'd8735, 16'd22259, 16'd65413});
	test_expansion(128'h065896de715909336b6b1199e31a48b7, {16'd57853, 16'd62214, 16'd14451, 16'd23507, 16'd60712, 16'd16954, 16'd13145, 16'd53902, 16'd31147, 16'd36591, 16'd5588, 16'd11497, 16'd10498, 16'd627, 16'd62589, 16'd26496, 16'd29910, 16'd26117, 16'd60304, 16'd28175, 16'd30111, 16'd56598, 16'd30800, 16'd9527, 16'd65417, 16'd12703});
	test_expansion(128'h3ab2589af159af020f90d3b48a288b4d, {16'd24179, 16'd17385, 16'd33018, 16'd22705, 16'd24374, 16'd52092, 16'd10925, 16'd62186, 16'd32390, 16'd13491, 16'd3051, 16'd29219, 16'd58168, 16'd63477, 16'd14250, 16'd37039, 16'd56638, 16'd36454, 16'd20396, 16'd5194, 16'd9144, 16'd62079, 16'd15640, 16'd53477, 16'd17192, 16'd3816});
	test_expansion(128'hfd41c30a86fa9761ed93e632e8dd45dd, {16'd48409, 16'd58797, 16'd59291, 16'd32327, 16'd63186, 16'd38193, 16'd23722, 16'd28656, 16'd45362, 16'd54342, 16'd63481, 16'd26515, 16'd958, 16'd60512, 16'd48236, 16'd16594, 16'd17462, 16'd58119, 16'd3562, 16'd44918, 16'd48047, 16'd33756, 16'd36909, 16'd53592, 16'd17899, 16'd43143});
	test_expansion(128'h03c324457d93ee01047cbdfbe952aa75, {16'd41013, 16'd15742, 16'd56301, 16'd17340, 16'd48312, 16'd64274, 16'd9555, 16'd27285, 16'd27615, 16'd12158, 16'd7679, 16'd15428, 16'd22977, 16'd51636, 16'd61526, 16'd64685, 16'd10066, 16'd56840, 16'd7196, 16'd3420, 16'd10339, 16'd28429, 16'd21245, 16'd5250, 16'd8281, 16'd60293});
	test_expansion(128'h7e82cc0fd6caf2616f5b1d1c62b77f7c, {16'd46024, 16'd13544, 16'd698, 16'd17478, 16'd7048, 16'd65204, 16'd51959, 16'd57495, 16'd18941, 16'd35111, 16'd36543, 16'd1076, 16'd51862, 16'd3127, 16'd58882, 16'd49681, 16'd61097, 16'd24938, 16'd44846, 16'd40733, 16'd22959, 16'd56485, 16'd63947, 16'd11661, 16'd36456, 16'd25957});
	test_expansion(128'h806de7de7beb993df2659003aadd1b38, {16'd64533, 16'd47159, 16'd16217, 16'd22626, 16'd5236, 16'd9179, 16'd52869, 16'd543, 16'd23377, 16'd9934, 16'd53830, 16'd24138, 16'd58495, 16'd9599, 16'd49109, 16'd5336, 16'd61228, 16'd36033, 16'd39430, 16'd59663, 16'd51068, 16'd12850, 16'd12000, 16'd15196, 16'd53312, 16'd12630});
	test_expansion(128'hf3c8f66e32006c4dc664b81b9a39be55, {16'd63710, 16'd24370, 16'd2481, 16'd14051, 16'd24050, 16'd54329, 16'd13265, 16'd32062, 16'd55316, 16'd22713, 16'd41176, 16'd8405, 16'd62054, 16'd14238, 16'd45615, 16'd2781, 16'd4374, 16'd39446, 16'd27143, 16'd44202, 16'd56328, 16'd58863, 16'd34922, 16'd16687, 16'd54408, 16'd28103});
	test_expansion(128'h7c37a1a1d5e6c27cf3286c579f8026f9, {16'd17403, 16'd25942, 16'd32721, 16'd20183, 16'd37556, 16'd63879, 16'd28427, 16'd16172, 16'd62928, 16'd7081, 16'd20691, 16'd57554, 16'd11384, 16'd28724, 16'd34599, 16'd23778, 16'd4277, 16'd18856, 16'd23016, 16'd27341, 16'd62977, 16'd43826, 16'd4212, 16'd53385, 16'd38625, 16'd62306});
	test_expansion(128'h9cfce7fe6e4e8f2e57c8b9b196f8674d, {16'd19561, 16'd17147, 16'd25816, 16'd25907, 16'd14351, 16'd52237, 16'd52628, 16'd33931, 16'd543, 16'd54289, 16'd46416, 16'd19352, 16'd61570, 16'd60010, 16'd52535, 16'd5097, 16'd33061, 16'd349, 16'd21794, 16'd40347, 16'd62210, 16'd24666, 16'd15678, 16'd44343, 16'd64818, 16'd48608});
	test_expansion(128'hdb2aee296ca98147e081ae6fdfe3fec0, {16'd42127, 16'd62322, 16'd33019, 16'd43556, 16'd14842, 16'd57661, 16'd18532, 16'd33221, 16'd53183, 16'd25034, 16'd33031, 16'd62010, 16'd44404, 16'd46380, 16'd36135, 16'd41177, 16'd36337, 16'd21126, 16'd31001, 16'd19639, 16'd42430, 16'd12194, 16'd19841, 16'd33446, 16'd35637, 16'd3166});
	test_expansion(128'hf002e268248fc3738035d3191f7247ea, {16'd5630, 16'd13134, 16'd31571, 16'd61414, 16'd22287, 16'd54067, 16'd20819, 16'd20111, 16'd26657, 16'd232, 16'd45808, 16'd53641, 16'd45334, 16'd33977, 16'd17464, 16'd56494, 16'd25962, 16'd37790, 16'd5092, 16'd54997, 16'd6773, 16'd55418, 16'd22675, 16'd42916, 16'd39042, 16'd1629});
	test_expansion(128'h937ce7e3dc7d1bc7b8d89a15ac8b55f1, {16'd11583, 16'd40802, 16'd282, 16'd23050, 16'd20359, 16'd54689, 16'd35388, 16'd34809, 16'd20460, 16'd11230, 16'd64193, 16'd54808, 16'd60330, 16'd40221, 16'd11587, 16'd28013, 16'd52880, 16'd54572, 16'd6054, 16'd30577, 16'd21087, 16'd40373, 16'd1707, 16'd65344, 16'd1537, 16'd59958});
	test_expansion(128'h097ab33c4ab9ad640f81b6ea3eaeed6f, {16'd31807, 16'd30249, 16'd17395, 16'd24446, 16'd23093, 16'd12203, 16'd64370, 16'd34018, 16'd21544, 16'd20819, 16'd9011, 16'd16046, 16'd30454, 16'd16896, 16'd34610, 16'd29607, 16'd8636, 16'd31732, 16'd44049, 16'd29404, 16'd48738, 16'd52023, 16'd22092, 16'd11989, 16'd20377, 16'd45509});
	test_expansion(128'hbc7da9d1b8eaf9cd39a315a9be872d9c, {16'd62989, 16'd2024, 16'd26867, 16'd65240, 16'd10862, 16'd56258, 16'd13700, 16'd51459, 16'd22003, 16'd63887, 16'd40234, 16'd59322, 16'd52689, 16'd60128, 16'd27151, 16'd36343, 16'd46060, 16'd2145, 16'd596, 16'd19668, 16'd21330, 16'd53839, 16'd60997, 16'd37234, 16'd1176, 16'd60906});
	test_expansion(128'hf0be3436bc9622dc4b2bb4c6d7b4aada, {16'd12992, 16'd38878, 16'd19139, 16'd46195, 16'd24296, 16'd58018, 16'd7563, 16'd20789, 16'd39293, 16'd14948, 16'd58242, 16'd59861, 16'd42810, 16'd44044, 16'd31095, 16'd19516, 16'd23600, 16'd21569, 16'd13436, 16'd2449, 16'd13353, 16'd36513, 16'd37324, 16'd51804, 16'd28754, 16'd61720});
	test_expansion(128'hae64d4a4e61b46e598d09cd103637623, {16'd34872, 16'd34048, 16'd8184, 16'd49216, 16'd38055, 16'd15640, 16'd62926, 16'd35035, 16'd14983, 16'd37100, 16'd2001, 16'd24064, 16'd61813, 16'd7362, 16'd62753, 16'd51150, 16'd2586, 16'd48734, 16'd13732, 16'd26505, 16'd12120, 16'd22067, 16'd28873, 16'd39658, 16'd53394, 16'd8558});
	test_expansion(128'h8325c5d5cebc72a6686e66027baa72b5, {16'd4451, 16'd61906, 16'd17462, 16'd21809, 16'd40159, 16'd37213, 16'd34011, 16'd11613, 16'd43187, 16'd50860, 16'd58995, 16'd39703, 16'd19193, 16'd55745, 16'd16831, 16'd23552, 16'd59680, 16'd47941, 16'd9946, 16'd21508, 16'd27648, 16'd28343, 16'd61317, 16'd8879, 16'd51983, 16'd25612});
	test_expansion(128'hd5ce46f121ebedcf50e61bf3129577fb, {16'd35509, 16'd28245, 16'd58850, 16'd49223, 16'd10736, 16'd41008, 16'd29243, 16'd316, 16'd45496, 16'd22410, 16'd1656, 16'd17146, 16'd49031, 16'd37494, 16'd60511, 16'd9958, 16'd50489, 16'd30725, 16'd7190, 16'd43110, 16'd49788, 16'd58619, 16'd46728, 16'd1939, 16'd33747, 16'd50936});
	test_expansion(128'h446f8c846c1169f0c067e5f953954a3d, {16'd40395, 16'd33807, 16'd16905, 16'd38819, 16'd51275, 16'd4830, 16'd62497, 16'd63608, 16'd20123, 16'd2983, 16'd18536, 16'd2446, 16'd56426, 16'd20605, 16'd58557, 16'd36354, 16'd44911, 16'd32184, 16'd15995, 16'd64743, 16'd41344, 16'd32599, 16'd65148, 16'd36773, 16'd22871, 16'd52465});
	test_expansion(128'h071e29df1923ef62464bea487ef92067, {16'd33721, 16'd62691, 16'd6355, 16'd40039, 16'd45274, 16'd42506, 16'd52209, 16'd953, 16'd11633, 16'd6223, 16'd13752, 16'd11422, 16'd9667, 16'd13629, 16'd14158, 16'd5793, 16'd25793, 16'd34879, 16'd7038, 16'd47850, 16'd23733, 16'd26854, 16'd9582, 16'd50196, 16'd12037, 16'd46436});
	test_expansion(128'hecb31c7abb9a8e768600ad400fde2fba, {16'd51480, 16'd27209, 16'd10073, 16'd23859, 16'd59739, 16'd17165, 16'd2845, 16'd13754, 16'd4775, 16'd39464, 16'd32770, 16'd52724, 16'd19532, 16'd57412, 16'd17376, 16'd58922, 16'd52505, 16'd48662, 16'd16620, 16'd31886, 16'd629, 16'd26766, 16'd64679, 16'd32893, 16'd59809, 16'd57146});
	test_expansion(128'ha76a1120160608c7f94a52cfc3fa8490, {16'd64769, 16'd57462, 16'd51293, 16'd38166, 16'd1299, 16'd29588, 16'd55926, 16'd47288, 16'd36146, 16'd49150, 16'd9955, 16'd32326, 16'd52710, 16'd4588, 16'd16255, 16'd42847, 16'd59259, 16'd29024, 16'd44519, 16'd12849, 16'd3902, 16'd8525, 16'd65407, 16'd37289, 16'd7287, 16'd29601});
	test_expansion(128'h7293d9f4198d49e3d9e40e1d3544f453, {16'd28612, 16'd16809, 16'd55786, 16'd28800, 16'd34765, 16'd2575, 16'd43738, 16'd46567, 16'd42039, 16'd38854, 16'd27399, 16'd54013, 16'd32087, 16'd25342, 16'd30745, 16'd26269, 16'd41236, 16'd35702, 16'd40444, 16'd46148, 16'd43547, 16'd41346, 16'd32880, 16'd34569, 16'd13747, 16'd50860});
	test_expansion(128'h3d696737fae29f90b9abd842297070bb, {16'd45945, 16'd48849, 16'd22940, 16'd439, 16'd9848, 16'd4026, 16'd62796, 16'd40775, 16'd20256, 16'd36752, 16'd10307, 16'd1418, 16'd44626, 16'd42169, 16'd53018, 16'd27690, 16'd64018, 16'd55033, 16'd44095, 16'd8964, 16'd23130, 16'd4383, 16'd43321, 16'd36256, 16'd29782, 16'd26387});
	test_expansion(128'h6099d913bf2aa7999dd6a167ddce460b, {16'd15108, 16'd17270, 16'd44021, 16'd15897, 16'd8595, 16'd65020, 16'd19566, 16'd16652, 16'd55264, 16'd48992, 16'd10167, 16'd56375, 16'd1921, 16'd42827, 16'd36115, 16'd10222, 16'd18700, 16'd17916, 16'd32130, 16'd25508, 16'd33080, 16'd19589, 16'd5902, 16'd27293, 16'd20103, 16'd35128});
	test_expansion(128'h5cb9c715ba10f541e4deeebd3a320b4b, {16'd2773, 16'd57522, 16'd62429, 16'd1486, 16'd17132, 16'd39709, 16'd57716, 16'd53523, 16'd53868, 16'd63371, 16'd59175, 16'd50427, 16'd30476, 16'd46704, 16'd47461, 16'd23514, 16'd55496, 16'd43493, 16'd3577, 16'd53708, 16'd34367, 16'd33677, 16'd25547, 16'd59427, 16'd30370, 16'd40952});
	test_expansion(128'he9c281626cf634f3de2d5730a1bc2fec, {16'd30923, 16'd46150, 16'd15386, 16'd9774, 16'd60412, 16'd31302, 16'd2574, 16'd59619, 16'd38630, 16'd23781, 16'd2194, 16'd62266, 16'd14069, 16'd18863, 16'd57741, 16'd14493, 16'd18759, 16'd5872, 16'd7019, 16'd53801, 16'd50331, 16'd24254, 16'd59347, 16'd50029, 16'd33720, 16'd63496});
	test_expansion(128'hab301659512d5d2d6a904c89d3fb51ae, {16'd61709, 16'd47645, 16'd26521, 16'd19, 16'd12908, 16'd15542, 16'd6197, 16'd62171, 16'd49122, 16'd49049, 16'd4745, 16'd37013, 16'd56858, 16'd62456, 16'd53978, 16'd51016, 16'd17929, 16'd3271, 16'd3560, 16'd56572, 16'd63483, 16'd39149, 16'd10445, 16'd48811, 16'd8756, 16'd65331});
	test_expansion(128'h92ff00b75c9a5c14f77a8ec8186eabf6, {16'd6452, 16'd24410, 16'd10498, 16'd43317, 16'd52845, 16'd14886, 16'd36771, 16'd60670, 16'd48527, 16'd60302, 16'd15397, 16'd25392, 16'd31465, 16'd50851, 16'd56431, 16'd12935, 16'd4653, 16'd3406, 16'd36130, 16'd59462, 16'd65059, 16'd28108, 16'd65301, 16'd2084, 16'd26709, 16'd31947});
	test_expansion(128'h09bb7ae8863aec88ef0aac1e6b7005c5, {16'd54167, 16'd52090, 16'd32303, 16'd22288, 16'd64060, 16'd2099, 16'd32917, 16'd2128, 16'd8150, 16'd7547, 16'd11082, 16'd43924, 16'd63991, 16'd32065, 16'd43166, 16'd24146, 16'd63629, 16'd42574, 16'd31950, 16'd6838, 16'd62901, 16'd41538, 16'd12435, 16'd61617, 16'd55239, 16'd3423});
	test_expansion(128'h998759537ed064d3970165b8288f9d28, {16'd52634, 16'd15229, 16'd48274, 16'd28, 16'd30979, 16'd45811, 16'd17341, 16'd32431, 16'd53317, 16'd37361, 16'd15251, 16'd50818, 16'd57349, 16'd46017, 16'd62392, 16'd758, 16'd54715, 16'd47255, 16'd11134, 16'd27723, 16'd4704, 16'd4787, 16'd12966, 16'd26663, 16'd11914, 16'd31673});
	test_expansion(128'h2b64562a559f9dd58ac0e7cf2d3b2516, {16'd46864, 16'd50027, 16'd54584, 16'd36445, 16'd16329, 16'd8408, 16'd1235, 16'd40289, 16'd39429, 16'd61294, 16'd44922, 16'd21372, 16'd22792, 16'd27931, 16'd36975, 16'd59460, 16'd14335, 16'd5571, 16'd29311, 16'd52640, 16'd46695, 16'd44015, 16'd53020, 16'd33947, 16'd32768, 16'd23046});
	test_expansion(128'hc9b4a4ae0d41e9ab7698bb2e4ee7e080, {16'd5120, 16'd29986, 16'd5805, 16'd14556, 16'd38361, 16'd34151, 16'd40546, 16'd5517, 16'd16643, 16'd57582, 16'd24397, 16'd54251, 16'd13267, 16'd38270, 16'd13571, 16'd54741, 16'd56964, 16'd33507, 16'd2180, 16'd54358, 16'd9396, 16'd31549, 16'd51770, 16'd15923, 16'd57726, 16'd29843});
	test_expansion(128'h8b84a49de7bb8aa1c3ced6af8a36ee1e, {16'd17794, 16'd65198, 16'd43000, 16'd48991, 16'd16992, 16'd33997, 16'd46207, 16'd2885, 16'd16492, 16'd9191, 16'd14771, 16'd24615, 16'd28085, 16'd51288, 16'd34108, 16'd3526, 16'd46870, 16'd43850, 16'd18456, 16'd35460, 16'd24739, 16'd4154, 16'd36519, 16'd22020, 16'd54105, 16'd35004});
	test_expansion(128'hc695e8d7030957962a415f3668444989, {16'd14411, 16'd56385, 16'd61276, 16'd36169, 16'd7720, 16'd26662, 16'd20862, 16'd54969, 16'd46834, 16'd34420, 16'd31210, 16'd60140, 16'd37665, 16'd59568, 16'd6995, 16'd21081, 16'd65295, 16'd13234, 16'd45176, 16'd18666, 16'd9755, 16'd37478, 16'd16899, 16'd32323, 16'd5539, 16'd25239});
	test_expansion(128'he54e1650a60ab9332a77c6e0952764ec, {16'd11822, 16'd47637, 16'd21168, 16'd47450, 16'd25760, 16'd22094, 16'd61415, 16'd4947, 16'd42957, 16'd8886, 16'd16933, 16'd56484, 16'd45173, 16'd64977, 16'd35181, 16'd51720, 16'd23660, 16'd25744, 16'd933, 16'd47665, 16'd44086, 16'd31665, 16'd10962, 16'd48508, 16'd60754, 16'd38612});
	test_expansion(128'h0e5a734a59bbe8d9cb6f51802c2064eb, {16'd35041, 16'd38183, 16'd61275, 16'd59006, 16'd27900, 16'd22419, 16'd29729, 16'd63294, 16'd35600, 16'd3296, 16'd49335, 16'd45315, 16'd30351, 16'd15232, 16'd27399, 16'd5604, 16'd24427, 16'd53327, 16'd40877, 16'd51676, 16'd61382, 16'd25492, 16'd39393, 16'd15526, 16'd63797, 16'd8039});
	test_expansion(128'h16d61be704c31b393b173a3352d74db7, {16'd22855, 16'd3036, 16'd43477, 16'd8216, 16'd56093, 16'd59189, 16'd61803, 16'd17317, 16'd64693, 16'd23250, 16'd59507, 16'd38919, 16'd18904, 16'd13722, 16'd54601, 16'd32142, 16'd35904, 16'd40805, 16'd49894, 16'd31946, 16'd64271, 16'd17192, 16'd8208, 16'd38752, 16'd44428, 16'd13340});
	test_expansion(128'hb344d420240a0692eab6c16083cbc358, {16'd51268, 16'd7510, 16'd8613, 16'd35856, 16'd34205, 16'd63494, 16'd39090, 16'd41491, 16'd57084, 16'd62158, 16'd16061, 16'd59127, 16'd53042, 16'd25012, 16'd17073, 16'd37723, 16'd25908, 16'd9459, 16'd36640, 16'd12338, 16'd17397, 16'd57242, 16'd26006, 16'd27071, 16'd22225, 16'd41222});
	test_expansion(128'h421972ca77e1e82da497e340e1bce6ae, {16'd41528, 16'd63381, 16'd44990, 16'd36094, 16'd40129, 16'd36049, 16'd61328, 16'd7126, 16'd39383, 16'd32364, 16'd55313, 16'd25135, 16'd42884, 16'd44832, 16'd49781, 16'd34267, 16'd25079, 16'd63257, 16'd3635, 16'd24465, 16'd3525, 16'd59695, 16'd40455, 16'd8907, 16'd3802, 16'd3008});
	test_expansion(128'hdafd22dc84c6658aadff251fe054255c, {16'd34619, 16'd55375, 16'd42548, 16'd31301, 16'd40385, 16'd38632, 16'd57171, 16'd59630, 16'd53138, 16'd18843, 16'd56133, 16'd36678, 16'd11271, 16'd47853, 16'd25037, 16'd5989, 16'd61969, 16'd32225, 16'd49291, 16'd23760, 16'd12325, 16'd51229, 16'd9470, 16'd39911, 16'd40096, 16'd764});
	test_expansion(128'ha625ad38300f9f653d0278b4df6a3d50, {16'd41140, 16'd44945, 16'd59095, 16'd682, 16'd48405, 16'd31446, 16'd35078, 16'd14830, 16'd64632, 16'd5654, 16'd31703, 16'd39085, 16'd36682, 16'd15225, 16'd39565, 16'd15044, 16'd16895, 16'd6680, 16'd23557, 16'd51190, 16'd54956, 16'd16585, 16'd16761, 16'd12364, 16'd54731, 16'd23185});
	test_expansion(128'h4bf4e629f3d31458734d12c30e328a75, {16'd54942, 16'd39367, 16'd63290, 16'd37502, 16'd25980, 16'd44828, 16'd32206, 16'd38265, 16'd12393, 16'd30255, 16'd17157, 16'd23471, 16'd10673, 16'd26410, 16'd42820, 16'd65271, 16'd42322, 16'd37852, 16'd11978, 16'd25925, 16'd31525, 16'd55183, 16'd24956, 16'd46362, 16'd38303, 16'd63440});
	test_expansion(128'h14f64e7722d40263a172bada849cd1e1, {16'd64496, 16'd40498, 16'd1497, 16'd25669, 16'd35880, 16'd13837, 16'd65478, 16'd8769, 16'd15055, 16'd18680, 16'd40077, 16'd49798, 16'd23173, 16'd23946, 16'd8066, 16'd33815, 16'd13493, 16'd47240, 16'd29277, 16'd1820, 16'd9252, 16'd21379, 16'd64646, 16'd28834, 16'd42977, 16'd62823});
	test_expansion(128'h0d6491f26da5b08176d208887426d528, {16'd4354, 16'd54726, 16'd53063, 16'd15934, 16'd44049, 16'd59870, 16'd14794, 16'd21737, 16'd42776, 16'd49119, 16'd53313, 16'd38943, 16'd51501, 16'd52710, 16'd2518, 16'd9026, 16'd47285, 16'd31910, 16'd7046, 16'd53213, 16'd53200, 16'd46186, 16'd26512, 16'd35370, 16'd11058, 16'd42229});
	test_expansion(128'h9aca1f57c4de4a48a007c0068499ff80, {16'd41909, 16'd41046, 16'd6135, 16'd28548, 16'd48117, 16'd18284, 16'd47203, 16'd33807, 16'd32093, 16'd45960, 16'd19621, 16'd55023, 16'd45588, 16'd17264, 16'd46628, 16'd37749, 16'd12505, 16'd53249, 16'd7941, 16'd61374, 16'd30438, 16'd20035, 16'd45736, 16'd13459, 16'd60212, 16'd11281});
	test_expansion(128'h90c73fdb5da372fc857284197844a7fd, {16'd28313, 16'd60936, 16'd43673, 16'd13792, 16'd58113, 16'd63961, 16'd63331, 16'd41449, 16'd59503, 16'd27104, 16'd27865, 16'd38490, 16'd47943, 16'd31222, 16'd36839, 16'd61285, 16'd38374, 16'd27074, 16'd41599, 16'd39055, 16'd7534, 16'd59976, 16'd7664, 16'd47072, 16'd7682, 16'd65273});
	test_expansion(128'haf19ad224b018a60b2a8829ea0762e15, {16'd19154, 16'd2082, 16'd40698, 16'd47950, 16'd21738, 16'd28291, 16'd27746, 16'd13227, 16'd49982, 16'd2730, 16'd53366, 16'd1095, 16'd21853, 16'd45333, 16'd17476, 16'd45111, 16'd28768, 16'd62691, 16'd65200, 16'd16050, 16'd16102, 16'd40167, 16'd14526, 16'd16369, 16'd54778, 16'd31804});
	test_expansion(128'hf8f1529773219ecaca1606fa1218c39a, {16'd61250, 16'd4170, 16'd64607, 16'd56491, 16'd62398, 16'd5863, 16'd15778, 16'd39870, 16'd59178, 16'd6500, 16'd37444, 16'd45522, 16'd60293, 16'd8353, 16'd26332, 16'd22392, 16'd28071, 16'd29545, 16'd41991, 16'd16550, 16'd2961, 16'd1191, 16'd47359, 16'd5231, 16'd36190, 16'd57586});
	test_expansion(128'hde8b48f5c17b2132654cb35b0f817d1b, {16'd52033, 16'd7928, 16'd59841, 16'd7493, 16'd9418, 16'd4490, 16'd33706, 16'd59097, 16'd51335, 16'd37379, 16'd8702, 16'd25111, 16'd44539, 16'd53024, 16'd60102, 16'd20866, 16'd5037, 16'd23965, 16'd43105, 16'd33054, 16'd58247, 16'd40015, 16'd14617, 16'd38722, 16'd15552, 16'd33393});
	test_expansion(128'h42cd5c880a9895e039f0a0b9b0a56164, {16'd51925, 16'd11582, 16'd22839, 16'd59188, 16'd44014, 16'd59674, 16'd23857, 16'd29027, 16'd45434, 16'd52437, 16'd12230, 16'd55526, 16'd20436, 16'd60276, 16'd47467, 16'd32391, 16'd1445, 16'd46356, 16'd53594, 16'd40720, 16'd36199, 16'd42091, 16'd51608, 16'd38587, 16'd45459, 16'd63033});
	test_expansion(128'h25a079906acf7e1fa32253284b751304, {16'd7195, 16'd32760, 16'd23441, 16'd23244, 16'd27501, 16'd24813, 16'd26612, 16'd46862, 16'd61168, 16'd49415, 16'd10695, 16'd29261, 16'd19005, 16'd52231, 16'd12705, 16'd6060, 16'd56312, 16'd64468, 16'd29217, 16'd30952, 16'd20615, 16'd18047, 16'd57953, 16'd30820, 16'd40800, 16'd24356});
	test_expansion(128'h47cc9fcac6b7455b8cc8292e8f880a93, {16'd43754, 16'd11390, 16'd58550, 16'd11378, 16'd64604, 16'd35862, 16'd11901, 16'd18918, 16'd47493, 16'd28420, 16'd36113, 16'd8842, 16'd30304, 16'd2714, 16'd42875, 16'd37803, 16'd50144, 16'd59588, 16'd9027, 16'd44807, 16'd57445, 16'd50068, 16'd58526, 16'd1905, 16'd27641, 16'd34497});
	test_expansion(128'h579ef869fab913f0d62604a5f7592619, {16'd58660, 16'd43170, 16'd34082, 16'd17341, 16'd52696, 16'd26759, 16'd21376, 16'd11511, 16'd9434, 16'd43739, 16'd4909, 16'd61751, 16'd55116, 16'd4059, 16'd43340, 16'd43053, 16'd56359, 16'd39724, 16'd40054, 16'd3228, 16'd31990, 16'd16214, 16'd18718, 16'd53824, 16'd2020, 16'd11700});
	test_expansion(128'hbed0ad2c1aeea285412d108590c19ae3, {16'd41550, 16'd54974, 16'd32676, 16'd12110, 16'd55114, 16'd27663, 16'd26495, 16'd34774, 16'd42899, 16'd3387, 16'd25815, 16'd112, 16'd51303, 16'd13681, 16'd56336, 16'd52232, 16'd16099, 16'd35862, 16'd64627, 16'd29947, 16'd3520, 16'd40516, 16'd30046, 16'd20766, 16'd15265, 16'd46469});
	test_expansion(128'hd3b61aa8bd43feec281ba1a84bc39856, {16'd5421, 16'd49917, 16'd49303, 16'd37326, 16'd41393, 16'd4181, 16'd58383, 16'd28800, 16'd39440, 16'd40059, 16'd40529, 16'd23636, 16'd22284, 16'd33315, 16'd19729, 16'd64976, 16'd51005, 16'd16898, 16'd31076, 16'd61682, 16'd24921, 16'd32156, 16'd61307, 16'd31074, 16'd26987, 16'd38722});
	test_expansion(128'hbef748bafe1ee3321e7937f63bbe1903, {16'd27199, 16'd62979, 16'd59725, 16'd60340, 16'd59227, 16'd9851, 16'd19041, 16'd49288, 16'd25754, 16'd51639, 16'd44953, 16'd46734, 16'd1236, 16'd14747, 16'd58766, 16'd14987, 16'd32356, 16'd55954, 16'd36080, 16'd55584, 16'd62846, 16'd862, 16'd35281, 16'd59509, 16'd12309, 16'd7450});
	test_expansion(128'hd4d64810fab0612a245bedc161b0cd01, {16'd50594, 16'd13568, 16'd63915, 16'd42673, 16'd53464, 16'd17418, 16'd28368, 16'd40373, 16'd45791, 16'd58835, 16'd18472, 16'd32037, 16'd53295, 16'd28559, 16'd50178, 16'd28646, 16'd31310, 16'd16679, 16'd63615, 16'd16114, 16'd24666, 16'd20491, 16'd42471, 16'd5385, 16'd14938, 16'd14806});
	test_expansion(128'h2608313729851ee57e09fe85c25cd4a8, {16'd23708, 16'd42254, 16'd26786, 16'd60876, 16'd22905, 16'd22624, 16'd51994, 16'd15015, 16'd30001, 16'd12568, 16'd45349, 16'd16045, 16'd18035, 16'd50601, 16'd48952, 16'd45785, 16'd21011, 16'd31837, 16'd64860, 16'd29759, 16'd11948, 16'd4114, 16'd9932, 16'd3022, 16'd24531, 16'd8462});
	test_expansion(128'h31e63178f5d02bf5fad68af40aa25d33, {16'd27813, 16'd5833, 16'd29537, 16'd48755, 16'd20918, 16'd33810, 16'd57179, 16'd28752, 16'd35870, 16'd35156, 16'd38606, 16'd53471, 16'd44713, 16'd45382, 16'd65304, 16'd31568, 16'd53414, 16'd50701, 16'd42728, 16'd38539, 16'd51179, 16'd59005, 16'd47823, 16'd26140, 16'd30169, 16'd2626});
	test_expansion(128'hfdf1e6e12b46a92968fded9e4302627e, {16'd7603, 16'd52928, 16'd44348, 16'd18505, 16'd53434, 16'd65255, 16'd46400, 16'd6016, 16'd23771, 16'd57512, 16'd45410, 16'd41638, 16'd42722, 16'd31323, 16'd27530, 16'd13924, 16'd47392, 16'd30440, 16'd58406, 16'd13149, 16'd23781, 16'd19962, 16'd7124, 16'd34761, 16'd40139, 16'd64598});
	test_expansion(128'h98e9cfa7ad12f9dfd9d9c21ada23b397, {16'd65211, 16'd20897, 16'd1715, 16'd45940, 16'd56665, 16'd60312, 16'd41790, 16'd5422, 16'd53731, 16'd58129, 16'd56729, 16'd14367, 16'd54583, 16'd26812, 16'd35950, 16'd26916, 16'd18931, 16'd792, 16'd43726, 16'd45012, 16'd2108, 16'd31904, 16'd33056, 16'd51980, 16'd35113, 16'd4187});
	test_expansion(128'hcc7992a59efb5c2b300bdbf535c8d0df, {16'd2280, 16'd64936, 16'd26816, 16'd14644, 16'd48059, 16'd35025, 16'd37369, 16'd61957, 16'd12217, 16'd18989, 16'd473, 16'd24740, 16'd27214, 16'd7555, 16'd60907, 16'd35029, 16'd43828, 16'd61233, 16'd39129, 16'd33305, 16'd2947, 16'd52712, 16'd41485, 16'd18059, 16'd56541, 16'd50089});
	test_expansion(128'hfa71d9b1e73576b23b4c6af529fd4fab, {16'd59153, 16'd59077, 16'd1312, 16'd1328, 16'd51041, 16'd20878, 16'd25618, 16'd31633, 16'd58284, 16'd20786, 16'd3696, 16'd55720, 16'd1661, 16'd15476, 16'd29755, 16'd29969, 16'd41741, 16'd34175, 16'd10844, 16'd31784, 16'd15247, 16'd5889, 16'd9730, 16'd8263, 16'd625, 16'd41441});
	test_expansion(128'he3ffc1ef1b56924531762aa5ce1a1081, {16'd45368, 16'd35391, 16'd22525, 16'd55297, 16'd5518, 16'd27605, 16'd6137, 16'd60823, 16'd16343, 16'd20400, 16'd32408, 16'd64275, 16'd47120, 16'd28923, 16'd5577, 16'd37170, 16'd63324, 16'd54471, 16'd10750, 16'd64198, 16'd27640, 16'd47485, 16'd22172, 16'd46349, 16'd29724, 16'd15397});
	test_expansion(128'hb6049257b30d29a178754496c4643869, {16'd34332, 16'd34781, 16'd28434, 16'd7796, 16'd43258, 16'd48051, 16'd10194, 16'd51510, 16'd34332, 16'd37210, 16'd4726, 16'd40843, 16'd14777, 16'd52012, 16'd11076, 16'd63936, 16'd23795, 16'd44901, 16'd8797, 16'd43098, 16'd28621, 16'd38030, 16'd3326, 16'd4418, 16'd49370, 16'd64529});
	test_expansion(128'h47b823c421b4ebabedabda71dd11b0f5, {16'd12208, 16'd32595, 16'd28162, 16'd11987, 16'd5771, 16'd19547, 16'd13707, 16'd40616, 16'd20821, 16'd62561, 16'd14479, 16'd34871, 16'd42466, 16'd10058, 16'd61923, 16'd17316, 16'd43743, 16'd3507, 16'd9606, 16'd47889, 16'd18299, 16'd20100, 16'd18766, 16'd38798, 16'd47434, 16'd38539});
	test_expansion(128'hf7de1a5ffb48c83c93d08e2a2179048d, {16'd51302, 16'd43823, 16'd41030, 16'd35310, 16'd6413, 16'd4541, 16'd22759, 16'd32744, 16'd38705, 16'd47011, 16'd20613, 16'd35260, 16'd6962, 16'd64262, 16'd56483, 16'd22271, 16'd13599, 16'd56941, 16'd26418, 16'd11504, 16'd30353, 16'd40069, 16'd60861, 16'd4021, 16'd61315, 16'd7017});
	test_expansion(128'h48e81e3fa567e6f567bf6ebaf7606dc4, {16'd19624, 16'd61395, 16'd8023, 16'd3051, 16'd47745, 16'd31509, 16'd31714, 16'd28145, 16'd64706, 16'd38893, 16'd65470, 16'd9872, 16'd41238, 16'd21147, 16'd33768, 16'd11938, 16'd2406, 16'd16191, 16'd39945, 16'd36293, 16'd22878, 16'd52698, 16'd30832, 16'd49875, 16'd30976, 16'd10313});
	test_expansion(128'h7496aa352055e94530c372ee9b2c0796, {16'd40989, 16'd56520, 16'd60877, 16'd15187, 16'd45279, 16'd56591, 16'd6097, 16'd34181, 16'd27304, 16'd9504, 16'd30183, 16'd17302, 16'd7548, 16'd60668, 16'd47124, 16'd31428, 16'd16049, 16'd37724, 16'd33098, 16'd40193, 16'd34226, 16'd13205, 16'd9927, 16'd13454, 16'd59392, 16'd49182});
	test_expansion(128'h9ed7a4ea3ba92f274063df17d6e1c797, {16'd47031, 16'd55896, 16'd8669, 16'd52575, 16'd38189, 16'd43314, 16'd22269, 16'd44917, 16'd38689, 16'd5139, 16'd52207, 16'd43679, 16'd14291, 16'd11410, 16'd48542, 16'd49964, 16'd65181, 16'd37222, 16'd52397, 16'd19639, 16'd42078, 16'd37913, 16'd11378, 16'd54474, 16'd5100, 16'd31476});
	test_expansion(128'ha27ead8cf23bfcfd55022685138cb2ff, {16'd29644, 16'd35634, 16'd50537, 16'd55723, 16'd46055, 16'd52518, 16'd11999, 16'd60964, 16'd14319, 16'd41422, 16'd56182, 16'd48025, 16'd30763, 16'd53795, 16'd8584, 16'd26067, 16'd10857, 16'd61262, 16'd28368, 16'd42634, 16'd22476, 16'd15810, 16'd18073, 16'd20303, 16'd27838, 16'd57549});
	test_expansion(128'ha79e629048cdccae0ffce728586b4fb4, {16'd56087, 16'd55013, 16'd38480, 16'd17296, 16'd44663, 16'd49534, 16'd25059, 16'd47088, 16'd42352, 16'd27959, 16'd43934, 16'd64563, 16'd14505, 16'd38389, 16'd57274, 16'd18150, 16'd44331, 16'd64510, 16'd32106, 16'd55672, 16'd37949, 16'd14754, 16'd56970, 16'd19442, 16'd51956, 16'd37920});
	test_expansion(128'he04735354d47f3fe6245d779e8dc9918, {16'd19575, 16'd15858, 16'd61173, 16'd15159, 16'd11569, 16'd18352, 16'd9271, 16'd21124, 16'd16183, 16'd24770, 16'd32740, 16'd11617, 16'd64372, 16'd6445, 16'd24980, 16'd10215, 16'd48456, 16'd19512, 16'd15840, 16'd44983, 16'd2691, 16'd32077, 16'd50494, 16'd12090, 16'd45324, 16'd62311});
	test_expansion(128'h486c4a66a8d850756728e8635748f94a, {16'd26596, 16'd6635, 16'd20722, 16'd25254, 16'd4396, 16'd62607, 16'd31610, 16'd65426, 16'd54597, 16'd29760, 16'd6648, 16'd32612, 16'd27488, 16'd9471, 16'd26927, 16'd32306, 16'd56249, 16'd58392, 16'd6460, 16'd42769, 16'd60719, 16'd33888, 16'd14857, 16'd2779, 16'd23810, 16'd62077});
	test_expansion(128'h0595056ea4193424a1f0a7bd8e58f208, {16'd31444, 16'd26379, 16'd11370, 16'd37592, 16'd9717, 16'd43532, 16'd54939, 16'd57962, 16'd52857, 16'd18716, 16'd54861, 16'd54262, 16'd32179, 16'd16211, 16'd33753, 16'd397, 16'd11801, 16'd20408, 16'd58091, 16'd49379, 16'd37161, 16'd20489, 16'd12787, 16'd25681, 16'd62513, 16'd14170});
	test_expansion(128'h542b1de6ab2b235d31e65ed58e9bf6e9, {16'd10176, 16'd36187, 16'd65103, 16'd36352, 16'd9902, 16'd52285, 16'd40581, 16'd57023, 16'd43627, 16'd34072, 16'd20610, 16'd43387, 16'd56924, 16'd51163, 16'd64082, 16'd51883, 16'd60133, 16'd11161, 16'd53219, 16'd31605, 16'd21033, 16'd49798, 16'd21841, 16'd14863, 16'd28832, 16'd15691});
	test_expansion(128'h8057467cae702eecfc1ff99e36dbe5bd, {16'd7720, 16'd29771, 16'd16453, 16'd9997, 16'd37276, 16'd57625, 16'd18092, 16'd33380, 16'd63611, 16'd9603, 16'd13272, 16'd56559, 16'd55243, 16'd47395, 16'd6647, 16'd56366, 16'd38855, 16'd21142, 16'd32940, 16'd35848, 16'd26031, 16'd22099, 16'd3471, 16'd30732, 16'd7090, 16'd1108});
	test_expansion(128'h9d41a74d04a369be4c30881633c2ffeb, {16'd22477, 16'd28693, 16'd42959, 16'd62119, 16'd21546, 16'd34523, 16'd65323, 16'd32486, 16'd15065, 16'd17512, 16'd30467, 16'd1254, 16'd52363, 16'd28966, 16'd12678, 16'd33208, 16'd1401, 16'd17632, 16'd18168, 16'd2641, 16'd23582, 16'd25406, 16'd34023, 16'd47477, 16'd12126, 16'd21940});
	test_expansion(128'h75700b4e9f744ae33d24cb80557076cb, {16'd9771, 16'd47706, 16'd28299, 16'd59658, 16'd60340, 16'd3023, 16'd52476, 16'd20292, 16'd16966, 16'd43405, 16'd6943, 16'd51956, 16'd16989, 16'd12792, 16'd28847, 16'd32738, 16'd53252, 16'd25714, 16'd9646, 16'd22262, 16'd22480, 16'd36196, 16'd62224, 16'd34544, 16'd62228, 16'd16355});
	test_expansion(128'h284fddf99a679385d181bc1b39627701, {16'd41263, 16'd58855, 16'd2678, 16'd57997, 16'd51353, 16'd10566, 16'd53841, 16'd6934, 16'd42977, 16'd65517, 16'd55863, 16'd46890, 16'd5838, 16'd60044, 16'd9895, 16'd2558, 16'd59345, 16'd47335, 16'd21863, 16'd29696, 16'd18087, 16'd6566, 16'd63691, 16'd41218, 16'd43396, 16'd23651});
	test_expansion(128'h07f1149f5468c6fec3fd65c69a434b8e, {16'd5464, 16'd21006, 16'd6039, 16'd38841, 16'd32979, 16'd29066, 16'd26104, 16'd8399, 16'd49012, 16'd27971, 16'd50106, 16'd43938, 16'd2437, 16'd62378, 16'd23752, 16'd31127, 16'd45740, 16'd8006, 16'd37300, 16'd35352, 16'd37312, 16'd7035, 16'd26748, 16'd2787, 16'd9278, 16'd44525});
	test_expansion(128'h901bffaf8e97c064a10226fd758f6587, {16'd57982, 16'd56965, 16'd59898, 16'd59496, 16'd8146, 16'd25679, 16'd31858, 16'd52260, 16'd45781, 16'd24059, 16'd49290, 16'd52600, 16'd35769, 16'd46526, 16'd32652, 16'd55325, 16'd50156, 16'd43770, 16'd36773, 16'd39020, 16'd21855, 16'd1871, 16'd13827, 16'd43331, 16'd51534, 16'd20427});
	test_expansion(128'h00e3ed51f7eba5d4c4f5d3dd0c3eaf3b, {16'd48911, 16'd32587, 16'd42913, 16'd39022, 16'd36938, 16'd31077, 16'd22285, 16'd1892, 16'd1956, 16'd40360, 16'd35577, 16'd10964, 16'd44333, 16'd31925, 16'd18289, 16'd52467, 16'd54559, 16'd63805, 16'd15196, 16'd32582, 16'd21671, 16'd25647, 16'd45665, 16'd50369, 16'd23005, 16'd36618});
	test_expansion(128'h4f424ec073b7a4389a9a5854e118b9eb, {16'd32238, 16'd9739, 16'd23273, 16'd45293, 16'd17096, 16'd17251, 16'd47176, 16'd40781, 16'd8928, 16'd16238, 16'd9113, 16'd1089, 16'd15072, 16'd13416, 16'd21671, 16'd19807, 16'd14670, 16'd52747, 16'd1179, 16'd57212, 16'd15908, 16'd61905, 16'd31643, 16'd61357, 16'd22095, 16'd53891});
	test_expansion(128'h5785a47b33db14ee41e629afd17787ce, {16'd19975, 16'd43987, 16'd8981, 16'd3768, 16'd65206, 16'd22511, 16'd52552, 16'd42668, 16'd8194, 16'd37946, 16'd14955, 16'd2212, 16'd6556, 16'd18831, 16'd37392, 16'd46728, 16'd13670, 16'd21008, 16'd56356, 16'd38409, 16'd60064, 16'd42872, 16'd54540, 16'd5015, 16'd7033, 16'd65311});
	test_expansion(128'h07e0a872f017a9d9641765add6b7ac8c, {16'd8321, 16'd32609, 16'd13794, 16'd4395, 16'd51513, 16'd30677, 16'd7799, 16'd4146, 16'd8424, 16'd14772, 16'd53164, 16'd19178, 16'd12693, 16'd27997, 16'd26913, 16'd6362, 16'd54691, 16'd30835, 16'd51525, 16'd34618, 16'd14395, 16'd7649, 16'd2567, 16'd14537, 16'd51900, 16'd8691});
	test_expansion(128'hf325d771660fdb484f430ba2129e225a, {16'd16687, 16'd61127, 16'd16181, 16'd54517, 16'd38744, 16'd10999, 16'd60348, 16'd1312, 16'd52916, 16'd19505, 16'd46942, 16'd47937, 16'd26197, 16'd3824, 16'd19505, 16'd50851, 16'd48925, 16'd63677, 16'd924, 16'd18634, 16'd37379, 16'd2614, 16'd5612, 16'd40697, 16'd40963, 16'd50778});
	test_expansion(128'hff2c0854601bff4dd7d995e76a3db103, {16'd19556, 16'd14211, 16'd56951, 16'd30063, 16'd14920, 16'd54477, 16'd37203, 16'd1542, 16'd57481, 16'd57242, 16'd63460, 16'd52932, 16'd33299, 16'd63830, 16'd44523, 16'd23813, 16'd28760, 16'd55687, 16'd18853, 16'd46036, 16'd9387, 16'd4507, 16'd4359, 16'd28179, 16'd20698, 16'd37572});
	test_expansion(128'h99ec59d83f4aeb23cf54c2995fb13b12, {16'd58732, 16'd35923, 16'd28947, 16'd52522, 16'd36946, 16'd40489, 16'd63513, 16'd22226, 16'd60334, 16'd19655, 16'd62833, 16'd44454, 16'd39007, 16'd59975, 16'd59170, 16'd8408, 16'd2654, 16'd14673, 16'd9912, 16'd12682, 16'd55573, 16'd14006, 16'd43914, 16'd52307, 16'd44474, 16'd29718});
	test_expansion(128'h97fb2eebefe175052773882150fcd35c, {16'd3360, 16'd54298, 16'd5600, 16'd19446, 16'd19136, 16'd7005, 16'd11852, 16'd43320, 16'd7348, 16'd43186, 16'd49715, 16'd11569, 16'd59963, 16'd20732, 16'd54727, 16'd1693, 16'd16918, 16'd23257, 16'd39837, 16'd32627, 16'd53277, 16'd50442, 16'd138, 16'd54291, 16'd19258, 16'd64575});
	test_expansion(128'hb21e1e5c0e5e636d2888a2a62b6d1a9e, {16'd44661, 16'd22902, 16'd61571, 16'd19846, 16'd15996, 16'd7466, 16'd1806, 16'd27161, 16'd5213, 16'd33719, 16'd23577, 16'd13120, 16'd8957, 16'd63658, 16'd64171, 16'd4980, 16'd11038, 16'd61509, 16'd56992, 16'd549, 16'd56587, 16'd4346, 16'd17954, 16'd3516, 16'd26026, 16'd17341});
	test_expansion(128'he72ad91dd531889edbfc3c0ca33965b0, {16'd39555, 16'd16899, 16'd23024, 16'd37901, 16'd5403, 16'd44759, 16'd8808, 16'd64101, 16'd43150, 16'd9953, 16'd1052, 16'd56535, 16'd9602, 16'd33064, 16'd11959, 16'd17634, 16'd61886, 16'd14500, 16'd3815, 16'd16569, 16'd40975, 16'd13683, 16'd12619, 16'd49065, 16'd48373, 16'd38900});
	test_expansion(128'h242142768a7464a686915e79cfa2e225, {16'd64641, 16'd12031, 16'd62221, 16'd22284, 16'd54295, 16'd34925, 16'd48333, 16'd40089, 16'd57677, 16'd17890, 16'd57928, 16'd29139, 16'd64460, 16'd24588, 16'd983, 16'd55884, 16'd34076, 16'd18481, 16'd16909, 16'd12272, 16'd57277, 16'd21312, 16'd33229, 16'd23764, 16'd48855, 16'd55726});
	test_expansion(128'ha052632c66ace5093b56a6e42e6f9b0d, {16'd43355, 16'd25617, 16'd12755, 16'd35641, 16'd61687, 16'd6134, 16'd27364, 16'd44449, 16'd36114, 16'd42848, 16'd62101, 16'd39961, 16'd40153, 16'd48199, 16'd52859, 16'd15917, 16'd21622, 16'd18296, 16'd7376, 16'd8455, 16'd25583, 16'd28611, 16'd44758, 16'd55710, 16'd33691, 16'd25317});
	test_expansion(128'h002c836d5ac49e6a609632bd37dc0fa7, {16'd56548, 16'd59178, 16'd56203, 16'd8222, 16'd28870, 16'd24446, 16'd17190, 16'd52103, 16'd36175, 16'd47193, 16'd30000, 16'd2719, 16'd39635, 16'd5368, 16'd37272, 16'd59599, 16'd53220, 16'd9056, 16'd46670, 16'd43805, 16'd6034, 16'd24505, 16'd65526, 16'd53680, 16'd41493, 16'd62873});
	test_expansion(128'h23c252455dfad2893a9bc7c02d3d54af, {16'd62986, 16'd52551, 16'd43292, 16'd11311, 16'd20137, 16'd50164, 16'd15575, 16'd48812, 16'd40598, 16'd26545, 16'd19010, 16'd37987, 16'd62174, 16'd33052, 16'd37775, 16'd50234, 16'd61162, 16'd47761, 16'd2763, 16'd56684, 16'd5911, 16'd5148, 16'd44727, 16'd43089, 16'd3544, 16'd22672});
	test_expansion(128'h8d86513ef692309dc5122ebcc5b9f269, {16'd5658, 16'd52736, 16'd24554, 16'd8871, 16'd37462, 16'd45787, 16'd63304, 16'd21903, 16'd36067, 16'd43727, 16'd8934, 16'd17017, 16'd32651, 16'd19577, 16'd18863, 16'd47143, 16'd55936, 16'd7087, 16'd53750, 16'd60664, 16'd3534, 16'd39235, 16'd59002, 16'd40803, 16'd26039, 16'd46651});
	test_expansion(128'h3c42b96abf143c012741f3a510066b2c, {16'd7076, 16'd29299, 16'd57203, 16'd5974, 16'd38074, 16'd40612, 16'd19974, 16'd44892, 16'd29614, 16'd14473, 16'd41192, 16'd30618, 16'd6400, 16'd21764, 16'd3367, 16'd38438, 16'd65363, 16'd29229, 16'd2050, 16'd25515, 16'd11578, 16'd47490, 16'd17684, 16'd60127, 16'd54348, 16'd15428});
	test_expansion(128'ha7087ad2ff903a35fd3610cc59431962, {16'd40786, 16'd27024, 16'd31521, 16'd50653, 16'd8761, 16'd28854, 16'd39689, 16'd51163, 16'd47184, 16'd13171, 16'd50138, 16'd35989, 16'd38433, 16'd28020, 16'd49758, 16'd30677, 16'd65298, 16'd60344, 16'd53873, 16'd35280, 16'd11851, 16'd62283, 16'd33303, 16'd35170, 16'd22708, 16'd34534});
	test_expansion(128'he745d6f3bc6a0eca329f460165b67dc8, {16'd51249, 16'd24241, 16'd41116, 16'd45968, 16'd41292, 16'd47616, 16'd62210, 16'd16015, 16'd18334, 16'd3476, 16'd52809, 16'd5712, 16'd30950, 16'd58372, 16'd26863, 16'd9076, 16'd26153, 16'd51483, 16'd16898, 16'd63449, 16'd10056, 16'd40044, 16'd48120, 16'd2020, 16'd62773, 16'd44967});
	test_expansion(128'h031409ef9015ee8c5a9db57d8a0b687c, {16'd31796, 16'd24667, 16'd61636, 16'd62575, 16'd50587, 16'd56175, 16'd47909, 16'd60092, 16'd63836, 16'd10630, 16'd42704, 16'd30647, 16'd42371, 16'd48931, 16'd1151, 16'd20783, 16'd48136, 16'd20457, 16'd29144, 16'd1176, 16'd18692, 16'd33184, 16'd55417, 16'd48594, 16'd53830, 16'd31110});
	test_expansion(128'h8b013223a33ef6c6a80b42141180d517, {16'd17066, 16'd7086, 16'd65151, 16'd19688, 16'd22052, 16'd13336, 16'd47341, 16'd5375, 16'd58218, 16'd18021, 16'd46718, 16'd55636, 16'd25587, 16'd31105, 16'd24994, 16'd57982, 16'd33597, 16'd53771, 16'd26222, 16'd10921, 16'd23712, 16'd54310, 16'd11689, 16'd16018, 16'd42344, 16'd25495});
	test_expansion(128'hed350a84f00c04318e84f4c35aecc0bb, {16'd58158, 16'd48330, 16'd49298, 16'd25805, 16'd49870, 16'd38314, 16'd3144, 16'd20030, 16'd4497, 16'd50740, 16'd54810, 16'd33120, 16'd62410, 16'd45409, 16'd7726, 16'd46905, 16'd30398, 16'd15592, 16'd26616, 16'd29113, 16'd9418, 16'd41935, 16'd12985, 16'd1651, 16'd56486, 16'd34205});
	test_expansion(128'h6a948ee7da74ccd8cffe946c008116fd, {16'd36308, 16'd17481, 16'd44702, 16'd14306, 16'd23827, 16'd3229, 16'd34497, 16'd52578, 16'd23913, 16'd22243, 16'd35254, 16'd26741, 16'd43468, 16'd19099, 16'd13264, 16'd6421, 16'd11739, 16'd50941, 16'd59001, 16'd54999, 16'd59978, 16'd34286, 16'd31966, 16'd37498, 16'd54066, 16'd41455});
	test_expansion(128'h000e97a390baecb7ec6fc782c5dbbbd4, {16'd41074, 16'd55203, 16'd56120, 16'd26665, 16'd26929, 16'd60586, 16'd33580, 16'd53995, 16'd240, 16'd2179, 16'd40361, 16'd22666, 16'd33013, 16'd35139, 16'd29978, 16'd7244, 16'd61811, 16'd25544, 16'd22692, 16'd50404, 16'd7098, 16'd2479, 16'd39863, 16'd57706, 16'd36855, 16'd42748});
	test_expansion(128'h9617bae31d7deb2c434d168a432c8de2, {16'd31244, 16'd7212, 16'd47368, 16'd5910, 16'd15448, 16'd45785, 16'd25186, 16'd58975, 16'd26218, 16'd50518, 16'd14432, 16'd13407, 16'd48802, 16'd11406, 16'd60648, 16'd17935, 16'd60431, 16'd25385, 16'd27372, 16'd24928, 16'd32652, 16'd7087, 16'd47635, 16'd16580, 16'd45431, 16'd50677});
	test_expansion(128'h0e5cf4be10e2de6567466ec97e2c5d3c, {16'd8281, 16'd58913, 16'd63656, 16'd13686, 16'd5158, 16'd43278, 16'd52876, 16'd24651, 16'd2740, 16'd7926, 16'd64926, 16'd33558, 16'd59455, 16'd13100, 16'd44137, 16'd15542, 16'd40456, 16'd19080, 16'd35390, 16'd41032, 16'd44720, 16'd11459, 16'd63366, 16'd58380, 16'd28536, 16'd12254});
	test_expansion(128'h7e17ee66d9dba602cc915ab191cac01e, {16'd53745, 16'd52484, 16'd58529, 16'd533, 16'd37155, 16'd3436, 16'd29759, 16'd35371, 16'd19418, 16'd18313, 16'd31710, 16'd34048, 16'd2136, 16'd5737, 16'd13226, 16'd8371, 16'd8782, 16'd30256, 16'd11921, 16'd62181, 16'd32228, 16'd14550, 16'd65205, 16'd30353, 16'd14499, 16'd12763});
	test_expansion(128'he43561b67d27d56fce8580bc051a7fe9, {16'd40423, 16'd31547, 16'd27337, 16'd7140, 16'd37556, 16'd52469, 16'd3450, 16'd47001, 16'd52050, 16'd25323, 16'd46397, 16'd43788, 16'd15275, 16'd31318, 16'd9079, 16'd47113, 16'd51142, 16'd52716, 16'd3560, 16'd1233, 16'd34083, 16'd11388, 16'd40244, 16'd59560, 16'd36316, 16'd12044});
	test_expansion(128'ha8ab368f74882cbc18a3bf8a89698c45, {16'd42662, 16'd10139, 16'd65038, 16'd71, 16'd40167, 16'd49535, 16'd37756, 16'd14642, 16'd29525, 16'd47830, 16'd2546, 16'd56102, 16'd6960, 16'd60823, 16'd15183, 16'd55153, 16'd10848, 16'd30822, 16'd4410, 16'd61538, 16'd6050, 16'd25286, 16'd40463, 16'd82, 16'd62718, 16'd5415});
	test_expansion(128'h62a33676978bc6278cb92e5aec34aab4, {16'd28415, 16'd60218, 16'd51772, 16'd29609, 16'd4017, 16'd5814, 16'd62198, 16'd8526, 16'd41439, 16'd26257, 16'd17987, 16'd23562, 16'd59887, 16'd29031, 16'd3799, 16'd62693, 16'd26158, 16'd5668, 16'd30155, 16'd39160, 16'd35946, 16'd2794, 16'd14260, 16'd1793, 16'd64513, 16'd29037});
	test_expansion(128'heb55a106ce31b441e6944b2cb6fa2958, {16'd24287, 16'd19279, 16'd26631, 16'd56861, 16'd57633, 16'd38615, 16'd32291, 16'd41903, 16'd38486, 16'd8979, 16'd47587, 16'd38341, 16'd56330, 16'd61190, 16'd61108, 16'd44711, 16'd8387, 16'd55660, 16'd29393, 16'd6164, 16'd57830, 16'd31444, 16'd5042, 16'd18867, 16'd31839, 16'd59959});
	test_expansion(128'h45fc12ce34e0801fa61f87cb547266c5, {16'd56341, 16'd22514, 16'd22718, 16'd33164, 16'd36892, 16'd35826, 16'd50604, 16'd48936, 16'd43704, 16'd15631, 16'd31586, 16'd44101, 16'd37243, 16'd44292, 16'd35350, 16'd49653, 16'd30814, 16'd38805, 16'd38593, 16'd30332, 16'd18016, 16'd65095, 16'd7504, 16'd57109, 16'd35753, 16'd22504});
	test_expansion(128'hcacbecd4f3727fe7c4606dab33b81e1b, {16'd24605, 16'd64158, 16'd32100, 16'd21300, 16'd38454, 16'd62747, 16'd64434, 16'd15528, 16'd15810, 16'd11090, 16'd28484, 16'd65322, 16'd40274, 16'd6948, 16'd62479, 16'd60612, 16'd33967, 16'd10804, 16'd7329, 16'd10987, 16'd21249, 16'd44428, 16'd30034, 16'd18731, 16'd40447, 16'd36585});
	test_expansion(128'h216455b7d0e43619be19bde647610146, {16'd47159, 16'd47595, 16'd56917, 16'd15, 16'd62253, 16'd43578, 16'd19368, 16'd22064, 16'd59648, 16'd7836, 16'd35828, 16'd1890, 16'd35918, 16'd60384, 16'd10792, 16'd27980, 16'd50086, 16'd27602, 16'd42182, 16'd18752, 16'd44678, 16'd10274, 16'd43366, 16'd46388, 16'd12495, 16'd8558});
	test_expansion(128'h830e7215748b7517f0133005eb876ff5, {16'd49001, 16'd39618, 16'd11984, 16'd4514, 16'd34412, 16'd65014, 16'd56062, 16'd183, 16'd36305, 16'd45308, 16'd59771, 16'd59716, 16'd11373, 16'd21701, 16'd43556, 16'd5087, 16'd23831, 16'd32096, 16'd38324, 16'd44369, 16'd43739, 16'd34743, 16'd47067, 16'd52124, 16'd37831, 16'd22979});
	test_expansion(128'hc8fdc270a814e10c5516196a0b11e8db, {16'd32960, 16'd18617, 16'd54214, 16'd32588, 16'd57772, 16'd38689, 16'd10251, 16'd37282, 16'd21879, 16'd57, 16'd42611, 16'd17897, 16'd14871, 16'd35531, 16'd28130, 16'd1574, 16'd17578, 16'd9184, 16'd17543, 16'd19490, 16'd45180, 16'd18912, 16'd28254, 16'd8274, 16'd18107, 16'd16233});
	test_expansion(128'ha192c53413a52cc42fd21d5d87ce0f10, {16'd58429, 16'd12536, 16'd8361, 16'd58742, 16'd65372, 16'd17971, 16'd9718, 16'd60918, 16'd56899, 16'd4888, 16'd14071, 16'd53654, 16'd24857, 16'd11829, 16'd10337, 16'd11354, 16'd59767, 16'd53928, 16'd21771, 16'd22252, 16'd13180, 16'd42187, 16'd30685, 16'd1032, 16'd39138, 16'd15863});
	test_expansion(128'hc22c980cf037a4058c5b55e960d22271, {16'd43231, 16'd56374, 16'd23864, 16'd45434, 16'd43758, 16'd24600, 16'd33213, 16'd14936, 16'd55811, 16'd3637, 16'd19849, 16'd21075, 16'd26525, 16'd51655, 16'd3681, 16'd41696, 16'd10283, 16'd32978, 16'd55713, 16'd8031, 16'd53500, 16'd23020, 16'd11586, 16'd31565, 16'd32907, 16'd24200});
	test_expansion(128'h0d4814ccddf61a8ba2646ad2e7c7b24b, {16'd46999, 16'd32359, 16'd34812, 16'd37423, 16'd44325, 16'd19386, 16'd2747, 16'd31825, 16'd17367, 16'd33649, 16'd22434, 16'd30648, 16'd1324, 16'd4799, 16'd38606, 16'd6463, 16'd15230, 16'd19858, 16'd31238, 16'd61427, 16'd25375, 16'd23869, 16'd38706, 16'd21145, 16'd44870, 16'd2786});
	test_expansion(128'he260794751a7deafda0b6bc9e8c6a293, {16'd48498, 16'd43018, 16'd1059, 16'd56367, 16'd32779, 16'd20050, 16'd19653, 16'd44133, 16'd11873, 16'd53405, 16'd16204, 16'd25058, 16'd30714, 16'd40597, 16'd33043, 16'd50580, 16'd4314, 16'd10827, 16'd37296, 16'd19743, 16'd39280, 16'd38602, 16'd53422, 16'd62555, 16'd48938, 16'd21662});
	test_expansion(128'heabe64dfa59cbb7e10ca8ca36dbb0e71, {16'd905, 16'd49305, 16'd44087, 16'd51932, 16'd1070, 16'd23672, 16'd19788, 16'd57456, 16'd26479, 16'd2671, 16'd35901, 16'd36935, 16'd49140, 16'd23162, 16'd19208, 16'd2258, 16'd48370, 16'd37988, 16'd42373, 16'd36364, 16'd17475, 16'd47727, 16'd47007, 16'd1894, 16'd31046, 16'd39939});
	test_expansion(128'h3351528d9b2bce20b78da193850a7350, {16'd13154, 16'd46470, 16'd2060, 16'd45522, 16'd40401, 16'd52817, 16'd52272, 16'd43214, 16'd58966, 16'd29375, 16'd52286, 16'd30364, 16'd41152, 16'd45371, 16'd40644, 16'd26939, 16'd44704, 16'd44427, 16'd2010, 16'd21464, 16'd65291, 16'd1336, 16'd2923, 16'd12032, 16'd37933, 16'd145});
	test_expansion(128'h22c0b5a8586d9636f9a824c81fabc926, {16'd37067, 16'd38697, 16'd13209, 16'd51946, 16'd43981, 16'd44113, 16'd31728, 16'd7981, 16'd17423, 16'd60595, 16'd53706, 16'd29010, 16'd7781, 16'd46767, 16'd281, 16'd45854, 16'd59969, 16'd43589, 16'd52980, 16'd23717, 16'd65215, 16'd44637, 16'd1972, 16'd21599, 16'd23326, 16'd22826});
	test_expansion(128'hca80df2afc5b2401eb31be27d65b8229, {16'd1345, 16'd31662, 16'd15536, 16'd22160, 16'd34317, 16'd51325, 16'd33399, 16'd43053, 16'd33826, 16'd47952, 16'd17362, 16'd35535, 16'd44904, 16'd58720, 16'd31272, 16'd54269, 16'd22612, 16'd6312, 16'd8808, 16'd25929, 16'd40230, 16'd54830, 16'd12650, 16'd43317, 16'd9871, 16'd45885});
	test_expansion(128'h7ad6d9d954ad4d62367759da36c35381, {16'd10395, 16'd16203, 16'd16693, 16'd55886, 16'd24034, 16'd21155, 16'd19366, 16'd22543, 16'd17984, 16'd57732, 16'd53866, 16'd54723, 16'd5783, 16'd62001, 16'd31792, 16'd56357, 16'd28983, 16'd45787, 16'd7492, 16'd10446, 16'd42182, 16'd29975, 16'd51475, 16'd51138, 16'd46418, 16'd25209});
	test_expansion(128'h05affeaccf68fd213ecf47a92820c9fb, {16'd14642, 16'd13627, 16'd2793, 16'd17746, 16'd14422, 16'd38425, 16'd59383, 16'd35920, 16'd431, 16'd6255, 16'd6622, 16'd7590, 16'd25331, 16'd19773, 16'd55264, 16'd50477, 16'd7265, 16'd12068, 16'd17985, 16'd32533, 16'd27314, 16'd56344, 16'd36399, 16'd8785, 16'd40785, 16'd32405});
	test_expansion(128'hab72031d60eef07a4153539c07d85eeb, {16'd44515, 16'd7664, 16'd19369, 16'd14931, 16'd17881, 16'd10667, 16'd6739, 16'd30508, 16'd35435, 16'd59092, 16'd13513, 16'd51516, 16'd34801, 16'd58910, 16'd5817, 16'd16439, 16'd50205, 16'd52532, 16'd50896, 16'd48058, 16'd65358, 16'd37075, 16'd11072, 16'd27936, 16'd12745, 16'd52646});
	test_expansion(128'h2b8fa691efcd71518c2f48057d06576f, {16'd13910, 16'd19586, 16'd3081, 16'd12353, 16'd58308, 16'd14339, 16'd56582, 16'd23363, 16'd15533, 16'd31098, 16'd35405, 16'd22958, 16'd55518, 16'd3686, 16'd39454, 16'd25540, 16'd16400, 16'd25761, 16'd52535, 16'd6947, 16'd15571, 16'd33391, 16'd12438, 16'd990, 16'd16396, 16'd4845});
	test_expansion(128'h27ed04ffc9a521b03d5a4aed30b477a7, {16'd63587, 16'd47300, 16'd50485, 16'd39457, 16'd37605, 16'd56405, 16'd50623, 16'd23122, 16'd47899, 16'd48050, 16'd3153, 16'd47353, 16'd6708, 16'd44626, 16'd57129, 16'd42372, 16'd45282, 16'd40117, 16'd39480, 16'd59348, 16'd42761, 16'd18242, 16'd53844, 16'd15597, 16'd41494, 16'd36877});
	test_expansion(128'h5f415bfe45f57501c158ea28d445e7af, {16'd53178, 16'd15242, 16'd16253, 16'd3916, 16'd41025, 16'd37080, 16'd62914, 16'd52427, 16'd23750, 16'd46585, 16'd9243, 16'd16757, 16'd65057, 16'd48784, 16'd40710, 16'd44076, 16'd32946, 16'd63466, 16'd9840, 16'd52335, 16'd8871, 16'd59801, 16'd40800, 16'd52998, 16'd30028, 16'd7280});
	test_expansion(128'h6fc2a3f4d1604987aea429b82e48f86a, {16'd20580, 16'd11528, 16'd24585, 16'd45946, 16'd12587, 16'd50353, 16'd27775, 16'd13377, 16'd7023, 16'd4247, 16'd50055, 16'd24262, 16'd40090, 16'd23698, 16'd599, 16'd54242, 16'd14224, 16'd9123, 16'd27237, 16'd29665, 16'd41978, 16'd13261, 16'd16998, 16'd5199, 16'd10485, 16'd19675});
	test_expansion(128'h07f3c4cb94d6c58a8bf641420a75ad0b, {16'd20394, 16'd65238, 16'd51512, 16'd53862, 16'd16158, 16'd57288, 16'd35819, 16'd44616, 16'd14666, 16'd45472, 16'd29805, 16'd28821, 16'd64104, 16'd12804, 16'd51952, 16'd9543, 16'd53804, 16'd22192, 16'd64009, 16'd10724, 16'd60187, 16'd36972, 16'd1053, 16'd3653, 16'd21835, 16'd59926});
	test_expansion(128'h56225c40bcb19d0d5a2232d83e87fcd5, {16'd4992, 16'd63397, 16'd56505, 16'd40575, 16'd9468, 16'd59883, 16'd31062, 16'd61916, 16'd28741, 16'd51877, 16'd47149, 16'd45440, 16'd21554, 16'd18689, 16'd50793, 16'd58765, 16'd52224, 16'd24272, 16'd21600, 16'd1663, 16'd24436, 16'd46487, 16'd43861, 16'd59296, 16'd56574, 16'd52564});
	test_expansion(128'hf01fd62532a078b9c670317b1a19d976, {16'd8873, 16'd43153, 16'd47462, 16'd21533, 16'd20250, 16'd16851, 16'd15846, 16'd36534, 16'd15510, 16'd42663, 16'd48601, 16'd34193, 16'd20776, 16'd24004, 16'd63085, 16'd20855, 16'd21201, 16'd15071, 16'd4944, 16'd47001, 16'd43729, 16'd45182, 16'd52804, 16'd12437, 16'd31892, 16'd20757});
	test_expansion(128'h38bab8b1cc41d62f3d4cdbe2343ca9b9, {16'd2817, 16'd60478, 16'd31216, 16'd18821, 16'd57681, 16'd29029, 16'd43444, 16'd23484, 16'd41051, 16'd57304, 16'd54044, 16'd24924, 16'd6845, 16'd46228, 16'd15736, 16'd65345, 16'd6498, 16'd44314, 16'd38519, 16'd45407, 16'd61399, 16'd59355, 16'd63346, 16'd33734, 16'd18662, 16'd65506});
	test_expansion(128'h8f5cea95903923448b228e2f41b72ad4, {16'd5814, 16'd28702, 16'd42, 16'd51263, 16'd60442, 16'd8245, 16'd65217, 16'd28628, 16'd34414, 16'd1832, 16'd2688, 16'd20729, 16'd43527, 16'd37618, 16'd10874, 16'd43683, 16'd9056, 16'd5391, 16'd64968, 16'd4227, 16'd49964, 16'd30080, 16'd61149, 16'd30336, 16'd59971, 16'd17962});
	test_expansion(128'h8e38c60276e74143bc6ae9653418eba6, {16'd51447, 16'd57991, 16'd27185, 16'd53405, 16'd2096, 16'd12979, 16'd24067, 16'd12821, 16'd871, 16'd48804, 16'd27442, 16'd22826, 16'd39203, 16'd8301, 16'd6640, 16'd2777, 16'd19342, 16'd39275, 16'd55494, 16'd36883, 16'd8762, 16'd19175, 16'd7353, 16'd21232, 16'd58347, 16'd2658});
	test_expansion(128'h6e34fdc4cfbd9c96d29d148d74330788, {16'd6490, 16'd43979, 16'd64156, 16'd25189, 16'd59185, 16'd15654, 16'd54024, 16'd29640, 16'd8559, 16'd61748, 16'd22957, 16'd11679, 16'd58190, 16'd7455, 16'd56143, 16'd38878, 16'd40014, 16'd7231, 16'd34592, 16'd54410, 16'd1498, 16'd23104, 16'd14284, 16'd35678, 16'd31656, 16'd49033});
	test_expansion(128'he82725e294be00762e4cc3a03ec0fcce, {16'd30064, 16'd24437, 16'd60550, 16'd34589, 16'd2248, 16'd7980, 16'd52545, 16'd198, 16'd48431, 16'd46953, 16'd52235, 16'd45698, 16'd10352, 16'd53612, 16'd52104, 16'd36701, 16'd54564, 16'd54373, 16'd59353, 16'd12897, 16'd44303, 16'd5927, 16'd30758, 16'd58801, 16'd43953, 16'd48754});
	test_expansion(128'hf8ae765a141069ead9aa1e2630e4715b, {16'd8134, 16'd10177, 16'd24277, 16'd3034, 16'd34419, 16'd18032, 16'd1158, 16'd52425, 16'd33831, 16'd45182, 16'd38243, 16'd17934, 16'd31099, 16'd55232, 16'd57407, 16'd58766, 16'd61211, 16'd19138, 16'd18253, 16'd58165, 16'd1543, 16'd24907, 16'd25115, 16'd53404, 16'd40427, 16'd38131});
	test_expansion(128'h1c24627123a5339e490da883664832e5, {16'd63648, 16'd57773, 16'd44471, 16'd38186, 16'd51748, 16'd12256, 16'd55417, 16'd10424, 16'd43453, 16'd45151, 16'd59522, 16'd54838, 16'd37359, 16'd1448, 16'd162, 16'd36395, 16'd24121, 16'd125, 16'd48214, 16'd43194, 16'd12614, 16'd54177, 16'd31301, 16'd8280, 16'd26585, 16'd47512});
	test_expansion(128'h9d207c030e0d703deb93b6d38b43aaa2, {16'd43428, 16'd24769, 16'd41921, 16'd27063, 16'd40206, 16'd38361, 16'd16923, 16'd608, 16'd57885, 16'd23248, 16'd42570, 16'd47791, 16'd59848, 16'd28236, 16'd65061, 16'd59866, 16'd62610, 16'd34844, 16'd43229, 16'd32134, 16'd49727, 16'd47945, 16'd16735, 16'd41349, 16'd62319, 16'd52343});
	test_expansion(128'hf60d42b435fccbb6f6418879cde220cd, {16'd38026, 16'd37812, 16'd26160, 16'd28475, 16'd60999, 16'd52459, 16'd14396, 16'd17224, 16'd59262, 16'd39527, 16'd1319, 16'd14740, 16'd1861, 16'd17682, 16'd15507, 16'd25296, 16'd37390, 16'd25733, 16'd62750, 16'd24011, 16'd45548, 16'd22200, 16'd55549, 16'd8401, 16'd30424, 16'd63239});
	test_expansion(128'h40ef90729a02f1dc0727dd76969413f6, {16'd58737, 16'd13938, 16'd27980, 16'd56698, 16'd19290, 16'd55826, 16'd3738, 16'd18995, 16'd64318, 16'd19641, 16'd16943, 16'd52108, 16'd63720, 16'd49115, 16'd49247, 16'd12497, 16'd20092, 16'd30719, 16'd10282, 16'd44085, 16'd3895, 16'd41522, 16'd61043, 16'd35813, 16'd64567, 16'd42099});
	test_expansion(128'hbc0eacc180d6454d24d763b8ab27999b, {16'd41866, 16'd4147, 16'd28226, 16'd64183, 16'd26742, 16'd300, 16'd47704, 16'd12464, 16'd38772, 16'd20164, 16'd2103, 16'd30382, 16'd11338, 16'd9282, 16'd29731, 16'd31345, 16'd15424, 16'd27336, 16'd27232, 16'd62519, 16'd41284, 16'd40590, 16'd26686, 16'd40586, 16'd24031, 16'd35302});
	test_expansion(128'hc052f24566f5e76233791b816f01bb5a, {16'd32692, 16'd17643, 16'd36675, 16'd34391, 16'd58809, 16'd63606, 16'd5812, 16'd45246, 16'd11578, 16'd10950, 16'd7652, 16'd56107, 16'd45005, 16'd25722, 16'd42327, 16'd53751, 16'd56359, 16'd47804, 16'd8392, 16'd35925, 16'd59955, 16'd17967, 16'd63363, 16'd53844, 16'd1260, 16'd20800});
	test_expansion(128'hb68b01719d100dafb6c2b3e4ce7ef2c1, {16'd2459, 16'd17665, 16'd6528, 16'd14052, 16'd55577, 16'd51792, 16'd58378, 16'd15407, 16'd47885, 16'd64571, 16'd11047, 16'd6979, 16'd33986, 16'd121, 16'd47747, 16'd10728, 16'd49666, 16'd48994, 16'd10774, 16'd29380, 16'd23419, 16'd1563, 16'd14399, 16'd61624, 16'd382, 16'd2282});
	test_expansion(128'h9a9927b60e270cd5f5e406db283071d0, {16'd48296, 16'd2617, 16'd5514, 16'd27184, 16'd54195, 16'd33851, 16'd3369, 16'd33715, 16'd53438, 16'd64373, 16'd33753, 16'd12970, 16'd33177, 16'd45745, 16'd2100, 16'd22473, 16'd23879, 16'd64325, 16'd56140, 16'd64220, 16'd2370, 16'd32788, 16'd6612, 16'd19972, 16'd12086, 16'd21008});
	test_expansion(128'hdd2dd83a5de4ca7125adfc5bcc6c8664, {16'd42607, 16'd64372, 16'd49404, 16'd4754, 16'd55655, 16'd31018, 16'd50966, 16'd47446, 16'd6882, 16'd34885, 16'd19493, 16'd19769, 16'd40786, 16'd21493, 16'd60343, 16'd56026, 16'd63500, 16'd13121, 16'd35472, 16'd28712, 16'd46249, 16'd34205, 16'd54600, 16'd55700, 16'd40609, 16'd26185});
	test_expansion(128'hde7d378dd128c56ea9273d90443eaf93, {16'd55504, 16'd63853, 16'd46163, 16'd12745, 16'd20888, 16'd60924, 16'd33670, 16'd56282, 16'd4400, 16'd9164, 16'd28132, 16'd33743, 16'd21713, 16'd43912, 16'd10094, 16'd23640, 16'd54232, 16'd60830, 16'd56589, 16'd63144, 16'd45662, 16'd46552, 16'd17711, 16'd11018, 16'd44615, 16'd25566});
	test_expansion(128'h2b724727c73acf3c9e74053e79cbd6c3, {16'd33633, 16'd50463, 16'd35800, 16'd20827, 16'd42104, 16'd28121, 16'd15634, 16'd63261, 16'd2368, 16'd24030, 16'd64160, 16'd53323, 16'd17067, 16'd38737, 16'd12082, 16'd35709, 16'd51630, 16'd15911, 16'd48505, 16'd45614, 16'd36484, 16'd9952, 16'd47671, 16'd62674, 16'd51911, 16'd63871});
	test_expansion(128'h192c4df1d8ae8c998075b6ee453373a5, {16'd16095, 16'd24163, 16'd28569, 16'd6187, 16'd30249, 16'd33139, 16'd48303, 16'd14588, 16'd51828, 16'd37264, 16'd40736, 16'd39464, 16'd18168, 16'd24856, 16'd16342, 16'd28329, 16'd62452, 16'd23489, 16'd24652, 16'd31437, 16'd48622, 16'd55771, 16'd43875, 16'd22167, 16'd54332, 16'd34299});
	test_expansion(128'h677dde71ccf367167eecc0ea784aaa94, {16'd60801, 16'd12566, 16'd15892, 16'd46454, 16'd18450, 16'd36476, 16'd9318, 16'd44310, 16'd20200, 16'd2484, 16'd33439, 16'd50152, 16'd34010, 16'd3895, 16'd16550, 16'd38434, 16'd27758, 16'd52561, 16'd18888, 16'd11481, 16'd56975, 16'd30059, 16'd21284, 16'd35205, 16'd5485, 16'd54798});
	test_expansion(128'h16c85f0c2cd22238a159eaccb573a13d, {16'd45794, 16'd39654, 16'd55794, 16'd37246, 16'd25442, 16'd1551, 16'd30606, 16'd6176, 16'd45445, 16'd63955, 16'd21788, 16'd2190, 16'd28219, 16'd17005, 16'd65373, 16'd42881, 16'd44758, 16'd45366, 16'd61813, 16'd40082, 16'd5666, 16'd30781, 16'd39185, 16'd15137, 16'd64112, 16'd13878});
	test_expansion(128'h013c3df1b9f4c821fee094a009063621, {16'd47342, 16'd758, 16'd22049, 16'd19160, 16'd14375, 16'd35251, 16'd53556, 16'd12781, 16'd42235, 16'd23530, 16'd4906, 16'd58572, 16'd47963, 16'd40700, 16'd55567, 16'd26398, 16'd9649, 16'd16712, 16'd13390, 16'd31769, 16'd19754, 16'd39340, 16'd32945, 16'd41077, 16'd37667, 16'd15319});
	test_expansion(128'h167b5cbcd12958f4b65be62916bf0e57, {16'd48731, 16'd39463, 16'd10569, 16'd27624, 16'd55002, 16'd19545, 16'd55338, 16'd65128, 16'd58939, 16'd35215, 16'd58322, 16'd58700, 16'd11751, 16'd60937, 16'd16481, 16'd51391, 16'd59076, 16'd17039, 16'd11749, 16'd24074, 16'd31053, 16'd16457, 16'd44212, 16'd27598, 16'd16567, 16'd11674});
	test_expansion(128'h36effd7e1ad74c6378fcb085055c94d6, {16'd39778, 16'd32763, 16'd49184, 16'd21339, 16'd52068, 16'd30434, 16'd37504, 16'd56653, 16'd21581, 16'd15011, 16'd21067, 16'd58139, 16'd50324, 16'd963, 16'd19773, 16'd8042, 16'd30885, 16'd22390, 16'd6566, 16'd54171, 16'd49566, 16'd32127, 16'd8749, 16'd26604, 16'd45171, 16'd33678});
	test_expansion(128'hf6750e13661ab826de5fac1c5d782a9d, {16'd13330, 16'd44477, 16'd61138, 16'd35940, 16'd2143, 16'd27731, 16'd45912, 16'd37929, 16'd9455, 16'd23084, 16'd8248, 16'd16849, 16'd43425, 16'd52572, 16'd27316, 16'd45673, 16'd6799, 16'd5792, 16'd43105, 16'd46519, 16'd53491, 16'd41888, 16'd28365, 16'd22920, 16'd71, 16'd21705});
	test_expansion(128'h1e564cba021a204a91bc99bed8fa87e0, {16'd40908, 16'd27252, 16'd60953, 16'd21267, 16'd41421, 16'd59855, 16'd35673, 16'd16674, 16'd59574, 16'd9212, 16'd29621, 16'd3167, 16'd55392, 16'd4534, 16'd50868, 16'd5172, 16'd47241, 16'd45996, 16'd58342, 16'd128, 16'd60741, 16'd4053, 16'd49428, 16'd41888, 16'd12432, 16'd50474});
	test_expansion(128'h349543d705391e3a609f75431e92de37, {16'd34921, 16'd25725, 16'd6809, 16'd10321, 16'd16298, 16'd17098, 16'd18270, 16'd42451, 16'd61831, 16'd33236, 16'd21656, 16'd50876, 16'd47431, 16'd29236, 16'd40402, 16'd23755, 16'd44805, 16'd35872, 16'd44909, 16'd8684, 16'd39626, 16'd44205, 16'd64901, 16'd64277, 16'd58542, 16'd25218});
	test_expansion(128'h368adbeda85affe21cc21c369fdb8b35, {16'd6523, 16'd11809, 16'd5111, 16'd41939, 16'd57340, 16'd8883, 16'd61997, 16'd15482, 16'd4072, 16'd35757, 16'd21437, 16'd40432, 16'd9485, 16'd55367, 16'd4939, 16'd6072, 16'd62471, 16'd61284, 16'd34535, 16'd56336, 16'd60735, 16'd45947, 16'd52730, 16'd34630, 16'd17212, 16'd48480});
	test_expansion(128'h9cd935287223c4c1199bfbce565b3bce, {16'd10559, 16'd56973, 16'd1584, 16'd29260, 16'd2275, 16'd28896, 16'd58962, 16'd62687, 16'd48248, 16'd44556, 16'd1834, 16'd25687, 16'd8980, 16'd20421, 16'd27936, 16'd26447, 16'd63939, 16'd37563, 16'd23167, 16'd60015, 16'd11330, 16'd52731, 16'd39464, 16'd32941, 16'd21749, 16'd52121});
	test_expansion(128'hfa5370971e9199b8821f226d85b4506c, {16'd47341, 16'd9257, 16'd27199, 16'd17572, 16'd11027, 16'd11728, 16'd37893, 16'd27282, 16'd52264, 16'd47877, 16'd48654, 16'd62866, 16'd50150, 16'd58777, 16'd41533, 16'd62249, 16'd1047, 16'd33349, 16'd30566, 16'd5542, 16'd11362, 16'd1507, 16'd59600, 16'd39228, 16'd57324, 16'd44734});
	test_expansion(128'h198f542f43fc636100718ff44ae03b69, {16'd15078, 16'd44443, 16'd8368, 16'd45917, 16'd20334, 16'd16721, 16'd51096, 16'd31080, 16'd49423, 16'd11768, 16'd34672, 16'd1408, 16'd23871, 16'd12998, 16'd53804, 16'd4168, 16'd32607, 16'd382, 16'd64464, 16'd22104, 16'd29187, 16'd48585, 16'd37589, 16'd10082, 16'd18913, 16'd22352});
	test_expansion(128'h6264907a1dee40d2259c2c9830be66e2, {16'd63254, 16'd24046, 16'd60267, 16'd4117, 16'd21179, 16'd1790, 16'd56812, 16'd18973, 16'd1999, 16'd10582, 16'd28351, 16'd23828, 16'd52669, 16'd56551, 16'd61482, 16'd25251, 16'd3365, 16'd10064, 16'd62201, 16'd9449, 16'd50284, 16'd27603, 16'd33173, 16'd55036, 16'd38374, 16'd48181});
	test_expansion(128'h524624e1d0800cc16c928d07083b4367, {16'd60911, 16'd33365, 16'd21189, 16'd23762, 16'd34055, 16'd48639, 16'd24676, 16'd44919, 16'd30192, 16'd1924, 16'd1542, 16'd20139, 16'd7973, 16'd20001, 16'd11718, 16'd27646, 16'd33048, 16'd3730, 16'd48635, 16'd29794, 16'd44356, 16'd41900, 16'd54259, 16'd59238, 16'd15541, 16'd39566});
	test_expansion(128'hd0667bedfdb87f0045650820a2435a94, {16'd61387, 16'd37030, 16'd49765, 16'd3409, 16'd64267, 16'd27730, 16'd57878, 16'd62769, 16'd15188, 16'd64400, 16'd6886, 16'd9351, 16'd52427, 16'd5700, 16'd38451, 16'd6902, 16'd20021, 16'd28499, 16'd44720, 16'd16609, 16'd20551, 16'd21999, 16'd43435, 16'd43604, 16'd56199, 16'd14101});
	test_expansion(128'h991477471ff9ca9c4db74e7d6ddaee50, {16'd12359, 16'd54035, 16'd30476, 16'd40111, 16'd13601, 16'd16768, 16'd31147, 16'd4873, 16'd28654, 16'd33209, 16'd13771, 16'd36036, 16'd28784, 16'd21846, 16'd55753, 16'd23845, 16'd39573, 16'd30782, 16'd3489, 16'd53050, 16'd9903, 16'd16911, 16'd39204, 16'd65376, 16'd51470, 16'd40130});
	test_expansion(128'h882004585d35cbee865ecea90592fc88, {16'd7066, 16'd20816, 16'd13259, 16'd47855, 16'd12879, 16'd14926, 16'd60936, 16'd25546, 16'd39771, 16'd37736, 16'd3104, 16'd40335, 16'd40081, 16'd56811, 16'd55701, 16'd32323, 16'd2056, 16'd7216, 16'd19276, 16'd36151, 16'd3536, 16'd29106, 16'd24052, 16'd35482, 16'd42146, 16'd55486});
	test_expansion(128'h76a1a8a9e4fc6850a499626adc8b637c, {16'd31058, 16'd20312, 16'd46399, 16'd28108, 16'd18309, 16'd10424, 16'd3583, 16'd32193, 16'd14184, 16'd424, 16'd50813, 16'd16163, 16'd15645, 16'd19774, 16'd5544, 16'd43475, 16'd61136, 16'd6933, 16'd42132, 16'd46690, 16'd53351, 16'd57171, 16'd10055, 16'd64891, 16'd3674, 16'd32350});
	test_expansion(128'he9072e06769fe6f6275ba5c61a62af75, {16'd48111, 16'd12908, 16'd49481, 16'd59200, 16'd18609, 16'd32584, 16'd46330, 16'd60592, 16'd47813, 16'd17693, 16'd49229, 16'd55391, 16'd64863, 16'd8172, 16'd31121, 16'd50287, 16'd8269, 16'd49936, 16'd7574, 16'd56901, 16'd38703, 16'd36030, 16'd45098, 16'd21334, 16'd13446, 16'd59732});
	test_expansion(128'hfd7279d010e3d8147aaa3c7b5aa36af2, {16'd45410, 16'd42839, 16'd23480, 16'd25708, 16'd15176, 16'd33015, 16'd48453, 16'd8862, 16'd48634, 16'd45190, 16'd61568, 16'd40588, 16'd59345, 16'd2106, 16'd15601, 16'd26452, 16'd5182, 16'd25649, 16'd43962, 16'd10087, 16'd19262, 16'd57495, 16'd57177, 16'd54941, 16'd8671, 16'd58700});
	test_expansion(128'hd83181bf4714fb1da64c5250355f3cf0, {16'd60304, 16'd64229, 16'd53056, 16'd31549, 16'd7709, 16'd23097, 16'd6150, 16'd34666, 16'd10281, 16'd59296, 16'd61171, 16'd12640, 16'd42407, 16'd49634, 16'd11022, 16'd53634, 16'd47037, 16'd16305, 16'd40978, 16'd43857, 16'd30140, 16'd30812, 16'd6884, 16'd52972, 16'd24699, 16'd24881});
	test_expansion(128'h5ccddf4f613c0ae81f460cddc0822753, {16'd59552, 16'd23249, 16'd56258, 16'd41663, 16'd31076, 16'd51860, 16'd34657, 16'd55353, 16'd47414, 16'd25330, 16'd34918, 16'd56277, 16'd35312, 16'd25974, 16'd57414, 16'd61117, 16'd35582, 16'd50707, 16'd53176, 16'd28071, 16'd15814, 16'd60698, 16'd41660, 16'd33875, 16'd28623, 16'd51308});
	test_expansion(128'h5b1638d03e5d11f9e5107b8d98b7c7cc, {16'd11796, 16'd58772, 16'd59444, 16'd16527, 16'd90, 16'd31973, 16'd47362, 16'd37970, 16'd39001, 16'd37343, 16'd20744, 16'd62513, 16'd42758, 16'd289, 16'd62770, 16'd59627, 16'd16347, 16'd22279, 16'd38472, 16'd59164, 16'd47719, 16'd4351, 16'd57282, 16'd60589, 16'd2957, 16'd33949});
	test_expansion(128'hf2919da02ed99934f74975cbc62c0b8b, {16'd62635, 16'd40232, 16'd9461, 16'd11983, 16'd47422, 16'd10586, 16'd49353, 16'd50786, 16'd29831, 16'd9679, 16'd54721, 16'd52039, 16'd22139, 16'd55783, 16'd64575, 16'd25299, 16'd52186, 16'd1468, 16'd56096, 16'd59281, 16'd2413, 16'd51208, 16'd39154, 16'd48470, 16'd62993, 16'd46155});
	test_expansion(128'h27841dae3c3674d494afd19a0e5700a6, {16'd1890, 16'd23868, 16'd61974, 16'd40157, 16'd55536, 16'd56965, 16'd22873, 16'd20843, 16'd51779, 16'd31480, 16'd16680, 16'd3095, 16'd6054, 16'd46159, 16'd33860, 16'd51565, 16'd2795, 16'd6870, 16'd5543, 16'd24481, 16'd23234, 16'd49958, 16'd19001, 16'd18975, 16'd57144, 16'd16145});
	test_expansion(128'hdeab7cd63071fb45cbbf917850ed3920, {16'd35470, 16'd38055, 16'd27147, 16'd54994, 16'd62827, 16'd32759, 16'd63466, 16'd59675, 16'd5446, 16'd63363, 16'd36417, 16'd17337, 16'd30307, 16'd23676, 16'd12930, 16'd22896, 16'd56992, 16'd59192, 16'd5357, 16'd5304, 16'd31923, 16'd65369, 16'd27438, 16'd59718, 16'd29848, 16'd52550});
	test_expansion(128'hff1604cea4b1fccc99d49a7972206866, {16'd42849, 16'd40644, 16'd54896, 16'd8987, 16'd31760, 16'd9202, 16'd3850, 16'd61164, 16'd41374, 16'd16231, 16'd1982, 16'd54877, 16'd12041, 16'd30681, 16'd2507, 16'd34020, 16'd3378, 16'd39403, 16'd4531, 16'd61142, 16'd13039, 16'd2542, 16'd31505, 16'd47204, 16'd63697, 16'd25158});
	test_expansion(128'h943907e90f45f06e94a2556a2751e259, {16'd28549, 16'd39435, 16'd4473, 16'd11839, 16'd34938, 16'd29262, 16'd30040, 16'd13718, 16'd59228, 16'd53161, 16'd31210, 16'd37422, 16'd42496, 16'd32865, 16'd53842, 16'd54860, 16'd16299, 16'd27090, 16'd58992, 16'd31325, 16'd51477, 16'd9203, 16'd49390, 16'd64206, 16'd14586, 16'd10464});
	test_expansion(128'h447671d2e04920586bfbb925840142e1, {16'd34140, 16'd15988, 16'd63877, 16'd33884, 16'd17085, 16'd56489, 16'd33641, 16'd58976, 16'd6357, 16'd30580, 16'd10380, 16'd44422, 16'd24269, 16'd54738, 16'd30503, 16'd20434, 16'd16742, 16'd28503, 16'd5696, 16'd16546, 16'd42993, 16'd43364, 16'd10053, 16'd19473, 16'd62283, 16'd55150});
	test_expansion(128'hb80f5ec2a95f6b32af63770e84291208, {16'd6284, 16'd3549, 16'd62809, 16'd61285, 16'd40776, 16'd31080, 16'd53362, 16'd12802, 16'd61686, 16'd58361, 16'd35163, 16'd928, 16'd54794, 16'd851, 16'd55638, 16'd56495, 16'd59713, 16'd52098, 16'd22030, 16'd59256, 16'd53802, 16'd59702, 16'd40181, 16'd31149, 16'd54155, 16'd53869});
	test_expansion(128'h9144073cd44f0585298f5835050030ee, {16'd33444, 16'd15752, 16'd37228, 16'd47488, 16'd61047, 16'd11119, 16'd18985, 16'd1902, 16'd21113, 16'd30535, 16'd37909, 16'd58058, 16'd28170, 16'd39026, 16'd43890, 16'd39085, 16'd60405, 16'd53665, 16'd23544, 16'd37835, 16'd21916, 16'd59896, 16'd47699, 16'd48314, 16'd60081, 16'd63663});
	test_expansion(128'hae8c3feca4c81db9d22f1227d413bef2, {16'd55855, 16'd21713, 16'd3850, 16'd56854, 16'd43070, 16'd15011, 16'd63128, 16'd36032, 16'd54094, 16'd38334, 16'd55915, 16'd27948, 16'd9382, 16'd26144, 16'd27467, 16'd2862, 16'd38413, 16'd56688, 16'd54224, 16'd21279, 16'd65454, 16'd52439, 16'd50972, 16'd50971, 16'd59279, 16'd57589});
	test_expansion(128'h4a33c373375a7dfa57d7d83c537aa690, {16'd34966, 16'd34933, 16'd42844, 16'd51440, 16'd49613, 16'd53895, 16'd15612, 16'd3653, 16'd56917, 16'd55623, 16'd22363, 16'd11448, 16'd32243, 16'd60220, 16'd26576, 16'd13462, 16'd30149, 16'd43538, 16'd26583, 16'd18726, 16'd51842, 16'd44053, 16'd12574, 16'd25937, 16'd65501, 16'd58128});
	test_expansion(128'hd45a9b2bc5cd3ea6659165c976a8a923, {16'd35009, 16'd45731, 16'd50229, 16'd22156, 16'd51500, 16'd55062, 16'd47184, 16'd4756, 16'd46553, 16'd46138, 16'd9391, 16'd43897, 16'd42577, 16'd2476, 16'd12265, 16'd15674, 16'd26014, 16'd28340, 16'd17346, 16'd44763, 16'd36302, 16'd9913, 16'd4883, 16'd55114, 16'd10958, 16'd65387});
	test_expansion(128'hee5355c00c4a10625a33f51840b246c4, {16'd24642, 16'd40354, 16'd47076, 16'd31787, 16'd43948, 16'd11693, 16'd41054, 16'd44133, 16'd10731, 16'd54202, 16'd52305, 16'd56842, 16'd39969, 16'd9662, 16'd17234, 16'd51960, 16'd39044, 16'd57036, 16'd51879, 16'd14982, 16'd16812, 16'd17908, 16'd54276, 16'd29824, 16'd47415, 16'd57992});
	test_expansion(128'hb65430d978ac03995ff949880299c922, {16'd41131, 16'd4234, 16'd23191, 16'd30745, 16'd62185, 16'd17199, 16'd17520, 16'd64388, 16'd33724, 16'd24999, 16'd38256, 16'd6537, 16'd32011, 16'd33326, 16'd36129, 16'd21410, 16'd5779, 16'd39855, 16'd65111, 16'd59968, 16'd2118, 16'd60139, 16'd46779, 16'd21759, 16'd52016, 16'd6411});
	test_expansion(128'h8174b876dad17b0134832a46cc79d86b, {16'd41020, 16'd12516, 16'd39609, 16'd62376, 16'd46488, 16'd5463, 16'd9965, 16'd43130, 16'd64034, 16'd54306, 16'd33400, 16'd20945, 16'd53224, 16'd44110, 16'd875, 16'd65163, 16'd45111, 16'd40696, 16'd37456, 16'd15671, 16'd45768, 16'd34643, 16'd32394, 16'd60332, 16'd13016, 16'd21043});
	test_expansion(128'hc343916f19d1113e0d6d8a2e74068980, {16'd49563, 16'd39516, 16'd63614, 16'd40522, 16'd51822, 16'd50225, 16'd37497, 16'd4424, 16'd7656, 16'd6307, 16'd40227, 16'd18426, 16'd53498, 16'd22895, 16'd47668, 16'd21202, 16'd42283, 16'd61480, 16'd46082, 16'd56707, 16'd58136, 16'd31859, 16'd57959, 16'd47931, 16'd51329, 16'd10486});
	test_expansion(128'h9da5d1025c549543add593bdd1b2efcd, {16'd4111, 16'd38139, 16'd13699, 16'd8459, 16'd54454, 16'd14361, 16'd50497, 16'd28710, 16'd20507, 16'd49096, 16'd58996, 16'd8315, 16'd24756, 16'd48485, 16'd20119, 16'd10536, 16'd31348, 16'd60622, 16'd38338, 16'd27451, 16'd38498, 16'd13072, 16'd17545, 16'd33091, 16'd10615, 16'd2808});
	test_expansion(128'hd317249d414a82707c175e7a9502be7b, {16'd9030, 16'd56184, 16'd46579, 16'd43616, 16'd53914, 16'd44428, 16'd36918, 16'd53908, 16'd13005, 16'd46087, 16'd40656, 16'd3325, 16'd57370, 16'd13872, 16'd12447, 16'd5165, 16'd7467, 16'd12025, 16'd54131, 16'd13993, 16'd54459, 16'd47677, 16'd53754, 16'd1340, 16'd2198, 16'd8073});
	test_expansion(128'h8ed8e5e3c13231d8a081f27660f092b5, {16'd32810, 16'd51550, 16'd59536, 16'd55665, 16'd26916, 16'd26176, 16'd6913, 16'd42390, 16'd2113, 16'd57983, 16'd56217, 16'd17991, 16'd57361, 16'd23315, 16'd42579, 16'd29975, 16'd29415, 16'd17652, 16'd1801, 16'd11564, 16'd28298, 16'd51000, 16'd9050, 16'd3467, 16'd1580, 16'd28423});
	test_expansion(128'he8b561d3ec82f225fd55e334754f4ce0, {16'd22825, 16'd37670, 16'd18588, 16'd43973, 16'd37543, 16'd59995, 16'd24238, 16'd39366, 16'd676, 16'd52486, 16'd40928, 16'd39799, 16'd28366, 16'd49145, 16'd22404, 16'd60339, 16'd33929, 16'd11519, 16'd5296, 16'd56863, 16'd39248, 16'd54224, 16'd2564, 16'd40969, 16'd26143, 16'd12068});
	test_expansion(128'h5f5d85a8cec57605d7a0726e7fba5b7c, {16'd63949, 16'd19061, 16'd51154, 16'd55055, 16'd42803, 16'd47527, 16'd31233, 16'd9395, 16'd5111, 16'd60830, 16'd60406, 16'd15027, 16'd18323, 16'd32396, 16'd42862, 16'd50621, 16'd3433, 16'd53471, 16'd22218, 16'd40456, 16'd44332, 16'd33189, 16'd39069, 16'd526, 16'd39933, 16'd30064});
	test_expansion(128'h2989bc6765aba5f048a0b71329649947, {16'd25935, 16'd25955, 16'd4922, 16'd18835, 16'd43992, 16'd58927, 16'd24659, 16'd17305, 16'd65008, 16'd34163, 16'd5299, 16'd61511, 16'd53030, 16'd21745, 16'd12951, 16'd4963, 16'd20675, 16'd36991, 16'd2332, 16'd21909, 16'd36122, 16'd404, 16'd41665, 16'd19177, 16'd46016, 16'd31615});
	test_expansion(128'h1eb37067150d1ec96668f38c58ecf9b1, {16'd27200, 16'd59598, 16'd38089, 16'd27935, 16'd40948, 16'd1881, 16'd9263, 16'd31283, 16'd34142, 16'd63209, 16'd5413, 16'd8317, 16'd59511, 16'd58087, 16'd51166, 16'd3749, 16'd33111, 16'd792, 16'd42597, 16'd4351, 16'd44236, 16'd54973, 16'd24670, 16'd50922, 16'd43731, 16'd20755});
	test_expansion(128'h63a1e1f1595af73342a8137a9050c03a, {16'd55327, 16'd31226, 16'd39645, 16'd50068, 16'd751, 16'd39915, 16'd22048, 16'd15696, 16'd62195, 16'd11068, 16'd57018, 16'd61987, 16'd64918, 16'd32777, 16'd5125, 16'd3684, 16'd28940, 16'd14690, 16'd49469, 16'd55387, 16'd46700, 16'd3439, 16'd30329, 16'd62248, 16'd20277, 16'd62473});
	test_expansion(128'h758d90dcc4fee7a821aff67382f9ab48, {16'd51178, 16'd5207, 16'd61305, 16'd49476, 16'd8821, 16'd64906, 16'd53528, 16'd56856, 16'd63611, 16'd2837, 16'd8187, 16'd20225, 16'd14378, 16'd56260, 16'd20036, 16'd15190, 16'd33496, 16'd23068, 16'd50212, 16'd2125, 16'd38276, 16'd33730, 16'd7665, 16'd19891, 16'd52845, 16'd61886});
	test_expansion(128'hbcbebc9975155e716cad56f971f7e6c5, {16'd41993, 16'd27357, 16'd43620, 16'd5898, 16'd64469, 16'd38984, 16'd35887, 16'd15120, 16'd34515, 16'd37206, 16'd12754, 16'd2096, 16'd46995, 16'd60755, 16'd30186, 16'd36090, 16'd61986, 16'd52150, 16'd65279, 16'd59468, 16'd25762, 16'd5770, 16'd51373, 16'd22806, 16'd6629, 16'd9983});
	test_expansion(128'h3ea86ffadb2e48caad46396b5089f799, {16'd40403, 16'd1485, 16'd18280, 16'd27417, 16'd10950, 16'd303, 16'd32062, 16'd18639, 16'd14611, 16'd61229, 16'd22821, 16'd50436, 16'd38898, 16'd61843, 16'd22855, 16'd16253, 16'd27316, 16'd60210, 16'd11002, 16'd1608, 16'd61089, 16'd57347, 16'd13100, 16'd7950, 16'd59616, 16'd5506});
	test_expansion(128'h5947a35b879bcaed20f0654124ed3983, {16'd40658, 16'd1638, 16'd47273, 16'd22680, 16'd28166, 16'd29217, 16'd10251, 16'd41595, 16'd37307, 16'd6613, 16'd49627, 16'd56628, 16'd15350, 16'd3525, 16'd20401, 16'd54844, 16'd8507, 16'd61739, 16'd27796, 16'd47164, 16'd23213, 16'd2949, 16'd35754, 16'd43102, 16'd59784, 16'd59308});
	test_expansion(128'hb5baffd7e3b8fc2b6922760d8efcec3f, {16'd56227, 16'd48232, 16'd21436, 16'd64135, 16'd14962, 16'd23334, 16'd17604, 16'd26352, 16'd16137, 16'd4506, 16'd50432, 16'd54877, 16'd12243, 16'd31144, 16'd44442, 16'd54124, 16'd23084, 16'd62424, 16'd49468, 16'd23662, 16'd56056, 16'd1142, 16'd53028, 16'd24554, 16'd45874, 16'd3768});
	test_expansion(128'h1e904949d14bdce5cad4163e0a984ef5, {16'd3980, 16'd46828, 16'd55318, 16'd39726, 16'd28775, 16'd46934, 16'd53065, 16'd40773, 16'd6894, 16'd6863, 16'd61112, 16'd45707, 16'd42060, 16'd24345, 16'd24336, 16'd34763, 16'd25330, 16'd57689, 16'd42426, 16'd30133, 16'd35659, 16'd46669, 16'd4399, 16'd64973, 16'd14882, 16'd58380});
	test_expansion(128'h7bd9c0531d8c136fc8b4322882b045bc, {16'd29423, 16'd12579, 16'd64411, 16'd14752, 16'd21916, 16'd39232, 16'd3920, 16'd45499, 16'd945, 16'd30712, 16'd64060, 16'd19619, 16'd5862, 16'd33818, 16'd56115, 16'd30911, 16'd33666, 16'd22867, 16'd13586, 16'd55651, 16'd65108, 16'd12259, 16'd11301, 16'd26150, 16'd44085, 16'd42907});
	test_expansion(128'hedec6dbc08d238d86c7c0dc5785f670c, {16'd3395, 16'd61904, 16'd10310, 16'd11518, 16'd37172, 16'd54461, 16'd49590, 16'd8259, 16'd52991, 16'd64262, 16'd8731, 16'd8445, 16'd54375, 16'd65362, 16'd3080, 16'd40080, 16'd60652, 16'd34922, 16'd15579, 16'd9477, 16'd19860, 16'd33902, 16'd8719, 16'd28670, 16'd47302, 16'd19067});
	test_expansion(128'h6f295b3f77d27ca177a0ba9883891e4a, {16'd45985, 16'd53508, 16'd50654, 16'd57065, 16'd41651, 16'd44014, 16'd60123, 16'd45100, 16'd3549, 16'd6483, 16'd10164, 16'd50473, 16'd57202, 16'd51229, 16'd49580, 16'd64181, 16'd39948, 16'd13444, 16'd47656, 16'd31646, 16'd28050, 16'd12494, 16'd41787, 16'd1764, 16'd64475, 16'd10472});
	test_expansion(128'h6935b5e4444718dcd7699ac11b891ccd, {16'd63396, 16'd5471, 16'd9776, 16'd5578, 16'd6077, 16'd46382, 16'd12223, 16'd50047, 16'd30774, 16'd60073, 16'd19617, 16'd13413, 16'd10120, 16'd25283, 16'd33076, 16'd24644, 16'd40410, 16'd7607, 16'd61177, 16'd1693, 16'd17489, 16'd11689, 16'd34410, 16'd16586, 16'd20463, 16'd41840});
	test_expansion(128'hab544fb7a061c62bd788677b1a6d2129, {16'd17410, 16'd56682, 16'd62275, 16'd30057, 16'd20507, 16'd38339, 16'd8626, 16'd21860, 16'd36191, 16'd32239, 16'd59655, 16'd16218, 16'd11509, 16'd5936, 16'd53289, 16'd50598, 16'd2790, 16'd43160, 16'd57788, 16'd55310, 16'd59032, 16'd37516, 16'd258, 16'd21754, 16'd56286, 16'd35576});
	test_expansion(128'hcc0d5b98e71e0a23db97e896c3c56460, {16'd4042, 16'd25141, 16'd49329, 16'd64103, 16'd49645, 16'd6426, 16'd21086, 16'd15169, 16'd40719, 16'd50821, 16'd14606, 16'd15214, 16'd19659, 16'd6197, 16'd983, 16'd1121, 16'd38701, 16'd57261, 16'd6087, 16'd24567, 16'd21661, 16'd45791, 16'd52740, 16'd55377, 16'd20434, 16'd30729});
	test_expansion(128'h1cd8ce781d762319174e879358b2f51f, {16'd33253, 16'd52333, 16'd28784, 16'd11523, 16'd31632, 16'd43424, 16'd65447, 16'd53363, 16'd7787, 16'd47354, 16'd17352, 16'd64798, 16'd52712, 16'd28763, 16'd42376, 16'd45084, 16'd13242, 16'd64749, 16'd29897, 16'd31946, 16'd691, 16'd50372, 16'd47018, 16'd65377, 16'd12341, 16'd9753});
	test_expansion(128'hb0a4eeca5edb8fc754d9de396b59b692, {16'd45928, 16'd64761, 16'd33265, 16'd38107, 16'd53804, 16'd49893, 16'd56622, 16'd53307, 16'd3548, 16'd4164, 16'd60990, 16'd29292, 16'd21575, 16'd37207, 16'd58211, 16'd55758, 16'd7646, 16'd39539, 16'd47935, 16'd30324, 16'd62957, 16'd42369, 16'd15395, 16'd28805, 16'd19277, 16'd56237});
	test_expansion(128'h3714f2fd9028125ad75f0a03e3d4d05d, {16'd52726, 16'd14622, 16'd48186, 16'd10552, 16'd6330, 16'd28409, 16'd56499, 16'd46513, 16'd7785, 16'd17299, 16'd58856, 16'd11167, 16'd5514, 16'd50122, 16'd57810, 16'd15301, 16'd47882, 16'd38350, 16'd10460, 16'd14692, 16'd25057, 16'd8357, 16'd15170, 16'd39061, 16'd1048, 16'd7601});
	test_expansion(128'h7f90b9dae619689bc510ec71ee72c1e3, {16'd60548, 16'd28230, 16'd16894, 16'd57239, 16'd55487, 16'd48446, 16'd55295, 16'd60173, 16'd40555, 16'd7328, 16'd29601, 16'd45840, 16'd8171, 16'd43672, 16'd12025, 16'd26690, 16'd19746, 16'd12766, 16'd47391, 16'd50156, 16'd31053, 16'd28491, 16'd8382, 16'd43265, 16'd39555, 16'd18233});
	test_expansion(128'h00c3be8ef6957c81ea46e405518b095d, {16'd28128, 16'd62010, 16'd945, 16'd25225, 16'd49465, 16'd37171, 16'd27124, 16'd52438, 16'd42202, 16'd2962, 16'd11026, 16'd55277, 16'd42652, 16'd31394, 16'd29656, 16'd14088, 16'd42246, 16'd51035, 16'd21437, 16'd279, 16'd36426, 16'd25585, 16'd867, 16'd16597, 16'd1015, 16'd36077});
	test_expansion(128'hfb16ed88c5b383b97cb93aafc21e280f, {16'd21134, 16'd4623, 16'd56149, 16'd4945, 16'd42088, 16'd8360, 16'd40004, 16'd26177, 16'd58542, 16'd26954, 16'd29481, 16'd18023, 16'd50859, 16'd32833, 16'd43616, 16'd46023, 16'd43162, 16'd20700, 16'd29433, 16'd40116, 16'd38790, 16'd32698, 16'd40863, 16'd6179, 16'd37102, 16'd42413});
	test_expansion(128'h5b9f35acdfd7698628ccc9cdf326fe1b, {16'd54961, 16'd62772, 16'd14813, 16'd27487, 16'd49562, 16'd42548, 16'd14934, 16'd44087, 16'd64598, 16'd49741, 16'd29413, 16'd11347, 16'd29697, 16'd37588, 16'd29327, 16'd32450, 16'd48875, 16'd1841, 16'd2924, 16'd64627, 16'd24281, 16'd2227, 16'd45300, 16'd27313, 16'd38504, 16'd2351});
	test_expansion(128'h3b573aa812e4984363a2f1ac0a8b8f30, {16'd53741, 16'd50109, 16'd2809, 16'd47324, 16'd48758, 16'd55442, 16'd32104, 16'd44807, 16'd57943, 16'd46066, 16'd14361, 16'd48071, 16'd29211, 16'd16934, 16'd21241, 16'd59867, 16'd36612, 16'd21320, 16'd3139, 16'd18836, 16'd12451, 16'd6225, 16'd50229, 16'd21912, 16'd44809, 16'd64158});
	test_expansion(128'h94eb09c6cd53bb43dabd71fdc0aa5874, {16'd52494, 16'd42589, 16'd49534, 16'd21683, 16'd3963, 16'd16815, 16'd45815, 16'd49743, 16'd61434, 16'd64252, 16'd10575, 16'd35777, 16'd60146, 16'd21956, 16'd28630, 16'd41854, 16'd49369, 16'd9415, 16'd65254, 16'd22252, 16'd62667, 16'd40644, 16'd47399, 16'd14382, 16'd49766, 16'd18808});
	test_expansion(128'h5035ea932965ff9d65d81b3cc65a3778, {16'd25052, 16'd34424, 16'd59588, 16'd57888, 16'd28902, 16'd36174, 16'd60315, 16'd46866, 16'd361, 16'd35732, 16'd22951, 16'd32903, 16'd37371, 16'd63788, 16'd64261, 16'd9724, 16'd29047, 16'd7608, 16'd29464, 16'd51061, 16'd28365, 16'd30980, 16'd31178, 16'd18664, 16'd12877, 16'd25735});
	test_expansion(128'h26710a1eea60a6e7270de22f5d89c301, {16'd1451, 16'd9961, 16'd12739, 16'd52740, 16'd44940, 16'd54685, 16'd32369, 16'd1599, 16'd49509, 16'd14859, 16'd25438, 16'd18706, 16'd25885, 16'd56334, 16'd52443, 16'd10490, 16'd46068, 16'd54288, 16'd27980, 16'd9061, 16'd61897, 16'd18905, 16'd24184, 16'd40288, 16'd62721, 16'd38919});
	test_expansion(128'hf5f637b6aa73b1f4da82aada0402881a, {16'd43058, 16'd58582, 16'd57383, 16'd57910, 16'd3529, 16'd2114, 16'd44983, 16'd49026, 16'd24055, 16'd12504, 16'd60676, 16'd11971, 16'd14882, 16'd625, 16'd39907, 16'd38358, 16'd19933, 16'd25131, 16'd48443, 16'd36198, 16'd15105, 16'd12706, 16'd14242, 16'd42507, 16'd37920, 16'd19333});
	test_expansion(128'h9f1ef5b83af376904b295f3b536e3cd6, {16'd35824, 16'd45044, 16'd17589, 16'd6884, 16'd48173, 16'd27214, 16'd19641, 16'd64170, 16'd7600, 16'd40330, 16'd26438, 16'd46848, 16'd4509, 16'd60974, 16'd3099, 16'd2757, 16'd42439, 16'd2984, 16'd17776, 16'd11943, 16'd18604, 16'd27661, 16'd13159, 16'd65327, 16'd9741, 16'd39795});
	test_expansion(128'h6e9c03e49597b379ca17183d4bbfd37e, {16'd24946, 16'd47335, 16'd43343, 16'd8394, 16'd16333, 16'd17165, 16'd53800, 16'd43922, 16'd59313, 16'd59076, 16'd42949, 16'd61567, 16'd32963, 16'd35065, 16'd18712, 16'd25348, 16'd56165, 16'd13503, 16'd23001, 16'd8711, 16'd63982, 16'd9827, 16'd31395, 16'd53849, 16'd7167, 16'd30953});
	test_expansion(128'h72a54478d1e7c81f3830ac240069b7c7, {16'd41745, 16'd40027, 16'd16025, 16'd7997, 16'd18282, 16'd3050, 16'd20313, 16'd65524, 16'd55684, 16'd52176, 16'd19940, 16'd30622, 16'd59993, 16'd64874, 16'd58121, 16'd28715, 16'd24360, 16'd47774, 16'd16566, 16'd31002, 16'd48261, 16'd52578, 16'd45408, 16'd12995, 16'd11464, 16'd12882});
	test_expansion(128'h15d87a7492bdede2d65ba4f9dde192aa, {16'd41963, 16'd19569, 16'd8968, 16'd50564, 16'd37621, 16'd54347, 16'd44142, 16'd6721, 16'd477, 16'd55057, 16'd19745, 16'd50213, 16'd20245, 16'd39466, 16'd21045, 16'd45357, 16'd1528, 16'd58344, 16'd12769, 16'd14182, 16'd19805, 16'd50271, 16'd34427, 16'd51534, 16'd54754, 16'd39741});
	test_expansion(128'h3e88e9b447c145e60cdfb68a2810bcf5, {16'd59645, 16'd6584, 16'd32869, 16'd1567, 16'd51005, 16'd22681, 16'd23841, 16'd13524, 16'd45153, 16'd56016, 16'd1233, 16'd58888, 16'd63579, 16'd1090, 16'd2865, 16'd18659, 16'd12267, 16'd49074, 16'd31197, 16'd14125, 16'd20286, 16'd47663, 16'd60016, 16'd45366, 16'd51309, 16'd22372});
	test_expansion(128'h90edf137aa5974574ca3fda90e63ba61, {16'd59930, 16'd35148, 16'd53890, 16'd17253, 16'd6491, 16'd5541, 16'd17877, 16'd7092, 16'd7819, 16'd17994, 16'd35225, 16'd38785, 16'd54878, 16'd35584, 16'd52397, 16'd36343, 16'd10836, 16'd55273, 16'd18830, 16'd7656, 16'd51110, 16'd15789, 16'd1224, 16'd49792, 16'd23873, 16'd24948});
	test_expansion(128'hb4eb3ecab9066d2eb177e95e95ff397b, {16'd1559, 16'd21554, 16'd56179, 16'd11626, 16'd35926, 16'd11910, 16'd29127, 16'd52047, 16'd8190, 16'd2412, 16'd31515, 16'd48721, 16'd38765, 16'd56967, 16'd45973, 16'd62509, 16'd2396, 16'd12229, 16'd40605, 16'd55902, 16'd61461, 16'd12941, 16'd46919, 16'd18317, 16'd62824, 16'd4150});
	test_expansion(128'h4db6ade44540789bfcb906a211470cb9, {16'd29330, 16'd17813, 16'd45290, 16'd30782, 16'd52768, 16'd3467, 16'd46969, 16'd57477, 16'd60177, 16'd35923, 16'd20580, 16'd42692, 16'd55448, 16'd38223, 16'd15161, 16'd1452, 16'd42190, 16'd52235, 16'd24794, 16'd11564, 16'd13699, 16'd8556, 16'd44726, 16'd21798, 16'd60560, 16'd17568});
	test_expansion(128'h6cfadc04fe7b5db423f18768f9353957, {16'd58012, 16'd905, 16'd58297, 16'd36220, 16'd6158, 16'd47928, 16'd26459, 16'd41802, 16'd12834, 16'd18047, 16'd49688, 16'd736, 16'd22678, 16'd12243, 16'd24911, 16'd27225, 16'd8837, 16'd39877, 16'd59332, 16'd44593, 16'd64356, 16'd44481, 16'd16694, 16'd64374, 16'd2848, 16'd57519});
	test_expansion(128'haf65a30cf9961d3247d0da742587c47f, {16'd57165, 16'd57964, 16'd49347, 16'd40284, 16'd48014, 16'd12065, 16'd30727, 16'd43159, 16'd63003, 16'd13769, 16'd8571, 16'd33051, 16'd52414, 16'd36048, 16'd34679, 16'd33896, 16'd53268, 16'd48061, 16'd36016, 16'd5871, 16'd20248, 16'd29823, 16'd27969, 16'd53592, 16'd3649, 16'd53901});
	test_expansion(128'hcb7d38b808336bf4555542bf7fae28d1, {16'd50163, 16'd20494, 16'd14076, 16'd42294, 16'd60437, 16'd56419, 16'd65304, 16'd32473, 16'd26331, 16'd18455, 16'd37720, 16'd8836, 16'd6342, 16'd33406, 16'd46848, 16'd48724, 16'd2340, 16'd34283, 16'd35258, 16'd21278, 16'd3622, 16'd22592, 16'd32991, 16'd31987, 16'd42560, 16'd20783});
	test_expansion(128'h939f71508eeb81c206ca00fe5c8df7ad, {16'd55721, 16'd41135, 16'd11355, 16'd11301, 16'd5973, 16'd3956, 16'd51717, 16'd46431, 16'd53857, 16'd35193, 16'd48790, 16'd54405, 16'd35905, 16'd58903, 16'd61236, 16'd51020, 16'd57800, 16'd63496, 16'd34357, 16'd28232, 16'd16963, 16'd7460, 16'd50142, 16'd37453, 16'd37594, 16'd25092});
	test_expansion(128'h7062edcb2334f592be394208e2de7610, {16'd60922, 16'd53589, 16'd36090, 16'd44975, 16'd53861, 16'd15286, 16'd32882, 16'd38224, 16'd53731, 16'd12635, 16'd35890, 16'd28258, 16'd32418, 16'd63443, 16'd31472, 16'd47599, 16'd5798, 16'd39709, 16'd41819, 16'd16030, 16'd56256, 16'd21544, 16'd33911, 16'd27442, 16'd14451, 16'd63847});
	test_expansion(128'h94b3a88ada5930caf97355901cfa595a, {16'd26081, 16'd8968, 16'd16577, 16'd13985, 16'd37707, 16'd35669, 16'd7093, 16'd25471, 16'd25792, 16'd30467, 16'd57727, 16'd38203, 16'd9456, 16'd23951, 16'd54232, 16'd35850, 16'd10759, 16'd50787, 16'd1454, 16'd18738, 16'd37666, 16'd17492, 16'd64059, 16'd33592, 16'd22611, 16'd51070});
	test_expansion(128'h0cec38f337bee7296efb2b178316bdfd, {16'd1905, 16'd2320, 16'd28227, 16'd26134, 16'd14127, 16'd59476, 16'd943, 16'd53962, 16'd56892, 16'd33884, 16'd16255, 16'd42301, 16'd40927, 16'd23234, 16'd12470, 16'd21271, 16'd22484, 16'd13495, 16'd8038, 16'd48092, 16'd4065, 16'd14852, 16'd29303, 16'd36566, 16'd57424, 16'd38682});
	test_expansion(128'hb63fc26b45aa4b2ef233415837dc0925, {16'd61807, 16'd3134, 16'd11869, 16'd60741, 16'd11275, 16'd19680, 16'd16309, 16'd41447, 16'd65151, 16'd20082, 16'd16347, 16'd49766, 16'd46326, 16'd25806, 16'd52936, 16'd50992, 16'd863, 16'd46343, 16'd33384, 16'd61325, 16'd39710, 16'd13513, 16'd40854, 16'd25731, 16'd62019, 16'd43878});
	test_expansion(128'h50357e07b7f49fff6689d8a57fe2828f, {16'd37593, 16'd63838, 16'd26354, 16'd29494, 16'd33928, 16'd39121, 16'd13685, 16'd12460, 16'd8032, 16'd11886, 16'd58161, 16'd58738, 16'd34749, 16'd36190, 16'd34587, 16'd10773, 16'd64295, 16'd19605, 16'd14772, 16'd40726, 16'd65328, 16'd25567, 16'd64812, 16'd52404, 16'd33304, 16'd27038});
	test_expansion(128'hfb314f8b268c574de64e2732e72a89ee, {16'd43073, 16'd28722, 16'd21906, 16'd61891, 16'd934, 16'd14866, 16'd4372, 16'd36388, 16'd47067, 16'd10665, 16'd56764, 16'd38550, 16'd3782, 16'd27881, 16'd43240, 16'd14628, 16'd39925, 16'd47986, 16'd37537, 16'd9177, 16'd25286, 16'd46074, 16'd31090, 16'd35028, 16'd16676, 16'd6978});
	test_expansion(128'h74776f7e6a32dfa76115d76df1448617, {16'd64504, 16'd65500, 16'd28266, 16'd38135, 16'd47534, 16'd33888, 16'd3742, 16'd37408, 16'd9083, 16'd55316, 16'd36601, 16'd37297, 16'd16234, 16'd49925, 16'd2897, 16'd11779, 16'd58831, 16'd62133, 16'd39595, 16'd16407, 16'd15958, 16'd8444, 16'd9057, 16'd36001, 16'd46508, 16'd35909});
	test_expansion(128'hb300c029ab4ae3cf65be75cc11456656, {16'd46423, 16'd43105, 16'd35756, 16'd61170, 16'd15916, 16'd37845, 16'd16889, 16'd42508, 16'd20589, 16'd5638, 16'd57643, 16'd6934, 16'd53721, 16'd53279, 16'd10103, 16'd2795, 16'd59572, 16'd65460, 16'd49904, 16'd14437, 16'd279, 16'd9567, 16'd58108, 16'd39748, 16'd33619, 16'd14377});
	test_expansion(128'h1c0281f4b78bb3c87b0293192e8dc807, {16'd1711, 16'd5973, 16'd5938, 16'd32891, 16'd55350, 16'd26382, 16'd38461, 16'd54301, 16'd62952, 16'd18304, 16'd52998, 16'd10191, 16'd19044, 16'd15861, 16'd10034, 16'd61487, 16'd54274, 16'd11191, 16'd35763, 16'd38981, 16'd1155, 16'd41369, 16'd10055, 16'd28430, 16'd46200, 16'd31627});
	test_expansion(128'h144965434f4f4b90e5b00a483b1ad616, {16'd9154, 16'd20288, 16'd34595, 16'd61, 16'd43103, 16'd58263, 16'd50473, 16'd42614, 16'd5065, 16'd25684, 16'd20674, 16'd22545, 16'd46885, 16'd12563, 16'd32197, 16'd19378, 16'd47517, 16'd10605, 16'd21588, 16'd65447, 16'd13752, 16'd13024, 16'd8818, 16'd33609, 16'd16993, 16'd33413});
	test_expansion(128'hb9a8b501457e3e0ab4c7526aa6778c17, {16'd10562, 16'd20322, 16'd18767, 16'd31237, 16'd45570, 16'd63763, 16'd47561, 16'd32348, 16'd41841, 16'd3219, 16'd13886, 16'd52026, 16'd22833, 16'd65057, 16'd33182, 16'd33085, 16'd49347, 16'd18747, 16'd32891, 16'd33408, 16'd47397, 16'd40734, 16'd28054, 16'd54341, 16'd26462, 16'd20103});
	test_expansion(128'h2f499963e9e60872165a19782225d553, {16'd27239, 16'd47220, 16'd58801, 16'd754, 16'd39665, 16'd13334, 16'd26682, 16'd19975, 16'd55828, 16'd52528, 16'd29014, 16'd11432, 16'd5929, 16'd7350, 16'd27291, 16'd5838, 16'd10006, 16'd60536, 16'd34030, 16'd8561, 16'd40825, 16'd6277, 16'd36551, 16'd58957, 16'd46695, 16'd14428});
	test_expansion(128'hd9c888eed6bb6c00095dcf0539541c94, {16'd25028, 16'd18351, 16'd53326, 16'd4352, 16'd23651, 16'd61769, 16'd27488, 16'd33676, 16'd52686, 16'd7206, 16'd63143, 16'd21140, 16'd40188, 16'd42282, 16'd46691, 16'd21452, 16'd28270, 16'd17426, 16'd23790, 16'd40422, 16'd29568, 16'd22389, 16'd13740, 16'd37921, 16'd719, 16'd8839});
	test_expansion(128'ha9786df3585b012a027e0b281eedf495, {16'd60368, 16'd798, 16'd44233, 16'd7225, 16'd46143, 16'd12473, 16'd44410, 16'd51403, 16'd39973, 16'd19134, 16'd5303, 16'd51442, 16'd57884, 16'd65386, 16'd26326, 16'd39022, 16'd8033, 16'd14569, 16'd10407, 16'd48774, 16'd3003, 16'd32361, 16'd20605, 16'd621, 16'd34235, 16'd15070});
	test_expansion(128'h14acceef48e2c1d52aba3fb053d6aa7a, {16'd18386, 16'd52423, 16'd42938, 16'd58631, 16'd39149, 16'd15349, 16'd32592, 16'd47603, 16'd8906, 16'd44462, 16'd44123, 16'd16098, 16'd14088, 16'd19719, 16'd24729, 16'd14236, 16'd2640, 16'd40595, 16'd17303, 16'd48582, 16'd7150, 16'd43960, 16'd60033, 16'd1771, 16'd44120, 16'd25299});
	test_expansion(128'h76896b59e0f2327264ed11ec587fb240, {16'd48924, 16'd45958, 16'd58174, 16'd25423, 16'd1606, 16'd50179, 16'd6675, 16'd19669, 16'd35461, 16'd6453, 16'd36176, 16'd51875, 16'd53215, 16'd33617, 16'd15484, 16'd44156, 16'd28492, 16'd34937, 16'd10330, 16'd12076, 16'd39327, 16'd3224, 16'd62116, 16'd65281, 16'd25107, 16'd48033});
	test_expansion(128'hd1ef484a1683cfbaf4d1f4b5b179ed6c, {16'd11877, 16'd29281, 16'd29943, 16'd44853, 16'd44965, 16'd28407, 16'd16955, 16'd27669, 16'd58620, 16'd52287, 16'd36460, 16'd15074, 16'd26768, 16'd23513, 16'd7128, 16'd36243, 16'd15040, 16'd24824, 16'd60673, 16'd27719, 16'd18547, 16'd8981, 16'd42905, 16'd50536, 16'd55827, 16'd5083});
	test_expansion(128'h4e2d6b59a26be9440b1d5a26cc8fb922, {16'd9100, 16'd7008, 16'd15876, 16'd29595, 16'd60633, 16'd22701, 16'd21830, 16'd44438, 16'd56916, 16'd24759, 16'd12064, 16'd49009, 16'd1978, 16'd11123, 16'd20321, 16'd27754, 16'd10305, 16'd1308, 16'd2717, 16'd23592, 16'd46775, 16'd47283, 16'd20235, 16'd4639, 16'd39299, 16'd65115});
	test_expansion(128'heae501855d41e8b1baef0b52fe8f6862, {16'd8807, 16'd41844, 16'd35411, 16'd57165, 16'd60287, 16'd1124, 16'd19541, 16'd26117, 16'd44515, 16'd35945, 16'd37372, 16'd43816, 16'd13292, 16'd42331, 16'd6747, 16'd40617, 16'd58949, 16'd12195, 16'd45081, 16'd8464, 16'd58374, 16'd51790, 16'd36191, 16'd9752, 16'd12887, 16'd1904});
	test_expansion(128'ha05fae822b57f2106e8ca1fa64f1a41c, {16'd51157, 16'd44409, 16'd60897, 16'd25552, 16'd44515, 16'd21613, 16'd44880, 16'd54478, 16'd57073, 16'd31158, 16'd9520, 16'd65509, 16'd46387, 16'd54332, 16'd20215, 16'd56118, 16'd13591, 16'd7584, 16'd55975, 16'd17194, 16'd12048, 16'd31743, 16'd46752, 16'd33022, 16'd60286, 16'd1577});
	test_expansion(128'hd2c19507a41185257022177c665ac1a5, {16'd64708, 16'd44108, 16'd7337, 16'd28225, 16'd27853, 16'd63803, 16'd42940, 16'd11143, 16'd23813, 16'd39529, 16'd60620, 16'd51777, 16'd16486, 16'd1705, 16'd40614, 16'd5047, 16'd54044, 16'd46608, 16'd12471, 16'd57770, 16'd33176, 16'd1729, 16'd61438, 16'd26793, 16'd64860, 16'd38498});
	test_expansion(128'ha2a9e27da6d636a8a12b19bec42b70c6, {16'd60981, 16'd25631, 16'd54372, 16'd16973, 16'd2897, 16'd865, 16'd48040, 16'd5605, 16'd11856, 16'd19807, 16'd9881, 16'd18518, 16'd61061, 16'd48605, 16'd25585, 16'd51720, 16'd65002, 16'd19160, 16'd30705, 16'd31393, 16'd24132, 16'd8839, 16'd3338, 16'd64882, 16'd56570, 16'd55273});
	test_expansion(128'h520d601b7f82f8e2478470a408cee019, {16'd37966, 16'd48527, 16'd4737, 16'd8474, 16'd27622, 16'd13046, 16'd7969, 16'd64079, 16'd23386, 16'd56161, 16'd41123, 16'd9233, 16'd38579, 16'd9300, 16'd44619, 16'd34517, 16'd52969, 16'd44488, 16'd16044, 16'd8157, 16'd4133, 16'd2430, 16'd61750, 16'd2463, 16'd34218, 16'd715});
	test_expansion(128'he1315de4ba7ebafdf8a7388de746d0e6, {16'd56404, 16'd28831, 16'd10089, 16'd32628, 16'd41642, 16'd30970, 16'd36096, 16'd1710, 16'd6204, 16'd32327, 16'd3399, 16'd3564, 16'd20843, 16'd41137, 16'd56094, 16'd53123, 16'd33681, 16'd59043, 16'd54465, 16'd44725, 16'd56662, 16'd28047, 16'd62025, 16'd43402, 16'd43843, 16'd27599});
	test_expansion(128'h1379262b29be0821ea08b2352bc63ff3, {16'd2677, 16'd12455, 16'd34427, 16'd43017, 16'd50906, 16'd30271, 16'd65120, 16'd29808, 16'd2001, 16'd32386, 16'd49881, 16'd360, 16'd26627, 16'd44417, 16'd32479, 16'd37506, 16'd56112, 16'd53338, 16'd59654, 16'd61095, 16'd64521, 16'd9474, 16'd33329, 16'd25214, 16'd41112, 16'd19065});
	test_expansion(128'hb7b186c0e43a91ffa672d8b42978aff9, {16'd60799, 16'd18006, 16'd63187, 16'd50932, 16'd2399, 16'd25717, 16'd65282, 16'd49314, 16'd61567, 16'd13148, 16'd660, 16'd47906, 16'd14215, 16'd21109, 16'd65436, 16'd23902, 16'd3101, 16'd5333, 16'd42589, 16'd7035, 16'd53341, 16'd3001, 16'd30804, 16'd17968, 16'd32468, 16'd61997});
	test_expansion(128'h70070080f6512f0f867e216194116d22, {16'd38109, 16'd33928, 16'd17121, 16'd59096, 16'd47179, 16'd38228, 16'd8628, 16'd54018, 16'd54359, 16'd41799, 16'd44912, 16'd64847, 16'd12205, 16'd29629, 16'd13787, 16'd13894, 16'd62612, 16'd54865, 16'd62521, 16'd1144, 16'd7828, 16'd21661, 16'd52198, 16'd35425, 16'd31570, 16'd58701});
	test_expansion(128'hd8e773339ef8110d435226f80a48e4f9, {16'd25879, 16'd12115, 16'd51093, 16'd46690, 16'd22594, 16'd48437, 16'd1646, 16'd57773, 16'd57747, 16'd1195, 16'd21548, 16'd31511, 16'd17294, 16'd4836, 16'd51673, 16'd26074, 16'd14349, 16'd23274, 16'd4646, 16'd36276, 16'd33168, 16'd10527, 16'd57940, 16'd23092, 16'd17961, 16'd18134});
	test_expansion(128'h5a175c751672bab2612429168a79ef34, {16'd8834, 16'd9886, 16'd19700, 16'd43044, 16'd47801, 16'd57821, 16'd29513, 16'd30408, 16'd44678, 16'd47118, 16'd21577, 16'd16594, 16'd51991, 16'd64407, 16'd56483, 16'd39156, 16'd33551, 16'd8729, 16'd27472, 16'd56879, 16'd29179, 16'd42236, 16'd2974, 16'd53183, 16'd14050, 16'd48011});
	test_expansion(128'hdde79a3e533d93e23ea4cb302507ee64, {16'd32490, 16'd28785, 16'd59578, 16'd19662, 16'd8612, 16'd28987, 16'd2766, 16'd57193, 16'd29630, 16'd7082, 16'd21881, 16'd11813, 16'd43727, 16'd8929, 16'd6038, 16'd25386, 16'd42408, 16'd63928, 16'd16785, 16'd36599, 16'd38563, 16'd40911, 16'd16229, 16'd50051, 16'd6367, 16'd54605});
	test_expansion(128'h22be8df76db12fae2dce4f31aced6264, {16'd10881, 16'd34460, 16'd45126, 16'd5646, 16'd57612, 16'd37019, 16'd17535, 16'd19194, 16'd43999, 16'd23069, 16'd5791, 16'd51645, 16'd15604, 16'd52005, 16'd51591, 16'd63271, 16'd44269, 16'd18277, 16'd53055, 16'd31633, 16'd56846, 16'd56690, 16'd37529, 16'd62044, 16'd26955, 16'd1536});
	test_expansion(128'he1452991816a685912f59fce3a57528f, {16'd29302, 16'd13707, 16'd56303, 16'd13098, 16'd61351, 16'd58309, 16'd58703, 16'd16568, 16'd45264, 16'd51553, 16'd24107, 16'd35812, 16'd62159, 16'd32739, 16'd65443, 16'd37300, 16'd5535, 16'd1068, 16'd21157, 16'd14687, 16'd51513, 16'd9621, 16'd20273, 16'd50962, 16'd60943, 16'd15907});
	test_expansion(128'hcae9324ac7f271eb828bf3442419c1a4, {16'd14791, 16'd25738, 16'd40687, 16'd11626, 16'd8317, 16'd44495, 16'd15655, 16'd23500, 16'd56803, 16'd16140, 16'd58671, 16'd20834, 16'd6218, 16'd63001, 16'd25814, 16'd51829, 16'd49252, 16'd3262, 16'd52460, 16'd50597, 16'd64515, 16'd9163, 16'd51702, 16'd7011, 16'd17200, 16'd23193});
	test_expansion(128'h0eda9e710780b835e8a3b46a75042a0b, {16'd34356, 16'd15, 16'd610, 16'd49678, 16'd18597, 16'd21428, 16'd54934, 16'd59576, 16'd36983, 16'd14988, 16'd49841, 16'd48852, 16'd370, 16'd45919, 16'd61754, 16'd54980, 16'd12077, 16'd49192, 16'd42626, 16'd64156, 16'd18570, 16'd7123, 16'd55501, 16'd46992, 16'd19926, 16'd54132});
	test_expansion(128'hdc53937c1f2258a17b64f39b569ad609, {16'd48563, 16'd7424, 16'd60483, 16'd64778, 16'd46844, 16'd34344, 16'd17239, 16'd34401, 16'd7350, 16'd6848, 16'd31820, 16'd40270, 16'd57456, 16'd50287, 16'd40897, 16'd49223, 16'd31354, 16'd41980, 16'd17596, 16'd59542, 16'd39334, 16'd53401, 16'd40197, 16'd507, 16'd37431, 16'd29371});
	test_expansion(128'hde82c3e62500fdeee4fdee3eb89c30d2, {16'd33845, 16'd35651, 16'd41574, 16'd202, 16'd55623, 16'd60723, 16'd45520, 16'd53477, 16'd25376, 16'd4541, 16'd44894, 16'd49835, 16'd9190, 16'd20158, 16'd24805, 16'd3422, 16'd34101, 16'd10732, 16'd28584, 16'd46260, 16'd4296, 16'd3271, 16'd32878, 16'd8861, 16'd2062, 16'd14175});
	test_expansion(128'hbb4b37a445a0afcce876c48da85977d3, {16'd63317, 16'd41063, 16'd14124, 16'd15960, 16'd18762, 16'd1271, 16'd7769, 16'd20018, 16'd8163, 16'd30926, 16'd45698, 16'd42639, 16'd26597, 16'd16747, 16'd32205, 16'd40515, 16'd17423, 16'd28432, 16'd39911, 16'd40511, 16'd41577, 16'd30451, 16'd24303, 16'd8200, 16'd48754, 16'd33091});
	test_expansion(128'h3a9a3d9aad4ed9d6c31f50b85b969317, {16'd12208, 16'd28743, 16'd44949, 16'd55222, 16'd15355, 16'd19382, 16'd34582, 16'd25031, 16'd57868, 16'd50000, 16'd27422, 16'd16334, 16'd52230, 16'd28548, 16'd38582, 16'd9535, 16'd50785, 16'd49603, 16'd5258, 16'd64570, 16'd51109, 16'd65393, 16'd64610, 16'd28429, 16'd33721, 16'd49999});
	test_expansion(128'hc49f47462501e229d9b154183e42d8e9, {16'd24999, 16'd19476, 16'd11850, 16'd11546, 16'd31377, 16'd14912, 16'd17925, 16'd6130, 16'd53937, 16'd26220, 16'd38573, 16'd49015, 16'd25168, 16'd56791, 16'd26267, 16'd31696, 16'd28451, 16'd11250, 16'd31103, 16'd39996, 16'd22687, 16'd56650, 16'd40098, 16'd6007, 16'd6275, 16'd20144});
	test_expansion(128'h5c623662cfc5ff82997c954a79fc99ac, {16'd39681, 16'd50289, 16'd61946, 16'd49498, 16'd58887, 16'd63661, 16'd34523, 16'd64205, 16'd36871, 16'd54803, 16'd62430, 16'd4398, 16'd19922, 16'd4254, 16'd19733, 16'd1035, 16'd1526, 16'd44451, 16'd42504, 16'd48966, 16'd18827, 16'd49997, 16'd30759, 16'd30479, 16'd19520, 16'd62143});
	test_expansion(128'h602f3e0cc137453654028d570fefc4bc, {16'd28974, 16'd10524, 16'd36220, 16'd6656, 16'd59826, 16'd34346, 16'd50970, 16'd17986, 16'd3483, 16'd17211, 16'd62804, 16'd57293, 16'd15608, 16'd54323, 16'd57961, 16'd3162, 16'd4805, 16'd16943, 16'd12817, 16'd44389, 16'd55884, 16'd2456, 16'd23401, 16'd40316, 16'd42908, 16'd33730});
	test_expansion(128'hde22f7aa82b328844d3ee09852d11667, {16'd3751, 16'd9887, 16'd14950, 16'd22017, 16'd2000, 16'd25948, 16'd7548, 16'd6442, 16'd21892, 16'd35535, 16'd53899, 16'd20365, 16'd10101, 16'd58379, 16'd13433, 16'd13752, 16'd691, 16'd17690, 16'd12740, 16'd56344, 16'd3329, 16'd9219, 16'd12061, 16'd43939, 16'd46690, 16'd41961});
	test_expansion(128'hb023bc9afd5f6c80fd26386ad951603e, {16'd11792, 16'd29159, 16'd60121, 16'd29371, 16'd35725, 16'd12345, 16'd54978, 16'd61418, 16'd42051, 16'd44788, 16'd56876, 16'd50521, 16'd19275, 16'd36572, 16'd31319, 16'd63114, 16'd19807, 16'd23205, 16'd57042, 16'd10442, 16'd4430, 16'd45700, 16'd35711, 16'd47192, 16'd8410, 16'd23868});
	test_expansion(128'h6ef908ec298a18d2e17fb3cf9049fc60, {16'd48113, 16'd27752, 16'd26968, 16'd41047, 16'd24725, 16'd64710, 16'd48408, 16'd42332, 16'd63094, 16'd10283, 16'd56447, 16'd46474, 16'd52781, 16'd11117, 16'd4648, 16'd23045, 16'd22272, 16'd56464, 16'd22019, 16'd53386, 16'd64782, 16'd55364, 16'd10303, 16'd61700, 16'd24530, 16'd25699});
	test_expansion(128'h4e7ec799e98645bdcbe12515e58b2498, {16'd60258, 16'd9696, 16'd63229, 16'd14645, 16'd52804, 16'd6196, 16'd735, 16'd63345, 16'd13348, 16'd52876, 16'd51370, 16'd24799, 16'd61065, 16'd16091, 16'd51411, 16'd13715, 16'd3125, 16'd12506, 16'd59700, 16'd45021, 16'd9739, 16'd28967, 16'd29296, 16'd54116, 16'd4498, 16'd42592});
	test_expansion(128'h776d00cbcd9835720806b67dd0d5590f, {16'd33925, 16'd55219, 16'd38549, 16'd50238, 16'd38538, 16'd28865, 16'd28358, 16'd49831, 16'd64083, 16'd20170, 16'd44477, 16'd47141, 16'd40764, 16'd31869, 16'd27958, 16'd7559, 16'd51182, 16'd55223, 16'd17209, 16'd41107, 16'd21569, 16'd58491, 16'd35659, 16'd8439, 16'd9477, 16'd34902});
	test_expansion(128'h38784ff4675a2cf13255120cdec61c63, {16'd46740, 16'd12058, 16'd28047, 16'd12186, 16'd15189, 16'd26633, 16'd59502, 16'd50962, 16'd28154, 16'd37775, 16'd62529, 16'd55918, 16'd7576, 16'd24835, 16'd41115, 16'd41823, 16'd24877, 16'd50520, 16'd59299, 16'd62821, 16'd9787, 16'd49744, 16'd19733, 16'd29617, 16'd5635, 16'd2146});
	test_expansion(128'hb93c3b8d502e8e2b9bae5db0bf013795, {16'd25956, 16'd56932, 16'd55878, 16'd62956, 16'd56876, 16'd35734, 16'd26436, 16'd11536, 16'd22400, 16'd26141, 16'd54372, 16'd60597, 16'd531, 16'd30855, 16'd60264, 16'd37515, 16'd26685, 16'd40000, 16'd18616, 16'd1263, 16'd55869, 16'd51860, 16'd4632, 16'd8835, 16'd11447, 16'd56379});
	test_expansion(128'h77bad688f227e287d55566cbe138c2c0, {16'd25557, 16'd12585, 16'd31422, 16'd1320, 16'd32525, 16'd140, 16'd61786, 16'd48076, 16'd47528, 16'd21070, 16'd2274, 16'd35794, 16'd34569, 16'd20407, 16'd15042, 16'd23221, 16'd49385, 16'd5278, 16'd37778, 16'd18234, 16'd61145, 16'd59635, 16'd47393, 16'd30468, 16'd45217, 16'd48329});
	test_expansion(128'h335344ca708b06a8349db2c932794909, {16'd19887, 16'd58218, 16'd24923, 16'd41355, 16'd4573, 16'd28950, 16'd56407, 16'd30007, 16'd14167, 16'd51831, 16'd57122, 16'd4128, 16'd41363, 16'd30472, 16'd60248, 16'd54047, 16'd51085, 16'd2467, 16'd44500, 16'd64453, 16'd60545, 16'd42277, 16'd5974, 16'd30421, 16'd12047, 16'd14490});
	test_expansion(128'hbbf36142e67e6e06cc8e4307e2b23ad5, {16'd59505, 16'd33270, 16'd9388, 16'd16659, 16'd2732, 16'd19897, 16'd2533, 16'd49136, 16'd4445, 16'd20758, 16'd12242, 16'd24782, 16'd32411, 16'd49846, 16'd52202, 16'd40682, 16'd57031, 16'd30725, 16'd25794, 16'd11027, 16'd23354, 16'd28952, 16'd17278, 16'd8674, 16'd57362, 16'd23374});
	test_expansion(128'he61e68e72c348dd34393871f9eb47f28, {16'd19610, 16'd64166, 16'd50037, 16'd10392, 16'd26294, 16'd53956, 16'd8744, 16'd38477, 16'd40913, 16'd16728, 16'd11958, 16'd58384, 16'd54811, 16'd25534, 16'd1442, 16'd49473, 16'd41121, 16'd59840, 16'd34133, 16'd24516, 16'd8367, 16'd18884, 16'd42420, 16'd3302, 16'd28723, 16'd32433});
	test_expansion(128'h9f5123b18b9d444b654fab9fa91bf2ea, {16'd22483, 16'd37138, 16'd22077, 16'd58007, 16'd32858, 16'd17712, 16'd41744, 16'd60048, 16'd50334, 16'd27360, 16'd7768, 16'd46322, 16'd19133, 16'd17372, 16'd54284, 16'd2206, 16'd10538, 16'd51652, 16'd33652, 16'd18359, 16'd50447, 16'd17615, 16'd23539, 16'd65133, 16'd53551, 16'd55822});
	test_expansion(128'h5bb80663bc8cdc009981f9ab68b87177, {16'd5180, 16'd55681, 16'd20892, 16'd45323, 16'd23848, 16'd41974, 16'd21129, 16'd42038, 16'd26549, 16'd41108, 16'd50058, 16'd28008, 16'd6625, 16'd42002, 16'd33770, 16'd48247, 16'd13163, 16'd25461, 16'd26340, 16'd11509, 16'd59640, 16'd46134, 16'd27449, 16'd64422, 16'd14875, 16'd13363});
	test_expansion(128'h551e750bbab020653f2d9c9d86ade576, {16'd44456, 16'd33917, 16'd38555, 16'd7178, 16'd49834, 16'd20549, 16'd63043, 16'd19055, 16'd60511, 16'd2866, 16'd37082, 16'd38096, 16'd36303, 16'd16502, 16'd54567, 16'd27277, 16'd55049, 16'd64561, 16'd12633, 16'd45073, 16'd49758, 16'd48513, 16'd46736, 16'd45547, 16'd23157, 16'd54684});
	test_expansion(128'h92c1a44220037fd341b5573ae7029375, {16'd33802, 16'd40325, 16'd26156, 16'd40559, 16'd4805, 16'd9864, 16'd55131, 16'd1363, 16'd3287, 16'd31124, 16'd62455, 16'd60306, 16'd19178, 16'd13491, 16'd23459, 16'd42393, 16'd46225, 16'd27187, 16'd21327, 16'd52670, 16'd27060, 16'd16282, 16'd64170, 16'd15258, 16'd57395, 16'd4863});
	test_expansion(128'h7addd3dd66fe23f45dafe0779512e252, {16'd31774, 16'd21144, 16'd14393, 16'd18941, 16'd59027, 16'd21763, 16'd6079, 16'd14608, 16'd53527, 16'd12547, 16'd61585, 16'd9125, 16'd42552, 16'd10251, 16'd38262, 16'd41860, 16'd9266, 16'd56804, 16'd6958, 16'd12574, 16'd827, 16'd58908, 16'd20937, 16'd35516, 16'd14509, 16'd16547});
	test_expansion(128'h632ec6230aebc51bf6dd22cbd0d15719, {16'd18175, 16'd22984, 16'd36284, 16'd8134, 16'd44849, 16'd53265, 16'd64265, 16'd34993, 16'd63137, 16'd42005, 16'd19788, 16'd24414, 16'd1932, 16'd34004, 16'd42539, 16'd6614, 16'd39394, 16'd9570, 16'd62879, 16'd12241, 16'd10839, 16'd19010, 16'd57785, 16'd1145, 16'd20151, 16'd3841});
	test_expansion(128'hcbaf3ec7b02e7a67c45a631b1c7eb4c6, {16'd27731, 16'd34303, 16'd41328, 16'd51723, 16'd16443, 16'd7264, 16'd107, 16'd10459, 16'd14869, 16'd36250, 16'd58999, 16'd50722, 16'd53948, 16'd6185, 16'd18194, 16'd12179, 16'd20325, 16'd23272, 16'd50157, 16'd32161, 16'd61616, 16'd33994, 16'd28260, 16'd16140, 16'd51687, 16'd25745});
	test_expansion(128'h1a23d35843ea0cbb5eea1818dc50c8b4, {16'd17048, 16'd1830, 16'd20611, 16'd63623, 16'd7029, 16'd12702, 16'd24634, 16'd23084, 16'd14658, 16'd22846, 16'd1738, 16'd22632, 16'd47987, 16'd7382, 16'd6147, 16'd60594, 16'd57347, 16'd48249, 16'd10087, 16'd17088, 16'd37459, 16'd44114, 16'd23408, 16'd8735, 16'd27886, 16'd9650});
	test_expansion(128'hadcc7fbe5bba0f8c088b9cb6ee46e146, {16'd7745, 16'd968, 16'd52272, 16'd24574, 16'd29360, 16'd17068, 16'd46614, 16'd3459, 16'd30428, 16'd36294, 16'd63257, 16'd31889, 16'd39820, 16'd20934, 16'd11725, 16'd48622, 16'd12756, 16'd64814, 16'd55778, 16'd34450, 16'd39434, 16'd37524, 16'd26955, 16'd45410, 16'd47110, 16'd24717});
	test_expansion(128'h688539c5d931e8f73ea7f326c7e5d919, {16'd11292, 16'd40194, 16'd20226, 16'd38635, 16'd22196, 16'd30237, 16'd37316, 16'd11284, 16'd48404, 16'd2692, 16'd35764, 16'd30731, 16'd41964, 16'd11792, 16'd65167, 16'd50554, 16'd51952, 16'd44024, 16'd41019, 16'd4196, 16'd13647, 16'd61779, 16'd8999, 16'd62575, 16'd29762, 16'd11467});
	test_expansion(128'hf883216bf546e45560363d940fdcd292, {16'd25307, 16'd22214, 16'd38109, 16'd875, 16'd60725, 16'd14071, 16'd17812, 16'd17716, 16'd59879, 16'd16021, 16'd14173, 16'd18355, 16'd5569, 16'd48672, 16'd10109, 16'd1798, 16'd52707, 16'd7986, 16'd43610, 16'd13407, 16'd34150, 16'd20981, 16'd50041, 16'd64343, 16'd13514, 16'd42244});
	test_expansion(128'h61d6ef11c9b5e7335882e1e8f1ef2d04, {16'd60408, 16'd28271, 16'd6913, 16'd23137, 16'd34986, 16'd34012, 16'd3614, 16'd45468, 16'd11364, 16'd10396, 16'd46148, 16'd60986, 16'd50176, 16'd18355, 16'd45468, 16'd36038, 16'd19903, 16'd54065, 16'd44192, 16'd32842, 16'd30593, 16'd21516, 16'd60428, 16'd63113, 16'd30522, 16'd23198});
	test_expansion(128'h3938fe2287073348f6ed0e66f591a517, {16'd9258, 16'd56243, 16'd54535, 16'd3925, 16'd62136, 16'd63075, 16'd33877, 16'd11990, 16'd59403, 16'd27644, 16'd12161, 16'd19890, 16'd51591, 16'd12426, 16'd45765, 16'd22627, 16'd39836, 16'd23286, 16'd12471, 16'd9365, 16'd12299, 16'd38831, 16'd37997, 16'd28946, 16'd41038, 16'd47718});
	test_expansion(128'h1f1fac91c1dbf50add505a1ac508bcb5, {16'd8479, 16'd57268, 16'd46772, 16'd31747, 16'd44488, 16'd62624, 16'd60664, 16'd58351, 16'd12888, 16'd48193, 16'd13204, 16'd1137, 16'd57181, 16'd45558, 16'd4995, 16'd52059, 16'd8907, 16'd30224, 16'd29866, 16'd16715, 16'd54150, 16'd6066, 16'd14096, 16'd59423, 16'd62032, 16'd47088});
	test_expansion(128'hc19ac6b1282ec6c6e5e82cfa85af7ce8, {16'd24406, 16'd243, 16'd13531, 16'd19185, 16'd49731, 16'd9618, 16'd56933, 16'd51702, 16'd64624, 16'd35269, 16'd12747, 16'd39241, 16'd31400, 16'd24339, 16'd250, 16'd53052, 16'd58047, 16'd27146, 16'd2303, 16'd49508, 16'd49393, 16'd49154, 16'd45159, 16'd36452, 16'd40282, 16'd10776});
	test_expansion(128'h2079953b6fe97acbae462bf364da0f05, {16'd22506, 16'd53253, 16'd13043, 16'd587, 16'd6100, 16'd13134, 16'd6726, 16'd38289, 16'd19558, 16'd58193, 16'd58993, 16'd38335, 16'd41362, 16'd59197, 16'd51224, 16'd6860, 16'd210, 16'd42500, 16'd35881, 16'd55698, 16'd8081, 16'd50768, 16'd51366, 16'd65383, 16'd13441, 16'd6521});
	test_expansion(128'h4fdd9c13d5b2ba18d9d1a5bae34e6626, {16'd34015, 16'd45006, 16'd18849, 16'd3585, 16'd60656, 16'd14768, 16'd6947, 16'd59891, 16'd20423, 16'd45668, 16'd15824, 16'd21494, 16'd22322, 16'd4385, 16'd21092, 16'd18741, 16'd54066, 16'd10875, 16'd18143, 16'd61439, 16'd5646, 16'd44426, 16'd14371, 16'd10606, 16'd63360, 16'd52654});
	test_expansion(128'hbf941ed5fc5ea6d4f63339f109c50fcd, {16'd62748, 16'd32898, 16'd24451, 16'd39499, 16'd59284, 16'd53863, 16'd35676, 16'd10471, 16'd41542, 16'd46852, 16'd8371, 16'd29563, 16'd13377, 16'd13972, 16'd48139, 16'd45400, 16'd4600, 16'd57475, 16'd17820, 16'd36894, 16'd194, 16'd8762, 16'd40586, 16'd35011, 16'd20620, 16'd43107});
	test_expansion(128'hde027705eff511f970c09b7ade46ac7e, {16'd28435, 16'd32010, 16'd45689, 16'd59998, 16'd54958, 16'd35497, 16'd55635, 16'd55110, 16'd32460, 16'd5154, 16'd25659, 16'd65292, 16'd1602, 16'd59577, 16'd50534, 16'd4335, 16'd24977, 16'd38917, 16'd45495, 16'd44908, 16'd26193, 16'd4545, 16'd30488, 16'd42984, 16'd18740, 16'd3331});
	test_expansion(128'h84fec071d9c3e9946470af9165ff513d, {16'd40481, 16'd48099, 16'd17772, 16'd56909, 16'd15280, 16'd38573, 16'd1396, 16'd5568, 16'd25153, 16'd35287, 16'd39882, 16'd30881, 16'd26193, 16'd15494, 16'd7493, 16'd5678, 16'd18690, 16'd18421, 16'd18499, 16'd6014, 16'd12947, 16'd33732, 16'd52423, 16'd6837, 16'd64629, 16'd8964});
	test_expansion(128'hd289a2c058a531615f67615464f72098, {16'd13409, 16'd11418, 16'd22142, 16'd27624, 16'd32608, 16'd444, 16'd1216, 16'd62007, 16'd21481, 16'd16393, 16'd29344, 16'd43320, 16'd54841, 16'd11352, 16'd17253, 16'd26408, 16'd31885, 16'd17461, 16'd56295, 16'd9890, 16'd21444, 16'd13760, 16'd22122, 16'd24632, 16'd22586, 16'd24063});
	test_expansion(128'h1818b8b7f23b508cb5edff0f7f455ed4, {16'd11132, 16'd22098, 16'd22703, 16'd61283, 16'd195, 16'd18210, 16'd21472, 16'd48843, 16'd12366, 16'd34351, 16'd57945, 16'd20627, 16'd13270, 16'd63617, 16'd24551, 16'd48620, 16'd24390, 16'd3164, 16'd63138, 16'd17950, 16'd42070, 16'd46460, 16'd24721, 16'd22598, 16'd10052, 16'd50747});
	test_expansion(128'h4f266ef29e26eaac079dea6ddda6f165, {16'd10602, 16'd16737, 16'd15474, 16'd47244, 16'd15537, 16'd27401, 16'd54975, 16'd8448, 16'd43648, 16'd40055, 16'd14696, 16'd38494, 16'd28112, 16'd63519, 16'd29944, 16'd54220, 16'd18879, 16'd15054, 16'd58815, 16'd14871, 16'd8134, 16'd27729, 16'd60324, 16'd42558, 16'd1502, 16'd53077});
	test_expansion(128'hf8d6dd8df9436fb5c2669249380d2133, {16'd46136, 16'd59899, 16'd20763, 16'd46656, 16'd40601, 16'd44532, 16'd39521, 16'd33316, 16'd52111, 16'd49021, 16'd28769, 16'd13522, 16'd35973, 16'd19577, 16'd27744, 16'd28268, 16'd7424, 16'd60551, 16'd20876, 16'd32960, 16'd23433, 16'd40049, 16'd59858, 16'd51003, 16'd37491, 16'd31815});
	test_expansion(128'h0fafdd0260bcc174051c0c76e3246838, {16'd15381, 16'd62920, 16'd49777, 16'd48600, 16'd43299, 16'd42136, 16'd17161, 16'd58517, 16'd44824, 16'd86, 16'd57981, 16'd2373, 16'd15288, 16'd3829, 16'd12301, 16'd3821, 16'd3873, 16'd34686, 16'd46119, 16'd41850, 16'd21125, 16'd61719, 16'd60809, 16'd20467, 16'd42850, 16'd6678});
	test_expansion(128'hdc7c41e4305c475464050091d9c219df, {16'd26356, 16'd63814, 16'd519, 16'd33417, 16'd30765, 16'd41853, 16'd22117, 16'd38596, 16'd3292, 16'd18661, 16'd43198, 16'd3299, 16'd18146, 16'd44530, 16'd4009, 16'd34874, 16'd7889, 16'd58552, 16'd59062, 16'd46739, 16'd22948, 16'd27796, 16'd63716, 16'd47879, 16'd42020, 16'd58054});
	test_expansion(128'h7e3fba7a97ee4de8a563e93577db60fc, {16'd64430, 16'd24323, 16'd49867, 16'd28070, 16'd58227, 16'd14723, 16'd55479, 16'd10551, 16'd19347, 16'd21062, 16'd10683, 16'd28479, 16'd10335, 16'd43988, 16'd58726, 16'd65181, 16'd30977, 16'd21813, 16'd1120, 16'd1244, 16'd61912, 16'd24392, 16'd35363, 16'd33467, 16'd19814, 16'd6292});
	test_expansion(128'heec0c955f7ea03ffa7612a9cbb4a1376, {16'd37008, 16'd1865, 16'd40029, 16'd19656, 16'd34495, 16'd4585, 16'd36964, 16'd11443, 16'd535, 16'd11818, 16'd30665, 16'd1948, 16'd9848, 16'd10226, 16'd49540, 16'd41689, 16'd44312, 16'd31380, 16'd5270, 16'd14865, 16'd51758, 16'd35603, 16'd42392, 16'd7615, 16'd44894, 16'd44797});
	test_expansion(128'h24c4e347a9a044b2ba398fed36022ad9, {16'd10121, 16'd40151, 16'd35732, 16'd11351, 16'd4073, 16'd24993, 16'd51432, 16'd20599, 16'd17112, 16'd40240, 16'd36658, 16'd7717, 16'd62583, 16'd38346, 16'd46189, 16'd20413, 16'd9865, 16'd2853, 16'd45707, 16'd48363, 16'd35814, 16'd12802, 16'd19487, 16'd28276, 16'd6188, 16'd44201});
	test_expansion(128'h0809260e0711b22bf8fd25f04adc959b, {16'd23157, 16'd46536, 16'd20942, 16'd13408, 16'd12091, 16'd7724, 16'd33376, 16'd40884, 16'd39843, 16'd7900, 16'd12837, 16'd59656, 16'd23019, 16'd1273, 16'd47430, 16'd8795, 16'd14910, 16'd18334, 16'd62560, 16'd46519, 16'd44708, 16'd47836, 16'd1946, 16'd7426, 16'd53914, 16'd12477});
	test_expansion(128'h392b7b37023f0b0b70e6ba516fa8b95b, {16'd21992, 16'd25470, 16'd29653, 16'd17800, 16'd15207, 16'd144, 16'd1892, 16'd6515, 16'd9406, 16'd60933, 16'd50862, 16'd25280, 16'd23194, 16'd32613, 16'd62632, 16'd36135, 16'd21421, 16'd27834, 16'd8882, 16'd55499, 16'd16881, 16'd34920, 16'd44597, 16'd32792, 16'd49633, 16'd44741});
	test_expansion(128'h2dd01b34a00e7ba11219838b03e1aebb, {16'd22702, 16'd1597, 16'd63352, 16'd14248, 16'd20172, 16'd2376, 16'd47668, 16'd29288, 16'd34597, 16'd40996, 16'd47359, 16'd27547, 16'd64537, 16'd18251, 16'd3122, 16'd38066, 16'd31656, 16'd13567, 16'd55862, 16'd56162, 16'd23037, 16'd54955, 16'd34254, 16'd55519, 16'd34788, 16'd29578});
	test_expansion(128'h66ff18c00c9d0ba12df1beb58f239a06, {16'd35898, 16'd24781, 16'd18919, 16'd61515, 16'd9350, 16'd22628, 16'd24503, 16'd39812, 16'd23161, 16'd35326, 16'd56404, 16'd13720, 16'd50702, 16'd57484, 16'd56937, 16'd5789, 16'd53731, 16'd61451, 16'd41988, 16'd18253, 16'd59742, 16'd41436, 16'd17478, 16'd59061, 16'd53377, 16'd62033});
	test_expansion(128'h3974069abd8ba9ac884f3edabee1f9f9, {16'd14784, 16'd37736, 16'd50894, 16'd42101, 16'd1622, 16'd61567, 16'd6144, 16'd53118, 16'd42058, 16'd44883, 16'd21346, 16'd56813, 16'd12462, 16'd53580, 16'd60885, 16'd18084, 16'd23441, 16'd27547, 16'd14057, 16'd42480, 16'd26067, 16'd64304, 16'd65027, 16'd3559, 16'd53, 16'd18323});
	test_expansion(128'ha5a61ab843c54514f7805fffcd8a7ecd, {16'd24203, 16'd15540, 16'd52248, 16'd39467, 16'd47958, 16'd34095, 16'd59755, 16'd43477, 16'd19571, 16'd32884, 16'd42544, 16'd1556, 16'd33628, 16'd17001, 16'd14934, 16'd46278, 16'd9632, 16'd494, 16'd9688, 16'd40205, 16'd30977, 16'd24814, 16'd747, 16'd23000, 16'd28796, 16'd64799});
	test_expansion(128'h4e83674742203b8a6e7f4cfcb4e30e85, {16'd52395, 16'd29482, 16'd3488, 16'd52617, 16'd17234, 16'd24784, 16'd55660, 16'd48830, 16'd46753, 16'd46306, 16'd5785, 16'd13044, 16'd30572, 16'd45374, 16'd14417, 16'd56931, 16'd54977, 16'd32831, 16'd62335, 16'd31614, 16'd7014, 16'd6074, 16'd32691, 16'd34784, 16'd27231, 16'd155});
	test_expansion(128'hc34f16e59b7482bd44805c757835240b, {16'd56304, 16'd27890, 16'd62118, 16'd41075, 16'd14315, 16'd21847, 16'd43185, 16'd41155, 16'd45932, 16'd32109, 16'd42729, 16'd17220, 16'd24004, 16'd55638, 16'd33542, 16'd40726, 16'd6292, 16'd26428, 16'd49499, 16'd60357, 16'd34215, 16'd42573, 16'd40782, 16'd40810, 16'd63548, 16'd50697});
	test_expansion(128'ha75ffd3d114baae49b727775329c1847, {16'd8745, 16'd5509, 16'd12163, 16'd57574, 16'd63022, 16'd28369, 16'd20865, 16'd58204, 16'd57989, 16'd58196, 16'd16171, 16'd5982, 16'd58964, 16'd47495, 16'd9709, 16'd20709, 16'd62481, 16'd37042, 16'd55238, 16'd61657, 16'd3986, 16'd30883, 16'd9247, 16'd11146, 16'd52997, 16'd17135});
	test_expansion(128'hafede5f57b1d98cc9f19a700ec69d132, {16'd50350, 16'd56071, 16'd37667, 16'd11862, 16'd12274, 16'd33605, 16'd20931, 16'd55502, 16'd45272, 16'd42874, 16'd51857, 16'd2696, 16'd8397, 16'd22024, 16'd55978, 16'd48695, 16'd38205, 16'd40169, 16'd18914, 16'd33079, 16'd31024, 16'd11880, 16'd51669, 16'd47120, 16'd19379, 16'd18391});
	test_expansion(128'hbf5077b043d065dce92dbfb0412ff8a1, {16'd19600, 16'd12146, 16'd49942, 16'd44582, 16'd31945, 16'd46539, 16'd62161, 16'd24758, 16'd15802, 16'd53422, 16'd59614, 16'd17495, 16'd28979, 16'd24264, 16'd2242, 16'd34975, 16'd39719, 16'd64465, 16'd33766, 16'd7993, 16'd46782, 16'd65123, 16'd59653, 16'd18419, 16'd31810, 16'd55340});
	test_expansion(128'h3d68f5fba826dded85c05d1d9944922e, {16'd5487, 16'd39907, 16'd45588, 16'd45740, 16'd20336, 16'd59723, 16'd19755, 16'd60068, 16'd6152, 16'd49537, 16'd49599, 16'd6263, 16'd16281, 16'd18984, 16'd38217, 16'd39371, 16'd4328, 16'd10649, 16'd38484, 16'd36902, 16'd60351, 16'd27282, 16'd13441, 16'd59288, 16'd47309, 16'd40215});
	test_expansion(128'h7e0e76889e6870e08025691b43ac1154, {16'd40484, 16'd62445, 16'd50765, 16'd10112, 16'd28833, 16'd22405, 16'd34521, 16'd6320, 16'd45395, 16'd61488, 16'd28015, 16'd13691, 16'd5709, 16'd41862, 16'd63783, 16'd18469, 16'd34519, 16'd31378, 16'd44793, 16'd37369, 16'd44375, 16'd56927, 16'd59720, 16'd49287, 16'd1026, 16'd52830});
	test_expansion(128'h1380b47dc15a9f2a275bfbd3f2492e80, {16'd46420, 16'd12102, 16'd28987, 16'd25177, 16'd8597, 16'd31221, 16'd7864, 16'd6710, 16'd15410, 16'd38793, 16'd61115, 16'd8073, 16'd65000, 16'd54265, 16'd28633, 16'd3291, 16'd3692, 16'd409, 16'd5524, 16'd8274, 16'd56261, 16'd11883, 16'd30975, 16'd17679, 16'd2034, 16'd63473});
	test_expansion(128'he282ea94cfdb61a6694dc0157836cbf9, {16'd26383, 16'd14162, 16'd45318, 16'd16775, 16'd15643, 16'd30559, 16'd1948, 16'd37430, 16'd20342, 16'd44677, 16'd59925, 16'd40274, 16'd2541, 16'd5740, 16'd18909, 16'd39850, 16'd28203, 16'd53290, 16'd50173, 16'd57704, 16'd37401, 16'd56113, 16'd19424, 16'd8551, 16'd38215, 16'd13810});
	test_expansion(128'h8dd6bf8d00c84ff15d1d8a981ad517c1, {16'd8115, 16'd22859, 16'd45909, 16'd62822, 16'd50587, 16'd18543, 16'd59698, 16'd38569, 16'd27058, 16'd32273, 16'd27066, 16'd11591, 16'd42955, 16'd3303, 16'd14743, 16'd24440, 16'd53362, 16'd30590, 16'd22897, 16'd35504, 16'd55227, 16'd31069, 16'd30015, 16'd63377, 16'd32958, 16'd34984});
	test_expansion(128'h0930dc77269b7cf45debc836723ba909, {16'd60103, 16'd17090, 16'd31538, 16'd57841, 16'd23651, 16'd28659, 16'd7817, 16'd48333, 16'd47342, 16'd50939, 16'd40784, 16'd62947, 16'd26362, 16'd32219, 16'd11898, 16'd225, 16'd30569, 16'd54784, 16'd64710, 16'd49026, 16'd24892, 16'd33730, 16'd58997, 16'd9709, 16'd52581, 16'd61289});
	test_expansion(128'hc430bcdeee6b1035aa7ec9b10e1a3789, {16'd50075, 16'd31942, 16'd28148, 16'd55647, 16'd33784, 16'd32844, 16'd51850, 16'd38598, 16'd30323, 16'd25270, 16'd60471, 16'd54135, 16'd34416, 16'd45699, 16'd27734, 16'd52732, 16'd38730, 16'd52308, 16'd56363, 16'd28448, 16'd48909, 16'd12246, 16'd10024, 16'd6536, 16'd14273, 16'd53428});
	test_expansion(128'h03eb7d26cae9b0bc5294959855440df5, {16'd47266, 16'd49044, 16'd51602, 16'd49397, 16'd61811, 16'd40023, 16'd58864, 16'd39202, 16'd53124, 16'd51030, 16'd49388, 16'd41785, 16'd51335, 16'd27287, 16'd21395, 16'd38747, 16'd55618, 16'd42516, 16'd14722, 16'd42085, 16'd59222, 16'd53716, 16'd47523, 16'd1047, 16'd61554, 16'd59014});
	test_expansion(128'hf85de800026ce63a21a23470323aa784, {16'd33877, 16'd61284, 16'd26701, 16'd20664, 16'd33084, 16'd57452, 16'd53444, 16'd57084, 16'd9571, 16'd32316, 16'd42506, 16'd49276, 16'd40929, 16'd44892, 16'd34293, 16'd44950, 16'd12984, 16'd17522, 16'd44498, 16'd46707, 16'd51045, 16'd63853, 16'd32719, 16'd56981, 16'd64422, 16'd24615});
	test_expansion(128'h2fc18cbfe48d0929dd82907cfcf81de9, {16'd61545, 16'd52857, 16'd47551, 16'd18648, 16'd16638, 16'd2348, 16'd45099, 16'd29865, 16'd33682, 16'd29512, 16'd3232, 16'd26227, 16'd15089, 16'd41208, 16'd26446, 16'd950, 16'd20700, 16'd51121, 16'd64, 16'd7725, 16'd58147, 16'd61187, 16'd38054, 16'd11644, 16'd59839, 16'd17646});
	test_expansion(128'h30c8fa1af3066a6cc29d3931b8d9473b, {16'd61130, 16'd65396, 16'd21889, 16'd5410, 16'd45856, 16'd27139, 16'd17776, 16'd10408, 16'd28079, 16'd13220, 16'd60090, 16'd56836, 16'd36094, 16'd4232, 16'd32281, 16'd60123, 16'd40711, 16'd927, 16'd11871, 16'd56448, 16'd33442, 16'd12490, 16'd55323, 16'd10466, 16'd25031, 16'd22113});
	test_expansion(128'h083f4bba1644fe1082ab51e38c0b100c, {16'd20533, 16'd50610, 16'd40975, 16'd38083, 16'd24158, 16'd31833, 16'd53083, 16'd15530, 16'd40732, 16'd21647, 16'd26316, 16'd32143, 16'd53885, 16'd9656, 16'd36858, 16'd30820, 16'd45656, 16'd36173, 16'd47730, 16'd8216, 16'd50924, 16'd41921, 16'd8156, 16'd2658, 16'd36821, 16'd61560});
	test_expansion(128'hf2adaabdb48a006341147ddcb9a4bd14, {16'd4164, 16'd42801, 16'd51635, 16'd58893, 16'd8059, 16'd44143, 16'd39056, 16'd18125, 16'd1331, 16'd29198, 16'd18559, 16'd53199, 16'd33329, 16'd53307, 16'd49922, 16'd4003, 16'd22869, 16'd47817, 16'd658, 16'd24759, 16'd7722, 16'd63723, 16'd36299, 16'd42421, 16'd39711, 16'd3151});
	test_expansion(128'h373d947be225242ecd7e6f2866a1f272, {16'd9732, 16'd1652, 16'd2650, 16'd60670, 16'd19837, 16'd38703, 16'd22020, 16'd26763, 16'd31762, 16'd65524, 16'd3816, 16'd1387, 16'd45459, 16'd6323, 16'd51645, 16'd1300, 16'd27227, 16'd38808, 16'd980, 16'd11554, 16'd32011, 16'd21676, 16'd26915, 16'd7887, 16'd43883, 16'd9092});
	test_expansion(128'hee8f64c7142113a370bb3f5ced22b847, {16'd50607, 16'd53571, 16'd8343, 16'd42388, 16'd10512, 16'd35165, 16'd14243, 16'd5908, 16'd64030, 16'd32657, 16'd53452, 16'd32513, 16'd36517, 16'd13894, 16'd13219, 16'd44048, 16'd47188, 16'd54521, 16'd16314, 16'd22489, 16'd23222, 16'd41328, 16'd13073, 16'd63252, 16'd16348, 16'd50905});
	test_expansion(128'hdcf509a90330bc2024d724e8d44ae83b, {16'd5861, 16'd27928, 16'd7089, 16'd6265, 16'd19739, 16'd64406, 16'd23527, 16'd57270, 16'd28137, 16'd14810, 16'd24646, 16'd10261, 16'd24470, 16'd61379, 16'd2199, 16'd14685, 16'd44038, 16'd44666, 16'd14783, 16'd7162, 16'd64483, 16'd32580, 16'd21002, 16'd63923, 16'd18696, 16'd7738});
	test_expansion(128'h521175dd0eaf155d9297b744f15e8c35, {16'd21463, 16'd64417, 16'd44266, 16'd43841, 16'd43576, 16'd43420, 16'd55793, 16'd28187, 16'd11057, 16'd37646, 16'd18315, 16'd54647, 16'd38499, 16'd60621, 16'd55404, 16'd60770, 16'd15407, 16'd6692, 16'd23642, 16'd45175, 16'd28202, 16'd31519, 16'd53801, 16'd5512, 16'd9790, 16'd42394});
	test_expansion(128'h87e7dea85f4bc8f8b536ed0cff6e991a, {16'd39148, 16'd24900, 16'd23819, 16'd6849, 16'd36194, 16'd21801, 16'd54921, 16'd18451, 16'd2982, 16'd29068, 16'd49983, 16'd18990, 16'd52887, 16'd20043, 16'd16345, 16'd42149, 16'd12029, 16'd18921, 16'd5847, 16'd22234, 16'd1696, 16'd65464, 16'd61068, 16'd28561, 16'd27808, 16'd28190});
	test_expansion(128'hd00a3a69c19b5d559464ee6f8395edc6, {16'd17014, 16'd8236, 16'd52698, 16'd41990, 16'd317, 16'd16148, 16'd50116, 16'd23075, 16'd41570, 16'd24998, 16'd14224, 16'd1702, 16'd12835, 16'd32907, 16'd28866, 16'd61879, 16'd57917, 16'd30337, 16'd7165, 16'd12693, 16'd19560, 16'd7373, 16'd47943, 16'd45776, 16'd4565, 16'd57366});
	test_expansion(128'h8b282e61dd815ba136a9ea6433e69245, {16'd34666, 16'd52546, 16'd46433, 16'd28397, 16'd58761, 16'd42943, 16'd15654, 16'd36606, 16'd36245, 16'd50236, 16'd44918, 16'd7136, 16'd38828, 16'd34614, 16'd8034, 16'd41256, 16'd64079, 16'd3732, 16'd32133, 16'd47662, 16'd52538, 16'd4939, 16'd23033, 16'd30922, 16'd49503, 16'd34950});
	test_expansion(128'h17247efda72f86e3cf7d3834528f712c, {16'd47415, 16'd25283, 16'd5129, 16'd21985, 16'd56675, 16'd397, 16'd51610, 16'd41241, 16'd41822, 16'd7945, 16'd31438, 16'd23012, 16'd64720, 16'd2098, 16'd60864, 16'd64897, 16'd43308, 16'd38101, 16'd23771, 16'd64807, 16'd12936, 16'd65254, 16'd4828, 16'd63280, 16'd19357, 16'd53280});
	test_expansion(128'h52fc17c6ac75d67cf68b5036b0a6ccad, {16'd42965, 16'd6072, 16'd49066, 16'd7309, 16'd59103, 16'd14109, 16'd47469, 16'd511, 16'd49356, 16'd376, 16'd64778, 16'd53248, 16'd50724, 16'd43039, 16'd29435, 16'd22497, 16'd24813, 16'd921, 16'd47178, 16'd35141, 16'd62527, 16'd21156, 16'd32214, 16'd50139, 16'd18661, 16'd47514});
	test_expansion(128'hb656e5aac649ba8a7cdecb48fa870283, {16'd51469, 16'd8348, 16'd63220, 16'd64341, 16'd23583, 16'd28195, 16'd58364, 16'd23075, 16'd35450, 16'd18888, 16'd32661, 16'd1976, 16'd3018, 16'd8297, 16'd7664, 16'd46746, 16'd13198, 16'd7294, 16'd15494, 16'd59617, 16'd1581, 16'd32029, 16'd61801, 16'd26749, 16'd2877, 16'd37658});
	test_expansion(128'h481afb8c71d9e28055027d611f320564, {16'd53643, 16'd2741, 16'd10406, 16'd40857, 16'd42163, 16'd35311, 16'd19847, 16'd34788, 16'd35680, 16'd9926, 16'd58642, 16'd63956, 16'd7214, 16'd41885, 16'd14623, 16'd39866, 16'd17734, 16'd4595, 16'd10836, 16'd33672, 16'd24426, 16'd32545, 16'd63829, 16'd52157, 16'd3658, 16'd52903});
	test_expansion(128'h364636402fcbe45038470b520612c537, {16'd46203, 16'd50672, 16'd57665, 16'd11853, 16'd957, 16'd13746, 16'd12082, 16'd939, 16'd49894, 16'd4740, 16'd8473, 16'd44289, 16'd18729, 16'd65032, 16'd13436, 16'd21579, 16'd7563, 16'd908, 16'd10416, 16'd46743, 16'd53371, 16'd9665, 16'd34267, 16'd29963, 16'd8759, 16'd10254});
	test_expansion(128'hcbadc78f50a50690ab5a674e1dc4d20d, {16'd27046, 16'd63752, 16'd14176, 16'd55384, 16'd64281, 16'd45015, 16'd26258, 16'd34235, 16'd4893, 16'd16548, 16'd34826, 16'd973, 16'd15567, 16'd33749, 16'd65321, 16'd47510, 16'd56506, 16'd28574, 16'd11983, 16'd60135, 16'd64979, 16'd63857, 16'd65086, 16'd14160, 16'd62200, 16'd54519});
	test_expansion(128'ha4df5d424ed366285f71f419b7cbfea1, {16'd24106, 16'd34365, 16'd34260, 16'd26687, 16'd19630, 16'd28506, 16'd43000, 16'd3110, 16'd890, 16'd47403, 16'd3490, 16'd64167, 16'd33000, 16'd23073, 16'd12782, 16'd3683, 16'd60810, 16'd36893, 16'd58266, 16'd42262, 16'd13905, 16'd53566, 16'd1172, 16'd65258, 16'd687, 16'd49681});
	test_expansion(128'h97f948b31eaccda21accceb033d43fa3, {16'd57638, 16'd43573, 16'd62165, 16'd5867, 16'd9892, 16'd10243, 16'd15773, 16'd52034, 16'd55453, 16'd440, 16'd63565, 16'd57886, 16'd11257, 16'd60294, 16'd25159, 16'd41044, 16'd25727, 16'd45345, 16'd41549, 16'd58108, 16'd47733, 16'd16935, 16'd35571, 16'd31448, 16'd14489, 16'd36615});
	test_expansion(128'h64450a5032ea054657d71fb635fcbdda, {16'd4893, 16'd28354, 16'd17789, 16'd52757, 16'd23291, 16'd5263, 16'd54730, 16'd18012, 16'd42414, 16'd30556, 16'd21621, 16'd15172, 16'd47479, 16'd8966, 16'd19664, 16'd21379, 16'd58518, 16'd31968, 16'd65167, 16'd33605, 16'd20776, 16'd7354, 16'd8648, 16'd46200, 16'd3601, 16'd32186});
	test_expansion(128'h1d814a6efe194468863885a2efa42425, {16'd39447, 16'd52194, 16'd7722, 16'd49244, 16'd47195, 16'd20664, 16'd42451, 16'd51258, 16'd7826, 16'd43785, 16'd21856, 16'd898, 16'd41843, 16'd48592, 16'd26804, 16'd39782, 16'd13517, 16'd36300, 16'd46141, 16'd46029, 16'd9195, 16'd48204, 16'd48169, 16'd20967, 16'd22530, 16'd36895});
	test_expansion(128'hb19da0fbd33acd606e0fbec6841f82c5, {16'd15882, 16'd25521, 16'd47367, 16'd21724, 16'd39658, 16'd29128, 16'd17287, 16'd50242, 16'd43976, 16'd2351, 16'd19772, 16'd28139, 16'd37695, 16'd62355, 16'd35870, 16'd6358, 16'd53505, 16'd16223, 16'd23028, 16'd14639, 16'd864, 16'd24798, 16'd52417, 16'd17060, 16'd47116, 16'd18256});
	test_expansion(128'h49b2fc19ed2615351dc50f779d66ec83, {16'd36936, 16'd55741, 16'd23928, 16'd24430, 16'd54159, 16'd10171, 16'd27822, 16'd12410, 16'd29792, 16'd14430, 16'd5520, 16'd64400, 16'd21300, 16'd26709, 16'd58329, 16'd4044, 16'd8434, 16'd2688, 16'd4715, 16'd57284, 16'd43766, 16'd30488, 16'd60633, 16'd20062, 16'd9290, 16'd63669});
	test_expansion(128'he3922792c1b40e59222afe30aade38b5, {16'd18547, 16'd13011, 16'd22385, 16'd48966, 16'd64154, 16'd36263, 16'd39175, 16'd53019, 16'd47093, 16'd9662, 16'd53856, 16'd58554, 16'd60241, 16'd11897, 16'd60005, 16'd14703, 16'd15309, 16'd44012, 16'd42282, 16'd43798, 16'd13896, 16'd53079, 16'd36060, 16'd15158, 16'd11544, 16'd63230});
	test_expansion(128'heaa982957ff10128388d5d65dc19fb81, {16'd29165, 16'd47832, 16'd9024, 16'd32412, 16'd19302, 16'd46118, 16'd2635, 16'd25089, 16'd24287, 16'd60821, 16'd60500, 16'd45109, 16'd8557, 16'd31991, 16'd53612, 16'd31752, 16'd24294, 16'd26109, 16'd50174, 16'd31315, 16'd2539, 16'd53513, 16'd52642, 16'd38000, 16'd17427, 16'd24600});
	test_expansion(128'h0dc3cf9da97e899bf05e9343e5af6c3f, {16'd1060, 16'd37220, 16'd10978, 16'd60161, 16'd18604, 16'd45737, 16'd6036, 16'd21125, 16'd44201, 16'd27145, 16'd19893, 16'd22880, 16'd47583, 16'd15767, 16'd30876, 16'd16407, 16'd44574, 16'd11460, 16'd977, 16'd48628, 16'd23892, 16'd44396, 16'd10453, 16'd23493, 16'd33057, 16'd53076});
	test_expansion(128'h6f4527933574fc5ed1a89299e354006b, {16'd6556, 16'd20147, 16'd41607, 16'd43202, 16'd38323, 16'd28748, 16'd10341, 16'd65071, 16'd3153, 16'd30693, 16'd1270, 16'd22625, 16'd62820, 16'd22893, 16'd47334, 16'd45042, 16'd50355, 16'd28815, 16'd54517, 16'd4735, 16'd32506, 16'd51946, 16'd25525, 16'd30278, 16'd11036, 16'd11130});
	test_expansion(128'h80e07aee19d51b5f5d7019261cf2fb5a, {16'd25759, 16'd37512, 16'd55302, 16'd7602, 16'd15543, 16'd49193, 16'd44105, 16'd5786, 16'd33395, 16'd55817, 16'd27759, 16'd50169, 16'd44083, 16'd37892, 16'd26098, 16'd6217, 16'd21037, 16'd30998, 16'd40687, 16'd969, 16'd26865, 16'd63591, 16'd46322, 16'd45988, 16'd47931, 16'd62280});
	test_expansion(128'h92c40eaabd2aac3691cec8cc746e8630, {16'd19324, 16'd47116, 16'd3825, 16'd55357, 16'd64299, 16'd12827, 16'd45841, 16'd51576, 16'd3160, 16'd29185, 16'd31614, 16'd49674, 16'd52743, 16'd44636, 16'd49771, 16'd59203, 16'd30520, 16'd47437, 16'd10655, 16'd40361, 16'd58147, 16'd61401, 16'd46338, 16'd41033, 16'd55254, 16'd27378});
	test_expansion(128'h5f55a3f2c3f41a4fcbb92c2df4fec365, {16'd40526, 16'd61354, 16'd22146, 16'd27989, 16'd9992, 16'd57350, 16'd61146, 16'd45102, 16'd56983, 16'd22302, 16'd8095, 16'd46862, 16'd16584, 16'd3699, 16'd63392, 16'd31817, 16'd16515, 16'd37645, 16'd12904, 16'd12840, 16'd4330, 16'd47144, 16'd45237, 16'd25354, 16'd25626, 16'd24207});
	test_expansion(128'he44b9764fb9161ac24f461d515648bf0, {16'd2812, 16'd14021, 16'd12662, 16'd25125, 16'd62599, 16'd29559, 16'd52947, 16'd58282, 16'd46222, 16'd33706, 16'd2198, 16'd44879, 16'd56938, 16'd63264, 16'd42963, 16'd36791, 16'd2130, 16'd2080, 16'd55766, 16'd56975, 16'd21555, 16'd63806, 16'd51492, 16'd15901, 16'd56504, 16'd17892});
	test_expansion(128'hf2fce63661b72fc70d6e8bde74488d41, {16'd11749, 16'd45582, 16'd24896, 16'd57603, 16'd1629, 16'd45992, 16'd26548, 16'd31347, 16'd51748, 16'd34028, 16'd1343, 16'd59510, 16'd23430, 16'd37680, 16'd45406, 16'd64336, 16'd42266, 16'd54817, 16'd19754, 16'd17834, 16'd23592, 16'd40228, 16'd2212, 16'd34132, 16'd3435, 16'd22281});
	test_expansion(128'h49c3bb1780a6c6553567f59c73989ac0, {16'd55957, 16'd28465, 16'd59700, 16'd18686, 16'd5639, 16'd49999, 16'd57243, 16'd37910, 16'd44140, 16'd19184, 16'd49319, 16'd46812, 16'd52737, 16'd51562, 16'd32310, 16'd6549, 16'd10822, 16'd64468, 16'd16047, 16'd57080, 16'd3272, 16'd47916, 16'd41741, 16'd4199, 16'd40179, 16'd35748});
	test_expansion(128'ha070dfe174c37c2369eb11574e9a72e4, {16'd63987, 16'd3503, 16'd38956, 16'd2631, 16'd55095, 16'd25509, 16'd3249, 16'd47306, 16'd6030, 16'd39963, 16'd14899, 16'd59980, 16'd29164, 16'd43391, 16'd53955, 16'd42924, 16'd24805, 16'd57121, 16'd63771, 16'd48383, 16'd45568, 16'd3546, 16'd40759, 16'd14067, 16'd42957, 16'd42723});
	test_expansion(128'h6c1539cac3e73ef226174b6eeb109ee6, {16'd41359, 16'd45603, 16'd54178, 16'd10178, 16'd16006, 16'd29076, 16'd60291, 16'd30926, 16'd37463, 16'd22282, 16'd49344, 16'd22549, 16'd20999, 16'd11683, 16'd31660, 16'd9054, 16'd48103, 16'd25247, 16'd8681, 16'd1985, 16'd5891, 16'd4001, 16'd20425, 16'd39256, 16'd64692, 16'd64721});
	test_expansion(128'h9badce08e4c20746f27c131af78ee66d, {16'd26420, 16'd42772, 16'd49400, 16'd17997, 16'd34393, 16'd11683, 16'd48968, 16'd16207, 16'd53322, 16'd39645, 16'd23350, 16'd48589, 16'd41935, 16'd34768, 16'd10202, 16'd18083, 16'd35761, 16'd35194, 16'd43741, 16'd40355, 16'd41808, 16'd21044, 16'd43929, 16'd44513, 16'd60627, 16'd15476});
	test_expansion(128'h3ecc2e715e6881edb630dcdb782cf4d5, {16'd23615, 16'd55200, 16'd64529, 16'd26786, 16'd175, 16'd54442, 16'd51809, 16'd50518, 16'd60753, 16'd10007, 16'd23161, 16'd37127, 16'd52451, 16'd33184, 16'd61588, 16'd41897, 16'd11333, 16'd5913, 16'd32507, 16'd40757, 16'd15157, 16'd39673, 16'd52641, 16'd63253, 16'd39572, 16'd45694});
	test_expansion(128'h6e5378084ad51d55d7f5e3c45c7c9bcd, {16'd57363, 16'd4994, 16'd43284, 16'd32729, 16'd53185, 16'd44645, 16'd40542, 16'd50997, 16'd41829, 16'd52206, 16'd38878, 16'd58352, 16'd51088, 16'd51147, 16'd45355, 16'd54475, 16'd54845, 16'd19584, 16'd36455, 16'd31029, 16'd4390, 16'd6798, 16'd57144, 16'd22137, 16'd11079, 16'd46920});
	test_expansion(128'he56641ec87067fa6815ae74fe79f7372, {16'd30968, 16'd60427, 16'd61813, 16'd61872, 16'd17175, 16'd24896, 16'd13294, 16'd12204, 16'd48817, 16'd46557, 16'd33576, 16'd50733, 16'd99, 16'd45935, 16'd7130, 16'd25110, 16'd14454, 16'd61903, 16'd167, 16'd56347, 16'd26275, 16'd38659, 16'd7316, 16'd18757, 16'd34708, 16'd12170});
	test_expansion(128'hcbbd593bfe79e1aca5eb2e794331c6cc, {16'd52896, 16'd3342, 16'd61691, 16'd15374, 16'd26675, 16'd14597, 16'd9293, 16'd45616, 16'd43660, 16'd10944, 16'd36391, 16'd56441, 16'd7636, 16'd49080, 16'd32020, 16'd7379, 16'd19568, 16'd40114, 16'd29159, 16'd38688, 16'd52964, 16'd57402, 16'd21267, 16'd22242, 16'd41784, 16'd38197});
	test_expansion(128'h86c95eb30437a8e4bafa61f1f0f2d25d, {16'd55759, 16'd54918, 16'd27074, 16'd11709, 16'd15076, 16'd26352, 16'd11724, 16'd31451, 16'd27663, 16'd11070, 16'd37442, 16'd48480, 16'd51714, 16'd64900, 16'd11182, 16'd21247, 16'd21113, 16'd61442, 16'd8998, 16'd5067, 16'd58582, 16'd49260, 16'd49281, 16'd30078, 16'd59521, 16'd43137});
	test_expansion(128'h6f51be8ce09fdcd9d2b7788ba574205c, {16'd27837, 16'd2033, 16'd1440, 16'd41428, 16'd32412, 16'd32892, 16'd58689, 16'd13813, 16'd59650, 16'd43925, 16'd53624, 16'd30783, 16'd43749, 16'd24329, 16'd45579, 16'd36016, 16'd28507, 16'd38293, 16'd14965, 16'd32642, 16'd45555, 16'd17004, 16'd21228, 16'd39893, 16'd37774, 16'd16043});
	test_expansion(128'h2a89902ff80c2b95ea0e2ddb7ebc429e, {16'd64749, 16'd60095, 16'd11800, 16'd4246, 16'd44812, 16'd63625, 16'd25204, 16'd25225, 16'd44510, 16'd49505, 16'd22234, 16'd28489, 16'd7996, 16'd55718, 16'd26762, 16'd9783, 16'd27753, 16'd1745, 16'd11124, 16'd54782, 16'd61711, 16'd12197, 16'd38558, 16'd43355, 16'd59182, 16'd54808});
	test_expansion(128'hc2a9e5495f9a66bdc1c470eaa3c484d4, {16'd27324, 16'd53363, 16'd36823, 16'd38176, 16'd63052, 16'd6166, 16'd61331, 16'd14037, 16'd46984, 16'd36334, 16'd48274, 16'd53079, 16'd25313, 16'd4066, 16'd50342, 16'd61027, 16'd59414, 16'd10272, 16'd15490, 16'd25881, 16'd43964, 16'd6435, 16'd61699, 16'd43510, 16'd22584, 16'd62721});
	test_expansion(128'h72769b037ed314b7ad5147c96a50cfba, {16'd37404, 16'd8445, 16'd5879, 16'd9411, 16'd56633, 16'd20937, 16'd54344, 16'd16654, 16'd5413, 16'd64617, 16'd45869, 16'd15567, 16'd56817, 16'd29976, 16'd23664, 16'd29291, 16'd34944, 16'd2179, 16'd1999, 16'd5661, 16'd2014, 16'd14450, 16'd9011, 16'd31365, 16'd14828, 16'd3338});
	test_expansion(128'hbfb113c866e25c69182bf0118b362328, {16'd2976, 16'd22652, 16'd20639, 16'd56659, 16'd44298, 16'd7759, 16'd24901, 16'd60082, 16'd21969, 16'd39320, 16'd53115, 16'd29477, 16'd56097, 16'd24710, 16'd54961, 16'd36571, 16'd38195, 16'd53924, 16'd13036, 16'd3507, 16'd39548, 16'd23637, 16'd64629, 16'd549, 16'd44386, 16'd46728});
	test_expansion(128'haa7269fa6550c77f3801e0efe6e451d6, {16'd8600, 16'd36186, 16'd42049, 16'd43010, 16'd15216, 16'd15627, 16'd33245, 16'd12139, 16'd1851, 16'd56562, 16'd32900, 16'd6254, 16'd63327, 16'd59777, 16'd65214, 16'd24466, 16'd47269, 16'd1344, 16'd23080, 16'd19569, 16'd19674, 16'd45694, 16'd33145, 16'd31196, 16'd1096, 16'd56298});
	test_expansion(128'he5fafc0665ead31c5d33ce6a73ffabfd, {16'd48303, 16'd45102, 16'd17149, 16'd49336, 16'd26338, 16'd30965, 16'd38124, 16'd62279, 16'd30678, 16'd25396, 16'd63990, 16'd64784, 16'd4845, 16'd20707, 16'd20677, 16'd50879, 16'd23672, 16'd8084, 16'd63967, 16'd2480, 16'd9086, 16'd33151, 16'd6748, 16'd52617, 16'd39673, 16'd46035});
	test_expansion(128'h0f2b4046d6a0d1429e4de5fece76f7f3, {16'd59547, 16'd3162, 16'd15486, 16'd58365, 16'd23424, 16'd40847, 16'd42463, 16'd37540, 16'd19754, 16'd6000, 16'd48232, 16'd14527, 16'd23789, 16'd16155, 16'd35647, 16'd4461, 16'd15232, 16'd48955, 16'd34086, 16'd20566, 16'd11009, 16'd28138, 16'd28924, 16'd4506, 16'd14443, 16'd37421});
	test_expansion(128'h0f44f389357ce5c3ee44e3293dea8c90, {16'd21637, 16'd2099, 16'd35850, 16'd58186, 16'd27875, 16'd45399, 16'd48185, 16'd18732, 16'd51913, 16'd63465, 16'd55113, 16'd34444, 16'd32085, 16'd23557, 16'd48462, 16'd56544, 16'd56431, 16'd21071, 16'd34146, 16'd9477, 16'd42435, 16'd20755, 16'd28200, 16'd44346, 16'd12680, 16'd24653});
	test_expansion(128'hbc349a2bbb233b8a47a5933ddb91de53, {16'd34354, 16'd16799, 16'd6259, 16'd50392, 16'd1638, 16'd61800, 16'd59506, 16'd55874, 16'd59566, 16'd55250, 16'd306, 16'd29118, 16'd41967, 16'd42751, 16'd28688, 16'd58920, 16'd51556, 16'd54579, 16'd22490, 16'd31735, 16'd35980, 16'd9093, 16'd13693, 16'd57396, 16'd65192, 16'd21362});
	test_expansion(128'hb8b59e86640cf81a78f3873b16a2efe1, {16'd28230, 16'd37475, 16'd35096, 16'd65291, 16'd15870, 16'd3399, 16'd64065, 16'd45572, 16'd60915, 16'd25965, 16'd64957, 16'd1433, 16'd39649, 16'd63967, 16'd19663, 16'd63404, 16'd3618, 16'd49642, 16'd2801, 16'd8240, 16'd13903, 16'd54233, 16'd48355, 16'd16075, 16'd1870, 16'd14455});
	test_expansion(128'h59de9164189532d4acc5be248618edc3, {16'd32534, 16'd27751, 16'd14815, 16'd18216, 16'd23364, 16'd19409, 16'd55033, 16'd47946, 16'd43168, 16'd33936, 16'd15575, 16'd31418, 16'd40434, 16'd61961, 16'd49776, 16'd10982, 16'd55836, 16'd50387, 16'd4728, 16'd30188, 16'd31260, 16'd24957, 16'd33008, 16'd15249, 16'd43199, 16'd19374});
	test_expansion(128'h2a7d327b747bb035702289c3159c1d51, {16'd16547, 16'd58675, 16'd16875, 16'd7622, 16'd3381, 16'd39497, 16'd7665, 16'd13917, 16'd35021, 16'd15355, 16'd8935, 16'd57897, 16'd48169, 16'd15947, 16'd27539, 16'd51489, 16'd25015, 16'd22530, 16'd51454, 16'd61158, 16'd36423, 16'd6599, 16'd53275, 16'd13053, 16'd12784, 16'd33192});
	test_expansion(128'h92c809dd215e13f38825bbb3b3eb521f, {16'd23240, 16'd14922, 16'd20036, 16'd37792, 16'd34165, 16'd46281, 16'd47017, 16'd30001, 16'd31506, 16'd42767, 16'd64879, 16'd7020, 16'd55050, 16'd8017, 16'd35686, 16'd13559, 16'd26121, 16'd10973, 16'd24734, 16'd53108, 16'd37990, 16'd36805, 16'd9436, 16'd37060, 16'd32781, 16'd44800});
	test_expansion(128'h311118cfd39df3e0df1c68eca75eedd7, {16'd8407, 16'd31791, 16'd40558, 16'd50837, 16'd54718, 16'd31170, 16'd45472, 16'd21111, 16'd40142, 16'd678, 16'd13547, 16'd63584, 16'd35177, 16'd8263, 16'd55997, 16'd47614, 16'd6105, 16'd11587, 16'd49056, 16'd65280, 16'd51341, 16'd50219, 16'd44693, 16'd60658, 16'd49740, 16'd51});
	test_expansion(128'h0a43231e2a62b7e2507d111dd62ada41, {16'd65454, 16'd26305, 16'd41661, 16'd33872, 16'd41855, 16'd55022, 16'd58753, 16'd21122, 16'd16606, 16'd12516, 16'd1135, 16'd19949, 16'd45303, 16'd26894, 16'd40113, 16'd29145, 16'd30569, 16'd47619, 16'd54504, 16'd51483, 16'd36050, 16'd64546, 16'd40203, 16'd57998, 16'd46387, 16'd17869});
	test_expansion(128'ha41fd408c8ac2778f8274d6aa69dc736, {16'd43514, 16'd27177, 16'd6256, 16'd38417, 16'd36671, 16'd45538, 16'd64922, 16'd61096, 16'd43990, 16'd33763, 16'd20751, 16'd17428, 16'd16866, 16'd28288, 16'd38247, 16'd39289, 16'd59815, 16'd6190, 16'd60366, 16'd34734, 16'd13601, 16'd14460, 16'd26401, 16'd16040, 16'd9277, 16'd14209});
	test_expansion(128'h6168979702a15a149f85846e0a196134, {16'd4088, 16'd16949, 16'd25202, 16'd25759, 16'd30191, 16'd45450, 16'd42613, 16'd52278, 16'd62403, 16'd21632, 16'd51729, 16'd37181, 16'd11138, 16'd11744, 16'd16851, 16'd23037, 16'd64173, 16'd37060, 16'd11662, 16'd30523, 16'd29682, 16'd13904, 16'd45246, 16'd44038, 16'd42648, 16'd45697});
	test_expansion(128'h87b32ec83e5492cdb032ae2dc8d25a73, {16'd36101, 16'd35593, 16'd25018, 16'd26319, 16'd45354, 16'd6688, 16'd59565, 16'd39047, 16'd57571, 16'd42363, 16'd47093, 16'd46762, 16'd48533, 16'd35033, 16'd29048, 16'd39387, 16'd29495, 16'd56696, 16'd62358, 16'd10406, 16'd12453, 16'd29912, 16'd15358, 16'd36275, 16'd10218, 16'd25129});
	test_expansion(128'hd7a604105bf718f9de67f66667a82bbc, {16'd38736, 16'd57314, 16'd25269, 16'd10162, 16'd27889, 16'd64461, 16'd38218, 16'd52406, 16'd32181, 16'd52280, 16'd31049, 16'd24650, 16'd33578, 16'd4584, 16'd63354, 16'd44647, 16'd33353, 16'd40942, 16'd64859, 16'd53023, 16'd56646, 16'd44034, 16'd46748, 16'd1666, 16'd10883, 16'd10606});
	test_expansion(128'h79f7e9b76e802c20d5f8eb174c394eb2, {16'd35436, 16'd35743, 16'd10576, 16'd21890, 16'd21040, 16'd34825, 16'd20087, 16'd27360, 16'd49590, 16'd58954, 16'd35394, 16'd26258, 16'd62115, 16'd17556, 16'd47162, 16'd30708, 16'd60110, 16'd24617, 16'd41865, 16'd1850, 16'd18583, 16'd8497, 16'd47451, 16'd40849, 16'd52355, 16'd19731});
	test_expansion(128'hae2b5e2a65268236345ec00525c4fe49, {16'd20068, 16'd64221, 16'd48733, 16'd15748, 16'd1294, 16'd10817, 16'd25164, 16'd38912, 16'd39892, 16'd50010, 16'd10410, 16'd1331, 16'd50528, 16'd53581, 16'd2187, 16'd55852, 16'd1539, 16'd9669, 16'd12602, 16'd9958, 16'd19235, 16'd1163, 16'd16164, 16'd16567, 16'd12879, 16'd39740});
	test_expansion(128'h20b01fed06089f51b74d06823ca2a3ea, {16'd63344, 16'd14673, 16'd3372, 16'd10475, 16'd26386, 16'd40949, 16'd30920, 16'd19489, 16'd45569, 16'd6586, 16'd36417, 16'd47474, 16'd58774, 16'd47679, 16'd41791, 16'd2950, 16'd21557, 16'd19513, 16'd3317, 16'd49029, 16'd50977, 16'd64662, 16'd4601, 16'd61002, 16'd14182, 16'd23046});
	test_expansion(128'ha4f2d42905dcfb7807406dca1368009c, {16'd52748, 16'd54693, 16'd53943, 16'd44612, 16'd2683, 16'd49149, 16'd29480, 16'd59071, 16'd36357, 16'd20574, 16'd58541, 16'd53903, 16'd62594, 16'd32549, 16'd56671, 16'd41461, 16'd7881, 16'd8234, 16'd22731, 16'd35371, 16'd15308, 16'd51356, 16'd50076, 16'd55887, 16'd9515, 16'd50416});
	test_expansion(128'h959fd0c4a12c14723bc82a1dfed13dd3, {16'd55874, 16'd53707, 16'd1043, 16'd3016, 16'd30667, 16'd40984, 16'd32227, 16'd58419, 16'd19629, 16'd14011, 16'd39001, 16'd44108, 16'd54247, 16'd1043, 16'd49887, 16'd64927, 16'd41596, 16'd12961, 16'd61527, 16'd43124, 16'd16445, 16'd37275, 16'd47141, 16'd19582, 16'd63328, 16'd6584});
	test_expansion(128'hbbfdeb2a4587e0528f409ae5ac7a1ebd, {16'd19641, 16'd30125, 16'd16218, 16'd46933, 16'd51556, 16'd13681, 16'd31904, 16'd20814, 16'd36439, 16'd24336, 16'd27426, 16'd11196, 16'd17700, 16'd61116, 16'd43715, 16'd3840, 16'd39101, 16'd8561, 16'd46352, 16'd16783, 16'd49356, 16'd4232, 16'd18112, 16'd33711, 16'd24811, 16'd3617});
	test_expansion(128'h2d913e8b16dc72f8d42f37be3775f1c9, {16'd52700, 16'd38998, 16'd60546, 16'd2920, 16'd16497, 16'd49312, 16'd61215, 16'd12217, 16'd23406, 16'd42470, 16'd56516, 16'd24907, 16'd57531, 16'd41465, 16'd47155, 16'd13437, 16'd37583, 16'd55892, 16'd58625, 16'd11746, 16'd40276, 16'd3455, 16'd6649, 16'd60707, 16'd29834, 16'd10161});
	test_expansion(128'h30d17a4330d408573ed65151d2dc1d22, {16'd40382, 16'd41476, 16'd64529, 16'd5188, 16'd46299, 16'd62877, 16'd22542, 16'd50488, 16'd49156, 16'd44199, 16'd11538, 16'd26587, 16'd14584, 16'd64771, 16'd36152, 16'd22903, 16'd19898, 16'd31192, 16'd45841, 16'd19537, 16'd43476, 16'd40325, 16'd27398, 16'd17593, 16'd20639, 16'd43501});
	test_expansion(128'h1b61d43b17e89968c3f841da583c883e, {16'd58264, 16'd10212, 16'd49780, 16'd10290, 16'd47713, 16'd19500, 16'd16845, 16'd4597, 16'd59420, 16'd37338, 16'd63387, 16'd23446, 16'd12885, 16'd1037, 16'd42701, 16'd3278, 16'd34634, 16'd41607, 16'd46140, 16'd8790, 16'd55972, 16'd60645, 16'd7063, 16'd19971, 16'd4630, 16'd50055});
	test_expansion(128'h799d68f9d03d2d3bdd9c8606c5c294af, {16'd48583, 16'd31770, 16'd1121, 16'd54506, 16'd11381, 16'd55603, 16'd1249, 16'd232, 16'd60428, 16'd3137, 16'd34092, 16'd34360, 16'd60551, 16'd21349, 16'd26161, 16'd26111, 16'd12341, 16'd14369, 16'd44099, 16'd19663, 16'd56642, 16'd42906, 16'd44269, 16'd5220, 16'd12964, 16'd34371});
	test_expansion(128'h5ee9244377d573c9270819829599e6a1, {16'd6870, 16'd32602, 16'd26608, 16'd55817, 16'd40848, 16'd59984, 16'd59822, 16'd44385, 16'd50737, 16'd38168, 16'd36199, 16'd42570, 16'd33660, 16'd6566, 16'd54034, 16'd44297, 16'd15072, 16'd25929, 16'd12844, 16'd60050, 16'd22972, 16'd2942, 16'd62413, 16'd41210, 16'd4953, 16'd47299});
	test_expansion(128'hc3f7033090b7b218cdeaf5da08a2bdf3, {16'd55700, 16'd37736, 16'd39640, 16'd2543, 16'd34756, 16'd29537, 16'd49421, 16'd3167, 16'd20860, 16'd40100, 16'd59628, 16'd42638, 16'd31919, 16'd12860, 16'd43203, 16'd30955, 16'd42731, 16'd8414, 16'd62752, 16'd60414, 16'd25837, 16'd17647, 16'd894, 16'd44680, 16'd50951, 16'd33389});
	test_expansion(128'he0d152383b0cebde51a56fadf65edc14, {16'd15758, 16'd64174, 16'd49561, 16'd15433, 16'd25912, 16'd45272, 16'd46604, 16'd60510, 16'd56575, 16'd38217, 16'd5955, 16'd9363, 16'd61362, 16'd29364, 16'd34311, 16'd24509, 16'd51997, 16'd59018, 16'd17598, 16'd14, 16'd54491, 16'd392, 16'd18077, 16'd45363, 16'd53201, 16'd16116});
	test_expansion(128'h6440fe8cdb69ffc3f0d8a2bee36a8e3e, {16'd40002, 16'd3027, 16'd25436, 16'd7640, 16'd15489, 16'd46174, 16'd51514, 16'd32365, 16'd21437, 16'd21365, 16'd25411, 16'd3518, 16'd37882, 16'd44133, 16'd23941, 16'd16389, 16'd11332, 16'd61817, 16'd5201, 16'd64364, 16'd33333, 16'd24404, 16'd193, 16'd41077, 16'd39796, 16'd3969});
	test_expansion(128'h8964e7afc4effb270a11d35fb74f1087, {16'd24774, 16'd38967, 16'd3261, 16'd40105, 16'd65324, 16'd62058, 16'd57088, 16'd58338, 16'd20033, 16'd59533, 16'd61839, 16'd3453, 16'd35957, 16'd14448, 16'd2648, 16'd40570, 16'd7101, 16'd34530, 16'd14911, 16'd53462, 16'd56462, 16'd56814, 16'd2564, 16'd57614, 16'd37519, 16'd32511});
	test_expansion(128'hfed87a1925ef0a9936536a736ddb3eab, {16'd50219, 16'd29736, 16'd56851, 16'd29989, 16'd56376, 16'd40970, 16'd39685, 16'd11753, 16'd7350, 16'd64619, 16'd8500, 16'd48224, 16'd920, 16'd24932, 16'd3537, 16'd50179, 16'd40148, 16'd50999, 16'd2258, 16'd18218, 16'd7986, 16'd58358, 16'd18203, 16'd27226, 16'd4526, 16'd8735});
	test_expansion(128'hf7d2a4e4a47c6647052930e27f286c35, {16'd51540, 16'd35487, 16'd57212, 16'd31607, 16'd15950, 16'd36123, 16'd5007, 16'd29621, 16'd63399, 16'd44686, 16'd59318, 16'd4832, 16'd42959, 16'd39793, 16'd60544, 16'd631, 16'd55052, 16'd29481, 16'd910, 16'd17753, 16'd54906, 16'd57692, 16'd4186, 16'd43007, 16'd25165, 16'd1803});
	test_expansion(128'h2f72eebce778484348a16e1400c8f887, {16'd12448, 16'd26402, 16'd24781, 16'd36985, 16'd15570, 16'd48808, 16'd8544, 16'd17264, 16'd56837, 16'd10806, 16'd34770, 16'd2760, 16'd46353, 16'd23958, 16'd21096, 16'd29056, 16'd31842, 16'd10289, 16'd61413, 16'd5714, 16'd2055, 16'd53582, 16'd45890, 16'd40565, 16'd9716, 16'd24832});
	test_expansion(128'h7a30597d0709dae36e234927c46650f6, {16'd4000, 16'd14216, 16'd5283, 16'd53452, 16'd9995, 16'd6116, 16'd49238, 16'd475, 16'd48385, 16'd47051, 16'd14343, 16'd10836, 16'd34678, 16'd4255, 16'd52638, 16'd7356, 16'd6912, 16'd62877, 16'd50272, 16'd23062, 16'd62736, 16'd37714, 16'd132, 16'd4937, 16'd20761, 16'd47378});
	test_expansion(128'h0769bac1dfc38b003f1badb9fc8c4164, {16'd23379, 16'd38527, 16'd7495, 16'd23179, 16'd15789, 16'd29236, 16'd58569, 16'd31542, 16'd43766, 16'd18076, 16'd58399, 16'd10057, 16'd26829, 16'd14152, 16'd57689, 16'd59234, 16'd41191, 16'd51744, 16'd61336, 16'd56433, 16'd42465, 16'd19749, 16'd57517, 16'd52419, 16'd60580, 16'd49887});
	test_expansion(128'h8ee2fbb8e9dd8fe35cd09959b68ab0a3, {16'd51919, 16'd33093, 16'd55538, 16'd42074, 16'd25801, 16'd25929, 16'd57984, 16'd25188, 16'd698, 16'd22795, 16'd11236, 16'd13340, 16'd23044, 16'd23476, 16'd28931, 16'd33953, 16'd53171, 16'd42130, 16'd47250, 16'd55696, 16'd9348, 16'd42391, 16'd23308, 16'd2968, 16'd34042, 16'd36351});
	test_expansion(128'h52341a3f3ad67cbe98d96ec215ca1fb4, {16'd33343, 16'd50066, 16'd4318, 16'd28469, 16'd64032, 16'd48014, 16'd13684, 16'd17926, 16'd28492, 16'd41678, 16'd15575, 16'd30488, 16'd30030, 16'd28853, 16'd12044, 16'd34042, 16'd58395, 16'd16036, 16'd36934, 16'd23151, 16'd59943, 16'd57223, 16'd57002, 16'd13042, 16'd46640, 16'd32477});
	test_expansion(128'h8ab661e762518ded7f44afcb10fa175d, {16'd22182, 16'd19820, 16'd38989, 16'd14993, 16'd57463, 16'd53070, 16'd40823, 16'd56342, 16'd6337, 16'd4322, 16'd20555, 16'd15158, 16'd35774, 16'd46336, 16'd17531, 16'd20546, 16'd20238, 16'd60106, 16'd3815, 16'd47331, 16'd41354, 16'd23622, 16'd36041, 16'd29971, 16'd65256, 16'd14031});
	test_expansion(128'ha04c30592b1a20d012b6eadfb7c1d5fd, {16'd35260, 16'd17814, 16'd24529, 16'd24127, 16'd3995, 16'd59056, 16'd27174, 16'd42875, 16'd11987, 16'd40137, 16'd24407, 16'd63238, 16'd59222, 16'd62697, 16'd37807, 16'd53770, 16'd27574, 16'd41044, 16'd20694, 16'd49527, 16'd122, 16'd63514, 16'd62681, 16'd59781, 16'd27888, 16'd62338});
	test_expansion(128'h5bba487286d43e09040becf7dc231256, {16'd44980, 16'd10336, 16'd47940, 16'd49456, 16'd36325, 16'd60251, 16'd3168, 16'd33278, 16'd33810, 16'd21754, 16'd55667, 16'd47424, 16'd9196, 16'd41838, 16'd32891, 16'd13927, 16'd22970, 16'd43209, 16'd63316, 16'd10012, 16'd51395, 16'd4771, 16'd1555, 16'd40684, 16'd58818, 16'd20695});
	test_expansion(128'h1a3d322e5738aecdbb419c176f4890f4, {16'd35310, 16'd22713, 16'd13234, 16'd7530, 16'd54540, 16'd19722, 16'd5153, 16'd28991, 16'd25046, 16'd36357, 16'd27456, 16'd53971, 16'd48703, 16'd3905, 16'd45977, 16'd37195, 16'd60065, 16'd11458, 16'd18765, 16'd7427, 16'd32723, 16'd22, 16'd36167, 16'd56155, 16'd20056, 16'd27851});
	test_expansion(128'h74055d72a2c6d5c8f21350ea9670c1fa, {16'd56625, 16'd7450, 16'd65268, 16'd5426, 16'd62280, 16'd10061, 16'd24843, 16'd52846, 16'd21297, 16'd45301, 16'd41531, 16'd62456, 16'd44936, 16'd280, 16'd59892, 16'd23492, 16'd45325, 16'd1091, 16'd26444, 16'd20950, 16'd17778, 16'd10301, 16'd40127, 16'd21894, 16'd38660, 16'd3612});
	test_expansion(128'hbaa229b8a27cc5eec5715473212221a8, {16'd29902, 16'd35856, 16'd63316, 16'd21087, 16'd61387, 16'd23596, 16'd31917, 16'd16209, 16'd49084, 16'd22451, 16'd38314, 16'd50256, 16'd19605, 16'd42028, 16'd16102, 16'd620, 16'd18096, 16'd25498, 16'd2443, 16'd20309, 16'd54291, 16'd16278, 16'd55432, 16'd46002, 16'd53319, 16'd61120});
	test_expansion(128'hfee67e1a1780826a6b61bb87ca21f06d, {16'd38100, 16'd27298, 16'd9801, 16'd32143, 16'd50629, 16'd7425, 16'd36977, 16'd32547, 16'd57490, 16'd48749, 16'd4533, 16'd15805, 16'd33996, 16'd26837, 16'd51090, 16'd3200, 16'd31300, 16'd50674, 16'd29675, 16'd25340, 16'd14615, 16'd56715, 16'd10263, 16'd51856, 16'd21982, 16'd29858});
	test_expansion(128'h180344a370aaa20ab4a737c4d462b9c7, {16'd8133, 16'd20534, 16'd26812, 16'd15834, 16'd27187, 16'd24805, 16'd62150, 16'd12205, 16'd33524, 16'd8493, 16'd42466, 16'd61445, 16'd45402, 16'd13279, 16'd3766, 16'd41885, 16'd11067, 16'd31039, 16'd12941, 16'd33191, 16'd60144, 16'd59652, 16'd12678, 16'd23341, 16'd34502, 16'd26107});
	test_expansion(128'h440d601095507e35aca70a0114ef1223, {16'd36070, 16'd51399, 16'd58361, 16'd48873, 16'd53792, 16'd50796, 16'd65420, 16'd48695, 16'd59693, 16'd26331, 16'd18441, 16'd62821, 16'd19700, 16'd41871, 16'd56586, 16'd40407, 16'd49591, 16'd32401, 16'd39902, 16'd5805, 16'd20166, 16'd59752, 16'd14592, 16'd51915, 16'd48034, 16'd64478});
	test_expansion(128'h7a2ccb314e323836ddef408eb3090248, {16'd65039, 16'd32675, 16'd29510, 16'd58564, 16'd47185, 16'd3718, 16'd60556, 16'd43705, 16'd14707, 16'd17118, 16'd18798, 16'd35705, 16'd21913, 16'd58283, 16'd37958, 16'd30156, 16'd3869, 16'd9369, 16'd55512, 16'd40415, 16'd19503, 16'd42285, 16'd48368, 16'd37863, 16'd44236, 16'd36351});
	test_expansion(128'hd0f1ad10a9444f0745c793fcc6b0cd74, {16'd44479, 16'd33103, 16'd50592, 16'd12743, 16'd26183, 16'd17949, 16'd51993, 16'd12306, 16'd50842, 16'd26249, 16'd1768, 16'd27146, 16'd59168, 16'd57883, 16'd21041, 16'd25264, 16'd5512, 16'd10333, 16'd28420, 16'd18929, 16'd2085, 16'd56811, 16'd1498, 16'd27257, 16'd42887, 16'd40479});
	test_expansion(128'hb5bee94904c46cf009b6e4fb6de58360, {16'd41658, 16'd15749, 16'd32194, 16'd58550, 16'd21618, 16'd31, 16'd54929, 16'd36730, 16'd35271, 16'd5463, 16'd61893, 16'd16631, 16'd34888, 16'd36708, 16'd41462, 16'd26267, 16'd13967, 16'd24505, 16'd9475, 16'd51170, 16'd22899, 16'd13780, 16'd64598, 16'd29460, 16'd22332, 16'd28072});
	test_expansion(128'h0b983bc13288b58d1c27cc665433bd6e, {16'd8985, 16'd53237, 16'd42883, 16'd40982, 16'd53980, 16'd44091, 16'd17633, 16'd8689, 16'd6599, 16'd24997, 16'd13888, 16'd33864, 16'd19570, 16'd27478, 16'd25034, 16'd56113, 16'd49280, 16'd587, 16'd56632, 16'd36819, 16'd23598, 16'd2275, 16'd52325, 16'd14015, 16'd44209, 16'd18676});
	test_expansion(128'hf4ac0f394e383c61d9770fbed9f2316a, {16'd45425, 16'd42065, 16'd54090, 16'd51855, 16'd9704, 16'd9674, 16'd51415, 16'd1678, 16'd42912, 16'd15250, 16'd61044, 16'd58975, 16'd11569, 16'd6532, 16'd37942, 16'd19736, 16'd52826, 16'd17778, 16'd62813, 16'd57937, 16'd43286, 16'd22888, 16'd61722, 16'd58047, 16'd12801, 16'd28990});
	test_expansion(128'h17fcc707ab7a9600bc0341eae099f096, {16'd52962, 16'd20843, 16'd40107, 16'd13758, 16'd58910, 16'd26742, 16'd61798, 16'd3473, 16'd594, 16'd2853, 16'd33388, 16'd30634, 16'd33211, 16'd11350, 16'd8855, 16'd23087, 16'd61994, 16'd22745, 16'd65042, 16'd4582, 16'd19949, 16'd3202, 16'd58698, 16'd50669, 16'd55662, 16'd57642});
	test_expansion(128'h5eae8f383257d3668964db4cd0f2b48c, {16'd7883, 16'd13816, 16'd27322, 16'd51975, 16'd21017, 16'd38028, 16'd47173, 16'd7722, 16'd14058, 16'd44411, 16'd19459, 16'd13907, 16'd60684, 16'd30526, 16'd59979, 16'd8813, 16'd39683, 16'd44952, 16'd30931, 16'd48494, 16'd51105, 16'd16465, 16'd28423, 16'd12506, 16'd64233, 16'd52358});
	test_expansion(128'hc1ed127afddca9abae2fe842c86e7720, {16'd8077, 16'd26192, 16'd46585, 16'd35997, 16'd9212, 16'd61551, 16'd48955, 16'd10039, 16'd28360, 16'd31970, 16'd51544, 16'd61846, 16'd54595, 16'd3671, 16'd34816, 16'd42893, 16'd46593, 16'd61724, 16'd9364, 16'd16738, 16'd18898, 16'd28962, 16'd53673, 16'd65304, 16'd53375, 16'd20396});
	test_expansion(128'hce9d7fa38b537caff9e105fe0e9df93c, {16'd31027, 16'd50855, 16'd56889, 16'd29727, 16'd26532, 16'd32813, 16'd51753, 16'd61400, 16'd10633, 16'd20693, 16'd53752, 16'd28140, 16'd47018, 16'd38933, 16'd24509, 16'd35630, 16'd26166, 16'd45233, 16'd53628, 16'd4442, 16'd26622, 16'd57475, 16'd50486, 16'd32870, 16'd62833, 16'd3712});
	test_expansion(128'h13eff89401ea16439612e076c177a181, {16'd54664, 16'd23367, 16'd3208, 16'd46859, 16'd44965, 16'd17403, 16'd46655, 16'd40055, 16'd7924, 16'd41610, 16'd31670, 16'd14468, 16'd9850, 16'd35115, 16'd21160, 16'd30400, 16'd64006, 16'd34514, 16'd55288, 16'd6034, 16'd21931, 16'd1616, 16'd20361, 16'd14560, 16'd7412, 16'd5012});
	test_expansion(128'hdd0b0f8f430b5bebdd222b68cda46b40, {16'd16470, 16'd20121, 16'd54901, 16'd35511, 16'd46550, 16'd15368, 16'd63785, 16'd9801, 16'd18815, 16'd30805, 16'd29772, 16'd8761, 16'd60563, 16'd9591, 16'd63348, 16'd18095, 16'd36589, 16'd30119, 16'd54300, 16'd58152, 16'd24260, 16'd41012, 16'd12881, 16'd35559, 16'd8564, 16'd11922});
	test_expansion(128'h35dbb679b46a607388cc876088869d8d, {16'd51301, 16'd52849, 16'd5516, 16'd50722, 16'd54205, 16'd25047, 16'd49687, 16'd57461, 16'd63735, 16'd52176, 16'd923, 16'd45725, 16'd11840, 16'd4578, 16'd49400, 16'd26814, 16'd13467, 16'd9745, 16'd4251, 16'd49461, 16'd2398, 16'd59479, 16'd24126, 16'd53649, 16'd16350, 16'd35643});
	test_expansion(128'h473e2ab3b4592e3f1c88cd6149139255, {16'd41853, 16'd3004, 16'd59153, 16'd14245, 16'd44090, 16'd41214, 16'd62081, 16'd65257, 16'd58662, 16'd60560, 16'd36698, 16'd29912, 16'd12959, 16'd21442, 16'd46323, 16'd16203, 16'd7759, 16'd35878, 16'd30675, 16'd9432, 16'd56940, 16'd28496, 16'd52511, 16'd57101, 16'd59575, 16'd16923});
	test_expansion(128'h755a4d024f8f1dcae0e05ab0985be138, {16'd33564, 16'd27606, 16'd8772, 16'd54957, 16'd11979, 16'd27462, 16'd17740, 16'd1400, 16'd47008, 16'd4455, 16'd49765, 16'd27469, 16'd26571, 16'd59694, 16'd49728, 16'd55768, 16'd41924, 16'd49527, 16'd33521, 16'd757, 16'd21742, 16'd31846, 16'd29870, 16'd20112, 16'd21719, 16'd6981});
	test_expansion(128'h9da415ff2d01bb88adb8bb18d036b5cb, {16'd4140, 16'd58501, 16'd63414, 16'd5300, 16'd27572, 16'd33301, 16'd32375, 16'd51442, 16'd38548, 16'd28056, 16'd40423, 16'd13884, 16'd52172, 16'd33699, 16'd56128, 16'd20801, 16'd25751, 16'd53515, 16'd8011, 16'd371, 16'd40149, 16'd16606, 16'd29584, 16'd57903, 16'd32136, 16'd18714});
	test_expansion(128'h766b036f15555047970a8624fdf720e4, {16'd51460, 16'd32856, 16'd26446, 16'd29136, 16'd43862, 16'd19349, 16'd21030, 16'd50855, 16'd25773, 16'd12729, 16'd37337, 16'd59667, 16'd18707, 16'd31003, 16'd46742, 16'd29533, 16'd4518, 16'd14683, 16'd4641, 16'd64212, 16'd36126, 16'd23522, 16'd56065, 16'd53464, 16'd61621, 16'd64155});
	test_expansion(128'hba9ef13451af6bd1292d32c31c17556f, {16'd1478, 16'd51878, 16'd2173, 16'd22692, 16'd29658, 16'd23849, 16'd43115, 16'd30155, 16'd8519, 16'd14872, 16'd19908, 16'd48489, 16'd53975, 16'd50236, 16'd39738, 16'd43646, 16'd7372, 16'd59488, 16'd58532, 16'd41662, 16'd49331, 16'd3116, 16'd37114, 16'd50879, 16'd51624, 16'd48093});
	test_expansion(128'h25c2d1933c7f1134ffe7c817d071883b, {16'd24525, 16'd21834, 16'd23411, 16'd43771, 16'd34625, 16'd45218, 16'd42782, 16'd60128, 16'd9401, 16'd38440, 16'd13866, 16'd19674, 16'd48522, 16'd15255, 16'd7433, 16'd26832, 16'd36240, 16'd45479, 16'd24595, 16'd10755, 16'd46012, 16'd55013, 16'd57984, 16'd40364, 16'd58186, 16'd49740});
	test_expansion(128'he95be8b5032c315eca4a0324963dc493, {16'd44987, 16'd13142, 16'd649, 16'd28857, 16'd58943, 16'd32054, 16'd53416, 16'd27714, 16'd6985, 16'd58067, 16'd28107, 16'd64250, 16'd17977, 16'd56063, 16'd37729, 16'd43114, 16'd30485, 16'd14902, 16'd24770, 16'd20026, 16'd37160, 16'd14915, 16'd32115, 16'd1599, 16'd21677, 16'd22169});
	test_expansion(128'hb6e5f2a5daeba4acf29ad2786401333e, {16'd31716, 16'd31062, 16'd54175, 16'd8057, 16'd60495, 16'd61318, 16'd47241, 16'd63440, 16'd15058, 16'd54623, 16'd21382, 16'd1372, 16'd52082, 16'd60007, 16'd48098, 16'd4822, 16'd29352, 16'd42033, 16'd47948, 16'd7298, 16'd20983, 16'd13783, 16'd19526, 16'd36467, 16'd5773, 16'd14972});
	test_expansion(128'hfb5848d54a1ff4d10978552afb0ae6f9, {16'd42433, 16'd55179, 16'd19212, 16'd18046, 16'd6793, 16'd32371, 16'd750, 16'd34087, 16'd30909, 16'd47754, 16'd3309, 16'd43680, 16'd1967, 16'd5584, 16'd51762, 16'd54522, 16'd41242, 16'd42196, 16'd60007, 16'd13125, 16'd3160, 16'd1644, 16'd32006, 16'd2961, 16'd35855, 16'd26478});
	test_expansion(128'h1a4af26eadf7d56ed3608eb7470a80cc, {16'd54941, 16'd51524, 16'd7496, 16'd47416, 16'd35098, 16'd10401, 16'd36448, 16'd27282, 16'd5805, 16'd25610, 16'd61557, 16'd31047, 16'd8897, 16'd28506, 16'd51516, 16'd33658, 16'd3658, 16'd42633, 16'd23519, 16'd32999, 16'd30391, 16'd36317, 16'd31981, 16'd17424, 16'd24332, 16'd42339});
	test_expansion(128'h6a60f7f052d17034ec74cc32e31071f4, {16'd28090, 16'd26932, 16'd24551, 16'd34889, 16'd32401, 16'd63972, 16'd2174, 16'd30467, 16'd40888, 16'd10505, 16'd43209, 16'd29072, 16'd63814, 16'd56593, 16'd42463, 16'd54904, 16'd40749, 16'd29728, 16'd47491, 16'd7943, 16'd38276, 16'd7257, 16'd54208, 16'd36030, 16'd7304, 16'd54182});
	test_expansion(128'hee140f64588483ee90dc97b82a5068e1, {16'd64536, 16'd62657, 16'd28974, 16'd15081, 16'd30490, 16'd60558, 16'd19479, 16'd40647, 16'd4427, 16'd58398, 16'd41041, 16'd14560, 16'd49323, 16'd23137, 16'd51482, 16'd48375, 16'd21242, 16'd8, 16'd15268, 16'd27470, 16'd64749, 16'd46836, 16'd33404, 16'd61374, 16'd15014, 16'd17340});
	test_expansion(128'h67c8638e30b70044380be558bfa926b1, {16'd58901, 16'd22422, 16'd18351, 16'd35919, 16'd12106, 16'd60492, 16'd28614, 16'd12616, 16'd41137, 16'd10382, 16'd1201, 16'd47148, 16'd37888, 16'd17627, 16'd18093, 16'd51256, 16'd45116, 16'd42298, 16'd63961, 16'd39861, 16'd42149, 16'd32916, 16'd54535, 16'd44364, 16'd45924, 16'd53425});
	test_expansion(128'hf2f954cfb51bdee186ba9e136b331cfb, {16'd2477, 16'd59535, 16'd14267, 16'd58605, 16'd49109, 16'd6793, 16'd30753, 16'd4710, 16'd37051, 16'd30271, 16'd1298, 16'd55815, 16'd9222, 16'd18462, 16'd17308, 16'd30953, 16'd36773, 16'd51058, 16'd36058, 16'd16591, 16'd43539, 16'd60857, 16'd32485, 16'd8296, 16'd33727, 16'd23738});
	test_expansion(128'h455c399e9ec90ae3e40eea78f9f5c304, {16'd24534, 16'd5723, 16'd45749, 16'd60688, 16'd60377, 16'd64215, 16'd44656, 16'd43266, 16'd6577, 16'd54612, 16'd31282, 16'd57091, 16'd37129, 16'd62230, 16'd60765, 16'd58153, 16'd40516, 16'd58113, 16'd41269, 16'd20687, 16'd25691, 16'd7840, 16'd30995, 16'd50226, 16'd12053, 16'd46887});
	test_expansion(128'hc5079fca831917d4613e9ec2fe70b346, {16'd49695, 16'd18357, 16'd14845, 16'd40470, 16'd29777, 16'd65344, 16'd61244, 16'd4026, 16'd20004, 16'd4067, 16'd13884, 16'd28616, 16'd10390, 16'd13984, 16'd42061, 16'd16419, 16'd42760, 16'd32218, 16'd2441, 16'd57302, 16'd47356, 16'd49340, 16'd3616, 16'd11644, 16'd20918, 16'd11454});
	test_expansion(128'h92acd20a6bc0a0230b9c875ce976f94e, {16'd51155, 16'd34596, 16'd8040, 16'd16737, 16'd63168, 16'd26340, 16'd26942, 16'd35033, 16'd14223, 16'd60956, 16'd13918, 16'd369, 16'd27819, 16'd37896, 16'd19368, 16'd51288, 16'd36386, 16'd17219, 16'd16156, 16'd50397, 16'd54168, 16'd33999, 16'd47862, 16'd58475, 16'd13842, 16'd2749});
	test_expansion(128'h47778ad01669e677b45d556800173b5f, {16'd51915, 16'd27135, 16'd6629, 16'd18323, 16'd8538, 16'd90, 16'd16461, 16'd2019, 16'd53447, 16'd58776, 16'd20574, 16'd57605, 16'd33661, 16'd13486, 16'd24795, 16'd10226, 16'd53608, 16'd10953, 16'd27143, 16'd57110, 16'd29393, 16'd9900, 16'd51448, 16'd38694, 16'd11806, 16'd5414});
	test_expansion(128'h09e7fa61f08aa0c0e1bab8e6dcb950d3, {16'd47382, 16'd43218, 16'd54748, 16'd60156, 16'd61627, 16'd53580, 16'd25529, 16'd8845, 16'd5594, 16'd26589, 16'd56177, 16'd33605, 16'd14373, 16'd26060, 16'd21932, 16'd41212, 16'd7412, 16'd888, 16'd44603, 16'd59086, 16'd49288, 16'd53954, 16'd41769, 16'd48084, 16'd27020, 16'd12503});
	test_expansion(128'hfdbb65d742d7e34071e4b7d1b595aaf5, {16'd38617, 16'd296, 16'd48343, 16'd47914, 16'd35505, 16'd30286, 16'd43118, 16'd21619, 16'd25320, 16'd55791, 16'd10340, 16'd50555, 16'd60650, 16'd6560, 16'd34843, 16'd63334, 16'd1901, 16'd59896, 16'd33707, 16'd11072, 16'd64820, 16'd56638, 16'd28748, 16'd12368, 16'd59623, 16'd24986});
	test_expansion(128'h52d739effd09fd2707ea9ab3d8692903, {16'd673, 16'd27455, 16'd47966, 16'd15667, 16'd20796, 16'd14733, 16'd36935, 16'd51711, 16'd49592, 16'd29592, 16'd37251, 16'd12582, 16'd33280, 16'd21917, 16'd11206, 16'd65035, 16'd1105, 16'd21098, 16'd32686, 16'd10543, 16'd65143, 16'd28970, 16'd22202, 16'd61656, 16'd26386, 16'd60508});
	test_expansion(128'h311e0ab3cdf1ad74bd7fa5df58aab07e, {16'd62129, 16'd13531, 16'd30649, 16'd20389, 16'd15880, 16'd16116, 16'd57619, 16'd45934, 16'd37612, 16'd39225, 16'd46001, 16'd27677, 16'd63324, 16'd48666, 16'd8679, 16'd59042, 16'd4004, 16'd64472, 16'd58041, 16'd41897, 16'd59460, 16'd65147, 16'd42132, 16'd51476, 16'd13957, 16'd25085});
	test_expansion(128'h0a8a715605a42a1fb02fdd8f7378d4f0, {16'd4077, 16'd17848, 16'd2383, 16'd33289, 16'd2977, 16'd43343, 16'd37101, 16'd7502, 16'd36021, 16'd25767, 16'd21360, 16'd51079, 16'd45980, 16'd15022, 16'd21241, 16'd15779, 16'd14008, 16'd57448, 16'd13191, 16'd61472, 16'd31307, 16'd36550, 16'd56114, 16'd39962, 16'd32593, 16'd55441});
	test_expansion(128'hec2c7bc2212e7ba7be087a4b7f905516, {16'd64005, 16'd15730, 16'd63086, 16'd6341, 16'd53792, 16'd49419, 16'd26488, 16'd28577, 16'd32749, 16'd35174, 16'd21286, 16'd13578, 16'd13833, 16'd13403, 16'd11190, 16'd1094, 16'd44261, 16'd15069, 16'd57928, 16'd47224, 16'd59474, 16'd4251, 16'd62455, 16'd22928, 16'd46371, 16'd15383});
	test_expansion(128'hf8c285ec7bb4c322e606258920a5e22a, {16'd51137, 16'd6893, 16'd38867, 16'd42067, 16'd3828, 16'd38129, 16'd57077, 16'd62329, 16'd12493, 16'd24966, 16'd10089, 16'd58604, 16'd29896, 16'd26836, 16'd59040, 16'd59134, 16'd40668, 16'd34313, 16'd24087, 16'd41966, 16'd22714, 16'd56985, 16'd2918, 16'd11591, 16'd19738, 16'd34701});
	test_expansion(128'h5a36bce8f2867a471c39971e5df3fa31, {16'd44247, 16'd5261, 16'd23957, 16'd24177, 16'd41546, 16'd33559, 16'd56784, 16'd10707, 16'd40453, 16'd38383, 16'd14503, 16'd49865, 16'd31085, 16'd9809, 16'd24671, 16'd59479, 16'd18091, 16'd62998, 16'd57526, 16'd39857, 16'd9441, 16'd59001, 16'd38608, 16'd43446, 16'd48331, 16'd62488});
	test_expansion(128'h04506f22859d94a1f06ae584937a5b6e, {16'd30122, 16'd35930, 16'd30006, 16'd55426, 16'd48147, 16'd54098, 16'd22922, 16'd30684, 16'd30746, 16'd31731, 16'd21915, 16'd9666, 16'd32394, 16'd35847, 16'd43493, 16'd41860, 16'd24269, 16'd22755, 16'd58126, 16'd48987, 16'd29179, 16'd33933, 16'd47099, 16'd16733, 16'd57243, 16'd52613});
	test_expansion(128'h59ec1eadfb2fb57993d78e5f592c76a6, {16'd22243, 16'd38216, 16'd50838, 16'd61450, 16'd1727, 16'd62132, 16'd31789, 16'd58161, 16'd12671, 16'd61147, 16'd17508, 16'd54839, 16'd50777, 16'd24124, 16'd22445, 16'd47015, 16'd60021, 16'd5541, 16'd27313, 16'd62427, 16'd34185, 16'd54333, 16'd30717, 16'd44008, 16'd61152, 16'd44308});
	test_expansion(128'h1a43e0b4942eb4cd2b4701cda42dd0b9, {16'd45587, 16'd31826, 16'd44018, 16'd4371, 16'd63459, 16'd61929, 16'd4777, 16'd9327, 16'd59424, 16'd63664, 16'd53854, 16'd64583, 16'd62871, 16'd36600, 16'd45412, 16'd25039, 16'd10309, 16'd46571, 16'd45901, 16'd24209, 16'd2607, 16'd23888, 16'd58678, 16'd14134, 16'd65144, 16'd1919});
	test_expansion(128'h01a3c1c6dd0cd39b49ffd067f5b25b33, {16'd26617, 16'd19239, 16'd5459, 16'd13727, 16'd31410, 16'd29092, 16'd31668, 16'd37567, 16'd7863, 16'd24515, 16'd59037, 16'd37979, 16'd4251, 16'd51273, 16'd45431, 16'd16401, 16'd26915, 16'd64182, 16'd3329, 16'd27386, 16'd16575, 16'd34428, 16'd23661, 16'd18339, 16'd44265, 16'd52783});
	test_expansion(128'h85ce4011edea4bc77640d67e52dda656, {16'd8990, 16'd26349, 16'd27529, 16'd45978, 16'd48210, 16'd27182, 16'd16549, 16'd55936, 16'd27335, 16'd49801, 16'd59974, 16'd56078, 16'd16089, 16'd51800, 16'd21646, 16'd28660, 16'd61132, 16'd49511, 16'd34572, 16'd7641, 16'd43374, 16'd64012, 16'd59928, 16'd63354, 16'd57174, 16'd45752});
	test_expansion(128'h3b6db6cfedc147252624eea0fef48180, {16'd27321, 16'd12194, 16'd23903, 16'd10966, 16'd13307, 16'd22282, 16'd64849, 16'd28641, 16'd22489, 16'd57100, 16'd33581, 16'd44299, 16'd32536, 16'd4960, 16'd3610, 16'd32318, 16'd19365, 16'd41637, 16'd29070, 16'd59685, 16'd21058, 16'd52584, 16'd42954, 16'd47879, 16'd16206, 16'd811});
	test_expansion(128'h5f5e1f008aeab9bfe38d6b89eb02af63, {16'd57500, 16'd23476, 16'd13732, 16'd38364, 16'd5175, 16'd17518, 16'd40410, 16'd11921, 16'd27303, 16'd58190, 16'd16464, 16'd60957, 16'd44592, 16'd9979, 16'd10322, 16'd56992, 16'd37051, 16'd17213, 16'd20881, 16'd40043, 16'd24557, 16'd51446, 16'd11619, 16'd25439, 16'd64712, 16'd29681});
	test_expansion(128'hff16fcddd86d4e034279cad19635f16e, {16'd29889, 16'd2201, 16'd16811, 16'd13465, 16'd46102, 16'd23525, 16'd49594, 16'd47641, 16'd24149, 16'd5625, 16'd10803, 16'd11472, 16'd1109, 16'd44004, 16'd52661, 16'd63770, 16'd62080, 16'd8514, 16'd60917, 16'd54760, 16'd38559, 16'd48367, 16'd36215, 16'd31027, 16'd24849, 16'd31932});
	test_expansion(128'h5de055b96f4f1f88aefc76e3e3f1ad41, {16'd56732, 16'd45298, 16'd64469, 16'd10211, 16'd15658, 16'd62218, 16'd58887, 16'd60743, 16'd34324, 16'd51452, 16'd42269, 16'd4234, 16'd38319, 16'd16136, 16'd13284, 16'd23103, 16'd46270, 16'd23627, 16'd16574, 16'd41819, 16'd61145, 16'd41178, 16'd25279, 16'd57013, 16'd20821, 16'd58894});
	test_expansion(128'hda686d5279bf209436b8eab44431902f, {16'd23729, 16'd50726, 16'd4163, 16'd51390, 16'd15131, 16'd3389, 16'd10211, 16'd64118, 16'd34939, 16'd32303, 16'd23605, 16'd58977, 16'd51283, 16'd31817, 16'd38751, 16'd21747, 16'd35906, 16'd49866, 16'd46807, 16'd60388, 16'd20406, 16'd36553, 16'd53229, 16'd21470, 16'd9224, 16'd61155});
	test_expansion(128'hdbe94ba8a4e63ebb8fa232168859db14, {16'd2447, 16'd5149, 16'd55231, 16'd58548, 16'd24861, 16'd62629, 16'd50250, 16'd2569, 16'd17380, 16'd53094, 16'd53507, 16'd2567, 16'd36010, 16'd64901, 16'd6443, 16'd35185, 16'd42577, 16'd8693, 16'd19669, 16'd20605, 16'd26143, 16'd20524, 16'd62612, 16'd30616, 16'd23673, 16'd17472});
	test_expansion(128'hebd865960b584e375c3ec1880e2d20b8, {16'd11218, 16'd32041, 16'd63295, 16'd2106, 16'd1904, 16'd32198, 16'd29002, 16'd9628, 16'd2587, 16'd3343, 16'd21637, 16'd11184, 16'd54330, 16'd7866, 16'd54350, 16'd7660, 16'd13721, 16'd21416, 16'd57198, 16'd52501, 16'd7143, 16'd42770, 16'd60000, 16'd55071, 16'd20241, 16'd39571});
	test_expansion(128'hca53d5e322bc1376718c245e662637b8, {16'd20151, 16'd45657, 16'd36369, 16'd53894, 16'd10431, 16'd34117, 16'd58231, 16'd47425, 16'd57355, 16'd15025, 16'd8205, 16'd46212, 16'd29282, 16'd2959, 16'd61168, 16'd57842, 16'd1805, 16'd40669, 16'd32440, 16'd51692, 16'd46004, 16'd63503, 16'd4213, 16'd62044, 16'd61477, 16'd45158});
	test_expansion(128'hadf68d5fa2961104344ffb54618a0490, {16'd39032, 16'd61023, 16'd55469, 16'd30292, 16'd57129, 16'd54590, 16'd21977, 16'd44651, 16'd55516, 16'd33852, 16'd36606, 16'd10932, 16'd33472, 16'd31209, 16'd40213, 16'd7748, 16'd40276, 16'd51909, 16'd51497, 16'd55798, 16'd65376, 16'd53258, 16'd56586, 16'd13404, 16'd23754, 16'd44631});
	test_expansion(128'h0f912504abd1510ef95faa8b35887f4d, {16'd20270, 16'd22883, 16'd542, 16'd26455, 16'd64480, 16'd52743, 16'd10662, 16'd57348, 16'd15555, 16'd5781, 16'd7371, 16'd54569, 16'd42833, 16'd15713, 16'd29261, 16'd53223, 16'd14294, 16'd48458, 16'd41008, 16'd56612, 16'd58343, 16'd22220, 16'd21167, 16'd44841, 16'd6507, 16'd60843});
	test_expansion(128'h7742cc993e80d713ec677417cec0775f, {16'd21103, 16'd50198, 16'd4018, 16'd31324, 16'd1776, 16'd19268, 16'd42047, 16'd55120, 16'd8128, 16'd2588, 16'd6340, 16'd35881, 16'd51596, 16'd1927, 16'd14374, 16'd6390, 16'd54340, 16'd2765, 16'd63439, 16'd41495, 16'd39851, 16'd43518, 16'd2521, 16'd43218, 16'd4726, 16'd42842});
	test_expansion(128'h6352a13c0a131fa276ab01cdb8321318, {16'd8149, 16'd59844, 16'd44189, 16'd2449, 16'd52619, 16'd18817, 16'd42242, 16'd10440, 16'd12992, 16'd10063, 16'd10424, 16'd20083, 16'd6542, 16'd53795, 16'd49342, 16'd29903, 16'd20823, 16'd29029, 16'd42850, 16'd59619, 16'd62885, 16'd7857, 16'd46789, 16'd56613, 16'd3086, 16'd2730});
	test_expansion(128'h8520fd36a38179bc044baacfa37bd66b, {16'd17901, 16'd53039, 16'd22380, 16'd16614, 16'd15902, 16'd14455, 16'd1505, 16'd26569, 16'd39349, 16'd27627, 16'd34913, 16'd52969, 16'd17951, 16'd33284, 16'd51168, 16'd61230, 16'd19642, 16'd34590, 16'd56992, 16'd52067, 16'd46713, 16'd25508, 16'd28117, 16'd7541, 16'd7399, 16'd33241});
	test_expansion(128'hfa475ec8e97efc0f75dcaaf8fc52b527, {16'd1415, 16'd46445, 16'd22807, 16'd11984, 16'd17806, 16'd30212, 16'd13016, 16'd57465, 16'd32363, 16'd32139, 16'd26471, 16'd10641, 16'd8482, 16'd55322, 16'd32444, 16'd48261, 16'd35677, 16'd46720, 16'd48218, 16'd52938, 16'd48611, 16'd53813, 16'd12409, 16'd33243, 16'd22584, 16'd52183});
	test_expansion(128'hf9e0e3d918b1f5040fb66748e938d324, {16'd4799, 16'd61837, 16'd62238, 16'd36520, 16'd51658, 16'd27212, 16'd52214, 16'd27112, 16'd8749, 16'd55026, 16'd36846, 16'd12100, 16'd51760, 16'd23598, 16'd36838, 16'd27971, 16'd17216, 16'd51032, 16'd16540, 16'd57623, 16'd18821, 16'd48281, 16'd60474, 16'd38867, 16'd35888, 16'd28600});
	test_expansion(128'h7979ebe74fff84a960269fbf8f0f4e37, {16'd62717, 16'd57427, 16'd5980, 16'd44107, 16'd26063, 16'd46979, 16'd1415, 16'd24757, 16'd14345, 16'd22018, 16'd48430, 16'd18901, 16'd42764, 16'd63027, 16'd32629, 16'd54230, 16'd45893, 16'd32289, 16'd62155, 16'd54229, 16'd23876, 16'd54963, 16'd6711, 16'd63452, 16'd7063, 16'd15055});
	test_expansion(128'h9a0d28d4d57dfa3bbf461cab91ae3339, {16'd42838, 16'd48935, 16'd57020, 16'd9067, 16'd5047, 16'd23775, 16'd56955, 16'd32062, 16'd59948, 16'd32424, 16'd46562, 16'd38332, 16'd3488, 16'd12589, 16'd3126, 16'd25216, 16'd57876, 16'd16802, 16'd26913, 16'd54471, 16'd46779, 16'd6376, 16'd28340, 16'd43631, 16'd58982, 16'd1440});
	test_expansion(128'h50e3e2e124247bf5dafabd21ca324f74, {16'd23054, 16'd32857, 16'd8442, 16'd16491, 16'd55619, 16'd13210, 16'd60308, 16'd5732, 16'd21079, 16'd49808, 16'd14698, 16'd16944, 16'd38417, 16'd55006, 16'd51536, 16'd41285, 16'd3589, 16'd10301, 16'd46952, 16'd2075, 16'd54297, 16'd14944, 16'd13516, 16'd6875, 16'd57659, 16'd23841});
	test_expansion(128'h88d63ea4d5cbcdcd844fdd1938535351, {16'd13084, 16'd48041, 16'd11594, 16'd24356, 16'd32602, 16'd18449, 16'd17688, 16'd35444, 16'd28726, 16'd32173, 16'd50562, 16'd10306, 16'd34060, 16'd53908, 16'd35777, 16'd15975, 16'd17381, 16'd42148, 16'd27340, 16'd55623, 16'd36852, 16'd60188, 16'd62826, 16'd64781, 16'd34650, 16'd28642});
	test_expansion(128'he98bc787d677c704c0e1dad7d4cb354c, {16'd32828, 16'd48188, 16'd50508, 16'd37020, 16'd32684, 16'd33255, 16'd59079, 16'd23891, 16'd63251, 16'd41244, 16'd56905, 16'd6549, 16'd2097, 16'd57781, 16'd10339, 16'd14993, 16'd29237, 16'd45808, 16'd41543, 16'd4139, 16'd36397, 16'd12595, 16'd52863, 16'd62187, 16'd21588, 16'd17817});
	test_expansion(128'he2277efc2159725a6b5905c89064f1dc, {16'd2586, 16'd39765, 16'd22573, 16'd29465, 16'd37006, 16'd32410, 16'd59825, 16'd65439, 16'd40669, 16'd34606, 16'd54264, 16'd13297, 16'd27162, 16'd61008, 16'd54987, 16'd5503, 16'd4535, 16'd34169, 16'd6326, 16'd40704, 16'd15933, 16'd46535, 16'd60351, 16'd53870, 16'd48118, 16'd6439});
	test_expansion(128'h46080d55caec812b63af3c29b9c6c885, {16'd14523, 16'd19042, 16'd1742, 16'd27472, 16'd44910, 16'd23874, 16'd55231, 16'd40858, 16'd12366, 16'd23910, 16'd15076, 16'd17722, 16'd22421, 16'd42250, 16'd14910, 16'd33009, 16'd30601, 16'd61101, 16'd44218, 16'd38121, 16'd16646, 16'd20313, 16'd43731, 16'd56246, 16'd45016, 16'd46442});
	test_expansion(128'h721fbb92a5654c54934a0e84a0f2a8db, {16'd34043, 16'd41018, 16'd10203, 16'd14409, 16'd3383, 16'd17853, 16'd65168, 16'd41101, 16'd57197, 16'd65487, 16'd37774, 16'd13780, 16'd55136, 16'd13036, 16'd5197, 16'd37439, 16'd31954, 16'd32667, 16'd58391, 16'd29465, 16'd55106, 16'd37712, 16'd30201, 16'd50914, 16'd18315, 16'd40112});
	test_expansion(128'h4bfcf9c13757a7dcaf695352b17358de, {16'd32507, 16'd37119, 16'd17798, 16'd58277, 16'd9754, 16'd61222, 16'd26427, 16'd39845, 16'd19826, 16'd48178, 16'd2837, 16'd29581, 16'd55554, 16'd23380, 16'd7744, 16'd62321, 16'd42554, 16'd18495, 16'd52729, 16'd13566, 16'd35187, 16'd35017, 16'd6967, 16'd59828, 16'd24719, 16'd63879});
	test_expansion(128'h927480804391c9aa834d1be6a5683186, {16'd62088, 16'd3945, 16'd28281, 16'd62273, 16'd50421, 16'd12920, 16'd21623, 16'd13446, 16'd51918, 16'd693, 16'd16519, 16'd13536, 16'd28502, 16'd1681, 16'd3801, 16'd18745, 16'd17110, 16'd24204, 16'd53640, 16'd8950, 16'd23136, 16'd19640, 16'd33353, 16'd62550, 16'd43603, 16'd4202});
	test_expansion(128'hdaaac9bdaa98730b57dbe04e321c65df, {16'd15211, 16'd24981, 16'd54170, 16'd49670, 16'd32504, 16'd27257, 16'd2881, 16'd30440, 16'd24325, 16'd1290, 16'd30133, 16'd6485, 16'd3994, 16'd56081, 16'd61462, 16'd56084, 16'd15177, 16'd5858, 16'd3668, 16'd9072, 16'd26028, 16'd56257, 16'd48955, 16'd49465, 16'd25675, 16'd17176});
	test_expansion(128'hbe7de47abe012a6b247462fe07bf113d, {16'd25476, 16'd56546, 16'd49474, 16'd18481, 16'd63877, 16'd48640, 16'd7860, 16'd12293, 16'd58715, 16'd53793, 16'd6703, 16'd13652, 16'd38978, 16'd57234, 16'd63140, 16'd46046, 16'd11442, 16'd38836, 16'd5657, 16'd8852, 16'd16835, 16'd10009, 16'd36299, 16'd17375, 16'd49804, 16'd56270});
	test_expansion(128'h5755da58b02fcc9d92a30a309534c2ee, {16'd7171, 16'd62113, 16'd38794, 16'd28140, 16'd28299, 16'd63240, 16'd7311, 16'd49761, 16'd7088, 16'd37750, 16'd9611, 16'd33756, 16'd40367, 16'd61547, 16'd9560, 16'd17064, 16'd42222, 16'd35633, 16'd49884, 16'd9884, 16'd27585, 16'd12714, 16'd36353, 16'd13677, 16'd55113, 16'd52566});
	test_expansion(128'h41b848c1a9d0de3250b104dc261c4ba8, {16'd59617, 16'd37459, 16'd56034, 16'd20009, 16'd47208, 16'd56523, 16'd50698, 16'd53688, 16'd386, 16'd14270, 16'd26278, 16'd18561, 16'd29713, 16'd58665, 16'd16985, 16'd2960, 16'd20333, 16'd54722, 16'd13324, 16'd60179, 16'd41888, 16'd41344, 16'd48465, 16'd10943, 16'd7142, 16'd32932});
	test_expansion(128'hb1d1d800aaa4adc485842ee59d2d226e, {16'd64952, 16'd17890, 16'd17153, 16'd63577, 16'd3757, 16'd29925, 16'd64599, 16'd54619, 16'd35350, 16'd18494, 16'd52118, 16'd186, 16'd44627, 16'd64618, 16'd14465, 16'd25503, 16'd33399, 16'd21570, 16'd10291, 16'd12659, 16'd6352, 16'd25279, 16'd3725, 16'd22498, 16'd57898, 16'd7376});
	test_expansion(128'h2f030eeb7ae12377269c2561be001daf, {16'd41925, 16'd12550, 16'd63542, 16'd32946, 16'd4641, 16'd32745, 16'd24767, 16'd10482, 16'd17332, 16'd18431, 16'd95, 16'd28589, 16'd19175, 16'd63023, 16'd31181, 16'd37735, 16'd7686, 16'd43777, 16'd16056, 16'd43771, 16'd45061, 16'd37372, 16'd29125, 16'd10774, 16'd29920, 16'd26395});
	test_expansion(128'hf059b8c16d9200c5e1e2d3b51abd2ec9, {16'd1139, 16'd51093, 16'd8513, 16'd11373, 16'd63979, 16'd37002, 16'd47580, 16'd64805, 16'd17979, 16'd59791, 16'd64586, 16'd11525, 16'd23126, 16'd40536, 16'd43512, 16'd2173, 16'd38886, 16'd13058, 16'd65091, 16'd31742, 16'd26242, 16'd62461, 16'd25328, 16'd21884, 16'd2864, 16'd36376});
	test_expansion(128'hfb6538ef2260cab208a981849336def5, {16'd4323, 16'd20047, 16'd65220, 16'd20812, 16'd4254, 16'd65237, 16'd9810, 16'd33800, 16'd23914, 16'd24735, 16'd55020, 16'd17492, 16'd15073, 16'd44447, 16'd7914, 16'd11315, 16'd46090, 16'd26991, 16'd5853, 16'd41672, 16'd30710, 16'd18652, 16'd15442, 16'd17223, 16'd22860, 16'd27642});
	test_expansion(128'h35c6fb4ba436eec3ca47e518871c51c6, {16'd54822, 16'd65064, 16'd41186, 16'd21304, 16'd55411, 16'd38350, 16'd52309, 16'd47860, 16'd38988, 16'd57285, 16'd29819, 16'd31499, 16'd65246, 16'd38148, 16'd63596, 16'd15004, 16'd7984, 16'd4389, 16'd46409, 16'd12849, 16'd18896, 16'd29536, 16'd56574, 16'd24349, 16'd7883, 16'd42});
	test_expansion(128'h2d8c828ac0e7b7421a68ec6b2cbdfbc2, {16'd12298, 16'd58359, 16'd17813, 16'd33087, 16'd42708, 16'd16059, 16'd41577, 16'd19735, 16'd40730, 16'd7195, 16'd16083, 16'd34859, 16'd1134, 16'd36558, 16'd33025, 16'd14375, 16'd2608, 16'd18314, 16'd27565, 16'd44898, 16'd20729, 16'd20896, 16'd24877, 16'd17834, 16'd47539, 16'd1945});
	test_expansion(128'ha4e89863857c14f0ec3ad06b95075127, {16'd2149, 16'd6909, 16'd60585, 16'd41929, 16'd6321, 16'd36037, 16'd55966, 16'd1235, 16'd33880, 16'd57397, 16'd12039, 16'd24197, 16'd6042, 16'd7201, 16'd1283, 16'd41508, 16'd5135, 16'd46062, 16'd6764, 16'd35777, 16'd26736, 16'd28943, 16'd46467, 16'd64014, 16'd56740, 16'd60135});
	test_expansion(128'he54f675790c21d1e82b4a74b42099237, {16'd44169, 16'd10105, 16'd50673, 16'd46432, 16'd24413, 16'd10642, 16'd60086, 16'd43904, 16'd38477, 16'd3956, 16'd57378, 16'd39970, 16'd50307, 16'd9139, 16'd48692, 16'd58626, 16'd63194, 16'd58524, 16'd6765, 16'd47111, 16'd51564, 16'd51251, 16'd60084, 16'd15542, 16'd24903, 16'd42305});
	test_expansion(128'hc4f827c6c16211ac53d46ebceeaf6656, {16'd16022, 16'd32590, 16'd38632, 16'd26897, 16'd1868, 16'd5992, 16'd366, 16'd17262, 16'd17152, 16'd20327, 16'd12324, 16'd23428, 16'd48777, 16'd40723, 16'd56084, 16'd22663, 16'd40252, 16'd14190, 16'd10795, 16'd33469, 16'd18447, 16'd8651, 16'd8892, 16'd34891, 16'd28549, 16'd33616});
	test_expansion(128'h9499f7f1eb487d9e842321c0b73ebe31, {16'd28859, 16'd29257, 16'd50827, 16'd64178, 16'd15453, 16'd39048, 16'd31337, 16'd22191, 16'd21146, 16'd54792, 16'd37151, 16'd8883, 16'd61843, 16'd7082, 16'd3393, 16'd10100, 16'd16828, 16'd15139, 16'd18311, 16'd8448, 16'd21093, 16'd50668, 16'd58615, 16'd37972, 16'd57090, 16'd5424});
	test_expansion(128'h5c147760e164e7b57ea6029b97b0bdb2, {16'd51118, 16'd44217, 16'd29179, 16'd30841, 16'd52378, 16'd63694, 16'd36606, 16'd47334, 16'd40687, 16'd22551, 16'd1306, 16'd52955, 16'd26421, 16'd29786, 16'd61745, 16'd27959, 16'd56399, 16'd52927, 16'd64395, 16'd19276, 16'd62585, 16'd26421, 16'd24170, 16'd18416, 16'd12375, 16'd18414});
	test_expansion(128'h786c485bba26140b0077d5207a9afb59, {16'd8444, 16'd49090, 16'd13933, 16'd59577, 16'd23533, 16'd14019, 16'd6540, 16'd60296, 16'd50021, 16'd49952, 16'd38805, 16'd37803, 16'd2313, 16'd29533, 16'd8496, 16'd36462, 16'd65405, 16'd56744, 16'd4567, 16'd15339, 16'd14942, 16'd6549, 16'd63468, 16'd19164, 16'd8936, 16'd16526});
	test_expansion(128'h1f6ad246d1b5bd3889b0e1f6469ae011, {16'd27055, 16'd59825, 16'd29802, 16'd11385, 16'd65427, 16'd8865, 16'd16310, 16'd5993, 16'd30661, 16'd33084, 16'd58581, 16'd9538, 16'd61837, 16'd13700, 16'd21274, 16'd44391, 16'd12565, 16'd6409, 16'd48858, 16'd39341, 16'd32864, 16'd59735, 16'd59355, 16'd3193, 16'd47915, 16'd4922});
	test_expansion(128'h72c596541674cd5d5700ff746c2de197, {16'd46470, 16'd22438, 16'd28254, 16'd13071, 16'd58456, 16'd25705, 16'd53263, 16'd24335, 16'd43301, 16'd60450, 16'd33015, 16'd21837, 16'd39620, 16'd50669, 16'd29783, 16'd35951, 16'd59543, 16'd1823, 16'd42058, 16'd35531, 16'd50958, 16'd49424, 16'd54428, 16'd8053, 16'd5640, 16'd29006});
	test_expansion(128'h8f61b5273ba38970da8bed380ad787a1, {16'd26182, 16'd24960, 16'd12630, 16'd3205, 16'd34767, 16'd1753, 16'd27568, 16'd12037, 16'd59351, 16'd27675, 16'd63873, 16'd65321, 16'd47076, 16'd53574, 16'd50166, 16'd7031, 16'd50635, 16'd32070, 16'd61424, 16'd10999, 16'd57265, 16'd19978, 16'd10057, 16'd35939, 16'd42171, 16'd30165});
	test_expansion(128'h1bfdbb9fafbcdc3fadf3da1935f9ccf1, {16'd7334, 16'd14563, 16'd34780, 16'd36902, 16'd43309, 16'd14330, 16'd51733, 16'd57671, 16'd1051, 16'd29917, 16'd41974, 16'd18814, 16'd49497, 16'd8328, 16'd41339, 16'd48636, 16'd51620, 16'd3839, 16'd32837, 16'd47226, 16'd52396, 16'd33078, 16'd23393, 16'd6666, 16'd61189, 16'd11263});
	test_expansion(128'hfd8e772e5436d640d669df12d9e10d99, {16'd36468, 16'd62954, 16'd14387, 16'd46232, 16'd27968, 16'd59276, 16'd20907, 16'd64518, 16'd13283, 16'd35385, 16'd40625, 16'd43372, 16'd41346, 16'd48359, 16'd62433, 16'd38414, 16'd30455, 16'd36393, 16'd46624, 16'd50885, 16'd2461, 16'd35246, 16'd65326, 16'd28248, 16'd64365, 16'd2663});
	test_expansion(128'h8ea1a4db4f2775e22dbf5c491f241923, {16'd3295, 16'd7975, 16'd54731, 16'd7407, 16'd58390, 16'd12143, 16'd11641, 16'd29037, 16'd1849, 16'd47188, 16'd58849, 16'd56151, 16'd50990, 16'd19915, 16'd22380, 16'd47434, 16'd17450, 16'd1660, 16'd44906, 16'd46226, 16'd34605, 16'd52079, 16'd11592, 16'd45433, 16'd34, 16'd53408});
	test_expansion(128'hf050a9aee8a41bf3961ebb03e577590f, {16'd30651, 16'd34675, 16'd20444, 16'd61231, 16'd19488, 16'd58959, 16'd61919, 16'd24951, 16'd5211, 16'd33390, 16'd33373, 16'd36934, 16'd36411, 16'd43350, 16'd26845, 16'd37900, 16'd34136, 16'd9980, 16'd40591, 16'd60959, 16'd56934, 16'd30043, 16'd36020, 16'd38551, 16'd41020, 16'd45408});
	test_expansion(128'h9732a0abf0946afe3ac9b28156e92743, {16'd8057, 16'd1048, 16'd36852, 16'd53476, 16'd19845, 16'd62411, 16'd28486, 16'd48955, 16'd41847, 16'd24253, 16'd36617, 16'd43221, 16'd50685, 16'd21025, 16'd10313, 16'd55867, 16'd39692, 16'd8425, 16'd58058, 16'd19154, 16'd14670, 16'd44078, 16'd47272, 16'd56734, 16'd35473, 16'd14680});
	test_expansion(128'h22148e63004bf40b396a29431e8ce2e1, {16'd23287, 16'd43047, 16'd65221, 16'd31183, 16'd62870, 16'd34339, 16'd30734, 16'd6406, 16'd8831, 16'd19260, 16'd8088, 16'd48227, 16'd57046, 16'd1069, 16'd14151, 16'd26739, 16'd31181, 16'd27559, 16'd34506, 16'd20879, 16'd46004, 16'd42688, 16'd18424, 16'd62334, 16'd14180, 16'd32464});
	test_expansion(128'h9036b26256eac6b111b3c5f72c8b6fff, {16'd48042, 16'd1357, 16'd29225, 16'd12751, 16'd35009, 16'd44347, 16'd16611, 16'd63267, 16'd8613, 16'd16897, 16'd23698, 16'd55588, 16'd10484, 16'd33710, 16'd1374, 16'd2117, 16'd56232, 16'd29927, 16'd61775, 16'd7195, 16'd9837, 16'd47214, 16'd28102, 16'd43076, 16'd22722, 16'd53679});
	test_expansion(128'hc9f1a07a6602c7ba7473d98d4cbe3353, {16'd65194, 16'd18870, 16'd5196, 16'd28368, 16'd2090, 16'd40191, 16'd12596, 16'd59413, 16'd53447, 16'd32216, 16'd50589, 16'd48166, 16'd59549, 16'd19402, 16'd36048, 16'd54964, 16'd63410, 16'd64058, 16'd59338, 16'd14618, 16'd40785, 16'd36116, 16'd22020, 16'd40692, 16'd50421, 16'd1420});
	test_expansion(128'h2a4ac4df245738ce9c28a1379c8d0357, {16'd47565, 16'd31949, 16'd20291, 16'd6924, 16'd47476, 16'd60625, 16'd62008, 16'd34433, 16'd40771, 16'd62419, 16'd43896, 16'd14743, 16'd42438, 16'd53666, 16'd40078, 16'd40320, 16'd55938, 16'd49272, 16'd55522, 16'd49954, 16'd58802, 16'd44135, 16'd39654, 16'd21805, 16'd28884, 16'd58401});
	test_expansion(128'h87b1340a4f93aff50f784a31a23c2213, {16'd4783, 16'd18356, 16'd61072, 16'd61238, 16'd62196, 16'd11071, 16'd64997, 16'd57125, 16'd61879, 16'd49729, 16'd32519, 16'd8618, 16'd8285, 16'd20312, 16'd56566, 16'd3261, 16'd1242, 16'd14884, 16'd500, 16'd51939, 16'd50798, 16'd64458, 16'd9901, 16'd56910, 16'd12611, 16'd21544});
	test_expansion(128'hb24ee3c9cdb52e51cad41a42193ab361, {16'd45164, 16'd44725, 16'd29913, 16'd6699, 16'd3222, 16'd61789, 16'd23445, 16'd52833, 16'd35196, 16'd562, 16'd15128, 16'd7614, 16'd56759, 16'd369, 16'd10985, 16'd17758, 16'd16420, 16'd8573, 16'd10451, 16'd35792, 16'd40948, 16'd306, 16'd10355, 16'd13800, 16'd57897, 16'd59048});
	test_expansion(128'h7eb36b002e118cad959448fef6bb9661, {16'd18592, 16'd30252, 16'd62446, 16'd48969, 16'd41155, 16'd5918, 16'd7630, 16'd5856, 16'd7429, 16'd63290, 16'd4736, 16'd14860, 16'd49314, 16'd36968, 16'd44826, 16'd9014, 16'd65105, 16'd16558, 16'd38167, 16'd62620, 16'd6900, 16'd34647, 16'd61931, 16'd1113, 16'd54269, 16'd28608});
	test_expansion(128'h44478361da0cdf4cae9dcaf3915d092a, {16'd51747, 16'd61486, 16'd33676, 16'd18736, 16'd1745, 16'd3370, 16'd60911, 16'd50224, 16'd18457, 16'd27574, 16'd56337, 16'd40010, 16'd59303, 16'd54049, 16'd8687, 16'd36964, 16'd7185, 16'd51782, 16'd24687, 16'd7568, 16'd57504, 16'd63118, 16'd548, 16'd37097, 16'd65305, 16'd38766});
	test_expansion(128'h3631b97fd2ad497a6296f30e3994db5f, {16'd25642, 16'd936, 16'd15724, 16'd60210, 16'd55402, 16'd36874, 16'd50398, 16'd9774, 16'd2682, 16'd55700, 16'd21078, 16'd65136, 16'd172, 16'd56033, 16'd53942, 16'd59024, 16'd45751, 16'd23247, 16'd1289, 16'd40542, 16'd17974, 16'd52809, 16'd47212, 16'd38873, 16'd31294, 16'd9262});
	test_expansion(128'hbd4c6d915b4e10122e022cbb8ff0ccb2, {16'd18551, 16'd1476, 16'd42913, 16'd10886, 16'd33504, 16'd30009, 16'd50602, 16'd4195, 16'd45173, 16'd890, 16'd44184, 16'd53083, 16'd4512, 16'd39096, 16'd16703, 16'd36454, 16'd41769, 16'd32010, 16'd25280, 16'd9523, 16'd15150, 16'd27702, 16'd41783, 16'd18280, 16'd54741, 16'd41366});
	test_expansion(128'h818475da52f2aa7d4f42bb95139fefb5, {16'd31177, 16'd39649, 16'd64702, 16'd26757, 16'd24855, 16'd49954, 16'd7603, 16'd6109, 16'd35569, 16'd25883, 16'd25930, 16'd31228, 16'd4768, 16'd23306, 16'd63711, 16'd27979, 16'd30828, 16'd21023, 16'd49257, 16'd3714, 16'd28320, 16'd25376, 16'd51411, 16'd43221, 16'd56952, 16'd45057});
	test_expansion(128'h170217d7a85f2ff3d10e7fb238305108, {16'd33633, 16'd29811, 16'd44338, 16'd39166, 16'd54659, 16'd16129, 16'd40291, 16'd11203, 16'd29771, 16'd20416, 16'd58802, 16'd43671, 16'd43117, 16'd32197, 16'd8603, 16'd54396, 16'd17734, 16'd29003, 16'd51299, 16'd30838, 16'd29514, 16'd27101, 16'd64673, 16'd53207, 16'd64967, 16'd14409});
	test_expansion(128'h02c57c65dd07b45969f355b8ecf628e8, {16'd41074, 16'd20613, 16'd29770, 16'd33291, 16'd9575, 16'd62920, 16'd43685, 16'd56041, 16'd9387, 16'd6586, 16'd33167, 16'd6900, 16'd44930, 16'd19986, 16'd64627, 16'd54155, 16'd8706, 16'd43294, 16'd18621, 16'd19433, 16'd6419, 16'd27764, 16'd57696, 16'd46726, 16'd15648, 16'd55283});
	test_expansion(128'h656de40e9d221a4b2862b8edae501891, {16'd44421, 16'd61014, 16'd55648, 16'd33173, 16'd42415, 16'd59637, 16'd61652, 16'd1432, 16'd32097, 16'd65086, 16'd60598, 16'd14125, 16'd12545, 16'd64933, 16'd57980, 16'd50917, 16'd41396, 16'd39589, 16'd8409, 16'd41527, 16'd57294, 16'd6812, 16'd49130, 16'd3683, 16'd7219, 16'd4926});
	test_expansion(128'hda34f1ad92a0cc414d0ee571e3c1b1a7, {16'd57799, 16'd57510, 16'd7565, 16'd24254, 16'd1851, 16'd54375, 16'd60307, 16'd37767, 16'd27360, 16'd58999, 16'd65215, 16'd56886, 16'd52332, 16'd58773, 16'd10481, 16'd27801, 16'd115, 16'd58084, 16'd12400, 16'd9705, 16'd1538, 16'd41343, 16'd1556, 16'd51025, 16'd44941, 16'd27408});
	test_expansion(128'hefe2342476cbef735602d37f9103ad5f, {16'd641, 16'd47688, 16'd12952, 16'd57299, 16'd22156, 16'd4582, 16'd60676, 16'd9363, 16'd8718, 16'd63833, 16'd57650, 16'd9850, 16'd52235, 16'd61184, 16'd12404, 16'd13005, 16'd43130, 16'd15975, 16'd45789, 16'd16279, 16'd37445, 16'd16120, 16'd64851, 16'd7376, 16'd11026, 16'd356});
	test_expansion(128'hbdee627c502a62256c2fe1f7942fb1ad, {16'd22248, 16'd14616, 16'd42944, 16'd36344, 16'd56749, 16'd419, 16'd34213, 16'd57355, 16'd18577, 16'd9584, 16'd41646, 16'd45767, 16'd55966, 16'd20093, 16'd54823, 16'd25823, 16'd25304, 16'd17120, 16'd34424, 16'd12561, 16'd39140, 16'd24998, 16'd45074, 16'd55503, 16'd40083, 16'd51500});
	test_expansion(128'h223084d3ef4cd0aecee69a2815475052, {16'd48147, 16'd48396, 16'd27696, 16'd23336, 16'd36778, 16'd26780, 16'd49130, 16'd25202, 16'd18974, 16'd33186, 16'd11358, 16'd46518, 16'd49944, 16'd49341, 16'd40423, 16'd63724, 16'd24744, 16'd61723, 16'd54606, 16'd63808, 16'd47836, 16'd48326, 16'd51452, 16'd30575, 16'd60083, 16'd39012});
	test_expansion(128'hd6ebe0130790db77de29ef13494d19f3, {16'd31786, 16'd35572, 16'd36762, 16'd9219, 16'd49205, 16'd34165, 16'd53594, 16'd16224, 16'd15098, 16'd54459, 16'd42891, 16'd5734, 16'd914, 16'd45130, 16'd47353, 16'd51257, 16'd57642, 16'd53006, 16'd45989, 16'd2789, 16'd15881, 16'd14211, 16'd55085, 16'd40051, 16'd40176, 16'd21217});
	test_expansion(128'h46f3dbcc443a8ca42fce7e1da70ddd4f, {16'd24169, 16'd53088, 16'd27404, 16'd1591, 16'd4658, 16'd10193, 16'd39430, 16'd55054, 16'd61050, 16'd63296, 16'd60959, 16'd18531, 16'd22117, 16'd38483, 16'd65350, 16'd32841, 16'd49103, 16'd54700, 16'd8216, 16'd62640, 16'd60167, 16'd27985, 16'd57950, 16'd51179, 16'd42748, 16'd19161});
	test_expansion(128'h5acb8d60a251beb4e726f176eb5376f0, {16'd53876, 16'd29164, 16'd33143, 16'd31616, 16'd27242, 16'd14806, 16'd34704, 16'd49580, 16'd17329, 16'd62107, 16'd47749, 16'd64770, 16'd60181, 16'd17673, 16'd57931, 16'd56616, 16'd24501, 16'd31270, 16'd15974, 16'd64698, 16'd24706, 16'd41436, 16'd62549, 16'd64551, 16'd65024, 16'd44296});
	test_expansion(128'h6977e9754a49f5b27d2d59c14826fad9, {16'd50544, 16'd62160, 16'd63866, 16'd55941, 16'd11613, 16'd24855, 16'd56297, 16'd16868, 16'd56554, 16'd51744, 16'd11549, 16'd17751, 16'd8805, 16'd10049, 16'd12064, 16'd34303, 16'd55230, 16'd24794, 16'd13171, 16'd15275, 16'd18731, 16'd47572, 16'd46470, 16'd47282, 16'd28997, 16'd8396});
	test_expansion(128'hfe7f65b0a92657ceed05fceeddf2b2d3, {16'd6007, 16'd19645, 16'd47002, 16'd57679, 16'd14618, 16'd25157, 16'd18725, 16'd41102, 16'd59478, 16'd17226, 16'd14288, 16'd48047, 16'd4468, 16'd52621, 16'd31457, 16'd35106, 16'd61893, 16'd20279, 16'd12819, 16'd65213, 16'd22827, 16'd47253, 16'd27835, 16'd65005, 16'd3448, 16'd2150});
	test_expansion(128'hf524becd2d6e6c09c0818a6fcef44920, {16'd5375, 16'd28465, 16'd20402, 16'd216, 16'd51368, 16'd48476, 16'd64677, 16'd8699, 16'd25348, 16'd23589, 16'd7345, 16'd38893, 16'd41797, 16'd44345, 16'd23010, 16'd54450, 16'd50290, 16'd41781, 16'd7453, 16'd55057, 16'd38208, 16'd23254, 16'd57653, 16'd6869, 16'd22452, 16'd12588});
	test_expansion(128'h38abe6758e591634ee062f0f5736faa6, {16'd36176, 16'd11379, 16'd1640, 16'd56632, 16'd14525, 16'd42857, 16'd57925, 16'd14515, 16'd41988, 16'd22417, 16'd26581, 16'd47415, 16'd39291, 16'd58135, 16'd50128, 16'd50814, 16'd31078, 16'd5185, 16'd6186, 16'd39516, 16'd51454, 16'd424, 16'd62276, 16'd6468, 16'd60908, 16'd54613});
	test_expansion(128'h31bea255cee8399b155273ecd11027d3, {16'd8281, 16'd44539, 16'd15396, 16'd29606, 16'd58515, 16'd19876, 16'd56799, 16'd40086, 16'd9778, 16'd56846, 16'd21207, 16'd17760, 16'd57866, 16'd7871, 16'd32890, 16'd59382, 16'd50249, 16'd441, 16'd25362, 16'd50491, 16'd22492, 16'd55202, 16'd11585, 16'd49496, 16'd63633, 16'd18605});
	test_expansion(128'h96b01fa9143da9c34a1e021d5306ade1, {16'd30153, 16'd10473, 16'd37077, 16'd22116, 16'd50933, 16'd1635, 16'd45836, 16'd30404, 16'd58196, 16'd9560, 16'd51849, 16'd61954, 16'd32265, 16'd7459, 16'd9684, 16'd57811, 16'd8958, 16'd19703, 16'd65151, 16'd45694, 16'd22172, 16'd59157, 16'd52903, 16'd36551, 16'd30431, 16'd22471});
	test_expansion(128'hecbdb52f4fd3d4004e3c32f8db21f2ec, {16'd9438, 16'd49924, 16'd36734, 16'd3847, 16'd40530, 16'd21743, 16'd44974, 16'd17745, 16'd8912, 16'd41551, 16'd13500, 16'd28554, 16'd60150, 16'd55939, 16'd15634, 16'd35752, 16'd17042, 16'd16185, 16'd43364, 16'd33607, 16'd27382, 16'd11758, 16'd43590, 16'd45420, 16'd11081, 16'd39606});
	test_expansion(128'ha9c84d90673a00a252b7f9bcd047a8a5, {16'd32464, 16'd35822, 16'd6011, 16'd24703, 16'd3394, 16'd58060, 16'd47650, 16'd60617, 16'd40586, 16'd52646, 16'd21554, 16'd22401, 16'd40982, 16'd14687, 16'd37561, 16'd65001, 16'd39229, 16'd18895, 16'd60662, 16'd24177, 16'd60759, 16'd26694, 16'd50168, 16'd35077, 16'd26552, 16'd36152});
	test_expansion(128'h36f1b32ef0c8e74197008f642ff57131, {16'd17062, 16'd54913, 16'd54371, 16'd56506, 16'd59944, 16'd31695, 16'd42430, 16'd1239, 16'd40068, 16'd58249, 16'd55890, 16'd29526, 16'd65497, 16'd1095, 16'd49395, 16'd54318, 16'd33844, 16'd53389, 16'd63520, 16'd34441, 16'd41852, 16'd25309, 16'd13347, 16'd54512, 16'd51969, 16'd1725});
	test_expansion(128'h9739b8db60a7bb4ee60ab1911c7602df, {16'd22065, 16'd24497, 16'd12353, 16'd6413, 16'd3503, 16'd20382, 16'd61208, 16'd46821, 16'd64377, 16'd43476, 16'd46910, 16'd37333, 16'd17453, 16'd63237, 16'd48234, 16'd34930, 16'd54698, 16'd23596, 16'd35730, 16'd41668, 16'd60898, 16'd17086, 16'd419, 16'd47936, 16'd53558, 16'd1768});
	test_expansion(128'hef46718bb4e26cfb7a93034ba53d0eee, {16'd43474, 16'd47386, 16'd37311, 16'd37533, 16'd59465, 16'd20035, 16'd40246, 16'd14804, 16'd49819, 16'd47148, 16'd63976, 16'd21169, 16'd39587, 16'd16780, 16'd6753, 16'd43182, 16'd5353, 16'd61680, 16'd64989, 16'd39929, 16'd24724, 16'd29685, 16'd33468, 16'd59788, 16'd5241, 16'd28362});
	test_expansion(128'h5b1e37e66e1541ccc78c91cd0fbb8534, {16'd18274, 16'd42139, 16'd24427, 16'd26656, 16'd23607, 16'd51083, 16'd17441, 16'd36533, 16'd56813, 16'd53946, 16'd51815, 16'd55834, 16'd362, 16'd10407, 16'd58646, 16'd455, 16'd36135, 16'd5316, 16'd8337, 16'd46269, 16'd52870, 16'd23635, 16'd35838, 16'd27700, 16'd10219, 16'd54225});
	test_expansion(128'he132b40383455901b55088afa6094247, {16'd37244, 16'd35119, 16'd234, 16'd16493, 16'd8889, 16'd18015, 16'd32481, 16'd55207, 16'd17394, 16'd54686, 16'd35879, 16'd1423, 16'd52066, 16'd56277, 16'd25470, 16'd9510, 16'd11960, 16'd56536, 16'd32241, 16'd14185, 16'd31443, 16'd1685, 16'd141, 16'd49522, 16'd50353, 16'd58302});
	test_expansion(128'hf8f1fb49d42897e1e2f9d7ff2b1e91bb, {16'd11819, 16'd17819, 16'd44173, 16'd10947, 16'd24270, 16'd54355, 16'd62843, 16'd36213, 16'd11957, 16'd25059, 16'd3676, 16'd37497, 16'd21110, 16'd6035, 16'd58508, 16'd38691, 16'd9548, 16'd61077, 16'd11678, 16'd5075, 16'd58792, 16'd41535, 16'd12764, 16'd15589, 16'd59205, 16'd40815});
	test_expansion(128'hc8c85fee3b0636e1cda1289be32d7d37, {16'd27383, 16'd3699, 16'd8053, 16'd11124, 16'd54635, 16'd38422, 16'd61320, 16'd9317, 16'd38228, 16'd24017, 16'd61957, 16'd32489, 16'd62515, 16'd33403, 16'd30893, 16'd57842, 16'd14781, 16'd32838, 16'd60954, 16'd2950, 16'd15896, 16'd9818, 16'd64708, 16'd42779, 16'd64466, 16'd38142});
	test_expansion(128'h23498db0cc23d1501e60f8fb1b7b3e51, {16'd30802, 16'd26824, 16'd45749, 16'd48979, 16'd56768, 16'd23722, 16'd39473, 16'd23251, 16'd32728, 16'd7724, 16'd2879, 16'd47048, 16'd15197, 16'd22645, 16'd35851, 16'd15615, 16'd18095, 16'd4126, 16'd43703, 16'd29479, 16'd51801, 16'd18899, 16'd44470, 16'd15105, 16'd13792, 16'd3409});
	test_expansion(128'h718ace072efc116f841839c29cb2ff18, {16'd64665, 16'd59272, 16'd49742, 16'd31322, 16'd48654, 16'd9704, 16'd28281, 16'd29111, 16'd10294, 16'd62630, 16'd57426, 16'd52986, 16'd31896, 16'd43128, 16'd9853, 16'd61209, 16'd38502, 16'd8018, 16'd30455, 16'd3361, 16'd47072, 16'd56833, 16'd27476, 16'd30465, 16'd22244, 16'd54492});
	test_expansion(128'h0a5444c7f307a9affe1fd6b1122cc14c, {16'd27150, 16'd41889, 16'd33378, 16'd43216, 16'd45018, 16'd64935, 16'd64328, 16'd28719, 16'd16948, 16'd12558, 16'd53940, 16'd634, 16'd51981, 16'd38521, 16'd58309, 16'd36284, 16'd4555, 16'd19502, 16'd46225, 16'd44515, 16'd25055, 16'd64239, 16'd30138, 16'd39813, 16'd11066, 16'd37010});
	test_expansion(128'hbc053656fa6979d8ef6d0db600821d7a, {16'd61300, 16'd44002, 16'd50438, 16'd62172, 16'd36246, 16'd1329, 16'd56491, 16'd37515, 16'd14235, 16'd4878, 16'd10363, 16'd36303, 16'd48177, 16'd22706, 16'd9547, 16'd61258, 16'd48418, 16'd53385, 16'd12318, 16'd25241, 16'd36373, 16'd28443, 16'd18558, 16'd29144, 16'd61987, 16'd60742});
	test_expansion(128'h6bd27eee52dc169575ef2e9a2d32be53, {16'd60197, 16'd53929, 16'd32092, 16'd23981, 16'd55629, 16'd55321, 16'd56626, 16'd57249, 16'd47080, 16'd52325, 16'd38223, 16'd51143, 16'd33431, 16'd62042, 16'd38741, 16'd27387, 16'd12371, 16'd62728, 16'd61582, 16'd4961, 16'd20074, 16'd30996, 16'd17290, 16'd36079, 16'd33396, 16'd51712});
	test_expansion(128'hab07a15dd83e14a49d78d1d524c0dcf1, {16'd7315, 16'd54718, 16'd12493, 16'd20574, 16'd1947, 16'd57708, 16'd48197, 16'd35543, 16'd44945, 16'd12198, 16'd6584, 16'd41498, 16'd28510, 16'd44565, 16'd5051, 16'd18758, 16'd21324, 16'd18162, 16'd44784, 16'd27670, 16'd7589, 16'd28368, 16'd8296, 16'd51380, 16'd60106, 16'd8964});
	test_expansion(128'h2cd63a876585e7b0b0f64cabcaa180f5, {16'd55776, 16'd59840, 16'd41830, 16'd28289, 16'd6952, 16'd20404, 16'd23881, 16'd60546, 16'd50892, 16'd10742, 16'd3765, 16'd2267, 16'd46628, 16'd64319, 16'd16472, 16'd39270, 16'd60676, 16'd19911, 16'd39586, 16'd8141, 16'd60311, 16'd45564, 16'd2217, 16'd63792, 16'd63763, 16'd47039});
	test_expansion(128'h5a4bd08ca19fb705735d25a7a734723e, {16'd31539, 16'd58231, 16'd31746, 16'd30930, 16'd26994, 16'd14003, 16'd31301, 16'd50665, 16'd1320, 16'd56324, 16'd39503, 16'd42297, 16'd25705, 16'd35700, 16'd30553, 16'd21776, 16'd14774, 16'd2384, 16'd35971, 16'd56953, 16'd25008, 16'd31898, 16'd22978, 16'd11960, 16'd26485, 16'd25379});
	test_expansion(128'h7a702a808a5a3b6adc8708fc5a85755b, {16'd8100, 16'd23239, 16'd48548, 16'd49461, 16'd35461, 16'd19946, 16'd40194, 16'd19789, 16'd38549, 16'd46741, 16'd63826, 16'd57486, 16'd20695, 16'd37387, 16'd33977, 16'd39276, 16'd63236, 16'd32260, 16'd33375, 16'd29323, 16'd29969, 16'd54795, 16'd30247, 16'd65349, 16'd62364, 16'd47027});
	test_expansion(128'h1c59db483e0e2a4dfefe91ccd53c5222, {16'd49830, 16'd22623, 16'd5777, 16'd33752, 16'd51087, 16'd63767, 16'd55949, 16'd53462, 16'd40842, 16'd24308, 16'd44271, 16'd29506, 16'd30724, 16'd32732, 16'd16052, 16'd60273, 16'd63385, 16'd51492, 16'd58276, 16'd37482, 16'd54151, 16'd32159, 16'd19120, 16'd34876, 16'd25511, 16'd4881});
	test_expansion(128'h879d0a9418b2bee7a7aa68d7f3730a14, {16'd61903, 16'd53688, 16'd49013, 16'd6084, 16'd29695, 16'd33618, 16'd34312, 16'd1257, 16'd10853, 16'd5876, 16'd23155, 16'd45656, 16'd25673, 16'd10543, 16'd3163, 16'd63871, 16'd9221, 16'd52905, 16'd52166, 16'd3636, 16'd14635, 16'd29175, 16'd35067, 16'd34566, 16'd56484, 16'd19116});
	test_expansion(128'hfceae3623bbc2f6a3bbb57b30b94ef9d, {16'd55803, 16'd46714, 16'd17124, 16'd61975, 16'd31658, 16'd40391, 16'd29071, 16'd46034, 16'd7399, 16'd57069, 16'd26399, 16'd32286, 16'd35879, 16'd49827, 16'd45631, 16'd29516, 16'd25, 16'd30708, 16'd20878, 16'd47059, 16'd30772, 16'd887, 16'd4341, 16'd64514, 16'd21257, 16'd6002});
	test_expansion(128'he04e08c573ada0da0eb5a79a5db01af0, {16'd61637, 16'd58423, 16'd48080, 16'd64420, 16'd15985, 16'd8271, 16'd58579, 16'd6927, 16'd49616, 16'd13415, 16'd39533, 16'd59517, 16'd47066, 16'd51683, 16'd62374, 16'd2185, 16'd53902, 16'd39225, 16'd21562, 16'd56721, 16'd2590, 16'd38249, 16'd47756, 16'd62383, 16'd42949, 16'd56340});
	test_expansion(128'h0e2d0c820e1f34853114f25e5ef75f2d, {16'd19255, 16'd48708, 16'd36878, 16'd52758, 16'd13450, 16'd63964, 16'd53032, 16'd6616, 16'd42301, 16'd47312, 16'd12203, 16'd26254, 16'd406, 16'd43278, 16'd59403, 16'd38880, 16'd28826, 16'd51308, 16'd28771, 16'd17589, 16'd24857, 16'd26404, 16'd43803, 16'd21139, 16'd25435, 16'd40187});
	test_expansion(128'h9356b9ffaed9f1be4694b7ba51b05648, {16'd25812, 16'd2368, 16'd42607, 16'd33615, 16'd30480, 16'd27908, 16'd61804, 16'd9184, 16'd51313, 16'd9251, 16'd939, 16'd39660, 16'd28756, 16'd16601, 16'd19744, 16'd47653, 16'd2999, 16'd49838, 16'd43125, 16'd26480, 16'd29098, 16'd26602, 16'd20121, 16'd46233, 16'd37647, 16'd54563});
	test_expansion(128'h256100dd3aa2cae0f88dfbace1465428, {16'd51165, 16'd10633, 16'd15354, 16'd33536, 16'd57963, 16'd33423, 16'd148, 16'd61450, 16'd57032, 16'd20060, 16'd23816, 16'd5781, 16'd42323, 16'd30074, 16'd24610, 16'd37342, 16'd7821, 16'd47360, 16'd35203, 16'd23230, 16'd40727, 16'd21793, 16'd59622, 16'd34098, 16'd28149, 16'd16745});
	test_expansion(128'hd7b0b22baeed36e5c9147a0ecc5b73f7, {16'd38420, 16'd7851, 16'd52503, 16'd33853, 16'd34724, 16'd7078, 16'd16680, 16'd3941, 16'd4456, 16'd46027, 16'd39637, 16'd64700, 16'd21730, 16'd22261, 16'd43689, 16'd20953, 16'd26971, 16'd57700, 16'd34381, 16'd45254, 16'd58562, 16'd42574, 16'd56332, 16'd27008, 16'd11268, 16'd2338});
	test_expansion(128'hc8c67c238edcf442ed8ffa7cbdbdf4c3, {16'd50071, 16'd30717, 16'd9715, 16'd25972, 16'd57226, 16'd27253, 16'd38386, 16'd8544, 16'd55785, 16'd56167, 16'd18841, 16'd28944, 16'd30458, 16'd42094, 16'd52307, 16'd60742, 16'd11565, 16'd59368, 16'd15301, 16'd43901, 16'd34226, 16'd47294, 16'd45118, 16'd56282, 16'd34348, 16'd35030});
	test_expansion(128'h24a090f1ff8606e1e504ed37501c9a2b, {16'd22978, 16'd6288, 16'd43234, 16'd17478, 16'd9287, 16'd50577, 16'd918, 16'd53133, 16'd3722, 16'd6995, 16'd15970, 16'd45849, 16'd13332, 16'd1780, 16'd46694, 16'd22733, 16'd51105, 16'd31263, 16'd65461, 16'd38275, 16'd39515, 16'd55864, 16'd53255, 16'd56495, 16'd60675, 16'd3769});
	test_expansion(128'h078b8e23a64afc4e5e34cee3add8fe17, {16'd15998, 16'd36309, 16'd63595, 16'd18316, 16'd31714, 16'd36752, 16'd20554, 16'd63780, 16'd34643, 16'd57204, 16'd8653, 16'd64508, 16'd54784, 16'd5308, 16'd53750, 16'd46856, 16'd17480, 16'd38668, 16'd32712, 16'd21599, 16'd33238, 16'd23784, 16'd47690, 16'd7344, 16'd17707, 16'd51733});
	test_expansion(128'h5e8f8a8d71fc255bf811e777921ff57d, {16'd31990, 16'd16797, 16'd16605, 16'd56718, 16'd39174, 16'd4245, 16'd14297, 16'd43582, 16'd51558, 16'd50822, 16'd43788, 16'd50219, 16'd49263, 16'd828, 16'd64591, 16'd58829, 16'd7237, 16'd56219, 16'd25518, 16'd28012, 16'd369, 16'd59528, 16'd17314, 16'd39034, 16'd17599, 16'd29192});
	test_expansion(128'hbb731d1f6cb10c08069bc1fa317f912c, {16'd13612, 16'd13719, 16'd63871, 16'd48314, 16'd53291, 16'd63993, 16'd45996, 16'd28150, 16'd30424, 16'd54272, 16'd42619, 16'd40936, 16'd29632, 16'd36702, 16'd61400, 16'd13495, 16'd39972, 16'd30805, 16'd42675, 16'd43307, 16'd8733, 16'd24761, 16'd7840, 16'd700, 16'd46399, 16'd63403});
	test_expansion(128'hf5300f61ab770d1150772f9e0173d9e2, {16'd17696, 16'd40705, 16'd30603, 16'd280, 16'd54316, 16'd5372, 16'd1418, 16'd44403, 16'd28639, 16'd29625, 16'd19311, 16'd30126, 16'd61813, 16'd18370, 16'd29447, 16'd49748, 16'd26282, 16'd9951, 16'd33699, 16'd39889, 16'd17238, 16'd38790, 16'd27211, 16'd56228, 16'd63395, 16'd15187});
	test_expansion(128'h22b5c179467b16c8c1fb936b3cb7292f, {16'd11301, 16'd39125, 16'd42095, 16'd35732, 16'd52588, 16'd29422, 16'd28432, 16'd58805, 16'd59071, 16'd54325, 16'd10264, 16'd38780, 16'd25135, 16'd65349, 16'd28117, 16'd5762, 16'd34650, 16'd33767, 16'd56155, 16'd16065, 16'd54155, 16'd49113, 16'd6528, 16'd45485, 16'd62605, 16'd52206});
	test_expansion(128'h7dcc5b7314a0f23c5081874a210e92d8, {16'd1764, 16'd5244, 16'd5055, 16'd43393, 16'd1241, 16'd15528, 16'd30463, 16'd6026, 16'd11532, 16'd17415, 16'd6885, 16'd40813, 16'd5975, 16'd30491, 16'd25615, 16'd55116, 16'd32374, 16'd28309, 16'd4055, 16'd3421, 16'd55800, 16'd40484, 16'd23376, 16'd17217, 16'd30883, 16'd41547});
	test_expansion(128'hbc473eb8f349880da01d1cfed4b2eff8, {16'd3329, 16'd25223, 16'd57639, 16'd56674, 16'd64379, 16'd61562, 16'd19354, 16'd22164, 16'd36725, 16'd6190, 16'd17854, 16'd56000, 16'd58920, 16'd64600, 16'd11537, 16'd42413, 16'd24591, 16'd15660, 16'd35268, 16'd3711, 16'd60307, 16'd33419, 16'd52687, 16'd19450, 16'd7536, 16'd60455});
	test_expansion(128'hc3dd90236a8df45053b2a7f8dc83cf9a, {16'd34369, 16'd18052, 16'd30873, 16'd35972, 16'd16874, 16'd62777, 16'd33831, 16'd64531, 16'd16174, 16'd15552, 16'd63103, 16'd59892, 16'd49286, 16'd48930, 16'd24301, 16'd25818, 16'd7167, 16'd17958, 16'd60999, 16'd32661, 16'd20860, 16'd30304, 16'd61348, 16'd49119, 16'd16395, 16'd31421});
	test_expansion(128'hcb1712e6354c5ab864bdba0238f86aa1, {16'd9139, 16'd44309, 16'd41406, 16'd51237, 16'd48141, 16'd61357, 16'd28129, 16'd13883, 16'd19140, 16'd49636, 16'd25899, 16'd13958, 16'd46634, 16'd21644, 16'd48254, 16'd28993, 16'd23032, 16'd13069, 16'd18932, 16'd32524, 16'd42725, 16'd39074, 16'd34343, 16'd39058, 16'd55921, 16'd13270});
	test_expansion(128'h630ebf2c34c66c3da37cf0be189003b8, {16'd22570, 16'd3966, 16'd9685, 16'd60249, 16'd26468, 16'd15135, 16'd36759, 16'd25351, 16'd58089, 16'd10598, 16'd4382, 16'd34573, 16'd57534, 16'd11880, 16'd41581, 16'd27279, 16'd26119, 16'd21194, 16'd25693, 16'd29041, 16'd33341, 16'd42853, 16'd37132, 16'd61911, 16'd5835, 16'd2456});
	test_expansion(128'hf68e2f9f9d6c99163858fbb6f0612d44, {16'd34892, 16'd51177, 16'd35536, 16'd47613, 16'd30708, 16'd42852, 16'd35171, 16'd43108, 16'd6924, 16'd35499, 16'd12214, 16'd14125, 16'd2655, 16'd22637, 16'd13369, 16'd47573, 16'd17119, 16'd41684, 16'd54009, 16'd55514, 16'd3623, 16'd56671, 16'd16521, 16'd6391, 16'd6445, 16'd64561});
	test_expansion(128'hae7fa255c92486adf114e3eaaf76bdf0, {16'd13723, 16'd39106, 16'd1427, 16'd8006, 16'd15903, 16'd13625, 16'd36173, 16'd27948, 16'd12984, 16'd36060, 16'd55206, 16'd58587, 16'd8332, 16'd5969, 16'd2723, 16'd25214, 16'd36102, 16'd14907, 16'd29489, 16'd6286, 16'd2472, 16'd25434, 16'd26297, 16'd63298, 16'd29321, 16'd61955});
	test_expansion(128'h47345c2f94eaf6639ff7b16726844d02, {16'd57337, 16'd57006, 16'd61661, 16'd1416, 16'd9542, 16'd1578, 16'd62077, 16'd20192, 16'd13261, 16'd32567, 16'd2097, 16'd14565, 16'd24159, 16'd60264, 16'd43106, 16'd127, 16'd59662, 16'd2422, 16'd59047, 16'd63585, 16'd13831, 16'd13249, 16'd55111, 16'd48660, 16'd64279, 16'd22588});
	test_expansion(128'h652f9ad760c963ed3f5a0477bccbf317, {16'd12068, 16'd37995, 16'd37683, 16'd3052, 16'd36100, 16'd50965, 16'd15511, 16'd41882, 16'd26403, 16'd59150, 16'd20190, 16'd21486, 16'd20055, 16'd51339, 16'd57504, 16'd10981, 16'd46000, 16'd42364, 16'd6244, 16'd856, 16'd5384, 16'd44879, 16'd4022, 16'd34108, 16'd29941, 16'd51835});
	test_expansion(128'hf7397007183cf5c14e29e4c49a151e74, {16'd61448, 16'd18107, 16'd12429, 16'd24345, 16'd27698, 16'd12005, 16'd43855, 16'd5850, 16'd50938, 16'd8189, 16'd736, 16'd14865, 16'd9598, 16'd57896, 16'd61828, 16'd42188, 16'd3975, 16'd4444, 16'd60719, 16'd34066, 16'd49586, 16'd16964, 16'd39611, 16'd36974, 16'd10290, 16'd35766});
	test_expansion(128'h96f67dde8e2cb9f7ebf76c367d322733, {16'd49622, 16'd1016, 16'd2516, 16'd39411, 16'd209, 16'd28475, 16'd65227, 16'd31970, 16'd62625, 16'd43530, 16'd40625, 16'd52856, 16'd26844, 16'd32166, 16'd39381, 16'd28631, 16'd365, 16'd62575, 16'd7365, 16'd5419, 16'd17203, 16'd8537, 16'd37086, 16'd12570, 16'd37375, 16'd34012});
	test_expansion(128'h7b0b647398a7863324e21029e346a47d, {16'd62917, 16'd22625, 16'd53275, 16'd36277, 16'd24622, 16'd39291, 16'd14316, 16'd48910, 16'd1025, 16'd62910, 16'd57989, 16'd54096, 16'd39795, 16'd1597, 16'd1508, 16'd46983, 16'd49100, 16'd24916, 16'd1745, 16'd1115, 16'd56735, 16'd2529, 16'd62627, 16'd53835, 16'd48430, 16'd35907});
	test_expansion(128'hfe209557b4c20428e21e03e66c8d3ef3, {16'd49124, 16'd27859, 16'd34652, 16'd22051, 16'd65068, 16'd35335, 16'd9148, 16'd41389, 16'd3084, 16'd44298, 16'd7695, 16'd59889, 16'd46266, 16'd20587, 16'd58582, 16'd13222, 16'd23056, 16'd24912, 16'd65308, 16'd31013, 16'd46882, 16'd41499, 16'd23635, 16'd1344, 16'd52012, 16'd51085});
	test_expansion(128'h7fb0d611ccc44e5ed292b1e47b0345b9, {16'd5421, 16'd64829, 16'd55067, 16'd8306, 16'd17592, 16'd43110, 16'd11732, 16'd3556, 16'd63900, 16'd20217, 16'd31878, 16'd7364, 16'd54503, 16'd62896, 16'd44455, 16'd30581, 16'd56370, 16'd20836, 16'd20739, 16'd53735, 16'd40094, 16'd8424, 16'd12709, 16'd4670, 16'd15819, 16'd31038});
	test_expansion(128'hf3ae055de56db1d76c3c91d1b3e79695, {16'd19224, 16'd63801, 16'd39262, 16'd10021, 16'd18543, 16'd55936, 16'd30308, 16'd7337, 16'd48255, 16'd33427, 16'd44662, 16'd3745, 16'd53360, 16'd44163, 16'd51611, 16'd38882, 16'd11118, 16'd8044, 16'd55008, 16'd14229, 16'd2688, 16'd39276, 16'd33487, 16'd17734, 16'd15384, 16'd5100});
	test_expansion(128'h6ea593df1041452442d328bfb461678e, {16'd15039, 16'd36923, 16'd63084, 16'd55927, 16'd24383, 16'd9926, 16'd3698, 16'd43169, 16'd30031, 16'd17588, 16'd56202, 16'd46877, 16'd59649, 16'd25832, 16'd14342, 16'd24964, 16'd4696, 16'd36410, 16'd53724, 16'd32761, 16'd21415, 16'd34691, 16'd26331, 16'd35953, 16'd6943, 16'd42605});
	test_expansion(128'hef18741ca730420cb80c8e86ac7009a8, {16'd44642, 16'd34524, 16'd61665, 16'd45942, 16'd43304, 16'd56841, 16'd60985, 16'd19272, 16'd38373, 16'd20918, 16'd998, 16'd7620, 16'd36930, 16'd59969, 16'd32021, 16'd60867, 16'd30489, 16'd16046, 16'd57056, 16'd51324, 16'd19973, 16'd26539, 16'd2281, 16'd44955, 16'd1672, 16'd22883});
	test_expansion(128'h1405d5839f4acbf7fa6b73a2083fe47c, {16'd55479, 16'd4015, 16'd26377, 16'd16602, 16'd801, 16'd49847, 16'd8291, 16'd13372, 16'd57021, 16'd60606, 16'd6958, 16'd50307, 16'd51326, 16'd3406, 16'd13075, 16'd36133, 16'd61500, 16'd23865, 16'd20515, 16'd53375, 16'd42672, 16'd32358, 16'd48549, 16'd47345, 16'd14295, 16'd4379});
	test_expansion(128'h221527d41de76704d22d6287c394c1d5, {16'd21001, 16'd45415, 16'd50483, 16'd21971, 16'd19067, 16'd2193, 16'd1758, 16'd14114, 16'd39798, 16'd46390, 16'd37556, 16'd31725, 16'd21155, 16'd24449, 16'd7079, 16'd64109, 16'd14415, 16'd3940, 16'd43570, 16'd51105, 16'd7904, 16'd14627, 16'd11617, 16'd34982, 16'd33444, 16'd56367});
	test_expansion(128'hedc5adab74184b10be41e46797f6bde0, {16'd36732, 16'd61017, 16'd8791, 16'd197, 16'd37007, 16'd12486, 16'd24765, 16'd50558, 16'd1905, 16'd36756, 16'd2105, 16'd28040, 16'd11775, 16'd39226, 16'd28716, 16'd54819, 16'd27992, 16'd2895, 16'd29578, 16'd31121, 16'd12333, 16'd37615, 16'd58233, 16'd10234, 16'd22341, 16'd22537});
	test_expansion(128'h79a372cf98296b6d20f630d1d2e98bf3, {16'd12693, 16'd55603, 16'd54377, 16'd59079, 16'd35843, 16'd48103, 16'd1042, 16'd48941, 16'd41572, 16'd62509, 16'd25449, 16'd49618, 16'd16357, 16'd4150, 16'd42038, 16'd57202, 16'd62953, 16'd22814, 16'd4832, 16'd26007, 16'd18505, 16'd16511, 16'd8658, 16'd60445, 16'd19165, 16'd9533});
	test_expansion(128'h2fe677790f9688edf2bfae97d6796a95, {16'd5830, 16'd15314, 16'd49553, 16'd16473, 16'd63657, 16'd17476, 16'd10998, 16'd18124, 16'd51869, 16'd63792, 16'd64284, 16'd53238, 16'd38858, 16'd2147, 16'd38338, 16'd62438, 16'd39566, 16'd63105, 16'd63946, 16'd63898, 16'd55551, 16'd52666, 16'd20367, 16'd45008, 16'd31963, 16'd49898});
	test_expansion(128'h401bd336c64bcdcc34ebac419e0d43a7, {16'd18683, 16'd65118, 16'd47534, 16'd15620, 16'd57718, 16'd49097, 16'd19943, 16'd56227, 16'd37146, 16'd17604, 16'd12662, 16'd17104, 16'd30426, 16'd1212, 16'd29503, 16'd45617, 16'd65247, 16'd45833, 16'd29882, 16'd40656, 16'd43771, 16'd1181, 16'd48660, 16'd40270, 16'd13800, 16'd53079});
	test_expansion(128'h221fe579d9e308ba372f3d5440432523, {16'd49074, 16'd31288, 16'd39728, 16'd15497, 16'd27979, 16'd28384, 16'd51392, 16'd5827, 16'd2732, 16'd45143, 16'd45411, 16'd54550, 16'd7049, 16'd29951, 16'd5449, 16'd25764, 16'd49113, 16'd9939, 16'd19655, 16'd5936, 16'd4168, 16'd54596, 16'd61309, 16'd50672, 16'd38414, 16'd52378});
	test_expansion(128'hd8a52ef8140c76d9e50cadbeec680ab8, {16'd48176, 16'd48502, 16'd60042, 16'd33374, 16'd42130, 16'd35243, 16'd42207, 16'd50233, 16'd5964, 16'd51280, 16'd1291, 16'd47734, 16'd575, 16'd16358, 16'd63382, 16'd2937, 16'd8858, 16'd4704, 16'd37981, 16'd13959, 16'd7306, 16'd50420, 16'd40520, 16'd23412, 16'd38274, 16'd2681});
	test_expansion(128'hdade1e63b4258bd6e4451ef416929e70, {16'd60709, 16'd58384, 16'd23106, 16'd43591, 16'd52064, 16'd52681, 16'd33140, 16'd20962, 16'd20284, 16'd58596, 16'd44464, 16'd21478, 16'd62834, 16'd52411, 16'd6588, 16'd39521, 16'd8479, 16'd10698, 16'd31656, 16'd15688, 16'd29113, 16'd64452, 16'd37480, 16'd10152, 16'd38735, 16'd38347});
	test_expansion(128'hf79adf45a986db5d245c507424c53b47, {16'd53256, 16'd4232, 16'd11475, 16'd24043, 16'd12728, 16'd14958, 16'd63593, 16'd39578, 16'd57482, 16'd18252, 16'd58496, 16'd658, 16'd50789, 16'd26624, 16'd17815, 16'd21028, 16'd35018, 16'd27962, 16'd7384, 16'd34146, 16'd21347, 16'd9093, 16'd22698, 16'd31157, 16'd25409, 16'd8967});
	test_expansion(128'h1047a7dfab589a40d77dab960cf2f89a, {16'd51801, 16'd21057, 16'd44687, 16'd28394, 16'd4962, 16'd59773, 16'd61070, 16'd5887, 16'd370, 16'd11304, 16'd7891, 16'd5056, 16'd21876, 16'd43091, 16'd23906, 16'd19154, 16'd34678, 16'd25441, 16'd61624, 16'd39846, 16'd5127, 16'd20806, 16'd12406, 16'd43287, 16'd49559, 16'd29698});
	test_expansion(128'h70391fb2c14779e07efdfb4153ddf100, {16'd20585, 16'd36869, 16'd57694, 16'd45985, 16'd14200, 16'd41841, 16'd47277, 16'd37873, 16'd6672, 16'd8420, 16'd64249, 16'd10234, 16'd19035, 16'd50190, 16'd29561, 16'd51738, 16'd23063, 16'd39331, 16'd57571, 16'd23687, 16'd47031, 16'd30928, 16'd26325, 16'd2784, 16'd55923, 16'd9840});
	test_expansion(128'h55d3f84e46f1c0842053b89ce1aa0b89, {16'd32004, 16'd14491, 16'd28410, 16'd5296, 16'd8467, 16'd60764, 16'd49403, 16'd36612, 16'd4866, 16'd2216, 16'd45338, 16'd7227, 16'd19512, 16'd44945, 16'd56032, 16'd47761, 16'd8923, 16'd26418, 16'd53549, 16'd23500, 16'd45139, 16'd36987, 16'd34571, 16'd27343, 16'd4109, 16'd3349});
	test_expansion(128'hdfe2b83c45797ddb6c4164a1dee6a1d0, {16'd10522, 16'd18477, 16'd50096, 16'd46035, 16'd61513, 16'd7631, 16'd8416, 16'd25232, 16'd18408, 16'd46616, 16'd58119, 16'd35317, 16'd27930, 16'd2109, 16'd49221, 16'd12744, 16'd37516, 16'd63239, 16'd13129, 16'd10529, 16'd8455, 16'd45486, 16'd52584, 16'd1624, 16'd22435, 16'd4057});
	test_expansion(128'h6527a3fa52fc5800a5b615e961c0078b, {16'd51077, 16'd42503, 16'd60913, 16'd19413, 16'd63505, 16'd4163, 16'd23163, 16'd21598, 16'd48372, 16'd10356, 16'd10917, 16'd8222, 16'd9756, 16'd41878, 16'd10331, 16'd52441, 16'd43882, 16'd15865, 16'd42547, 16'd44978, 16'd57004, 16'd51441, 16'd37710, 16'd9382, 16'd16201, 16'd10473});
	test_expansion(128'hef411f0654a810e0e0c14a7d62dda1c9, {16'd57449, 16'd14531, 16'd28519, 16'd28870, 16'd22301, 16'd28666, 16'd20936, 16'd61856, 16'd59851, 16'd8338, 16'd2393, 16'd24120, 16'd5665, 16'd3749, 16'd56862, 16'd38292, 16'd16030, 16'd51185, 16'd63096, 16'd55578, 16'd13396, 16'd36098, 16'd29027, 16'd12296, 16'd61888, 16'd43599});
	test_expansion(128'h3fe5b47899cd2e66efb136d74c1a1800, {16'd28689, 16'd57530, 16'd57697, 16'd5964, 16'd31233, 16'd5911, 16'd50692, 16'd49921, 16'd919, 16'd56694, 16'd13976, 16'd49891, 16'd5030, 16'd14188, 16'd49769, 16'd18981, 16'd39726, 16'd11231, 16'd51436, 16'd52983, 16'd965, 16'd64723, 16'd7973, 16'd965, 16'd18442, 16'd28025});
	test_expansion(128'he0c3c96782661fb584480f14c5c88298, {16'd46802, 16'd39692, 16'd27002, 16'd44900, 16'd8538, 16'd9093, 16'd35387, 16'd46141, 16'd12564, 16'd64801, 16'd53983, 16'd13255, 16'd12748, 16'd30382, 16'd10734, 16'd43483, 16'd23950, 16'd22035, 16'd23730, 16'd18, 16'd36016, 16'd32136, 16'd39287, 16'd532, 16'd34481, 16'd3183});
	test_expansion(128'h276f336d83d94d3fbb874c1bbfe70694, {16'd32312, 16'd42247, 16'd11843, 16'd8499, 16'd50209, 16'd12567, 16'd64953, 16'd56338, 16'd53953, 16'd48196, 16'd16232, 16'd31664, 16'd41846, 16'd36282, 16'd54891, 16'd53187, 16'd39120, 16'd3443, 16'd31154, 16'd53657, 16'd47395, 16'd56256, 16'd44586, 16'd48574, 16'd27277, 16'd9716});
	test_expansion(128'h9e11ae3274a38078df19909ffc3ce706, {16'd46775, 16'd33130, 16'd35760, 16'd41421, 16'd31373, 16'd27609, 16'd18207, 16'd31839, 16'd43083, 16'd35154, 16'd54685, 16'd1746, 16'd1818, 16'd24216, 16'd2455, 16'd40542, 16'd28825, 16'd29200, 16'd39045, 16'd36703, 16'd61028, 16'd57432, 16'd40121, 16'd63209, 16'd38172, 16'd28909});
	test_expansion(128'hf07d874c9642c47fef1381cd46b64cc5, {16'd24063, 16'd22413, 16'd1414, 16'd17869, 16'd25288, 16'd54764, 16'd24011, 16'd32061, 16'd32093, 16'd64652, 16'd4239, 16'd10992, 16'd33403, 16'd47228, 16'd42931, 16'd24954, 16'd45568, 16'd60907, 16'd32321, 16'd28402, 16'd32996, 16'd26683, 16'd16325, 16'd57883, 16'd31646, 16'd60165});
	test_expansion(128'h59a9a9acf2f2729c5f636e7ee53707b1, {16'd37818, 16'd10087, 16'd62177, 16'd33199, 16'd50667, 16'd41204, 16'd2388, 16'd13372, 16'd51363, 16'd29464, 16'd36112, 16'd4154, 16'd59258, 16'd25590, 16'd11868, 16'd25986, 16'd54853, 16'd50732, 16'd5385, 16'd57407, 16'd49309, 16'd26087, 16'd31795, 16'd35867, 16'd22844, 16'd49462});
	test_expansion(128'h46a43dd9d8c2092099df8b3ca925f878, {16'd32342, 16'd50246, 16'd34587, 16'd25772, 16'd34387, 16'd174, 16'd48769, 16'd5541, 16'd54700, 16'd36229, 16'd40344, 16'd24309, 16'd11838, 16'd46007, 16'd55203, 16'd39750, 16'd24774, 16'd10511, 16'd19967, 16'd26318, 16'd63263, 16'd20171, 16'd24282, 16'd63816, 16'd46458, 16'd41249});
	test_expansion(128'h3dc4f0e4323d2d16b2b44e300a00e4ea, {16'd7539, 16'd46089, 16'd33757, 16'd64561, 16'd37014, 16'd63371, 16'd49660, 16'd5395, 16'd41526, 16'd19200, 16'd18248, 16'd53584, 16'd30682, 16'd35647, 16'd17753, 16'd13581, 16'd20936, 16'd48070, 16'd40452, 16'd61946, 16'd49738, 16'd3770, 16'd47948, 16'd17819, 16'd48766, 16'd25662});
	test_expansion(128'hfe4b649c8474ab4ea746ee7235e5e771, {16'd58377, 16'd31238, 16'd22076, 16'd60862, 16'd42081, 16'd38836, 16'd47336, 16'd698, 16'd36999, 16'd52032, 16'd43851, 16'd32959, 16'd64447, 16'd40025, 16'd42574, 16'd6558, 16'd47254, 16'd56390, 16'd54015, 16'd60969, 16'd2802, 16'd30329, 16'd37431, 16'd18179, 16'd53755, 16'd38667});
	test_expansion(128'h3314e1e24b15cd82ee279c7476c2fb62, {16'd20566, 16'd41658, 16'd45247, 16'd15969, 16'd42082, 16'd40386, 16'd13542, 16'd2975, 16'd50198, 16'd52405, 16'd10466, 16'd8689, 16'd35667, 16'd16105, 16'd19202, 16'd47444, 16'd14469, 16'd52656, 16'd36374, 16'd24504, 16'd31642, 16'd20607, 16'd27712, 16'd54495, 16'd43378, 16'd51729});
	test_expansion(128'h1f10110de3ace61b47c5b4c237c4f943, {16'd20665, 16'd13031, 16'd63399, 16'd20503, 16'd15312, 16'd25367, 16'd53739, 16'd7496, 16'd48479, 16'd1360, 16'd19198, 16'd31610, 16'd47989, 16'd42444, 16'd60955, 16'd10525, 16'd34952, 16'd10109, 16'd54981, 16'd34665, 16'd15698, 16'd62932, 16'd54199, 16'd54716, 16'd49830, 16'd53511});
	test_expansion(128'hb04350dae98a9e02ec41a37d0a684425, {16'd29817, 16'd2926, 16'd31280, 16'd14652, 16'd3781, 16'd26655, 16'd9703, 16'd20885, 16'd29783, 16'd32040, 16'd45682, 16'd25213, 16'd61918, 16'd1806, 16'd30654, 16'd55135, 16'd8054, 16'd2561, 16'd12649, 16'd4751, 16'd60868, 16'd20009, 16'd31405, 16'd51865, 16'd37570, 16'd846});
	test_expansion(128'h8d5b625229e3c99ffb9e7ec5ed6b32a8, {16'd31699, 16'd26960, 16'd37588, 16'd3375, 16'd8815, 16'd60120, 16'd14956, 16'd47009, 16'd36180, 16'd46912, 16'd42314, 16'd29444, 16'd56025, 16'd60745, 16'd14648, 16'd30757, 16'd33038, 16'd25578, 16'd25421, 16'd12496, 16'd34440, 16'd2820, 16'd34166, 16'd21296, 16'd50658, 16'd44678});
	test_expansion(128'hc423fbd39e847ff2c855f5a7eafbedb6, {16'd7126, 16'd36689, 16'd59225, 16'd27012, 16'd40797, 16'd27068, 16'd32181, 16'd31163, 16'd4657, 16'd28377, 16'd21387, 16'd63241, 16'd49433, 16'd22891, 16'd17877, 16'd17864, 16'd60241, 16'd42524, 16'd29855, 16'd53836, 16'd54354, 16'd35554, 16'd53353, 16'd52795, 16'd50746, 16'd31775});
	test_expansion(128'h849ee45ffa6c68b8524b69ed4369bca6, {16'd19692, 16'd28582, 16'd56429, 16'd56638, 16'd33086, 16'd5021, 16'd25438, 16'd60937, 16'd51644, 16'd20422, 16'd36559, 16'd5602, 16'd34721, 16'd28325, 16'd39699, 16'd5322, 16'd53896, 16'd58360, 16'd47502, 16'd62949, 16'd8993, 16'd9079, 16'd61055, 16'd5867, 16'd56603, 16'd62826});
	test_expansion(128'h67b2185020ca97e13b6d6d9fdec9d3f8, {16'd13234, 16'd59518, 16'd43273, 16'd62904, 16'd51377, 16'd32280, 16'd28948, 16'd5394, 16'd28871, 16'd15591, 16'd32097, 16'd38690, 16'd51960, 16'd56655, 16'd45038, 16'd10715, 16'd1013, 16'd62332, 16'd25712, 16'd46181, 16'd51349, 16'd19623, 16'd29900, 16'd26666, 16'd64743, 16'd19802});
	test_expansion(128'h40b581f6052cd77c38f52539eb2c243a, {16'd33549, 16'd30504, 16'd2987, 16'd56168, 16'd29028, 16'd3061, 16'd33111, 16'd46221, 16'd10053, 16'd57602, 16'd35755, 16'd14853, 16'd62932, 16'd13939, 16'd42634, 16'd31658, 16'd35846, 16'd23303, 16'd43637, 16'd28547, 16'd26323, 16'd9899, 16'd58451, 16'd24147, 16'd57405, 16'd19947});
	test_expansion(128'h3eca652f62edf05dec776cdd1e6bca1c, {16'd22806, 16'd53877, 16'd28723, 16'd30385, 16'd42381, 16'd5025, 16'd55673, 16'd11059, 16'd57167, 16'd22985, 16'd18152, 16'd38887, 16'd23038, 16'd8036, 16'd42607, 16'd35012, 16'd21032, 16'd20508, 16'd42606, 16'd25688, 16'd47472, 16'd7456, 16'd34774, 16'd36381, 16'd57941, 16'd23731});
	test_expansion(128'hd6cdcba01592c1ec78da34a416d372ab, {16'd6462, 16'd28495, 16'd36067, 16'd47247, 16'd21891, 16'd34145, 16'd16832, 16'd9937, 16'd57325, 16'd42456, 16'd28406, 16'd44621, 16'd8664, 16'd22251, 16'd1509, 16'd59272, 16'd48728, 16'd5979, 16'd32416, 16'd14232, 16'd7567, 16'd6607, 16'd44984, 16'd25353, 16'd38844, 16'd23968});
	test_expansion(128'h928f826b1f930262005819c1a311b0db, {16'd14293, 16'd27235, 16'd15877, 16'd2169, 16'd61364, 16'd22309, 16'd3600, 16'd65018, 16'd18937, 16'd46595, 16'd35013, 16'd42333, 16'd60073, 16'd32524, 16'd63740, 16'd58020, 16'd16467, 16'd55321, 16'd11100, 16'd25979, 16'd2129, 16'd28387, 16'd31162, 16'd3823, 16'd30470, 16'd23159});
	test_expansion(128'h2dd18e494a90ae05eeb6291ade81195c, {16'd32102, 16'd55127, 16'd12788, 16'd5470, 16'd42511, 16'd36596, 16'd31997, 16'd1159, 16'd5559, 16'd54420, 16'd64839, 16'd26312, 16'd23538, 16'd4605, 16'd61454, 16'd47670, 16'd26471, 16'd5058, 16'd45518, 16'd23259, 16'd55476, 16'd28231, 16'd34065, 16'd52536, 16'd59494, 16'd54430});
	test_expansion(128'h258e8f7d98888b9c534a665c2f474147, {16'd43836, 16'd30722, 16'd58796, 16'd3726, 16'd9671, 16'd13727, 16'd24344, 16'd22835, 16'd4538, 16'd35599, 16'd12510, 16'd49259, 16'd22439, 16'd56588, 16'd8547, 16'd48954, 16'd23128, 16'd19049, 16'd28523, 16'd24617, 16'd28090, 16'd51671, 16'd38363, 16'd29419, 16'd41541, 16'd49374});
	test_expansion(128'hb8767cde9763357d00f4d2c4daff5f51, {16'd23089, 16'd25364, 16'd51863, 16'd26423, 16'd10036, 16'd8664, 16'd48746, 16'd47148, 16'd28848, 16'd64291, 16'd48615, 16'd32714, 16'd37066, 16'd57780, 16'd15657, 16'd30118, 16'd6931, 16'd19263, 16'd34809, 16'd51025, 16'd33476, 16'd49021, 16'd20174, 16'd58789, 16'd27826, 16'd48420});
	test_expansion(128'hddb1b45072c57df7200db03d3603bb92, {16'd7931, 16'd36173, 16'd54071, 16'd8289, 16'd14339, 16'd15451, 16'd9140, 16'd61125, 16'd52655, 16'd64018, 16'd10629, 16'd31953, 16'd7371, 16'd40992, 16'd46985, 16'd6642, 16'd28619, 16'd46042, 16'd55070, 16'd36263, 16'd58192, 16'd11294, 16'd12439, 16'd31681, 16'd43272, 16'd47608});
	test_expansion(128'h02ce5bfae94a7ea028cc3441f5f31183, {16'd64517, 16'd35845, 16'd8948, 16'd47582, 16'd56790, 16'd14219, 16'd662, 16'd58769, 16'd42819, 16'd22531, 16'd37663, 16'd6930, 16'd35977, 16'd12397, 16'd36672, 16'd5493, 16'd4077, 16'd62492, 16'd42439, 16'd33893, 16'd40641, 16'd41281, 16'd5601, 16'd61263, 16'd8875, 16'd27970});
	test_expansion(128'hea7d5e5f217d8b4c6ab0393dc34a8685, {16'd16348, 16'd32905, 16'd65053, 16'd41580, 16'd10070, 16'd56218, 16'd57028, 16'd34980, 16'd64886, 16'd18847, 16'd36938, 16'd18385, 16'd45371, 16'd17436, 16'd31434, 16'd32269, 16'd22912, 16'd1550, 16'd11535, 16'd11999, 16'd15712, 16'd44692, 16'd57238, 16'd37811, 16'd48584, 16'd21316});
	test_expansion(128'hd12d5df801e84586d5d362d62261836f, {16'd21060, 16'd25690, 16'd48424, 16'd50225, 16'd13482, 16'd60502, 16'd2036, 16'd3517, 16'd9725, 16'd40171, 16'd64568, 16'd37007, 16'd33583, 16'd27697, 16'd51233, 16'd65248, 16'd12095, 16'd1211, 16'd25779, 16'd5173, 16'd13056, 16'd27092, 16'd22842, 16'd22759, 16'd9042, 16'd30307});
	test_expansion(128'h6435600f01b7f274eba1ce6b7a1ef3cc, {16'd30236, 16'd16466, 16'd5791, 16'd36254, 16'd27734, 16'd23485, 16'd5795, 16'd63023, 16'd40666, 16'd49036, 16'd25913, 16'd39085, 16'd4971, 16'd24024, 16'd42120, 16'd48472, 16'd24977, 16'd60076, 16'd47498, 16'd42023, 16'd54088, 16'd59706, 16'd46065, 16'd42515, 16'd51036, 16'd16590});
	test_expansion(128'h4b99aa496ceddb5161bea9bf0f6d1209, {16'd27789, 16'd1963, 16'd35080, 16'd47561, 16'd23155, 16'd55393, 16'd20758, 16'd30484, 16'd2753, 16'd57420, 16'd53504, 16'd62656, 16'd23696, 16'd6495, 16'd13122, 16'd49084, 16'd41816, 16'd42235, 16'd22614, 16'd52051, 16'd21656, 16'd44720, 16'd11774, 16'd4415, 16'd43199, 16'd9858});
	test_expansion(128'h914d827f3b24a0ddc3d0e5e7d8258072, {16'd26115, 16'd13771, 16'd60186, 16'd7837, 16'd61051, 16'd2362, 16'd7714, 16'd44790, 16'd13858, 16'd52383, 16'd43111, 16'd46859, 16'd17702, 16'd52974, 16'd19084, 16'd11141, 16'd239, 16'd51650, 16'd52775, 16'd26934, 16'd13224, 16'd31942, 16'd6082, 16'd39116, 16'd49156, 16'd56019});
	test_expansion(128'hfdbd705ba0140aa4f72b90d11d4bde4f, {16'd57282, 16'd20702, 16'd56638, 16'd3880, 16'd47384, 16'd46772, 16'd13807, 16'd43197, 16'd51334, 16'd47343, 16'd47662, 16'd45510, 16'd34529, 16'd47060, 16'd2923, 16'd18474, 16'd16866, 16'd23218, 16'd37015, 16'd25740, 16'd56942, 16'd44706, 16'd63214, 16'd22345, 16'd43919, 16'd12253});
	test_expansion(128'hbe064f848ad3cd26835ba85e396a192f, {16'd61265, 16'd23467, 16'd31468, 16'd20229, 16'd40964, 16'd1882, 16'd43701, 16'd27165, 16'd6820, 16'd58306, 16'd62460, 16'd56203, 16'd37864, 16'd40598, 16'd18908, 16'd20283, 16'd31252, 16'd1957, 16'd57839, 16'd58445, 16'd41346, 16'd2142, 16'd43518, 16'd54577, 16'd32794, 16'd51420});
	test_expansion(128'hc70e99c0815f004ceb5eeb195aa16db8, {16'd45077, 16'd56706, 16'd25845, 16'd15664, 16'd716, 16'd24716, 16'd58897, 16'd8201, 16'd44522, 16'd50528, 16'd38725, 16'd11049, 16'd15899, 16'd11756, 16'd38313, 16'd7091, 16'd31417, 16'd28830, 16'd26437, 16'd9425, 16'd7140, 16'd31559, 16'd15508, 16'd59958, 16'd51873, 16'd54744});
	test_expansion(128'hd4a703c58156fc7cf35ab0c1bb378c87, {16'd26498, 16'd30570, 16'd65432, 16'd60439, 16'd50512, 16'd21423, 16'd44077, 16'd44120, 16'd1989, 16'd8684, 16'd32328, 16'd21197, 16'd20859, 16'd36112, 16'd9584, 16'd30256, 16'd27883, 16'd49205, 16'd31624, 16'd11361, 16'd40690, 16'd48764, 16'd11829, 16'd59092, 16'd16401, 16'd24801});
	test_expansion(128'h54dba3a77df6735b32795dec57e9ce03, {16'd20696, 16'd1096, 16'd50313, 16'd14326, 16'd46013, 16'd8155, 16'd4997, 16'd56325, 16'd63712, 16'd28989, 16'd60335, 16'd51773, 16'd36226, 16'd54241, 16'd14956, 16'd51317, 16'd36932, 16'd2743, 16'd32707, 16'd2997, 16'd64780, 16'd30204, 16'd54889, 16'd10670, 16'd352, 16'd32284});
	test_expansion(128'h1f71d3faf3a8ad35b94a55349d4b2f38, {16'd47458, 16'd20733, 16'd1824, 16'd48634, 16'd50807, 16'd17602, 16'd50853, 16'd34100, 16'd43080, 16'd10743, 16'd36894, 16'd36329, 16'd55231, 16'd37442, 16'd56244, 16'd37319, 16'd53546, 16'd36220, 16'd36292, 16'd63989, 16'd32818, 16'd5649, 16'd6832, 16'd23192, 16'd13421, 16'd37577});
	test_expansion(128'h4c278d7d3776ee48628a20297116a504, {16'd26183, 16'd6377, 16'd34299, 16'd22351, 16'd47175, 16'd47582, 16'd11825, 16'd59864, 16'd20634, 16'd8841, 16'd27115, 16'd64246, 16'd32117, 16'd45798, 16'd8963, 16'd60274, 16'd38761, 16'd30753, 16'd18663, 16'd60947, 16'd52610, 16'd45197, 16'd6556, 16'd59815, 16'd45825, 16'd61690});
	test_expansion(128'hef7df18ac85e0ae62184c3766daa60a0, {16'd16776, 16'd17828, 16'd29223, 16'd18218, 16'd6774, 16'd58923, 16'd59376, 16'd52061, 16'd12624, 16'd11877, 16'd50486, 16'd63928, 16'd50894, 16'd28662, 16'd30988, 16'd7709, 16'd17980, 16'd16990, 16'd60225, 16'd28389, 16'd48103, 16'd39813, 16'd30136, 16'd18465, 16'd24216, 16'd36783});
	test_expansion(128'h2ca5f8282f9bbd7a682caa67ddf80ae6, {16'd26879, 16'd61021, 16'd31627, 16'd10661, 16'd20256, 16'd30339, 16'd3957, 16'd39125, 16'd61360, 16'd64369, 16'd9161, 16'd695, 16'd45290, 16'd57721, 16'd56558, 16'd44558, 16'd40739, 16'd39780, 16'd55420, 16'd3032, 16'd17753, 16'd41471, 16'd33109, 16'd949, 16'd24675, 16'd12971});
	test_expansion(128'h1b36e09fa1d9c62685f9b6a982ab60d9, {16'd28789, 16'd8295, 16'd4991, 16'd10699, 16'd28369, 16'd39035, 16'd57029, 16'd57126, 16'd28037, 16'd4221, 16'd12858, 16'd40889, 16'd32589, 16'd41962, 16'd33714, 16'd15772, 16'd45768, 16'd61521, 16'd49944, 16'd56805, 16'd8748, 16'd23393, 16'd59401, 16'd57574, 16'd14854, 16'd15304});
	test_expansion(128'h4bb1ec95c6875df6fc085eb5bc015529, {16'd36112, 16'd5133, 16'd47594, 16'd51294, 16'd63320, 16'd44106, 16'd13450, 16'd11402, 16'd18494, 16'd46486, 16'd49408, 16'd18265, 16'd50913, 16'd12092, 16'd19735, 16'd5624, 16'd30429, 16'd48283, 16'd13984, 16'd5996, 16'd51563, 16'd374, 16'd63183, 16'd34315, 16'd14505, 16'd10909});
	test_expansion(128'h6adbda9c84662818e6b29d643cfd8230, {16'd14932, 16'd61135, 16'd58744, 16'd36761, 16'd41257, 16'd13220, 16'd60257, 16'd34749, 16'd33501, 16'd59309, 16'd13358, 16'd40005, 16'd13834, 16'd28532, 16'd58138, 16'd21107, 16'd54814, 16'd29609, 16'd32545, 16'd55022, 16'd62035, 16'd15608, 16'd54183, 16'd54109, 16'd34544, 16'd11049});
	test_expansion(128'h744fdc0b8b9da106ee68b09ede156d1b, {16'd54316, 16'd64078, 16'd49148, 16'd32719, 16'd18537, 16'd2519, 16'd40160, 16'd35424, 16'd28416, 16'd54695, 16'd48844, 16'd32538, 16'd53400, 16'd46898, 16'd33773, 16'd55464, 16'd61189, 16'd56700, 16'd20177, 16'd50175, 16'd11949, 16'd44717, 16'd32336, 16'd62239, 16'd51419, 16'd36129});
	test_expansion(128'h505b72fa0b0a67464414014d55d97972, {16'd64214, 16'd15875, 16'd34944, 16'd30165, 16'd7404, 16'd12402, 16'd34322, 16'd29947, 16'd60840, 16'd4393, 16'd53658, 16'd4664, 16'd12104, 16'd30858, 16'd34264, 16'd60992, 16'd29099, 16'd19398, 16'd58588, 16'd62511, 16'd20334, 16'd42673, 16'd10460, 16'd36548, 16'd9021, 16'd4085});
	test_expansion(128'h285329322e91f2d6dd9372d4265acbee, {16'd37253, 16'd7243, 16'd58200, 16'd55222, 16'd33446, 16'd48094, 16'd19939, 16'd40369, 16'd63485, 16'd48059, 16'd30683, 16'd45952, 16'd15514, 16'd52447, 16'd12385, 16'd23492, 16'd22827, 16'd5839, 16'd49130, 16'd37801, 16'd58719, 16'd51446, 16'd60315, 16'd29187, 16'd8339, 16'd25230});
	test_expansion(128'hb3981616cb40f257d7ab4abbe49c57d2, {16'd39054, 16'd49324, 16'd53384, 16'd28766, 16'd32852, 16'd11180, 16'd62956, 16'd9297, 16'd28632, 16'd32679, 16'd49076, 16'd43272, 16'd59359, 16'd45483, 16'd42439, 16'd60220, 16'd9611, 16'd6985, 16'd18425, 16'd17329, 16'd53794, 16'd53953, 16'd28339, 16'd4601, 16'd12490, 16'd29664});
	test_expansion(128'h5a0d41085c0788baba6401517d350de3, {16'd61472, 16'd42194, 16'd45, 16'd40907, 16'd43845, 16'd41811, 16'd32050, 16'd55360, 16'd38771, 16'd41184, 16'd14826, 16'd19317, 16'd36457, 16'd57091, 16'd59070, 16'd7286, 16'd27803, 16'd2049, 16'd38066, 16'd34056, 16'd21037, 16'd26922, 16'd28056, 16'd22062, 16'd39811, 16'd30549});
	test_expansion(128'h45f23f38c430855b412c3a8730922c2a, {16'd38477, 16'd20289, 16'd26520, 16'd4454, 16'd60383, 16'd29200, 16'd57896, 16'd50989, 16'd43885, 16'd18277, 16'd17032, 16'd47382, 16'd13780, 16'd54662, 16'd43346, 16'd31549, 16'd6639, 16'd13654, 16'd1412, 16'd6898, 16'd2398, 16'd8471, 16'd64014, 16'd48168, 16'd63638, 16'd57893});
	test_expansion(128'h0b4be27601fe4703fd8019699bbee6a9, {16'd2791, 16'd3690, 16'd46022, 16'd44232, 16'd36987, 16'd41261, 16'd39579, 16'd18014, 16'd40928, 16'd53690, 16'd5535, 16'd21892, 16'd50571, 16'd63401, 16'd22730, 16'd63881, 16'd11275, 16'd58120, 16'd44037, 16'd16913, 16'd56452, 16'd60321, 16'd45675, 16'd61506, 16'd9275, 16'd20881});
	test_expansion(128'h6d93db7ba84ef86ffafd0317f1da5c81, {16'd48778, 16'd50017, 16'd13484, 16'd49552, 16'd40194, 16'd48660, 16'd17276, 16'd22592, 16'd16071, 16'd3269, 16'd15439, 16'd4396, 16'd4087, 16'd47452, 16'd60224, 16'd51746, 16'd62549, 16'd1526, 16'd52340, 16'd22580, 16'd28252, 16'd20784, 16'd1505, 16'd35013, 16'd41549, 16'd34204});
	test_expansion(128'h9b3948e7c099e4fbca495f96ba7c1228, {16'd46661, 16'd10378, 16'd60728, 16'd13003, 16'd63359, 16'd8676, 16'd51008, 16'd39020, 16'd56807, 16'd50113, 16'd47873, 16'd25933, 16'd31589, 16'd19466, 16'd31610, 16'd49071, 16'd52564, 16'd56434, 16'd4683, 16'd50291, 16'd12852, 16'd63711, 16'd43570, 16'd39081, 16'd12669, 16'd14739});
	test_expansion(128'h7837bf2be8469323804be2f98e9ad298, {16'd40949, 16'd18248, 16'd20403, 16'd46165, 16'd43314, 16'd63661, 16'd55979, 16'd24539, 16'd62122, 16'd17621, 16'd38820, 16'd24761, 16'd34982, 16'd23273, 16'd43360, 16'd16023, 16'd34890, 16'd62325, 16'd33818, 16'd42611, 16'd47135, 16'd5481, 16'd26792, 16'd15125, 16'd64576, 16'd21793});
	test_expansion(128'h5e24ca909834dd65e2646bd0bac73810, {16'd28684, 16'd35869, 16'd42395, 16'd64419, 16'd41707, 16'd13202, 16'd8565, 16'd36622, 16'd2330, 16'd47958, 16'd53159, 16'd5502, 16'd17464, 16'd30811, 16'd19482, 16'd58518, 16'd60199, 16'd36990, 16'd20584, 16'd42019, 16'd28199, 16'd15015, 16'd4851, 16'd29259, 16'd23681, 16'd5206});
	test_expansion(128'h6bb5fd8056c382ddb17c0b889a852a8c, {16'd32905, 16'd32580, 16'd6995, 16'd34897, 16'd2386, 16'd15131, 16'd14664, 16'd23133, 16'd42127, 16'd8577, 16'd18790, 16'd43522, 16'd60859, 16'd853, 16'd44680, 16'd55874, 16'd3093, 16'd47688, 16'd25481, 16'd18292, 16'd56195, 16'd14325, 16'd31391, 16'd62906, 16'd13297, 16'd38698});
	test_expansion(128'h8e7a2d0a25e41694d23334e8e02ba298, {16'd11391, 16'd61353, 16'd15563, 16'd6414, 16'd48852, 16'd12576, 16'd23240, 16'd7756, 16'd29042, 16'd60843, 16'd52301, 16'd64802, 16'd56361, 16'd27780, 16'd11531, 16'd35826, 16'd40924, 16'd42433, 16'd47197, 16'd18695, 16'd63404, 16'd62170, 16'd21252, 16'd1749, 16'd51276, 16'd31277});
	test_expansion(128'h7a6ad3cd63101abef8f7788c6945284a, {16'd53988, 16'd23424, 16'd34308, 16'd1761, 16'd11616, 16'd52837, 16'd54277, 16'd27776, 16'd32970, 16'd12557, 16'd51220, 16'd32521, 16'd16151, 16'd5146, 16'd27995, 16'd32872, 16'd18383, 16'd7973, 16'd6746, 16'd62190, 16'd5046, 16'd7859, 16'd57382, 16'd15209, 16'd29057, 16'd23298});
	test_expansion(128'h374875235daef17a03e78907f1f35d2d, {16'd15211, 16'd19923, 16'd47234, 16'd56814, 16'd52151, 16'd10361, 16'd60365, 16'd36311, 16'd7774, 16'd40111, 16'd32897, 16'd34617, 16'd32378, 16'd53047, 16'd30894, 16'd36248, 16'd23528, 16'd55667, 16'd52772, 16'd60885, 16'd34755, 16'd14011, 16'd49660, 16'd52987, 16'd16176, 16'd41795});
	test_expansion(128'hf6cf1e6408f94e7c436ddc5c42ceb2d8, {16'd49190, 16'd36157, 16'd7766, 16'd58776, 16'd42479, 16'd16931, 16'd63976, 16'd7402, 16'd59418, 16'd39501, 16'd52557, 16'd21943, 16'd36279, 16'd37509, 16'd12172, 16'd28939, 16'd58203, 16'd24403, 16'd23459, 16'd38559, 16'd52278, 16'd35376, 16'd65515, 16'd1341, 16'd46548, 16'd1210});
	test_expansion(128'he04558ee2dc362d87d15e7f616f327e2, {16'd3722, 16'd30821, 16'd64005, 16'd49518, 16'd4748, 16'd16154, 16'd59222, 16'd1152, 16'd58063, 16'd35571, 16'd42920, 16'd24393, 16'd33535, 16'd44630, 16'd39103, 16'd47327, 16'd30176, 16'd39199, 16'd43184, 16'd673, 16'd18161, 16'd9901, 16'd16992, 16'd32028, 16'd21376, 16'd7855});
	test_expansion(128'h457d88c8a0553bedf53685cf6679fa1c, {16'd26087, 16'd7807, 16'd25333, 16'd2254, 16'd64246, 16'd62763, 16'd19218, 16'd39415, 16'd56496, 16'd6712, 16'd35966, 16'd631, 16'd25079, 16'd37286, 16'd33241, 16'd59239, 16'd19310, 16'd32917, 16'd42193, 16'd45562, 16'd34129, 16'd41198, 16'd26024, 16'd26068, 16'd27892, 16'd31010});
	test_expansion(128'haedb01dc9e648ba81d667f9b6af898ad, {16'd4558, 16'd49514, 16'd39450, 16'd47888, 16'd38342, 16'd40237, 16'd64302, 16'd9001, 16'd46611, 16'd63842, 16'd11210, 16'd57513, 16'd31747, 16'd39382, 16'd13088, 16'd32687, 16'd57121, 16'd26200, 16'd58284, 16'd61179, 16'd7606, 16'd52542, 16'd36887, 16'd25466, 16'd52835, 16'd52328});
	test_expansion(128'hfc2c90fba6f4a1137d9cf834a6350722, {16'd37170, 16'd23821, 16'd30131, 16'd47470, 16'd39935, 16'd40102, 16'd9681, 16'd44646, 16'd11130, 16'd41561, 16'd46999, 16'd59301, 16'd17122, 16'd51996, 16'd60283, 16'd13576, 16'd50854, 16'd54601, 16'd42949, 16'd43802, 16'd23194, 16'd55398, 16'd23093, 16'd7611, 16'd26448, 16'd51281});
	test_expansion(128'ha5b6041924d8b065ffcfb8b20b32316d, {16'd13447, 16'd43785, 16'd25665, 16'd43367, 16'd37100, 16'd40731, 16'd7871, 16'd24925, 16'd63738, 16'd57507, 16'd50674, 16'd29757, 16'd41359, 16'd51882, 16'd35347, 16'd40649, 16'd59040, 16'd18170, 16'd21362, 16'd31001, 16'd43515, 16'd10022, 16'd29094, 16'd42110, 16'd37830, 16'd28293});
	test_expansion(128'hb0b23062086c956566c934c73cb2daed, {16'd21319, 16'd38128, 16'd24759, 16'd15961, 16'd61618, 16'd33510, 16'd15223, 16'd34757, 16'd8473, 16'd64438, 16'd22475, 16'd36916, 16'd50654, 16'd37914, 16'd5359, 16'd52126, 16'd24971, 16'd25943, 16'd37257, 16'd8795, 16'd46348, 16'd44506, 16'd63302, 16'd18732, 16'd13572, 16'd53797});
	test_expansion(128'h6a73498929dea4370644090bb08b513b, {16'd39511, 16'd7497, 16'd5494, 16'd59799, 16'd6192, 16'd53325, 16'd26371, 16'd1658, 16'd28665, 16'd25519, 16'd52111, 16'd27254, 16'd25459, 16'd8560, 16'd8318, 16'd7337, 16'd59615, 16'd47537, 16'd46605, 16'd40078, 16'd37615, 16'd6595, 16'd61469, 16'd61935, 16'd47562, 16'd28675});
	test_expansion(128'hee1723d8bde1b5424dc159ffc252cd9d, {16'd53907, 16'd783, 16'd8269, 16'd28384, 16'd2308, 16'd51998, 16'd26865, 16'd34485, 16'd41828, 16'd7498, 16'd8319, 16'd51907, 16'd7369, 16'd18526, 16'd27679, 16'd25724, 16'd34832, 16'd17100, 16'd24228, 16'd249, 16'd46239, 16'd40552, 16'd34534, 16'd3220, 16'd56208, 16'd38406});
	test_expansion(128'h318e81ae058d39a98a9761ac594c691a, {16'd57757, 16'd980, 16'd58947, 16'd8497, 16'd50425, 16'd36073, 16'd18299, 16'd36788, 16'd19773, 16'd9477, 16'd16233, 16'd61651, 16'd35698, 16'd35845, 16'd12370, 16'd22678, 16'd8230, 16'd13536, 16'd25449, 16'd1548, 16'd33399, 16'd2969, 16'd41466, 16'd57896, 16'd29620, 16'd43606});
	test_expansion(128'h54a15aff19fb0b651367253b4b5565b4, {16'd12121, 16'd53469, 16'd62158, 16'd13003, 16'd4236, 16'd43675, 16'd45653, 16'd51393, 16'd34441, 16'd38253, 16'd5936, 16'd14658, 16'd8130, 16'd16750, 16'd44493, 16'd60733, 16'd53627, 16'd40710, 16'd36814, 16'd34344, 16'd13408, 16'd57602, 16'd52650, 16'd50291, 16'd5405, 16'd21575});
	test_expansion(128'h274baccf9629e6ecb0c0f741b80844e0, {16'd58650, 16'd27558, 16'd21217, 16'd60490, 16'd57482, 16'd5778, 16'd48415, 16'd23250, 16'd20416, 16'd62640, 16'd866, 16'd41685, 16'd41015, 16'd26612, 16'd63464, 16'd38237, 16'd4537, 16'd44182, 16'd10624, 16'd62099, 16'd58354, 16'd7674, 16'd31595, 16'd6377, 16'd19296, 16'd60400});
	test_expansion(128'h616bc42cd266dac8122227b8122875ae, {16'd35281, 16'd62843, 16'd51654, 16'd61883, 16'd23718, 16'd9423, 16'd5791, 16'd45884, 16'd4199, 16'd28840, 16'd44389, 16'd5032, 16'd62481, 16'd48488, 16'd45190, 16'd22634, 16'd15146, 16'd2634, 16'd6846, 16'd11585, 16'd48091, 16'd31103, 16'd4024, 16'd4737, 16'd15695, 16'd38396});
	test_expansion(128'h273bfe49bd8a106d99af42a473123a54, {16'd48498, 16'd45519, 16'd32233, 16'd57488, 16'd18150, 16'd53745, 16'd10338, 16'd50497, 16'd39298, 16'd53859, 16'd60800, 16'd44424, 16'd63221, 16'd23213, 16'd12020, 16'd22258, 16'd58539, 16'd7651, 16'd47701, 16'd39727, 16'd34767, 16'd34881, 16'd33592, 16'd21389, 16'd46649, 16'd61444});
	test_expansion(128'h1e6a8b423a48d544838b94412a83a78e, {16'd26612, 16'd53868, 16'd44093, 16'd6317, 16'd28651, 16'd59065, 16'd42081, 16'd22438, 16'd2367, 16'd31133, 16'd42859, 16'd64962, 16'd57825, 16'd35341, 16'd48403, 16'd37904, 16'd39987, 16'd58118, 16'd20121, 16'd12311, 16'd38652, 16'd12625, 16'd2232, 16'd56506, 16'd4408, 16'd58226});
	test_expansion(128'hb0df13dade59fad8081547e406b4efeb, {16'd30837, 16'd47337, 16'd57571, 16'd29433, 16'd51913, 16'd20958, 16'd25259, 16'd44965, 16'd9042, 16'd41582, 16'd6016, 16'd40601, 16'd63011, 16'd17826, 16'd22393, 16'd36009, 16'd4834, 16'd47103, 16'd30226, 16'd36205, 16'd30638, 16'd18103, 16'd45549, 16'd10890, 16'd60898, 16'd10050});
	test_expansion(128'h48bdcc158463e922270c8a47b89afbf0, {16'd38203, 16'd10488, 16'd46162, 16'd39971, 16'd6526, 16'd59545, 16'd18193, 16'd56791, 16'd18475, 16'd24291, 16'd388, 16'd19002, 16'd49488, 16'd13873, 16'd10563, 16'd30758, 16'd56987, 16'd30291, 16'd45958, 16'd15012, 16'd37669, 16'd35914, 16'd37709, 16'd42341, 16'd51899, 16'd48820});
	test_expansion(128'h8d6400672c8827d28462635c4ad8bda2, {16'd37651, 16'd19426, 16'd12172, 16'd56927, 16'd9827, 16'd20292, 16'd43310, 16'd31703, 16'd6500, 16'd4072, 16'd7341, 16'd50914, 16'd46237, 16'd53111, 16'd33635, 16'd20383, 16'd24424, 16'd24001, 16'd28684, 16'd13929, 16'd28323, 16'd30812, 16'd47612, 16'd23886, 16'd32822, 16'd3402});
	test_expansion(128'h6da7ce2efb887d27fec3d04e629152c1, {16'd9028, 16'd55141, 16'd49539, 16'd27576, 16'd50100, 16'd33863, 16'd36035, 16'd42165, 16'd20454, 16'd61500, 16'd20010, 16'd17050, 16'd17724, 16'd45202, 16'd45870, 16'd37170, 16'd42952, 16'd31789, 16'd43616, 16'd40696, 16'd43506, 16'd56227, 16'd1912, 16'd56557, 16'd31540, 16'd48007});
	test_expansion(128'h964f8ead55b71f807f43c20de1f74e3f, {16'd44933, 16'd5810, 16'd22988, 16'd12707, 16'd9783, 16'd53010, 16'd40579, 16'd20883, 16'd14304, 16'd40022, 16'd7262, 16'd9459, 16'd22287, 16'd36039, 16'd44997, 16'd48751, 16'd56024, 16'd23446, 16'd62800, 16'd34377, 16'd23385, 16'd16856, 16'd63512, 16'd47324, 16'd14112, 16'd37855});
	test_expansion(128'hbeafa2779f3d3b60035cf74bfca1b730, {16'd11019, 16'd12121, 16'd64636, 16'd46586, 16'd57518, 16'd15321, 16'd64060, 16'd42856, 16'd48121, 16'd42655, 16'd32346, 16'd11013, 16'd42930, 16'd12859, 16'd51514, 16'd53422, 16'd30279, 16'd4637, 16'd21369, 16'd43173, 16'd18980, 16'd54922, 16'd31318, 16'd36765, 16'd25146, 16'd39233});
	test_expansion(128'hf76b81fa247489ae8f1e3ae4c394a59d, {16'd27120, 16'd51687, 16'd49743, 16'd63550, 16'd49803, 16'd59716, 16'd19739, 16'd26095, 16'd28511, 16'd46372, 16'd22412, 16'd11563, 16'd32053, 16'd17056, 16'd43129, 16'd64585, 16'd65296, 16'd41833, 16'd59285, 16'd10476, 16'd35603, 16'd14700, 16'd253, 16'd36664, 16'd19086, 16'd45157});
	test_expansion(128'h86318d73609a87ceaa39555c98251426, {16'd3425, 16'd17744, 16'd44570, 16'd56359, 16'd7969, 16'd37205, 16'd44286, 16'd57978, 16'd21035, 16'd31516, 16'd25296, 16'd8096, 16'd7131, 16'd7546, 16'd9564, 16'd14096, 16'd46698, 16'd37736, 16'd14518, 16'd57024, 16'd23737, 16'd23349, 16'd35671, 16'd41970, 16'd14940, 16'd50858});
	test_expansion(128'he0dfb8720ca460af7f45c3af60afcd88, {16'd50549, 16'd22534, 16'd4259, 16'd25908, 16'd59615, 16'd55435, 16'd17421, 16'd40765, 16'd38920, 16'd44498, 16'd55874, 16'd55554, 16'd43622, 16'd15245, 16'd16208, 16'd60067, 16'd33427, 16'd4515, 16'd12872, 16'd18700, 16'd54421, 16'd65166, 16'd55714, 16'd55716, 16'd3833, 16'd33250});
	test_expansion(128'h3aa85c894711e290e8dfa77b141dd5c4, {16'd19655, 16'd6087, 16'd23298, 16'd23859, 16'd11442, 16'd56894, 16'd36937, 16'd58743, 16'd51069, 16'd56618, 16'd25380, 16'd36186, 16'd55196, 16'd47797, 16'd60482, 16'd10184, 16'd16756, 16'd54102, 16'd19406, 16'd53018, 16'd34429, 16'd23561, 16'd56828, 16'd36972, 16'd16736, 16'd45167});
	test_expansion(128'h14434426cdc2337ff71f914a6a8eae26, {16'd62273, 16'd56086, 16'd42464, 16'd6780, 16'd34838, 16'd54167, 16'd61279, 16'd57109, 16'd28196, 16'd38976, 16'd51348, 16'd2369, 16'd12010, 16'd2896, 16'd47673, 16'd62018, 16'd27475, 16'd49727, 16'd58686, 16'd48226, 16'd35331, 16'd3519, 16'd40201, 16'd37985, 16'd23863, 16'd11296});
	test_expansion(128'hf7fe487928a626618d9cbcaeeff864fb, {16'd3958, 16'd50263, 16'd15372, 16'd62148, 16'd24869, 16'd13904, 16'd57824, 16'd42892, 16'd56533, 16'd25083, 16'd58616, 16'd40781, 16'd16258, 16'd3719, 16'd5161, 16'd53582, 16'd25180, 16'd35989, 16'd61468, 16'd19020, 16'd11452, 16'd23060, 16'd45263, 16'd37166, 16'd26512, 16'd14011});
	test_expansion(128'hd95b37a4200b057433c469710825990e, {16'd18982, 16'd50350, 16'd31752, 16'd62455, 16'd55103, 16'd41346, 16'd18205, 16'd61711, 16'd22119, 16'd49055, 16'd15096, 16'd37819, 16'd36203, 16'd65111, 16'd10735, 16'd9860, 16'd47855, 16'd31976, 16'd23995, 16'd22601, 16'd21556, 16'd44622, 16'd24934, 16'd47172, 16'd26431, 16'd16362});
	test_expansion(128'h3034bfeee12df14e8187ec51728f3aa8, {16'd3048, 16'd8420, 16'd8576, 16'd4620, 16'd45016, 16'd60060, 16'd52121, 16'd9953, 16'd63351, 16'd56194, 16'd32191, 16'd18449, 16'd38353, 16'd12502, 16'd670, 16'd29101, 16'd50386, 16'd54887, 16'd18669, 16'd57798, 16'd53128, 16'd43078, 16'd63215, 16'd50114, 16'd10612, 16'd65444});
	test_expansion(128'h7ed6cd51df8ce4abf55e2da2289b3298, {16'd8495, 16'd8562, 16'd51567, 16'd10412, 16'd36571, 16'd17789, 16'd4458, 16'd4414, 16'd64255, 16'd52873, 16'd12739, 16'd34477, 16'd35179, 16'd29965, 16'd27399, 16'd52458, 16'd45823, 16'd11993, 16'd61461, 16'd33162, 16'd1955, 16'd25003, 16'd25662, 16'd65126, 16'd60688, 16'd7171});
	test_expansion(128'heb071dff1ebe2b7336733dd264c3e9b4, {16'd24460, 16'd14558, 16'd20741, 16'd63736, 16'd7596, 16'd17080, 16'd39661, 16'd15778, 16'd18406, 16'd6413, 16'd28609, 16'd17660, 16'd37541, 16'd40245, 16'd58417, 16'd2871, 16'd31061, 16'd29714, 16'd37765, 16'd48685, 16'd13203, 16'd38400, 16'd25807, 16'd64534, 16'd59654, 16'd32670});
	test_expansion(128'h2f23a71a721d4e5baa041eaa7d9e051e, {16'd565, 16'd19293, 16'd32997, 16'd36501, 16'd60261, 16'd38782, 16'd12409, 16'd1399, 16'd19803, 16'd14911, 16'd12743, 16'd19702, 16'd36035, 16'd45162, 16'd14176, 16'd38349, 16'd18249, 16'd48800, 16'd63783, 16'd590, 16'd9262, 16'd63547, 16'd56798, 16'd44547, 16'd13720, 16'd16039});
	test_expansion(128'h013df7fd710ef980610270d12ee9eb97, {16'd39857, 16'd40753, 16'd52937, 16'd53453, 16'd51971, 16'd9826, 16'd55590, 16'd25894, 16'd8320, 16'd23531, 16'd62987, 16'd6485, 16'd48460, 16'd34361, 16'd60763, 16'd16693, 16'd47782, 16'd28205, 16'd771, 16'd53888, 16'd63038, 16'd64747, 16'd51240, 16'd9903, 16'd5703, 16'd56488});
	test_expansion(128'h3ba08bdaf3905592dced0e9f6a7a5705, {16'd44025, 16'd41007, 16'd22389, 16'd29199, 16'd2156, 16'd55343, 16'd51210, 16'd61031, 16'd58039, 16'd57489, 16'd27303, 16'd49305, 16'd1365, 16'd17139, 16'd42929, 16'd52419, 16'd56909, 16'd22651, 16'd12287, 16'd1627, 16'd28149, 16'd46991, 16'd33398, 16'd41567, 16'd22460, 16'd5845});
	test_expansion(128'hc330e168dee072f13970208560040942, {16'd39481, 16'd60196, 16'd1076, 16'd13875, 16'd10286, 16'd48086, 16'd43522, 16'd18105, 16'd9792, 16'd2789, 16'd37325, 16'd23860, 16'd30821, 16'd55262, 16'd29504, 16'd46404, 16'd11007, 16'd7491, 16'd17317, 16'd2744, 16'd63713, 16'd1048, 16'd7628, 16'd31005, 16'd47371, 16'd48023});
	test_expansion(128'h60a537081d101af3e9e2c4a82de2dc87, {16'd28054, 16'd19746, 16'd11950, 16'd25631, 16'd30310, 16'd14814, 16'd58852, 16'd12883, 16'd48712, 16'd41521, 16'd42935, 16'd54759, 16'd59931, 16'd4880, 16'd53388, 16'd50535, 16'd15982, 16'd24675, 16'd11459, 16'd27593, 16'd50850, 16'd33733, 16'd55989, 16'd39934, 16'd29800, 16'd50434});
	test_expansion(128'hfd80ff390a42714e236dba55a2841aab, {16'd58441, 16'd44008, 16'd53583, 16'd59842, 16'd23303, 16'd32811, 16'd32904, 16'd28428, 16'd65430, 16'd40023, 16'd52913, 16'd47789, 16'd15900, 16'd34018, 16'd29197, 16'd52958, 16'd50663, 16'd29051, 16'd48123, 16'd8291, 16'd57545, 16'd61191, 16'd60183, 16'd35563, 16'd33845, 16'd13620});
	test_expansion(128'h948d28e6b82c1d6827494aba44b95b15, {16'd1008, 16'd50034, 16'd29875, 16'd5366, 16'd49064, 16'd28537, 16'd64589, 16'd8457, 16'd16872, 16'd32640, 16'd22457, 16'd29114, 16'd17204, 16'd2732, 16'd18968, 16'd9272, 16'd25554, 16'd36392, 16'd28790, 16'd54029, 16'd63185, 16'd17879, 16'd64212, 16'd2092, 16'd8354, 16'd37879});
	test_expansion(128'h822fac97e896d0a5913967b41721317a, {16'd4582, 16'd40896, 16'd17045, 16'd61493, 16'd14430, 16'd47197, 16'd59962, 16'd46980, 16'd17227, 16'd29100, 16'd3498, 16'd60881, 16'd20997, 16'd34003, 16'd13005, 16'd7151, 16'd23952, 16'd6048, 16'd34618, 16'd9595, 16'd16196, 16'd5077, 16'd15778, 16'd5771, 16'd28244, 16'd9611});
	test_expansion(128'h04b5d3dab7e25ced952a0d13d337e77d, {16'd20922, 16'd64579, 16'd26288, 16'd24264, 16'd16104, 16'd63789, 16'd12568, 16'd16586, 16'd52231, 16'd42312, 16'd39367, 16'd50092, 16'd18500, 16'd33368, 16'd42231, 16'd42690, 16'd43094, 16'd33413, 16'd43707, 16'd26744, 16'd4219, 16'd39856, 16'd63380, 16'd1757, 16'd3989, 16'd2748});
	test_expansion(128'h5d6ce9bbda04ac866cb0a537baca3f40, {16'd7349, 16'd59513, 16'd17365, 16'd53499, 16'd33142, 16'd25039, 16'd5501, 16'd48044, 16'd26838, 16'd60608, 16'd24681, 16'd57979, 16'd8848, 16'd35352, 16'd60989, 16'd30174, 16'd61591, 16'd34709, 16'd25009, 16'd12400, 16'd4579, 16'd59503, 16'd31372, 16'd4929, 16'd3677, 16'd39731});
	test_expansion(128'h25c1e24be2f4d919f5b8a27477aabbe1, {16'd39183, 16'd34768, 16'd41302, 16'd61497, 16'd51256, 16'd15172, 16'd7340, 16'd52314, 16'd29687, 16'd58441, 16'd18076, 16'd49384, 16'd61067, 16'd48265, 16'd61291, 16'd47946, 16'd10181, 16'd19163, 16'd41895, 16'd34689, 16'd24693, 16'd52609, 16'd43933, 16'd7969, 16'd59548, 16'd63508});
	test_expansion(128'hb9506665db144fc130b7e52579edbe65, {16'd44890, 16'd26432, 16'd58530, 16'd2711, 16'd13717, 16'd44498, 16'd15450, 16'd31966, 16'd8064, 16'd36790, 16'd62017, 16'd63164, 16'd5059, 16'd30135, 16'd4938, 16'd46203, 16'd3350, 16'd1362, 16'd45724, 16'd952, 16'd46253, 16'd19784, 16'd16659, 16'd54602, 16'd24275, 16'd11549});
	test_expansion(128'h3b63187ac70cd493ef5785dcb144e628, {16'd15301, 16'd64734, 16'd16812, 16'd50661, 16'd13389, 16'd61989, 16'd36658, 16'd2247, 16'd12293, 16'd30590, 16'd33947, 16'd5058, 16'd3525, 16'd35177, 16'd41095, 16'd14921, 16'd5032, 16'd20539, 16'd286, 16'd42574, 16'd14401, 16'd42002, 16'd49016, 16'd18066, 16'd35063, 16'd50820});
	test_expansion(128'he2d781f2d9a8e54765d3642556e9fad3, {16'd13249, 16'd49709, 16'd17045, 16'd56613, 16'd49914, 16'd45681, 16'd47752, 16'd59401, 16'd1462, 16'd6236, 16'd4956, 16'd40579, 16'd23027, 16'd42506, 16'd31385, 16'd23943, 16'd48319, 16'd20019, 16'd63159, 16'd35418, 16'd38677, 16'd44437, 16'd2011, 16'd25517, 16'd43705, 16'd31199});
	test_expansion(128'h5e08d1b4d786313b992846bee0864226, {16'd2065, 16'd29439, 16'd43142, 16'd30707, 16'd9001, 16'd16241, 16'd50075, 16'd57158, 16'd4115, 16'd34521, 16'd12620, 16'd5351, 16'd11883, 16'd9245, 16'd18747, 16'd46140, 16'd18660, 16'd52639, 16'd59056, 16'd60219, 16'd56247, 16'd53718, 16'd37375, 16'd54284, 16'd18120, 16'd1380});
	test_expansion(128'h61ef2ddc4b93c3092ebafd2e7ee365e7, {16'd43086, 16'd22215, 16'd56740, 16'd17390, 16'd18895, 16'd17335, 16'd11581, 16'd20944, 16'd36952, 16'd39477, 16'd41649, 16'd65268, 16'd43172, 16'd63653, 16'd30402, 16'd52488, 16'd61402, 16'd10195, 16'd55838, 16'd50820, 16'd46791, 16'd22117, 16'd33147, 16'd1765, 16'd57914, 16'd16003});
	test_expansion(128'h0bd738526c554603e6891eef5e59e8b5, {16'd51584, 16'd34309, 16'd19008, 16'd28127, 16'd11708, 16'd40355, 16'd25292, 16'd59364, 16'd10569, 16'd59940, 16'd49105, 16'd6246, 16'd40767, 16'd48243, 16'd46817, 16'd26818, 16'd16319, 16'd15580, 16'd34688, 16'd35906, 16'd30588, 16'd49801, 16'd36068, 16'd26102, 16'd12260, 16'd49032});
	test_expansion(128'h31c578909c04e8f7a2780c8942f920b7, {16'd53392, 16'd6929, 16'd44927, 16'd14149, 16'd8361, 16'd18769, 16'd4332, 16'd3917, 16'd32688, 16'd35590, 16'd43113, 16'd21383, 16'd55050, 16'd43632, 16'd32525, 16'd39297, 16'd13628, 16'd30021, 16'd22071, 16'd25691, 16'd55628, 16'd4733, 16'd37951, 16'd48898, 16'd35499, 16'd17448});
	test_expansion(128'h795f041567f0688b746c14d498790246, {16'd49995, 16'd60125, 16'd42208, 16'd38259, 16'd57151, 16'd28756, 16'd28846, 16'd4850, 16'd20472, 16'd3506, 16'd1533, 16'd40855, 16'd44900, 16'd59422, 16'd53241, 16'd55526, 16'd21039, 16'd28917, 16'd37069, 16'd60065, 16'd42617, 16'd59553, 16'd11172, 16'd33059, 16'd55582, 16'd43470});
	test_expansion(128'hc608f0e2d50505baec59197f8e93043a, {16'd39609, 16'd36277, 16'd61615, 16'd12645, 16'd10146, 16'd11062, 16'd13681, 16'd6294, 16'd45146, 16'd50429, 16'd13829, 16'd60451, 16'd17319, 16'd11233, 16'd19857, 16'd58665, 16'd12981, 16'd62223, 16'd33496, 16'd58511, 16'd55811, 16'd9401, 16'd45666, 16'd22178, 16'd52600, 16'd27690});
	test_expansion(128'h3ce42dac584f0f847865d0f71d26dbe2, {16'd32032, 16'd54465, 16'd41364, 16'd19225, 16'd50478, 16'd37899, 16'd56819, 16'd64681, 16'd27274, 16'd7360, 16'd43272, 16'd31150, 16'd32539, 16'd26912, 16'd25400, 16'd51110, 16'd39557, 16'd22962, 16'd23333, 16'd15354, 16'd11269, 16'd9520, 16'd39662, 16'd65090, 16'd20638, 16'd14978});
	test_expansion(128'hbf4d969a50e678369aced8f141c5c803, {16'd13335, 16'd62412, 16'd11485, 16'd42857, 16'd41007, 16'd33066, 16'd34484, 16'd50809, 16'd16723, 16'd55702, 16'd18600, 16'd3481, 16'd31930, 16'd41760, 16'd46036, 16'd17398, 16'd53684, 16'd8273, 16'd56823, 16'd32093, 16'd30205, 16'd24070, 16'd25721, 16'd37469, 16'd50938, 16'd15785});
	test_expansion(128'h5959c4b8e6334794bb9580307057c819, {16'd18398, 16'd8653, 16'd13628, 16'd32195, 16'd12985, 16'd30705, 16'd20413, 16'd28337, 16'd56063, 16'd56004, 16'd256, 16'd59871, 16'd15413, 16'd21746, 16'd27319, 16'd29782, 16'd16076, 16'd48977, 16'd53561, 16'd27856, 16'd22238, 16'd3548, 16'd60087, 16'd7554, 16'd21197, 16'd44643});
	test_expansion(128'h2c3e6ed53f78895c0e25bc6cbbee0300, {16'd54143, 16'd3816, 16'd5166, 16'd49310, 16'd60914, 16'd52424, 16'd27548, 16'd33635, 16'd44382, 16'd15028, 16'd26724, 16'd28831, 16'd54861, 16'd45506, 16'd8057, 16'd23136, 16'd19149, 16'd18910, 16'd15584, 16'd63202, 16'd46031, 16'd52639, 16'd31204, 16'd40412, 16'd45992, 16'd62195});
	test_expansion(128'h45b1c9af5e005bb8303f9fcea318ef80, {16'd64681, 16'd45098, 16'd36948, 16'd48555, 16'd41923, 16'd42583, 16'd26964, 16'd45104, 16'd13046, 16'd56499, 16'd28040, 16'd6464, 16'd11077, 16'd19264, 16'd57857, 16'd19415, 16'd37273, 16'd53908, 16'd36787, 16'd18647, 16'd29756, 16'd3662, 16'd60412, 16'd32335, 16'd6524, 16'd30148});
	test_expansion(128'h325a607e78301c60efd90fedfa5e0c67, {16'd48756, 16'd8893, 16'd7635, 16'd27137, 16'd59337, 16'd31014, 16'd56972, 16'd2458, 16'd16901, 16'd14440, 16'd50918, 16'd37254, 16'd58723, 16'd13049, 16'd48708, 16'd55082, 16'd38518, 16'd4038, 16'd51267, 16'd53492, 16'd45397, 16'd64543, 16'd3101, 16'd20316, 16'd27487, 16'd57294});
	test_expansion(128'h8142f2d189beeafc9ff34037b983b095, {16'd52386, 16'd24783, 16'd60681, 16'd33661, 16'd12112, 16'd10807, 16'd54480, 16'd8849, 16'd22514, 16'd30008, 16'd14581, 16'd14335, 16'd22699, 16'd30992, 16'd24043, 16'd61062, 16'd13722, 16'd5629, 16'd20619, 16'd29600, 16'd1846, 16'd63539, 16'd28473, 16'd18644, 16'd46589, 16'd52970});
	test_expansion(128'h3af9b7efe2e0d78613fa7ec7470321c0, {16'd62301, 16'd2825, 16'd18375, 16'd15841, 16'd63759, 16'd41531, 16'd450, 16'd62541, 16'd53378, 16'd41362, 16'd18557, 16'd6552, 16'd10543, 16'd23384, 16'd8957, 16'd56410, 16'd11926, 16'd63521, 16'd56059, 16'd47425, 16'd7476, 16'd1439, 16'd54297, 16'd49482, 16'd57286, 16'd23736});
	test_expansion(128'h6a1323519536b154b09a49bbcf6dc326, {16'd35984, 16'd51039, 16'd41477, 16'd41888, 16'd39076, 16'd41252, 16'd2781, 16'd12177, 16'd61131, 16'd62577, 16'd34127, 16'd41849, 16'd46324, 16'd46924, 16'd48052, 16'd14677, 16'd24327, 16'd7602, 16'd1754, 16'd4170, 16'd38601, 16'd43931, 16'd40500, 16'd25250, 16'd56299, 16'd56170});
	test_expansion(128'h50eb4bf5742cd0b37b2c367a3370cb4d, {16'd31858, 16'd3426, 16'd1297, 16'd62457, 16'd20243, 16'd16518, 16'd4053, 16'd34126, 16'd7018, 16'd36597, 16'd51192, 16'd9866, 16'd57698, 16'd30107, 16'd49248, 16'd7743, 16'd26089, 16'd58230, 16'd44569, 16'd26525, 16'd11597, 16'd32805, 16'd21742, 16'd5562, 16'd23834, 16'd62809});
	test_expansion(128'h4164bd1fdf4cc7842f4fdb5d402627d8, {16'd31339, 16'd13222, 16'd58046, 16'd760, 16'd61430, 16'd48959, 16'd30267, 16'd38863, 16'd37926, 16'd22959, 16'd52434, 16'd20770, 16'd2449, 16'd50038, 16'd50867, 16'd46138, 16'd19449, 16'd5503, 16'd5123, 16'd15421, 16'd9761, 16'd42727, 16'd30440, 16'd38341, 16'd23810, 16'd11775});
	test_expansion(128'hd71ea548f5827c8bea2fb1884970b484, {16'd21917, 16'd36594, 16'd38928, 16'd4881, 16'd57313, 16'd48517, 16'd62931, 16'd44923, 16'd50320, 16'd53595, 16'd4258, 16'd6691, 16'd32353, 16'd20684, 16'd30819, 16'd63232, 16'd32582, 16'd2090, 16'd46979, 16'd64714, 16'd10729, 16'd14715, 16'd34605, 16'd57174, 16'd56682, 16'd46158});
	test_expansion(128'he379d6493a84856cf8f6d82c5df6c59f, {16'd46683, 16'd22828, 16'd14255, 16'd7162, 16'd51706, 16'd28976, 16'd29291, 16'd18671, 16'd56941, 16'd17071, 16'd58286, 16'd10733, 16'd18353, 16'd22075, 16'd56380, 16'd46033, 16'd23187, 16'd45997, 16'd57157, 16'd12741, 16'd15573, 16'd49674, 16'd7286, 16'd28483, 16'd51426, 16'd24823});
	test_expansion(128'hc409109db0611082381be6c0e8fb21cd, {16'd6554, 16'd36064, 16'd14460, 16'd62297, 16'd8223, 16'd31546, 16'd20217, 16'd18897, 16'd11801, 16'd9123, 16'd46617, 16'd15804, 16'd14953, 16'd48783, 16'd5627, 16'd63559, 16'd53477, 16'd3540, 16'd42557, 16'd38414, 16'd30617, 16'd57035, 16'd41243, 16'd41055, 16'd60388, 16'd33657});
	test_expansion(128'h2e7723d02653d5bb2d42023f66e4d49c, {16'd64206, 16'd16211, 16'd11168, 16'd23734, 16'd3293, 16'd54777, 16'd19790, 16'd59229, 16'd42046, 16'd26702, 16'd57142, 16'd49257, 16'd52697, 16'd57798, 16'd27621, 16'd14772, 16'd23957, 16'd44005, 16'd63069, 16'd61234, 16'd48755, 16'd61650, 16'd10507, 16'd63742, 16'd63196, 16'd40461});
	test_expansion(128'h77fe9149efb5028474f0fbc81dd78b01, {16'd28776, 16'd30337, 16'd4529, 16'd65234, 16'd59202, 16'd3104, 16'd60758, 16'd53786, 16'd45374, 16'd51508, 16'd6671, 16'd20059, 16'd22990, 16'd40830, 16'd4254, 16'd23831, 16'd38825, 16'd40246, 16'd64835, 16'd23942, 16'd58802, 16'd57044, 16'd8580, 16'd52265, 16'd64770, 16'd20899});
	test_expansion(128'h910f786918bbb9233228e30bab9cd685, {16'd17594, 16'd31193, 16'd13230, 16'd6005, 16'd9792, 16'd17664, 16'd20887, 16'd64963, 16'd23, 16'd6891, 16'd19065, 16'd10155, 16'd40059, 16'd53183, 16'd47104, 16'd49895, 16'd61562, 16'd46539, 16'd27189, 16'd16068, 16'd13374, 16'd11759, 16'd26857, 16'd12861, 16'd48289, 16'd38059});
	test_expansion(128'h8a0cb56e706de5adf1c657b3b863d5a8, {16'd62640, 16'd27108, 16'd26375, 16'd49353, 16'd38437, 16'd20985, 16'd23946, 16'd18262, 16'd22196, 16'd42408, 16'd16912, 16'd6806, 16'd20291, 16'd7144, 16'd57753, 16'd3368, 16'd37909, 16'd6809, 16'd51038, 16'd15714, 16'd45614, 16'd55110, 16'd10510, 16'd22511, 16'd45226, 16'd54434});
	test_expansion(128'hf46b1aac6a48d9d0ffc523a211082c1e, {16'd9592, 16'd4328, 16'd23712, 16'd14613, 16'd4587, 16'd63070, 16'd27766, 16'd64341, 16'd42591, 16'd43651, 16'd44876, 16'd24642, 16'd62047, 16'd20135, 16'd34176, 16'd58638, 16'd24878, 16'd18078, 16'd28337, 16'd12705, 16'd731, 16'd22027, 16'd47789, 16'd19862, 16'd22568, 16'd37251});
	test_expansion(128'hb455098c86aa591aafcfd61a594548c5, {16'd55946, 16'd42373, 16'd18575, 16'd7975, 16'd30150, 16'd51666, 16'd14486, 16'd47549, 16'd32192, 16'd59457, 16'd30190, 16'd10852, 16'd3557, 16'd3644, 16'd63585, 16'd56341, 16'd7645, 16'd31528, 16'd28435, 16'd2108, 16'd55906, 16'd57746, 16'd10009, 16'd11956, 16'd47268, 16'd4709});
	test_expansion(128'h1935f61048aedc02d82b488080d982f4, {16'd4857, 16'd13680, 16'd43220, 16'd47893, 16'd15037, 16'd51528, 16'd1332, 16'd16224, 16'd55516, 16'd6102, 16'd16713, 16'd52789, 16'd6616, 16'd45987, 16'd33803, 16'd11781, 16'd3631, 16'd7901, 16'd19396, 16'd62788, 16'd53400, 16'd37512, 16'd662, 16'd41433, 16'd21767, 16'd25005});
	test_expansion(128'h547253c5d1344aa14622321ca5517b36, {16'd43557, 16'd33711, 16'd14442, 16'd52046, 16'd18927, 16'd21820, 16'd17012, 16'd53972, 16'd31717, 16'd12640, 16'd16191, 16'd26727, 16'd64740, 16'd36993, 16'd40516, 16'd36460, 16'd25638, 16'd50201, 16'd62427, 16'd46098, 16'd8876, 16'd14663, 16'd58345, 16'd16370, 16'd56608, 16'd31375});
	test_expansion(128'h5395d7138f907860ef99181816aad76f, {16'd65199, 16'd19079, 16'd48474, 16'd59136, 16'd48799, 16'd52476, 16'd53567, 16'd27018, 16'd19819, 16'd3940, 16'd21867, 16'd6050, 16'd58204, 16'd61973, 16'd9187, 16'd59012, 16'd51638, 16'd10431, 16'd18038, 16'd47958, 16'd37784, 16'd49107, 16'd17894, 16'd37847, 16'd61813, 16'd36256});
	test_expansion(128'h893d47b03ba810f558ac0efdddb99554, {16'd21606, 16'd49641, 16'd54268, 16'd8386, 16'd22355, 16'd29923, 16'd10422, 16'd39195, 16'd28612, 16'd21083, 16'd41097, 16'd56432, 16'd18359, 16'd8808, 16'd24365, 16'd54726, 16'd32355, 16'd22522, 16'd28137, 16'd17971, 16'd15582, 16'd3404, 16'd33988, 16'd17574, 16'd11820, 16'd5511});
	test_expansion(128'hb9398c2e5a772fb81bc50d24f0d41337, {16'd21239, 16'd39159, 16'd33700, 16'd11465, 16'd35831, 16'd46940, 16'd12604, 16'd53528, 16'd36732, 16'd61775, 16'd56552, 16'd34878, 16'd24758, 16'd59299, 16'd4634, 16'd2212, 16'd61524, 16'd36187, 16'd13107, 16'd12373, 16'd1339, 16'd34279, 16'd15714, 16'd20993, 16'd45511, 16'd41042});
	test_expansion(128'h49a5a429996318251e3b795b3f494c7f, {16'd8714, 16'd37405, 16'd14676, 16'd39690, 16'd13614, 16'd62095, 16'd41022, 16'd6849, 16'd12633, 16'd29148, 16'd31179, 16'd1968, 16'd10940, 16'd61614, 16'd16933, 16'd16325, 16'd21045, 16'd64418, 16'd28103, 16'd52978, 16'd11084, 16'd28229, 16'd41467, 16'd63612, 16'd37770, 16'd41160});
	test_expansion(128'h97d239622fbe5d899dde43422cb08470, {16'd44659, 16'd32158, 16'd49180, 16'd50594, 16'd3467, 16'd9427, 16'd50590, 16'd8720, 16'd63019, 16'd42033, 16'd2178, 16'd63121, 16'd57026, 16'd61352, 16'd40997, 16'd33526, 16'd9341, 16'd3119, 16'd11936, 16'd19686, 16'd44390, 16'd29169, 16'd19707, 16'd63955, 16'd20167, 16'd17005});
	test_expansion(128'h04bab2c5af45c765a976d052b65f38c7, {16'd39429, 16'd3750, 16'd53769, 16'd9001, 16'd5290, 16'd8797, 16'd53739, 16'd21920, 16'd1567, 16'd38081, 16'd41297, 16'd60665, 16'd33993, 16'd57047, 16'd59913, 16'd62651, 16'd3591, 16'd45372, 16'd10370, 16'd58953, 16'd739, 16'd34483, 16'd13703, 16'd10456, 16'd52185, 16'd38858});
	test_expansion(128'hb3bec002fb948761d2f6a0a34ff60f52, {16'd23116, 16'd61132, 16'd30857, 16'd26810, 16'd56302, 16'd26220, 16'd27156, 16'd27023, 16'd27875, 16'd57244, 16'd43583, 16'd60272, 16'd10145, 16'd11227, 16'd3330, 16'd15525, 16'd25603, 16'd61100, 16'd57215, 16'd50228, 16'd16413, 16'd48111, 16'd41775, 16'd22654, 16'd9179, 16'd9910});
	test_expansion(128'hd08b28cbd739dcc39e808faab137990f, {16'd37105, 16'd55086, 16'd45996, 16'd14822, 16'd4154, 16'd62259, 16'd58521, 16'd54034, 16'd36090, 16'd59746, 16'd502, 16'd43986, 16'd18940, 16'd28008, 16'd19334, 16'd62340, 16'd11141, 16'd31818, 16'd21766, 16'd17920, 16'd48279, 16'd48257, 16'd30123, 16'd44117, 16'd35543, 16'd24065});
	test_expansion(128'h5b8e55e5c80642370024021502909455, {16'd16324, 16'd5409, 16'd13720, 16'd55137, 16'd59678, 16'd19021, 16'd7437, 16'd23814, 16'd6467, 16'd846, 16'd34444, 16'd28367, 16'd25302, 16'd13873, 16'd40450, 16'd59545, 16'd50880, 16'd47458, 16'd60614, 16'd50100, 16'd28691, 16'd19432, 16'd60487, 16'd16127, 16'd9909, 16'd14716});
	test_expansion(128'h023151cbff8694ede62eec12cce7875a, {16'd16119, 16'd37229, 16'd32210, 16'd31388, 16'd50543, 16'd65280, 16'd12404, 16'd44102, 16'd7685, 16'd18229, 16'd16570, 16'd19632, 16'd64954, 16'd8221, 16'd4200, 16'd52201, 16'd3184, 16'd18919, 16'd912, 16'd52234, 16'd65099, 16'd13094, 16'd2872, 16'd39620, 16'd12335, 16'd758});
	test_expansion(128'h5c174d094b4bf74b964959e1139f6b66, {16'd22696, 16'd55914, 16'd46979, 16'd23824, 16'd9053, 16'd45905, 16'd27812, 16'd7549, 16'd11435, 16'd3168, 16'd48880, 16'd41422, 16'd24776, 16'd41993, 16'd21322, 16'd31752, 16'd59405, 16'd64728, 16'd32240, 16'd32145, 16'd52972, 16'd46344, 16'd32541, 16'd57464, 16'd13012, 16'd65057});
	test_expansion(128'ha71713405c524874142ce68a7586d401, {16'd32560, 16'd19678, 16'd61278, 16'd19406, 16'd22839, 16'd15945, 16'd57988, 16'd55881, 16'd47436, 16'd44207, 16'd33042, 16'd4928, 16'd35630, 16'd26896, 16'd42469, 16'd3536, 16'd4583, 16'd44244, 16'd38341, 16'd173, 16'd64201, 16'd45520, 16'd43883, 16'd26555, 16'd15099, 16'd26846});
	test_expansion(128'he84ff2377aafaf473d6ef52f971ef651, {16'd56680, 16'd47605, 16'd11230, 16'd9554, 16'd23307, 16'd20940, 16'd44017, 16'd59633, 16'd4314, 16'd34710, 16'd6051, 16'd1280, 16'd42704, 16'd38740, 16'd36223, 16'd54739, 16'd17709, 16'd15170, 16'd27970, 16'd44055, 16'd20667, 16'd839, 16'd57960, 16'd55687, 16'd63091, 16'd6971});
	test_expansion(128'h3adf56db34bdf3ac9402f9e0cf05d9ff, {16'd39721, 16'd11291, 16'd10479, 16'd14737, 16'd31464, 16'd38888, 16'd14339, 16'd57222, 16'd35296, 16'd39305, 16'd47431, 16'd30071, 16'd53780, 16'd5391, 16'd60473, 16'd30506, 16'd26619, 16'd24934, 16'd55594, 16'd54966, 16'd55479, 16'd48296, 16'd25328, 16'd55303, 16'd9633, 16'd1466});
	test_expansion(128'h9f34648bb27c9b12e35a9c7fffdbc05e, {16'd64751, 16'd63854, 16'd56509, 16'd57686, 16'd14210, 16'd14055, 16'd3746, 16'd57064, 16'd1613, 16'd23980, 16'd28453, 16'd7358, 16'd756, 16'd40541, 16'd20652, 16'd22758, 16'd4381, 16'd64670, 16'd11459, 16'd30568, 16'd10403, 16'd5505, 16'd15669, 16'd33192, 16'd52066, 16'd28836});
	test_expansion(128'ha5a8ff3f42b4ca833bb4a92b703c1bca, {16'd54283, 16'd18820, 16'd29817, 16'd45323, 16'd25090, 16'd36992, 16'd18189, 16'd57082, 16'd62538, 16'd62710, 16'd34384, 16'd19028, 16'd36835, 16'd11665, 16'd49579, 16'd22870, 16'd29215, 16'd6552, 16'd51156, 16'd24953, 16'd3067, 16'd39508, 16'd11180, 16'd55754, 16'd23301, 16'd65364});
	test_expansion(128'h84c34aea343b028977c491eb5e24a1d3, {16'd21329, 16'd22288, 16'd59798, 16'd24491, 16'd36891, 16'd60908, 16'd37823, 16'd29550, 16'd50416, 16'd2474, 16'd11870, 16'd32815, 16'd3496, 16'd32030, 16'd32944, 16'd57572, 16'd33686, 16'd63210, 16'd14229, 16'd7368, 16'd49316, 16'd14120, 16'd63, 16'd22226, 16'd8806, 16'd23897});
	test_expansion(128'h7718b6f42aa09c796c5b215af1c03fd6, {16'd13603, 16'd43950, 16'd64392, 16'd42016, 16'd17921, 16'd29754, 16'd34936, 16'd41303, 16'd40177, 16'd44723, 16'd15183, 16'd42287, 16'd27332, 16'd52510, 16'd20701, 16'd26819, 16'd31430, 16'd44813, 16'd8488, 16'd60625, 16'd5326, 16'd56541, 16'd40717, 16'd29841, 16'd3847, 16'd64920});
	test_expansion(128'h8c53fe65f737533d0f90fd6c5b7cdde7, {16'd51444, 16'd27912, 16'd37602, 16'd15759, 16'd61347, 16'd22902, 16'd3244, 16'd39108, 16'd55106, 16'd8298, 16'd62203, 16'd59801, 16'd61004, 16'd13775, 16'd4944, 16'd42142, 16'd43099, 16'd24398, 16'd63009, 16'd21377, 16'd5593, 16'd31054, 16'd64993, 16'd1945, 16'd35291, 16'd37241});
	test_expansion(128'h262a2f8e2a3689ba035b3362f9ff3175, {16'd2271, 16'd11412, 16'd53039, 16'd21234, 16'd3559, 16'd20556, 16'd54679, 16'd30573, 16'd51353, 16'd11174, 16'd26051, 16'd57081, 16'd53886, 16'd41045, 16'd47750, 16'd25425, 16'd10204, 16'd10029, 16'd33285, 16'd65489, 16'd22953, 16'd52972, 16'd46966, 16'd44948, 16'd11276, 16'd26263});
	test_expansion(128'h4dab2ff17239f9345ef1ae8363aa211d, {16'd59330, 16'd29893, 16'd36412, 16'd33343, 16'd24282, 16'd21904, 16'd24540, 16'd46594, 16'd34580, 16'd257, 16'd42176, 16'd46989, 16'd44411, 16'd62922, 16'd43626, 16'd49824, 16'd33181, 16'd41239, 16'd1777, 16'd64714, 16'd50847, 16'd27009, 16'd49240, 16'd23489, 16'd31518, 16'd16252});
	test_expansion(128'hd6e6a381d9de9ab9938fd89528842c46, {16'd35957, 16'd25522, 16'd34219, 16'd839, 16'd24237, 16'd50399, 16'd31857, 16'd59200, 16'd9768, 16'd31009, 16'd5197, 16'd61980, 16'd28687, 16'd49977, 16'd22309, 16'd4720, 16'd35069, 16'd1606, 16'd37759, 16'd18235, 16'd17370, 16'd63055, 16'd36463, 16'd14071, 16'd12660, 16'd40333});
	test_expansion(128'h6ab0cac4ce504eef2a0b06c7b8f2f791, {16'd2834, 16'd11710, 16'd15033, 16'd20445, 16'd367, 16'd35383, 16'd3682, 16'd40988, 16'd6092, 16'd22999, 16'd8358, 16'd53695, 16'd24017, 16'd9652, 16'd45717, 16'd26191, 16'd59604, 16'd12034, 16'd31849, 16'd64926, 16'd43471, 16'd33439, 16'd8042, 16'd59649, 16'd44768, 16'd55417});
	test_expansion(128'h3a565c5ac540efca6fb0fbd1922aff21, {16'd14659, 16'd18706, 16'd5554, 16'd13853, 16'd52195, 16'd52656, 16'd6082, 16'd29573, 16'd53981, 16'd25752, 16'd13975, 16'd51694, 16'd58295, 16'd22593, 16'd15922, 16'd20439, 16'd44588, 16'd39203, 16'd29624, 16'd12290, 16'd10860, 16'd27732, 16'd55553, 16'd36146, 16'd32610, 16'd38349});
	test_expansion(128'hb185af52f52dd2e5fd61e49e37c78fb5, {16'd62086, 16'd45981, 16'd51177, 16'd34276, 16'd24270, 16'd43065, 16'd21247, 16'd13570, 16'd5430, 16'd61567, 16'd43402, 16'd45688, 16'd57156, 16'd6028, 16'd373, 16'd54521, 16'd7762, 16'd3567, 16'd20794, 16'd33865, 16'd46721, 16'd39989, 16'd35347, 16'd33585, 16'd58098, 16'd60835});
	test_expansion(128'hc50c526454bef2c0e01dc0bece32c069, {16'd21849, 16'd39249, 16'd124, 16'd62272, 16'd57810, 16'd25063, 16'd10042, 16'd19588, 16'd8926, 16'd33830, 16'd13713, 16'd63409, 16'd57338, 16'd12122, 16'd26791, 16'd47246, 16'd41740, 16'd50618, 16'd11021, 16'd49438, 16'd42893, 16'd35388, 16'd5300, 16'd54349, 16'd4109, 16'd65352});
	test_expansion(128'hc096785305a536363fe9041be235ad23, {16'd45239, 16'd93, 16'd20376, 16'd60977, 16'd45558, 16'd36136, 16'd34862, 16'd63218, 16'd17981, 16'd38871, 16'd42329, 16'd54386, 16'd8495, 16'd14464, 16'd648, 16'd36878, 16'd59859, 16'd3553, 16'd51672, 16'd57758, 16'd38502, 16'd35392, 16'd14134, 16'd34567, 16'd51081, 16'd62162});
	test_expansion(128'h18805d5693f88f110e43764c0d745ed7, {16'd35451, 16'd48556, 16'd53255, 16'd14776, 16'd17329, 16'd36826, 16'd15735, 16'd60618, 16'd10523, 16'd21893, 16'd262, 16'd60939, 16'd5382, 16'd10004, 16'd54526, 16'd41670, 16'd688, 16'd1260, 16'd18338, 16'd127, 16'd22814, 16'd18627, 16'd51029, 16'd38309, 16'd27401, 16'd17934});
	test_expansion(128'h611c3396b7357b2c310ddedd5aaee9f0, {16'd25177, 16'd53663, 16'd26248, 16'd58281, 16'd58460, 16'd8406, 16'd30473, 16'd7264, 16'd32901, 16'd48449, 16'd25950, 16'd18829, 16'd64881, 16'd39082, 16'd14197, 16'd53179, 16'd63438, 16'd4807, 16'd56661, 16'd28022, 16'd55658, 16'd51828, 16'd59654, 16'd39168, 16'd47021, 16'd30193});
	test_expansion(128'h41e40718c6be97e664cdc6b9103b4fdc, {16'd11347, 16'd19984, 16'd12258, 16'd8266, 16'd58808, 16'd63882, 16'd9340, 16'd10741, 16'd837, 16'd49276, 16'd40861, 16'd2079, 16'd46191, 16'd46071, 16'd15922, 16'd52152, 16'd26518, 16'd26111, 16'd34502, 16'd52924, 16'd61165, 16'd11007, 16'd62969, 16'd33270, 16'd29281, 16'd22310});
	test_expansion(128'h44f02de62bf960c2d401dc036ba979ab, {16'd6926, 16'd45687, 16'd34924, 16'd43125, 16'd55757, 16'd24885, 16'd47883, 16'd26482, 16'd9537, 16'd4043, 16'd55930, 16'd62336, 16'd32032, 16'd2617, 16'd62581, 16'd45282, 16'd31837, 16'd56529, 16'd59732, 16'd62349, 16'd57878, 16'd32388, 16'd28047, 16'd49287, 16'd42117, 16'd33229});
	test_expansion(128'h9a42af3391e05b1f12004b362759474c, {16'd1293, 16'd4607, 16'd32096, 16'd5681, 16'd23679, 16'd61844, 16'd56978, 16'd49956, 16'd31539, 16'd33757, 16'd52916, 16'd39832, 16'd61551, 16'd36673, 16'd57273, 16'd42365, 16'd55401, 16'd25594, 16'd57673, 16'd63050, 16'd48199, 16'd38127, 16'd33521, 16'd30874, 16'd43299, 16'd46333});
	test_expansion(128'hfedf2ad21702d5498e659aa23b9cc9b3, {16'd58752, 16'd1396, 16'd58669, 16'd52451, 16'd53953, 16'd32732, 16'd30923, 16'd60403, 16'd24702, 16'd16947, 16'd50038, 16'd14918, 16'd11354, 16'd17357, 16'd54335, 16'd12334, 16'd14910, 16'd1902, 16'd17880, 16'd243, 16'd45655, 16'd7588, 16'd63969, 16'd2373, 16'd32684, 16'd2558});
	test_expansion(128'h3398c88a8ea40fff5e7957da0979eced, {16'd5503, 16'd55217, 16'd20180, 16'd47079, 16'd14291, 16'd22814, 16'd13119, 16'd17271, 16'd45950, 16'd187, 16'd13674, 16'd34898, 16'd32358, 16'd57461, 16'd23045, 16'd38583, 16'd36904, 16'd31118, 16'd41987, 16'd25358, 16'd64571, 16'd737, 16'd52814, 16'd22796, 16'd33891, 16'd4373});
	test_expansion(128'h89ac4fe12591554933cfd313c4de0237, {16'd38648, 16'd34494, 16'd62310, 16'd49013, 16'd18099, 16'd21965, 16'd58886, 16'd7554, 16'd37758, 16'd27994, 16'd11698, 16'd61762, 16'd19873, 16'd53379, 16'd7270, 16'd26464, 16'd20375, 16'd15962, 16'd45558, 16'd63288, 16'd20024, 16'd8072, 16'd14008, 16'd453, 16'd11760, 16'd64723});
	test_expansion(128'h3c97769158f387b3111a8255624f55e0, {16'd46065, 16'd58215, 16'd62752, 16'd5360, 16'd35938, 16'd60197, 16'd63279, 16'd17699, 16'd43436, 16'd21650, 16'd21947, 16'd54268, 16'd7953, 16'd61395, 16'd13448, 16'd29954, 16'd3489, 16'd4982, 16'd8213, 16'd47402, 16'd55588, 16'd34111, 16'd50767, 16'd54516, 16'd1672, 16'd18445});
	test_expansion(128'h8226739c882603af77ba5a4896b839e3, {16'd27209, 16'd15941, 16'd58875, 16'd56812, 16'd26394, 16'd338, 16'd41016, 16'd55784, 16'd64084, 16'd61597, 16'd63577, 16'd64177, 16'd8536, 16'd31617, 16'd2448, 16'd60615, 16'd39159, 16'd56507, 16'd21239, 16'd16675, 16'd58111, 16'd49743, 16'd40389, 16'd36435, 16'd18754, 16'd10814});
	test_expansion(128'hf097b1a9f7571be0d10b8e2f40667c88, {16'd52196, 16'd10919, 16'd45274, 16'd53566, 16'd59557, 16'd30000, 16'd14272, 16'd52661, 16'd20682, 16'd42596, 16'd46656, 16'd46904, 16'd43825, 16'd65382, 16'd35972, 16'd52961, 16'd64192, 16'd9990, 16'd39207, 16'd37470, 16'd14095, 16'd33000, 16'd33901, 16'd21815, 16'd55509, 16'd58671});
	test_expansion(128'h3edd2a6f7eba660cdba721ce51ca9e65, {16'd35515, 16'd16889, 16'd22768, 16'd49792, 16'd19093, 16'd30518, 16'd32085, 16'd14667, 16'd45613, 16'd21248, 16'd54609, 16'd43848, 16'd21896, 16'd11522, 16'd40248, 16'd46760, 16'd54802, 16'd37269, 16'd52994, 16'd64292, 16'd42236, 16'd60896, 16'd65187, 16'd37114, 16'd43282, 16'd44134});
	test_expansion(128'h51554de21657ad9d0bf3864ef94d75a7, {16'd60050, 16'd62185, 16'd45712, 16'd17365, 16'd14941, 16'd32239, 16'd5581, 16'd23084, 16'd49157, 16'd32557, 16'd46971, 16'd64101, 16'd52740, 16'd49628, 16'd22102, 16'd53481, 16'd23069, 16'd46617, 16'd51413, 16'd62500, 16'd27257, 16'd49525, 16'd23822, 16'd17194, 16'd35468, 16'd18055});
	test_expansion(128'h4893992d11201c58f38f6cfacb7e474f, {16'd15447, 16'd59208, 16'd43896, 16'd20689, 16'd32826, 16'd60920, 16'd25513, 16'd49888, 16'd34065, 16'd56107, 16'd21634, 16'd49631, 16'd47915, 16'd56557, 16'd52020, 16'd24965, 16'd62728, 16'd12856, 16'd18190, 16'd63432, 16'd62299, 16'd51363, 16'd51835, 16'd30874, 16'd36740, 16'd38671});
	test_expansion(128'h5a9a98b21a9f6392bf72296b6ad1d813, {16'd48152, 16'd45753, 16'd41607, 16'd14879, 16'd18713, 16'd60757, 16'd14150, 16'd42379, 16'd49235, 16'd26990, 16'd24359, 16'd39726, 16'd57297, 16'd58908, 16'd28865, 16'd10775, 16'd56192, 16'd35490, 16'd57027, 16'd55271, 16'd53551, 16'd58994, 16'd31780, 16'd34163, 16'd59095, 16'd16816});
	test_expansion(128'h162ab7757670013a01ac601ed18c54ef, {16'd52902, 16'd5649, 16'd63789, 16'd48111, 16'd20883, 16'd2956, 16'd13258, 16'd28338, 16'd33354, 16'd13520, 16'd40794, 16'd47895, 16'd51748, 16'd54709, 16'd61530, 16'd2998, 16'd10212, 16'd25121, 16'd950, 16'd61687, 16'd11701, 16'd25423, 16'd45040, 16'd51887, 16'd65173, 16'd7788});
	test_expansion(128'ha798e1c09539ac36d527ead8d23c5e45, {16'd62209, 16'd61246, 16'd26893, 16'd29875, 16'd32183, 16'd63507, 16'd11949, 16'd59502, 16'd33857, 16'd13577, 16'd28143, 16'd50308, 16'd28950, 16'd31450, 16'd24518, 16'd7180, 16'd33061, 16'd50795, 16'd8730, 16'd61220, 16'd13666, 16'd59428, 16'd1641, 16'd26775, 16'd49230, 16'd54846});
	test_expansion(128'h503eb2d508c4b14ed379938bd3d9a96b, {16'd9344, 16'd54885, 16'd57445, 16'd2296, 16'd54011, 16'd52677, 16'd3863, 16'd23810, 16'd36584, 16'd43458, 16'd35058, 16'd59415, 16'd5239, 16'd59717, 16'd5455, 16'd60076, 16'd6239, 16'd52658, 16'd63647, 16'd21970, 16'd37967, 16'd38264, 16'd26481, 16'd4745, 16'd9732, 16'd60432});
	test_expansion(128'hd1625b3735bf1c72d15516bf2a98d252, {16'd63208, 16'd39228, 16'd31735, 16'd12495, 16'd818, 16'd48306, 16'd35315, 16'd16467, 16'd31354, 16'd49711, 16'd29091, 16'd62741, 16'd32684, 16'd16060, 16'd21478, 16'd55486, 16'd7686, 16'd22565, 16'd6582, 16'd8587, 16'd60674, 16'd33665, 16'd49112, 16'd17569, 16'd2877, 16'd16045});
	test_expansion(128'h8c297bb2284fa81f9585cdd0b9cee709, {16'd62064, 16'd47775, 16'd38048, 16'd64304, 16'd18789, 16'd52835, 16'd58028, 16'd59662, 16'd35333, 16'd39322, 16'd50439, 16'd7149, 16'd23064, 16'd50741, 16'd15610, 16'd54788, 16'd6205, 16'd32264, 16'd20749, 16'd54021, 16'd17203, 16'd49734, 16'd57241, 16'd39951, 16'd34735, 16'd61260});
	test_expansion(128'h261cd6a5f6a6fb3c1be92d49463f37aa, {16'd43202, 16'd14457, 16'd6371, 16'd41749, 16'd6101, 16'd27354, 16'd62956, 16'd12406, 16'd13314, 16'd24998, 16'd11963, 16'd9501, 16'd54611, 16'd882, 16'd27648, 16'd61967, 16'd19873, 16'd53676, 16'd27602, 16'd57908, 16'd21345, 16'd8216, 16'd34099, 16'd44050, 16'd2551, 16'd59512});
	test_expansion(128'he1006ed73f86817b6252d548ab7c3ea8, {16'd43502, 16'd48266, 16'd17386, 16'd47188, 16'd64660, 16'd2788, 16'd63484, 16'd62682, 16'd49125, 16'd14238, 16'd43932, 16'd38725, 16'd49809, 16'd45667, 16'd29525, 16'd283, 16'd56734, 16'd38742, 16'd32779, 16'd21873, 16'd44253, 16'd57288, 16'd50630, 16'd279, 16'd48168, 16'd52641});
	test_expansion(128'hd048070e255b2fbcd2ec1a352d27c2ee, {16'd24247, 16'd60462, 16'd44780, 16'd32609, 16'd59580, 16'd40581, 16'd1531, 16'd40358, 16'd21438, 16'd44920, 16'd30053, 16'd38240, 16'd49806, 16'd55898, 16'd56107, 16'd23837, 16'd15817, 16'd6452, 16'd53781, 16'd22367, 16'd31197, 16'd60303, 16'd60768, 16'd57579, 16'd11205, 16'd51437});
	test_expansion(128'h2cc5e13fe3d41403ae775d263810eb75, {16'd21132, 16'd57523, 16'd14809, 16'd56081, 16'd11138, 16'd40623, 16'd7865, 16'd29228, 16'd28312, 16'd33252, 16'd60378, 16'd57467, 16'd53079, 16'd38244, 16'd25799, 16'd29340, 16'd40749, 16'd31719, 16'd38284, 16'd191, 16'd62371, 16'd25388, 16'd54392, 16'd48359, 16'd55661, 16'd62461});
	test_expansion(128'h1626c3ea4580846490b0c69dba5a5e4a, {16'd60505, 16'd62929, 16'd3513, 16'd58189, 16'd11995, 16'd13983, 16'd14666, 16'd38067, 16'd34239, 16'd13002, 16'd46852, 16'd62137, 16'd62739, 16'd12385, 16'd60377, 16'd54617, 16'd18383, 16'd31252, 16'd7033, 16'd34331, 16'd25273, 16'd63100, 16'd40632, 16'd31553, 16'd31095, 16'd17801});
	test_expansion(128'hec640bfd4ea6aae3abab9c5f0e695a03, {16'd14200, 16'd59981, 16'd61958, 16'd36484, 16'd5089, 16'd23261, 16'd2886, 16'd62766, 16'd58165, 16'd41877, 16'd30939, 16'd25030, 16'd43114, 16'd13413, 16'd56183, 16'd49864, 16'd34725, 16'd59584, 16'd58894, 16'd56062, 16'd37075, 16'd15750, 16'd48364, 16'd41094, 16'd43446, 16'd7863});
	test_expansion(128'h757b7c05e2e58022784b111b53a43302, {16'd12354, 16'd51054, 16'd25687, 16'd33594, 16'd23365, 16'd53487, 16'd60674, 16'd18805, 16'd51845, 16'd21280, 16'd63155, 16'd39127, 16'd17660, 16'd3930, 16'd25315, 16'd26003, 16'd41635, 16'd55745, 16'd8534, 16'd18073, 16'd17521, 16'd13284, 16'd60441, 16'd28020, 16'd9254, 16'd35357});
	test_expansion(128'ha0fb6d2cc33175f118c61da1d044a44b, {16'd58373, 16'd25126, 16'd50593, 16'd37814, 16'd5645, 16'd25390, 16'd176, 16'd45087, 16'd26885, 16'd39485, 16'd63638, 16'd64844, 16'd7383, 16'd25760, 16'd37041, 16'd40147, 16'd33154, 16'd37064, 16'd11804, 16'd62849, 16'd30965, 16'd22350, 16'd61839, 16'd11946, 16'd1158, 16'd57068});
	test_expansion(128'h01366f970da6fc2fb788eb6cdb607dde, {16'd32663, 16'd60729, 16'd13525, 16'd30181, 16'd36948, 16'd58915, 16'd7333, 16'd14155, 16'd46371, 16'd64900, 16'd63394, 16'd37202, 16'd3971, 16'd64031, 16'd35117, 16'd11560, 16'd5768, 16'd50822, 16'd16633, 16'd23229, 16'd64867, 16'd49337, 16'd30436, 16'd32341, 16'd39881, 16'd13154});
	test_expansion(128'h6fa4068cdb4a2c79fd679fcbc6dc522c, {16'd30962, 16'd27744, 16'd12509, 16'd16183, 16'd34176, 16'd15623, 16'd45797, 16'd35824, 16'd17085, 16'd10692, 16'd4807, 16'd52464, 16'd25490, 16'd50098, 16'd24168, 16'd59501, 16'd38424, 16'd20702, 16'd65477, 16'd35031, 16'd50869, 16'd43708, 16'd57055, 16'd8065, 16'd21268, 16'd23777});
	test_expansion(128'h865ded14173aa0a0ddc77be4a329211e, {16'd16049, 16'd35636, 16'd40778, 16'd39862, 16'd27851, 16'd26587, 16'd23108, 16'd42726, 16'd63808, 16'd37021, 16'd20865, 16'd40057, 16'd12991, 16'd46507, 16'd16388, 16'd22168, 16'd9419, 16'd42482, 16'd26005, 16'd52877, 16'd4523, 16'd41197, 16'd60383, 16'd44114, 16'd53585, 16'd40016});
	test_expansion(128'h6931b9ce252cbb0125f7ad551de07e32, {16'd20508, 16'd17312, 16'd5784, 16'd7516, 16'd50850, 16'd62165, 16'd62665, 16'd15014, 16'd41470, 16'd29195, 16'd49920, 16'd53740, 16'd58696, 16'd15991, 16'd31869, 16'd15875, 16'd57961, 16'd36167, 16'd49748, 16'd3618, 16'd6265, 16'd13780, 16'd48656, 16'd19925, 16'd62529, 16'd41609});
	test_expansion(128'he7afd65259e88c6d1261fa6b7137461c, {16'd45725, 16'd47838, 16'd55071, 16'd20653, 16'd49353, 16'd39943, 16'd5759, 16'd54221, 16'd16873, 16'd38626, 16'd4501, 16'd58764, 16'd35924, 16'd21413, 16'd54341, 16'd3301, 16'd38576, 16'd61913, 16'd35693, 16'd18343, 16'd34752, 16'd22274, 16'd44886, 16'd23761, 16'd482, 16'd35942});
	test_expansion(128'h12bad9240378a632e54476d787a9c7e0, {16'd43383, 16'd58460, 16'd56099, 16'd7299, 16'd42846, 16'd18432, 16'd45536, 16'd62881, 16'd10359, 16'd2048, 16'd13900, 16'd10936, 16'd20310, 16'd3796, 16'd11463, 16'd40935, 16'd12198, 16'd32462, 16'd38968, 16'd53428, 16'd37959, 16'd23795, 16'd50523, 16'd10445, 16'd26437, 16'd35050});
	test_expansion(128'hf78b8c09e9af208d172345d62c1ec8a6, {16'd36397, 16'd10434, 16'd46400, 16'd32800, 16'd25679, 16'd43876, 16'd26053, 16'd28400, 16'd63004, 16'd1306, 16'd26506, 16'd36634, 16'd8724, 16'd52664, 16'd3430, 16'd50779, 16'd17134, 16'd4151, 16'd13444, 16'd1076, 16'd36449, 16'd443, 16'd3343, 16'd29480, 16'd13854, 16'd9190});
	test_expansion(128'h66be6b6838d97f7b8932d5b29bd4e7bc, {16'd36619, 16'd30112, 16'd1734, 16'd34329, 16'd11615, 16'd1219, 16'd5489, 16'd25663, 16'd24915, 16'd61333, 16'd34199, 16'd7918, 16'd19160, 16'd7219, 16'd50526, 16'd13371, 16'd41263, 16'd44688, 16'd8126, 16'd47258, 16'd37352, 16'd30710, 16'd27615, 16'd18903, 16'd16959, 16'd44685});
	test_expansion(128'h9f43ce1e29ec5303e8013ce5e530c305, {16'd9929, 16'd14991, 16'd51734, 16'd10856, 16'd13219, 16'd25296, 16'd62654, 16'd41000, 16'd21435, 16'd2055, 16'd22278, 16'd36749, 16'd46307, 16'd15784, 16'd35348, 16'd3932, 16'd13266, 16'd46116, 16'd38962, 16'd51249, 16'd48719, 16'd61589, 16'd29747, 16'd31853, 16'd23306, 16'd32033});
	test_expansion(128'hd0c4496d05a02b6700656799b5e1acf6, {16'd35068, 16'd48126, 16'd58952, 16'd35722, 16'd14496, 16'd42292, 16'd22224, 16'd62712, 16'd24217, 16'd8962, 16'd55418, 16'd18523, 16'd49481, 16'd21877, 16'd34342, 16'd29347, 16'd19818, 16'd40201, 16'd59584, 16'd7206, 16'd59127, 16'd36532, 16'd16670, 16'd25388, 16'd64918, 16'd46082});
	test_expansion(128'hae226af44a59672ddedffd7335bb54f6, {16'd20202, 16'd38248, 16'd33554, 16'd15822, 16'd3734, 16'd14806, 16'd9377, 16'd51780, 16'd13309, 16'd65493, 16'd2412, 16'd12056, 16'd18817, 16'd35095, 16'd51650, 16'd58006, 16'd63335, 16'd46948, 16'd3469, 16'd50166, 16'd6524, 16'd1982, 16'd42805, 16'd7659, 16'd20888, 16'd35040});
	test_expansion(128'h3378759e53d73ef835bf97595625682b, {16'd28234, 16'd1353, 16'd14745, 16'd30601, 16'd64858, 16'd20188, 16'd29271, 16'd13111, 16'd29473, 16'd53460, 16'd26641, 16'd43226, 16'd56784, 16'd12047, 16'd14266, 16'd3459, 16'd40524, 16'd7250, 16'd61231, 16'd44418, 16'd20261, 16'd57524, 16'd6083, 16'd61705, 16'd62500, 16'd47611});
	test_expansion(128'h5a949f2dc5623014cb89f7379e4b4031, {16'd59287, 16'd64609, 16'd64562, 16'd32706, 16'd46395, 16'd37335, 16'd59194, 16'd45476, 16'd20308, 16'd483, 16'd9703, 16'd64387, 16'd16873, 16'd63422, 16'd62208, 16'd21945, 16'd3557, 16'd10210, 16'd1166, 16'd57906, 16'd59814, 16'd3593, 16'd19216, 16'd17788, 16'd59889, 16'd802});
	test_expansion(128'hf542f76446025bf6c336fa7de273a1e4, {16'd5891, 16'd6220, 16'd37166, 16'd32137, 16'd38150, 16'd14177, 16'd43623, 16'd55418, 16'd35070, 16'd63964, 16'd23840, 16'd45544, 16'd49001, 16'd24892, 16'd38766, 16'd50356, 16'd29223, 16'd5009, 16'd36267, 16'd32187, 16'd28212, 16'd30700, 16'd4324, 16'd4798, 16'd53470, 16'd38784});
	test_expansion(128'h7d9f927efcde26a36b75dd3c4fbbdf94, {16'd12695, 16'd41959, 16'd12564, 16'd31260, 16'd35680, 16'd36823, 16'd39091, 16'd25173, 16'd1834, 16'd35285, 16'd55991, 16'd63920, 16'd4715, 16'd58551, 16'd59821, 16'd32031, 16'd21058, 16'd21487, 16'd6641, 16'd14582, 16'd27585, 16'd55466, 16'd54886, 16'd7683, 16'd23476, 16'd56116});
	test_expansion(128'h7e6a1082b5a09bdacfa1682db910b540, {16'd62833, 16'd32603, 16'd23967, 16'd21115, 16'd22482, 16'd51091, 16'd33711, 16'd42168, 16'd18206, 16'd39625, 16'd30801, 16'd47247, 16'd60197, 16'd42843, 16'd55254, 16'd65445, 16'd47766, 16'd15614, 16'd64568, 16'd51773, 16'd4936, 16'd14186, 16'd21669, 16'd17148, 16'd43989, 16'd13231});
	test_expansion(128'hd5572da33b08e5788d8d7f76cc08da0b, {16'd26472, 16'd43790, 16'd14298, 16'd46802, 16'd48419, 16'd3649, 16'd4690, 16'd41825, 16'd57857, 16'd48466, 16'd4091, 16'd46926, 16'd42762, 16'd19860, 16'd1288, 16'd24794, 16'd28666, 16'd64454, 16'd43582, 16'd37, 16'd57132, 16'd4175, 16'd14073, 16'd19107, 16'd4656, 16'd14049});
	test_expansion(128'h6277d8ce589651802903150d81abc658, {16'd7459, 16'd36786, 16'd28460, 16'd55239, 16'd4609, 16'd9433, 16'd2468, 16'd46059, 16'd30299, 16'd13794, 16'd16496, 16'd42145, 16'd18769, 16'd5053, 16'd55393, 16'd32260, 16'd65500, 16'd62782, 16'd16068, 16'd27424, 16'd31435, 16'd48432, 16'd49226, 16'd25119, 16'd505, 16'd15024});
	test_expansion(128'he6e4a2b7741ba5c0684f2282652696c2, {16'd26665, 16'd48631, 16'd65159, 16'd49342, 16'd8128, 16'd3482, 16'd10915, 16'd5861, 16'd12030, 16'd3054, 16'd33202, 16'd17852, 16'd9882, 16'd50173, 16'd62188, 16'd4261, 16'd21299, 16'd51070, 16'd14853, 16'd62061, 16'd32133, 16'd48247, 16'd35084, 16'd2647, 16'd58778, 16'd48582});
	test_expansion(128'ha98040e3077a3c746900d6bfc4c18126, {16'd35111, 16'd1765, 16'd21335, 16'd53165, 16'd349, 16'd57529, 16'd57964, 16'd34535, 16'd40868, 16'd50698, 16'd50359, 16'd58945, 16'd63307, 16'd13749, 16'd9012, 16'd2751, 16'd37446, 16'd49453, 16'd775, 16'd8132, 16'd55788, 16'd12080, 16'd30843, 16'd44434, 16'd65465, 16'd47451});
	test_expansion(128'hc21e2e824718e872ace27f227b141edf, {16'd63441, 16'd49867, 16'd20556, 16'd13436, 16'd49661, 16'd33519, 16'd52435, 16'd30695, 16'd29673, 16'd41348, 16'd33406, 16'd62089, 16'd50918, 16'd23836, 16'd28632, 16'd732, 16'd44054, 16'd35122, 16'd41347, 16'd30284, 16'd21590, 16'd62320, 16'd54411, 16'd29848, 16'd50003, 16'd62085});
	test_expansion(128'hcf3ba0c1b8808e8b21ee6b8ad24b57a1, {16'd33131, 16'd51787, 16'd35327, 16'd10154, 16'd19366, 16'd42857, 16'd15323, 16'd4224, 16'd22350, 16'd36001, 16'd53432, 16'd58901, 16'd42629, 16'd4047, 16'd40130, 16'd33939, 16'd40763, 16'd10884, 16'd20571, 16'd38020, 16'd37171, 16'd65174, 16'd15666, 16'd14148, 16'd25136, 16'd62040});
	test_expansion(128'h5e445fd41535691b1b9c2fd7bd3bf4a3, {16'd28543, 16'd33172, 16'd43160, 16'd61802, 16'd23693, 16'd11372, 16'd32524, 16'd22080, 16'd2333, 16'd140, 16'd17942, 16'd43585, 16'd62713, 16'd14273, 16'd60813, 16'd53188, 16'd38603, 16'd25631, 16'd49907, 16'd16933, 16'd28416, 16'd42105, 16'd38941, 16'd18518, 16'd49155, 16'd19881});
	test_expansion(128'h03d07a0873f6700b73e0c1d236f43889, {16'd44101, 16'd51463, 16'd4355, 16'd31938, 16'd55060, 16'd58454, 16'd58651, 16'd44826, 16'd29014, 16'd17977, 16'd44545, 16'd18037, 16'd43961, 16'd41640, 16'd58091, 16'd23377, 16'd23611, 16'd42133, 16'd61156, 16'd22982, 16'd47590, 16'd1266, 16'd13305, 16'd1363, 16'd57866, 16'd61506});
	test_expansion(128'h7b8170403875aa17b20ee08b35108cba, {16'd38584, 16'd44166, 16'd56150, 16'd64528, 16'd62541, 16'd37607, 16'd41833, 16'd5195, 16'd23837, 16'd64544, 16'd47844, 16'd6260, 16'd14717, 16'd64939, 16'd56909, 16'd40458, 16'd55979, 16'd6887, 16'd36306, 16'd61915, 16'd18186, 16'd28641, 16'd35765, 16'd15237, 16'd27452, 16'd29086});
	test_expansion(128'h341d6bebce4e63e99e6c1271b87969a4, {16'd4028, 16'd50482, 16'd64396, 16'd55149, 16'd3025, 16'd28963, 16'd4995, 16'd4876, 16'd31584, 16'd59242, 16'd27558, 16'd29231, 16'd57724, 16'd60616, 16'd47380, 16'd53890, 16'd26762, 16'd53167, 16'd9371, 16'd62182, 16'd37103, 16'd18156, 16'd21051, 16'd28526, 16'd2996, 16'd43683});
	test_expansion(128'h71dbd67fdd28dcb83f0c294907941d3b, {16'd37830, 16'd52068, 16'd51401, 16'd55760, 16'd8578, 16'd31645, 16'd52676, 16'd42787, 16'd43555, 16'd5262, 16'd45361, 16'd56097, 16'd31906, 16'd17176, 16'd21961, 16'd37471, 16'd27385, 16'd18062, 16'd47281, 16'd59388, 16'd48442, 16'd24841, 16'd41661, 16'd8922, 16'd15603, 16'd6558});
	test_expansion(128'h2184735c04235ac200eb31ede3a2c571, {16'd41475, 16'd33544, 16'd9859, 16'd59154, 16'd23993, 16'd21878, 16'd25107, 16'd22045, 16'd57467, 16'd54476, 16'd27687, 16'd45866, 16'd18337, 16'd5491, 16'd56652, 16'd49255, 16'd2289, 16'd8588, 16'd45619, 16'd53221, 16'd31503, 16'd43957, 16'd37753, 16'd38775, 16'd60854, 16'd28187});
	test_expansion(128'h44b1d8b74507a6ecedcbdcea9a7720e7, {16'd12018, 16'd44757, 16'd47537, 16'd31638, 16'd25988, 16'd58650, 16'd63754, 16'd39302, 16'd52700, 16'd19807, 16'd62537, 16'd6462, 16'd51651, 16'd10637, 16'd24027, 16'd28685, 16'd54286, 16'd18994, 16'd51118, 16'd31966, 16'd56967, 16'd42658, 16'd19602, 16'd13447, 16'd60969, 16'd16162});
	test_expansion(128'h4f5fdd83e6689857692d4a9c89aded2b, {16'd16177, 16'd5541, 16'd58378, 16'd56766, 16'd27562, 16'd29866, 16'd22431, 16'd56286, 16'd25859, 16'd13604, 16'd63297, 16'd55705, 16'd56644, 16'd33471, 16'd5767, 16'd55517, 16'd27334, 16'd44877, 16'd11234, 16'd17133, 16'd34342, 16'd49947, 16'd32713, 16'd7157, 16'd42719, 16'd15182});
	test_expansion(128'h9fbc2ea733c46c0839edfbfe6715258d, {16'd457, 16'd33458, 16'd32289, 16'd23247, 16'd36289, 16'd55369, 16'd30907, 16'd31522, 16'd21701, 16'd16117, 16'd35558, 16'd32183, 16'd22265, 16'd40869, 16'd55847, 16'd6661, 16'd41127, 16'd54501, 16'd60359, 16'd43241, 16'd50457, 16'd35996, 16'd12355, 16'd57473, 16'd60613, 16'd35857});
	test_expansion(128'hc4b5f7c9409e8c205132b4c403e9650e, {16'd27664, 16'd46211, 16'd48087, 16'd24282, 16'd33820, 16'd29960, 16'd38642, 16'd17202, 16'd25158, 16'd60496, 16'd11715, 16'd61531, 16'd54504, 16'd11332, 16'd37346, 16'd40592, 16'd29523, 16'd44096, 16'd35223, 16'd52793, 16'd32825, 16'd9434, 16'd10841, 16'd26634, 16'd21391, 16'd50164});
	test_expansion(128'h41e20670c6766867a71edd1f4869f83c, {16'd40943, 16'd46496, 16'd33280, 16'd60505, 16'd25815, 16'd7084, 16'd5262, 16'd36463, 16'd5801, 16'd15728, 16'd3722, 16'd13205, 16'd57537, 16'd19152, 16'd50402, 16'd14027, 16'd56986, 16'd1004, 16'd47879, 16'd30406, 16'd33202, 16'd35017, 16'd640, 16'd17676, 16'd4125, 16'd61648});
	test_expansion(128'ha6ae9a1ad4f6bcf62287bed69ef0619d, {16'd60239, 16'd13406, 16'd32953, 16'd25994, 16'd12803, 16'd47500, 16'd37033, 16'd57998, 16'd17660, 16'd55177, 16'd21876, 16'd62351, 16'd32594, 16'd29583, 16'd62651, 16'd20011, 16'd56753, 16'd13493, 16'd25959, 16'd21185, 16'd59969, 16'd64981, 16'd53394, 16'd7165, 16'd6919, 16'd49970});
	test_expansion(128'h782cccee3538f4b32a003597f6b1f521, {16'd29131, 16'd47947, 16'd11126, 16'd53448, 16'd23842, 16'd51053, 16'd8531, 16'd2612, 16'd6247, 16'd29326, 16'd58201, 16'd14734, 16'd24770, 16'd19614, 16'd64028, 16'd46836, 16'd42371, 16'd58505, 16'd7775, 16'd16838, 16'd9407, 16'd10137, 16'd756, 16'd38215, 16'd44967, 16'd28008});
	test_expansion(128'hb47eac917ded92f8d0408805b01a8810, {16'd32679, 16'd31876, 16'd13118, 16'd31856, 16'd39286, 16'd37067, 16'd3240, 16'd62219, 16'd28614, 16'd16399, 16'd12342, 16'd10387, 16'd50645, 16'd8151, 16'd56651, 16'd61862, 16'd58801, 16'd10510, 16'd46282, 16'd4308, 16'd16491, 16'd38878, 16'd25430, 16'd44042, 16'd32171, 16'd56716});
	test_expansion(128'h6cc7c0e48ab43476d71a768e4834a879, {16'd14403, 16'd18345, 16'd21807, 16'd23908, 16'd52852, 16'd59426, 16'd29097, 16'd40629, 16'd35314, 16'd25985, 16'd370, 16'd51433, 16'd38070, 16'd11318, 16'd22776, 16'd65110, 16'd24078, 16'd23941, 16'd35593, 16'd43455, 16'd27525, 16'd30219, 16'd12807, 16'd44349, 16'd15791, 16'd7562});
	test_expansion(128'hcb2429442afe12b021766e0e16a085fc, {16'd26650, 16'd9689, 16'd30198, 16'd46778, 16'd7806, 16'd7957, 16'd48005, 16'd29317, 16'd29412, 16'd30645, 16'd47457, 16'd44864, 16'd9984, 16'd48077, 16'd40922, 16'd21368, 16'd52035, 16'd4729, 16'd31972, 16'd56706, 16'd18299, 16'd41352, 16'd58609, 16'd61847, 16'd11607, 16'd34214});
	test_expansion(128'h285025e897de998d5c22403e80a7a6e8, {16'd41698, 16'd57954, 16'd5807, 16'd15690, 16'd5685, 16'd32459, 16'd25719, 16'd43210, 16'd43916, 16'd14873, 16'd24642, 16'd25732, 16'd26198, 16'd1663, 16'd51451, 16'd9013, 16'd30299, 16'd19715, 16'd54371, 16'd23852, 16'd16116, 16'd17567, 16'd6957, 16'd12686, 16'd40792, 16'd14201});
	test_expansion(128'h87f36a0438b2ee9679078b352be47873, {16'd3949, 16'd6174, 16'd60975, 16'd42578, 16'd62992, 16'd53627, 16'd58647, 16'd32354, 16'd17142, 16'd43076, 16'd22896, 16'd42387, 16'd65062, 16'd65227, 16'd27038, 16'd47880, 16'd13458, 16'd4207, 16'd49603, 16'd54015, 16'd15753, 16'd32234, 16'd44756, 16'd40057, 16'd26758, 16'd15229});
	test_expansion(128'hca6bcafa7bce6fa913eccc47f2ed7a9e, {16'd60584, 16'd19648, 16'd32373, 16'd26082, 16'd11088, 16'd19657, 16'd47601, 16'd7016, 16'd53069, 16'd38131, 16'd36019, 16'd45187, 16'd27568, 16'd18909, 16'd41291, 16'd1665, 16'd56017, 16'd32555, 16'd14162, 16'd195, 16'd41313, 16'd19106, 16'd54879, 16'd49977, 16'd35845, 16'd11077});
	test_expansion(128'hda4f967a4ea57c83044bf8e4772294d9, {16'd53707, 16'd27951, 16'd63678, 16'd55720, 16'd24072, 16'd44353, 16'd7694, 16'd49743, 16'd56656, 16'd13083, 16'd43099, 16'd55025, 16'd13400, 16'd54822, 16'd59600, 16'd22842, 16'd41773, 16'd3490, 16'd49476, 16'd6051, 16'd12286, 16'd44742, 16'd12891, 16'd4242, 16'd55133, 16'd36124});
	test_expansion(128'h99f0b57c6c5c323dc833a656561b2807, {16'd33061, 16'd20514, 16'd42419, 16'd35041, 16'd7182, 16'd19784, 16'd21063, 16'd47692, 16'd7040, 16'd13006, 16'd63624, 16'd52901, 16'd6592, 16'd8947, 16'd7310, 16'd1957, 16'd26264, 16'd28198, 16'd8158, 16'd54339, 16'd8903, 16'd21568, 16'd8752, 16'd24376, 16'd8480, 16'd2164});
	test_expansion(128'h74e9d25a647063bad8dc2131ff37bc3e, {16'd10429, 16'd340, 16'd54304, 16'd57102, 16'd60889, 16'd33099, 16'd25297, 16'd45061, 16'd9107, 16'd53784, 16'd57945, 16'd8889, 16'd543, 16'd26074, 16'd27730, 16'd2763, 16'd41969, 16'd33404, 16'd15807, 16'd2317, 16'd12143, 16'd59826, 16'd52802, 16'd37569, 16'd33261, 16'd63372});
	test_expansion(128'h810acd9469898741fa83de6a41af2c71, {16'd17707, 16'd39288, 16'd52305, 16'd21515, 16'd46136, 16'd63553, 16'd32352, 16'd60271, 16'd27812, 16'd63349, 16'd65132, 16'd15860, 16'd17319, 16'd44986, 16'd65208, 16'd29181, 16'd46371, 16'd52479, 16'd16994, 16'd42140, 16'd24850, 16'd45883, 16'd45352, 16'd47751, 16'd25502, 16'd40660});
	test_expansion(128'h14e9282226af862b6ca8f1d5ca9a1915, {16'd18421, 16'd62672, 16'd37400, 16'd43695, 16'd28653, 16'd7811, 16'd27887, 16'd49506, 16'd1178, 16'd39317, 16'd42838, 16'd37957, 16'd44665, 16'd33604, 16'd49403, 16'd24788, 16'd4894, 16'd25020, 16'd24300, 16'd19292, 16'd37709, 16'd9471, 16'd34679, 16'd43332, 16'd28292, 16'd22297});
	test_expansion(128'hf9e25b4bd1e58b8851a487bb5f1df65f, {16'd34726, 16'd2321, 16'd2834, 16'd32051, 16'd921, 16'd25038, 16'd64165, 16'd22273, 16'd64195, 16'd11350, 16'd16229, 16'd28036, 16'd1061, 16'd21124, 16'd45145, 16'd5641, 16'd63387, 16'd51917, 16'd22711, 16'd19494, 16'd39107, 16'd27993, 16'd50033, 16'd34334, 16'd50012, 16'd31388});
	test_expansion(128'h3ff9519714b47d7840387d20a9d56fbc, {16'd18628, 16'd56171, 16'd590, 16'd4483, 16'd25394, 16'd39738, 16'd37729, 16'd10718, 16'd25609, 16'd60507, 16'd56706, 16'd17396, 16'd13360, 16'd21611, 16'd31698, 16'd30331, 16'd31908, 16'd5191, 16'd26076, 16'd39179, 16'd52652, 16'd43310, 16'd37595, 16'd30246, 16'd29441, 16'd44543});
	test_expansion(128'h96df22121b649d1875b20ba39e2827b8, {16'd9449, 16'd6898, 16'd62846, 16'd32240, 16'd37621, 16'd12347, 16'd7285, 16'd12838, 16'd41951, 16'd62658, 16'd64190, 16'd42237, 16'd52417, 16'd14618, 16'd28636, 16'd52939, 16'd55162, 16'd59017, 16'd24911, 16'd39004, 16'd5782, 16'd56687, 16'd47693, 16'd17747, 16'd9328, 16'd42307});
	test_expansion(128'hfe2307df2ee150aaa242091349f55a35, {16'd54449, 16'd12804, 16'd10364, 16'd58760, 16'd28345, 16'd5784, 16'd10223, 16'd44171, 16'd58543, 16'd17407, 16'd59103, 16'd14679, 16'd45080, 16'd27958, 16'd6467, 16'd22687, 16'd43639, 16'd29223, 16'd65380, 16'd56153, 16'd53058, 16'd39860, 16'd12563, 16'd52410, 16'd22947, 16'd38081});
	test_expansion(128'ha597ad19f489f5a54f700abd4f2baf2c, {16'd12587, 16'd8696, 16'd23969, 16'd34186, 16'd14350, 16'd61929, 16'd3745, 16'd30738, 16'd60880, 16'd11790, 16'd58111, 16'd25360, 16'd40962, 16'd26201, 16'd37537, 16'd7558, 16'd5527, 16'd59895, 16'd36539, 16'd32407, 16'd42532, 16'd25020, 16'd25776, 16'd38209, 16'd58399, 16'd21663});
	test_expansion(128'h26788a75f3fde254adcddde6aa9f30ce, {16'd44061, 16'd25444, 16'd17518, 16'd20342, 16'd52041, 16'd24980, 16'd48570, 16'd29093, 16'd46478, 16'd33183, 16'd28048, 16'd37936, 16'd49716, 16'd40691, 16'd915, 16'd29370, 16'd5628, 16'd4879, 16'd17949, 16'd30841, 16'd52773, 16'd703, 16'd32282, 16'd22469, 16'd1899, 16'd35288});
	test_expansion(128'h0cad2156f2265a049980cd4029a5b182, {16'd29396, 16'd52637, 16'd19793, 16'd42237, 16'd12464, 16'd5464, 16'd39766, 16'd42236, 16'd38869, 16'd41080, 16'd26280, 16'd57798, 16'd53976, 16'd13275, 16'd53226, 16'd54720, 16'd20806, 16'd65535, 16'd28290, 16'd46060, 16'd21489, 16'd57733, 16'd38504, 16'd337, 16'd57078, 16'd9712});
	test_expansion(128'h6625c936485e54fc34866ec41fff7051, {16'd30030, 16'd41885, 16'd24571, 16'd60427, 16'd48423, 16'd25884, 16'd31911, 16'd25914, 16'd25981, 16'd63893, 16'd9572, 16'd40596, 16'd29958, 16'd19687, 16'd45246, 16'd333, 16'd50097, 16'd26090, 16'd27623, 16'd17290, 16'd58482, 16'd52984, 16'd26710, 16'd17483, 16'd8024, 16'd23719});
	test_expansion(128'h15c057a19f968f19ab0ca716ea02769b, {16'd41626, 16'd33119, 16'd8699, 16'd31290, 16'd6980, 16'd62847, 16'd45917, 16'd45697, 16'd64983, 16'd35751, 16'd6259, 16'd41434, 16'd12848, 16'd26912, 16'd36630, 16'd1353, 16'd56208, 16'd56131, 16'd51801, 16'd23891, 16'd5103, 16'd53494, 16'd64668, 16'd46339, 16'd16597, 16'd18828});
	test_expansion(128'h617b7869257c9570d7d857e9c9010c38, {16'd16893, 16'd36174, 16'd55722, 16'd57649, 16'd21806, 16'd45480, 16'd61463, 16'd63674, 16'd14486, 16'd48608, 16'd1398, 16'd39250, 16'd22114, 16'd51394, 16'd33487, 16'd27099, 16'd14136, 16'd62528, 16'd25299, 16'd48203, 16'd2003, 16'd42363, 16'd20165, 16'd50842, 16'd57499, 16'd61933});
	test_expansion(128'h45baf60dc82e5ab9daf59b72a56f2793, {16'd19858, 16'd52686, 16'd16575, 16'd51685, 16'd23304, 16'd40743, 16'd17517, 16'd47081, 16'd50713, 16'd40709, 16'd44378, 16'd29868, 16'd5105, 16'd9462, 16'd19127, 16'd56454, 16'd9323, 16'd48569, 16'd28215, 16'd19455, 16'd54410, 16'd21410, 16'd21562, 16'd54978, 16'd6294, 16'd16723});
	test_expansion(128'h49bb844a66e6d4a18b39556a9098839b, {16'd26499, 16'd62471, 16'd44503, 16'd9273, 16'd19806, 16'd17991, 16'd64971, 16'd50164, 16'd41633, 16'd40998, 16'd27723, 16'd40267, 16'd59643, 16'd25276, 16'd38303, 16'd4689, 16'd29578, 16'd4701, 16'd38024, 16'd35225, 16'd36284, 16'd9825, 16'd64958, 16'd51686, 16'd20426, 16'd34701});
	test_expansion(128'h3464083eecbd918efdbc915286aeb658, {16'd38372, 16'd9843, 16'd53765, 16'd61388, 16'd49426, 16'd38272, 16'd50193, 16'd41508, 16'd28587, 16'd56285, 16'd56773, 16'd8104, 16'd56137, 16'd49180, 16'd49705, 16'd30250, 16'd7658, 16'd42686, 16'd63345, 16'd2522, 16'd424, 16'd63065, 16'd10602, 16'd26865, 16'd45370, 16'd2319});
	test_expansion(128'h818e5de024823b385e4c458a5a293f97, {16'd59021, 16'd43869, 16'd50717, 16'd60952, 16'd12454, 16'd50031, 16'd488, 16'd30922, 16'd22227, 16'd21296, 16'd63588, 16'd51069, 16'd22038, 16'd26491, 16'd63245, 16'd55629, 16'd37284, 16'd50998, 16'd54418, 16'd1911, 16'd25319, 16'd64000, 16'd40706, 16'd37571, 16'd11300, 16'd20498});
	test_expansion(128'h650d85adf293e3a95193e1f148b09ff0, {16'd19183, 16'd61689, 16'd180, 16'd21314, 16'd11117, 16'd57756, 16'd14408, 16'd51489, 16'd13434, 16'd39374, 16'd15406, 16'd7039, 16'd54309, 16'd6829, 16'd54082, 16'd41862, 16'd60624, 16'd9612, 16'd21796, 16'd32509, 16'd61396, 16'd8244, 16'd62368, 16'd28044, 16'd31445, 16'd1415});
	test_expansion(128'hc991568d21e6d560b026b2e050958232, {16'd24104, 16'd508, 16'd31977, 16'd59123, 16'd31782, 16'd51469, 16'd15567, 16'd19240, 16'd59770, 16'd39932, 16'd24818, 16'd63859, 16'd17520, 16'd6813, 16'd2049, 16'd59892, 16'd23316, 16'd33427, 16'd47745, 16'd137, 16'd50869, 16'd53968, 16'd19191, 16'd56048, 16'd20247, 16'd28600});
	test_expansion(128'h6cfd902f9ddf368f2bdb9b66c6e20b7a, {16'd21479, 16'd6178, 16'd50867, 16'd50254, 16'd912, 16'd16901, 16'd51123, 16'd25348, 16'd23834, 16'd59981, 16'd44706, 16'd11679, 16'd8824, 16'd54833, 16'd29782, 16'd25306, 16'd23830, 16'd34707, 16'd22799, 16'd45632, 16'd57038, 16'd30664, 16'd48494, 16'd7457, 16'd60522, 16'd29690});
	test_expansion(128'h8ea4671f53831ff714a4fa2ffef4719d, {16'd18993, 16'd57987, 16'd49838, 16'd26540, 16'd59684, 16'd39664, 16'd60878, 16'd49109, 16'd34794, 16'd16304, 16'd43608, 16'd39077, 16'd37240, 16'd42000, 16'd13351, 16'd33100, 16'd37027, 16'd27745, 16'd56073, 16'd16078, 16'd65181, 16'd24422, 16'd49584, 16'd9749, 16'd26617, 16'd3794});
	test_expansion(128'he537698bfff0a0f8013a5cc2f75783ab, {16'd28989, 16'd48698, 16'd34335, 16'd8850, 16'd8877, 16'd64438, 16'd2835, 16'd35147, 16'd58932, 16'd50777, 16'd41324, 16'd56514, 16'd1828, 16'd49386, 16'd5599, 16'd8413, 16'd49643, 16'd37812, 16'd41929, 16'd53875, 16'd18388, 16'd36076, 16'd25843, 16'd19396, 16'd45942, 16'd24288});
	test_expansion(128'h89054dcb12c3156c794975883257623d, {16'd53785, 16'd20702, 16'd58518, 16'd59068, 16'd58163, 16'd14525, 16'd24781, 16'd15584, 16'd32957, 16'd64726, 16'd26812, 16'd6691, 16'd63813, 16'd12851, 16'd45450, 16'd55702, 16'd7888, 16'd2138, 16'd35385, 16'd56657, 16'd52265, 16'd51902, 16'd46552, 16'd32585, 16'd52759, 16'd7390});
	test_expansion(128'h1210e0202f34567576807652e9fb7038, {16'd43144, 16'd47920, 16'd52962, 16'd8125, 16'd23311, 16'd35696, 16'd54564, 16'd58919, 16'd24715, 16'd9633, 16'd27539, 16'd32461, 16'd19647, 16'd58202, 16'd58781, 16'd13445, 16'd43643, 16'd56420, 16'd3008, 16'd4404, 16'd41923, 16'd31572, 16'd56556, 16'd44754, 16'd29787, 16'd14836});
	test_expansion(128'h40f6c5eb72413196ddf64625e1ade710, {16'd28961, 16'd10902, 16'd13488, 16'd63425, 16'd53416, 16'd16886, 16'd5677, 16'd47090, 16'd15117, 16'd50411, 16'd56259, 16'd22294, 16'd3822, 16'd4062, 16'd9615, 16'd32725, 16'd16793, 16'd31026, 16'd43715, 16'd43248, 16'd61971, 16'd18914, 16'd33997, 16'd13154, 16'd44942, 16'd7293});
	test_expansion(128'hd7dabd78937f5e705b0c85fb0951c78b, {16'd22971, 16'd65034, 16'd3223, 16'd41757, 16'd26909, 16'd57667, 16'd16923, 16'd28028, 16'd24694, 16'd64470, 16'd55081, 16'd17050, 16'd35560, 16'd13619, 16'd4207, 16'd16849, 16'd31902, 16'd38051, 16'd53293, 16'd35404, 16'd7824, 16'd54577, 16'd4141, 16'd6049, 16'd8006, 16'd6822});
	test_expansion(128'h53ef2ffb4499bf5537ca39fe4d9c76e4, {16'd9403, 16'd21496, 16'd48575, 16'd23810, 16'd16802, 16'd11006, 16'd16175, 16'd41435, 16'd5937, 16'd63442, 16'd30129, 16'd49313, 16'd21919, 16'd2117, 16'd55900, 16'd20684, 16'd41775, 16'd25083, 16'd46629, 16'd53214, 16'd54421, 16'd47561, 16'd50950, 16'd45638, 16'd16706, 16'd32574});
	test_expansion(128'hb54bcf88b213b4cb2c8b55464008748c, {16'd22682, 16'd49328, 16'd57600, 16'd59695, 16'd7211, 16'd59154, 16'd54740, 16'd14187, 16'd15460, 16'd49624, 16'd20584, 16'd64223, 16'd36512, 16'd60699, 16'd60901, 16'd62035, 16'd16800, 16'd30430, 16'd44058, 16'd26937, 16'd2675, 16'd8101, 16'd11466, 16'd1581, 16'd17499, 16'd42809});
	test_expansion(128'h8bf69f3647ef67cbd8ebbb4d91781b28, {16'd20260, 16'd6474, 16'd18508, 16'd27847, 16'd55649, 16'd64871, 16'd42284, 16'd18303, 16'd13584, 16'd3920, 16'd41953, 16'd15363, 16'd49493, 16'd27806, 16'd25938, 16'd5843, 16'd58255, 16'd55859, 16'd24341, 16'd22961, 16'd27028, 16'd12288, 16'd58371, 16'd27825, 16'd52411, 16'd34003});
	test_expansion(128'h091e5246ff336bdc9ae1b1e25320201e, {16'd35365, 16'd16423, 16'd41572, 16'd45072, 16'd49937, 16'd61066, 16'd34821, 16'd53465, 16'd6575, 16'd4135, 16'd20077, 16'd29651, 16'd31032, 16'd11163, 16'd2049, 16'd57003, 16'd21053, 16'd10980, 16'd18162, 16'd796, 16'd21755, 16'd904, 16'd13772, 16'd64083, 16'd8919, 16'd59959});
	test_expansion(128'h36fa757730b3dea592d60b23d33f79c1, {16'd18357, 16'd27785, 16'd6771, 16'd50796, 16'd39160, 16'd4332, 16'd58374, 16'd52625, 16'd50669, 16'd49144, 16'd53024, 16'd9233, 16'd23065, 16'd6844, 16'd18105, 16'd59061, 16'd9387, 16'd13053, 16'd37585, 16'd34192, 16'd38785, 16'd31038, 16'd44539, 16'd15547, 16'd25775, 16'd46081});
	test_expansion(128'h4cbbaa96e6dc5f7262d93366058b2b73, {16'd54434, 16'd21417, 16'd26288, 16'd54627, 16'd8696, 16'd12279, 16'd5661, 16'd57494, 16'd29456, 16'd5980, 16'd36600, 16'd61076, 16'd13934, 16'd61491, 16'd47207, 16'd45660, 16'd54516, 16'd18239, 16'd36300, 16'd28139, 16'd2582, 16'd60415, 16'd24162, 16'd39684, 16'd5631, 16'd37537});
	test_expansion(128'h2895e1c4669994e2bdbbe775f496030e, {16'd57772, 16'd18640, 16'd8315, 16'd14745, 16'd15133, 16'd31113, 16'd37218, 16'd62239, 16'd60970, 16'd54555, 16'd19682, 16'd58910, 16'd59413, 16'd9053, 16'd31868, 16'd63632, 16'd30508, 16'd38019, 16'd34550, 16'd40268, 16'd59163, 16'd38825, 16'd33897, 16'd14702, 16'd33776, 16'd38787});
	test_expansion(128'hbebd76350cc3812429d8ee77e8fa5744, {16'd59914, 16'd46128, 16'd25658, 16'd39041, 16'd19796, 16'd6256, 16'd6735, 16'd45354, 16'd6397, 16'd10837, 16'd305, 16'd8685, 16'd18862, 16'd1927, 16'd32024, 16'd21024, 16'd65258, 16'd54980, 16'd39781, 16'd25307, 16'd45140, 16'd41877, 16'd6654, 16'd41715, 16'd55586, 16'd23151});
	test_expansion(128'h1651f7dd041f1456fe803ac53a9ce0b6, {16'd25318, 16'd2715, 16'd43807, 16'd1090, 16'd19612, 16'd51470, 16'd50690, 16'd6720, 16'd8699, 16'd5022, 16'd1279, 16'd12468, 16'd23427, 16'd15109, 16'd9033, 16'd8487, 16'd31246, 16'd23977, 16'd46054, 16'd43320, 16'd1061, 16'd31360, 16'd35963, 16'd48649, 16'd52421, 16'd5120});
	test_expansion(128'hdde3d70e7be1892ba674b0f598de9707, {16'd51803, 16'd33173, 16'd18307, 16'd3509, 16'd41944, 16'd10444, 16'd43445, 16'd20062, 16'd16778, 16'd58687, 16'd45667, 16'd48584, 16'd52211, 16'd52253, 16'd22709, 16'd4886, 16'd37574, 16'd47603, 16'd57328, 16'd41171, 16'd41727, 16'd62182, 16'd41411, 16'd49845, 16'd15318, 16'd32490});
	test_expansion(128'h5eed8b44b55350715c8ca5889ba25986, {16'd57222, 16'd61236, 16'd30726, 16'd6994, 16'd55819, 16'd5675, 16'd8375, 16'd14917, 16'd17231, 16'd55654, 16'd62907, 16'd49910, 16'd1099, 16'd27479, 16'd34772, 16'd1264, 16'd48857, 16'd12614, 16'd2729, 16'd6200, 16'd657, 16'd60001, 16'd59389, 16'd44836, 16'd34859, 16'd58057});
	test_expansion(128'h3798ca132bfcc6eab755d4097394dd37, {16'd54029, 16'd47605, 16'd47334, 16'd2340, 16'd38847, 16'd53586, 16'd1610, 16'd48900, 16'd42005, 16'd65061, 16'd45166, 16'd44550, 16'd38211, 16'd32515, 16'd42525, 16'd12211, 16'd17450, 16'd53609, 16'd32633, 16'd47028, 16'd15306, 16'd17193, 16'd34036, 16'd18678, 16'd12549, 16'd44808});
	test_expansion(128'h7842d572de9bc7139f5817e5f4517169, {16'd59268, 16'd24453, 16'd63680, 16'd56006, 16'd38787, 16'd34809, 16'd37396, 16'd14645, 16'd27632, 16'd14346, 16'd38935, 16'd13577, 16'd1715, 16'd20171, 16'd59239, 16'd6635, 16'd26426, 16'd60011, 16'd60923, 16'd39952, 16'd24991, 16'd38002, 16'd6509, 16'd14907, 16'd49077, 16'd31557});
	test_expansion(128'hd5bdf7766f15576a12b3f60a9d395b87, {16'd7627, 16'd59917, 16'd31424, 16'd32582, 16'd26224, 16'd45475, 16'd14390, 16'd20254, 16'd55632, 16'd27577, 16'd35558, 16'd51995, 16'd46718, 16'd48368, 16'd1264, 16'd43428, 16'd33613, 16'd10246, 16'd56792, 16'd27442, 16'd54703, 16'd11387, 16'd50388, 16'd64338, 16'd9764, 16'd42792});
	test_expansion(128'h7dcc5837ee112060a2f3d301937eed5a, {16'd37126, 16'd43841, 16'd3399, 16'd58442, 16'd48871, 16'd34277, 16'd43256, 16'd538, 16'd26042, 16'd54633, 16'd54482, 16'd36050, 16'd53684, 16'd20158, 16'd26288, 16'd30147, 16'd38372, 16'd14898, 16'd52451, 16'd14349, 16'd16772, 16'd60997, 16'd34364, 16'd47559, 16'd9340, 16'd9598});
	test_expansion(128'h4169463189472c45a579c9830a8af470, {16'd39888, 16'd26673, 16'd16123, 16'd22994, 16'd9053, 16'd65371, 16'd35453, 16'd38340, 16'd61397, 16'd17774, 16'd49256, 16'd15835, 16'd2383, 16'd29554, 16'd49854, 16'd52745, 16'd11890, 16'd27564, 16'd52327, 16'd49471, 16'd52168, 16'd5744, 16'd54337, 16'd28936, 16'd58268, 16'd37793});
	test_expansion(128'h218fb9bb9860244a640ef9818bce3e1f, {16'd37950, 16'd10468, 16'd11291, 16'd61000, 16'd20312, 16'd27518, 16'd59275, 16'd25381, 16'd41465, 16'd7648, 16'd23325, 16'd60038, 16'd22987, 16'd18686, 16'd57898, 16'd48431, 16'd3173, 16'd24613, 16'd33548, 16'd4733, 16'd15875, 16'd45069, 16'd26751, 16'd30769, 16'd41984, 16'd53738});
	test_expansion(128'h411e0a0da1380349d3c750fee31e26d3, {16'd31932, 16'd14446, 16'd30918, 16'd40075, 16'd56958, 16'd62392, 16'd56035, 16'd48460, 16'd60547, 16'd8845, 16'd802, 16'd59361, 16'd52421, 16'd59433, 16'd23213, 16'd28243, 16'd20215, 16'd1764, 16'd28713, 16'd5102, 16'd42201, 16'd18104, 16'd45407, 16'd9179, 16'd9281, 16'd33506});
	test_expansion(128'hdef86f6b9a4e6b8478e1486652aab421, {16'd48224, 16'd23671, 16'd40997, 16'd20263, 16'd42845, 16'd8713, 16'd10807, 16'd17676, 16'd16474, 16'd52423, 16'd21962, 16'd26499, 16'd55315, 16'd41371, 16'd60556, 16'd10346, 16'd54517, 16'd3747, 16'd61835, 16'd47955, 16'd54726, 16'd1329, 16'd19715, 16'd42910, 16'd29285, 16'd52734});
	test_expansion(128'hea4d740aeb3442204b883fdd18547824, {16'd52777, 16'd5540, 16'd63214, 16'd26401, 16'd65444, 16'd17783, 16'd51341, 16'd15910, 16'd30445, 16'd7251, 16'd20429, 16'd26601, 16'd50253, 16'd25071, 16'd9952, 16'd54818, 16'd58373, 16'd46576, 16'd7116, 16'd45969, 16'd18099, 16'd40184, 16'd46384, 16'd51420, 16'd61105, 16'd27368});
	test_expansion(128'h458eb93fa0f8b8db4e74aee11ad808d1, {16'd38182, 16'd44799, 16'd37712, 16'd10792, 16'd10845, 16'd54426, 16'd60757, 16'd30564, 16'd43001, 16'd40137, 16'd24332, 16'd8218, 16'd1881, 16'd58234, 16'd29877, 16'd5593, 16'd58966, 16'd12734, 16'd58575, 16'd28842, 16'd34062, 16'd43875, 16'd60854, 16'd62486, 16'd23407, 16'd43698});
	test_expansion(128'h2de0a79874537104b2e8e07c5027a588, {16'd55353, 16'd29899, 16'd24301, 16'd47680, 16'd8877, 16'd19008, 16'd19092, 16'd50492, 16'd5071, 16'd58084, 16'd57079, 16'd17389, 16'd24729, 16'd37284, 16'd48886, 16'd31883, 16'd53697, 16'd29170, 16'd32533, 16'd3283, 16'd26407, 16'd28960, 16'd44164, 16'd53444, 16'd54121, 16'd45884});
	test_expansion(128'h1924a171310b06c2c82891db9974b76d, {16'd14382, 16'd6626, 16'd47282, 16'd16854, 16'd37480, 16'd51447, 16'd63498, 16'd42281, 16'd32435, 16'd18170, 16'd28470, 16'd39306, 16'd3670, 16'd314, 16'd62621, 16'd59109, 16'd41259, 16'd51657, 16'd7638, 16'd43129, 16'd56550, 16'd64784, 16'd64252, 16'd44322, 16'd55848, 16'd44827});
	test_expansion(128'h64e5d3fc8d5bc9cd2f51a6f25c315f2f, {16'd15657, 16'd44494, 16'd18559, 16'd1593, 16'd41242, 16'd428, 16'd59323, 16'd34787, 16'd4121, 16'd57011, 16'd39758, 16'd42724, 16'd50666, 16'd41216, 16'd59943, 16'd61753, 16'd62822, 16'd16191, 16'd33767, 16'd24045, 16'd9640, 16'd3103, 16'd22713, 16'd32316, 16'd36270, 16'd2672});
	test_expansion(128'h2fa8bdea09b21b7872378870e0482500, {16'd5298, 16'd20689, 16'd47526, 16'd685, 16'd33808, 16'd1589, 16'd20018, 16'd34895, 16'd33982, 16'd56200, 16'd23518, 16'd39096, 16'd1485, 16'd14256, 16'd31678, 16'd33424, 16'd42465, 16'd37992, 16'd9473, 16'd45333, 16'd1959, 16'd32889, 16'd5969, 16'd8528, 16'd45320, 16'd36914});
	test_expansion(128'h6ff4ad7a13b655d602762496481fbb5e, {16'd13132, 16'd61875, 16'd39138, 16'd35421, 16'd23235, 16'd8439, 16'd8998, 16'd60807, 16'd60446, 16'd65273, 16'd59835, 16'd29552, 16'd37338, 16'd31677, 16'd62540, 16'd18439, 16'd34538, 16'd27704, 16'd57276, 16'd38299, 16'd46719, 16'd61263, 16'd11014, 16'd43921, 16'd50247, 16'd3283});
	test_expansion(128'hbce159388b64b8da9390a1d39132c592, {16'd5104, 16'd6201, 16'd39661, 16'd5891, 16'd23043, 16'd56698, 16'd40310, 16'd64574, 16'd60556, 16'd52057, 16'd29590, 16'd48447, 16'd3797, 16'd12738, 16'd32736, 16'd15735, 16'd58529, 16'd1968, 16'd49519, 16'd6739, 16'd49290, 16'd46447, 16'd15771, 16'd65450, 16'd29542, 16'd45888});
	test_expansion(128'h03622fc6cb8f8016e178506a6e4cd3e3, {16'd1361, 16'd5662, 16'd29593, 16'd19818, 16'd45397, 16'd36265, 16'd6787, 16'd37334, 16'd33498, 16'd1321, 16'd40520, 16'd39271, 16'd9441, 16'd43016, 16'd48146, 16'd60852, 16'd44464, 16'd50595, 16'd47003, 16'd44807, 16'd61846, 16'd11588, 16'd8771, 16'd9325, 16'd44564, 16'd18744});
	test_expansion(128'hc583bfe552b36248963cfd8f5e2f579a, {16'd47741, 16'd39692, 16'd32584, 16'd44423, 16'd18277, 16'd12998, 16'd5081, 16'd49496, 16'd29823, 16'd29259, 16'd7607, 16'd41426, 16'd54403, 16'd21902, 16'd21828, 16'd30309, 16'd4301, 16'd22864, 16'd54798, 16'd56247, 16'd60338, 16'd48854, 16'd18530, 16'd8881, 16'd45184, 16'd6901});
	test_expansion(128'hb3ac406c8208a844a2c254c8b6988aa2, {16'd30145, 16'd9501, 16'd22410, 16'd44581, 16'd9771, 16'd7887, 16'd1024, 16'd7202, 16'd18485, 16'd27816, 16'd45788, 16'd45079, 16'd56196, 16'd30558, 16'd50642, 16'd51043, 16'd57571, 16'd29109, 16'd6373, 16'd27495, 16'd33054, 16'd31096, 16'd42346, 16'd56728, 16'd26645, 16'd33874});
	test_expansion(128'h63aed749eb42ce51d72f9985dc35e04e, {16'd40206, 16'd7476, 16'd27852, 16'd34498, 16'd39739, 16'd7966, 16'd61385, 16'd16931, 16'd39545, 16'd10369, 16'd32515, 16'd13022, 16'd63495, 16'd34466, 16'd44446, 16'd11539, 16'd63028, 16'd41452, 16'd19101, 16'd51385, 16'd5983, 16'd34109, 16'd568, 16'd44871, 16'd35980, 16'd17854});
	test_expansion(128'hd8188a3def12d24f0b0a7cabf721148e, {16'd14950, 16'd34158, 16'd9219, 16'd36219, 16'd37104, 16'd27725, 16'd57379, 16'd17245, 16'd62656, 16'd10287, 16'd44109, 16'd14356, 16'd25319, 16'd17639, 16'd25058, 16'd53580, 16'd58688, 16'd21368, 16'd12153, 16'd54702, 16'd50010, 16'd24067, 16'd15715, 16'd57243, 16'd5687, 16'd39757});
	test_expansion(128'heb0d0157756bc0842f7dd5aa9ce21c6e, {16'd55806, 16'd28296, 16'd16568, 16'd37174, 16'd58469, 16'd35766, 16'd57708, 16'd40544, 16'd48757, 16'd27149, 16'd18889, 16'd32467, 16'd9960, 16'd52028, 16'd21380, 16'd46463, 16'd19789, 16'd4483, 16'd39940, 16'd800, 16'd35766, 16'd54243, 16'd39022, 16'd3706, 16'd50831, 16'd30137});
	test_expansion(128'hf162e70b6b22455cc5d93d139a473698, {16'd62048, 16'd41484, 16'd958, 16'd7592, 16'd14876, 16'd10064, 16'd64588, 16'd18257, 16'd63728, 16'd62620, 16'd5118, 16'd15346, 16'd8329, 16'd49020, 16'd5823, 16'd61262, 16'd43684, 16'd29322, 16'd24382, 16'd54053, 16'd25184, 16'd60441, 16'd42819, 16'd34415, 16'd22644, 16'd16447});
	test_expansion(128'hb272b6eea51dfcc083733347f1ea5816, {16'd14712, 16'd63633, 16'd39962, 16'd17924, 16'd35345, 16'd25852, 16'd10789, 16'd19249, 16'd56129, 16'd22947, 16'd17129, 16'd52235, 16'd27985, 16'd39157, 16'd48202, 16'd54975, 16'd64793, 16'd10229, 16'd50076, 16'd3113, 16'd25280, 16'd23317, 16'd23304, 16'd6199, 16'd60500, 16'd30220});
	test_expansion(128'h32f31ff14820d1b951571b0495970229, {16'd57070, 16'd10898, 16'd33664, 16'd21236, 16'd30926, 16'd30842, 16'd34651, 16'd25701, 16'd22984, 16'd5849, 16'd2580, 16'd59204, 16'd7930, 16'd60191, 16'd45002, 16'd4231, 16'd15513, 16'd39574, 16'd18147, 16'd12489, 16'd39681, 16'd26825, 16'd27996, 16'd5360, 16'd22498, 16'd30883});
	test_expansion(128'ha6302425bbce2813f1575763a4ae94ac, {16'd54710, 16'd47088, 16'd1137, 16'd56049, 16'd60275, 16'd45733, 16'd62590, 16'd25903, 16'd14970, 16'd45564, 16'd13698, 16'd32523, 16'd49181, 16'd42418, 16'd21470, 16'd33566, 16'd57345, 16'd40927, 16'd13519, 16'd34238, 16'd51300, 16'd41210, 16'd33738, 16'd6150, 16'd19168, 16'd36185});
	test_expansion(128'h5ffea9c17f42319d5266553fcd3de9cc, {16'd21223, 16'd60216, 16'd26645, 16'd27713, 16'd7776, 16'd59053, 16'd3756, 16'd64448, 16'd1083, 16'd17776, 16'd42558, 16'd23446, 16'd45539, 16'd33059, 16'd31501, 16'd5568, 16'd47260, 16'd27226, 16'd11970, 16'd17695, 16'd12777, 16'd48181, 16'd41396, 16'd57079, 16'd22865, 16'd37146});
	test_expansion(128'hd5b2f65ec7b05fd32a81428e097f797c, {16'd28657, 16'd6222, 16'd9282, 16'd289, 16'd63842, 16'd25531, 16'd380, 16'd7368, 16'd16527, 16'd29980, 16'd31439, 16'd9865, 16'd36398, 16'd39871, 16'd56025, 16'd37032, 16'd33885, 16'd12909, 16'd3503, 16'd19261, 16'd63111, 16'd61430, 16'd57604, 16'd54633, 16'd43465, 16'd48021});
	test_expansion(128'hed2c10350dbdbd9c0ff2b88c0bbb9a29, {16'd17751, 16'd4478, 16'd9972, 16'd25572, 16'd3469, 16'd24600, 16'd6187, 16'd46368, 16'd9093, 16'd53962, 16'd8234, 16'd42000, 16'd65232, 16'd53867, 16'd32620, 16'd648, 16'd46688, 16'd1946, 16'd28288, 16'd39110, 16'd8273, 16'd9461, 16'd25752, 16'd25319, 16'd19919, 16'd53565});
	test_expansion(128'h3522c802420af264db5006368c4896fc, {16'd52940, 16'd1903, 16'd10836, 16'd10929, 16'd31848, 16'd13445, 16'd23024, 16'd33548, 16'd64850, 16'd25017, 16'd32940, 16'd34103, 16'd2092, 16'd36829, 16'd1047, 16'd63294, 16'd64076, 16'd65098, 16'd37690, 16'd17770, 16'd14091, 16'd22686, 16'd61301, 16'd20595, 16'd38897, 16'd45709});
	test_expansion(128'hdc3905afe107ec2f93e66169bd37598e, {16'd27171, 16'd13713, 16'd2560, 16'd23261, 16'd58845, 16'd51433, 16'd39274, 16'd32752, 16'd5213, 16'd25759, 16'd19554, 16'd63498, 16'd48263, 16'd18131, 16'd5233, 16'd38441, 16'd46415, 16'd50316, 16'd48431, 16'd59045, 16'd41725, 16'd15858, 16'd12400, 16'd30585, 16'd50400, 16'd10743});
	test_expansion(128'hb056ddad549e80fec989f4a9c490517c, {16'd65461, 16'd6814, 16'd63760, 16'd20547, 16'd49841, 16'd53902, 16'd38192, 16'd7182, 16'd22683, 16'd59256, 16'd52988, 16'd20470, 16'd10063, 16'd9452, 16'd16420, 16'd24278, 16'd7870, 16'd49574, 16'd19664, 16'd21699, 16'd30037, 16'd2340, 16'd20765, 16'd35488, 16'd47784, 16'd45937});
	test_expansion(128'hfd56f5b975c14ab00590c789bee23587, {16'd18781, 16'd45483, 16'd13516, 16'd19148, 16'd65194, 16'd45880, 16'd23648, 16'd15423, 16'd33561, 16'd5110, 16'd51250, 16'd62141, 16'd61183, 16'd39102, 16'd34284, 16'd47193, 16'd57281, 16'd59774, 16'd55896, 16'd45805, 16'd22274, 16'd37918, 16'd16971, 16'd26138, 16'd48504, 16'd55342});
	test_expansion(128'h2ccc6de7c8e5e63fe821388f53bf42b2, {16'd24538, 16'd53879, 16'd28905, 16'd60765, 16'd18078, 16'd42472, 16'd44422, 16'd61996, 16'd24682, 16'd20218, 16'd31595, 16'd31309, 16'd53461, 16'd55545, 16'd56745, 16'd51611, 16'd40883, 16'd37713, 16'd4307, 16'd17512, 16'd53899, 16'd47757, 16'd28095, 16'd63708, 16'd32085, 16'd43340});
	test_expansion(128'hf55ef142cc181cdb9b32d243ade74fae, {16'd49280, 16'd27945, 16'd5004, 16'd52340, 16'd37553, 16'd52869, 16'd57041, 16'd15697, 16'd56657, 16'd27651, 16'd5173, 16'd53677, 16'd13978, 16'd60468, 16'd34781, 16'd34526, 16'd58680, 16'd14181, 16'd46281, 16'd19639, 16'd59990, 16'd61185, 16'd29161, 16'd58312, 16'd16563, 16'd24841});
	test_expansion(128'hd32e3805b6137f75b2971a24f28a8a6f, {16'd10252, 16'd4429, 16'd24984, 16'd40028, 16'd60973, 16'd12712, 16'd12032, 16'd37373, 16'd8119, 16'd62039, 16'd24900, 16'd11810, 16'd52591, 16'd35151, 16'd8564, 16'd33922, 16'd36575, 16'd53200, 16'd9576, 16'd43618, 16'd23768, 16'd14553, 16'd64896, 16'd13784, 16'd27907, 16'd47485});
	test_expansion(128'h0c1221359f12f360d82c8cdc87d89617, {16'd47739, 16'd17976, 16'd6647, 16'd30717, 16'd49117, 16'd55770, 16'd31834, 16'd38151, 16'd768, 16'd5429, 16'd30012, 16'd57328, 16'd26594, 16'd53248, 16'd36146, 16'd53122, 16'd33781, 16'd3223, 16'd18481, 16'd61824, 16'd16796, 16'd33717, 16'd24572, 16'd20238, 16'd41235, 16'd25057});
	test_expansion(128'ha5779620f1c1ca5b2a1b96c533a7af94, {16'd37110, 16'd45089, 16'd41950, 16'd38494, 16'd1846, 16'd49320, 16'd41113, 16'd55532, 16'd41047, 16'd25036, 16'd1665, 16'd54216, 16'd12480, 16'd36195, 16'd3613, 16'd12959, 16'd34174, 16'd43560, 16'd16601, 16'd10354, 16'd42377, 16'd7566, 16'd54165, 16'd20186, 16'd55905, 16'd63666});
	test_expansion(128'ha626f6843a23acfeb1c21ce352ba6d6c, {16'd41198, 16'd3984, 16'd45217, 16'd51403, 16'd55209, 16'd18152, 16'd36967, 16'd22727, 16'd47955, 16'd23003, 16'd46367, 16'd49729, 16'd30534, 16'd49435, 16'd49722, 16'd5785, 16'd12754, 16'd27538, 16'd1215, 16'd39829, 16'd20525, 16'd39427, 16'd36525, 16'd63172, 16'd54642, 16'd53999});
	test_expansion(128'h99e07eb6da5117986bd819b03143f179, {16'd8234, 16'd2481, 16'd26378, 16'd52718, 16'd10619, 16'd55606, 16'd5032, 16'd29857, 16'd60007, 16'd43110, 16'd50287, 16'd26103, 16'd26630, 16'd12179, 16'd31432, 16'd25795, 16'd36371, 16'd59226, 16'd56463, 16'd46507, 16'd29938, 16'd47726, 16'd25878, 16'd43762, 16'd29953, 16'd32002});
	test_expansion(128'h41c132992ac7616709551965ee5d6c46, {16'd52414, 16'd48103, 16'd39986, 16'd39102, 16'd38787, 16'd18070, 16'd59714, 16'd24977, 16'd8859, 16'd48390, 16'd22785, 16'd15921, 16'd57168, 16'd40204, 16'd29772, 16'd32411, 16'd39948, 16'd17753, 16'd2883, 16'd58142, 16'd27263, 16'd17622, 16'd12344, 16'd16551, 16'd14709, 16'd3061});
	test_expansion(128'he599fea739cab612ee3d609a8c6029d6, {16'd64470, 16'd12105, 16'd28723, 16'd6204, 16'd15126, 16'd61117, 16'd1458, 16'd35437, 16'd48135, 16'd19901, 16'd21970, 16'd35221, 16'd18715, 16'd187, 16'd4422, 16'd23989, 16'd5991, 16'd44994, 16'd36766, 16'd1144, 16'd21307, 16'd42967, 16'd44521, 16'd36443, 16'd52523, 16'd32561});
	test_expansion(128'h47c0d4c89477a35f8945644e463f450d, {16'd42706, 16'd47694, 16'd10153, 16'd50932, 16'd53159, 16'd34293, 16'd43112, 16'd62170, 16'd60991, 16'd2406, 16'd24487, 16'd64712, 16'd51440, 16'd10456, 16'd22019, 16'd2995, 16'd29190, 16'd34383, 16'd4248, 16'd44682, 16'd20716, 16'd3085, 16'd40156, 16'd21796, 16'd65483, 16'd62912});
	test_expansion(128'h7884cae4534dd149eade1631076bdf1d, {16'd46705, 16'd26657, 16'd64943, 16'd19479, 16'd46526, 16'd31363, 16'd10711, 16'd30915, 16'd35504, 16'd62824, 16'd50150, 16'd32643, 16'd15265, 16'd26003, 16'd56365, 16'd39724, 16'd49018, 16'd28420, 16'd55391, 16'd40865, 16'd29075, 16'd9520, 16'd25092, 16'd46881, 16'd575, 16'd62329});
	test_expansion(128'hb9d0d6bd300c0d03fd4314dc2aa8d537, {16'd32279, 16'd55784, 16'd9962, 16'd2363, 16'd38185, 16'd8590, 16'd3356, 16'd37545, 16'd55658, 16'd33723, 16'd44795, 16'd53385, 16'd33886, 16'd33536, 16'd4889, 16'd37278, 16'd26415, 16'd29641, 16'd30225, 16'd24134, 16'd31065, 16'd56594, 16'd21, 16'd21676, 16'd44187, 16'd56125});
	test_expansion(128'h659bd9b44d03c540ed494fe07b36f57c, {16'd30724, 16'd43365, 16'd47635, 16'd48124, 16'd46618, 16'd24864, 16'd54609, 16'd6783, 16'd54056, 16'd15359, 16'd53357, 16'd35054, 16'd2846, 16'd4731, 16'd17127, 16'd27118, 16'd1978, 16'd61672, 16'd29772, 16'd22417, 16'd48916, 16'd6406, 16'd57166, 16'd38088, 16'd47602, 16'd25577});
	test_expansion(128'hd3aa882ff84c151f77d7b9398d7a75de, {16'd27520, 16'd34899, 16'd2323, 16'd63498, 16'd14094, 16'd53922, 16'd11725, 16'd51818, 16'd62377, 16'd39581, 16'd39525, 16'd1641, 16'd9772, 16'd14419, 16'd595, 16'd10566, 16'd38618, 16'd58796, 16'd12076, 16'd2901, 16'd50495, 16'd45196, 16'd30961, 16'd65471, 16'd46607, 16'd3572});
	test_expansion(128'h9f49d0a2de828f05f5f227d918de217a, {16'd44052, 16'd51245, 16'd35308, 16'd18472, 16'd34028, 16'd43558, 16'd55169, 16'd18210, 16'd7928, 16'd8788, 16'd63875, 16'd38251, 16'd22174, 16'd35578, 16'd10202, 16'd49032, 16'd29987, 16'd26344, 16'd59257, 16'd2696, 16'd20197, 16'd57903, 16'd59328, 16'd32968, 16'd44785, 16'd64300});
	test_expansion(128'h6469f5ebf2999c30bf03cdda71564393, {16'd61767, 16'd4422, 16'd1832, 16'd60775, 16'd47645, 16'd296, 16'd1502, 16'd43922, 16'd18620, 16'd23994, 16'd26121, 16'd10552, 16'd47565, 16'd37686, 16'd37578, 16'd33405, 16'd452, 16'd15908, 16'd35951, 16'd19953, 16'd47176, 16'd58947, 16'd59656, 16'd11468, 16'd4231, 16'd26442});
	test_expansion(128'hb10d70dcede9eb955c18fd2ff73c6eed, {16'd53850, 16'd29771, 16'd25104, 16'd19839, 16'd55568, 16'd56003, 16'd33991, 16'd30585, 16'd13283, 16'd19550, 16'd15428, 16'd12024, 16'd39004, 16'd43886, 16'd44882, 16'd11443, 16'd50020, 16'd41728, 16'd12583, 16'd60422, 16'd60541, 16'd35522, 16'd43252, 16'd63479, 16'd25164, 16'd12757});
	test_expansion(128'h16645049f722c08fe92c55164388d26c, {16'd53841, 16'd57235, 16'd21312, 16'd61269, 16'd19733, 16'd6376, 16'd42550, 16'd38414, 16'd36988, 16'd54705, 16'd9528, 16'd32821, 16'd41430, 16'd31236, 16'd50183, 16'd30599, 16'd14515, 16'd39910, 16'd22026, 16'd15027, 16'd28992, 16'd54175, 16'd11458, 16'd42994, 16'd28373, 16'd58326});
	test_expansion(128'h01a37f4580d940113c485ccb16e99016, {16'd29726, 16'd60533, 16'd39250, 16'd34319, 16'd3597, 16'd4499, 16'd57730, 16'd9020, 16'd31180, 16'd24101, 16'd9616, 16'd43867, 16'd48504, 16'd18529, 16'd19915, 16'd49493, 16'd41298, 16'd52345, 16'd12375, 16'd20460, 16'd27119, 16'd12374, 16'd63713, 16'd13805, 16'd49858, 16'd14126});
	test_expansion(128'ha7683f5063f398ebeee618a5c288779b, {16'd7776, 16'd34445, 16'd38593, 16'd8477, 16'd46570, 16'd31231, 16'd56198, 16'd62680, 16'd42479, 16'd51458, 16'd11529, 16'd35510, 16'd29540, 16'd51371, 16'd10386, 16'd32672, 16'd61658, 16'd6364, 16'd47779, 16'd50085, 16'd35090, 16'd25015, 16'd1764, 16'd31109, 16'd17420, 16'd56542});
	test_expansion(128'h88c5458de63808033e00f8f7056b5977, {16'd48242, 16'd55263, 16'd54179, 16'd4771, 16'd56233, 16'd45633, 16'd9404, 16'd50590, 16'd38245, 16'd1977, 16'd29629, 16'd30622, 16'd27247, 16'd20823, 16'd29112, 16'd7455, 16'd19347, 16'd37212, 16'd53279, 16'd55671, 16'd50794, 16'd15616, 16'd31518, 16'd5160, 16'd28467, 16'd61830});
	test_expansion(128'h221af9c660435364a2ea6da79cc7c5e9, {16'd51640, 16'd15474, 16'd728, 16'd59303, 16'd8334, 16'd28795, 16'd48401, 16'd13893, 16'd10247, 16'd50951, 16'd34919, 16'd38749, 16'd59556, 16'd4646, 16'd44856, 16'd41267, 16'd61026, 16'd32798, 16'd17551, 16'd52463, 16'd62490, 16'd41085, 16'd55298, 16'd24347, 16'd28722, 16'd5469});
	test_expansion(128'h84ed611a567fb9d4092bb2c70c1e1f63, {16'd61763, 16'd17256, 16'd54015, 16'd23021, 16'd2265, 16'd42197, 16'd27321, 16'd6834, 16'd32554, 16'd9418, 16'd52960, 16'd60309, 16'd48456, 16'd28598, 16'd37652, 16'd58269, 16'd9341, 16'd40026, 16'd5130, 16'd43895, 16'd11963, 16'd40500, 16'd58411, 16'd24176, 16'd38148, 16'd10314});
	test_expansion(128'h7b65af92224b525e97c8006807e0ae19, {16'd5757, 16'd41522, 16'd28317, 16'd4571, 16'd25768, 16'd10114, 16'd22504, 16'd48221, 16'd35699, 16'd59952, 16'd32926, 16'd2965, 16'd27311, 16'd2905, 16'd35366, 16'd40639, 16'd55187, 16'd9606, 16'd62476, 16'd30111, 16'd21157, 16'd25311, 16'd20102, 16'd42885, 16'd22200, 16'd8534});
	test_expansion(128'hd139926d4fa4b2005047d17f346d6933, {16'd12198, 16'd61815, 16'd26613, 16'd29458, 16'd36457, 16'd65341, 16'd33528, 16'd31806, 16'd62516, 16'd1712, 16'd28984, 16'd35219, 16'd9260, 16'd22595, 16'd62748, 16'd14575, 16'd63387, 16'd24901, 16'd59929, 16'd527, 16'd12233, 16'd11434, 16'd8612, 16'd41543, 16'd22099, 16'd11180});
	test_expansion(128'h5af8723a8371ba41e758a05876322e94, {16'd54056, 16'd9647, 16'd38456, 16'd34718, 16'd47418, 16'd59110, 16'd21770, 16'd53415, 16'd56427, 16'd17399, 16'd6122, 16'd2587, 16'd63797, 16'd48325, 16'd54579, 16'd18599, 16'd1936, 16'd44447, 16'd41486, 16'd3408, 16'd2891, 16'd34265, 16'd4519, 16'd18539, 16'd19731, 16'd23657});
	test_expansion(128'h073becab5bc8cf7c561c78b175bf7f14, {16'd29309, 16'd11937, 16'd14153, 16'd31887, 16'd64810, 16'd43111, 16'd62008, 16'd41515, 16'd61237, 16'd62409, 16'd23031, 16'd39733, 16'd51818, 16'd50435, 16'd34078, 16'd53059, 16'd21769, 16'd7844, 16'd56985, 16'd15302, 16'd44070, 16'd40075, 16'd48082, 16'd51625, 16'd13090, 16'd35020});
	test_expansion(128'h1abda5715ca3f9b42b56b0341593cb33, {16'd1551, 16'd58959, 16'd43069, 16'd57247, 16'd32740, 16'd61143, 16'd40679, 16'd11491, 16'd1165, 16'd16057, 16'd65349, 16'd51865, 16'd55298, 16'd5980, 16'd6554, 16'd32640, 16'd4737, 16'd57627, 16'd61324, 16'd53248, 16'd11497, 16'd3908, 16'd1846, 16'd17029, 16'd21078, 16'd7414});
	test_expansion(128'h0f446235da6ffd1ab0d9335e04b74c11, {16'd55758, 16'd55067, 16'd64126, 16'd34140, 16'd46669, 16'd58133, 16'd58737, 16'd24515, 16'd43070, 16'd34629, 16'd14142, 16'd31841, 16'd40895, 16'd31366, 16'd28736, 16'd65397, 16'd39089, 16'd1024, 16'd57698, 16'd44552, 16'd47755, 16'd24961, 16'd47360, 16'd468, 16'd9007, 16'd37033});
	test_expansion(128'hdf93dc34f9acf3d54e6367a3d85181b0, {16'd1174, 16'd12745, 16'd41174, 16'd64405, 16'd39633, 16'd25753, 16'd36139, 16'd8489, 16'd23321, 16'd46857, 16'd28011, 16'd10108, 16'd29451, 16'd21862, 16'd35183, 16'd41295, 16'd20311, 16'd4869, 16'd2154, 16'd40078, 16'd13409, 16'd50862, 16'd42924, 16'd49249, 16'd45631, 16'd38470});
	test_expansion(128'hbdece9cdf667adc85d63bdeb39f4dcdf, {16'd28698, 16'd46035, 16'd2064, 16'd22264, 16'd36894, 16'd29970, 16'd45533, 16'd39346, 16'd14010, 16'd10196, 16'd56682, 16'd33189, 16'd48452, 16'd19294, 16'd34637, 16'd19310, 16'd13294, 16'd62907, 16'd3789, 16'd50124, 16'd42016, 16'd11061, 16'd11551, 16'd41364, 16'd56407, 16'd29503});
	test_expansion(128'h8981d0a1011b182894a60a9e0cdbe178, {16'd42773, 16'd39384, 16'd42705, 16'd56978, 16'd21255, 16'd13741, 16'd55441, 16'd39456, 16'd52035, 16'd60835, 16'd47242, 16'd10865, 16'd43673, 16'd3125, 16'd23486, 16'd18787, 16'd62440, 16'd58552, 16'd58616, 16'd24581, 16'd14031, 16'd63879, 16'd49878, 16'd46569, 16'd36346, 16'd18642});
	test_expansion(128'h89a8a3c8ffa197ac398d7f6b9e4f77c2, {16'd8919, 16'd60872, 16'd34178, 16'd4335, 16'd3002, 16'd14534, 16'd60895, 16'd13796, 16'd23584, 16'd12522, 16'd154, 16'd29143, 16'd24246, 16'd57099, 16'd50776, 16'd25502, 16'd22556, 16'd61913, 16'd50089, 16'd58129, 16'd30688, 16'd39125, 16'd15153, 16'd31794, 16'd44470, 16'd39231});
	test_expansion(128'h4bd97d08deaea413ea9e87746e615415, {16'd48195, 16'd59810, 16'd5080, 16'd38345, 16'd63000, 16'd47854, 16'd51090, 16'd63705, 16'd32861, 16'd12906, 16'd43265, 16'd36344, 16'd10648, 16'd24545, 16'd28389, 16'd61317, 16'd5152, 16'd31910, 16'd63700, 16'd58067, 16'd59695, 16'd33368, 16'd32336, 16'd26637, 16'd54280, 16'd36474});
	test_expansion(128'h3e90328d3b2b24eca3871203e3b18dac, {16'd50534, 16'd30281, 16'd35100, 16'd44121, 16'd31481, 16'd8852, 16'd41616, 16'd20394, 16'd23498, 16'd29522, 16'd44454, 16'd35068, 16'd49976, 16'd27023, 16'd24967, 16'd22150, 16'd22435, 16'd2458, 16'd1257, 16'd37986, 16'd63478, 16'd19216, 16'd36724, 16'd10652, 16'd39335, 16'd43204});
	test_expansion(128'ha77cb4b0c35071942e6efdcdccd6592d, {16'd24037, 16'd3670, 16'd61506, 16'd18146, 16'd62910, 16'd6751, 16'd24551, 16'd47302, 16'd57979, 16'd29226, 16'd41222, 16'd37802, 16'd52509, 16'd37082, 16'd12453, 16'd415, 16'd51976, 16'd47806, 16'd53296, 16'd39156, 16'd18610, 16'd60264, 16'd45462, 16'd34274, 16'd37752, 16'd61382});
	test_expansion(128'hcc945a9a20be5963f5a767dd60b6a097, {16'd29395, 16'd11231, 16'd29688, 16'd30003, 16'd904, 16'd39389, 16'd32035, 16'd22858, 16'd21728, 16'd13550, 16'd41614, 16'd17825, 16'd29876, 16'd28676, 16'd50458, 16'd31391, 16'd38302, 16'd39978, 16'd5769, 16'd13148, 16'd28070, 16'd43289, 16'd44296, 16'd36458, 16'd29491, 16'd26516});
	test_expansion(128'hfacb7f89b5bd5e200d9213ef18530e23, {16'd46893, 16'd50453, 16'd61872, 16'd28485, 16'd54407, 16'd2497, 16'd4853, 16'd5309, 16'd39537, 16'd36511, 16'd63171, 16'd46594, 16'd59766, 16'd25084, 16'd39556, 16'd39182, 16'd63578, 16'd48998, 16'd46305, 16'd41317, 16'd36608, 16'd36032, 16'd3839, 16'd3457, 16'd60537, 16'd64520});
	test_expansion(128'heb9ae9908b84b67e2de0116cc38224ea, {16'd55218, 16'd33000, 16'd16976, 16'd33829, 16'd7434, 16'd46356, 16'd13054, 16'd62960, 16'd25512, 16'd43901, 16'd37112, 16'd2268, 16'd58271, 16'd24543, 16'd33187, 16'd27753, 16'd1271, 16'd50740, 16'd25069, 16'd16351, 16'd20191, 16'd41177, 16'd20960, 16'd18692, 16'd1272, 16'd38420});
	test_expansion(128'h13816566d0f842d175bf5872826b54e2, {16'd44149, 16'd8049, 16'd48619, 16'd52678, 16'd62519, 16'd53352, 16'd31942, 16'd3703, 16'd1819, 16'd38645, 16'd59006, 16'd27308, 16'd22515, 16'd26938, 16'd6938, 16'd61223, 16'd637, 16'd43044, 16'd49761, 16'd64614, 16'd6272, 16'd56516, 16'd21296, 16'd9237, 16'd15826, 16'd63742});
	test_expansion(128'h154439076f5c4e6845730fe6e193d125, {16'd31543, 16'd6682, 16'd40131, 16'd40207, 16'd51385, 16'd62859, 16'd20115, 16'd31221, 16'd10723, 16'd25776, 16'd49420, 16'd42270, 16'd35730, 16'd39994, 16'd44625, 16'd60169, 16'd35680, 16'd60283, 16'd35627, 16'd55945, 16'd21908, 16'd35644, 16'd6737, 16'd4730, 16'd64991, 16'd58838});
	test_expansion(128'hd94ddb54cebebf44e6f8ab89e1234759, {16'd29707, 16'd40263, 16'd49073, 16'd61918, 16'd4469, 16'd25088, 16'd15694, 16'd30615, 16'd39376, 16'd25281, 16'd57570, 16'd4766, 16'd28741, 16'd11223, 16'd31788, 16'd22215, 16'd27737, 16'd27741, 16'd54009, 16'd3871, 16'd52327, 16'd60424, 16'd34890, 16'd48516, 16'd6750, 16'd15349});
	test_expansion(128'h569e2c6fec016814249c042e85a261a1, {16'd38916, 16'd56247, 16'd65013, 16'd56303, 16'd40438, 16'd15608, 16'd43744, 16'd55058, 16'd14960, 16'd11535, 16'd57173, 16'd3758, 16'd63566, 16'd60356, 16'd32771, 16'd52963, 16'd58296, 16'd61740, 16'd34371, 16'd31144, 16'd53689, 16'd59276, 16'd19509, 16'd36773, 16'd10629, 16'd39550});
	test_expansion(128'h3cd8b89b0ff0200ad862f42bbc6d59e5, {16'd21156, 16'd16086, 16'd930, 16'd19919, 16'd32113, 16'd39454, 16'd25701, 16'd11319, 16'd8326, 16'd11787, 16'd15722, 16'd33559, 16'd2125, 16'd44960, 16'd38669, 16'd25394, 16'd5958, 16'd14222, 16'd22572, 16'd20267, 16'd2268, 16'd45642, 16'd7821, 16'd14215, 16'd27718, 16'd40690});
	test_expansion(128'h58714ff901833296bbe1ca8f36a4a2d9, {16'd40669, 16'd24735, 16'd24345, 16'd20399, 16'd36645, 16'd29741, 16'd13713, 16'd1667, 16'd40763, 16'd34811, 16'd8189, 16'd34023, 16'd5430, 16'd6991, 16'd61933, 16'd53551, 16'd9461, 16'd25100, 16'd3877, 16'd18066, 16'd6833, 16'd48258, 16'd13540, 16'd3082, 16'd52096, 16'd32521});
	test_expansion(128'he7d043c5dd3bf875b58cd70aaf40bb9b, {16'd52699, 16'd64823, 16'd33067, 16'd34003, 16'd36185, 16'd3139, 16'd17930, 16'd14475, 16'd58171, 16'd27997, 16'd29981, 16'd50909, 16'd45920, 16'd46287, 16'd36265, 16'd57007, 16'd19973, 16'd43321, 16'd8906, 16'd37872, 16'd53978, 16'd16974, 16'd56572, 16'd63289, 16'd36786, 16'd1529});
	test_expansion(128'h77731ccbdb460259b420febe9da587c1, {16'd30522, 16'd37771, 16'd60487, 16'd63120, 16'd7880, 16'd17606, 16'd20226, 16'd11174, 16'd27856, 16'd10769, 16'd31717, 16'd32586, 16'd13800, 16'd6737, 16'd17554, 16'd1898, 16'd42279, 16'd56485, 16'd45808, 16'd59647, 16'd42422, 16'd8, 16'd46251, 16'd25322, 16'd32778, 16'd12846});
	test_expansion(128'ha68ea97aa98b11290561a757cc746ba7, {16'd53420, 16'd10776, 16'd27231, 16'd23964, 16'd58729, 16'd49779, 16'd18995, 16'd481, 16'd55320, 16'd23881, 16'd37785, 16'd22013, 16'd38652, 16'd51076, 16'd37062, 16'd19827, 16'd7504, 16'd15708, 16'd766, 16'd9938, 16'd50954, 16'd12696, 16'd20292, 16'd12772, 16'd35821, 16'd36073});
	test_expansion(128'h736f304b1104e66fdc2d3b9b93d8accf, {16'd10748, 16'd15451, 16'd16914, 16'd8959, 16'd34013, 16'd38128, 16'd621, 16'd23947, 16'd18549, 16'd43924, 16'd18101, 16'd14114, 16'd50219, 16'd59409, 16'd43629, 16'd44558, 16'd42589, 16'd25157, 16'd39515, 16'd699, 16'd34638, 16'd926, 16'd7352, 16'd41164, 16'd23562, 16'd57338});
	test_expansion(128'h889191373f23bebdf8960bc7d7c819b0, {16'd34360, 16'd13585, 16'd27077, 16'd52280, 16'd5973, 16'd38899, 16'd55248, 16'd57526, 16'd33115, 16'd2075, 16'd53050, 16'd27706, 16'd41112, 16'd60191, 16'd49700, 16'd16453, 16'd5643, 16'd11222, 16'd22135, 16'd29027, 16'd20112, 16'd33162, 16'd41042, 16'd50950, 16'd43365, 16'd23459});
	test_expansion(128'heed1e9e04938e597e1dcf00b82393f39, {16'd30010, 16'd64786, 16'd17108, 16'd49792, 16'd48235, 16'd52391, 16'd51249, 16'd39873, 16'd46, 16'd23754, 16'd5053, 16'd32515, 16'd341, 16'd62656, 16'd50026, 16'd50054, 16'd27653, 16'd45015, 16'd51720, 16'd8251, 16'd35649, 16'd28234, 16'd1863, 16'd58587, 16'd23767, 16'd3695});
	test_expansion(128'he85c9268f0cc7b51f990f646244d64b3, {16'd19484, 16'd26242, 16'd40000, 16'd40169, 16'd3692, 16'd13017, 16'd6129, 16'd30070, 16'd21004, 16'd1843, 16'd25989, 16'd62933, 16'd30178, 16'd40869, 16'd43931, 16'd61427, 16'd56778, 16'd54589, 16'd12257, 16'd10125, 16'd700, 16'd61239, 16'd2947, 16'd57947, 16'd21817, 16'd32184});
	test_expansion(128'hd897878a315be537b1aa33ea788a5ac7, {16'd48760, 16'd58640, 16'd57244, 16'd58604, 16'd59217, 16'd3692, 16'd11980, 16'd20625, 16'd40458, 16'd53130, 16'd19246, 16'd34018, 16'd30304, 16'd11296, 16'd40274, 16'd42677, 16'd49446, 16'd61380, 16'd41081, 16'd41615, 16'd39305, 16'd58288, 16'd39566, 16'd4214, 16'd42528, 16'd53134});
	test_expansion(128'hc8dfee90710c9696489d1d4f6e672349, {16'd59728, 16'd34634, 16'd36591, 16'd39554, 16'd46510, 16'd5989, 16'd36570, 16'd14546, 16'd21417, 16'd52579, 16'd56426, 16'd52004, 16'd46794, 16'd32902, 16'd56710, 16'd55024, 16'd59512, 16'd24834, 16'd27678, 16'd20373, 16'd65147, 16'd6268, 16'd5051, 16'd16678, 16'd45487, 16'd587});
	test_expansion(128'h2bc462cf610084a1035b42b52d9924e5, {16'd31358, 16'd52187, 16'd9410, 16'd58888, 16'd6982, 16'd9322, 16'd12089, 16'd9088, 16'd48730, 16'd1863, 16'd39479, 16'd55642, 16'd64275, 16'd64824, 16'd56655, 16'd21025, 16'd39559, 16'd54173, 16'd17810, 16'd28993, 16'd9934, 16'd1400, 16'd10253, 16'd26538, 16'd38543, 16'd33760});
	test_expansion(128'h1268f072d7592b109eb0dd530e6426d0, {16'd29713, 16'd40941, 16'd64363, 16'd2765, 16'd48230, 16'd13942, 16'd59082, 16'd60491, 16'd39430, 16'd1865, 16'd33589, 16'd15654, 16'd25240, 16'd5017, 16'd22696, 16'd52081, 16'd29805, 16'd9465, 16'd24224, 16'd5064, 16'd36430, 16'd13524, 16'd63230, 16'd9016, 16'd53290, 16'd40801});
	test_expansion(128'hdce78b35a92b07d61ffa525d5544272d, {16'd61723, 16'd6024, 16'd3368, 16'd35455, 16'd34844, 16'd9672, 16'd55743, 16'd25955, 16'd34712, 16'd35352, 16'd58942, 16'd40600, 16'd2024, 16'd30193, 16'd2883, 16'd32831, 16'd60697, 16'd57462, 16'd2586, 16'd61727, 16'd26385, 16'd40287, 16'd55324, 16'd65008, 16'd19740, 16'd56343});
	test_expansion(128'h7a7bd2d467acc36627961fb8f9f3b297, {16'd36883, 16'd61211, 16'd40751, 16'd18644, 16'd4624, 16'd37358, 16'd8802, 16'd16363, 16'd50655, 16'd24697, 16'd13076, 16'd55579, 16'd27265, 16'd54845, 16'd61590, 16'd41022, 16'd51614, 16'd10453, 16'd13976, 16'd24912, 16'd28926, 16'd21008, 16'd27843, 16'd31453, 16'd46864, 16'd37134});
	test_expansion(128'haf831e51604f717fbb79eaf17d091385, {16'd57169, 16'd48033, 16'd18460, 16'd52186, 16'd45511, 16'd65277, 16'd61246, 16'd2614, 16'd44665, 16'd55822, 16'd556, 16'd38927, 16'd27552, 16'd39988, 16'd49833, 16'd40419, 16'd14015, 16'd15632, 16'd22910, 16'd50938, 16'd11057, 16'd51378, 16'd50691, 16'd45400, 16'd32825, 16'd24341});
	test_expansion(128'hfd6609341efb27126248f0815e3945b4, {16'd15912, 16'd59588, 16'd21834, 16'd57904, 16'd5535, 16'd9211, 16'd42210, 16'd22297, 16'd64714, 16'd747, 16'd52393, 16'd5612, 16'd32675, 16'd31946, 16'd34438, 16'd40698, 16'd65292, 16'd46931, 16'd60667, 16'd9887, 16'd62670, 16'd7937, 16'd13244, 16'd26459, 16'd40940, 16'd62695});
	test_expansion(128'h1f4d21fa6dc2a62e07170ca0053e0adc, {16'd29967, 16'd39726, 16'd27725, 16'd30849, 16'd37300, 16'd59027, 16'd61114, 16'd43262, 16'd53876, 16'd25693, 16'd24362, 16'd41960, 16'd53442, 16'd59919, 16'd45316, 16'd36724, 16'd33786, 16'd26058, 16'd47485, 16'd49127, 16'd48373, 16'd57230, 16'd1328, 16'd2388, 16'd26104, 16'd88});
	test_expansion(128'h07ba28b52ca9de62a3d20edaa5549923, {16'd25528, 16'd41389, 16'd21908, 16'd49007, 16'd23159, 16'd21377, 16'd43569, 16'd50627, 16'd20790, 16'd63482, 16'd34358, 16'd2098, 16'd26657, 16'd36946, 16'd58285, 16'd13483, 16'd59907, 16'd40070, 16'd11646, 16'd36994, 16'd22141, 16'd44497, 16'd38810, 16'd47615, 16'd34382, 16'd7012});
	test_expansion(128'h1349535ddcb513c62f5455722892d678, {16'd29165, 16'd45720, 16'd19975, 16'd24379, 16'd38372, 16'd27681, 16'd14704, 16'd52173, 16'd29083, 16'd21521, 16'd17758, 16'd8317, 16'd20768, 16'd4180, 16'd54312, 16'd31265, 16'd33076, 16'd22555, 16'd60165, 16'd2991, 16'd52593, 16'd56345, 16'd6365, 16'd32733, 16'd61453, 16'd20127});
	test_expansion(128'hc8dc098d00fe4485be3f5b590bba1288, {16'd36711, 16'd49254, 16'd7963, 16'd60249, 16'd52969, 16'd26808, 16'd39285, 16'd36919, 16'd29736, 16'd42085, 16'd34887, 16'd35103, 16'd26159, 16'd11944, 16'd36804, 16'd57593, 16'd53095, 16'd133, 16'd6284, 16'd29215, 16'd46824, 16'd24333, 16'd34981, 16'd40760, 16'd63925, 16'd37831});
	test_expansion(128'hb7b15e54d0831c3672df899631086932, {16'd28128, 16'd16074, 16'd37981, 16'd21496, 16'd60341, 16'd17411, 16'd60343, 16'd8587, 16'd416, 16'd20541, 16'd19156, 16'd49342, 16'd18307, 16'd3179, 16'd43816, 16'd19999, 16'd49158, 16'd13796, 16'd64751, 16'd15396, 16'd24947, 16'd21048, 16'd40938, 16'd43273, 16'd31500, 16'd24857});
	test_expansion(128'h9232b1bcf74c69d999030c3f15a437fd, {16'd1691, 16'd56967, 16'd18676, 16'd1492, 16'd23268, 16'd1293, 16'd30493, 16'd13766, 16'd54795, 16'd52946, 16'd59136, 16'd10733, 16'd44694, 16'd44542, 16'd889, 16'd25231, 16'd40742, 16'd24158, 16'd59094, 16'd9805, 16'd26315, 16'd22935, 16'd49830, 16'd32918, 16'd11523, 16'd1534});
	test_expansion(128'h4064c9923ffcef7e3a2bef019fa4cf9d, {16'd28525, 16'd59174, 16'd62339, 16'd20808, 16'd34950, 16'd4409, 16'd21825, 16'd39096, 16'd34106, 16'd42543, 16'd32160, 16'd58709, 16'd55737, 16'd12746, 16'd47027, 16'd15377, 16'd59699, 16'd64836, 16'd61726, 16'd21830, 16'd44770, 16'd5470, 16'd55876, 16'd61934, 16'd16258, 16'd13615});
	test_expansion(128'h862604f883fdb65be809c38d0f1a03e5, {16'd20603, 16'd13904, 16'd25220, 16'd32838, 16'd11758, 16'd20316, 16'd61653, 16'd2097, 16'd27485, 16'd59580, 16'd42824, 16'd7069, 16'd49512, 16'd41648, 16'd32995, 16'd42607, 16'd16624, 16'd55445, 16'd8238, 16'd45657, 16'd12474, 16'd5388, 16'd10136, 16'd42670, 16'd44033, 16'd1257});
	test_expansion(128'hcbde4d6eacfd64b86ee4874eb4396164, {16'd58186, 16'd50697, 16'd4156, 16'd7136, 16'd18154, 16'd10188, 16'd26783, 16'd49449, 16'd44201, 16'd14950, 16'd48760, 16'd51219, 16'd27635, 16'd662, 16'd44505, 16'd58391, 16'd7954, 16'd31032, 16'd15362, 16'd5496, 16'd48983, 16'd57832, 16'd23144, 16'd64334, 16'd39308, 16'd21151});
	test_expansion(128'h1606553f7811306d67ac02eb46592f6c, {16'd15944, 16'd61227, 16'd20346, 16'd60597, 16'd12881, 16'd50946, 16'd11196, 16'd2157, 16'd63299, 16'd3691, 16'd49772, 16'd13524, 16'd31049, 16'd15918, 16'd54423, 16'd63497, 16'd11457, 16'd56002, 16'd15110, 16'd60324, 16'd4571, 16'd15700, 16'd61016, 16'd31906, 16'd13027, 16'd60746});
	test_expansion(128'ha3dd056313b2f98bff7fcf7ba1af6165, {16'd44923, 16'd34982, 16'd18384, 16'd8057, 16'd54903, 16'd64064, 16'd42040, 16'd37149, 16'd44136, 16'd40033, 16'd55116, 16'd38542, 16'd27300, 16'd42897, 16'd58196, 16'd47839, 16'd10440, 16'd6290, 16'd51780, 16'd64160, 16'd27533, 16'd57027, 16'd45545, 16'd9845, 16'd44030, 16'd58324});
	test_expansion(128'hbbe13d34e7c662f079f28a738b3a5aae, {16'd58309, 16'd23229, 16'd58652, 16'd42105, 16'd26012, 16'd58236, 16'd5621, 16'd56501, 16'd26886, 16'd65443, 16'd31639, 16'd61796, 16'd13234, 16'd64664, 16'd43419, 16'd52100, 16'd8134, 16'd64892, 16'd64527, 16'd23597, 16'd15307, 16'd6107, 16'd64380, 16'd36874, 16'd23945, 16'd16088});
	test_expansion(128'h8171888ceb2e17f1938fd2fd51341e52, {16'd62601, 16'd62633, 16'd57399, 16'd20643, 16'd64013, 16'd19789, 16'd45643, 16'd27333, 16'd7258, 16'd61248, 16'd58916, 16'd21517, 16'd19381, 16'd21665, 16'd47316, 16'd33632, 16'd50387, 16'd39094, 16'd6331, 16'd58688, 16'd13393, 16'd14874, 16'd63413, 16'd31403, 16'd42616, 16'd29426});
	test_expansion(128'hb317ec990ef19d417ae181dd2275472e, {16'd3899, 16'd16514, 16'd28622, 16'd23526, 16'd11180, 16'd47899, 16'd28988, 16'd19588, 16'd35868, 16'd30030, 16'd42751, 16'd21581, 16'd11531, 16'd5017, 16'd23980, 16'd61683, 16'd14092, 16'd30416, 16'd55880, 16'd47471, 16'd41513, 16'd65535, 16'd61729, 16'd54717, 16'd14355, 16'd64959});
	test_expansion(128'h6438cdc0f43d504ed24108398844addb, {16'd50567, 16'd31051, 16'd55695, 16'd36787, 16'd37688, 16'd14096, 16'd37436, 16'd46358, 16'd27963, 16'd39688, 16'd32160, 16'd28414, 16'd6818, 16'd29929, 16'd15, 16'd33600, 16'd1042, 16'd47520, 16'd48882, 16'd63725, 16'd42247, 16'd52228, 16'd11044, 16'd45423, 16'd17483, 16'd7371});
	test_expansion(128'h32df14931e4ea003b3c027a13417b434, {16'd40933, 16'd12454, 16'd49015, 16'd23657, 16'd9608, 16'd191, 16'd4548, 16'd16569, 16'd50859, 16'd23216, 16'd44673, 16'd45306, 16'd50912, 16'd43362, 16'd28484, 16'd38727, 16'd61643, 16'd12230, 16'd65268, 16'd11242, 16'd43676, 16'd30753, 16'd28724, 16'd63653, 16'd35694, 16'd54629});
	test_expansion(128'ha748a05efe1f6bb2deb64a8419935694, {16'd25843, 16'd22705, 16'd48160, 16'd43656, 16'd65045, 16'd25523, 16'd62572, 16'd35042, 16'd43944, 16'd20704, 16'd44110, 16'd19890, 16'd31766, 16'd43692, 16'd59484, 16'd39528, 16'd43001, 16'd27968, 16'd32870, 16'd63720, 16'd10471, 16'd53430, 16'd44205, 16'd48093, 16'd17599, 16'd28568});
	test_expansion(128'h6835ac3862e5a275e4a916474d094d6a, {16'd28765, 16'd47927, 16'd37337, 16'd34613, 16'd13658, 16'd23834, 16'd62749, 16'd2348, 16'd32317, 16'd39810, 16'd34155, 16'd64550, 16'd31453, 16'd52039, 16'd35422, 16'd5411, 16'd188, 16'd45576, 16'd50640, 16'd63645, 16'd14411, 16'd50727, 16'd15809, 16'd50558, 16'd59527, 16'd12118});
	test_expansion(128'h1329d1d026af252392fe0fac70af158f, {16'd55212, 16'd57259, 16'd45931, 16'd60059, 16'd6761, 16'd36248, 16'd30097, 16'd14425, 16'd45723, 16'd37782, 16'd31692, 16'd23572, 16'd11806, 16'd37278, 16'd40627, 16'd52193, 16'd28429, 16'd47078, 16'd9938, 16'd1927, 16'd61258, 16'd62211, 16'd56205, 16'd56176, 16'd55688, 16'd45770});
	test_expansion(128'h916b9244f1bde29ac76e6e212770c7a5, {16'd45765, 16'd5576, 16'd18622, 16'd5528, 16'd61400, 16'd33654, 16'd56185, 16'd12378, 16'd3586, 16'd60818, 16'd32178, 16'd3602, 16'd39767, 16'd41189, 16'd15206, 16'd60982, 16'd18855, 16'd22287, 16'd6309, 16'd20080, 16'd43574, 16'd45882, 16'd2788, 16'd48796, 16'd52346, 16'd57402});
	test_expansion(128'h56c72363f7423aa30d5b73d7a5019a48, {16'd61510, 16'd58210, 16'd10343, 16'd41002, 16'd15738, 16'd9892, 16'd8793, 16'd61318, 16'd17186, 16'd2973, 16'd19745, 16'd2868, 16'd29192, 16'd57752, 16'd59653, 16'd55195, 16'd26217, 16'd58949, 16'd55578, 16'd13726, 16'd21401, 16'd61601, 16'd61554, 16'd33470, 16'd20192, 16'd58859});
	test_expansion(128'h61e6e9b03ab20e5b62ddaf2717bf7061, {16'd35370, 16'd37710, 16'd43709, 16'd11070, 16'd53474, 16'd29439, 16'd45300, 16'd46284, 16'd13798, 16'd64603, 16'd35967, 16'd58743, 16'd25370, 16'd12677, 16'd51283, 16'd31982, 16'd44678, 16'd57541, 16'd57063, 16'd35826, 16'd24387, 16'd47223, 16'd19231, 16'd12953, 16'd59336, 16'd13047});
	test_expansion(128'h2acae05aeb1efb6c4f41b7c1d96c3823, {16'd60682, 16'd54609, 16'd37281, 16'd34193, 16'd62617, 16'd48647, 16'd25026, 16'd27982, 16'd50037, 16'd61170, 16'd7650, 16'd27788, 16'd23465, 16'd3212, 16'd12231, 16'd16056, 16'd16983, 16'd52498, 16'd11552, 16'd47967, 16'd61386, 16'd55411, 16'd9804, 16'd49317, 16'd13527, 16'd44773});
	test_expansion(128'h11e11b8e74a68ebaf8d6a9453726f9f4, {16'd53192, 16'd65053, 16'd24435, 16'd60366, 16'd30218, 16'd60456, 16'd45851, 16'd3082, 16'd58590, 16'd24626, 16'd33991, 16'd21535, 16'd42740, 16'd65423, 16'd42272, 16'd27549, 16'd2507, 16'd10128, 16'd40158, 16'd38714, 16'd6020, 16'd45583, 16'd21933, 16'd35928, 16'd28522, 16'd12095});
	test_expansion(128'hd898af670cc72dd33a08b51a167b7552, {16'd45993, 16'd14398, 16'd53783, 16'd43096, 16'd17927, 16'd26341, 16'd55347, 16'd50643, 16'd57336, 16'd11865, 16'd37949, 16'd20240, 16'd59132, 16'd29161, 16'd37437, 16'd11393, 16'd14129, 16'd3363, 16'd47014, 16'd19284, 16'd43086, 16'd55861, 16'd33917, 16'd21101, 16'd29351, 16'd19790});
	test_expansion(128'h69b8e24ff07a4cb79c126dc53430188e, {16'd33015, 16'd7582, 16'd44898, 16'd48406, 16'd40080, 16'd35867, 16'd46225, 16'd42789, 16'd26883, 16'd26152, 16'd3566, 16'd60632, 16'd5503, 16'd51418, 16'd40507, 16'd1554, 16'd144, 16'd32221, 16'd7382, 16'd18423, 16'd10904, 16'd33918, 16'd20667, 16'd13664, 16'd32510, 16'd32114});
	test_expansion(128'h5fdbaed29a368bce0f3fbec4f35cf7be, {16'd4417, 16'd24539, 16'd39777, 16'd40559, 16'd52013, 16'd36878, 16'd48411, 16'd59784, 16'd50110, 16'd5297, 16'd48288, 16'd8629, 16'd37999, 16'd52322, 16'd44844, 16'd21656, 16'd63835, 16'd12713, 16'd37706, 16'd63507, 16'd29117, 16'd45523, 16'd24668, 16'd640, 16'd62001, 16'd45410});
	test_expansion(128'h20533e18338f44c2e995ebc4f0a4391b, {16'd15697, 16'd53625, 16'd20466, 16'd22685, 16'd55299, 16'd29741, 16'd46963, 16'd44498, 16'd48878, 16'd24016, 16'd14543, 16'd53158, 16'd40288, 16'd14798, 16'd45513, 16'd1825, 16'd28149, 16'd27666, 16'd20045, 16'd23472, 16'd35286, 16'd15438, 16'd5249, 16'd20633, 16'd16234, 16'd53358});
	test_expansion(128'hc34c9244bb5b16438414a3d958349e13, {16'd49888, 16'd11989, 16'd51628, 16'd16604, 16'd927, 16'd52399, 16'd42341, 16'd56317, 16'd10778, 16'd27998, 16'd30905, 16'd42339, 16'd16507, 16'd37029, 16'd62474, 16'd6991, 16'd61850, 16'd34846, 16'd59367, 16'd25666, 16'd13224, 16'd5791, 16'd58984, 16'd13845, 16'd27709, 16'd55882});
	test_expansion(128'h8d3716e1d46f2873058c3efb9a89c737, {16'd57690, 16'd47125, 16'd36264, 16'd31845, 16'd13891, 16'd40837, 16'd54660, 16'd55726, 16'd3633, 16'd44397, 16'd20533, 16'd6964, 16'd44058, 16'd1706, 16'd37215, 16'd14725, 16'd65289, 16'd42768, 16'd58253, 16'd57681, 16'd4088, 16'd9045, 16'd12684, 16'd63493, 16'd18385, 16'd37886});
	test_expansion(128'hc74b0ee7868c32c8c5ec467e69992af9, {16'd30218, 16'd54470, 16'd37773, 16'd43384, 16'd25808, 16'd27678, 16'd25219, 16'd19208, 16'd33214, 16'd39333, 16'd12474, 16'd5556, 16'd31992, 16'd11756, 16'd5365, 16'd17442, 16'd44898, 16'd63328, 16'd54774, 16'd62359, 16'd24289, 16'd22011, 16'd8784, 16'd62913, 16'd21215, 16'd39307});
	test_expansion(128'hb63524151947d17ba23f966eb34d0af6, {16'd58155, 16'd499, 16'd6974, 16'd57262, 16'd45854, 16'd59538, 16'd62049, 16'd25273, 16'd13503, 16'd60496, 16'd45771, 16'd30821, 16'd28639, 16'd4884, 16'd60355, 16'd37261, 16'd39494, 16'd26135, 16'd47066, 16'd58776, 16'd47132, 16'd63695, 16'd60733, 16'd56460, 16'd4177, 16'd18630});
	test_expansion(128'hf93bc367a9014c8e4a4bc83c4827e824, {16'd819, 16'd24039, 16'd41866, 16'd34108, 16'd29470, 16'd34767, 16'd26273, 16'd64903, 16'd19825, 16'd21188, 16'd46452, 16'd12018, 16'd13595, 16'd40756, 16'd42461, 16'd62564, 16'd54355, 16'd61840, 16'd22100, 16'd9934, 16'd7261, 16'd54914, 16'd48290, 16'd22873, 16'd46819, 16'd40601});
	test_expansion(128'h584af9e46ff9ac6c3865a8830ea16423, {16'd47951, 16'd18855, 16'd32422, 16'd8037, 16'd3482, 16'd38095, 16'd14469, 16'd40718, 16'd27060, 16'd12127, 16'd45713, 16'd44332, 16'd12678, 16'd18965, 16'd59163, 16'd16899, 16'd50483, 16'd29912, 16'd50310, 16'd38881, 16'd26046, 16'd35163, 16'd12795, 16'd27250, 16'd1327, 16'd35138});
	test_expansion(128'hfd89792e159ef197b5d9505f288ddecc, {16'd36106, 16'd58815, 16'd5441, 16'd55344, 16'd1188, 16'd16006, 16'd64129, 16'd23583, 16'd44005, 16'd42752, 16'd33889, 16'd59266, 16'd35005, 16'd30085, 16'd41155, 16'd27664, 16'd33701, 16'd62352, 16'd23923, 16'd35624, 16'd10578, 16'd60272, 16'd32422, 16'd56196, 16'd60187, 16'd52568});
	test_expansion(128'hf884d7b9c26d06f0aed70629ec33c732, {16'd38938, 16'd37711, 16'd60796, 16'd64704, 16'd41766, 16'd40591, 16'd27509, 16'd51047, 16'd57896, 16'd21387, 16'd1772, 16'd38175, 16'd40758, 16'd59592, 16'd21458, 16'd52033, 16'd54899, 16'd28379, 16'd43020, 16'd13765, 16'd26819, 16'd33642, 16'd3837, 16'd10931, 16'd8639, 16'd23117});
	test_expansion(128'h6bd08d66ba95f52dfc807c5d3fbe878c, {16'd46669, 16'd62485, 16'd52041, 16'd33151, 16'd27643, 16'd8219, 16'd50945, 16'd65307, 16'd16111, 16'd53624, 16'd25235, 16'd44973, 16'd46554, 16'd48467, 16'd17197, 16'd22610, 16'd31179, 16'd4346, 16'd22102, 16'd51735, 16'd56519, 16'd13827, 16'd143, 16'd29558, 16'd14576, 16'd45752});
	test_expansion(128'hef56ac71e5987f390719fad15033101a, {16'd22048, 16'd41743, 16'd17875, 16'd13653, 16'd37330, 16'd61680, 16'd47712, 16'd15262, 16'd58892, 16'd32768, 16'd31164, 16'd34331, 16'd17163, 16'd65057, 16'd20231, 16'd47676, 16'd61803, 16'd37858, 16'd57841, 16'd59862, 16'd32968, 16'd5611, 16'd38633, 16'd54600, 16'd33429, 16'd13296});
	test_expansion(128'hbc957b63275cba372fb10c733da18825, {16'd49409, 16'd42342, 16'd17005, 16'd36086, 16'd44431, 16'd47822, 16'd4333, 16'd54614, 16'd57329, 16'd5592, 16'd44221, 16'd41318, 16'd17816, 16'd9104, 16'd480, 16'd10925, 16'd45835, 16'd14926, 16'd15227, 16'd1038, 16'd15814, 16'd51941, 16'd11555, 16'd62500, 16'd39823, 16'd87});
	test_expansion(128'h065f4933d226e73ab9d04e2449b7adfa, {16'd21042, 16'd26742, 16'd10434, 16'd1159, 16'd3609, 16'd20287, 16'd8323, 16'd6995, 16'd29062, 16'd63574, 16'd15801, 16'd10428, 16'd41047, 16'd63026, 16'd46713, 16'd26255, 16'd45091, 16'd31894, 16'd26741, 16'd62259, 16'd12544, 16'd56728, 16'd15397, 16'd11067, 16'd50922, 16'd44800});
	test_expansion(128'h8f27688b4b9640d2c61dd6a86e94fef9, {16'd15135, 16'd45872, 16'd34972, 16'd50913, 16'd60147, 16'd47950, 16'd63631, 16'd26374, 16'd48762, 16'd16303, 16'd437, 16'd38497, 16'd27520, 16'd38430, 16'd40232, 16'd37890, 16'd8816, 16'd58932, 16'd49335, 16'd34847, 16'd65464, 16'd21738, 16'd6610, 16'd46855, 16'd3678, 16'd61699});
	test_expansion(128'hcbaea997a1262f2c51b7901a9029ccd0, {16'd15859, 16'd10947, 16'd43578, 16'd39542, 16'd65317, 16'd28962, 16'd40487, 16'd57699, 16'd58133, 16'd57628, 16'd52195, 16'd35747, 16'd13784, 16'd58444, 16'd63531, 16'd6248, 16'd63663, 16'd23545, 16'd31653, 16'd21881, 16'd49581, 16'd31082, 16'd52961, 16'd19510, 16'd8330, 16'd20875});
	test_expansion(128'h39f22f215fa8bf96ece4528d7e97a720, {16'd47112, 16'd28332, 16'd37649, 16'd46640, 16'd9480, 16'd54654, 16'd13467, 16'd1245, 16'd50073, 16'd32979, 16'd51253, 16'd20598, 16'd34140, 16'd24554, 16'd52654, 16'd37416, 16'd49174, 16'd59432, 16'd14230, 16'd63452, 16'd55162, 16'd14552, 16'd5591, 16'd23119, 16'd35796, 16'd21454});
	test_expansion(128'ha3991be3bfeeaff11f39e8d5b1f95949, {16'd29219, 16'd41800, 16'd61116, 16'd53633, 16'd28079, 16'd2314, 16'd26411, 16'd27778, 16'd26571, 16'd62394, 16'd33152, 16'd4471, 16'd17609, 16'd16184, 16'd28171, 16'd41378, 16'd62777, 16'd21233, 16'd31374, 16'd32285, 16'd9199, 16'd10528, 16'd19643, 16'd37344, 16'd1733, 16'd31119});
	test_expansion(128'he78727aa470e8b34625bd849de52e43d, {16'd40482, 16'd2835, 16'd62125, 16'd60064, 16'd27579, 16'd462, 16'd34837, 16'd29502, 16'd46194, 16'd31421, 16'd9825, 16'd57870, 16'd35435, 16'd33973, 16'd15530, 16'd12768, 16'd63257, 16'd16027, 16'd47504, 16'd36999, 16'd47936, 16'd46186, 16'd65005, 16'd12965, 16'd50650, 16'd9002});
	test_expansion(128'h61b597d797b530e785f16a8a02e5a20a, {16'd40807, 16'd12723, 16'd64266, 16'd33633, 16'd52918, 16'd34675, 16'd58513, 16'd14281, 16'd11751, 16'd47064, 16'd62648, 16'd13961, 16'd2325, 16'd35190, 16'd6504, 16'd54901, 16'd64823, 16'd58874, 16'd20242, 16'd17298, 16'd50742, 16'd63076, 16'd9279, 16'd14562, 16'd37577, 16'd33569});
	test_expansion(128'h892505e76f0052ad63f5e75469d31aaa, {16'd43285, 16'd27897, 16'd47792, 16'd50401, 16'd39380, 16'd2858, 16'd9338, 16'd1403, 16'd53842, 16'd11944, 16'd21574, 16'd55506, 16'd9997, 16'd16674, 16'd18018, 16'd61117, 16'd49021, 16'd1607, 16'd59318, 16'd43978, 16'd35253, 16'd31671, 16'd53170, 16'd28158, 16'd34671, 16'd58976});
	test_expansion(128'hc02606d68fec2acb6c47e0de1ba1bcd0, {16'd53303, 16'd10645, 16'd52879, 16'd11082, 16'd14118, 16'd35747, 16'd32695, 16'd29588, 16'd35326, 16'd11521, 16'd48958, 16'd25055, 16'd61995, 16'd7887, 16'd15222, 16'd37152, 16'd20465, 16'd37751, 16'd5650, 16'd11480, 16'd7523, 16'd20200, 16'd5961, 16'd49380, 16'd29495, 16'd17351});
	test_expansion(128'h45263e7dea786d2ea7b4384d9127a306, {16'd11587, 16'd34644, 16'd17873, 16'd3504, 16'd32613, 16'd62641, 16'd5307, 16'd43091, 16'd7618, 16'd19025, 16'd51335, 16'd37875, 16'd16296, 16'd47884, 16'd34818, 16'd11597, 16'd13865, 16'd4454, 16'd26139, 16'd30437, 16'd5191, 16'd4119, 16'd62125, 16'd36791, 16'd4129, 16'd16660});
	test_expansion(128'h184c99dd8b81884ec1ee497b7909f0fb, {16'd57589, 16'd8007, 16'd30528, 16'd47717, 16'd11175, 16'd63551, 16'd34030, 16'd42567, 16'd61027, 16'd55280, 16'd59447, 16'd21548, 16'd36188, 16'd39729, 16'd2942, 16'd52518, 16'd36412, 16'd48029, 16'd15089, 16'd31953, 16'd18445, 16'd15679, 16'd21663, 16'd3089, 16'd4793, 16'd37985});
	test_expansion(128'h648c6ef5b9f510a9f3b5d10dda28f702, {16'd37454, 16'd48768, 16'd58066, 16'd64573, 16'd14501, 16'd62081, 16'd8357, 16'd45161, 16'd11902, 16'd34809, 16'd52886, 16'd56152, 16'd46633, 16'd359, 16'd59139, 16'd5810, 16'd25142, 16'd21474, 16'd41851, 16'd57871, 16'd20299, 16'd24795, 16'd17442, 16'd44982, 16'd39466, 16'd44054});
	test_expansion(128'h42d6f046e9deb7f292f5e0c0374197d0, {16'd52384, 16'd37955, 16'd21144, 16'd32022, 16'd23313, 16'd60544, 16'd47782, 16'd4821, 16'd24466, 16'd19238, 16'd54265, 16'd26766, 16'd12118, 16'd8330, 16'd21096, 16'd36513, 16'd62380, 16'd21009, 16'd44415, 16'd9531, 16'd5948, 16'd22993, 16'd15286, 16'd54757, 16'd4683, 16'd60655});
	test_expansion(128'h73729b8e5756e8bb71b477c82bebbd19, {16'd5602, 16'd28207, 16'd55441, 16'd31363, 16'd2894, 16'd50232, 16'd52498, 16'd41515, 16'd44224, 16'd43080, 16'd3024, 16'd14060, 16'd64472, 16'd19584, 16'd42973, 16'd26837, 16'd38152, 16'd56170, 16'd16780, 16'd27222, 16'd23611, 16'd43505, 16'd11495, 16'd34574, 16'd387, 16'd64818});
	test_expansion(128'hca889e7410a0a41482550e1153a4b3aa, {16'd54792, 16'd49596, 16'd13808, 16'd14871, 16'd30658, 16'd47442, 16'd64908, 16'd42048, 16'd39688, 16'd49614, 16'd60484, 16'd44974, 16'd11623, 16'd17537, 16'd11366, 16'd39677, 16'd36524, 16'd63651, 16'd14351, 16'd28307, 16'd44600, 16'd5067, 16'd50185, 16'd48017, 16'd23334, 16'd29331});
	test_expansion(128'h4b6a5c11962b36fbff24674bf92eec98, {16'd36295, 16'd41982, 16'd4438, 16'd54446, 16'd27409, 16'd57178, 16'd48209, 16'd11693, 16'd41274, 16'd61088, 16'd59967, 16'd22281, 16'd44418, 16'd59381, 16'd31043, 16'd38106, 16'd47333, 16'd22074, 16'd41452, 16'd3928, 16'd28502, 16'd32638, 16'd41581, 16'd38644, 16'd25680, 16'd45373});
	test_expansion(128'h78a80f4fbd989708bc61c0811413330a, {16'd19923, 16'd40643, 16'd49523, 16'd7715, 16'd19510, 16'd41755, 16'd6888, 16'd32509, 16'd64756, 16'd15884, 16'd48444, 16'd57336, 16'd60419, 16'd43451, 16'd61129, 16'd13455, 16'd1143, 16'd53801, 16'd23287, 16'd61149, 16'd13750, 16'd534, 16'd51357, 16'd35568, 16'd14182, 16'd23197});
	test_expansion(128'h773ddb607d798658ab33936adb5a601e, {16'd29706, 16'd19581, 16'd64014, 16'd35993, 16'd28025, 16'd35920, 16'd462, 16'd57394, 16'd10156, 16'd43059, 16'd29914, 16'd63505, 16'd30293, 16'd22832, 16'd53893, 16'd13716, 16'd7253, 16'd6306, 16'd37534, 16'd28523, 16'd29350, 16'd14477, 16'd13198, 16'd48629, 16'd51197, 16'd64551});
	test_expansion(128'h91758506892c59d4ad25cc7d2ca07d23, {16'd53642, 16'd57129, 16'd52590, 16'd19908, 16'd31910, 16'd53370, 16'd47550, 16'd56909, 16'd58064, 16'd46608, 16'd63739, 16'd26653, 16'd37025, 16'd56734, 16'd50660, 16'd56254, 16'd24184, 16'd4776, 16'd5648, 16'd59736, 16'd18928, 16'd17202, 16'd16495, 16'd30952, 16'd59729, 16'd4055});
	test_expansion(128'hcd962b7755f15ef8eee1bb5b3735b403, {16'd15541, 16'd14098, 16'd7549, 16'd29584, 16'd35863, 16'd10823, 16'd4129, 16'd58757, 16'd59481, 16'd24313, 16'd32176, 16'd52684, 16'd23957, 16'd63360, 16'd23007, 16'd16548, 16'd57840, 16'd56138, 16'd3190, 16'd32323, 16'd55420, 16'd59577, 16'd7522, 16'd42964, 16'd25357, 16'd38535});
	test_expansion(128'h405fcd7e8c26df23efa4a007735f4c84, {16'd63346, 16'd23824, 16'd56550, 16'd19775, 16'd5538, 16'd54669, 16'd1127, 16'd25530, 16'd45257, 16'd44778, 16'd24099, 16'd19840, 16'd52435, 16'd28534, 16'd54744, 16'd49035, 16'd25648, 16'd6493, 16'd8428, 16'd21527, 16'd11571, 16'd55280, 16'd60352, 16'd15693, 16'd29192, 16'd14265});
	test_expansion(128'h23442c9b590797486738ca65c8a7d5ee, {16'd8042, 16'd18702, 16'd33886, 16'd44873, 16'd23160, 16'd14447, 16'd41016, 16'd5796, 16'd16571, 16'd19055, 16'd53988, 16'd34647, 16'd48360, 16'd12988, 16'd17274, 16'd18256, 16'd33372, 16'd21260, 16'd34657, 16'd21817, 16'd7804, 16'd49369, 16'd19522, 16'd33215, 16'd31905, 16'd6139});
	test_expansion(128'hb7e7b8df4c10641c44a84d19217c2c1e, {16'd37609, 16'd39449, 16'd23984, 16'd32200, 16'd38330, 16'd36080, 16'd10336, 16'd38055, 16'd40312, 16'd52203, 16'd36990, 16'd1620, 16'd60608, 16'd60866, 16'd11538, 16'd42503, 16'd30165, 16'd29528, 16'd18279, 16'd45960, 16'd30363, 16'd57052, 16'd33819, 16'd2510, 16'd55527, 16'd29283});
	test_expansion(128'h65afaaf3801b9706fab77a68f24d8b31, {16'd26547, 16'd9818, 16'd29409, 16'd7803, 16'd14971, 16'd22604, 16'd24804, 16'd5593, 16'd35531, 16'd8138, 16'd29569, 16'd33228, 16'd45926, 16'd58492, 16'd22073, 16'd54414, 16'd3758, 16'd2260, 16'd3619, 16'd37319, 16'd21970, 16'd28265, 16'd34344, 16'd17040, 16'd24822, 16'd61264});
	test_expansion(128'h2ade49b0f214d58d8e1c41ddc6a997b9, {16'd39761, 16'd53291, 16'd18405, 16'd31067, 16'd1395, 16'd31561, 16'd1501, 16'd46899, 16'd45583, 16'd33953, 16'd21189, 16'd49392, 16'd31357, 16'd31636, 16'd33879, 16'd1311, 16'd32548, 16'd3548, 16'd56989, 16'd39082, 16'd41996, 16'd41758, 16'd20215, 16'd20015, 16'd25660, 16'd12106});
	test_expansion(128'h5124cfb3df21729ab03b8badda22e63d, {16'd48126, 16'd3672, 16'd32537, 16'd28961, 16'd47074, 16'd12311, 16'd58211, 16'd64216, 16'd34140, 16'd7165, 16'd19200, 16'd41968, 16'd55521, 16'd21477, 16'd42121, 16'd15967, 16'd38459, 16'd22838, 16'd50659, 16'd45398, 16'd32278, 16'd5383, 16'd6145, 16'd10917, 16'd4127, 16'd58181});
	test_expansion(128'h3a8d40ca0d1efecfd05632a016a6eb9a, {16'd33306, 16'd14691, 16'd49229, 16'd40802, 16'd20890, 16'd31788, 16'd32184, 16'd24174, 16'd23502, 16'd45548, 16'd56725, 16'd33762, 16'd48270, 16'd41605, 16'd47501, 16'd31075, 16'd37512, 16'd22675, 16'd38650, 16'd21394, 16'd35908, 16'd10629, 16'd28669, 16'd34472, 16'd29227, 16'd33395});
	test_expansion(128'h9638200e7493daa31e7d421e411cb0eb, {16'd26934, 16'd58746, 16'd60746, 16'd9448, 16'd30368, 16'd8776, 16'd34301, 16'd60852, 16'd34806, 16'd13003, 16'd8695, 16'd29010, 16'd43896, 16'd48055, 16'd20427, 16'd36607, 16'd6525, 16'd13191, 16'd32644, 16'd35074, 16'd6080, 16'd18159, 16'd44673, 16'd13285, 16'd31402, 16'd780});
	test_expansion(128'hbf6e21b3a522cec7467d816bcf9eb7b1, {16'd28546, 16'd7119, 16'd30055, 16'd43219, 16'd51698, 16'd33242, 16'd10754, 16'd52088, 16'd35594, 16'd7792, 16'd23034, 16'd6231, 16'd24265, 16'd6222, 16'd38, 16'd55479, 16'd45913, 16'd51042, 16'd255, 16'd38800, 16'd60827, 16'd36051, 16'd9428, 16'd39866, 16'd24083, 16'd32265});
	test_expansion(128'h418b27417aa8bc514ef9f2c8a606f5dc, {16'd31842, 16'd37102, 16'd64994, 16'd29906, 16'd6044, 16'd4885, 16'd39920, 16'd60007, 16'd38963, 16'd21567, 16'd27684, 16'd1849, 16'd65376, 16'd11961, 16'd34545, 16'd5809, 16'd19755, 16'd18670, 16'd27867, 16'd64897, 16'd32165, 16'd12154, 16'd32194, 16'd22989, 16'd5696, 16'd44602});
	test_expansion(128'ha1440cd711a4ea8bdbd8f9299ed2b60e, {16'd40281, 16'd13843, 16'd35231, 16'd6184, 16'd19928, 16'd5856, 16'd750, 16'd25202, 16'd33149, 16'd10558, 16'd25327, 16'd2068, 16'd20305, 16'd48857, 16'd17043, 16'd32604, 16'd57611, 16'd7329, 16'd64239, 16'd20019, 16'd21344, 16'd45781, 16'd12060, 16'd19444, 16'd51968, 16'd1171});
	test_expansion(128'h6959acb2470ac551483eb1d529ff96ac, {16'd23198, 16'd57597, 16'd50463, 16'd12251, 16'd19384, 16'd14156, 16'd10840, 16'd31890, 16'd40959, 16'd19341, 16'd14437, 16'd41483, 16'd30117, 16'd34495, 16'd20482, 16'd19177, 16'd12688, 16'd62420, 16'd42767, 16'd53104, 16'd2475, 16'd8706, 16'd30458, 16'd24407, 16'd56278, 16'd55417});
	test_expansion(128'h864aa8806ff17249102ef050540bb516, {16'd15155, 16'd36783, 16'd32322, 16'd51866, 16'd14454, 16'd46392, 16'd22530, 16'd50189, 16'd34986, 16'd23730, 16'd23274, 16'd38329, 16'd58347, 16'd11013, 16'd4996, 16'd60930, 16'd63645, 16'd17568, 16'd38996, 16'd48256, 16'd61620, 16'd1340, 16'd40766, 16'd7521, 16'd4357, 16'd31959});
	test_expansion(128'hf18f6cbc07499fe2fe42346b28d884cd, {16'd58774, 16'd52888, 16'd38561, 16'd42253, 16'd40696, 16'd1311, 16'd27136, 16'd4687, 16'd19390, 16'd17515, 16'd21851, 16'd61575, 16'd29146, 16'd2382, 16'd44264, 16'd10862, 16'd60876, 16'd57178, 16'd54363, 16'd51957, 16'd46118, 16'd37437, 16'd15641, 16'd33502, 16'd9246, 16'd58571});
	test_expansion(128'hf763042c19a242dcaabcc2e7d73bc0d1, {16'd4521, 16'd8839, 16'd61413, 16'd46847, 16'd49905, 16'd43318, 16'd60684, 16'd19283, 16'd57229, 16'd56745, 16'd15988, 16'd22049, 16'd30422, 16'd60674, 16'd44246, 16'd23173, 16'd34424, 16'd7690, 16'd36882, 16'd45192, 16'd62663, 16'd2412, 16'd59421, 16'd62501, 16'd2582, 16'd30358});
	test_expansion(128'h1064e94ccefa3549323680c3a7fc4f41, {16'd24496, 16'd31030, 16'd9843, 16'd40304, 16'd44182, 16'd28155, 16'd21738, 16'd5073, 16'd19494, 16'd42646, 16'd56080, 16'd27895, 16'd29122, 16'd40387, 16'd15272, 16'd7349, 16'd59074, 16'd6149, 16'd40387, 16'd53599, 16'd49005, 16'd15276, 16'd17328, 16'd54575, 16'd37208, 16'd42962});
	test_expansion(128'h99f82ce0ed36c12ee0d5404a22d05ecb, {16'd7600, 16'd16285, 16'd6573, 16'd31715, 16'd58181, 16'd1217, 16'd21101, 16'd5861, 16'd41177, 16'd55704, 16'd12023, 16'd10234, 16'd49655, 16'd49959, 16'd60839, 16'd1050, 16'd37467, 16'd28330, 16'd60774, 16'd13976, 16'd28357, 16'd38387, 16'd28137, 16'd38097, 16'd37337, 16'd56631});
	test_expansion(128'h2d7cffa885735155a466714f6707f8f6, {16'd43405, 16'd36535, 16'd6401, 16'd36442, 16'd54174, 16'd50275, 16'd23486, 16'd19818, 16'd29164, 16'd37657, 16'd55725, 16'd16262, 16'd27870, 16'd47383, 16'd59646, 16'd16250, 16'd57779, 16'd35949, 16'd15762, 16'd25344, 16'd7412, 16'd47633, 16'd14172, 16'd4788, 16'd14445, 16'd29039});
	test_expansion(128'h5476664a84cc592ee77c5ca1bd627894, {16'd46438, 16'd21742, 16'd41967, 16'd43022, 16'd61814, 16'd5792, 16'd60429, 16'd37025, 16'd24638, 16'd62842, 16'd47591, 16'd9879, 16'd58565, 16'd58820, 16'd52350, 16'd22815, 16'd22197, 16'd46011, 16'd905, 16'd10820, 16'd49083, 16'd46344, 16'd23355, 16'd63514, 16'd61821, 16'd10429});
	test_expansion(128'h214c2d697fe8775666edb89cb944a3a7, {16'd48970, 16'd48097, 16'd28882, 16'd34176, 16'd56967, 16'd5443, 16'd7428, 16'd18101, 16'd63303, 16'd23967, 16'd60345, 16'd48277, 16'd314, 16'd33389, 16'd33623, 16'd53413, 16'd47754, 16'd21428, 16'd18023, 16'd24225, 16'd57077, 16'd39546, 16'd16319, 16'd55069, 16'd16063, 16'd36876});
	test_expansion(128'h9f80122f8b91cb55b7abff975ce88109, {16'd24224, 16'd13052, 16'd20839, 16'd9302, 16'd57706, 16'd49404, 16'd51934, 16'd30043, 16'd35278, 16'd35645, 16'd40100, 16'd45828, 16'd36705, 16'd15262, 16'd35872, 16'd64983, 16'd25805, 16'd25204, 16'd28847, 16'd30788, 16'd63823, 16'd31291, 16'd54297, 16'd30086, 16'd45870, 16'd33412});
	test_expansion(128'h4165bb77f65f051833cfba5170bd4013, {16'd51095, 16'd59951, 16'd9337, 16'd15626, 16'd25999, 16'd24070, 16'd41627, 16'd218, 16'd38713, 16'd4379, 16'd58193, 16'd49900, 16'd363, 16'd54663, 16'd33790, 16'd62198, 16'd42524, 16'd4160, 16'd33848, 16'd44763, 16'd2626, 16'd42627, 16'd7323, 16'd61401, 16'd12822, 16'd10313});
	test_expansion(128'h47e08b364d9abc09f04fd7f1b37f6f57, {16'd25399, 16'd22063, 16'd36521, 16'd37092, 16'd29771, 16'd12217, 16'd54404, 16'd6369, 16'd27819, 16'd38272, 16'd46274, 16'd15437, 16'd30494, 16'd15552, 16'd35882, 16'd63241, 16'd40613, 16'd37197, 16'd36684, 16'd47076, 16'd51315, 16'd31504, 16'd37404, 16'd22168, 16'd56463, 16'd17663});
	test_expansion(128'h1a882029730c2c8c0f464dd93a2ac9e0, {16'd56353, 16'd47422, 16'd48583, 16'd1233, 16'd9268, 16'd25878, 16'd44088, 16'd61493, 16'd56745, 16'd50224, 16'd28547, 16'd6264, 16'd35402, 16'd31152, 16'd8763, 16'd260, 16'd21779, 16'd2667, 16'd53898, 16'd26421, 16'd9324, 16'd47891, 16'd21350, 16'd21821, 16'd33528, 16'd2042});
	test_expansion(128'hdba8449369ae5be9bfa0db0513341c86, {16'd14935, 16'd36735, 16'd4189, 16'd52849, 16'd53639, 16'd30830, 16'd7, 16'd52221, 16'd24990, 16'd2958, 16'd64705, 16'd4648, 16'd19755, 16'd39194, 16'd49370, 16'd61739, 16'd24148, 16'd26824, 16'd20103, 16'd15366, 16'd60017, 16'd57519, 16'd46805, 16'd26950, 16'd27994, 16'd2343});
	test_expansion(128'hf086f5aa4c6214ae0a7628cf2478f258, {16'd7529, 16'd12975, 16'd3525, 16'd32341, 16'd47983, 16'd6043, 16'd14877, 16'd61803, 16'd29662, 16'd33924, 16'd6787, 16'd10472, 16'd64770, 16'd42996, 16'd2336, 16'd2737, 16'd26021, 16'd64244, 16'd13582, 16'd39573, 16'd41800, 16'd3378, 16'd17244, 16'd39347, 16'd49803, 16'd63680});
	test_expansion(128'h482b7aeef0d05621f5b20ae9c6276a66, {16'd29973, 16'd16810, 16'd25872, 16'd8403, 16'd57165, 16'd39891, 16'd27833, 16'd23518, 16'd65472, 16'd21382, 16'd51950, 16'd44396, 16'd11708, 16'd7613, 16'd38715, 16'd56625, 16'd47314, 16'd42712, 16'd29535, 16'd30368, 16'd13175, 16'd24070, 16'd45643, 16'd37766, 16'd25990, 16'd5438});
	test_expansion(128'hea339dbde12030014120d089b3cd1674, {16'd56111, 16'd59854, 16'd16231, 16'd14747, 16'd6421, 16'd26573, 16'd16396, 16'd49354, 16'd4378, 16'd53422, 16'd21463, 16'd53581, 16'd6758, 16'd52912, 16'd52688, 16'd5270, 16'd14661, 16'd61255, 16'd14839, 16'd29934, 16'd37518, 16'd46818, 16'd44033, 16'd29865, 16'd2361, 16'd21268});
	test_expansion(128'h8d380eb62d2dba8eae90d3f875af229b, {16'd10549, 16'd28276, 16'd3980, 16'd58257, 16'd63578, 16'd57986, 16'd56069, 16'd25482, 16'd14978, 16'd50468, 16'd17302, 16'd18887, 16'd15031, 16'd34415, 16'd1713, 16'd37392, 16'd41458, 16'd58933, 16'd36466, 16'd11695, 16'd17550, 16'd38634, 16'd56226, 16'd56339, 16'd37520, 16'd58557});
	test_expansion(128'h2f366702e0bc7a25d9ccaa756541e522, {16'd46212, 16'd54972, 16'd16338, 16'd59857, 16'd63842, 16'd56415, 16'd28425, 16'd53406, 16'd15691, 16'd15654, 16'd11169, 16'd34486, 16'd18955, 16'd14763, 16'd38927, 16'd60211, 16'd43262, 16'd58531, 16'd19856, 16'd39968, 16'd27858, 16'd23131, 16'd15742, 16'd32258, 16'd57491, 16'd14529});
	test_expansion(128'haa863cf6caa0277661f80ac2d4885f57, {16'd2870, 16'd1822, 16'd49458, 16'd1778, 16'd10918, 16'd10612, 16'd52774, 16'd58081, 16'd40169, 16'd55642, 16'd57698, 16'd11092, 16'd5532, 16'd19273, 16'd44438, 16'd47091, 16'd15573, 16'd51276, 16'd18123, 16'd30375, 16'd20540, 16'd24266, 16'd59928, 16'd62619, 16'd34268, 16'd41169});
	test_expansion(128'hb80df25445124b5fb675683062ff3bdc, {16'd33820, 16'd61798, 16'd37636, 16'd55455, 16'd3850, 16'd60567, 16'd5369, 16'd16456, 16'd44432, 16'd44735, 16'd57349, 16'd7997, 16'd10068, 16'd51818, 16'd64274, 16'd36671, 16'd51639, 16'd45835, 16'd31289, 16'd55253, 16'd63286, 16'd61346, 16'd10896, 16'd508, 16'd55841, 16'd64094});
	test_expansion(128'h56768be4ab7ea004ab74095696bbb98a, {16'd61177, 16'd22534, 16'd884, 16'd5620, 16'd8343, 16'd23403, 16'd47359, 16'd50961, 16'd46246, 16'd34426, 16'd31572, 16'd36515, 16'd7714, 16'd11501, 16'd46073, 16'd27078, 16'd29056, 16'd42637, 16'd36368, 16'd50863, 16'd11775, 16'd62924, 16'd26824, 16'd54863, 16'd26141, 16'd47857});
	test_expansion(128'hdf3de7648c97a0ffa38f39fb9f1dc062, {16'd26820, 16'd59037, 16'd47870, 16'd16976, 16'd7482, 16'd13286, 16'd59446, 16'd37188, 16'd56193, 16'd29746, 16'd39720, 16'd3133, 16'd41841, 16'd12604, 16'd22845, 16'd57817, 16'd57474, 16'd40016, 16'd44035, 16'd4877, 16'd39367, 16'd52458, 16'd2864, 16'd1174, 16'd23360, 16'd27975});
	test_expansion(128'h23505082c0820985a9cd0213fbc70c93, {16'd32046, 16'd59102, 16'd53829, 16'd60338, 16'd19451, 16'd13860, 16'd9897, 16'd33739, 16'd10271, 16'd29861, 16'd39424, 16'd459, 16'd26829, 16'd10428, 16'd32467, 16'd32751, 16'd51849, 16'd60947, 16'd25335, 16'd28251, 16'd15724, 16'd14481, 16'd55294, 16'd60889, 16'd34784, 16'd62513});
	test_expansion(128'h0d00530d39f8e18e63d48a4751fd7b80, {16'd63724, 16'd43175, 16'd25483, 16'd64589, 16'd19168, 16'd13253, 16'd4967, 16'd51711, 16'd50946, 16'd59605, 16'd23383, 16'd39141, 16'd12385, 16'd33599, 16'd30388, 16'd27392, 16'd17496, 16'd22514, 16'd16770, 16'd636, 16'd45677, 16'd10853, 16'd12700, 16'd59726, 16'd41301, 16'd31337});
	test_expansion(128'h2f0d933812fbde681b8676be4698eb91, {16'd1512, 16'd42847, 16'd46534, 16'd8712, 16'd12853, 16'd14284, 16'd25739, 16'd58560, 16'd32134, 16'd12562, 16'd41163, 16'd4679, 16'd50694, 16'd57739, 16'd16692, 16'd45583, 16'd57363, 16'd11802, 16'd41611, 16'd32427, 16'd56997, 16'd6850, 16'd38992, 16'd26922, 16'd63300, 16'd40551});
	test_expansion(128'hca224c3279c4f24785ac0ad980217fa3, {16'd2743, 16'd53734, 16'd38072, 16'd59849, 16'd62819, 16'd27028, 16'd43702, 16'd20589, 16'd4655, 16'd23080, 16'd59272, 16'd24440, 16'd21556, 16'd11439, 16'd58395, 16'd58405, 16'd56600, 16'd30339, 16'd14654, 16'd32202, 16'd32933, 16'd31101, 16'd42354, 16'd31144, 16'd64046, 16'd46900});
	test_expansion(128'heb49ef1464a0c079005d0a5d6f446bd4, {16'd55100, 16'd21905, 16'd55516, 16'd4923, 16'd19093, 16'd57318, 16'd36171, 16'd21477, 16'd46917, 16'd427, 16'd53051, 16'd54684, 16'd40422, 16'd1471, 16'd61502, 16'd26172, 16'd58211, 16'd40676, 16'd8413, 16'd8760, 16'd65061, 16'd21041, 16'd55377, 16'd59148, 16'd42056, 16'd45433});
	test_expansion(128'hc4ae99777970ddca969058ddea1b8b32, {16'd12474, 16'd16347, 16'd62823, 16'd62670, 16'd52207, 16'd30497, 16'd31809, 16'd4765, 16'd14615, 16'd28583, 16'd33700, 16'd15815, 16'd62635, 16'd13482, 16'd40004, 16'd47158, 16'd3114, 16'd6278, 16'd14936, 16'd19319, 16'd38064, 16'd59154, 16'd585, 16'd29452, 16'd3057, 16'd56312});
	test_expansion(128'h711450cd8e5a0ee8ad772bb503c38efd, {16'd65127, 16'd19995, 16'd51541, 16'd52979, 16'd16066, 16'd36953, 16'd19684, 16'd43190, 16'd41950, 16'd58985, 16'd40916, 16'd33625, 16'd21122, 16'd25414, 16'd60187, 16'd26273, 16'd32561, 16'd48212, 16'd26336, 16'd33664, 16'd42938, 16'd6818, 16'd54893, 16'd50900, 16'd57575, 16'd17513});
	test_expansion(128'h4860aef7e23bccd630055c7caa30c226, {16'd25815, 16'd42980, 16'd56792, 16'd7542, 16'd57676, 16'd55819, 16'd54212, 16'd24375, 16'd57764, 16'd55300, 16'd31937, 16'd41653, 16'd4, 16'd19634, 16'd38078, 16'd24189, 16'd63515, 16'd36461, 16'd22623, 16'd17866, 16'd43351, 16'd61349, 16'd42889, 16'd24259, 16'd24543, 16'd22597});
	test_expansion(128'hf4c0f0828aed22fb9a0435717e5e7ca4, {16'd2314, 16'd57438, 16'd47279, 16'd30351, 16'd55220, 16'd40418, 16'd56203, 16'd40575, 16'd48665, 16'd3833, 16'd53763, 16'd55130, 16'd38627, 16'd7459, 16'd43015, 16'd9733, 16'd59949, 16'd18939, 16'd60934, 16'd40316, 16'd36365, 16'd25254, 16'd8335, 16'd38895, 16'd24923, 16'd43163});
	test_expansion(128'hf6772a2d5ac5710b9a6c9bcd79679f30, {16'd49986, 16'd56734, 16'd53981, 16'd8121, 16'd35092, 16'd49478, 16'd65050, 16'd35431, 16'd56110, 16'd44065, 16'd24212, 16'd4367, 16'd4358, 16'd2039, 16'd39912, 16'd1689, 16'd48505, 16'd16082, 16'd234, 16'd43338, 16'd50010, 16'd13752, 16'd62888, 16'd21796, 16'd56137, 16'd56461});
	test_expansion(128'hcbbbf07d6ea0fe412ec77348b153a293, {16'd45899, 16'd46777, 16'd40206, 16'd4828, 16'd42736, 16'd46755, 16'd15261, 16'd47525, 16'd23003, 16'd17943, 16'd47853, 16'd1913, 16'd58942, 16'd44876, 16'd19832, 16'd14495, 16'd21728, 16'd12207, 16'd40422, 16'd28163, 16'd52024, 16'd24128, 16'd7177, 16'd26968, 16'd56293, 16'd17317});
	test_expansion(128'hde49bfec81ed359388dfb89fe0095d2b, {16'd57970, 16'd23258, 16'd39271, 16'd54790, 16'd63447, 16'd16598, 16'd42970, 16'd27128, 16'd35001, 16'd45676, 16'd42729, 16'd55946, 16'd1635, 16'd195, 16'd40536, 16'd31473, 16'd2934, 16'd2056, 16'd37057, 16'd46618, 16'd21290, 16'd17000, 16'd43915, 16'd9388, 16'd44166, 16'd63643});
	test_expansion(128'h7d8d2049232f20caf1f0a6ad6838945c, {16'd43405, 16'd63222, 16'd51343, 16'd65052, 16'd14790, 16'd51911, 16'd26171, 16'd57350, 16'd49778, 16'd32062, 16'd43387, 16'd29922, 16'd24211, 16'd16736, 16'd16747, 16'd38087, 16'd49831, 16'd4117, 16'd52662, 16'd16007, 16'd171, 16'd10202, 16'd52432, 16'd57567, 16'd60600, 16'd42881});
	test_expansion(128'h7fc02dcf793614e1f2420111f8322124, {16'd33741, 16'd25273, 16'd16179, 16'd25527, 16'd40241, 16'd15962, 16'd14489, 16'd3811, 16'd36135, 16'd3355, 16'd27552, 16'd41212, 16'd2184, 16'd49735, 16'd31799, 16'd10936, 16'd44446, 16'd62349, 16'd63479, 16'd42553, 16'd41320, 16'd53239, 16'd2164, 16'd24590, 16'd17941, 16'd56497});
	test_expansion(128'hef5a7b34a476cb910b0732439528e648, {16'd47049, 16'd60342, 16'd58671, 16'd44217, 16'd3606, 16'd58686, 16'd35577, 16'd3091, 16'd55667, 16'd59599, 16'd16835, 16'd5944, 16'd31025, 16'd14248, 16'd64424, 16'd42434, 16'd6580, 16'd58913, 16'd61541, 16'd15984, 16'd29645, 16'd30244, 16'd5353, 16'd1485, 16'd6692, 16'd52641});
	test_expansion(128'h1eba8cc30937d180c6c9d335d634b0d4, {16'd56027, 16'd38806, 16'd16238, 16'd34204, 16'd30059, 16'd59726, 16'd25093, 16'd61487, 16'd50059, 16'd11005, 16'd48141, 16'd34967, 16'd19867, 16'd44932, 16'd4701, 16'd15103, 16'd40179, 16'd2058, 16'd8464, 16'd4207, 16'd37934, 16'd56370, 16'd8604, 16'd20803, 16'd63772, 16'd33132});
	test_expansion(128'h529dfa4b186090c7a880d8e2fabbf4fd, {16'd58223, 16'd25034, 16'd35735, 16'd9651, 16'd23741, 16'd8197, 16'd10677, 16'd53249, 16'd43645, 16'd17590, 16'd53187, 16'd15014, 16'd1021, 16'd64084, 16'd23213, 16'd7570, 16'd9095, 16'd38050, 16'd8014, 16'd48816, 16'd52312, 16'd61547, 16'd24594, 16'd9031, 16'd57186, 16'd26683});
	test_expansion(128'ha34d30757a2287cffb61386f01ac3309, {16'd13485, 16'd2493, 16'd19693, 16'd10342, 16'd23669, 16'd11, 16'd48794, 16'd60538, 16'd14425, 16'd21550, 16'd10764, 16'd6889, 16'd41987, 16'd48643, 16'd2463, 16'd11254, 16'd11127, 16'd49030, 16'd18682, 16'd53929, 16'd56825, 16'd25994, 16'd44972, 16'd36087, 16'd55499, 16'd28217});
	test_expansion(128'h06680968d66a93755234cc62e7bd66ce, {16'd28500, 16'd33713, 16'd60256, 16'd3934, 16'd18361, 16'd31106, 16'd5778, 16'd14459, 16'd37659, 16'd61722, 16'd33093, 16'd46762, 16'd24476, 16'd17410, 16'd25741, 16'd29567, 16'd64063, 16'd35477, 16'd28724, 16'd21173, 16'd4944, 16'd62000, 16'd25586, 16'd62992, 16'd35382, 16'd8085});
	test_expansion(128'hc09b0994e066df8bde6ecb6c923a9677, {16'd59589, 16'd31625, 16'd24970, 16'd5230, 16'd22624, 16'd61255, 16'd35497, 16'd11356, 16'd46873, 16'd48681, 16'd15694, 16'd53140, 16'd32970, 16'd434, 16'd23559, 16'd64031, 16'd12079, 16'd32683, 16'd46018, 16'd56489, 16'd52028, 16'd12050, 16'd50132, 16'd19432, 16'd30776, 16'd57247});
	test_expansion(128'hc03ae17ed0bd1be14db0f25e753d3d18, {16'd14171, 16'd2071, 16'd29488, 16'd4408, 16'd44110, 16'd39598, 16'd4552, 16'd54484, 16'd59743, 16'd27978, 16'd44453, 16'd40022, 16'd6861, 16'd3781, 16'd15953, 16'd42966, 16'd30841, 16'd23944, 16'd31723, 16'd19394, 16'd59480, 16'd33077, 16'd57134, 16'd33780, 16'd6456, 16'd43235});
	test_expansion(128'h4cf30aadb2f2e81cadec9c879efe5447, {16'd31717, 16'd12421, 16'd5780, 16'd47867, 16'd53630, 16'd24771, 16'd41959, 16'd64898, 16'd63295, 16'd1127, 16'd53360, 16'd46289, 16'd45480, 16'd26491, 16'd63860, 16'd44692, 16'd16676, 16'd42997, 16'd57309, 16'd61415, 16'd20059, 16'd36281, 16'd57640, 16'd1662, 16'd43811, 16'd68});
	test_expansion(128'h346cfea4d15c7bdce2f3a35c30e0cfeb, {16'd59740, 16'd50306, 16'd30707, 16'd2316, 16'd64475, 16'd52722, 16'd23217, 16'd13635, 16'd15687, 16'd57661, 16'd6226, 16'd47547, 16'd48659, 16'd16653, 16'd8762, 16'd22952, 16'd57306, 16'd54015, 16'd45505, 16'd17517, 16'd38771, 16'd23430, 16'd32479, 16'd16484, 16'd64913, 16'd50433});
	test_expansion(128'hd88732621c576c50674a4ad650a38f6a, {16'd6172, 16'd48598, 16'd22324, 16'd56551, 16'd65249, 16'd21097, 16'd62027, 16'd65170, 16'd22651, 16'd48618, 16'd10490, 16'd53366, 16'd12920, 16'd36061, 16'd2014, 16'd28511, 16'd59919, 16'd34457, 16'd44706, 16'd43655, 16'd38321, 16'd22161, 16'd54295, 16'd56338, 16'd41711, 16'd29976});
	test_expansion(128'h3d4fc191a8764e1dfaeb7118f07e740e, {16'd46522, 16'd48265, 16'd19350, 16'd16595, 16'd41197, 16'd25541, 16'd2032, 16'd7528, 16'd27613, 16'd47958, 16'd59594, 16'd61891, 16'd43090, 16'd46743, 16'd21537, 16'd62676, 16'd45891, 16'd37499, 16'd16082, 16'd49492, 16'd1719, 16'd64999, 16'd47779, 16'd13528, 16'd48995, 16'd38279});
	test_expansion(128'h0f5b4490f7157f8c1f965ff6d8d70827, {16'd26679, 16'd34965, 16'd45865, 16'd50023, 16'd11788, 16'd42325, 16'd22523, 16'd20125, 16'd61963, 16'd30471, 16'd35910, 16'd26060, 16'd7873, 16'd24779, 16'd15757, 16'd61855, 16'd48767, 16'd59341, 16'd55323, 16'd61337, 16'd20249, 16'd42895, 16'd8761, 16'd5317, 16'd43952, 16'd28112});
	test_expansion(128'h892a1d28efa2accd489472e6faf94468, {16'd8954, 16'd58042, 16'd38607, 16'd34179, 16'd4272, 16'd14767, 16'd36217, 16'd61091, 16'd17909, 16'd1698, 16'd49583, 16'd29524, 16'd25626, 16'd4317, 16'd40051, 16'd52170, 16'd46130, 16'd56548, 16'd22036, 16'd50503, 16'd16495, 16'd57413, 16'd43073, 16'd35554, 16'd1912, 16'd35104});
	test_expansion(128'h73399b71cde1a02ed23840ff4250fb53, {16'd43542, 16'd34034, 16'd47381, 16'd5872, 16'd20360, 16'd43780, 16'd55664, 16'd7093, 16'd10858, 16'd65466, 16'd50272, 16'd27693, 16'd9118, 16'd28402, 16'd54004, 16'd17404, 16'd63643, 16'd6113, 16'd44689, 16'd56872, 16'd14796, 16'd134, 16'd64199, 16'd46490, 16'd15947, 16'd19147});
	test_expansion(128'h6fdc07b85ed6e74fa232a7af669f33c7, {16'd11390, 16'd31758, 16'd25924, 16'd56991, 16'd51857, 16'd61638, 16'd54455, 16'd50141, 16'd52801, 16'd43186, 16'd10472, 16'd31495, 16'd61213, 16'd65505, 16'd8993, 16'd62105, 16'd3066, 16'd5609, 16'd57669, 16'd2832, 16'd49293, 16'd19802, 16'd21387, 16'd30976, 16'd56599, 16'd45560});
	test_expansion(128'h9019b4198cdcaf98caf343fb4fb88002, {16'd12145, 16'd59393, 16'd12857, 16'd52895, 16'd22414, 16'd38342, 16'd26586, 16'd31387, 16'd17418, 16'd54385, 16'd7393, 16'd64814, 16'd12072, 16'd52132, 16'd25245, 16'd50387, 16'd19910, 16'd49159, 16'd8067, 16'd31845, 16'd16910, 16'd11941, 16'd685, 16'd13784, 16'd39992, 16'd63316});
	test_expansion(128'h35544ade79507f90306364c7ac1e1520, {16'd25866, 16'd1966, 16'd7827, 16'd21838, 16'd56526, 16'd8516, 16'd56151, 16'd46056, 16'd35267, 16'd43323, 16'd26751, 16'd50148, 16'd37404, 16'd14481, 16'd5072, 16'd64908, 16'd64062, 16'd32512, 16'd65491, 16'd3727, 16'd53019, 16'd37135, 16'd1455, 16'd3988, 16'd16032, 16'd55440});
	test_expansion(128'h6718c967a886ec1f9695942ea8fde51d, {16'd49808, 16'd20087, 16'd56384, 16'd59543, 16'd36753, 16'd16654, 16'd7972, 16'd58237, 16'd10803, 16'd64457, 16'd51320, 16'd17169, 16'd60008, 16'd36423, 16'd41205, 16'd63423, 16'd64755, 16'd57354, 16'd1462, 16'd43310, 16'd29271, 16'd4494, 16'd33761, 16'd63987, 16'd63726, 16'd63983});
	test_expansion(128'h60374e6927275eece98fbce382eac851, {16'd44854, 16'd2011, 16'd63280, 16'd30361, 16'd48652, 16'd48798, 16'd2974, 16'd4830, 16'd50274, 16'd42962, 16'd62, 16'd53300, 16'd51881, 16'd46140, 16'd61945, 16'd43632, 16'd11771, 16'd30169, 16'd25265, 16'd15812, 16'd25636, 16'd3821, 16'd58491, 16'd56364, 16'd53384, 16'd48153});
	test_expansion(128'hc31874b42e00ee25fb4fdaee3b27fafb, {16'd27717, 16'd4970, 16'd17046, 16'd16346, 16'd46678, 16'd14845, 16'd41109, 16'd3428, 16'd38120, 16'd29907, 16'd58759, 16'd28163, 16'd29697, 16'd9289, 16'd44330, 16'd59777, 16'd50668, 16'd61532, 16'd36151, 16'd11808, 16'd13966, 16'd36952, 16'd47561, 16'd49502, 16'd12386, 16'd7192});
	test_expansion(128'h370a12ed0759196d974b7cead7ec4687, {16'd64030, 16'd51977, 16'd13276, 16'd51515, 16'd40853, 16'd25386, 16'd1852, 16'd18156, 16'd48766, 16'd26672, 16'd21235, 16'd45384, 16'd42918, 16'd31623, 16'd7325, 16'd9716, 16'd29982, 16'd20919, 16'd20173, 16'd43428, 16'd58355, 16'd18301, 16'd8973, 16'd11768, 16'd59421, 16'd62848});
	test_expansion(128'he505f473551212b6387fc9dc5e6c3d34, {16'd40835, 16'd52731, 16'd13615, 16'd17387, 16'd53464, 16'd29144, 16'd3056, 16'd48099, 16'd43389, 16'd31815, 16'd24602, 16'd33835, 16'd57366, 16'd49985, 16'd5332, 16'd65484, 16'd29696, 16'd29967, 16'd3409, 16'd16636, 16'd49940, 16'd17695, 16'd8228, 16'd43166, 16'd59044, 16'd31134});
	test_expansion(128'h49424ad6060791ff939317b7d45a1a6a, {16'd59681, 16'd18154, 16'd49948, 16'd35478, 16'd59963, 16'd24715, 16'd19592, 16'd5384, 16'd7792, 16'd24245, 16'd27643, 16'd57793, 16'd21423, 16'd61223, 16'd41472, 16'd47022, 16'd20468, 16'd61716, 16'd25488, 16'd216, 16'd50376, 16'd51624, 16'd13883, 16'd50795, 16'd33157, 16'd38515});
	test_expansion(128'h092034a8fc2c5575f9fafcc21125c497, {16'd14858, 16'd40460, 16'd19325, 16'd18157, 16'd64405, 16'd5481, 16'd33628, 16'd47175, 16'd60235, 16'd61157, 16'd48229, 16'd8236, 16'd31921, 16'd20981, 16'd39122, 16'd63391, 16'd23912, 16'd46350, 16'd64348, 16'd46634, 16'd3488, 16'd57453, 16'd13655, 16'd13838, 16'd10156, 16'd6586});
	test_expansion(128'h2cc1fce76eb73423558d2ded72556d1b, {16'd4237, 16'd33544, 16'd5459, 16'd25307, 16'd44251, 16'd55428, 16'd43314, 16'd11160, 16'd2325, 16'd29252, 16'd16474, 16'd54300, 16'd44384, 16'd31417, 16'd44660, 16'd43555, 16'd40787, 16'd55579, 16'd21003, 16'd27, 16'd37608, 16'd28901, 16'd11953, 16'd12807, 16'd3051, 16'd1104});
	test_expansion(128'h98305feab76d7c5a931d50b3a9d923eb, {16'd53034, 16'd26207, 16'd47304, 16'd61501, 16'd6786, 16'd20497, 16'd5307, 16'd26833, 16'd58503, 16'd16119, 16'd58324, 16'd31710, 16'd7288, 16'd8976, 16'd57096, 16'd42428, 16'd53043, 16'd64918, 16'd43633, 16'd1858, 16'd9511, 16'd21231, 16'd33361, 16'd2340, 16'd34245, 16'd44043});
	test_expansion(128'h2a1633e04174815e43d84400f1e7bf80, {16'd55246, 16'd15355, 16'd17255, 16'd5126, 16'd55907, 16'd24140, 16'd37427, 16'd30144, 16'd58016, 16'd31978, 16'd27115, 16'd16279, 16'd35589, 16'd56368, 16'd2420, 16'd34279, 16'd29476, 16'd11962, 16'd23554, 16'd38106, 16'd5739, 16'd49597, 16'd34339, 16'd1726, 16'd18847, 16'd26264});
	test_expansion(128'he8c70d484e197be7442c3c80d6ddd37e, {16'd45601, 16'd4577, 16'd12371, 16'd40177, 16'd5672, 16'd1093, 16'd7044, 16'd33643, 16'd30791, 16'd64588, 16'd27242, 16'd13405, 16'd58987, 16'd6653, 16'd24351, 16'd3572, 16'd31823, 16'd47705, 16'd56766, 16'd31152, 16'd28670, 16'd24323, 16'd662, 16'd28054, 16'd51557, 16'd11669});
	test_expansion(128'h53782244d70c1681584beeb65e8d7083, {16'd58411, 16'd64897, 16'd2437, 16'd37860, 16'd61211, 16'd7133, 16'd63122, 16'd6253, 16'd53751, 16'd21199, 16'd14003, 16'd60672, 16'd63743, 16'd58618, 16'd58988, 16'd53498, 16'd53462, 16'd60013, 16'd40303, 16'd35983, 16'd29258, 16'd3028, 16'd46003, 16'd2892, 16'd300, 16'd35984});
	test_expansion(128'h08f0a73337c1001a2acbb47b55a66708, {16'd43404, 16'd44822, 16'd18310, 16'd46363, 16'd26097, 16'd59327, 16'd41989, 16'd43284, 16'd36535, 16'd38749, 16'd54254, 16'd10771, 16'd51102, 16'd21658, 16'd43177, 16'd14163, 16'd29419, 16'd12292, 16'd45782, 16'd40661, 16'd28260, 16'd5304, 16'd47135, 16'd62114, 16'd11793, 16'd13903});
	test_expansion(128'ha927ba21b0a4a831251d05923a63634b, {16'd59632, 16'd2486, 16'd40111, 16'd49032, 16'd18772, 16'd38762, 16'd54110, 16'd2907, 16'd35280, 16'd43951, 16'd40979, 16'd51265, 16'd60557, 16'd6879, 16'd4860, 16'd51291, 16'd62241, 16'd49518, 16'd27900, 16'd33121, 16'd37892, 16'd44840, 16'd64423, 16'd63427, 16'd42905, 16'd32465});
	test_expansion(128'h7e4fc3c36007f366a9e697ecb8d15992, {16'd58023, 16'd63714, 16'd53701, 16'd29277, 16'd34077, 16'd38259, 16'd10800, 16'd8304, 16'd53271, 16'd38886, 16'd42989, 16'd55202, 16'd11069, 16'd52001, 16'd37450, 16'd16324, 16'd24413, 16'd15896, 16'd55358, 16'd61890, 16'd11269, 16'd8507, 16'd61833, 16'd43407, 16'd649, 16'd7062});
	test_expansion(128'haf578ec7eab382708e4426ccc4604de9, {16'd39705, 16'd444, 16'd12398, 16'd3692, 16'd37639, 16'd59598, 16'd11831, 16'd57011, 16'd60420, 16'd917, 16'd32573, 16'd32484, 16'd62019, 16'd16724, 16'd1265, 16'd45292, 16'd54451, 16'd12680, 16'd55242, 16'd41573, 16'd50194, 16'd34360, 16'd5403, 16'd42736, 16'd52607, 16'd24681});
	test_expansion(128'h390fa44949eaef69f3087cb4eed68b94, {16'd30577, 16'd4567, 16'd59442, 16'd34415, 16'd19090, 16'd51150, 16'd9980, 16'd50146, 16'd27461, 16'd42259, 16'd56723, 16'd1104, 16'd43643, 16'd46317, 16'd44377, 16'd40384, 16'd25089, 16'd32163, 16'd15469, 16'd36245, 16'd28197, 16'd51940, 16'd62726, 16'd43423, 16'd11479, 16'd47274});
	test_expansion(128'ha046e08f18bc186a14beaf7b97eee132, {16'd38589, 16'd14643, 16'd31984, 16'd34676, 16'd9945, 16'd40816, 16'd21373, 16'd25630, 16'd54433, 16'd19211, 16'd13047, 16'd45239, 16'd45497, 16'd12683, 16'd45971, 16'd23904, 16'd25490, 16'd52236, 16'd14291, 16'd4598, 16'd12953, 16'd40446, 16'd43028, 16'd43152, 16'd37132, 16'd18585});
	test_expansion(128'he89977004d24863512adb7ab56a4a3fd, {16'd3384, 16'd58245, 16'd58743, 16'd12177, 16'd41091, 16'd11840, 16'd6535, 16'd27924, 16'd37716, 16'd56190, 16'd64467, 16'd54832, 16'd27020, 16'd2288, 16'd33580, 16'd4379, 16'd2435, 16'd7376, 16'd43104, 16'd18331, 16'd51076, 16'd51775, 16'd43879, 16'd63151, 16'd58668, 16'd33608});
	test_expansion(128'h35b663f62deb583541ceed5bbfcfc745, {16'd11963, 16'd58552, 16'd3013, 16'd16095, 16'd9867, 16'd8025, 16'd41834, 16'd58812, 16'd34256, 16'd39649, 16'd22643, 16'd54741, 16'd65243, 16'd49826, 16'd5134, 16'd47854, 16'd62573, 16'd43707, 16'd30372, 16'd22020, 16'd47705, 16'd27122, 16'd62262, 16'd18111, 16'd65473, 16'd62436});
	test_expansion(128'h344f8b7b914d4c9faaf25950784ba6e5, {16'd13810, 16'd54637, 16'd8324, 16'd37771, 16'd14713, 16'd37154, 16'd21847, 16'd22836, 16'd51204, 16'd45031, 16'd5839, 16'd26313, 16'd33308, 16'd25833, 16'd37389, 16'd29574, 16'd6901, 16'd61907, 16'd17424, 16'd4823, 16'd25456, 16'd28078, 16'd3894, 16'd44515, 16'd19902, 16'd54433});
	test_expansion(128'h1608c2b3fd71465b76fe0bdb122009e6, {16'd49378, 16'd38081, 16'd38407, 16'd17473, 16'd63747, 16'd36395, 16'd6436, 16'd61495, 16'd6712, 16'd14212, 16'd40475, 16'd33451, 16'd279, 16'd31808, 16'd62895, 16'd1908, 16'd52297, 16'd8395, 16'd49112, 16'd10263, 16'd29092, 16'd61224, 16'd1443, 16'd63407, 16'd42250, 16'd48581});
	test_expansion(128'h2d74f912db8252c4e6f99ef17d56d912, {16'd55416, 16'd94, 16'd12076, 16'd37466, 16'd42649, 16'd2018, 16'd17600, 16'd57167, 16'd1464, 16'd57171, 16'd41350, 16'd55153, 16'd61954, 16'd11805, 16'd38034, 16'd19647, 16'd61701, 16'd53046, 16'd10611, 16'd63594, 16'd18968, 16'd29072, 16'd29325, 16'd53566, 16'd33005, 16'd38391});
	test_expansion(128'hbeaa449126d4a1c5738282361b3488ed, {16'd62931, 16'd7573, 16'd62017, 16'd53617, 16'd30105, 16'd7194, 16'd12295, 16'd5747, 16'd5988, 16'd16449, 16'd13473, 16'd35233, 16'd15960, 16'd12297, 16'd19916, 16'd57863, 16'd43563, 16'd42091, 16'd9170, 16'd37796, 16'd53356, 16'd42469, 16'd40576, 16'd21233, 16'd6790, 16'd59386});
	test_expansion(128'hd213a2041387de5c5f527d7b2f6b7fc7, {16'd3040, 16'd23088, 16'd11976, 16'd53503, 16'd3540, 16'd31628, 16'd48601, 16'd53042, 16'd12233, 16'd20348, 16'd44729, 16'd11870, 16'd47901, 16'd64549, 16'd2834, 16'd10768, 16'd5665, 16'd55136, 16'd7237, 16'd2, 16'd13298, 16'd44545, 16'd52085, 16'd39229, 16'd36197, 16'd45529});
	test_expansion(128'h52f8909cc15cc6ed5ef86df54a4b151c, {16'd24819, 16'd9863, 16'd62739, 16'd60930, 16'd2826, 16'd62013, 16'd45173, 16'd56177, 16'd14245, 16'd61232, 16'd45032, 16'd58830, 16'd2312, 16'd25079, 16'd3498, 16'd44868, 16'd51116, 16'd34447, 16'd13465, 16'd54439, 16'd5519, 16'd21002, 16'd18305, 16'd63645, 16'd59342, 16'd33810});
	test_expansion(128'h12a4a8057eba9576ac2f6988f0075012, {16'd22742, 16'd58553, 16'd36779, 16'd55314, 16'd48235, 16'd59452, 16'd24603, 16'd1401, 16'd42199, 16'd20283, 16'd5616, 16'd48880, 16'd55343, 16'd18270, 16'd7078, 16'd1114, 16'd46028, 16'd13969, 16'd3733, 16'd37076, 16'd15722, 16'd10402, 16'd25783, 16'd27104, 16'd6158, 16'd15379});
	test_expansion(128'hfd92abfb5917754ca01fa29f58f1ad7c, {16'd50934, 16'd14084, 16'd58023, 16'd16099, 16'd61032, 16'd52655, 16'd64249, 16'd17407, 16'd47117, 16'd19192, 16'd20379, 16'd48420, 16'd58099, 16'd27605, 16'd49291, 16'd26288, 16'd48043, 16'd47984, 16'd54532, 16'd32067, 16'd60506, 16'd60192, 16'd38959, 16'd27022, 16'd6266, 16'd44414});
	test_expansion(128'h030c8903983c978cece32d7204763e29, {16'd15561, 16'd776, 16'd8998, 16'd32565, 16'd61419, 16'd16057, 16'd43031, 16'd11486, 16'd8408, 16'd63881, 16'd53179, 16'd19620, 16'd23271, 16'd1613, 16'd51492, 16'd28539, 16'd17452, 16'd29947, 16'd37788, 16'd42976, 16'd27962, 16'd31940, 16'd6662, 16'd50107, 16'd24051, 16'd57900});
	test_expansion(128'hca2a9271d3e01662fb646565778f8eb8, {16'd64998, 16'd50335, 16'd22470, 16'd23300, 16'd40713, 16'd13957, 16'd14163, 16'd60602, 16'd27537, 16'd15552, 16'd57006, 16'd28150, 16'd41680, 16'd38100, 16'd8818, 16'd11809, 16'd923, 16'd20238, 16'd41988, 16'd44680, 16'd6708, 16'd21789, 16'd24874, 16'd50504, 16'd56066, 16'd24892});
	test_expansion(128'hac3bf9a76f6f9834af755d4e7aa9a1df, {16'd45010, 16'd14058, 16'd31985, 16'd61483, 16'd11451, 16'd54173, 16'd10093, 16'd24223, 16'd29344, 16'd4483, 16'd55716, 16'd33233, 16'd38607, 16'd19131, 16'd28820, 16'd63799, 16'd63232, 16'd43560, 16'd54134, 16'd54078, 16'd57239, 16'd28202, 16'd59481, 16'd60251, 16'd48416, 16'd44570});
	test_expansion(128'he62e372156299669e3de658143f448b6, {16'd14590, 16'd22736, 16'd23501, 16'd35431, 16'd38843, 16'd17895, 16'd23988, 16'd59389, 16'd4412, 16'd15786, 16'd857, 16'd22690, 16'd7645, 16'd36223, 16'd47136, 16'd33702, 16'd13309, 16'd6793, 16'd60602, 16'd15983, 16'd20003, 16'd23957, 16'd61310, 16'd8166, 16'd5755, 16'd49071});
	test_expansion(128'hc86561aa0021249e460092e60660af4a, {16'd14434, 16'd688, 16'd32538, 16'd9205, 16'd39580, 16'd58291, 16'd58355, 16'd12734, 16'd44606, 16'd34774, 16'd47872, 16'd50700, 16'd30695, 16'd24369, 16'd33541, 16'd64360, 16'd17638, 16'd50881, 16'd9789, 16'd22740, 16'd60654, 16'd28228, 16'd10825, 16'd48985, 16'd23743, 16'd63659});
	test_expansion(128'h354938d62b4adfe4dd3dec1b2cb70765, {16'd15549, 16'd6566, 16'd13543, 16'd25686, 16'd19379, 16'd9441, 16'd19498, 16'd14598, 16'd11040, 16'd52849, 16'd26275, 16'd27961, 16'd1743, 16'd15200, 16'd24157, 16'd12411, 16'd64104, 16'd62806, 16'd34274, 16'd2122, 16'd43263, 16'd11547, 16'd36156, 16'd5340, 16'd45284, 16'd20114});
	test_expansion(128'h8894483375063a58e7426d19bfb3f814, {16'd35964, 16'd31735, 16'd57017, 16'd19830, 16'd51410, 16'd56951, 16'd1808, 16'd6659, 16'd63057, 16'd40957, 16'd60424, 16'd658, 16'd57202, 16'd64656, 16'd43637, 16'd39605, 16'd18602, 16'd1702, 16'd25511, 16'd14988, 16'd28816, 16'd11881, 16'd39436, 16'd27539, 16'd6776, 16'd6191});
	test_expansion(128'h73a939077005f4869b73ad0004cb68a2, {16'd24664, 16'd52459, 16'd32535, 16'd5047, 16'd16036, 16'd4234, 16'd21095, 16'd34059, 16'd48851, 16'd61845, 16'd13467, 16'd59536, 16'd21994, 16'd3330, 16'd56691, 16'd42008, 16'd61021, 16'd48654, 16'd51928, 16'd31726, 16'd16660, 16'd57462, 16'd55757, 16'd33800, 16'd33388, 16'd57912});
	test_expansion(128'hee1d9e8f47e65d01057c49d9fdfa580e, {16'd46444, 16'd55796, 16'd62602, 16'd37599, 16'd20936, 16'd34230, 16'd32932, 16'd30523, 16'd28201, 16'd8916, 16'd4532, 16'd6527, 16'd17271, 16'd62873, 16'd56606, 16'd44544, 16'd26186, 16'd12796, 16'd15005, 16'd42885, 16'd18848, 16'd37535, 16'd10142, 16'd46482, 16'd52882, 16'd25582});
	test_expansion(128'h45c85cd6971521ecc1d75229da5199d7, {16'd40122, 16'd17259, 16'd41301, 16'd12354, 16'd33466, 16'd47757, 16'd44567, 16'd27160, 16'd57010, 16'd53092, 16'd3351, 16'd24813, 16'd63663, 16'd32071, 16'd50991, 16'd3051, 16'd18981, 16'd23782, 16'd44394, 16'd46721, 16'd57037, 16'd6794, 16'd2450, 16'd16038, 16'd12057, 16'd49880});
	test_expansion(128'he54bd753c645afa75656829c579ea4e3, {16'd7303, 16'd5858, 16'd40990, 16'd25656, 16'd26016, 16'd40789, 16'd10873, 16'd15628, 16'd2203, 16'd49107, 16'd26379, 16'd21093, 16'd14494, 16'd1711, 16'd36648, 16'd55890, 16'd43115, 16'd8876, 16'd48553, 16'd65039, 16'd44840, 16'd4075, 16'd15170, 16'd25952, 16'd4050, 16'd54568});
	test_expansion(128'hb73fbe72b591be6b4aed1dd05c00de44, {16'd304, 16'd56944, 16'd55429, 16'd48955, 16'd52986, 16'd6813, 16'd27253, 16'd44399, 16'd19573, 16'd57913, 16'd33422, 16'd32712, 16'd46116, 16'd48604, 16'd52475, 16'd18054, 16'd39503, 16'd58323, 16'd56131, 16'd60742, 16'd24344, 16'd62562, 16'd52207, 16'd38115, 16'd14804, 16'd22971});
	test_expansion(128'h5e97570682cf63f2a293f6f10933ec9a, {16'd1181, 16'd21831, 16'd18065, 16'd43711, 16'd13315, 16'd39192, 16'd21482, 16'd1321, 16'd41273, 16'd58109, 16'd58895, 16'd58338, 16'd12849, 16'd35888, 16'd20562, 16'd16834, 16'd9015, 16'd54710, 16'd2619, 16'd51469, 16'd62099, 16'd22864, 16'd48495, 16'd25215, 16'd44950, 16'd56138});
	test_expansion(128'hba8e20b510ecd70b4c23cca26bfe57c9, {16'd15875, 16'd402, 16'd45211, 16'd53845, 16'd12493, 16'd50122, 16'd59001, 16'd62814, 16'd10791, 16'd63012, 16'd64954, 16'd39182, 16'd45134, 16'd11266, 16'd31451, 16'd4254, 16'd25803, 16'd62427, 16'd54208, 16'd51133, 16'd10030, 16'd61024, 16'd36147, 16'd59428, 16'd2015, 16'd43760});
	test_expansion(128'h97a977e7ef8681bf14d3a854a3d060f4, {16'd4632, 16'd3852, 16'd34928, 16'd37865, 16'd37146, 16'd60840, 16'd30307, 16'd62595, 16'd20095, 16'd43910, 16'd48155, 16'd5006, 16'd39827, 16'd22790, 16'd35580, 16'd4597, 16'd28918, 16'd934, 16'd1637, 16'd10246, 16'd15746, 16'd30443, 16'd59833, 16'd47679, 16'd15017, 16'd58023});
	test_expansion(128'h288f36611d892cb841e0cfa4cac79a7b, {16'd56581, 16'd11935, 16'd30680, 16'd36854, 16'd27263, 16'd38592, 16'd3691, 16'd3811, 16'd26218, 16'd49292, 16'd22858, 16'd8034, 16'd4987, 16'd8782, 16'd40319, 16'd58207, 16'd42788, 16'd14749, 16'd31904, 16'd3658, 16'd47786, 16'd42219, 16'd62450, 16'd10645, 16'd25517, 16'd23313});
	test_expansion(128'he0906daaae06a16c0123247e20d9cc05, {16'd26491, 16'd13880, 16'd1033, 16'd2610, 16'd41315, 16'd46240, 16'd17774, 16'd60460, 16'd3377, 16'd19138, 16'd22863, 16'd64374, 16'd49593, 16'd53362, 16'd57752, 16'd61614, 16'd47440, 16'd32153, 16'd39518, 16'd16967, 16'd18526, 16'd38628, 16'd60157, 16'd62870, 16'd13260, 16'd65315});
	test_expansion(128'h0f03e986fee779fd109e81d0bae63c12, {16'd6080, 16'd26555, 16'd61148, 16'd2559, 16'd3198, 16'd6852, 16'd22672, 16'd7336, 16'd41891, 16'd10371, 16'd50747, 16'd42832, 16'd35710, 16'd16603, 16'd24348, 16'd15839, 16'd61065, 16'd19038, 16'd20032, 16'd47146, 16'd49403, 16'd61513, 16'd37870, 16'd28817, 16'd51852, 16'd25449});
	test_expansion(128'h9faffca1f270c8aaa7bc3300db061bac, {16'd21874, 16'd41433, 16'd45511, 16'd65156, 16'd65355, 16'd57846, 16'd46167, 16'd27141, 16'd17968, 16'd22707, 16'd55440, 16'd31295, 16'd1634, 16'd58346, 16'd7936, 16'd6020, 16'd27777, 16'd50293, 16'd53620, 16'd33916, 16'd54235, 16'd3483, 16'd59599, 16'd27039, 16'd2223, 16'd18130});
	test_expansion(128'he5733be26055e19f669f3cd2605d0fba, {16'd35813, 16'd50153, 16'd6669, 16'd59372, 16'd43395, 16'd20189, 16'd35779, 16'd27321, 16'd42056, 16'd39610, 16'd4051, 16'd62621, 16'd36950, 16'd34740, 16'd56748, 16'd35755, 16'd1579, 16'd62014, 16'd58972, 16'd46537, 16'd25494, 16'd10666, 16'd17001, 16'd7272, 16'd17638, 16'd17911});
	test_expansion(128'had0f375086021b36cf93356da7ee556a, {16'd5577, 16'd41189, 16'd24322, 16'd7120, 16'd33530, 16'd32601, 16'd5276, 16'd14895, 16'd11993, 16'd18406, 16'd29558, 16'd39296, 16'd46267, 16'd29839, 16'd29600, 16'd48195, 16'd11576, 16'd44522, 16'd51338, 16'd44411, 16'd1584, 16'd64203, 16'd17178, 16'd60581, 16'd5899, 16'd61289});
	test_expansion(128'h2a424dd23d54be1b38ff5df589d42c58, {16'd45051, 16'd26017, 16'd20439, 16'd60490, 16'd544, 16'd14009, 16'd41744, 16'd61955, 16'd816, 16'd59619, 16'd16501, 16'd62938, 16'd40907, 16'd12985, 16'd33401, 16'd24905, 16'd47732, 16'd59583, 16'd24244, 16'd26460, 16'd46730, 16'd49304, 16'd58052, 16'd28496, 16'd62400, 16'd47096});
	test_expansion(128'h6245405945a9c32b613da52c0c75eb23, {16'd25727, 16'd44316, 16'd11766, 16'd48590, 16'd34599, 16'd59702, 16'd10257, 16'd61098, 16'd51962, 16'd5932, 16'd28295, 16'd28199, 16'd33856, 16'd39314, 16'd54720, 16'd62657, 16'd6694, 16'd36319, 16'd13148, 16'd19941, 16'd5830, 16'd33180, 16'd54151, 16'd41341, 16'd19554, 16'd24343});
	test_expansion(128'h85281ae6716d2c659bf24434e76d3c04, {16'd15879, 16'd14898, 16'd55131, 16'd35411, 16'd31538, 16'd51347, 16'd63005, 16'd35566, 16'd5439, 16'd257, 16'd423, 16'd18401, 16'd47461, 16'd5705, 16'd60846, 16'd15924, 16'd14818, 16'd12158, 16'd6973, 16'd10528, 16'd22547, 16'd57275, 16'd46316, 16'd4837, 16'd26902, 16'd11611});
	test_expansion(128'h43b2c3c342e84a1a0ccd9f3962abca22, {16'd29597, 16'd7363, 16'd2215, 16'd19615, 16'd40962, 16'd24262, 16'd865, 16'd8198, 16'd30167, 16'd19895, 16'd23246, 16'd36171, 16'd65463, 16'd50395, 16'd45040, 16'd51861, 16'd21651, 16'd47514, 16'd62816, 16'd38900, 16'd33091, 16'd20162, 16'd24445, 16'd57596, 16'd44056, 16'd14798});
	test_expansion(128'h67d23a307eb5b867a0881ecdc1fea0fe, {16'd21044, 16'd6418, 16'd26418, 16'd6006, 16'd572, 16'd31202, 16'd54467, 16'd45327, 16'd8168, 16'd56536, 16'd10722, 16'd23639, 16'd25663, 16'd56902, 16'd48606, 16'd46176, 16'd46611, 16'd38954, 16'd41205, 16'd3398, 16'd24107, 16'd46342, 16'd33835, 16'd40266, 16'd35921, 16'd1541});
	test_expansion(128'h32efae199c8fa227d98031dca829673e, {16'd57749, 16'd40902, 16'd49600, 16'd22963, 16'd40576, 16'd7257, 16'd57102, 16'd39979, 16'd12762, 16'd21179, 16'd649, 16'd35536, 16'd63613, 16'd36378, 16'd30888, 16'd1845, 16'd27621, 16'd53102, 16'd47954, 16'd19450, 16'd11467, 16'd4784, 16'd13880, 16'd35656, 16'd47143, 16'd1514});
	test_expansion(128'h333a0f3e142c66144ec468ab04d9ffb8, {16'd57455, 16'd10745, 16'd49849, 16'd6683, 16'd44467, 16'd61428, 16'd45505, 16'd38147, 16'd5368, 16'd54479, 16'd44247, 16'd54524, 16'd61853, 16'd51546, 16'd59078, 16'd31162, 16'd43536, 16'd48783, 16'd15865, 16'd43254, 16'd25370, 16'd9399, 16'd55598, 16'd54346, 16'd1885, 16'd12960});
	test_expansion(128'h51ec816d3d4313177d8cd7ba7370524f, {16'd42408, 16'd20000, 16'd25152, 16'd44236, 16'd20350, 16'd61591, 16'd60806, 16'd62792, 16'd46586, 16'd11530, 16'd37154, 16'd51588, 16'd53282, 16'd14813, 16'd47010, 16'd63652, 16'd15227, 16'd122, 16'd50011, 16'd32209, 16'd52211, 16'd35880, 16'd64431, 16'd941, 16'd29299, 16'd15482});
	test_expansion(128'h136245883ca74ff8980ebb2d99d62049, {16'd33152, 16'd21310, 16'd26022, 16'd40974, 16'd50379, 16'd8567, 16'd47629, 16'd9922, 16'd50556, 16'd22864, 16'd37029, 16'd29902, 16'd2008, 16'd27465, 16'd22964, 16'd38960, 16'd41281, 16'd11195, 16'd29399, 16'd45826, 16'd17580, 16'd46497, 16'd59995, 16'd43901, 16'd36214, 16'd55687});
	test_expansion(128'h3c43dd4c1629df02e99c7b8eca42fb14, {16'd40789, 16'd59227, 16'd62088, 16'd25134, 16'd15789, 16'd43396, 16'd29344, 16'd804, 16'd29033, 16'd64399, 16'd64473, 16'd37150, 16'd58595, 16'd60519, 16'd28705, 16'd764, 16'd23087, 16'd1015, 16'd63563, 16'd62594, 16'd4180, 16'd43429, 16'd30111, 16'd52709, 16'd42945, 16'd18691});
	test_expansion(128'h1e24595eea98fa47c91f47ecb3c13d54, {16'd55333, 16'd34122, 16'd11967, 16'd43891, 16'd29932, 16'd49155, 16'd1627, 16'd32679, 16'd61253, 16'd31609, 16'd34996, 16'd51252, 16'd17987, 16'd46790, 16'd10824, 16'd401, 16'd56555, 16'd50595, 16'd3715, 16'd32489, 16'd49266, 16'd54865, 16'd25671, 16'd52459, 16'd372, 16'd3919});
	test_expansion(128'hce98146ce0179a040983631deb88df3a, {16'd57986, 16'd13636, 16'd63420, 16'd33454, 16'd53104, 16'd21577, 16'd4238, 16'd64929, 16'd58617, 16'd40622, 16'd47151, 16'd53065, 16'd58333, 16'd2644, 16'd1423, 16'd5687, 16'd27650, 16'd1458, 16'd32844, 16'd53552, 16'd50647, 16'd20975, 16'd21469, 16'd60306, 16'd34870, 16'd24718});
	test_expansion(128'ha235e01a83f09c4d8a05cf1882b1b3b4, {16'd21356, 16'd36365, 16'd29352, 16'd2623, 16'd55525, 16'd28427, 16'd31892, 16'd18073, 16'd21165, 16'd18864, 16'd46259, 16'd35186, 16'd24421, 16'd33602, 16'd46154, 16'd10685, 16'd7192, 16'd57644, 16'd6624, 16'd58834, 16'd35250, 16'd41385, 16'd60537, 16'd27634, 16'd20207, 16'd56914});
	test_expansion(128'hc3f077e69be3d31090ea24eef7ab8541, {16'd34959, 16'd43451, 16'd35623, 16'd59396, 16'd32979, 16'd27038, 16'd1387, 16'd35624, 16'd49920, 16'd65523, 16'd42276, 16'd38517, 16'd7493, 16'd35642, 16'd44924, 16'd59815, 16'd4537, 16'd58804, 16'd47713, 16'd25878, 16'd43476, 16'd34565, 16'd47684, 16'd12020, 16'd22038, 16'd30313});
	test_expansion(128'hd2ab8719b3c0b061c7b827db70703538, {16'd21806, 16'd44726, 16'd57456, 16'd57785, 16'd42848, 16'd36839, 16'd61024, 16'd46442, 16'd9290, 16'd36671, 16'd63234, 16'd33683, 16'd27746, 16'd62009, 16'd36409, 16'd46301, 16'd23553, 16'd34085, 16'd26304, 16'd61548, 16'd60152, 16'd6334, 16'd22272, 16'd65065, 16'd43044, 16'd43450});
	test_expansion(128'h47ce9905d74ad90a879b752d74c0028b, {16'd45131, 16'd56812, 16'd62807, 16'd15843, 16'd10117, 16'd42201, 16'd16639, 16'd29860, 16'd9467, 16'd38933, 16'd7985, 16'd46438, 16'd5343, 16'd10713, 16'd6151, 16'd892, 16'd13231, 16'd58753, 16'd25432, 16'd55419, 16'd21067, 16'd29958, 16'd746, 16'd53762, 16'd52732, 16'd18920});
	test_expansion(128'hf28362e0940bb2b1ee16bda2ce1fb3ba, {16'd1089, 16'd5313, 16'd51683, 16'd16382, 16'd19604, 16'd53726, 16'd17856, 16'd35608, 16'd39817, 16'd1473, 16'd35962, 16'd3746, 16'd53718, 16'd1856, 16'd4227, 16'd50680, 16'd22813, 16'd51883, 16'd48955, 16'd40193, 16'd49753, 16'd32831, 16'd7828, 16'd64661, 16'd33674, 16'd55278});
	test_expansion(128'ha95ac6dac5dda17d9f988d7dd3dbde5c, {16'd56990, 16'd39645, 16'd58714, 16'd62357, 16'd47593, 16'd5223, 16'd25823, 16'd34628, 16'd38943, 16'd49183, 16'd14240, 16'd24050, 16'd56996, 16'd56978, 16'd45028, 16'd8673, 16'd24757, 16'd56310, 16'd52684, 16'd45200, 16'd11533, 16'd58345, 16'd22117, 16'd48843, 16'd36937, 16'd48578});
	test_expansion(128'hbade0cdd487ec101e457d69f3ee74c2e, {16'd28381, 16'd43413, 16'd34549, 16'd30099, 16'd37585, 16'd28483, 16'd49977, 16'd22954, 16'd59719, 16'd18536, 16'd21401, 16'd7932, 16'd27993, 16'd7426, 16'd63411, 16'd49630, 16'd21583, 16'd32315, 16'd39865, 16'd31350, 16'd38579, 16'd51709, 16'd16068, 16'd18276, 16'd27579, 16'd8358});
	test_expansion(128'hfcfb73f0af6b47b0fc0d89fdab9f4c90, {16'd13145, 16'd12634, 16'd54089, 16'd26160, 16'd44134, 16'd6936, 16'd59891, 16'd35377, 16'd53213, 16'd27857, 16'd53372, 16'd54689, 16'd52421, 16'd59911, 16'd10432, 16'd22530, 16'd2451, 16'd28971, 16'd40890, 16'd21504, 16'd46412, 16'd7866, 16'd57551, 16'd46932, 16'd7928, 16'd27846});
	test_expansion(128'ha6cf8124a2b2365dca8efcc733ecb9a5, {16'd25488, 16'd41787, 16'd15257, 16'd12191, 16'd48403, 16'd15880, 16'd15431, 16'd33656, 16'd9146, 16'd32621, 16'd40368, 16'd64014, 16'd8604, 16'd26235, 16'd48510, 16'd13922, 16'd61429, 16'd61000, 16'd61841, 16'd27200, 16'd59975, 16'd21215, 16'd27593, 16'd46124, 16'd29342, 16'd35330});
	test_expansion(128'hfceb57437b107dc00f84837c647a21e4, {16'd22774, 16'd59107, 16'd59168, 16'd57073, 16'd65405, 16'd11362, 16'd60496, 16'd3655, 16'd52421, 16'd58088, 16'd38247, 16'd51545, 16'd61895, 16'd47226, 16'd49807, 16'd14584, 16'd33474, 16'd6849, 16'd39970, 16'd51481, 16'd64773, 16'd59043, 16'd45538, 16'd55050, 16'd50059, 16'd46009});
	test_expansion(128'h6c20473431f7f38f266542b605edf69f, {16'd22181, 16'd43984, 16'd37862, 16'd45988, 16'd8227, 16'd13160, 16'd21021, 16'd63153, 16'd49026, 16'd53036, 16'd19091, 16'd4261, 16'd8359, 16'd33320, 16'd62922, 16'd63516, 16'd64887, 16'd35409, 16'd3910, 16'd6494, 16'd35055, 16'd47412, 16'd33985, 16'd28421, 16'd11874, 16'd54531});
	test_expansion(128'h80c98ebe12129f51f318179a471ca295, {16'd41165, 16'd37286, 16'd37847, 16'd50815, 16'd5480, 16'd61808, 16'd63435, 16'd58963, 16'd16720, 16'd36787, 16'd51007, 16'd38812, 16'd44589, 16'd28186, 16'd44281, 16'd5348, 16'd3202, 16'd30073, 16'd768, 16'd6499, 16'd16633, 16'd14431, 16'd11255, 16'd16861, 16'd44383, 16'd6371});
	test_expansion(128'hac84b61e9ef399307cf8a34112ce6dae, {16'd36271, 16'd56604, 16'd4355, 16'd21555, 16'd58133, 16'd48844, 16'd32126, 16'd17479, 16'd44347, 16'd50038, 16'd252, 16'd30623, 16'd17565, 16'd48703, 16'd58039, 16'd44569, 16'd47032, 16'd50021, 16'd11987, 16'd28117, 16'd2021, 16'd59243, 16'd50368, 16'd41151, 16'd6359, 16'd21026});
	test_expansion(128'he1f1187475d0a2686f3a73432c82107e, {16'd25082, 16'd41007, 16'd61797, 16'd59548, 16'd33056, 16'd26568, 16'd39218, 16'd47430, 16'd14499, 16'd40623, 16'd27151, 16'd1722, 16'd59412, 16'd23902, 16'd53927, 16'd61670, 16'd26074, 16'd41080, 16'd29885, 16'd19412, 16'd22534, 16'd61317, 16'd37187, 16'd64921, 16'd49805, 16'd34703});
	test_expansion(128'hb768aad6e4b1c7b4a4a5fcb1d135c5a6, {16'd51240, 16'd3308, 16'd3180, 16'd54516, 16'd50312, 16'd57899, 16'd13208, 16'd37637, 16'd53987, 16'd34685, 16'd58719, 16'd3703, 16'd32228, 16'd60681, 16'd29229, 16'd43363, 16'd31393, 16'd7028, 16'd25973, 16'd23379, 16'd47110, 16'd26524, 16'd59932, 16'd2336, 16'd7019, 16'd25505});
	test_expansion(128'hdd65c21dd89535584458bcfbaeb00c5d, {16'd60942, 16'd9617, 16'd18831, 16'd723, 16'd23154, 16'd47266, 16'd4733, 16'd41827, 16'd1032, 16'd52042, 16'd22003, 16'd17246, 16'd38774, 16'd204, 16'd7350, 16'd17134, 16'd17988, 16'd4518, 16'd43257, 16'd46196, 16'd61321, 16'd16745, 16'd61524, 16'd3902, 16'd23881, 16'd35508});
	test_expansion(128'h769239dcbef79dfa5afd86c1bb632b1c, {16'd32138, 16'd19440, 16'd29248, 16'd17977, 16'd39829, 16'd44761, 16'd13421, 16'd37489, 16'd45946, 16'd60452, 16'd60991, 16'd24844, 16'd55161, 16'd2039, 16'd29660, 16'd15476, 16'd45938, 16'd44263, 16'd11405, 16'd55672, 16'd40116, 16'd27383, 16'd52817, 16'd41079, 16'd42128, 16'd41211});
	test_expansion(128'h3f6f700a5db4dd2811f7bc161ba273ec, {16'd16871, 16'd7821, 16'd59902, 16'd26052, 16'd64887, 16'd58763, 16'd46015, 16'd57006, 16'd33569, 16'd8967, 16'd9807, 16'd35334, 16'd1503, 16'd56818, 16'd60947, 16'd11390, 16'd36620, 16'd8157, 16'd17024, 16'd13990, 16'd1640, 16'd31696, 16'd12127, 16'd28303, 16'd20391, 16'd64848});
	test_expansion(128'h2999fc0be2bb5b755f4159d84776eb06, {16'd35173, 16'd2682, 16'd46549, 16'd5854, 16'd37776, 16'd18336, 16'd36560, 16'd15212, 16'd28388, 16'd63937, 16'd50294, 16'd5063, 16'd28776, 16'd19746, 16'd58453, 16'd63884, 16'd56593, 16'd13586, 16'd53329, 16'd53933, 16'd47475, 16'd55349, 16'd24140, 16'd4397, 16'd12446, 16'd20928});
	test_expansion(128'h0014909f1d73906c6023377c2408d6e0, {16'd57346, 16'd21532, 16'd26409, 16'd62348, 16'd22686, 16'd39513, 16'd11688, 16'd2779, 16'd11894, 16'd24443, 16'd41512, 16'd32246, 16'd29320, 16'd42251, 16'd63510, 16'd35962, 16'd63074, 16'd31833, 16'd61353, 16'd28652, 16'd27373, 16'd54665, 16'd49089, 16'd18251, 16'd22517, 16'd51518});
	test_expansion(128'h5ca5df27c29e6597b008927954394585, {16'd32487, 16'd61545, 16'd46365, 16'd36448, 16'd41567, 16'd8682, 16'd3165, 16'd59360, 16'd24216, 16'd30994, 16'd36263, 16'd29372, 16'd25315, 16'd29678, 16'd48907, 16'd10224, 16'd18918, 16'd18238, 16'd35148, 16'd14542, 16'd4536, 16'd30487, 16'd20728, 16'd55680, 16'd50964, 16'd9739});
	test_expansion(128'ha73186d405655df6e55eddf8bf0c5e2a, {16'd22765, 16'd50334, 16'd2683, 16'd20082, 16'd29896, 16'd12554, 16'd16646, 16'd996, 16'd12011, 16'd34560, 16'd39119, 16'd9851, 16'd44857, 16'd64660, 16'd59754, 16'd42866, 16'd36881, 16'd62825, 16'd56316, 16'd43581, 16'd29627, 16'd40799, 16'd26126, 16'd41919, 16'd25215, 16'd22360});
	test_expansion(128'h129d8aaaa99cbc9a0006afb94b5236d9, {16'd47495, 16'd29927, 16'd55537, 16'd46457, 16'd46664, 16'd54411, 16'd7452, 16'd25439, 16'd50521, 16'd57214, 16'd59585, 16'd30150, 16'd48482, 16'd60000, 16'd24218, 16'd62255, 16'd48382, 16'd30283, 16'd10178, 16'd63257, 16'd15367, 16'd17446, 16'd34901, 16'd30953, 16'd12167, 16'd5419});
	test_expansion(128'h1cdb3534616c48045a6db13814e1a24a, {16'd59718, 16'd12366, 16'd62894, 16'd19320, 16'd20910, 16'd31536, 16'd53726, 16'd62952, 16'd39809, 16'd18090, 16'd53331, 16'd1978, 16'd40963, 16'd13995, 16'd1115, 16'd42606, 16'd45575, 16'd41343, 16'd60085, 16'd61055, 16'd59509, 16'd5268, 16'd26337, 16'd11367, 16'd28791, 16'd6639});
	test_expansion(128'he245226522ca3cf833325f53bf733000, {16'd11681, 16'd11020, 16'd40911, 16'd9917, 16'd60426, 16'd22596, 16'd35099, 16'd945, 16'd21128, 16'd23292, 16'd3702, 16'd6451, 16'd32824, 16'd11511, 16'd59821, 16'd45326, 16'd36736, 16'd10080, 16'd46544, 16'd25054, 16'd22158, 16'd50455, 16'd44169, 16'd7302, 16'd30258, 16'd24212});
	test_expansion(128'h9b1aba00e898c196fe94b436dd95d69e, {16'd64641, 16'd23197, 16'd29659, 16'd37432, 16'd25871, 16'd51253, 16'd38534, 16'd41067, 16'd11586, 16'd60285, 16'd2804, 16'd56544, 16'd4747, 16'd24434, 16'd26217, 16'd30393, 16'd41852, 16'd17720, 16'd62111, 16'd58282, 16'd2110, 16'd32988, 16'd13062, 16'd3269, 16'd39326, 16'd35476});
	test_expansion(128'h2f28cb4fc4e334ec5830ce043b74f699, {16'd2628, 16'd64893, 16'd57712, 16'd616, 16'd33213, 16'd34385, 16'd7242, 16'd29905, 16'd10967, 16'd10048, 16'd35358, 16'd44544, 16'd39806, 16'd16082, 16'd34184, 16'd54284, 16'd44760, 16'd24791, 16'd4350, 16'd61204, 16'd16331, 16'd13450, 16'd39902, 16'd28737, 16'd46781, 16'd37429});
	test_expansion(128'h3b7905f5a930b3ff95d9ed2f10f88358, {16'd36249, 16'd61039, 16'd46728, 16'd54845, 16'd43692, 16'd11971, 16'd20302, 16'd38858, 16'd1505, 16'd9082, 16'd24814, 16'd9752, 16'd54857, 16'd10049, 16'd49782, 16'd15889, 16'd17624, 16'd55876, 16'd34863, 16'd4358, 16'd44314, 16'd10166, 16'd52557, 16'd28899, 16'd21490, 16'd30286});
	test_expansion(128'hc7bbc1984d4c32ab49f5c1881e179570, {16'd3444, 16'd61426, 16'd58207, 16'd13673, 16'd8679, 16'd47238, 16'd48525, 16'd56612, 16'd41464, 16'd37252, 16'd23778, 16'd4153, 16'd15808, 16'd52485, 16'd39231, 16'd23418, 16'd27174, 16'd17169, 16'd35929, 16'd55696, 16'd9406, 16'd10861, 16'd48980, 16'd38687, 16'd25678, 16'd20353});
	test_expansion(128'h3ff7933bec70355a48bc0a187cf6b048, {16'd21316, 16'd28419, 16'd20436, 16'd3251, 16'd41334, 16'd51778, 16'd48157, 16'd12859, 16'd51866, 16'd33166, 16'd62030, 16'd26495, 16'd9646, 16'd8450, 16'd50055, 16'd43159, 16'd6389, 16'd16671, 16'd7048, 16'd41351, 16'd19910, 16'd58840, 16'd38823, 16'd12117, 16'd29588, 16'd14665});
	test_expansion(128'hd4ae202895ceb578649e2dbbea428708, {16'd30958, 16'd24954, 16'd472, 16'd60945, 16'd49658, 16'd28145, 16'd1457, 16'd60133, 16'd44712, 16'd40417, 16'd24648, 16'd46998, 16'd51109, 16'd58215, 16'd54729, 16'd34374, 16'd31776, 16'd54400, 16'd57293, 16'd41197, 16'd29053, 16'd59285, 16'd58027, 16'd2095, 16'd57587, 16'd9188});
	test_expansion(128'h8d2a6ca8097c4351f900f1c6f66b29c1, {16'd53363, 16'd63769, 16'd27075, 16'd55750, 16'd17837, 16'd11548, 16'd48978, 16'd4427, 16'd10692, 16'd6635, 16'd54799, 16'd59742, 16'd61579, 16'd30894, 16'd63347, 16'd47427, 16'd2400, 16'd22751, 16'd59439, 16'd38800, 16'd61454, 16'd13470, 16'd39202, 16'd58810, 16'd31967, 16'd36384});
	test_expansion(128'hb43994a1dc029064580bad143308c09a, {16'd47000, 16'd7311, 16'd46900, 16'd17050, 16'd21221, 16'd47479, 16'd44200, 16'd56455, 16'd21642, 16'd15071, 16'd32656, 16'd1091, 16'd12406, 16'd30844, 16'd56167, 16'd23371, 16'd44031, 16'd22725, 16'd18597, 16'd38809, 16'd33320, 16'd59706, 16'd25737, 16'd116, 16'd55364, 16'd59191});
	test_expansion(128'h63faebcd07346d7786c0cb5e0602e1d1, {16'd32139, 16'd10003, 16'd61022, 16'd13931, 16'd27369, 16'd60028, 16'd51710, 16'd3050, 16'd28053, 16'd10679, 16'd25715, 16'd64274, 16'd29332, 16'd63217, 16'd13252, 16'd63172, 16'd24099, 16'd24074, 16'd51753, 16'd11933, 16'd9885, 16'd32250, 16'd60912, 16'd63517, 16'd20220, 16'd24063});
	test_expansion(128'hecf8f7be9e71b15c16b3d0ec8afb6a0d, {16'd17294, 16'd25765, 16'd34365, 16'd47024, 16'd5899, 16'd16082, 16'd53625, 16'd26154, 16'd59927, 16'd4467, 16'd25502, 16'd21625, 16'd31723, 16'd65467, 16'd25068, 16'd56587, 16'd50980, 16'd31156, 16'd28156, 16'd25342, 16'd46245, 16'd54395, 16'd4782, 16'd52598, 16'd24230, 16'd28636});
	test_expansion(128'hfc00336772b3b1fd87f2cca3b10fe67e, {16'd5859, 16'd33128, 16'd38788, 16'd4880, 16'd41937, 16'd34920, 16'd14816, 16'd33712, 16'd50951, 16'd28917, 16'd33110, 16'd39126, 16'd20607, 16'd46132, 16'd43690, 16'd43744, 16'd17864, 16'd32575, 16'd53720, 16'd52470, 16'd58572, 16'd58989, 16'd55425, 16'd11948, 16'd61171, 16'd33839});
	test_expansion(128'h79c424a66b89ad1fcb74c3fe2b82bb8a, {16'd10181, 16'd34777, 16'd8915, 16'd27316, 16'd16062, 16'd56922, 16'd64599, 16'd295, 16'd52442, 16'd1850, 16'd12106, 16'd25139, 16'd64442, 16'd52455, 16'd20423, 16'd51525, 16'd48360, 16'd39897, 16'd65043, 16'd14261, 16'd62201, 16'd56862, 16'd56593, 16'd16030, 16'd34842, 16'd3283});
	test_expansion(128'h035d015f6037648ad6eba3b9e3cea72e, {16'd37708, 16'd48214, 16'd4438, 16'd32385, 16'd18071, 16'd20359, 16'd26194, 16'd46913, 16'd18190, 16'd41585, 16'd63113, 16'd48348, 16'd57133, 16'd2751, 16'd32535, 16'd58333, 16'd22437, 16'd26868, 16'd26651, 16'd36011, 16'd61963, 16'd62550, 16'd53656, 16'd23626, 16'd58773, 16'd58161});
	test_expansion(128'h802d981a060c8070ea05ecfd02fc4adc, {16'd38669, 16'd35063, 16'd10016, 16'd49739, 16'd62485, 16'd30925, 16'd64931, 16'd25562, 16'd27344, 16'd53922, 16'd57224, 16'd33460, 16'd11724, 16'd19808, 16'd8220, 16'd45937, 16'd36812, 16'd64838, 16'd14296, 16'd2226, 16'd24539, 16'd18834, 16'd32135, 16'd27911, 16'd11290, 16'd60924});
	test_expansion(128'h4e6e3d0ad58e34491a6d10896a252387, {16'd16078, 16'd36030, 16'd64563, 16'd17511, 16'd22351, 16'd34967, 16'd32891, 16'd28943, 16'd39259, 16'd27458, 16'd58235, 16'd61663, 16'd29274, 16'd34067, 16'd38632, 16'd42280, 16'd59554, 16'd11041, 16'd53468, 16'd19191, 16'd7849, 16'd11559, 16'd63370, 16'd54296, 16'd47163, 16'd58898});
	test_expansion(128'h7760e77d0d1507c8f3d332bd101992d7, {16'd62789, 16'd39444, 16'd35089, 16'd29491, 16'd5960, 16'd35862, 16'd60247, 16'd49903, 16'd57203, 16'd34327, 16'd4459, 16'd12659, 16'd26402, 16'd64931, 16'd12550, 16'd6880, 16'd6329, 16'd3184, 16'd41117, 16'd46026, 16'd22725, 16'd44441, 16'd54313, 16'd54911, 16'd33826, 16'd17808});
	test_expansion(128'hb6250b8e55049c2b46d9f807d8f23097, {16'd27156, 16'd54646, 16'd53180, 16'd48631, 16'd15767, 16'd30268, 16'd5848, 16'd5247, 16'd1470, 16'd14887, 16'd42533, 16'd62521, 16'd42635, 16'd61165, 16'd6082, 16'd39769, 16'd34021, 16'd23179, 16'd15072, 16'd47239, 16'd42958, 16'd20640, 16'd24765, 16'd24355, 16'd41511, 16'd46074});
	test_expansion(128'h679f36a85a3d4c3b6f351278908d148f, {16'd24160, 16'd62318, 16'd56587, 16'd17285, 16'd7645, 16'd54227, 16'd10820, 16'd45279, 16'd44720, 16'd13876, 16'd43436, 16'd50489, 16'd5351, 16'd28052, 16'd50842, 16'd26440, 16'd33234, 16'd42392, 16'd38838, 16'd36659, 16'd60384, 16'd60690, 16'd35938, 16'd14770, 16'd40869, 16'd8104});
	test_expansion(128'h277054d7f6e6e3b77ae0e75321066a20, {16'd37124, 16'd6313, 16'd24278, 16'd30847, 16'd64734, 16'd5952, 16'd49043, 16'd50375, 16'd10451, 16'd11876, 16'd4790, 16'd45128, 16'd13075, 16'd9285, 16'd6457, 16'd17625, 16'd52920, 16'd6672, 16'd43420, 16'd32394, 16'd29186, 16'd2003, 16'd60100, 16'd55839, 16'd46037, 16'd56536});
	test_expansion(128'h5d48c996f4d8cb2e5cebab2b3236cc1d, {16'd64894, 16'd32347, 16'd43648, 16'd14528, 16'd38858, 16'd42413, 16'd45933, 16'd8251, 16'd62317, 16'd407, 16'd55862, 16'd5303, 16'd56575, 16'd20087, 16'd56200, 16'd19599, 16'd45137, 16'd50584, 16'd22052, 16'd21329, 16'd53694, 16'd19806, 16'd51510, 16'd43944, 16'd10876, 16'd16542});
	test_expansion(128'hf394b4a1d2e0c716c05c302028026be6, {16'd32757, 16'd26488, 16'd41768, 16'd29652, 16'd26482, 16'd17476, 16'd29324, 16'd45378, 16'd21166, 16'd45591, 16'd6309, 16'd45586, 16'd45805, 16'd22672, 16'd12213, 16'd61547, 16'd37622, 16'd40960, 16'd62726, 16'd27343, 16'd32164, 16'd63197, 16'd9743, 16'd61032, 16'd53624, 16'd9357});
	test_expansion(128'h718bbc3354651c0a0f12c293997643ad, {16'd58542, 16'd52878, 16'd32865, 16'd19895, 16'd40666, 16'd60492, 16'd33880, 16'd48355, 16'd45057, 16'd19624, 16'd53089, 16'd10049, 16'd12028, 16'd24882, 16'd33786, 16'd32496, 16'd57830, 16'd28192, 16'd57730, 16'd4816, 16'd35302, 16'd5654, 16'd55617, 16'd13402, 16'd6221, 16'd48536});
	test_expansion(128'h79b2a8812e190a8c83fc590e7ab742e0, {16'd36083, 16'd27777, 16'd30663, 16'd27268, 16'd62591, 16'd12388, 16'd51588, 16'd12729, 16'd41155, 16'd24629, 16'd1352, 16'd23499, 16'd33673, 16'd46400, 16'd44769, 16'd41031, 16'd56770, 16'd8298, 16'd40629, 16'd14929, 16'd57790, 16'd50849, 16'd51553, 16'd5051, 16'd39041, 16'd59990});
	test_expansion(128'h4b09921c57f6e37588312c3cba3f6dfe, {16'd19412, 16'd51474, 16'd52193, 16'd38170, 16'd33807, 16'd6841, 16'd63354, 16'd5435, 16'd47818, 16'd56066, 16'd53792, 16'd55639, 16'd18660, 16'd2046, 16'd22094, 16'd5036, 16'd44563, 16'd47375, 16'd26743, 16'd2432, 16'd22809, 16'd61796, 16'd25948, 16'd39832, 16'd42106, 16'd35326});
	test_expansion(128'ha17a0de91578d88883e17cb83cdbc132, {16'd20153, 16'd27304, 16'd14001, 16'd32902, 16'd32303, 16'd27361, 16'd3890, 16'd46642, 16'd62716, 16'd28558, 16'd24828, 16'd54652, 16'd36711, 16'd14163, 16'd64157, 16'd43461, 16'd26320, 16'd19565, 16'd34305, 16'd42515, 16'd30228, 16'd57055, 16'd10994, 16'd15278, 16'd35186, 16'd57725});
	test_expansion(128'hc2b5385bbee637ecd2ee85e5e4280775, {16'd63683, 16'd12407, 16'd11409, 16'd18450, 16'd36140, 16'd15574, 16'd53108, 16'd54624, 16'd44540, 16'd6858, 16'd20578, 16'd58613, 16'd57521, 16'd37867, 16'd30258, 16'd48184, 16'd24102, 16'd37973, 16'd30834, 16'd36876, 16'd40760, 16'd13227, 16'd4078, 16'd28655, 16'd62002, 16'd40282});
	test_expansion(128'hefc4eefbd65b18b10ad86af130d16a6f, {16'd23698, 16'd12419, 16'd53988, 16'd53698, 16'd41481, 16'd8701, 16'd38682, 16'd1678, 16'd47004, 16'd45567, 16'd42844, 16'd64308, 16'd56043, 16'd11532, 16'd5441, 16'd11568, 16'd1586, 16'd9866, 16'd5957, 16'd18475, 16'd3929, 16'd6489, 16'd52945, 16'd44230, 16'd31820, 16'd53462});
	test_expansion(128'h1c27b767ac12fda8ff548cfb44b4ff0a, {16'd21102, 16'd43150, 16'd8743, 16'd62236, 16'd61032, 16'd7255, 16'd24736, 16'd26544, 16'd3198, 16'd2539, 16'd46592, 16'd53100, 16'd6576, 16'd30934, 16'd24270, 16'd41353, 16'd65417, 16'd42444, 16'd20222, 16'd25454, 16'd20706, 16'd4890, 16'd54408, 16'd34668, 16'd35616, 16'd45365});
	test_expansion(128'h532177369aded68eae5fe3b7a27b8a16, {16'd28386, 16'd41267, 16'd35035, 16'd42760, 16'd10583, 16'd50313, 16'd8404, 16'd27791, 16'd30533, 16'd27507, 16'd63285, 16'd36724, 16'd40373, 16'd20086, 16'd43164, 16'd27876, 16'd19982, 16'd29727, 16'd47489, 16'd35973, 16'd27457, 16'd52864, 16'd23659, 16'd43761, 16'd12486, 16'd35636});
	test_expansion(128'haadecc8c98ecd94c9c31105ad246e304, {16'd4991, 16'd56832, 16'd55156, 16'd41305, 16'd28632, 16'd8854, 16'd720, 16'd43455, 16'd11639, 16'd22203, 16'd27196, 16'd59017, 16'd31545, 16'd28997, 16'd62906, 16'd5698, 16'd57918, 16'd2303, 16'd5545, 16'd31004, 16'd64290, 16'd51792, 16'd14901, 16'd56823, 16'd5869, 16'd2878});
	test_expansion(128'h7048277edd5d1a5f2bc150c819a537d0, {16'd64915, 16'd62026, 16'd52300, 16'd34995, 16'd8218, 16'd55580, 16'd34587, 16'd23139, 16'd58706, 16'd36682, 16'd35043, 16'd38881, 16'd54337, 16'd59872, 16'd32314, 16'd44849, 16'd29313, 16'd36907, 16'd48360, 16'd29625, 16'd4886, 16'd7287, 16'd47408, 16'd28005, 16'd16255, 16'd23560});
	test_expansion(128'h412305919a89508cbc6ee4f604edfdbe, {16'd6350, 16'd56556, 16'd34283, 16'd58968, 16'd51179, 16'd46374, 16'd41133, 16'd23783, 16'd55848, 16'd50715, 16'd3694, 16'd18141, 16'd23962, 16'd25117, 16'd65319, 16'd48225, 16'd29348, 16'd10535, 16'd39313, 16'd1821, 16'd32018, 16'd33498, 16'd48024, 16'd51405, 16'd25743, 16'd12373});
	test_expansion(128'hc8c3d8df324e9a6b2504038a5595300b, {16'd21828, 16'd14357, 16'd41192, 16'd46089, 16'd65007, 16'd55352, 16'd47139, 16'd58631, 16'd38410, 16'd39533, 16'd1609, 16'd61258, 16'd4079, 16'd54233, 16'd21617, 16'd41761, 16'd23336, 16'd60939, 16'd24463, 16'd54528, 16'd58263, 16'd17880, 16'd15167, 16'd46327, 16'd14520, 16'd19332});
	test_expansion(128'h9dd21043986f71a9d0f19c7c36b822e1, {16'd51935, 16'd17588, 16'd1130, 16'd63349, 16'd17579, 16'd29486, 16'd48443, 16'd58443, 16'd35254, 16'd24048, 16'd18143, 16'd6973, 16'd52054, 16'd43230, 16'd9647, 16'd21108, 16'd50957, 16'd38314, 16'd13199, 16'd62414, 16'd34372, 16'd62282, 16'd60155, 16'd19929, 16'd48790, 16'd12247});
	test_expansion(128'h4f354a6853773ad1fcd6118606e6738a, {16'd29717, 16'd13720, 16'd25521, 16'd59106, 16'd38744, 16'd41081, 16'd2939, 16'd15732, 16'd13364, 16'd50156, 16'd52832, 16'd50186, 16'd62861, 16'd5316, 16'd46883, 16'd774, 16'd22054, 16'd27614, 16'd2144, 16'd22733, 16'd54104, 16'd32312, 16'd12855, 16'd40137, 16'd40529, 16'd42982});
	test_expansion(128'h649045ec2bbbba8f27809c8c6045624e, {16'd48128, 16'd46258, 16'd65427, 16'd20665, 16'd49320, 16'd51833, 16'd63676, 16'd45430, 16'd57883, 16'd44156, 16'd25123, 16'd61422, 16'd26837, 16'd30944, 16'd40473, 16'd24177, 16'd21145, 16'd41299, 16'd19659, 16'd56648, 16'd29505, 16'd60650, 16'd6817, 16'd32927, 16'd59075, 16'd49760});
	test_expansion(128'h1328bb4a7d9faba457a2d23593cd57ad, {16'd12547, 16'd30171, 16'd30680, 16'd46299, 16'd14004, 16'd21373, 16'd50838, 16'd15521, 16'd2448, 16'd25236, 16'd14134, 16'd41778, 16'd47145, 16'd39564, 16'd6636, 16'd64184, 16'd55501, 16'd59987, 16'd40780, 16'd44302, 16'd33413, 16'd43956, 16'd39401, 16'd58048, 16'd43952, 16'd18838});
	test_expansion(128'hbec399d6775b920d3108ebb669e19d18, {16'd24113, 16'd1531, 16'd4346, 16'd14874, 16'd3992, 16'd36671, 16'd51188, 16'd5612, 16'd20085, 16'd46953, 16'd13881, 16'd41224, 16'd56871, 16'd33487, 16'd17276, 16'd47516, 16'd16439, 16'd27435, 16'd62573, 16'd46531, 16'd63997, 16'd31513, 16'd18248, 16'd28815, 16'd59488, 16'd34221});
	test_expansion(128'h72775394396743628f76ed989fd4ba90, {16'd59432, 16'd52280, 16'd11895, 16'd15835, 16'd19725, 16'd46151, 16'd46020, 16'd31818, 16'd5386, 16'd1194, 16'd23795, 16'd5135, 16'd60541, 16'd22880, 16'd55428, 16'd11622, 16'd49700, 16'd21633, 16'd44414, 16'd10844, 16'd4562, 16'd25975, 16'd59760, 16'd49802, 16'd57309, 16'd32901});
	test_expansion(128'h559c3de3607d0f23d58db3371d5abd94, {16'd60739, 16'd21659, 16'd9326, 16'd443, 16'd56802, 16'd32418, 16'd3945, 16'd19905, 16'd56020, 16'd33065, 16'd55722, 16'd9702, 16'd41253, 16'd10400, 16'd1452, 16'd6236, 16'd62893, 16'd56254, 16'd17212, 16'd28581, 16'd13313, 16'd57736, 16'd10965, 16'd57774, 16'd43491, 16'd54685});
	test_expansion(128'h03df78dd721e457a25f28b54721a84e5, {16'd31657, 16'd40098, 16'd25468, 16'd40064, 16'd5982, 16'd13471, 16'd17560, 16'd44987, 16'd10005, 16'd44650, 16'd29198, 16'd20679, 16'd5408, 16'd39178, 16'd46201, 16'd63856, 16'd28372, 16'd16240, 16'd10316, 16'd49280, 16'd49633, 16'd20831, 16'd31281, 16'd17210, 16'd37044, 16'd37554});
	test_expansion(128'h1b6a5c84fd3a36e77e6e9cfcb3c5ca75, {16'd36440, 16'd59833, 16'd2161, 16'd28693, 16'd50595, 16'd46083, 16'd26130, 16'd8596, 16'd28027, 16'd39739, 16'd49263, 16'd11, 16'd26878, 16'd6368, 16'd18467, 16'd43844, 16'd13595, 16'd49101, 16'd62758, 16'd46559, 16'd22155, 16'd18780, 16'd18677, 16'd36491, 16'd32475, 16'd54630});
	test_expansion(128'h1b36a52021bccd05a527990ca5141127, {16'd19160, 16'd54043, 16'd12483, 16'd8779, 16'd17018, 16'd11683, 16'd58272, 16'd38435, 16'd56116, 16'd43750, 16'd1399, 16'd55774, 16'd54750, 16'd26707, 16'd63943, 16'd34867, 16'd44419, 16'd45426, 16'd2464, 16'd13344, 16'd28862, 16'd14184, 16'd52433, 16'd61023, 16'd17068, 16'd12797});
	test_expansion(128'hcbec0ceb6bb2102a5f0234997ee0d9dc, {16'd57355, 16'd11639, 16'd44693, 16'd26051, 16'd29113, 16'd21771, 16'd45468, 16'd58193, 16'd45348, 16'd47963, 16'd4222, 16'd35717, 16'd63949, 16'd43811, 16'd22300, 16'd41673, 16'd61250, 16'd32220, 16'd43337, 16'd49573, 16'd12010, 16'd10756, 16'd20791, 16'd60900, 16'd971, 16'd14818});
	test_expansion(128'haac19a25616c07b3fe3dfb8ac637cebd, {16'd59515, 16'd683, 16'd39001, 16'd9245, 16'd12561, 16'd49737, 16'd39609, 16'd42523, 16'd7506, 16'd23050, 16'd65136, 16'd26383, 16'd61778, 16'd33905, 16'd64695, 16'd19466, 16'd2332, 16'd46170, 16'd1201, 16'd25919, 16'd8135, 16'd22017, 16'd25971, 16'd26070, 16'd65404, 16'd12692});
	test_expansion(128'hb94c9e44001e158a3a65e21c0f8a6a80, {16'd50382, 16'd20056, 16'd44573, 16'd23993, 16'd54629, 16'd2848, 16'd20375, 16'd27638, 16'd61256, 16'd21205, 16'd57080, 16'd41942, 16'd36537, 16'd38337, 16'd12564, 16'd12210, 16'd59998, 16'd13083, 16'd52393, 16'd57516, 16'd36661, 16'd46652, 16'd45941, 16'd1634, 16'd198, 16'd29675});
	test_expansion(128'h10d3a9f91c713a21a789c2c1c312857e, {16'd1897, 16'd35314, 16'd61829, 16'd18427, 16'd10027, 16'd26328, 16'd26693, 16'd14525, 16'd1564, 16'd57575, 16'd60122, 16'd63217, 16'd44548, 16'd10277, 16'd60137, 16'd63889, 16'd35524, 16'd6416, 16'd47156, 16'd34979, 16'd19995, 16'd237, 16'd51250, 16'd36404, 16'd46774, 16'd33526});
	test_expansion(128'hca129f932b63ed263434465c605b31f7, {16'd3842, 16'd13197, 16'd37876, 16'd6893, 16'd24651, 16'd19241, 16'd60883, 16'd30914, 16'd21054, 16'd2968, 16'd45335, 16'd61557, 16'd56435, 16'd45770, 16'd50449, 16'd47341, 16'd17339, 16'd22078, 16'd15776, 16'd34006, 16'd49176, 16'd8417, 16'd58949, 16'd31216, 16'd61749, 16'd38698});
	test_expansion(128'h0e859f472adf89f649c9901af3255ff2, {16'd12744, 16'd19277, 16'd59335, 16'd57270, 16'd239, 16'd16882, 16'd14740, 16'd32976, 16'd42349, 16'd58272, 16'd15081, 16'd22233, 16'd43282, 16'd6878, 16'd20204, 16'd16348, 16'd14822, 16'd61965, 16'd13911, 16'd15326, 16'd7302, 16'd58802, 16'd58066, 16'd25846, 16'd48849, 16'd39771});
	test_expansion(128'hcde7a95e802f0e5f414b409152bb6f75, {16'd38660, 16'd33867, 16'd8645, 16'd54421, 16'd9839, 16'd16301, 16'd266, 16'd14138, 16'd59485, 16'd26822, 16'd197, 16'd25001, 16'd55913, 16'd32761, 16'd10359, 16'd37034, 16'd7359, 16'd55362, 16'd7485, 16'd3298, 16'd53752, 16'd65349, 16'd24540, 16'd51191, 16'd64396, 16'd22948});
	test_expansion(128'h7942e687283cfabe0ef7b89fd6559328, {16'd63603, 16'd44452, 16'd31133, 16'd42495, 16'd11296, 16'd32856, 16'd16698, 16'd35701, 16'd47789, 16'd23246, 16'd58391, 16'd32971, 16'd1014, 16'd49673, 16'd12499, 16'd7190, 16'd61628, 16'd28030, 16'd29318, 16'd59540, 16'd59234, 16'd40897, 16'd14933, 16'd29331, 16'd36231, 16'd13715});
	test_expansion(128'hb2b6ab7b1cbf18f892e13b1899986552, {16'd50490, 16'd22425, 16'd25530, 16'd38676, 16'd65381, 16'd60487, 16'd2843, 16'd11572, 16'd33962, 16'd19481, 16'd16552, 16'd52007, 16'd59993, 16'd10557, 16'd28017, 16'd15951, 16'd55923, 16'd23414, 16'd29855, 16'd50356, 16'd22060, 16'd6034, 16'd141, 16'd57462, 16'd49794, 16'd53873});
	test_expansion(128'ha5e5ee39f1687db558413a8319b98657, {16'd46171, 16'd63027, 16'd55288, 16'd12890, 16'd2658, 16'd52005, 16'd44634, 16'd418, 16'd48771, 16'd26192, 16'd23106, 16'd23935, 16'd27930, 16'd19583, 16'd18678, 16'd25961, 16'd3460, 16'd14875, 16'd41182, 16'd14386, 16'd53965, 16'd37939, 16'd43184, 16'd59068, 16'd52690, 16'd2433});
	test_expansion(128'h162458b8fbc2378f9f8c1a1168f241fb, {16'd38786, 16'd34039, 16'd7621, 16'd48189, 16'd12557, 16'd55505, 16'd13336, 16'd25708, 16'd15869, 16'd38023, 16'd43791, 16'd15413, 16'd45302, 16'd48705, 16'd31400, 16'd56828, 16'd24456, 16'd28487, 16'd22653, 16'd14012, 16'd47422, 16'd45371, 16'd38573, 16'd50249, 16'd10186, 16'd20383});
	test_expansion(128'hf39f1fb6b6130ee177ce7195e54a5d59, {16'd8282, 16'd38835, 16'd56242, 16'd30807, 16'd20703, 16'd20054, 16'd53387, 16'd22203, 16'd47263, 16'd8261, 16'd26610, 16'd23492, 16'd48818, 16'd52635, 16'd55362, 16'd35568, 16'd12803, 16'd24146, 16'd30151, 16'd28332, 16'd9121, 16'd31420, 16'd11197, 16'd55473, 16'd35126, 16'd24526});
	test_expansion(128'h6835744767627c39c1eee33ef6affc72, {16'd28788, 16'd10925, 16'd24449, 16'd38257, 16'd15298, 16'd61223, 16'd26745, 16'd26246, 16'd38553, 16'd36402, 16'd11928, 16'd47462, 16'd10659, 16'd49862, 16'd55973, 16'd29076, 16'd58791, 16'd26132, 16'd38650, 16'd39857, 16'd4330, 16'd37798, 16'd21557, 16'd6711, 16'd29089, 16'd58668});
	test_expansion(128'hebf3c725d9e6c4c7d6031ddcc0b48ffe, {16'd23530, 16'd45590, 16'd15993, 16'd57364, 16'd9035, 16'd64307, 16'd23039, 16'd22860, 16'd30967, 16'd51689, 16'd47958, 16'd32325, 16'd35805, 16'd41315, 16'd30516, 16'd59990, 16'd45018, 16'd58774, 16'd21766, 16'd57413, 16'd47979, 16'd37705, 16'd5367, 16'd14086, 16'd1296, 16'd29084});
	test_expansion(128'had9c8b07b776bfbbee4b37ad800f832a, {16'd57600, 16'd65383, 16'd77, 16'd32864, 16'd54720, 16'd8539, 16'd4077, 16'd4679, 16'd353, 16'd11728, 16'd54293, 16'd17354, 16'd17649, 16'd39402, 16'd24143, 16'd32692, 16'd42832, 16'd46098, 16'd62480, 16'd5321, 16'd49441, 16'd4725, 16'd45975, 16'd21080, 16'd25223, 16'd16909});
	test_expansion(128'hce4f17f94e3e89cf3214e86b33db4e93, {16'd35712, 16'd8689, 16'd2633, 16'd15560, 16'd57921, 16'd48952, 16'd18112, 16'd46463, 16'd60789, 16'd32675, 16'd55239, 16'd53563, 16'd14255, 16'd5824, 16'd34590, 16'd59840, 16'd25935, 16'd25188, 16'd10489, 16'd23890, 16'd27069, 16'd51619, 16'd46600, 16'd39712, 16'd8553, 16'd49576});
	test_expansion(128'h126835db81224c2184f8acf600937ff0, {16'd64267, 16'd13664, 16'd54153, 16'd28787, 16'd36377, 16'd45845, 16'd11134, 16'd51371, 16'd57818, 16'd39538, 16'd16657, 16'd9419, 16'd46854, 16'd27912, 16'd54377, 16'd39820, 16'd3185, 16'd12091, 16'd33433, 16'd41475, 16'd41498, 16'd50322, 16'd13714, 16'd32643, 16'd36983, 16'd22416});
	test_expansion(128'he40c3db097fdc8d5d13a93940f9ea5fe, {16'd11519, 16'd29474, 16'd2094, 16'd46420, 16'd24240, 16'd22738, 16'd19908, 16'd28994, 16'd29519, 16'd7238, 16'd61101, 16'd35101, 16'd13080, 16'd12677, 16'd160, 16'd23519, 16'd32223, 16'd8334, 16'd54895, 16'd59151, 16'd35477, 16'd47478, 16'd16665, 16'd56022, 16'd56733, 16'd47174});
	test_expansion(128'h4d0d41cef4e9ad8d16412fb27188050f, {16'd45818, 16'd51369, 16'd22648, 16'd21420, 16'd14129, 16'd52030, 16'd16502, 16'd11664, 16'd35588, 16'd32930, 16'd31987, 16'd52727, 16'd9577, 16'd31810, 16'd19823, 16'd52087, 16'd47198, 16'd22001, 16'd23264, 16'd25107, 16'd35720, 16'd6237, 16'd47046, 16'd15818, 16'd10267, 16'd36524});
	test_expansion(128'h0a0eaacd31dd5d2d615e3e53a9d9ef87, {16'd63364, 16'd53870, 16'd5864, 16'd51575, 16'd29432, 16'd52830, 16'd52446, 16'd41590, 16'd24691, 16'd14475, 16'd16685, 16'd15276, 16'd65334, 16'd6020, 16'd39735, 16'd2698, 16'd30190, 16'd65203, 16'd42661, 16'd22650, 16'd50925, 16'd8456, 16'd45294, 16'd54762, 16'd36936, 16'd61705});
	test_expansion(128'h82467d823288a6e352459bbad9d3cacd, {16'd13780, 16'd63942, 16'd46767, 16'd64360, 16'd54368, 16'd25150, 16'd48310, 16'd58989, 16'd59213, 16'd62634, 16'd21717, 16'd47828, 16'd14528, 16'd51042, 16'd20396, 16'd64319, 16'd40203, 16'd17670, 16'd5842, 16'd54255, 16'd24128, 16'd45571, 16'd33065, 16'd34875, 16'd53858, 16'd54278});
	test_expansion(128'h16907b8401d960ce102dc0279ddeb2bf, {16'd15952, 16'd8132, 16'd19568, 16'd7131, 16'd20303, 16'd55111, 16'd4385, 16'd43477, 16'd19375, 16'd27481, 16'd58347, 16'd192, 16'd13881, 16'd37593, 16'd55296, 16'd27756, 16'd20757, 16'd21930, 16'd19810, 16'd52250, 16'd13318, 16'd63268, 16'd29865, 16'd56638, 16'd4496, 16'd57134});
	test_expansion(128'h8479d23b8704940db7ebaf247f2a708c, {16'd707, 16'd18745, 16'd11366, 16'd25169, 16'd11590, 16'd53020, 16'd40107, 16'd14705, 16'd65120, 16'd9132, 16'd65427, 16'd61939, 16'd49420, 16'd7732, 16'd10269, 16'd53374, 16'd18416, 16'd62210, 16'd56534, 16'd58072, 16'd31439, 16'd37759, 16'd45873, 16'd59880, 16'd36786, 16'd18923});
	test_expansion(128'hc98f644fd510f8912bf278e6ae23c069, {16'd40959, 16'd16623, 16'd282, 16'd31958, 16'd36177, 16'd22167, 16'd38320, 16'd41367, 16'd44620, 16'd22692, 16'd9295, 16'd208, 16'd40666, 16'd20773, 16'd2242, 16'd11412, 16'd44992, 16'd39931, 16'd64896, 16'd41340, 16'd27895, 16'd6233, 16'd5593, 16'd55826, 16'd6537, 16'd31679});
	test_expansion(128'h71003c9edb510280d1d14fd22edf4528, {16'd30131, 16'd34326, 16'd26085, 16'd60472, 16'd11114, 16'd38778, 16'd21175, 16'd41092, 16'd6931, 16'd26945, 16'd45470, 16'd30025, 16'd6788, 16'd41077, 16'd54137, 16'd6813, 16'd6700, 16'd32098, 16'd14846, 16'd59883, 16'd7703, 16'd46885, 16'd15831, 16'd46287, 16'd50706, 16'd40023});
	test_expansion(128'h9e5e10f78ce8dce73bc62265d531878e, {16'd5313, 16'd4365, 16'd16226, 16'd1467, 16'd50856, 16'd33837, 16'd38478, 16'd31238, 16'd11499, 16'd44669, 16'd51342, 16'd50447, 16'd47253, 16'd8295, 16'd56159, 16'd45124, 16'd60946, 16'd52851, 16'd38236, 16'd20470, 16'd1427, 16'd16849, 16'd46559, 16'd53341, 16'd6158, 16'd30298});
	test_expansion(128'h74989933615f9825bb61bc5cb4c43007, {16'd3004, 16'd36240, 16'd59236, 16'd42740, 16'd6054, 16'd61694, 16'd14677, 16'd9427, 16'd42586, 16'd22118, 16'd39325, 16'd27593, 16'd18288, 16'd31953, 16'd47534, 16'd60501, 16'd60162, 16'd28785, 16'd29906, 16'd10660, 16'd39270, 16'd61733, 16'd58319, 16'd30994, 16'd43303, 16'd38474});
	test_expansion(128'h5edd725e60fa66a2488a5c0820c64434, {16'd25978, 16'd14677, 16'd31394, 16'd22705, 16'd22966, 16'd719, 16'd14221, 16'd6262, 16'd24866, 16'd40527, 16'd52366, 16'd39813, 16'd32147, 16'd1321, 16'd35823, 16'd39096, 16'd49809, 16'd63342, 16'd24164, 16'd56733, 16'd61362, 16'd49243, 16'd23457, 16'd19965, 16'd19469, 16'd52369});
	test_expansion(128'ha8e111961c5105354bf8a9f0c90aa2a4, {16'd18105, 16'd47432, 16'd35000, 16'd18399, 16'd34563, 16'd51550, 16'd62302, 16'd27203, 16'd6800, 16'd64495, 16'd32481, 16'd33486, 16'd60830, 16'd31930, 16'd6554, 16'd43519, 16'd4181, 16'd15355, 16'd60194, 16'd27854, 16'd1722, 16'd21156, 16'd1905, 16'd31851, 16'd5388, 16'd43122});
	test_expansion(128'hfb7d1d513a0da59936af9b0824eb0e52, {16'd38316, 16'd6506, 16'd43778, 16'd17152, 16'd20313, 16'd30884, 16'd3163, 16'd22523, 16'd39315, 16'd29948, 16'd29804, 16'd60451, 16'd52485, 16'd50341, 16'd27397, 16'd55799, 16'd45770, 16'd45841, 16'd43839, 16'd10897, 16'd50482, 16'd61682, 16'd58702, 16'd6755, 16'd10775, 16'd48816});
	test_expansion(128'hd09d42230d57e40b244eb6c31296000a, {16'd42065, 16'd59777, 16'd34431, 16'd51106, 16'd24276, 16'd9433, 16'd19755, 16'd19866, 16'd15976, 16'd62005, 16'd23033, 16'd52022, 16'd14740, 16'd60953, 16'd22863, 16'd3657, 16'd14191, 16'd62916, 16'd63816, 16'd39980, 16'd352, 16'd7774, 16'd3327, 16'd52519, 16'd6728, 16'd55619});
	test_expansion(128'hc9320d4ac07fb78d2abed178d325fe44, {16'd15966, 16'd11372, 16'd39467, 16'd43629, 16'd42907, 16'd64217, 16'd57280, 16'd33189, 16'd36743, 16'd20566, 16'd2838, 16'd58589, 16'd6028, 16'd53451, 16'd8214, 16'd26889, 16'd43912, 16'd44106, 16'd58504, 16'd33566, 16'd15185, 16'd31851, 16'd43127, 16'd35087, 16'd60094, 16'd6867});
	test_expansion(128'h80cc760376cd67056e974500ac9c91ef, {16'd5655, 16'd30419, 16'd13719, 16'd52545, 16'd50872, 16'd1714, 16'd21175, 16'd34582, 16'd56416, 16'd45299, 16'd9005, 16'd14962, 16'd18323, 16'd24768, 16'd44017, 16'd59705, 16'd10365, 16'd9023, 16'd17936, 16'd2929, 16'd52665, 16'd51001, 16'd15037, 16'd1369, 16'd34207, 16'd24547});
	test_expansion(128'hf8e4221469a8782ab10f3b5589b71575, {16'd42753, 16'd56463, 16'd35272, 16'd65213, 16'd25535, 16'd8602, 16'd47099, 16'd14120, 16'd12319, 16'd19320, 16'd30961, 16'd48402, 16'd12576, 16'd49973, 16'd16397, 16'd61453, 16'd48993, 16'd27314, 16'd30030, 16'd59172, 16'd9520, 16'd59387, 16'd4663, 16'd9584, 16'd47884, 16'd41206});
	test_expansion(128'h9b2cc2994e51470e758f48a1137e2827, {16'd41759, 16'd31486, 16'd53420, 16'd22933, 16'd30859, 16'd33563, 16'd41109, 16'd11808, 16'd49193, 16'd20715, 16'd52353, 16'd65210, 16'd13789, 16'd54677, 16'd3297, 16'd9665, 16'd60258, 16'd37391, 16'd11493, 16'd36414, 16'd57266, 16'd62326, 16'd20482, 16'd7822, 16'd11440, 16'd36412});
	test_expansion(128'hfb0d140cb4070620e8618c7ead79d45b, {16'd1505, 16'd33853, 16'd56076, 16'd43540, 16'd52379, 16'd40085, 16'd17895, 16'd25048, 16'd46339, 16'd21246, 16'd24399, 16'd34734, 16'd25606, 16'd47539, 16'd58147, 16'd50258, 16'd57227, 16'd50028, 16'd23128, 16'd64554, 16'd36057, 16'd8889, 16'd16599, 16'd39727, 16'd58457, 16'd33304});
	test_expansion(128'h0158b06c06b283db0071df9506041cf8, {16'd4327, 16'd35212, 16'd59221, 16'd35312, 16'd38760, 16'd62367, 16'd5618, 16'd46611, 16'd51350, 16'd22885, 16'd27345, 16'd13838, 16'd36844, 16'd20909, 16'd23937, 16'd31456, 16'd19905, 16'd40174, 16'd2636, 16'd24093, 16'd54236, 16'd2924, 16'd15694, 16'd48297, 16'd41260, 16'd3685});
	test_expansion(128'h4693a99c9cf8078f71e0517c8074cfe7, {16'd6094, 16'd56285, 16'd36481, 16'd31959, 16'd838, 16'd35136, 16'd15215, 16'd3933, 16'd64469, 16'd41180, 16'd3519, 16'd34744, 16'd19064, 16'd42118, 16'd48129, 16'd33781, 16'd26882, 16'd25189, 16'd20313, 16'd43166, 16'd31625, 16'd26673, 16'd41102, 16'd65478, 16'd50507, 16'd47374});
	test_expansion(128'h8f30540c0f4f07a8dea48d688a328876, {16'd40458, 16'd1136, 16'd22428, 16'd38166, 16'd5384, 16'd53965, 16'd33354, 16'd42416, 16'd46143, 16'd57364, 16'd45836, 16'd31050, 16'd59258, 16'd55515, 16'd27629, 16'd25095, 16'd54807, 16'd32603, 16'd54382, 16'd22169, 16'd55630, 16'd38312, 16'd49309, 16'd52220, 16'd29349, 16'd23261});
	test_expansion(128'h3a2a7c264528576043840149d0b66c5a, {16'd22376, 16'd27023, 16'd43112, 16'd1996, 16'd7796, 16'd1321, 16'd53828, 16'd26943, 16'd21473, 16'd62035, 16'd34090, 16'd64137, 16'd49952, 16'd32887, 16'd21741, 16'd41266, 16'd3155, 16'd11524, 16'd14627, 16'd29176, 16'd44323, 16'd26887, 16'd42706, 16'd11853, 16'd29264, 16'd15785});
	test_expansion(128'hd934bf90526d17688f024ba84cb66b1d, {16'd15600, 16'd17752, 16'd5032, 16'd37458, 16'd58666, 16'd19978, 16'd50517, 16'd36807, 16'd6660, 16'd50961, 16'd9890, 16'd16758, 16'd59936, 16'd15623, 16'd7255, 16'd20192, 16'd50593, 16'd46106, 16'd34644, 16'd39212, 16'd39537, 16'd63857, 16'd193, 16'd53914, 16'd28443, 16'd26253});
	test_expansion(128'hf1e8b3a589d1d5de0c3052da837b6c98, {16'd13410, 16'd17963, 16'd31776, 16'd8946, 16'd17238, 16'd22280, 16'd22270, 16'd53593, 16'd52322, 16'd65392, 16'd63381, 16'd52629, 16'd44534, 16'd56753, 16'd37965, 16'd62469, 16'd36917, 16'd51179, 16'd35520, 16'd7693, 16'd29341, 16'd31050, 16'd870, 16'd43168, 16'd13977, 16'd54704});
	test_expansion(128'h78fd1b1d4e80e026b7eaccc3f8ae4d2a, {16'd27072, 16'd40182, 16'd35926, 16'd27869, 16'd5859, 16'd31108, 16'd32866, 16'd20818, 16'd57370, 16'd25288, 16'd42038, 16'd27012, 16'd63630, 16'd58075, 16'd3970, 16'd65223, 16'd56257, 16'd45604, 16'd24323, 16'd57118, 16'd11737, 16'd4544, 16'd61943, 16'd6289, 16'd16510, 16'd15107});
	test_expansion(128'haeeee1e30845fc3a9b136ed4afb97b76, {16'd60469, 16'd9727, 16'd13179, 16'd32993, 16'd245, 16'd59685, 16'd62758, 16'd11546, 16'd11842, 16'd61529, 16'd4651, 16'd38557, 16'd11995, 16'd53714, 16'd54012, 16'd13288, 16'd21521, 16'd63612, 16'd54339, 16'd29484, 16'd6637, 16'd27082, 16'd31428, 16'd37341, 16'd20958, 16'd59687});
	test_expansion(128'h4ed78d0f7b2de4fa71510c0d86ae86ce, {16'd17949, 16'd47965, 16'd62006, 16'd816, 16'd48111, 16'd67, 16'd52106, 16'd40927, 16'd30136, 16'd57957, 16'd18876, 16'd62492, 16'd58058, 16'd8101, 16'd30965, 16'd9125, 16'd25979, 16'd33137, 16'd4007, 16'd32013, 16'd43991, 16'd20091, 16'd59627, 16'd2125, 16'd8319, 16'd35305});
	test_expansion(128'h43d21045c93f6aa15d621a00eb920cfd, {16'd28552, 16'd15141, 16'd58812, 16'd43825, 16'd6920, 16'd48977, 16'd16478, 16'd24554, 16'd58806, 16'd16362, 16'd28201, 16'd51199, 16'd12071, 16'd22846, 16'd4042, 16'd9036, 16'd46905, 16'd7096, 16'd18941, 16'd63537, 16'd26152, 16'd4269, 16'd20612, 16'd48328, 16'd58124, 16'd42311});
	test_expansion(128'h77c4d64ac8456a39d08d322ccf0cdf04, {16'd31123, 16'd17855, 16'd52855, 16'd19266, 16'd50927, 16'd28147, 16'd20381, 16'd576, 16'd48182, 16'd29125, 16'd40468, 16'd11511, 16'd20653, 16'd56773, 16'd24993, 16'd24984, 16'd52393, 16'd15819, 16'd4586, 16'd33204, 16'd14930, 16'd25921, 16'd49727, 16'd9379, 16'd33917, 16'd59663});
	test_expansion(128'h5cecc3b70e3c254ca603e9087645f23b, {16'd14309, 16'd52298, 16'd48659, 16'd29866, 16'd58043, 16'd1346, 16'd18081, 16'd49254, 16'd27365, 16'd50253, 16'd50767, 16'd64686, 16'd57689, 16'd63532, 16'd30829, 16'd1054, 16'd40284, 16'd62605, 16'd31333, 16'd30143, 16'd64677, 16'd35492, 16'd59583, 16'd23687, 16'd63765, 16'd4905});
	test_expansion(128'he0772cf004ce81768159cc66a9833f6d, {16'd11515, 16'd63141, 16'd31075, 16'd46735, 16'd38725, 16'd23439, 16'd29411, 16'd55683, 16'd61542, 16'd34184, 16'd43473, 16'd54521, 16'd29691, 16'd54536, 16'd9028, 16'd47075, 16'd19346, 16'd10982, 16'd42147, 16'd61246, 16'd40646, 16'd56863, 16'd33505, 16'd16350, 16'd9699, 16'd26187});
	test_expansion(128'h053a861eb62227bcf489fe07d413ccfc, {16'd33791, 16'd9767, 16'd58781, 16'd54172, 16'd18153, 16'd21173, 16'd47639, 16'd30947, 16'd54761, 16'd26049, 16'd3728, 16'd39441, 16'd38970, 16'd50245, 16'd23936, 16'd47761, 16'd20369, 16'd38232, 16'd21931, 16'd1342, 16'd3098, 16'd37754, 16'd11805, 16'd8220, 16'd41017, 16'd53936});
	test_expansion(128'hd0f1cdcd2befc1d5b502f981c33fa7ed, {16'd36013, 16'd41182, 16'd63641, 16'd64268, 16'd33824, 16'd21232, 16'd28159, 16'd25791, 16'd65093, 16'd30892, 16'd754, 16'd516, 16'd25821, 16'd23406, 16'd22942, 16'd12045, 16'd6453, 16'd17791, 16'd57625, 16'd35210, 16'd60539, 16'd13428, 16'd34610, 16'd58631, 16'd51338, 16'd10960});
	test_expansion(128'h8de1fddb88d622bb2a4b2ed09cd5fc61, {16'd22297, 16'd64580, 16'd50023, 16'd6805, 16'd57243, 16'd14798, 16'd61667, 16'd61110, 16'd26863, 16'd63125, 16'd10943, 16'd35557, 16'd62415, 16'd19339, 16'd56558, 16'd17112, 16'd16343, 16'd12939, 16'd19163, 16'd38446, 16'd22984, 16'd50188, 16'd26921, 16'd32819, 16'd25205, 16'd8770});
	test_expansion(128'hd5b340cbafcea976e5cc2eb803b0bbac, {16'd61679, 16'd34083, 16'd55389, 16'd48110, 16'd44742, 16'd37606, 16'd3416, 16'd45719, 16'd22667, 16'd54530, 16'd37357, 16'd56206, 16'd18380, 16'd15566, 16'd34190, 16'd9586, 16'd63049, 16'd59616, 16'd31790, 16'd33285, 16'd18529, 16'd62339, 16'd56622, 16'd63670, 16'd12400, 16'd44909});
	test_expansion(128'hf98dcc0282787dea2b730aea79543aa0, {16'd49623, 16'd40798, 16'd15174, 16'd12505, 16'd56985, 16'd17396, 16'd56190, 16'd31412, 16'd6068, 16'd2180, 16'd18764, 16'd7629, 16'd36956, 16'd1562, 16'd30140, 16'd17582, 16'd59959, 16'd8453, 16'd15016, 16'd61702, 16'd56562, 16'd38503, 16'd21308, 16'd17031, 16'd22822, 16'd45670});
	test_expansion(128'h0926ae525b69575669f430476c6d9b52, {16'd44859, 16'd34733, 16'd1792, 16'd30317, 16'd16258, 16'd60851, 16'd47752, 16'd55157, 16'd58073, 16'd47811, 16'd15182, 16'd64249, 16'd11883, 16'd55712, 16'd7152, 16'd33500, 16'd50617, 16'd1935, 16'd20482, 16'd63156, 16'd19229, 16'd19663, 16'd26057, 16'd10086, 16'd13872, 16'd41437});
	test_expansion(128'hfeed2e86dc722bfdc8bc3df749f1fb7b, {16'd37548, 16'd14723, 16'd30674, 16'd26058, 16'd5029, 16'd2252, 16'd7448, 16'd39455, 16'd55568, 16'd63752, 16'd60298, 16'd39499, 16'd11933, 16'd49518, 16'd42302, 16'd44614, 16'd52865, 16'd61912, 16'd22071, 16'd44733, 16'd51307, 16'd35147, 16'd16767, 16'd28041, 16'd46646, 16'd60786});
	test_expansion(128'h55f488275365b90b0a240ba622066dbd, {16'd18045, 16'd12274, 16'd53630, 16'd29826, 16'd31384, 16'd2229, 16'd40358, 16'd39400, 16'd6788, 16'd47148, 16'd18680, 16'd14681, 16'd32516, 16'd6136, 16'd47277, 16'd14326, 16'd41410, 16'd30994, 16'd26722, 16'd35823, 16'd7082, 16'd9349, 16'd30137, 16'd15697, 16'd26219, 16'd48957});
	test_expansion(128'he6ebaeac345b6d1a2cc17e8cde7a01a6, {16'd11738, 16'd53748, 16'd28789, 16'd53892, 16'd57234, 16'd39569, 16'd27126, 16'd34978, 16'd33655, 16'd820, 16'd23516, 16'd31797, 16'd42891, 16'd8857, 16'd19000, 16'd7320, 16'd57669, 16'd22441, 16'd3303, 16'd3478, 16'd11774, 16'd29089, 16'd15854, 16'd33164, 16'd64951, 16'd53380});
	test_expansion(128'h3cf7f01dadb1f3a5979451cbeaace9c5, {16'd3118, 16'd44517, 16'd39962, 16'd8234, 16'd57652, 16'd41446, 16'd39900, 16'd28200, 16'd64752, 16'd60189, 16'd18935, 16'd36947, 16'd28821, 16'd56342, 16'd2730, 16'd62134, 16'd22126, 16'd26471, 16'd43068, 16'd53002, 16'd37754, 16'd49153, 16'd59667, 16'd3136, 16'd24196, 16'd64794});
	test_expansion(128'h876e3c05fd71b3194f506bd6928eb44b, {16'd56562, 16'd13412, 16'd55818, 16'd40384, 16'd715, 16'd58781, 16'd51150, 16'd6765, 16'd45599, 16'd30771, 16'd37086, 16'd21208, 16'd46921, 16'd44928, 16'd2947, 16'd54682, 16'd8303, 16'd54104, 16'd59939, 16'd28661, 16'd38436, 16'd9743, 16'd27406, 16'd48698, 16'd58898, 16'd42318});
	test_expansion(128'h0d95380c922ca32646f7900d05e3a8f2, {16'd35686, 16'd57321, 16'd51294, 16'd19245, 16'd31615, 16'd37065, 16'd29879, 16'd50256, 16'd26934, 16'd30541, 16'd24383, 16'd47176, 16'd11601, 16'd51156, 16'd14190, 16'd49759, 16'd29731, 16'd22342, 16'd48961, 16'd54748, 16'd11019, 16'd43008, 16'd29334, 16'd17277, 16'd11698, 16'd555});
	test_expansion(128'hb11da6561e6e6e015015f56d5283d5fd, {16'd47359, 16'd20873, 16'd9707, 16'd58340, 16'd10000, 16'd60576, 16'd31513, 16'd36261, 16'd25996, 16'd22746, 16'd8045, 16'd6846, 16'd43678, 16'd32884, 16'd12571, 16'd48176, 16'd40274, 16'd16775, 16'd53182, 16'd27274, 16'd47005, 16'd34632, 16'd2804, 16'd22526, 16'd5982, 16'd61165});
	test_expansion(128'had71bdf49dbe6a3a9267b2b52e794906, {16'd2436, 16'd18628, 16'd49277, 16'd37472, 16'd37087, 16'd60729, 16'd47081, 16'd16818, 16'd52213, 16'd20850, 16'd29869, 16'd45831, 16'd53890, 16'd22281, 16'd58464, 16'd2097, 16'd7904, 16'd29097, 16'd30246, 16'd64515, 16'd46570, 16'd23716, 16'd54281, 16'd62270, 16'd32269, 16'd58475});
	test_expansion(128'h67051f273f15a1139c915266a7a3fbe5, {16'd35414, 16'd51484, 16'd32544, 16'd31673, 16'd32290, 16'd7502, 16'd59012, 16'd6045, 16'd27463, 16'd25787, 16'd64348, 16'd14298, 16'd5485, 16'd30744, 16'd49538, 16'd46931, 16'd21709, 16'd39935, 16'd14619, 16'd65004, 16'd47704, 16'd42089, 16'd43940, 16'd12345, 16'd1265, 16'd39539});
	test_expansion(128'h207c0bc410508dcb6c9282f40155f4dc, {16'd17489, 16'd41145, 16'd57978, 16'd199, 16'd10372, 16'd57476, 16'd15693, 16'd33988, 16'd49043, 16'd34835, 16'd20109, 16'd22723, 16'd6510, 16'd53603, 16'd55224, 16'd37823, 16'd4123, 16'd27054, 16'd27599, 16'd40487, 16'd20862, 16'd41784, 16'd6056, 16'd2609, 16'd45078, 16'd48448});
	test_expansion(128'h597f48942a7f113eceb72b2d1c2282cc, {16'd53810, 16'd47759, 16'd62613, 16'd57824, 16'd56545, 16'd32951, 16'd33880, 16'd25255, 16'd50569, 16'd34254, 16'd56625, 16'd63063, 16'd36948, 16'd20411, 16'd50483, 16'd46725, 16'd16617, 16'd28203, 16'd36153, 16'd32601, 16'd18463, 16'd5159, 16'd35680, 16'd10200, 16'd59189, 16'd7387});
	test_expansion(128'h133627e7f75c1e8358b64b03fcb5b119, {16'd25239, 16'd8801, 16'd37475, 16'd31050, 16'd19461, 16'd61059, 16'd62598, 16'd15063, 16'd38095, 16'd64972, 16'd32189, 16'd23098, 16'd324, 16'd22881, 16'd7654, 16'd30964, 16'd1002, 16'd36747, 16'd9350, 16'd14776, 16'd25597, 16'd9462, 16'd52055, 16'd25950, 16'd38787, 16'd2894});
	test_expansion(128'h599208c4221ea4c45c8ae0f8de51686a, {16'd15098, 16'd47757, 16'd43758, 16'd48845, 16'd29135, 16'd46338, 16'd6569, 16'd58658, 16'd65082, 16'd64566, 16'd20624, 16'd13575, 16'd5011, 16'd59871, 16'd52871, 16'd18457, 16'd257, 16'd64564, 16'd40085, 16'd40793, 16'd3232, 16'd55846, 16'd44415, 16'd52859, 16'd5744, 16'd7697});
	test_expansion(128'h6f3c2ce76de9acc099e0b1489174c78e, {16'd51604, 16'd17270, 16'd52322, 16'd1490, 16'd25320, 16'd13750, 16'd20989, 16'd47918, 16'd37396, 16'd45719, 16'd24424, 16'd39967, 16'd29442, 16'd48425, 16'd54944, 16'd2182, 16'd18303, 16'd38498, 16'd24629, 16'd1034, 16'd8753, 16'd39041, 16'd18078, 16'd10426, 16'd24237, 16'd53108});
	test_expansion(128'he95980cfc82fb2860180b1fc89eb3e20, {16'd29428, 16'd30188, 16'd21407, 16'd14537, 16'd45664, 16'd5844, 16'd20852, 16'd64006, 16'd484, 16'd6642, 16'd46576, 16'd21044, 16'd2271, 16'd58235, 16'd36153, 16'd53773, 16'd46930, 16'd34190, 16'd39437, 16'd47643, 16'd28789, 16'd33149, 16'd3485, 16'd27067, 16'd22128, 16'd31412});
	test_expansion(128'h1d83c0c7cbdf51a8fb787ccb86193f4f, {16'd8792, 16'd22020, 16'd36260, 16'd56858, 16'd33839, 16'd13624, 16'd56468, 16'd48448, 16'd58847, 16'd6054, 16'd60838, 16'd25731, 16'd28229, 16'd60474, 16'd13572, 16'd47481, 16'd38352, 16'd18864, 16'd49418, 16'd52367, 16'd42854, 16'd1447, 16'd34805, 16'd27860, 16'd4181, 16'd37298});
	test_expansion(128'hdddb3d448c6b761fff4b0e5e71b51842, {16'd11041, 16'd9436, 16'd19415, 16'd13632, 16'd9814, 16'd29617, 16'd43860, 16'd61086, 16'd16354, 16'd34162, 16'd27152, 16'd36175, 16'd34194, 16'd49428, 16'd5412, 16'd23768, 16'd18265, 16'd27555, 16'd49446, 16'd42041, 16'd55217, 16'd48355, 16'd20327, 16'd25160, 16'd30783, 16'd46355});
	test_expansion(128'hb9c758256060fa096100ee6abc719750, {16'd30234, 16'd53748, 16'd40490, 16'd28567, 16'd63063, 16'd47901, 16'd17499, 16'd45688, 16'd61982, 16'd64791, 16'd6794, 16'd35465, 16'd9350, 16'd10528, 16'd722, 16'd59028, 16'd35915, 16'd34085, 16'd2218, 16'd3107, 16'd22264, 16'd17033, 16'd18148, 16'd62322, 16'd39295, 16'd2204});
	test_expansion(128'h6c0fca14178b9505bddcf31ac156c820, {16'd188, 16'd64795, 16'd19864, 16'd57296, 16'd5111, 16'd33760, 16'd20500, 16'd45846, 16'd53470, 16'd963, 16'd10841, 16'd11318, 16'd33959, 16'd35623, 16'd13243, 16'd32570, 16'd55869, 16'd17355, 16'd39696, 16'd37719, 16'd47241, 16'd60574, 16'd12861, 16'd41404, 16'd34819, 16'd47416});
	test_expansion(128'h5bb0a313eceb64472c5a962a906bc763, {16'd56584, 16'd41778, 16'd41651, 16'd14247, 16'd46719, 16'd50753, 16'd24872, 16'd16943, 16'd27199, 16'd37735, 16'd52521, 16'd12382, 16'd54075, 16'd38402, 16'd6494, 16'd15467, 16'd46697, 16'd54224, 16'd57854, 16'd58260, 16'd63015, 16'd61678, 16'd34881, 16'd61267, 16'd20522, 16'd55656});
	test_expansion(128'h563f1872b0cb97ffca69cc17e482a60a, {16'd14017, 16'd63908, 16'd22316, 16'd12647, 16'd25443, 16'd9945, 16'd35581, 16'd6922, 16'd33380, 16'd62373, 16'd45802, 16'd59200, 16'd37939, 16'd20326, 16'd57753, 16'd12559, 16'd32186, 16'd13300, 16'd1860, 16'd12805, 16'd54114, 16'd14912, 16'd8599, 16'd50422, 16'd13136, 16'd18253});
	test_expansion(128'hed52adff5a7298bc1eb8db4c0e50f1f9, {16'd9189, 16'd16601, 16'd62033, 16'd45415, 16'd979, 16'd752, 16'd58165, 16'd2558, 16'd51467, 16'd18179, 16'd48322, 16'd36329, 16'd41329, 16'd27327, 16'd13778, 16'd62996, 16'd11567, 16'd61428, 16'd39187, 16'd43756, 16'd28853, 16'd641, 16'd30719, 16'd57697, 16'd37150, 16'd29197});
	test_expansion(128'h5dd4a0a1fadb2212878f7f5cf33b5ebb, {16'd10797, 16'd55450, 16'd13262, 16'd5373, 16'd56579, 16'd53299, 16'd35221, 16'd64518, 16'd64940, 16'd32639, 16'd50708, 16'd39956, 16'd41050, 16'd16064, 16'd58120, 16'd28069, 16'd39513, 16'd16108, 16'd27019, 16'd36577, 16'd25297, 16'd41702, 16'd27706, 16'd21232, 16'd14091, 16'd39245});
	test_expansion(128'he0be742186157321966291ecd364f4e7, {16'd35793, 16'd32684, 16'd6615, 16'd25984, 16'd14604, 16'd60276, 16'd44158, 16'd37137, 16'd21976, 16'd56288, 16'd36993, 16'd6161, 16'd33700, 16'd18980, 16'd43706, 16'd21089, 16'd46506, 16'd16626, 16'd29277, 16'd53460, 16'd10543, 16'd1434, 16'd1406, 16'd59578, 16'd10249, 16'd10432});
	test_expansion(128'h6f037a08a2396c00d612fde4232c5758, {16'd23785, 16'd42334, 16'd25049, 16'd47713, 16'd7978, 16'd21599, 16'd19923, 16'd8158, 16'd32363, 16'd24965, 16'd14675, 16'd47175, 16'd56766, 16'd61166, 16'd48067, 16'd63800, 16'd8533, 16'd61811, 16'd17779, 16'd3092, 16'd1204, 16'd57828, 16'd51782, 16'd11754, 16'd60992, 16'd20629});
	test_expansion(128'h7c9d2d488cf9d1bfb59dc1bdeeb9a54c, {16'd24069, 16'd18993, 16'd64699, 16'd54942, 16'd12207, 16'd31209, 16'd22061, 16'd20110, 16'd23736, 16'd38247, 16'd35391, 16'd48294, 16'd19416, 16'd10213, 16'd1379, 16'd11503, 16'd63345, 16'd55457, 16'd32141, 16'd53440, 16'd15728, 16'd11894, 16'd56086, 16'd31644, 16'd43157, 16'd18787});
	test_expansion(128'h28c280e3629f3712e5edcc022b10dcb3, {16'd44066, 16'd24712, 16'd6464, 16'd31047, 16'd4731, 16'd49111, 16'd30009, 16'd60285, 16'd59823, 16'd45291, 16'd54322, 16'd28951, 16'd42331, 16'd29245, 16'd38900, 16'd40576, 16'd51687, 16'd31466, 16'd49598, 16'd40912, 16'd21519, 16'd2966, 16'd4764, 16'd27850, 16'd22107, 16'd11809});
	test_expansion(128'h15393f3a1905abdf6bd6ccf4ae934000, {16'd24194, 16'd15223, 16'd6931, 16'd37059, 16'd38903, 16'd29385, 16'd28326, 16'd30430, 16'd58942, 16'd28191, 16'd7906, 16'd34793, 16'd51587, 16'd56575, 16'd45948, 16'd58504, 16'd23045, 16'd48333, 16'd23344, 16'd35350, 16'd64387, 16'd25254, 16'd44847, 16'd30303, 16'd13309, 16'd25913});
	test_expansion(128'hb4f0a2237eec0bfcc8d4c47ae92f125b, {16'd53799, 16'd32746, 16'd48191, 16'd60678, 16'd49251, 16'd61533, 16'd9247, 16'd29886, 16'd3591, 16'd44892, 16'd31704, 16'd45098, 16'd19034, 16'd28065, 16'd50490, 16'd15008, 16'd40084, 16'd1126, 16'd11754, 16'd31076, 16'd8441, 16'd17667, 16'd55991, 16'd62722, 16'd45447, 16'd61306});
	test_expansion(128'h702c5691bf511104ba0e015b7237404e, {16'd18725, 16'd7665, 16'd35522, 16'd47098, 16'd28657, 16'd3352, 16'd40692, 16'd47831, 16'd53374, 16'd41284, 16'd23539, 16'd45236, 16'd23553, 16'd50087, 16'd51946, 16'd57613, 16'd34615, 16'd33946, 16'd62294, 16'd33407, 16'd12552, 16'd52572, 16'd806, 16'd8417, 16'd57285, 16'd46501});
	test_expansion(128'h87dc9d2d4b4ff4e7e141b3f0cfaedd6c, {16'd36491, 16'd21907, 16'd32485, 16'd42637, 16'd55053, 16'd2902, 16'd2809, 16'd17463, 16'd10485, 16'd33761, 16'd43778, 16'd40027, 16'd15279, 16'd34820, 16'd10781, 16'd50424, 16'd49160, 16'd60061, 16'd55210, 16'd6994, 16'd26069, 16'd32865, 16'd17888, 16'd12567, 16'd19650, 16'd13487});
	test_expansion(128'hc116375e746a8b596616c7410f791330, {16'd17081, 16'd25561, 16'd56720, 16'd14696, 16'd36805, 16'd47259, 16'd35373, 16'd52548, 16'd27095, 16'd34966, 16'd15805, 16'd22314, 16'd771, 16'd42485, 16'd47900, 16'd46051, 16'd65107, 16'd46209, 16'd48481, 16'd4674, 16'd44411, 16'd15761, 16'd9325, 16'd45792, 16'd56830, 16'd38915});
	test_expansion(128'h39900a46cb94814251c158f1229c7bd1, {16'd58283, 16'd4521, 16'd8623, 16'd39555, 16'd34890, 16'd12069, 16'd8862, 16'd4920, 16'd32019, 16'd45478, 16'd63854, 16'd54446, 16'd17724, 16'd24625, 16'd27345, 16'd29005, 16'd14186, 16'd49648, 16'd54130, 16'd33249, 16'd62202, 16'd27061, 16'd59440, 16'd26208, 16'd52910, 16'd1453});
	test_expansion(128'h94de8d66b2f23cdd398b8b1837cb0aae, {16'd3507, 16'd33457, 16'd18153, 16'd35543, 16'd25307, 16'd7010, 16'd6166, 16'd59142, 16'd33075, 16'd20091, 16'd56869, 16'd15586, 16'd53052, 16'd11835, 16'd18967, 16'd38208, 16'd43601, 16'd33907, 16'd44973, 16'd42687, 16'd16567, 16'd47044, 16'd25453, 16'd19481, 16'd16427, 16'd32025});
	test_expansion(128'h7083f8b4442381b66e8218efccc01591, {16'd29037, 16'd59164, 16'd19894, 16'd22757, 16'd21255, 16'd710, 16'd1456, 16'd13283, 16'd49134, 16'd1620, 16'd39614, 16'd17289, 16'd23017, 16'd9128, 16'd33741, 16'd31796, 16'd52945, 16'd63384, 16'd6882, 16'd44150, 16'd52515, 16'd32290, 16'd4257, 16'd43991, 16'd37178, 16'd16676});
	test_expansion(128'h9b71a650c1c25a96a72c043faeaa8f7f, {16'd47259, 16'd25978, 16'd11381, 16'd24301, 16'd37836, 16'd64461, 16'd24076, 16'd59891, 16'd9245, 16'd54902, 16'd55025, 16'd46549, 16'd36795, 16'd14461, 16'd33098, 16'd18776, 16'd6142, 16'd60985, 16'd42403, 16'd60756, 16'd59426, 16'd16800, 16'd13780, 16'd20968, 16'd29989, 16'd3131});
	test_expansion(128'h89e703945ed5a30437ad547a44af5b8f, {16'd65518, 16'd45425, 16'd48785, 16'd9102, 16'd54580, 16'd51666, 16'd24498, 16'd46222, 16'd26769, 16'd56623, 16'd42737, 16'd21142, 16'd41672, 16'd32920, 16'd48357, 16'd27626, 16'd62076, 16'd24695, 16'd62479, 16'd24852, 16'd20009, 16'd62725, 16'd45042, 16'd36366, 16'd47218, 16'd14354});
	test_expansion(128'h345cf1343771508ed527df9595d53758, {16'd57895, 16'd1323, 16'd6209, 16'd43558, 16'd43501, 16'd56112, 16'd16058, 16'd44378, 16'd59967, 16'd15439, 16'd21904, 16'd36648, 16'd64312, 16'd15695, 16'd32638, 16'd363, 16'd27733, 16'd18906, 16'd8142, 16'd45909, 16'd60338, 16'd58508, 16'd49091, 16'd60226, 16'd35098, 16'd49264});
	test_expansion(128'hcb2fa7fac9696f2bc9fddb90ddfe2a23, {16'd39552, 16'd58505, 16'd13803, 16'd30247, 16'd14167, 16'd59141, 16'd29751, 16'd45959, 16'd12022, 16'd26144, 16'd16410, 16'd45148, 16'd22607, 16'd48928, 16'd45503, 16'd29179, 16'd26208, 16'd21755, 16'd53789, 16'd31574, 16'd28225, 16'd37621, 16'd20656, 16'd21883, 16'd12722, 16'd47350});
	test_expansion(128'hab188cc294465bb61a92e28272c2f518, {16'd28714, 16'd45285, 16'd11614, 16'd27399, 16'd63518, 16'd25577, 16'd32036, 16'd36532, 16'd38643, 16'd36008, 16'd25965, 16'd27088, 16'd22707, 16'd9066, 16'd46539, 16'd32659, 16'd3046, 16'd47612, 16'd5289, 16'd47051, 16'd5982, 16'd65525, 16'd32811, 16'd36548, 16'd19577, 16'd10863});
	test_expansion(128'h2d97dd31849215aabab2c2aedb4a65f2, {16'd5615, 16'd62473, 16'd50915, 16'd43766, 16'd25979, 16'd32897, 16'd59570, 16'd57019, 16'd49186, 16'd6106, 16'd29723, 16'd27917, 16'd34645, 16'd1896, 16'd2681, 16'd52259, 16'd50440, 16'd4900, 16'd65134, 16'd44299, 16'd59266, 16'd25055, 16'd36023, 16'd57785, 16'd53802, 16'd60287});
	test_expansion(128'hd600769df4120c3c8da09421e7b04819, {16'd11813, 16'd9042, 16'd29480, 16'd47472, 16'd48112, 16'd7025, 16'd42935, 16'd4361, 16'd55274, 16'd65262, 16'd37531, 16'd21708, 16'd49543, 16'd36945, 16'd27859, 16'd15616, 16'd11086, 16'd58751, 16'd53138, 16'd50626, 16'd45731, 16'd34690, 16'd5306, 16'd40593, 16'd24224, 16'd946});
	test_expansion(128'h601460fc428575f75011dccd6998dd19, {16'd26467, 16'd36384, 16'd60528, 16'd39368, 16'd19255, 16'd22029, 16'd47226, 16'd63817, 16'd14728, 16'd3498, 16'd39130, 16'd61913, 16'd7300, 16'd15833, 16'd17646, 16'd23783, 16'd52953, 16'd49308, 16'd40522, 16'd26687, 16'd62336, 16'd34930, 16'd45005, 16'd47276, 16'd15647, 16'd64478});
	test_expansion(128'he9ca65f3ea147ceec502630ac15cf561, {16'd16303, 16'd8595, 16'd56092, 16'd13910, 16'd45801, 16'd36296, 16'd58661, 16'd11760, 16'd18654, 16'd22874, 16'd651, 16'd24259, 16'd56325, 16'd19304, 16'd26099, 16'd42957, 16'd1206, 16'd5218, 16'd49363, 16'd32607, 16'd26365, 16'd3496, 16'd21037, 16'd25462, 16'd15928, 16'd49801});
	test_expansion(128'h7c76c5e5f95d2e705a6fa0979487e860, {16'd42645, 16'd2083, 16'd38273, 16'd38037, 16'd54888, 16'd26616, 16'd13526, 16'd447, 16'd16156, 16'd49821, 16'd35873, 16'd53486, 16'd38794, 16'd39009, 16'd60877, 16'd32489, 16'd3484, 16'd1442, 16'd17102, 16'd4020, 16'd9633, 16'd46603, 16'd28619, 16'd6644, 16'd10396, 16'd64831});
	test_expansion(128'h2e85701923607ad0789f6210dc317f03, {16'd44077, 16'd64125, 16'd8797, 16'd11632, 16'd52702, 16'd48544, 16'd54739, 16'd47451, 16'd17892, 16'd52724, 16'd56538, 16'd12371, 16'd31034, 16'd18765, 16'd17534, 16'd41786, 16'd21740, 16'd45593, 16'd12962, 16'd29590, 16'd29516, 16'd56874, 16'd17234, 16'd29655, 16'd51679, 16'd21413});
	test_expansion(128'h96620c243ca02b4cb46794228b4c341c, {16'd41790, 16'd17639, 16'd54795, 16'd5019, 16'd38187, 16'd26776, 16'd38789, 16'd5928, 16'd33139, 16'd11484, 16'd38606, 16'd22361, 16'd35873, 16'd36682, 16'd8791, 16'd23939, 16'd5147, 16'd49580, 16'd1631, 16'd27162, 16'd32639, 16'd1006, 16'd23422, 16'd23018, 16'd31136, 16'd57984});
	test_expansion(128'hf090ad144006e2c2acc898709c2efbf2, {16'd31384, 16'd54002, 16'd55475, 16'd52932, 16'd48744, 16'd19896, 16'd58041, 16'd16089, 16'd1624, 16'd49878, 16'd39622, 16'd19887, 16'd59574, 16'd36776, 16'd19377, 16'd43821, 16'd64468, 16'd17485, 16'd15984, 16'd15597, 16'd295, 16'd6442, 16'd18470, 16'd55913, 16'd50053, 16'd28358});
	test_expansion(128'h243210c82b76de4983697727d94b6bf0, {16'd34681, 16'd28599, 16'd59033, 16'd35883, 16'd31672, 16'd53111, 16'd17692, 16'd13472, 16'd8760, 16'd10099, 16'd17085, 16'd9165, 16'd15212, 16'd48405, 16'd20949, 16'd6870, 16'd26803, 16'd35136, 16'd2802, 16'd29809, 16'd44694, 16'd55092, 16'd33784, 16'd56720, 16'd65063, 16'd4960});
	test_expansion(128'h873e63852f94e3b9eab316a0b30b7b3e, {16'd53768, 16'd11967, 16'd53926, 16'd44358, 16'd31605, 16'd59913, 16'd9355, 16'd13603, 16'd8339, 16'd1698, 16'd60224, 16'd25388, 16'd18765, 16'd15430, 16'd42316, 16'd9809, 16'd148, 16'd49968, 16'd29218, 16'd18946, 16'd53690, 16'd19764, 16'd17732, 16'd53771, 16'd24912, 16'd65024});
	test_expansion(128'heed4a7c28bb142e636ca24b19c90edd5, {16'd35508, 16'd47173, 16'd11911, 16'd32582, 16'd14929, 16'd32409, 16'd12740, 16'd36920, 16'd10124, 16'd10433, 16'd25163, 16'd7836, 16'd32331, 16'd34818, 16'd11693, 16'd46701, 16'd46165, 16'd15595, 16'd30240, 16'd36966, 16'd20900, 16'd4665, 16'd10907, 16'd4711, 16'd12362, 16'd26348});
	test_expansion(128'h7f3a28ca859365e6e723e444b946fbd9, {16'd15369, 16'd53837, 16'd26150, 16'd22642, 16'd17320, 16'd14728, 16'd59086, 16'd56035, 16'd53728, 16'd37987, 16'd7753, 16'd41947, 16'd35206, 16'd50046, 16'd4586, 16'd41037, 16'd7642, 16'd3863, 16'd2364, 16'd26212, 16'd43774, 16'd22426, 16'd34798, 16'd59006, 16'd13438, 16'd13382});
	test_expansion(128'h5d0a2d11bde2d05c946e343d7ad8097d, {16'd31678, 16'd47492, 16'd24520, 16'd58478, 16'd42411, 16'd62165, 16'd5227, 16'd2553, 16'd10224, 16'd31196, 16'd61306, 16'd16692, 16'd3538, 16'd35769, 16'd30863, 16'd29145, 16'd5484, 16'd48016, 16'd42370, 16'd60170, 16'd48134, 16'd40845, 16'd54969, 16'd6213, 16'd26379, 16'd31473});
	test_expansion(128'h0a194da193c32d202728af754416e90a, {16'd1282, 16'd35515, 16'd60817, 16'd59316, 16'd49230, 16'd53413, 16'd48608, 16'd57095, 16'd31498, 16'd54160, 16'd60111, 16'd22669, 16'd18819, 16'd49782, 16'd15880, 16'd16061, 16'd2006, 16'd51700, 16'd51447, 16'd21016, 16'd27792, 16'd31781, 16'd63445, 16'd12381, 16'd56044, 16'd52365});
	test_expansion(128'hc36886f0cd653acbed974cd208616eb3, {16'd7936, 16'd50166, 16'd4946, 16'd47799, 16'd36746, 16'd24806, 16'd5912, 16'd8408, 16'd1778, 16'd59809, 16'd3782, 16'd51371, 16'd40018, 16'd22800, 16'd28516, 16'd25579, 16'd27161, 16'd21172, 16'd33214, 16'd26404, 16'd49312, 16'd2376, 16'd2373, 16'd30681, 16'd6417, 16'd9586});
	test_expansion(128'h134e367f01752ae823224365573c0231, {16'd21356, 16'd2592, 16'd59824, 16'd55623, 16'd64364, 16'd41927, 16'd11563, 16'd52490, 16'd34502, 16'd64114, 16'd61353, 16'd60178, 16'd63707, 16'd51415, 16'd18713, 16'd40880, 16'd63849, 16'd1034, 16'd56531, 16'd5266, 16'd21035, 16'd5018, 16'd49840, 16'd36870, 16'd58011, 16'd22309});
	test_expansion(128'h9d19cd2f5e355436e42fb3da7a2a7b44, {16'd17641, 16'd8846, 16'd43851, 16'd60651, 16'd58927, 16'd4095, 16'd19154, 16'd52044, 16'd39814, 16'd34823, 16'd3742, 16'd15022, 16'd50979, 16'd38424, 16'd14513, 16'd9131, 16'd19062, 16'd6780, 16'd39193, 16'd51434, 16'd55587, 16'd45854, 16'd11811, 16'd31687, 16'd43341, 16'd31802});
	test_expansion(128'hb8d0c0a7f4712f5d517ca8fc99604b60, {16'd940, 16'd35345, 16'd17408, 16'd64442, 16'd58439, 16'd42041, 16'd49478, 16'd3170, 16'd35113, 16'd32396, 16'd13318, 16'd60211, 16'd52661, 16'd12318, 16'd27012, 16'd5795, 16'd17105, 16'd242, 16'd33292, 16'd30403, 16'd60937, 16'd48887, 16'd46441, 16'd60282, 16'd22144, 16'd16349});
	test_expansion(128'hbfe8132c791bb8b213f12f777dd4221a, {16'd38737, 16'd47082, 16'd22911, 16'd52961, 16'd24112, 16'd43726, 16'd59624, 16'd28091, 16'd58066, 16'd8042, 16'd30367, 16'd46776, 16'd34631, 16'd64888, 16'd62247, 16'd34736, 16'd31884, 16'd17728, 16'd35049, 16'd36448, 16'd51631, 16'd30486, 16'd44309, 16'd39629, 16'd42843, 16'd39801});
	test_expansion(128'h5b149448aabc58ea736e04b47d969737, {16'd51652, 16'd14271, 16'd62654, 16'd61352, 16'd45699, 16'd3046, 16'd53006, 16'd27596, 16'd29063, 16'd52596, 16'd5252, 16'd26854, 16'd24317, 16'd28147, 16'd54383, 16'd35336, 16'd35925, 16'd17071, 16'd63307, 16'd2846, 16'd33624, 16'd63548, 16'd13690, 16'd6478, 16'd32733, 16'd37321});
	test_expansion(128'ha329244830b55374f95d9797cc19c160, {16'd12065, 16'd35877, 16'd12597, 16'd3567, 16'd40468, 16'd27461, 16'd17160, 16'd23136, 16'd7964, 16'd44038, 16'd59634, 16'd25006, 16'd60479, 16'd4894, 16'd37115, 16'd26297, 16'd40725, 16'd23812, 16'd16491, 16'd44754, 16'd35469, 16'd39285, 16'd35722, 16'd56202, 16'd8698, 16'd8366});
	test_expansion(128'he050332e45c24d3e56a21f124f6e97a9, {16'd65378, 16'd50339, 16'd6091, 16'd36107, 16'd31833, 16'd32176, 16'd10660, 16'd43435, 16'd46569, 16'd43097, 16'd42387, 16'd5306, 16'd35018, 16'd2202, 16'd56216, 16'd16110, 16'd19133, 16'd1011, 16'd5144, 16'd7329, 16'd31338, 16'd3632, 16'd2353, 16'd5055, 16'd13574, 16'd12834});
	test_expansion(128'h6a110543676b9cebd555ce3878403aa7, {16'd9872, 16'd34780, 16'd13878, 16'd38090, 16'd14728, 16'd45628, 16'd30264, 16'd38884, 16'd2496, 16'd45152, 16'd2575, 16'd43249, 16'd35101, 16'd19262, 16'd23535, 16'd60887, 16'd10800, 16'd33632, 16'd212, 16'd20233, 16'd38660, 16'd24164, 16'd2005, 16'd48664, 16'd48260, 16'd41825});
	test_expansion(128'hb50b9e5edfaa9c1900217364eaceb054, {16'd48347, 16'd26583, 16'd65418, 16'd16965, 16'd63560, 16'd58786, 16'd10381, 16'd52494, 16'd50217, 16'd11949, 16'd51728, 16'd55583, 16'd55398, 16'd46798, 16'd64645, 16'd55071, 16'd58469, 16'd8489, 16'd32012, 16'd32091, 16'd14891, 16'd49004, 16'd30100, 16'd17078, 16'd3977, 16'd27493});
	test_expansion(128'h48caff812fcae29d8b56dd8ce37e7e5c, {16'd60253, 16'd62254, 16'd12073, 16'd65344, 16'd57345, 16'd53821, 16'd35502, 16'd3991, 16'd39803, 16'd26499, 16'd10055, 16'd10164, 16'd18008, 16'd64303, 16'd29987, 16'd31683, 16'd16712, 16'd49170, 16'd37118, 16'd63170, 16'd15115, 16'd22053, 16'd48024, 16'd30521, 16'd26894, 16'd43900});
	test_expansion(128'hbb10ca339596e455a12cf5c823381e20, {16'd52912, 16'd37499, 16'd14431, 16'd63799, 16'd17232, 16'd31660, 16'd2152, 16'd13861, 16'd35128, 16'd43033, 16'd37720, 16'd35600, 16'd32348, 16'd15473, 16'd20816, 16'd61153, 16'd54118, 16'd652, 16'd62330, 16'd4279, 16'd54026, 16'd3635, 16'd37262, 16'd41665, 16'd49860, 16'd21778});
	test_expansion(128'h1dd7b195f451b3bbc6ea786ac2002a17, {16'd20199, 16'd23901, 16'd41544, 16'd2549, 16'd34320, 16'd42255, 16'd18729, 16'd30947, 16'd33181, 16'd26222, 16'd17532, 16'd13377, 16'd10083, 16'd50532, 16'd58457, 16'd5436, 16'd48381, 16'd49503, 16'd64785, 16'd2766, 16'd54496, 16'd2637, 16'd7907, 16'd13304, 16'd10826, 16'd33650});
	test_expansion(128'h29d21e2bba51205c7be83d1dbddbf8fa, {16'd23030, 16'd6148, 16'd24943, 16'd25644, 16'd11389, 16'd28157, 16'd62805, 16'd43526, 16'd56225, 16'd15580, 16'd15172, 16'd18574, 16'd7086, 16'd28429, 16'd12625, 16'd6972, 16'd51470, 16'd21538, 16'd26809, 16'd37884, 16'd26173, 16'd61545, 16'd37277, 16'd11915, 16'd31755, 16'd27005});
	test_expansion(128'h0b0d9c4863e0d5151224fe83fa2a2d3d, {16'd50973, 16'd64558, 16'd50540, 16'd59, 16'd36028, 16'd34672, 16'd2728, 16'd34362, 16'd52306, 16'd60593, 16'd7953, 16'd55255, 16'd22025, 16'd17710, 16'd50865, 16'd44669, 16'd26362, 16'd5582, 16'd13896, 16'd1094, 16'd11870, 16'd1547, 16'd45424, 16'd36528, 16'd58852, 16'd61269});
	test_expansion(128'hc65b745ed9493932f2e5c010d103efc5, {16'd46004, 16'd49226, 16'd4265, 16'd36435, 16'd59190, 16'd15463, 16'd28973, 16'd55975, 16'd346, 16'd57382, 16'd27805, 16'd34942, 16'd50059, 16'd27844, 16'd59492, 16'd15209, 16'd41237, 16'd48044, 16'd58394, 16'd29856, 16'd9287, 16'd42956, 16'd65360, 16'd14425, 16'd4900, 16'd19379});
	test_expansion(128'h076c44a318fe3179dc99f09bc8a2af6c, {16'd11569, 16'd37238, 16'd65221, 16'd2036, 16'd54286, 16'd6396, 16'd47322, 16'd50213, 16'd44907, 16'd49829, 16'd52600, 16'd38926, 16'd22479, 16'd37605, 16'd10819, 16'd47258, 16'd12281, 16'd47570, 16'd22780, 16'd60972, 16'd46088, 16'd32767, 16'd59688, 16'd55143, 16'd24917, 16'd19715});
	test_expansion(128'h907e4970f3b0b0d4e075359a8b650332, {16'd28172, 16'd33276, 16'd6102, 16'd32318, 16'd28848, 16'd24791, 16'd54096, 16'd31701, 16'd46977, 16'd61861, 16'd42981, 16'd26079, 16'd1313, 16'd53589, 16'd20965, 16'd33823, 16'd46496, 16'd61970, 16'd5056, 16'd20861, 16'd43110, 16'd64414, 16'd41109, 16'd56573, 16'd59521, 16'd38855});
	test_expansion(128'hf2a5f7f416de689e9258ce372b6e9684, {16'd7182, 16'd42826, 16'd42415, 16'd4557, 16'd31493, 16'd44691, 16'd62696, 16'd33873, 16'd21516, 16'd16028, 16'd22592, 16'd51713, 16'd3442, 16'd40802, 16'd48014, 16'd3346, 16'd7100, 16'd1280, 16'd55669, 16'd41200, 16'd1901, 16'd43451, 16'd45587, 16'd43647, 16'd35395, 16'd8183});
	test_expansion(128'h922faa2bcc759540d570d24d79930263, {16'd30845, 16'd43563, 16'd56676, 16'd38093, 16'd28481, 16'd13237, 16'd55828, 16'd4636, 16'd9833, 16'd9707, 16'd23281, 16'd35865, 16'd6300, 16'd29311, 16'd27214, 16'd25654, 16'd35580, 16'd8291, 16'd21613, 16'd48233, 16'd60056, 16'd171, 16'd57386, 16'd599, 16'd21893, 16'd51600});
	test_expansion(128'h3bc647ec480ffc82b6930df95e3eea03, {16'd57980, 16'd4285, 16'd22423, 16'd37215, 16'd44411, 16'd49510, 16'd59095, 16'd19757, 16'd28571, 16'd64000, 16'd41743, 16'd13117, 16'd16953, 16'd15355, 16'd20839, 16'd999, 16'd21997, 16'd13311, 16'd36189, 16'd6864, 16'd24418, 16'd26485, 16'd34879, 16'd20238, 16'd58985, 16'd63513});
	test_expansion(128'h59f1529fc8a3d2a29f180b2ae8e215fb, {16'd56662, 16'd48576, 16'd21508, 16'd59370, 16'd7063, 16'd45563, 16'd42102, 16'd49100, 16'd58246, 16'd45926, 16'd43260, 16'd43302, 16'd27337, 16'd44451, 16'd6706, 16'd15475, 16'd2469, 16'd38841, 16'd13934, 16'd34059, 16'd39278, 16'd45266, 16'd892, 16'd2302, 16'd6128, 16'd4793});
	test_expansion(128'hc3427d964014e258ffbe59cdd142f181, {16'd29249, 16'd45987, 16'd21865, 16'd17692, 16'd19410, 16'd36856, 16'd38019, 16'd29820, 16'd34477, 16'd62570, 16'd42623, 16'd7970, 16'd32738, 16'd61573, 16'd27327, 16'd26520, 16'd5070, 16'd47537, 16'd17692, 16'd25919, 16'd16434, 16'd18967, 16'd5798, 16'd54898, 16'd53312, 16'd55047});
	test_expansion(128'h89a29391dd6296635688ecb5d0ed63d5, {16'd49306, 16'd64994, 16'd50321, 16'd4066, 16'd7877, 16'd39350, 16'd206, 16'd28659, 16'd10736, 16'd61643, 16'd43621, 16'd41102, 16'd18213, 16'd48820, 16'd41694, 16'd13435, 16'd8247, 16'd37973, 16'd24502, 16'd62219, 16'd42530, 16'd46503, 16'd64208, 16'd40689, 16'd2371, 16'd51123});
	test_expansion(128'h7b8a508860faf40420e0ade23c484854, {16'd11330, 16'd56533, 16'd12953, 16'd39091, 16'd51998, 16'd54120, 16'd58202, 16'd44845, 16'd7392, 16'd31409, 16'd61245, 16'd31712, 16'd47446, 16'd54766, 16'd21562, 16'd51313, 16'd16114, 16'd30890, 16'd48527, 16'd54909, 16'd17038, 16'd26136, 16'd29283, 16'd56198, 16'd63280, 16'd32434});
	test_expansion(128'h501759138a23ef6eec12c1e952ed750c, {16'd61317, 16'd23568, 16'd44856, 16'd27257, 16'd12592, 16'd12155, 16'd21596, 16'd2965, 16'd47797, 16'd19875, 16'd31245, 16'd59789, 16'd34009, 16'd17699, 16'd6370, 16'd4732, 16'd16837, 16'd59645, 16'd1084, 16'd45576, 16'd46904, 16'd60571, 16'd31549, 16'd20797, 16'd58856, 16'd47305});
	test_expansion(128'hbe8ddb1f2572695a36b7bd6c1bf0bfc8, {16'd61414, 16'd39678, 16'd52800, 16'd835, 16'd36846, 16'd35551, 16'd31553, 16'd57180, 16'd54196, 16'd46138, 16'd50739, 16'd36307, 16'd51438, 16'd56018, 16'd6996, 16'd26340, 16'd35141, 16'd28911, 16'd41642, 16'd12091, 16'd1692, 16'd28430, 16'd43763, 16'd6850, 16'd10219, 16'd18298});
	test_expansion(128'h1bb7388ea85b77b340a6b9235f864c3d, {16'd27323, 16'd49549, 16'd21782, 16'd63618, 16'd8441, 16'd21367, 16'd61005, 16'd19005, 16'd40297, 16'd33168, 16'd49443, 16'd35593, 16'd16979, 16'd12954, 16'd5902, 16'd46179, 16'd28738, 16'd15334, 16'd14848, 16'd25223, 16'd52049, 16'd55014, 16'd31874, 16'd10987, 16'd17721, 16'd31447});
	test_expansion(128'h3f523ccf5ef7cf2cb2b2ca20c2070d82, {16'd59772, 16'd51554, 16'd12319, 16'd21555, 16'd1499, 16'd4611, 16'd58699, 16'd16248, 16'd48713, 16'd56039, 16'd47259, 16'd8243, 16'd52780, 16'd671, 16'd59887, 16'd43288, 16'd39389, 16'd62073, 16'd63842, 16'd51302, 16'd9107, 16'd21539, 16'd8105, 16'd26958, 16'd56741, 16'd17724});
	test_expansion(128'h23b189fec07ad420b906c15401db7bcd, {16'd36790, 16'd11820, 16'd30677, 16'd11763, 16'd56633, 16'd32515, 16'd36084, 16'd23980, 16'd3991, 16'd50723, 16'd37222, 16'd13677, 16'd61991, 16'd61811, 16'd16456, 16'd11822, 16'd10657, 16'd26977, 16'd46401, 16'd36875, 16'd22854, 16'd32868, 16'd48454, 16'd51553, 16'd29476, 16'd33667});
	test_expansion(128'h5b5df9cfc5d486f9742eafa8fcc0df2f, {16'd14281, 16'd40904, 16'd13826, 16'd8731, 16'd55313, 16'd46627, 16'd57001, 16'd26490, 16'd31464, 16'd59017, 16'd31016, 16'd44825, 16'd30111, 16'd8849, 16'd56733, 16'd38175, 16'd15124, 16'd42975, 16'd17913, 16'd19275, 16'd40830, 16'd55056, 16'd26637, 16'd8068, 16'd18583, 16'd59170});
	test_expansion(128'h044c56e2a2afdbd490eca36674b2b710, {16'd6729, 16'd6723, 16'd41073, 16'd42846, 16'd9277, 16'd9626, 16'd27717, 16'd29172, 16'd15538, 16'd35928, 16'd3204, 16'd43694, 16'd26427, 16'd64714, 16'd11756, 16'd64372, 16'd35140, 16'd37564, 16'd23978, 16'd42547, 16'd47950, 16'd21491, 16'd45261, 16'd50578, 16'd59062, 16'd48798});
	test_expansion(128'h2d2e4523a5d2ac1f8d0bce7fd2758e3a, {16'd14209, 16'd3691, 16'd50, 16'd19566, 16'd28951, 16'd43112, 16'd7123, 16'd41482, 16'd3735, 16'd12454, 16'd41574, 16'd22703, 16'd32920, 16'd6986, 16'd50703, 16'd44191, 16'd45925, 16'd499, 16'd20541, 16'd59428, 16'd16057, 16'd14948, 16'd12363, 16'd28237, 16'd35388, 16'd22828});
	test_expansion(128'ha51402095ca8afc3480dba0bdc42ae99, {16'd47713, 16'd48699, 16'd7520, 16'd8030, 16'd31915, 16'd17690, 16'd63762, 16'd4414, 16'd30723, 16'd42436, 16'd4536, 16'd8235, 16'd49862, 16'd35244, 16'd64278, 16'd60396, 16'd22480, 16'd50017, 16'd677, 16'd48971, 16'd39744, 16'd18322, 16'd38539, 16'd62235, 16'd14599, 16'd22687});
	test_expansion(128'h2107284cb8ce1d59ec0befba3cb38cf0, {16'd61210, 16'd3283, 16'd42139, 16'd44755, 16'd7635, 16'd63355, 16'd12983, 16'd35767, 16'd23079, 16'd64664, 16'd34361, 16'd34325, 16'd40956, 16'd25045, 16'd23226, 16'd64278, 16'd18976, 16'd42352, 16'd7160, 16'd48738, 16'd458, 16'd45109, 16'd61572, 16'd54082, 16'd64177, 16'd19008});
	test_expansion(128'h88b67485bb03ebc8c25d97d9d02a9461, {16'd28714, 16'd34487, 16'd1082, 16'd54882, 16'd1692, 16'd19358, 16'd37095, 16'd3724, 16'd40935, 16'd46690, 16'd595, 16'd31738, 16'd46391, 16'd64346, 16'd48480, 16'd43495, 16'd48782, 16'd27418, 16'd38046, 16'd41890, 16'd48375, 16'd19174, 16'd29270, 16'd48056, 16'd51299, 16'd58445});
	test_expansion(128'hb82f8ef93b8e246e6fff65dbc3cf4334, {16'd37668, 16'd8099, 16'd39625, 16'd27021, 16'd64019, 16'd47960, 16'd7257, 16'd61031, 16'd51005, 16'd58392, 16'd63816, 16'd58114, 16'd44165, 16'd50102, 16'd63789, 16'd52617, 16'd41707, 16'd58533, 16'd4215, 16'd2291, 16'd64429, 16'd44942, 16'd22246, 16'd4787, 16'd55499, 16'd35891});
	test_expansion(128'he0f110e41451e84bad127bf2cf40e27d, {16'd45417, 16'd4143, 16'd33485, 16'd58799, 16'd32057, 16'd37642, 16'd54735, 16'd26267, 16'd62749, 16'd35213, 16'd14368, 16'd1002, 16'd37892, 16'd4388, 16'd27494, 16'd58277, 16'd27523, 16'd12554, 16'd31648, 16'd54026, 16'd19601, 16'd11311, 16'd19600, 16'd61481, 16'd12975, 16'd42935});
	test_expansion(128'h233d47d6cbae832b2629529a2087e0db, {16'd20230, 16'd10791, 16'd45009, 16'd26701, 16'd47128, 16'd20455, 16'd50709, 16'd12400, 16'd42725, 16'd4209, 16'd30604, 16'd51901, 16'd44933, 16'd54615, 16'd34638, 16'd34450, 16'd33670, 16'd61126, 16'd37134, 16'd20971, 16'd21605, 16'd63571, 16'd43578, 16'd35783, 16'd58729, 16'd11141});
	test_expansion(128'h6a1a6a54a9bdb2488a2f2280afef7655, {16'd25435, 16'd3568, 16'd11281, 16'd48653, 16'd37341, 16'd58998, 16'd35294, 16'd34173, 16'd43815, 16'd11131, 16'd52189, 16'd9927, 16'd18867, 16'd54138, 16'd28335, 16'd65299, 16'd27501, 16'd40785, 16'd40165, 16'd51738, 16'd26961, 16'd29579, 16'd38410, 16'd2234, 16'd57081, 16'd57446});
	test_expansion(128'h9ae74b3ea1573185289c4cc8322bd14b, {16'd41566, 16'd3838, 16'd46210, 16'd64661, 16'd562, 16'd29317, 16'd42058, 16'd46707, 16'd38564, 16'd21281, 16'd34669, 16'd24333, 16'd62941, 16'd45585, 16'd57117, 16'd24943, 16'd32710, 16'd21284, 16'd53391, 16'd63090, 16'd25073, 16'd21860, 16'd11016, 16'd49225, 16'd10446, 16'd63207});
	test_expansion(128'h702343b409b45fceeca55d03deb1d788, {16'd32009, 16'd8630, 16'd38746, 16'd7809, 16'd28272, 16'd52610, 16'd47467, 16'd10068, 16'd52745, 16'd22596, 16'd6304, 16'd28969, 16'd39800, 16'd12994, 16'd16177, 16'd12461, 16'd45981, 16'd49616, 16'd15201, 16'd55457, 16'd5303, 16'd46613, 16'd38895, 16'd34755, 16'd52350, 16'd24086});
	test_expansion(128'hf9f4d6ad67d0ab84a750392aeab15934, {16'd6283, 16'd42985, 16'd14516, 16'd10853, 16'd8138, 16'd9057, 16'd25582, 16'd63279, 16'd20370, 16'd38328, 16'd18810, 16'd5231, 16'd37871, 16'd21345, 16'd30690, 16'd15052, 16'd31326, 16'd5938, 16'd19440, 16'd46296, 16'd23247, 16'd25253, 16'd37722, 16'd12481, 16'd3947, 16'd30862});
	test_expansion(128'h4282659d89223c3fd46469e1ca38a692, {16'd55912, 16'd3436, 16'd61550, 16'd57007, 16'd29606, 16'd53593, 16'd14366, 16'd3136, 16'd35412, 16'd38258, 16'd25577, 16'd27037, 16'd42246, 16'd18686, 16'd62941, 16'd32267, 16'd34044, 16'd16082, 16'd51554, 16'd23431, 16'd26204, 16'd38456, 16'd1492, 16'd39471, 16'd54600, 16'd37806});
	test_expansion(128'h395733b5ff255624fbe26ef734c6bc08, {16'd3569, 16'd9670, 16'd61504, 16'd33782, 16'd57070, 16'd30137, 16'd16505, 16'd9839, 16'd8926, 16'd33586, 16'd55826, 16'd29608, 16'd51028, 16'd19933, 16'd48076, 16'd34063, 16'd30909, 16'd27218, 16'd59118, 16'd5700, 16'd40768, 16'd51878, 16'd22065, 16'd14134, 16'd32083, 16'd51280});
	test_expansion(128'h5fef6b5db4f73e475c223103943fea7f, {16'd57632, 16'd22113, 16'd28497, 16'd43200, 16'd11070, 16'd6795, 16'd53518, 16'd4450, 16'd42085, 16'd11538, 16'd26512, 16'd6450, 16'd49895, 16'd25450, 16'd46719, 16'd47945, 16'd8724, 16'd51206, 16'd2519, 16'd21957, 16'd57641, 16'd46757, 16'd2497, 16'd39358, 16'd31758, 16'd44359});
	test_expansion(128'h08ef6188ba30ea95a2b9fcd8ceccf9a4, {16'd58253, 16'd34659, 16'd18252, 16'd2163, 16'd31458, 16'd20743, 16'd45877, 16'd19266, 16'd10170, 16'd3365, 16'd14159, 16'd57434, 16'd53813, 16'd14527, 16'd28389, 16'd35613, 16'd23345, 16'd27117, 16'd37473, 16'd1803, 16'd2454, 16'd2776, 16'd1262, 16'd53646, 16'd6402, 16'd5194});
	test_expansion(128'h70fe3bf8a0ef2e1694e965bae5e00fcf, {16'd16063, 16'd8223, 16'd15453, 16'd26373, 16'd28057, 16'd46819, 16'd40155, 16'd58507, 16'd36894, 16'd58135, 16'd46533, 16'd5568, 16'd54706, 16'd53445, 16'd35532, 16'd1877, 16'd8550, 16'd35958, 16'd52618, 16'd36325, 16'd28729, 16'd30428, 16'd27915, 16'd42730, 16'd61733, 16'd31513});
	test_expansion(128'h9a62e778d21d8d79612b903717b99b3f, {16'd31384, 16'd32424, 16'd40976, 16'd35291, 16'd65077, 16'd39403, 16'd35123, 16'd32458, 16'd44535, 16'd12962, 16'd19201, 16'd24766, 16'd40402, 16'd25869, 16'd65122, 16'd53795, 16'd33518, 16'd2245, 16'd24688, 16'd53450, 16'd5888, 16'd4525, 16'd14613, 16'd48573, 16'd36149, 16'd37535});
	test_expansion(128'hfbbfa8aaadc5e299f61e69321a456caf, {16'd42329, 16'd30230, 16'd1939, 16'd17667, 16'd31041, 16'd55749, 16'd50564, 16'd3419, 16'd62648, 16'd24848, 16'd5709, 16'd8441, 16'd3528, 16'd29439, 16'd45387, 16'd50882, 16'd49085, 16'd61584, 16'd63306, 16'd6104, 16'd52125, 16'd43472, 16'd56715, 16'd49560, 16'd18315, 16'd3515});
	test_expansion(128'hfc2d18fb95d8d07b3089c3a52f172015, {16'd1253, 16'd33370, 16'd39449, 16'd55036, 16'd25971, 16'd58909, 16'd42338, 16'd28060, 16'd4905, 16'd60689, 16'd14049, 16'd55197, 16'd29713, 16'd3451, 16'd17597, 16'd29197, 16'd19017, 16'd1924, 16'd17913, 16'd14818, 16'd56191, 16'd42203, 16'd1746, 16'd19003, 16'd56420, 16'd57123});
	test_expansion(128'h34fc728aa85f27a2638e7f78cdef51d2, {16'd22377, 16'd11554, 16'd55610, 16'd16124, 16'd37442, 16'd27577, 16'd56080, 16'd50249, 16'd29933, 16'd6017, 16'd56272, 16'd54791, 16'd58587, 16'd47417, 16'd65109, 16'd4989, 16'd54326, 16'd23380, 16'd6547, 16'd62652, 16'd37461, 16'd51223, 16'd54482, 16'd47314, 16'd2587, 16'd64310});
	test_expansion(128'h28e1da8e32b29409c3cb650341ec0c20, {16'd14935, 16'd9048, 16'd39011, 16'd62216, 16'd16245, 16'd52643, 16'd40639, 16'd50548, 16'd49666, 16'd12032, 16'd36309, 16'd55545, 16'd46243, 16'd13196, 16'd27336, 16'd23254, 16'd43172, 16'd63966, 16'd31224, 16'd61506, 16'd62040, 16'd19881, 16'd10441, 16'd2700, 16'd32444, 16'd64477});
	test_expansion(128'h566ec4ab61d3a47fed21562c961277a9, {16'd47678, 16'd38010, 16'd55831, 16'd10396, 16'd8443, 16'd52456, 16'd27220, 16'd3895, 16'd11872, 16'd23862, 16'd6919, 16'd24498, 16'd51436, 16'd45922, 16'd27869, 16'd16953, 16'd17005, 16'd16053, 16'd2351, 16'd23097, 16'd48319, 16'd47165, 16'd27943, 16'd20262, 16'd7393, 16'd53919});
	test_expansion(128'h346a364ec8e56f4f9d897d71a34371d2, {16'd33078, 16'd21739, 16'd48701, 16'd55085, 16'd20929, 16'd795, 16'd50839, 16'd35878, 16'd29006, 16'd49116, 16'd39515, 16'd55995, 16'd63691, 16'd42108, 16'd26050, 16'd46466, 16'd19313, 16'd60037, 16'd51238, 16'd4304, 16'd12978, 16'd26247, 16'd38775, 16'd58006, 16'd40187, 16'd38597});
	test_expansion(128'hf61d2a73490f56c3c66cc2eef5152977, {16'd40357, 16'd35240, 16'd13275, 16'd24919, 16'd47380, 16'd55480, 16'd61812, 16'd58136, 16'd17746, 16'd8044, 16'd64944, 16'd44229, 16'd46276, 16'd39780, 16'd6101, 16'd11943, 16'd22654, 16'd53200, 16'd61581, 16'd1957, 16'd65348, 16'd44051, 16'd54085, 16'd50611, 16'd7800, 16'd32300});
	test_expansion(128'h3474d1375f157827140dc2e30732fb83, {16'd43719, 16'd1200, 16'd2485, 16'd23094, 16'd5632, 16'd391, 16'd12711, 16'd48709, 16'd23775, 16'd14571, 16'd25149, 16'd38035, 16'd1272, 16'd38633, 16'd15513, 16'd33830, 16'd13601, 16'd27688, 16'd61085, 16'd54712, 16'd23803, 16'd13914, 16'd34009, 16'd29807, 16'd60752, 16'd4647});
	test_expansion(128'h3438f557e0d5ba6e74e66a86b89e3609, {16'd35841, 16'd9290, 16'd35681, 16'd52509, 16'd46934, 16'd56796, 16'd50518, 16'd22155, 16'd31309, 16'd40600, 16'd41253, 16'd26527, 16'd46500, 16'd35845, 16'd32909, 16'd56372, 16'd22147, 16'd7303, 16'd33016, 16'd42931, 16'd36306, 16'd2074, 16'd37839, 16'd5347, 16'd59346, 16'd8447});
	test_expansion(128'hbcc7cc74e226909ca98fbb79b6c4e26e, {16'd10872, 16'd12670, 16'd1491, 16'd39431, 16'd28948, 16'd19070, 16'd2449, 16'd6999, 16'd52160, 16'd28229, 16'd43204, 16'd17014, 16'd5127, 16'd18304, 16'd44636, 16'd55790, 16'd62463, 16'd35527, 16'd53815, 16'd33218, 16'd7513, 16'd25317, 16'd50190, 16'd39059, 16'd42171, 16'd15617});
	test_expansion(128'had3776252b84d61c6902f2e01e252e27, {16'd20859, 16'd30736, 16'd60220, 16'd7571, 16'd23490, 16'd20701, 16'd15052, 16'd31515, 16'd32513, 16'd62017, 16'd20865, 16'd23214, 16'd25172, 16'd17237, 16'd7850, 16'd23074, 16'd65042, 16'd32954, 16'd2655, 16'd4987, 16'd23842, 16'd30164, 16'd52598, 16'd53080, 16'd34574, 16'd25220});
	test_expansion(128'h0534c779c55a803ef029fea2b5f3b233, {16'd61291, 16'd42448, 16'd2813, 16'd26227, 16'd19008, 16'd62447, 16'd1328, 16'd12569, 16'd21114, 16'd60730, 16'd2922, 16'd11320, 16'd20566, 16'd11543, 16'd41618, 16'd10704, 16'd24278, 16'd18719, 16'd58392, 16'd22853, 16'd36755, 16'd11442, 16'd46853, 16'd18535, 16'd43596, 16'd9088});
	test_expansion(128'h3d5006a4db2f750c25b6145e532f196c, {16'd57337, 16'd50283, 16'd18030, 16'd43707, 16'd52975, 16'd27857, 16'd20485, 16'd41611, 16'd14473, 16'd33661, 16'd56391, 16'd28399, 16'd24025, 16'd48752, 16'd32974, 16'd64282, 16'd45884, 16'd65287, 16'd20957, 16'd50913, 16'd55189, 16'd40297, 16'd64039, 16'd12631, 16'd29782, 16'd57849});
	test_expansion(128'h6a6d802f2dcfb76ad0471b1347472a1a, {16'd5844, 16'd48307, 16'd41269, 16'd27064, 16'd23879, 16'd25628, 16'd57167, 16'd26326, 16'd16093, 16'd14902, 16'd13614, 16'd28005, 16'd29540, 16'd26021, 16'd26764, 16'd52671, 16'd46002, 16'd62957, 16'd58546, 16'd38967, 16'd32940, 16'd16118, 16'd13882, 16'd17707, 16'd15388, 16'd35863});
	test_expansion(128'h7134b8c5f572a8eb746b671fd71d1808, {16'd22873, 16'd32620, 16'd50831, 16'd15992, 16'd12496, 16'd22791, 16'd32845, 16'd57178, 16'd25365, 16'd25658, 16'd7490, 16'd24947, 16'd56965, 16'd32309, 16'd27145, 16'd54676, 16'd51114, 16'd56290, 16'd34227, 16'd59460, 16'd57448, 16'd31910, 16'd19330, 16'd62426, 16'd16261, 16'd31558});
	test_expansion(128'h8c5d0dd8474e731892319547f1a4029f, {16'd13345, 16'd2498, 16'd30026, 16'd12693, 16'd38734, 16'd42053, 16'd10638, 16'd47329, 16'd63182, 16'd49444, 16'd65037, 16'd8493, 16'd59264, 16'd20762, 16'd19587, 16'd42650, 16'd14430, 16'd56326, 16'd38581, 16'd65021, 16'd41973, 16'd46435, 16'd17479, 16'd5028, 16'd48097, 16'd34502});
	test_expansion(128'h34cab673655fe1a7085ea4882b40b1aa, {16'd3192, 16'd19249, 16'd2929, 16'd52083, 16'd23575, 16'd5221, 16'd58116, 16'd30638, 16'd38117, 16'd61758, 16'd63568, 16'd49765, 16'd23835, 16'd41972, 16'd3895, 16'd12642, 16'd47074, 16'd41619, 16'd25256, 16'd37537, 16'd7671, 16'd49665, 16'd29769, 16'd44262, 16'd50830, 16'd603});
	test_expansion(128'h783c9debd85461b871a4abe8178adfec, {16'd30716, 16'd56008, 16'd5177, 16'd46178, 16'd51531, 16'd61760, 16'd16618, 16'd10764, 16'd54784, 16'd46292, 16'd12220, 16'd33655, 16'd39999, 16'd39436, 16'd11328, 16'd40572, 16'd62369, 16'd39649, 16'd18123, 16'd17289, 16'd2477, 16'd27185, 16'd8467, 16'd24947, 16'd54139, 16'd14458});
	test_expansion(128'h8174445bf30acae11e3879fa77953c73, {16'd1713, 16'd15080, 16'd55995, 16'd32247, 16'd62046, 16'd678, 16'd55114, 16'd23908, 16'd11406, 16'd24128, 16'd62012, 16'd25826, 16'd54801, 16'd16059, 16'd16712, 16'd48799, 16'd53775, 16'd41683, 16'd64713, 16'd35334, 16'd39181, 16'd62123, 16'd30738, 16'd60506, 16'd22239, 16'd34504});
	test_expansion(128'h76cb65c1606e7d468ec4d688b324eb03, {16'd59874, 16'd12027, 16'd31713, 16'd32381, 16'd56812, 16'd24586, 16'd20964, 16'd64735, 16'd54544, 16'd34922, 16'd40436, 16'd58869, 16'd18540, 16'd52660, 16'd4449, 16'd51441, 16'd6275, 16'd20325, 16'd58509, 16'd55677, 16'd34976, 16'd33482, 16'd30037, 16'd26455, 16'd40250, 16'd28250});
	test_expansion(128'h48fb61b33996c1c127f0ceace108d200, {16'd10429, 16'd2853, 16'd39245, 16'd10633, 16'd10402, 16'd62201, 16'd22775, 16'd14901, 16'd2376, 16'd4700, 16'd37218, 16'd52233, 16'd20571, 16'd41602, 16'd40367, 16'd52211, 16'd26189, 16'd39685, 16'd27996, 16'd5378, 16'd37073, 16'd10633, 16'd17521, 16'd31408, 16'd10116, 16'd62726});
	test_expansion(128'h06d303910c1445e31013807d3d48baab, {16'd33239, 16'd64724, 16'd53760, 16'd39551, 16'd38894, 16'd19724, 16'd51407, 16'd32848, 16'd31610, 16'd46766, 16'd44982, 16'd3973, 16'd50495, 16'd42429, 16'd15939, 16'd44331, 16'd56212, 16'd24945, 16'd63264, 16'd16279, 16'd47513, 16'd14731, 16'd8568, 16'd63116, 16'd61735, 16'd31973});
	test_expansion(128'hbd69a00498a954e980b5c16d3427433e, {16'd40571, 16'd7412, 16'd45735, 16'd33150, 16'd16058, 16'd56534, 16'd33860, 16'd23221, 16'd7151, 16'd34690, 16'd51255, 16'd19647, 16'd10202, 16'd22832, 16'd4400, 16'd44971, 16'd52826, 16'd7762, 16'd57735, 16'd11389, 16'd14978, 16'd19095, 16'd15854, 16'd16299, 16'd35201, 16'd62545});
	test_expansion(128'h0c60b406448863807e74eba64e88b459, {16'd30653, 16'd24441, 16'd24885, 16'd19739, 16'd14650, 16'd452, 16'd42836, 16'd60201, 16'd45654, 16'd47054, 16'd50834, 16'd6467, 16'd7667, 16'd45459, 16'd21975, 16'd48348, 16'd45710, 16'd53271, 16'd49496, 16'd4650, 16'd62068, 16'd59321, 16'd53648, 16'd33471, 16'd46458, 16'd5267});
	test_expansion(128'h05a59dc0e8e5ee565538bc07332aed00, {16'd39360, 16'd23756, 16'd16072, 16'd54624, 16'd54203, 16'd41270, 16'd41161, 16'd17485, 16'd30857, 16'd16674, 16'd23033, 16'd30205, 16'd40843, 16'd61810, 16'd59438, 16'd57812, 16'd55440, 16'd51889, 16'd7445, 16'd13348, 16'd38401, 16'd3014, 16'd8349, 16'd60718, 16'd38279, 16'd15558});
	test_expansion(128'hc6e649aba2819cc5b246ca9e6dab93e9, {16'd36722, 16'd51336, 16'd31012, 16'd32497, 16'd32903, 16'd29985, 16'd51569, 16'd15165, 16'd10055, 16'd17842, 16'd47056, 16'd13194, 16'd23439, 16'd51030, 16'd49187, 16'd4821, 16'd27467, 16'd25128, 16'd763, 16'd11157, 16'd3513, 16'd47603, 16'd8133, 16'd7655, 16'd37051, 16'd27273});
	test_expansion(128'h416d7d9f83f58acc448b2273f380eec7, {16'd27113, 16'd24639, 16'd51488, 16'd63561, 16'd54173, 16'd14863, 16'd44004, 16'd47961, 16'd41127, 16'd41825, 16'd14502, 16'd15363, 16'd16428, 16'd18827, 16'd4445, 16'd34203, 16'd20541, 16'd55132, 16'd3690, 16'd9541, 16'd11002, 16'd6930, 16'd38719, 16'd39699, 16'd22152, 16'd28853});
	test_expansion(128'h11022ba8a78fb0908b78a4300cd77dac, {16'd22698, 16'd32907, 16'd27146, 16'd61478, 16'd64225, 16'd54900, 16'd50541, 16'd41894, 16'd61435, 16'd55449, 16'd21954, 16'd39847, 16'd24311, 16'd25880, 16'd20518, 16'd32158, 16'd32946, 16'd46484, 16'd27524, 16'd4172, 16'd1449, 16'd21331, 16'd42169, 16'd26357, 16'd51318, 16'd53002});
	test_expansion(128'h87815ee41b9f14e682476bd715c8b386, {16'd51746, 16'd33696, 16'd40654, 16'd60005, 16'd36847, 16'd21430, 16'd64514, 16'd15030, 16'd28295, 16'd7513, 16'd31986, 16'd18525, 16'd27051, 16'd42813, 16'd29087, 16'd60817, 16'd16946, 16'd63034, 16'd49610, 16'd16396, 16'd922, 16'd27072, 16'd17592, 16'd43647, 16'd36239, 16'd5638});
	test_expansion(128'h1d0dc79e8f6fd73197e71013abe1d0b3, {16'd19154, 16'd2741, 16'd29756, 16'd61045, 16'd65342, 16'd21835, 16'd57331, 16'd33326, 16'd45884, 16'd49646, 16'd14449, 16'd12669, 16'd6196, 16'd22053, 16'd53082, 16'd34155, 16'd15111, 16'd24395, 16'd56825, 16'd42840, 16'd6004, 16'd39521, 16'd19081, 16'd36324, 16'd10532, 16'd48246});
	test_expansion(128'h6334fe9f7567a14f63af11e138a4638d, {16'd38716, 16'd34175, 16'd6575, 16'd65255, 16'd56255, 16'd30514, 16'd54907, 16'd35563, 16'd35138, 16'd41274, 16'd13648, 16'd38949, 16'd59843, 16'd52728, 16'd59035, 16'd3949, 16'd60464, 16'd24340, 16'd33173, 16'd41057, 16'd44048, 16'd57965, 16'd8574, 16'd40675, 16'd61644, 16'd49523});
	test_expansion(128'he794e095e8a46f11baafda3afe038cea, {16'd19124, 16'd30038, 16'd54918, 16'd25045, 16'd4907, 16'd3200, 16'd56508, 16'd27223, 16'd34009, 16'd18183, 16'd37175, 16'd60625, 16'd56034, 16'd39862, 16'd55267, 16'd35471, 16'd18110, 16'd46702, 16'd15397, 16'd54150, 16'd26724, 16'd58141, 16'd52093, 16'd38938, 16'd28694, 16'd13230});
	test_expansion(128'h9230c050462d83ea560542fda867af83, {16'd39970, 16'd205, 16'd12201, 16'd16963, 16'd2947, 16'd53528, 16'd64718, 16'd15115, 16'd40342, 16'd29871, 16'd47439, 16'd45905, 16'd2710, 16'd45713, 16'd43941, 16'd50004, 16'd3329, 16'd20824, 16'd52040, 16'd5011, 16'd20308, 16'd52033, 16'd34684, 16'd47599, 16'd10907, 16'd27825});
	test_expansion(128'hbc951452a0af51f8425ff0af6da5e41c, {16'd64879, 16'd18153, 16'd8302, 16'd35530, 16'd30857, 16'd52313, 16'd4880, 16'd17388, 16'd42648, 16'd43685, 16'd37574, 16'd18368, 16'd61368, 16'd52439, 16'd11453, 16'd41739, 16'd42706, 16'd51197, 16'd17687, 16'd16580, 16'd40656, 16'd25064, 16'd27326, 16'd31916, 16'd936, 16'd17228});
	test_expansion(128'h31139e678f6624ae99c90bdd06344a40, {16'd27986, 16'd5265, 16'd26579, 16'd14577, 16'd50343, 16'd4441, 16'd37790, 16'd51946, 16'd54947, 16'd52907, 16'd31168, 16'd32594, 16'd64039, 16'd5062, 16'd47909, 16'd19646, 16'd64307, 16'd41821, 16'd55752, 16'd28954, 16'd22485, 16'd360, 16'd41099, 16'd4718, 16'd12428, 16'd5464});
	test_expansion(128'h10c124b3c3b8bb3fa0cecb91164325ef, {16'd40647, 16'd24924, 16'd65460, 16'd2681, 16'd56249, 16'd30542, 16'd47835, 16'd59751, 16'd20022, 16'd57298, 16'd39859, 16'd64592, 16'd19906, 16'd14146, 16'd18488, 16'd37271, 16'd22461, 16'd48921, 16'd47208, 16'd30127, 16'd57631, 16'd46296, 16'd43608, 16'd2088, 16'd7332, 16'd46374});
	test_expansion(128'h0561289a311ebf95ff577475b7d70cfa, {16'd50538, 16'd43525, 16'd11502, 16'd55686, 16'd44220, 16'd54541, 16'd14288, 16'd25794, 16'd26591, 16'd48775, 16'd58072, 16'd59562, 16'd34944, 16'd61852, 16'd55748, 16'd35135, 16'd40182, 16'd48724, 16'd15788, 16'd17884, 16'd31329, 16'd31968, 16'd63563, 16'd25316, 16'd34893, 16'd7646});
	test_expansion(128'h6c142c061b948a4551b379855e8638d0, {16'd24791, 16'd36412, 16'd59688, 16'd53783, 16'd4322, 16'd45274, 16'd23311, 16'd5812, 16'd34220, 16'd57108, 16'd61494, 16'd42694, 16'd61853, 16'd26648, 16'd15779, 16'd8020, 16'd47100, 16'd56431, 16'd26164, 16'd31361, 16'd19686, 16'd19347, 16'd45798, 16'd35142, 16'd61032, 16'd64299});
	test_expansion(128'hb002e0d6cea9d7ff6b1712b09fc9e4ba, {16'd9446, 16'd23726, 16'd64851, 16'd21403, 16'd4113, 16'd20103, 16'd59552, 16'd27186, 16'd34842, 16'd39124, 16'd58837, 16'd40249, 16'd18196, 16'd22756, 16'd38913, 16'd52755, 16'd3549, 16'd64933, 16'd42138, 16'd16897, 16'd25557, 16'd13030, 16'd53253, 16'd7461, 16'd2249, 16'd24282});
	test_expansion(128'hf07af7ab98de0f6a47a100b0058224f7, {16'd27044, 16'd47138, 16'd53260, 16'd21689, 16'd58675, 16'd7107, 16'd51773, 16'd59218, 16'd48373, 16'd32556, 16'd12195, 16'd12276, 16'd48739, 16'd28283, 16'd58624, 16'd2562, 16'd50296, 16'd7683, 16'd62286, 16'd54433, 16'd34286, 16'd42091, 16'd29672, 16'd16732, 16'd18537, 16'd20487});
	test_expansion(128'ha5c63c41731e2d97cfb8a13369c79542, {16'd37165, 16'd48999, 16'd51716, 16'd14799, 16'd52142, 16'd47873, 16'd32364, 16'd58669, 16'd59478, 16'd61805, 16'd23056, 16'd51811, 16'd354, 16'd62878, 16'd5068, 16'd65230, 16'd4691, 16'd58038, 16'd36886, 16'd55940, 16'd21925, 16'd54036, 16'd33016, 16'd30515, 16'd63015, 16'd58622});
	test_expansion(128'ha9bf703782f90ca5d7de6369bc51d126, {16'd9997, 16'd19790, 16'd43457, 16'd33152, 16'd18212, 16'd38273, 16'd9302, 16'd3539, 16'd37905, 16'd43123, 16'd23761, 16'd17219, 16'd16143, 16'd62488, 16'd2516, 16'd49587, 16'd57181, 16'd55011, 16'd31182, 16'd42186, 16'd54383, 16'd31966, 16'd60521, 16'd25623, 16'd40543, 16'd11028});
	test_expansion(128'h3bbd22fa4ecaea21045fbe8f4035470a, {16'd33459, 16'd47345, 16'd31949, 16'd63317, 16'd2800, 16'd37638, 16'd10692, 16'd34537, 16'd47486, 16'd29853, 16'd54460, 16'd25359, 16'd9320, 16'd30291, 16'd34451, 16'd10561, 16'd30218, 16'd36251, 16'd43836, 16'd60316, 16'd49906, 16'd27108, 16'd34756, 16'd46168, 16'd40671, 16'd5980});
	test_expansion(128'h71cb189ac2b16b059db452c774a4809a, {16'd63429, 16'd48442, 16'd25362, 16'd25580, 16'd64334, 16'd45586, 16'd55738, 16'd51032, 16'd31694, 16'd35895, 16'd56154, 16'd14093, 16'd30157, 16'd63195, 16'd34824, 16'd20018, 16'd37795, 16'd9192, 16'd28418, 16'd61186, 16'd3999, 16'd15894, 16'd18489, 16'd52120, 16'd29579, 16'd12509});
	test_expansion(128'h4c3e8ebbe6bd14131e877056666d097e, {16'd5538, 16'd6537, 16'd19298, 16'd52649, 16'd5351, 16'd53229, 16'd49767, 16'd20429, 16'd38480, 16'd36681, 16'd1776, 16'd13934, 16'd38851, 16'd55324, 16'd22657, 16'd43372, 16'd11360, 16'd7524, 16'd26935, 16'd43875, 16'd52480, 16'd22574, 16'd24963, 16'd46939, 16'd39471, 16'd31265});
	test_expansion(128'hc69e83da502467e566b47db7f423dbd7, {16'd43164, 16'd39978, 16'd7276, 16'd48361, 16'd43308, 16'd5235, 16'd55064, 16'd29412, 16'd53747, 16'd56811, 16'd51150, 16'd32990, 16'd55755, 16'd22978, 16'd48615, 16'd34580, 16'd45383, 16'd44018, 16'd10734, 16'd24985, 16'd29099, 16'd41865, 16'd20255, 16'd22701, 16'd41553, 16'd3360});
	test_expansion(128'hb0751e0029e4691d802d88eee44a8749, {16'd63060, 16'd60815, 16'd39854, 16'd37428, 16'd42132, 16'd65279, 16'd47945, 16'd42806, 16'd11877, 16'd39013, 16'd9879, 16'd57980, 16'd21278, 16'd39947, 16'd36614, 16'd8927, 16'd55375, 16'd58651, 16'd31859, 16'd3854, 16'd6826, 16'd15243, 16'd35652, 16'd15833, 16'd20231, 16'd8043});
	test_expansion(128'h3af9ed7a8463c3b6211d4ca24ab5a583, {16'd34980, 16'd2079, 16'd44061, 16'd26277, 16'd56703, 16'd8594, 16'd9803, 16'd36758, 16'd44776, 16'd38023, 16'd10804, 16'd58146, 16'd31183, 16'd29843, 16'd32399, 16'd21995, 16'd64634, 16'd26946, 16'd14313, 16'd42134, 16'd19667, 16'd47531, 16'd42177, 16'd54345, 16'd19855, 16'd31979});
	test_expansion(128'h950d4f0df2d9045c62f63e36537d4bda, {16'd37477, 16'd2109, 16'd61108, 16'd65360, 16'd28535, 16'd47433, 16'd18138, 16'd30772, 16'd42857, 16'd14002, 16'd23884, 16'd20847, 16'd27097, 16'd42477, 16'd41738, 16'd19484, 16'd27570, 16'd52049, 16'd49424, 16'd17912, 16'd62360, 16'd32275, 16'd7376, 16'd26506, 16'd13739, 16'd11627});
	test_expansion(128'h68f94e8cf5684e6933e92a042e36cdbb, {16'd12749, 16'd13640, 16'd14773, 16'd35914, 16'd63120, 16'd33247, 16'd23335, 16'd55226, 16'd23012, 16'd21546, 16'd61478, 16'd21485, 16'd5605, 16'd17839, 16'd6946, 16'd56477, 16'd50992, 16'd41141, 16'd51162, 16'd12540, 16'd16966, 16'd29216, 16'd56522, 16'd59029, 16'd27667, 16'd14645});
	test_expansion(128'h6fc4ee844f01cf54c83a3689c8ecf280, {16'd18117, 16'd13114, 16'd54783, 16'd53286, 16'd19056, 16'd12514, 16'd41734, 16'd4168, 16'd20298, 16'd28022, 16'd20003, 16'd59685, 16'd18537, 16'd62348, 16'd31455, 16'd22206, 16'd21294, 16'd15690, 16'd44109, 16'd62246, 16'd6498, 16'd63087, 16'd12654, 16'd46828, 16'd3214, 16'd1162});
	test_expansion(128'h0f076b8c6ac4885686ef3c5c07107312, {16'd24472, 16'd4910, 16'd42328, 16'd59579, 16'd39225, 16'd32566, 16'd60045, 16'd7516, 16'd23777, 16'd38066, 16'd51554, 16'd56899, 16'd65520, 16'd55805, 16'd50485, 16'd22400, 16'd4906, 16'd2709, 16'd50228, 16'd9805, 16'd23059, 16'd35439, 16'd50403, 16'd14600, 16'd3068, 16'd36214});
	test_expansion(128'h3b981e965d2fba0427e132565ca0bd31, {16'd39795, 16'd36250, 16'd58437, 16'd59519, 16'd35448, 16'd25599, 16'd53685, 16'd49964, 16'd21538, 16'd45503, 16'd37053, 16'd64562, 16'd38268, 16'd22256, 16'd17080, 16'd40408, 16'd53343, 16'd52706, 16'd42386, 16'd62301, 16'd10518, 16'd43514, 16'd44003, 16'd9103, 16'd25077, 16'd59541});
	test_expansion(128'hbd1bc4c0d8bc5781997815b3548b4975, {16'd31294, 16'd17825, 16'd41818, 16'd3120, 16'd292, 16'd1480, 16'd24499, 16'd21498, 16'd2120, 16'd31828, 16'd14308, 16'd12933, 16'd48676, 16'd39822, 16'd34179, 16'd53474, 16'd33182, 16'd40396, 16'd37142, 16'd7650, 16'd57707, 16'd33787, 16'd203, 16'd63083, 16'd11342, 16'd27178});
	test_expansion(128'h45c9ea3dcd6ed90678d332801e106fd9, {16'd19805, 16'd47463, 16'd19709, 16'd41924, 16'd43793, 16'd47920, 16'd62673, 16'd2135, 16'd55043, 16'd36711, 16'd36204, 16'd23658, 16'd63898, 16'd4113, 16'd62358, 16'd34324, 16'd42128, 16'd34017, 16'd34931, 16'd18417, 16'd32820, 16'd25692, 16'd61214, 16'd7710, 16'd33412, 16'd7288});
	test_expansion(128'h7024f957ac65ba149320cc7777d5029c, {16'd2346, 16'd48141, 16'd35496, 16'd21501, 16'd27238, 16'd33667, 16'd37308, 16'd10440, 16'd22959, 16'd63367, 16'd30103, 16'd50602, 16'd53753, 16'd4798, 16'd59113, 16'd54026, 16'd63217, 16'd882, 16'd43874, 16'd61981, 16'd5233, 16'd29647, 16'd4584, 16'd27491, 16'd44420, 16'd38760});
	test_expansion(128'hfa02f4dd95680bef6f2a1ddb6099f33c, {16'd11798, 16'd36268, 16'd11808, 16'd21659, 16'd56823, 16'd51732, 16'd62459, 16'd55517, 16'd47337, 16'd19084, 16'd53850, 16'd25980, 16'd18636, 16'd9824, 16'd19205, 16'd43318, 16'd40972, 16'd10144, 16'd30270, 16'd31298, 16'd52054, 16'd13177, 16'd54705, 16'd22495, 16'd43436, 16'd8040});
	test_expansion(128'h5483bd5094580f79749f19eaa6918ae4, {16'd57913, 16'd16393, 16'd62932, 16'd28361, 16'd51996, 16'd24515, 16'd62147, 16'd27788, 16'd16924, 16'd61069, 16'd30781, 16'd28160, 16'd35157, 16'd40296, 16'd2590, 16'd35163, 16'd47698, 16'd63677, 16'd37061, 16'd8115, 16'd26924, 16'd17576, 16'd56631, 16'd23050, 16'd51758, 16'd10823});
	test_expansion(128'hf7c2be38ab9a8b17eecdb956631f3e6f, {16'd30522, 16'd48686, 16'd13456, 16'd21590, 16'd32040, 16'd5324, 16'd56299, 16'd20782, 16'd28200, 16'd33176, 16'd32617, 16'd29617, 16'd34724, 16'd35211, 16'd40930, 16'd7548, 16'd63349, 16'd19256, 16'd44233, 16'd61412, 16'd61591, 16'd21320, 16'd14673, 16'd21858, 16'd53954, 16'd51409});
	test_expansion(128'hfbc9c3a77d7c61d85f1d6070d94036fa, {16'd15847, 16'd6804, 16'd807, 16'd34190, 16'd21763, 16'd30211, 16'd26624, 16'd26601, 16'd50724, 16'd35463, 16'd37697, 16'd16190, 16'd18972, 16'd54088, 16'd20864, 16'd15728, 16'd42964, 16'd55908, 16'd9389, 16'd33978, 16'd35165, 16'd42736, 16'd388, 16'd61223, 16'd9308, 16'd51222});
	test_expansion(128'h09d70d121702e7aee98fe986c5f5f523, {16'd26877, 16'd41202, 16'd14631, 16'd61523, 16'd63430, 16'd23403, 16'd54437, 16'd39709, 16'd5337, 16'd44633, 16'd50857, 16'd33411, 16'd55531, 16'd60187, 16'd35560, 16'd61233, 16'd48882, 16'd27534, 16'd36275, 16'd43123, 16'd13890, 16'd32799, 16'd2738, 16'd64226, 16'd691, 16'd39108});
	test_expansion(128'hdd291eaf1e3e4a69c250c9c985fcbd89, {16'd36251, 16'd56624, 16'd52561, 16'd50666, 16'd60596, 16'd15470, 16'd57494, 16'd32335, 16'd54503, 16'd56247, 16'd41309, 16'd36004, 16'd47577, 16'd57676, 16'd51046, 16'd211, 16'd48272, 16'd16052, 16'd29346, 16'd48411, 16'd48738, 16'd50247, 16'd5952, 16'd56209, 16'd38334, 16'd4331});
	test_expansion(128'h4b2ef4abce504d6e9458fd503c8adbb6, {16'd18765, 16'd5189, 16'd42271, 16'd34984, 16'd51872, 16'd47612, 16'd7945, 16'd28396, 16'd24073, 16'd59967, 16'd17176, 16'd16023, 16'd52488, 16'd5326, 16'd21965, 16'd37261, 16'd51621, 16'd48222, 16'd21993, 16'd23152, 16'd6527, 16'd21551, 16'd1955, 16'd61507, 16'd23835, 16'd19060});
	test_expansion(128'h16fd521ac6017f846ab1f15b83a76dc5, {16'd4655, 16'd36596, 16'd56988, 16'd34692, 16'd57954, 16'd1300, 16'd26285, 16'd9344, 16'd16584, 16'd23279, 16'd37931, 16'd62382, 16'd56800, 16'd37826, 16'd8411, 16'd31880, 16'd19921, 16'd46185, 16'd42579, 16'd1774, 16'd33876, 16'd2747, 16'd16353, 16'd44622, 16'd48113, 16'd38774});
	test_expansion(128'h34a7639727904716cbbc66f91310ab14, {16'd37881, 16'd33956, 16'd14321, 16'd36211, 16'd24190, 16'd3145, 16'd39462, 16'd59604, 16'd25954, 16'd19210, 16'd32865, 16'd12881, 16'd49448, 16'd10202, 16'd42183, 16'd43184, 16'd64780, 16'd45097, 16'd20024, 16'd53361, 16'd30437, 16'd13726, 16'd42502, 16'd49844, 16'd40955, 16'd28637});
	test_expansion(128'h3d2c3855cbe1bf5efeacbb1f69015e9a, {16'd2384, 16'd19137, 16'd6407, 16'd29986, 16'd20548, 16'd48680, 16'd46895, 16'd32156, 16'd19583, 16'd58884, 16'd23039, 16'd27679, 16'd5036, 16'd59993, 16'd2882, 16'd23429, 16'd9732, 16'd44415, 16'd54247, 16'd8629, 16'd2417, 16'd43036, 16'd12769, 16'd36210, 16'd41741, 16'd37966});
	test_expansion(128'h00cf4c1596e0812834d217ecb21cc901, {16'd25141, 16'd3216, 16'd39348, 16'd1021, 16'd44492, 16'd1153, 16'd20066, 16'd408, 16'd44874, 16'd27139, 16'd11684, 16'd32053, 16'd29236, 16'd40934, 16'd644, 16'd41368, 16'd20792, 16'd18446, 16'd47945, 16'd8965, 16'd26590, 16'd41074, 16'd16319, 16'd11904, 16'd50795, 16'd48228});
	test_expansion(128'h323a929a91555cc28bddfd954ae8c8f9, {16'd25280, 16'd3766, 16'd62853, 16'd40373, 16'd44825, 16'd31132, 16'd43212, 16'd45305, 16'd60258, 16'd24729, 16'd34233, 16'd64195, 16'd3090, 16'd45711, 16'd40532, 16'd41172, 16'd28901, 16'd24998, 16'd46213, 16'd13932, 16'd17324, 16'd22137, 16'd23732, 16'd29034, 16'd58145, 16'd24775});
	test_expansion(128'h7d44858d85825261ed3090d35549a990, {16'd13049, 16'd24543, 16'd55726, 16'd29874, 16'd50169, 16'd40301, 16'd63627, 16'd36763, 16'd56912, 16'd24628, 16'd31657, 16'd59818, 16'd63250, 16'd50744, 16'd43293, 16'd12179, 16'd19137, 16'd23562, 16'd59994, 16'd13734, 16'd32676, 16'd53918, 16'd33453, 16'd42640, 16'd22273, 16'd31333});
	test_expansion(128'hb9ddb21affdc189bb3ed16f70b9fed16, {16'd3495, 16'd24659, 16'd12753, 16'd58349, 16'd58179, 16'd54404, 16'd25258, 16'd20927, 16'd47130, 16'd18654, 16'd32394, 16'd51917, 16'd1757, 16'd13509, 16'd20507, 16'd14872, 16'd29563, 16'd27819, 16'd40189, 16'd6068, 16'd45705, 16'd38414, 16'd55508, 16'd13081, 16'd8073, 16'd14000});
	test_expansion(128'he93eabb73691e80eedf2c6e015ae3b39, {16'd2549, 16'd18465, 16'd6209, 16'd63639, 16'd27897, 16'd51909, 16'd37054, 16'd50816, 16'd15786, 16'd49436, 16'd25342, 16'd57948, 16'd30691, 16'd30808, 16'd3846, 16'd16782, 16'd45775, 16'd38336, 16'd55156, 16'd59233, 16'd11351, 16'd27106, 16'd4725, 16'd6351, 16'd30077, 16'd21731});
	test_expansion(128'h4eefdef5f99ec725fca3a8f1a41d98c8, {16'd27930, 16'd16992, 16'd64267, 16'd7392, 16'd61286, 16'd59622, 16'd9626, 16'd32318, 16'd31552, 16'd30874, 16'd48678, 16'd63171, 16'd50804, 16'd10888, 16'd60596, 16'd51626, 16'd42256, 16'd18645, 16'd55290, 16'd24334, 16'd56868, 16'd32509, 16'd18710, 16'd2410, 16'd10709, 16'd58023});
	test_expansion(128'heaa5062110065284d5b730a23c47bb06, {16'd51419, 16'd59042, 16'd54659, 16'd3674, 16'd1092, 16'd49839, 16'd64888, 16'd62319, 16'd49968, 16'd3252, 16'd49177, 16'd52273, 16'd46523, 16'd49721, 16'd24103, 16'd1349, 16'd7451, 16'd31716, 16'd63915, 16'd54075, 16'd30290, 16'd4134, 16'd13304, 16'd41413, 16'd30856, 16'd5684});
	test_expansion(128'h56e915ce9bed5aa12e49113cc6016f78, {16'd7610, 16'd2367, 16'd43073, 16'd55350, 16'd51133, 16'd52044, 16'd47754, 16'd8471, 16'd34012, 16'd15884, 16'd14906, 16'd56457, 16'd35338, 16'd36460, 16'd37240, 16'd48397, 16'd23619, 16'd64579, 16'd42762, 16'd7057, 16'd26129, 16'd18855, 16'd15472, 16'd42682, 16'd52108, 16'd35954});
	test_expansion(128'hc142d978a295320b6eb4e2a6bad71891, {16'd31428, 16'd10025, 16'd22417, 16'd12450, 16'd61651, 16'd10959, 16'd56051, 16'd21109, 16'd4738, 16'd29306, 16'd19045, 16'd5665, 16'd25753, 16'd31757, 16'd50575, 16'd56279, 16'd4394, 16'd23872, 16'd3226, 16'd36793, 16'd137, 16'd22327, 16'd536, 16'd52896, 16'd7819, 16'd50551});
	test_expansion(128'h2318980e5f490ac8ff0784c46b71ceed, {16'd18507, 16'd11386, 16'd3972, 16'd29437, 16'd19831, 16'd34975, 16'd20748, 16'd64823, 16'd59004, 16'd59608, 16'd65044, 16'd13060, 16'd56523, 16'd63001, 16'd54198, 16'd40156, 16'd31549, 16'd18572, 16'd5989, 16'd56632, 16'd33006, 16'd10290, 16'd21682, 16'd8499, 16'd10451, 16'd37549});
	test_expansion(128'he989c9e0c3cdd395296483187593051d, {16'd26750, 16'd38571, 16'd30382, 16'd53627, 16'd8594, 16'd44237, 16'd15277, 16'd45929, 16'd35683, 16'd39945, 16'd60174, 16'd33402, 16'd24087, 16'd40952, 16'd59386, 16'd59536, 16'd28013, 16'd10097, 16'd40485, 16'd36629, 16'd57818, 16'd61962, 16'd34642, 16'd10689, 16'd1694, 16'd20612});
	test_expansion(128'h4c90eb79a950bb05f203474f4d4704d8, {16'd10671, 16'd63730, 16'd58239, 16'd1628, 16'd6577, 16'd46634, 16'd12246, 16'd44964, 16'd4729, 16'd1249, 16'd15770, 16'd17992, 16'd27767, 16'd13327, 16'd61938, 16'd28397, 16'd6645, 16'd42238, 16'd65360, 16'd36432, 16'd55011, 16'd55445, 16'd7733, 16'd11739, 16'd41893, 16'd34258});
	test_expansion(128'he8336c6ed21c0aade5262dd5ed14744c, {16'd31588, 16'd12543, 16'd11092, 16'd1746, 16'd52055, 16'd27950, 16'd38293, 16'd8793, 16'd33319, 16'd17914, 16'd52861, 16'd6135, 16'd27305, 16'd11476, 16'd64136, 16'd50034, 16'd48292, 16'd101, 16'd63708, 16'd41537, 16'd21624, 16'd7768, 16'd55099, 16'd53775, 16'd26847, 16'd27927});
	test_expansion(128'h7b8603903a713ed04276149708b6a30e, {16'd52728, 16'd15129, 16'd22309, 16'd49821, 16'd60458, 16'd56387, 16'd46575, 16'd55780, 16'd48349, 16'd24864, 16'd46670, 16'd5587, 16'd34279, 16'd41347, 16'd19570, 16'd62809, 16'd13838, 16'd29080, 16'd24649, 16'd52751, 16'd60416, 16'd59771, 16'd3659, 16'd4231, 16'd51465, 16'd55274});
	test_expansion(128'h34c4d2b1564559dab07a8ca3d273cc61, {16'd34296, 16'd33315, 16'd59019, 16'd32399, 16'd29306, 16'd30650, 16'd26291, 16'd21096, 16'd39587, 16'd17061, 16'd54787, 16'd10688, 16'd38243, 16'd59549, 16'd57532, 16'd15809, 16'd2950, 16'd20767, 16'd2731, 16'd22158, 16'd45805, 16'd49526, 16'd6954, 16'd51090, 16'd6097, 16'd38170});
	test_expansion(128'hfc38b80961a68ba56b1b49bfa44be2cb, {16'd12623, 16'd321, 16'd57176, 16'd7878, 16'd31317, 16'd57296, 16'd51750, 16'd29456, 16'd31049, 16'd43194, 16'd22505, 16'd16885, 16'd13335, 16'd48305, 16'd17302, 16'd33581, 16'd53059, 16'd35267, 16'd9840, 16'd11509, 16'd16198, 16'd24692, 16'd10451, 16'd28775, 16'd29854, 16'd58995});
	test_expansion(128'hbb07d15d8489bc3aed649d4bf6d8c925, {16'd44494, 16'd46748, 16'd63077, 16'd28683, 16'd3183, 16'd15349, 16'd17158, 16'd3480, 16'd53870, 16'd40229, 16'd16172, 16'd49435, 16'd29323, 16'd26810, 16'd52764, 16'd6428, 16'd41226, 16'd18433, 16'd47714, 16'd8724, 16'd41822, 16'd44870, 16'd2045, 16'd5747, 16'd24616, 16'd11477});
	test_expansion(128'h4b28b08267a963fb2a97accb93da5670, {16'd7807, 16'd47576, 16'd5777, 16'd10511, 16'd40298, 16'd19114, 16'd9423, 16'd46871, 16'd6202, 16'd1806, 16'd20123, 16'd56348, 16'd26783, 16'd12267, 16'd12882, 16'd58354, 16'd49034, 16'd18970, 16'd18349, 16'd47285, 16'd2386, 16'd48686, 16'd3788, 16'd34164, 16'd42965, 16'd14396});
	test_expansion(128'h11198ab86348b4d9046d065ea122fed1, {16'd38437, 16'd6216, 16'd65053, 16'd43376, 16'd15131, 16'd37749, 16'd39604, 16'd46750, 16'd6706, 16'd9770, 16'd48354, 16'd45931, 16'd45783, 16'd1317, 16'd60158, 16'd63726, 16'd2791, 16'd34965, 16'd39010, 16'd32178, 16'd13633, 16'd57517, 16'd2524, 16'd11983, 16'd23554, 16'd10655});
	test_expansion(128'h9495a1d156a25095805cb4821206ce94, {16'd61778, 16'd5582, 16'd42799, 16'd51483, 16'd37887, 16'd24958, 16'd5034, 16'd18715, 16'd59637, 16'd7331, 16'd45209, 16'd16308, 16'd34056, 16'd51462, 16'd58290, 16'd8663, 16'd28206, 16'd27141, 16'd4826, 16'd48880, 16'd27003, 16'd42953, 16'd36576, 16'd12872, 16'd48410, 16'd19391});
	test_expansion(128'h6540a2ab04b60ead29f42d42166803d2, {16'd43853, 16'd43028, 16'd34496, 16'd64359, 16'd57924, 16'd43684, 16'd8108, 16'd30549, 16'd43845, 16'd20345, 16'd32416, 16'd32156, 16'd41240, 16'd1173, 16'd532, 16'd21699, 16'd36587, 16'd54421, 16'd11096, 16'd55150, 16'd53076, 16'd24141, 16'd33118, 16'd27664, 16'd14977, 16'd23176});
	test_expansion(128'h0a718a734c64c20d35e1f15190f14cfc, {16'd31334, 16'd18877, 16'd43150, 16'd45526, 16'd9642, 16'd31754, 16'd23080, 16'd27061, 16'd30545, 16'd19250, 16'd52057, 16'd44786, 16'd4210, 16'd60463, 16'd32254, 16'd49687, 16'd45485, 16'd375, 16'd48554, 16'd8541, 16'd52561, 16'd18165, 16'd64259, 16'd63964, 16'd33625, 16'd54252});
	test_expansion(128'ha6eab4072f615f40d9d26a88a13b7f4d, {16'd4281, 16'd14081, 16'd5780, 16'd43973, 16'd53695, 16'd24940, 16'd1594, 16'd54119, 16'd59913, 16'd12161, 16'd34855, 16'd51465, 16'd33628, 16'd6028, 16'd43099, 16'd4071, 16'd56211, 16'd27527, 16'd10063, 16'd31364, 16'd38062, 16'd47992, 16'd31495, 16'd28280, 16'd8284, 16'd11731});
	test_expansion(128'h0a8fbb0ebe6d8fd2a28ef2487362c5e7, {16'd25174, 16'd59639, 16'd48862, 16'd5086, 16'd29427, 16'd17607, 16'd20965, 16'd57321, 16'd13852, 16'd59965, 16'd31762, 16'd10469, 16'd33352, 16'd41824, 16'd32152, 16'd43151, 16'd20453, 16'd3953, 16'd31155, 16'd31974, 16'd21990, 16'd38363, 16'd876, 16'd24342, 16'd58863, 16'd7468});
	test_expansion(128'hd28115836f628d22be4096f0f38041b6, {16'd38258, 16'd16549, 16'd3532, 16'd17025, 16'd18641, 16'd40416, 16'd1333, 16'd16034, 16'd58285, 16'd7842, 16'd12495, 16'd31082, 16'd45989, 16'd43671, 16'd40474, 16'd41101, 16'd56937, 16'd60248, 16'd33981, 16'd50926, 16'd25853, 16'd38609, 16'd25425, 16'd11048, 16'd23908, 16'd59491});
	test_expansion(128'h0de222d60daa5ae2720ca7e79f44d72c, {16'd19442, 16'd61140, 16'd28801, 16'd58489, 16'd41996, 16'd10393, 16'd37742, 16'd15699, 16'd50360, 16'd30053, 16'd29306, 16'd31726, 16'd22078, 16'd34407, 16'd31466, 16'd32587, 16'd57702, 16'd54693, 16'd47670, 16'd1369, 16'd61105, 16'd45602, 16'd37450, 16'd30075, 16'd28120, 16'd55262});
	test_expansion(128'h01acbb3f80e9d6248e386dbc7316240b, {16'd11814, 16'd18387, 16'd20474, 16'd52447, 16'd61645, 16'd25713, 16'd65263, 16'd58758, 16'd1661, 16'd601, 16'd6296, 16'd6216, 16'd55075, 16'd50187, 16'd44315, 16'd52931, 16'd30439, 16'd26146, 16'd20287, 16'd58727, 16'd7488, 16'd52343, 16'd34657, 16'd22420, 16'd49426, 16'd24019});
	test_expansion(128'hac6f33c3f076fd782371de655ef798b1, {16'd65259, 16'd31337, 16'd33443, 16'd60467, 16'd28242, 16'd64172, 16'd4942, 16'd49722, 16'd639, 16'd53425, 16'd21395, 16'd18192, 16'd39076, 16'd9055, 16'd28757, 16'd19039, 16'd48939, 16'd6401, 16'd61503, 16'd42291, 16'd40879, 16'd57660, 16'd1465, 16'd28183, 16'd19540, 16'd65486});
	test_expansion(128'h5b0ad6a900b62135c0576826c2672796, {16'd15148, 16'd39644, 16'd41600, 16'd30777, 16'd62323, 16'd13993, 16'd22617, 16'd47859, 16'd13847, 16'd32030, 16'd11509, 16'd43727, 16'd17855, 16'd11381, 16'd19764, 16'd56732, 16'd8095, 16'd27866, 16'd30456, 16'd41437, 16'd18314, 16'd56292, 16'd52851, 16'd28959, 16'd30366, 16'd4140});
	test_expansion(128'h81ab5e081993a7e884f7598e4bafb5ec, {16'd3875, 16'd52193, 16'd61822, 16'd19697, 16'd56821, 16'd63458, 16'd44808, 16'd31708, 16'd45489, 16'd32271, 16'd3961, 16'd13484, 16'd54625, 16'd16787, 16'd1603, 16'd34124, 16'd19619, 16'd25390, 16'd1406, 16'd48427, 16'd38663, 16'd1374, 16'd40021, 16'd8005, 16'd33407, 16'd4269});
	test_expansion(128'h16a495d32ca9a083eaef1c05a1af8a9f, {16'd58017, 16'd62599, 16'd1837, 16'd38537, 16'd27836, 16'd31859, 16'd16813, 16'd39654, 16'd15370, 16'd59919, 16'd3040, 16'd19109, 16'd1249, 16'd51082, 16'd10514, 16'd41385, 16'd61253, 16'd37698, 16'd9268, 16'd12004, 16'd40546, 16'd3789, 16'd58952, 16'd56045, 16'd2630, 16'd21202});
	test_expansion(128'h386a44a329036f49741b038d0f333048, {16'd20503, 16'd59930, 16'd4514, 16'd11325, 16'd12818, 16'd28463, 16'd253, 16'd34386, 16'd51908, 16'd47649, 16'd35603, 16'd35853, 16'd38703, 16'd18937, 16'd5922, 16'd65486, 16'd20131, 16'd1683, 16'd50570, 16'd35302, 16'd7650, 16'd2341, 16'd45645, 16'd26118, 16'd41728, 16'd31724});
	test_expansion(128'h0ea30b45fef2d64ef7ce437b990ac5d5, {16'd62180, 16'd44224, 16'd45034, 16'd11277, 16'd43294, 16'd14846, 16'd25626, 16'd20900, 16'd16505, 16'd13650, 16'd27258, 16'd19094, 16'd59634, 16'd57616, 16'd4405, 16'd58032, 16'd22741, 16'd27384, 16'd2612, 16'd39272, 16'd59445, 16'd13663, 16'd22272, 16'd9231, 16'd6602, 16'd64903});
	test_expansion(128'hde36cd33cf59a8aed8df6e6565c99fac, {16'd24569, 16'd60389, 16'd38904, 16'd45786, 16'd49820, 16'd13933, 16'd33819, 16'd4035, 16'd42302, 16'd9728, 16'd4658, 16'd62694, 16'd45585, 16'd38885, 16'd37625, 16'd43602, 16'd43325, 16'd15337, 16'd2048, 16'd29434, 16'd4850, 16'd13442, 16'd12666, 16'd24085, 16'd8924, 16'd32886});
	test_expansion(128'h770eb8f3eca4004c5fc3ab672f269c4c, {16'd37392, 16'd44815, 16'd16410, 16'd32555, 16'd13530, 16'd37518, 16'd35509, 16'd17000, 16'd52560, 16'd23330, 16'd38174, 16'd17828, 16'd3702, 16'd4324, 16'd8000, 16'd44253, 16'd27294, 16'd61992, 16'd33909, 16'd46679, 16'd62081, 16'd34619, 16'd10770, 16'd62392, 16'd56513, 16'd40513});
	test_expansion(128'h3fcca940b7043eea58f112e7ffd362ae, {16'd26837, 16'd798, 16'd57217, 16'd33222, 16'd53683, 16'd30674, 16'd16023, 16'd42448, 16'd5175, 16'd33559, 16'd28949, 16'd28786, 16'd46985, 16'd30053, 16'd29167, 16'd58675, 16'd9223, 16'd37508, 16'd27090, 16'd64074, 16'd18220, 16'd7197, 16'd23745, 16'd1782, 16'd13706, 16'd60553});
	test_expansion(128'h4ce69af82c8b23365990ee79d1d728fb, {16'd49013, 16'd4627, 16'd44663, 16'd43418, 16'd1485, 16'd47791, 16'd40206, 16'd27709, 16'd48426, 16'd60923, 16'd35343, 16'd19727, 16'd20803, 16'd62094, 16'd33614, 16'd2004, 16'd42420, 16'd40433, 16'd55527, 16'd17895, 16'd54313, 16'd26441, 16'd5629, 16'd31893, 16'd28228, 16'd34111});
	test_expansion(128'he392431fbae28de7ecfc4759f9d701db, {16'd45357, 16'd39444, 16'd21490, 16'd11469, 16'd56429, 16'd21361, 16'd19785, 16'd55323, 16'd61893, 16'd2493, 16'd27735, 16'd32325, 16'd12945, 16'd47578, 16'd29610, 16'd32220, 16'd4123, 16'd42154, 16'd10922, 16'd47158, 16'd40483, 16'd28951, 16'd47430, 16'd42127, 16'd64550, 16'd60840});
	test_expansion(128'hfdc4016a6b65ebaedee4027e083b49e7, {16'd18920, 16'd65163, 16'd23144, 16'd49681, 16'd52297, 16'd49862, 16'd47959, 16'd20482, 16'd3216, 16'd23641, 16'd5529, 16'd50789, 16'd64532, 16'd39349, 16'd64018, 16'd25020, 16'd29137, 16'd51502, 16'd64046, 16'd11674, 16'd59918, 16'd51563, 16'd28078, 16'd39213, 16'd50450, 16'd40345});
	test_expansion(128'hf951bc944658641a767c4be210d5caba, {16'd55900, 16'd34449, 16'd23013, 16'd49013, 16'd43372, 16'd12272, 16'd60091, 16'd57747, 16'd15852, 16'd44509, 16'd60244, 16'd15587, 16'd35212, 16'd46980, 16'd56013, 16'd47367, 16'd18428, 16'd40170, 16'd48964, 16'd44759, 16'd47316, 16'd7820, 16'd33216, 16'd6521, 16'd4977, 16'd28177});
	test_expansion(128'h006aee88bf56c23f02d5a67d1848ce28, {16'd14625, 16'd42026, 16'd3108, 16'd52860, 16'd19326, 16'd32185, 16'd14216, 16'd23606, 16'd5870, 16'd38072, 16'd23169, 16'd42937, 16'd7002, 16'd52754, 16'd38740, 16'd61408, 16'd59402, 16'd44888, 16'd28240, 16'd22233, 16'd61376, 16'd52311, 16'd58488, 16'd48522, 16'd9238, 16'd13});
	test_expansion(128'hb83ed04595cafd907eda218c67952607, {16'd46429, 16'd4322, 16'd52596, 16'd18879, 16'd33683, 16'd13138, 16'd52839, 16'd22195, 16'd53832, 16'd2654, 16'd27705, 16'd36981, 16'd56712, 16'd25167, 16'd24742, 16'd32455, 16'd15956, 16'd57882, 16'd35955, 16'd4583, 16'd58706, 16'd58312, 16'd40496, 16'd30196, 16'd22287, 16'd48762});
	test_expansion(128'h748ec2867cc93ebf81ccd31f0dce85c7, {16'd5616, 16'd56605, 16'd59337, 16'd9082, 16'd46115, 16'd5674, 16'd4540, 16'd19859, 16'd40430, 16'd59169, 16'd9977, 16'd57103, 16'd16704, 16'd59345, 16'd42547, 16'd7281, 16'd52557, 16'd18817, 16'd9703, 16'd28196, 16'd3836, 16'd30164, 16'd63438, 16'd13713, 16'd56963, 16'd1380});
	test_expansion(128'h96ad2eae526d390bd992620821a4b9ae, {16'd47179, 16'd2287, 16'd19892, 16'd21402, 16'd21946, 16'd59197, 16'd3190, 16'd57978, 16'd23845, 16'd57859, 16'd17619, 16'd47630, 16'd60624, 16'd12323, 16'd11689, 16'd1515, 16'd61694, 16'd42691, 16'd10717, 16'd34987, 16'd37195, 16'd9205, 16'd26187, 16'd56403, 16'd65518, 16'd40006});
	test_expansion(128'ha05adbcf036718a4d110fe6a1dc35763, {16'd31272, 16'd58729, 16'd30398, 16'd45994, 16'd53277, 16'd9902, 16'd44144, 16'd29863, 16'd58850, 16'd25437, 16'd37129, 16'd16953, 16'd6911, 16'd24728, 16'd15652, 16'd38198, 16'd4556, 16'd27675, 16'd28121, 16'd33355, 16'd35960, 16'd54122, 16'd47904, 16'd3948, 16'd37900, 16'd18475});
	test_expansion(128'h9f4951fc1447b1ee37b81c99807d90ce, {16'd53415, 16'd15195, 16'd59517, 16'd17800, 16'd16148, 16'd34802, 16'd11930, 16'd58514, 16'd13550, 16'd6056, 16'd22822, 16'd43349, 16'd24644, 16'd28582, 16'd26857, 16'd62295, 16'd615, 16'd59420, 16'd45147, 16'd57969, 16'd51337, 16'd16229, 16'd27713, 16'd13348, 16'd32146, 16'd63957});
	test_expansion(128'hd1274ae861e6478e01746b299722434b, {16'd27273, 16'd18099, 16'd63946, 16'd51587, 16'd35792, 16'd36345, 16'd15, 16'd24660, 16'd33982, 16'd22290, 16'd65312, 16'd49782, 16'd14155, 16'd28273, 16'd59448, 16'd16426, 16'd56532, 16'd31910, 16'd40166, 16'd19035, 16'd16908, 16'd62111, 16'd46041, 16'd31949, 16'd29046, 16'd1590});
	test_expansion(128'h3f2fdc54cc8fc4a6c2d62bbff5cdffdb, {16'd17074, 16'd55599, 16'd17191, 16'd24222, 16'd50515, 16'd47362, 16'd11488, 16'd24840, 16'd43092, 16'd50784, 16'd6925, 16'd54287, 16'd21169, 16'd30455, 16'd40134, 16'd50971, 16'd62972, 16'd47713, 16'd58621, 16'd53395, 16'd54492, 16'd59326, 16'd64559, 16'd8989, 16'd62717, 16'd53271});
	test_expansion(128'h91a6e8414e40fab3b6ab2d0dd749d4e4, {16'd62960, 16'd52152, 16'd37137, 16'd10831, 16'd2432, 16'd65330, 16'd24280, 16'd28903, 16'd54211, 16'd36573, 16'd13224, 16'd9578, 16'd37070, 16'd10484, 16'd5091, 16'd23729, 16'd32160, 16'd14315, 16'd63721, 16'd1158, 16'd25947, 16'd64632, 16'd62813, 16'd36248, 16'd58555, 16'd13644});
	test_expansion(128'hab90c3c4ff27262510e7f630cd5fce12, {16'd26720, 16'd26952, 16'd38476, 16'd28971, 16'd50674, 16'd23742, 16'd12508, 16'd21027, 16'd62501, 16'd25912, 16'd59460, 16'd42966, 16'd29153, 16'd28025, 16'd56485, 16'd10602, 16'd7529, 16'd14357, 16'd46766, 16'd35424, 16'd54000, 16'd41453, 16'd28963, 16'd50806, 16'd16062, 16'd39768});
	test_expansion(128'h87a17ae45000032a1722f537ed9f435e, {16'd24611, 16'd3581, 16'd25750, 16'd41365, 16'd14213, 16'd46081, 16'd11239, 16'd19475, 16'd18245, 16'd21994, 16'd6080, 16'd12920, 16'd64175, 16'd30480, 16'd41255, 16'd58141, 16'd577, 16'd60571, 16'd24655, 16'd65471, 16'd21650, 16'd996, 16'd9501, 16'd6781, 16'd54307, 16'd60275});
	test_expansion(128'h6c0058261db5818f317cf08eb4af518f, {16'd61439, 16'd4806, 16'd2904, 16'd20124, 16'd63184, 16'd63294, 16'd17049, 16'd40505, 16'd6154, 16'd9559, 16'd3038, 16'd36451, 16'd63771, 16'd7759, 16'd55702, 16'd29780, 16'd12525, 16'd55902, 16'd64943, 16'd5228, 16'd58498, 16'd19169, 16'd62487, 16'd29716, 16'd26572, 16'd33435});
	test_expansion(128'ha2327e47c981e7b5a1543dfc04a23bf8, {16'd39586, 16'd14380, 16'd17728, 16'd64222, 16'd15196, 16'd14366, 16'd12004, 16'd4357, 16'd60879, 16'd62826, 16'd42003, 16'd60279, 16'd51293, 16'd24635, 16'd52333, 16'd59466, 16'd21579, 16'd32505, 16'd57258, 16'd44314, 16'd50432, 16'd21152, 16'd357, 16'd17815, 16'd25928, 16'd31903});
	test_expansion(128'h5f1a6a7c78280886ba20a4fecf39d283, {16'd4594, 16'd42753, 16'd25437, 16'd65387, 16'd42831, 16'd6965, 16'd3764, 16'd40848, 16'd32055, 16'd38862, 16'd7467, 16'd16094, 16'd33784, 16'd15591, 16'd46166, 16'd19426, 16'd15368, 16'd53801, 16'd25697, 16'd58934, 16'd46247, 16'd48115, 16'd53982, 16'd37281, 16'd53456, 16'd15768});
	test_expansion(128'h6e8b5a6e561e0ac02e582d31d7da11e5, {16'd59669, 16'd32140, 16'd47210, 16'd51614, 16'd15181, 16'd16616, 16'd24282, 16'd12697, 16'd42906, 16'd19741, 16'd13112, 16'd35142, 16'd23310, 16'd52837, 16'd37316, 16'd58729, 16'd52087, 16'd31417, 16'd6139, 16'd44459, 16'd9740, 16'd60897, 16'd3232, 16'd59975, 16'd22295, 16'd63257});
	test_expansion(128'h51491ff3fd60d6a4de03b91cab2a59af, {16'd62919, 16'd41638, 16'd63327, 16'd54373, 16'd3538, 16'd24469, 16'd41233, 16'd57535, 16'd33697, 16'd30851, 16'd54569, 16'd27903, 16'd17847, 16'd4642, 16'd55492, 16'd45622, 16'd33274, 16'd18953, 16'd49328, 16'd46479, 16'd11251, 16'd23000, 16'd8599, 16'd28292, 16'd23530, 16'd19462});
	test_expansion(128'hbc679c3154235734d4fb3cb067ca4a1d, {16'd5832, 16'd45361, 16'd28658, 16'd6829, 16'd35120, 16'd45711, 16'd56607, 16'd52311, 16'd4652, 16'd8250, 16'd51635, 16'd23783, 16'd22248, 16'd64652, 16'd5634, 16'd52039, 16'd61118, 16'd26368, 16'd35676, 16'd4396, 16'd55727, 16'd10254, 16'd32173, 16'd22333, 16'd6461, 16'd2187});
	test_expansion(128'h5804c28520d2138c92357979d55f61ab, {16'd27507, 16'd59599, 16'd32185, 16'd30894, 16'd43158, 16'd64584, 16'd19119, 16'd42602, 16'd14046, 16'd37497, 16'd60272, 16'd17256, 16'd40901, 16'd12159, 16'd16506, 16'd62151, 16'd4664, 16'd62845, 16'd33508, 16'd49831, 16'd26581, 16'd45651, 16'd27216, 16'd44280, 16'd29048, 16'd8608});
	test_expansion(128'h73c22f054e8a2bdded1354c82acee1bf, {16'd63905, 16'd22595, 16'd4200, 16'd61277, 16'd47894, 16'd22220, 16'd30597, 16'd28495, 16'd29707, 16'd58864, 16'd57949, 16'd167, 16'd10267, 16'd5653, 16'd9405, 16'd47671, 16'd34727, 16'd60238, 16'd4766, 16'd59322, 16'd29947, 16'd53392, 16'd52499, 16'd56753, 16'd2593, 16'd5115});
	test_expansion(128'h042e5bf46190a32f3192c643b391ec73, {16'd57244, 16'd3594, 16'd15556, 16'd39307, 16'd54731, 16'd46726, 16'd24689, 16'd52157, 16'd3683, 16'd34651, 16'd47386, 16'd43973, 16'd4444, 16'd13963, 16'd11571, 16'd18157, 16'd19199, 16'd3019, 16'd52343, 16'd56403, 16'd47279, 16'd62193, 16'd53969, 16'd52508, 16'd14556, 16'd58764});
	test_expansion(128'h43c95686d8d43b14e4a232b712d9a6ad, {16'd41288, 16'd59449, 16'd44413, 16'd2677, 16'd14439, 16'd3468, 16'd10138, 16'd2116, 16'd51785, 16'd12707, 16'd25052, 16'd35985, 16'd9901, 16'd45538, 16'd29663, 16'd39864, 16'd50763, 16'd53549, 16'd29083, 16'd63879, 16'd16204, 16'd19186, 16'd29899, 16'd48913, 16'd55760, 16'd37161});
	test_expansion(128'h375a21b7c7678842767c1fa1d5cd07b1, {16'd33879, 16'd63364, 16'd30424, 16'd31260, 16'd47538, 16'd54605, 16'd47519, 16'd22753, 16'd10080, 16'd3322, 16'd26183, 16'd41469, 16'd41637, 16'd25606, 16'd35973, 16'd51502, 16'd41628, 16'd54472, 16'd8883, 16'd3322, 16'd1022, 16'd5422, 16'd32114, 16'd32879, 16'd63333, 16'd26257});
	test_expansion(128'h7007b70e32db89babeb27a2f9a000814, {16'd29442, 16'd29009, 16'd41321, 16'd50507, 16'd55237, 16'd51952, 16'd51009, 16'd15599, 16'd43613, 16'd15147, 16'd39638, 16'd40045, 16'd386, 16'd18878, 16'd36187, 16'd43035, 16'd16516, 16'd34364, 16'd15488, 16'd39530, 16'd6828, 16'd46190, 16'd25257, 16'd11919, 16'd34542, 16'd22352});
	test_expansion(128'h35e035a8276e55dfdd2d1f5a46539026, {16'd434, 16'd6632, 16'd47192, 16'd22498, 16'd7040, 16'd24030, 16'd39293, 16'd30604, 16'd5942, 16'd28894, 16'd60284, 16'd60549, 16'd46067, 16'd63624, 16'd54268, 16'd17232, 16'd6762, 16'd7134, 16'd16026, 16'd31789, 16'd46886, 16'd16117, 16'd42147, 16'd39496, 16'd32744, 16'd33755});
	test_expansion(128'h9d27a53b28ae8d3b9032b9dba0b8bb8b, {16'd28167, 16'd17477, 16'd23302, 16'd6930, 16'd110, 16'd6520, 16'd426, 16'd10681, 16'd12035, 16'd11054, 16'd34461, 16'd27651, 16'd51892, 16'd65533, 16'd60505, 16'd20224, 16'd56336, 16'd26796, 16'd45022, 16'd63044, 16'd34401, 16'd27377, 16'd13418, 16'd7681, 16'd55336, 16'd43473});
	test_expansion(128'h6acdc41c0627b850747d9ea4590308e5, {16'd47121, 16'd62379, 16'd5107, 16'd30329, 16'd107, 16'd27467, 16'd4923, 16'd65284, 16'd17850, 16'd3985, 16'd54617, 16'd34427, 16'd57768, 16'd54040, 16'd41863, 16'd43366, 16'd17773, 16'd33109, 16'd41643, 16'd44571, 16'd12584, 16'd29924, 16'd54445, 16'd60549, 16'd64920, 16'd20414});
	test_expansion(128'h65b32a164a6405e06cecd3d9087595ce, {16'd19755, 16'd44125, 16'd32920, 16'd16015, 16'd2415, 16'd45073, 16'd21787, 16'd51615, 16'd17672, 16'd21279, 16'd46052, 16'd1501, 16'd29912, 16'd54498, 16'd47894, 16'd18777, 16'd57366, 16'd19649, 16'd46066, 16'd15520, 16'd9679, 16'd64977, 16'd55981, 16'd6150, 16'd47674, 16'd61974});
	test_expansion(128'h137f86cbfe57724397dcb01144261c62, {16'd55056, 16'd51492, 16'd27384, 16'd7101, 16'd13224, 16'd4541, 16'd51246, 16'd31086, 16'd55017, 16'd53955, 16'd5730, 16'd44394, 16'd40362, 16'd13351, 16'd533, 16'd26720, 16'd27541, 16'd20740, 16'd1688, 16'd49829, 16'd1824, 16'd58893, 16'd57959, 16'd29931, 16'd49989, 16'd37909});
	test_expansion(128'h1e5338337a93c5dc32e775a1da7f728b, {16'd18056, 16'd65060, 16'd2993, 16'd26681, 16'd59168, 16'd7657, 16'd20749, 16'd52751, 16'd27282, 16'd50308, 16'd34390, 16'd31142, 16'd21233, 16'd51164, 16'd38561, 16'd28693, 16'd29569, 16'd1629, 16'd31046, 16'd52944, 16'd42731, 16'd44142, 16'd42060, 16'd5222, 16'd62725, 16'd10764});
	test_expansion(128'hc5a42ccc142b44ec3ccedc00306370ea, {16'd62214, 16'd20351, 16'd47225, 16'd52418, 16'd13916, 16'd46281, 16'd34756, 16'd22969, 16'd35941, 16'd59080, 16'd46351, 16'd58323, 16'd32327, 16'd4846, 16'd26277, 16'd6471, 16'd26498, 16'd29401, 16'd18080, 16'd37421, 16'd47926, 16'd52924, 16'd21855, 16'd34447, 16'd15128, 16'd46021});
	test_expansion(128'h3c8a45353e811bf9af7adec741841d04, {16'd50760, 16'd57331, 16'd55159, 16'd51843, 16'd45100, 16'd29501, 16'd13659, 16'd26097, 16'd11137, 16'd58301, 16'd33271, 16'd55349, 16'd56811, 16'd21352, 16'd63405, 16'd11938, 16'd3658, 16'd6324, 16'd11534, 16'd19952, 16'd57812, 16'd21547, 16'd18270, 16'd39062, 16'd32122, 16'd41172});
	test_expansion(128'hf29123ea6f3b1d73ad9326c5302bffe1, {16'd31373, 16'd64745, 16'd61811, 16'd46604, 16'd54639, 16'd27509, 16'd3963, 16'd44677, 16'd54414, 16'd16704, 16'd44340, 16'd12973, 16'd16373, 16'd27725, 16'd21309, 16'd15662, 16'd38576, 16'd38726, 16'd61408, 16'd7885, 16'd29143, 16'd42169, 16'd24041, 16'd39733, 16'd35259, 16'd61326});
	test_expansion(128'hb5d7b46df80c79c353909cc01c930311, {16'd33401, 16'd14271, 16'd1478, 16'd32879, 16'd35998, 16'd3510, 16'd1962, 16'd10100, 16'd21512, 16'd18052, 16'd24304, 16'd49898, 16'd39850, 16'd25253, 16'd62775, 16'd27464, 16'd11611, 16'd15256, 16'd21383, 16'd39706, 16'd42761, 16'd14779, 16'd57729, 16'd16636, 16'd21365, 16'd9033});
	test_expansion(128'h9595a788ffd0bd5e2388f86a5fdfb422, {16'd10746, 16'd19281, 16'd60217, 16'd6327, 16'd60963, 16'd117, 16'd22465, 16'd4503, 16'd43649, 16'd40630, 16'd52593, 16'd43492, 16'd23062, 16'd59265, 16'd55646, 16'd25699, 16'd29912, 16'd57017, 16'd25766, 16'd51429, 16'd50073, 16'd40105, 16'd30816, 16'd52700, 16'd5114, 16'd60008});
	test_expansion(128'h94cfd97a5f4fbace067e008065b7450e, {16'd1466, 16'd31457, 16'd25686, 16'd14587, 16'd44581, 16'd60744, 16'd25466, 16'd49137, 16'd38137, 16'd62084, 16'd37142, 16'd40861, 16'd36119, 16'd50427, 16'd41809, 16'd46463, 16'd12946, 16'd10243, 16'd29512, 16'd32492, 16'd28679, 16'd23936, 16'd9680, 16'd36752, 16'd44720, 16'd15352});
	test_expansion(128'h3d756b4110d79db63a129148007fd1f5, {16'd34354, 16'd37791, 16'd21526, 16'd61760, 16'd1461, 16'd26026, 16'd61467, 16'd1872, 16'd65528, 16'd35815, 16'd16609, 16'd13630, 16'd33917, 16'd55931, 16'd8979, 16'd19105, 16'd36752, 16'd45407, 16'd18756, 16'd14142, 16'd15273, 16'd60264, 16'd5246, 16'd48036, 16'd24806, 16'd4746});
	test_expansion(128'h0b721700d844fe96cdf84ee19d0ce684, {16'd7908, 16'd9407, 16'd22083, 16'd15791, 16'd6889, 16'd25079, 16'd27240, 16'd62849, 16'd48755, 16'd57996, 16'd60466, 16'd50505, 16'd5596, 16'd9306, 16'd64394, 16'd58901, 16'd5006, 16'd60025, 16'd47011, 16'd3129, 16'd1654, 16'd3887, 16'd28147, 16'd15671, 16'd65390, 16'd5169});
	test_expansion(128'h3c687b677ba753af253e7b9b03310a55, {16'd11285, 16'd20244, 16'd32537, 16'd9173, 16'd1719, 16'd4934, 16'd32265, 16'd58035, 16'd2701, 16'd51141, 16'd15683, 16'd51970, 16'd33226, 16'd39772, 16'd62391, 16'd8975, 16'd37186, 16'd33391, 16'd54053, 16'd42419, 16'd20711, 16'd5060, 16'd38939, 16'd57964, 16'd23888, 16'd58348});
	test_expansion(128'h1198d9d4919bdbaf1a74fe91a44525f5, {16'd44696, 16'd15011, 16'd9565, 16'd60558, 16'd24781, 16'd20613, 16'd18576, 16'd39333, 16'd3604, 16'd54960, 16'd11603, 16'd5479, 16'd53431, 16'd58580, 16'd35199, 16'd45568, 16'd15647, 16'd55040, 16'd21500, 16'd25172, 16'd19716, 16'd55175, 16'd15768, 16'd27663, 16'd26245, 16'd34130});
	test_expansion(128'h8a8e6abcfb04a62310c779284c6b7d82, {16'd9240, 16'd8780, 16'd26864, 16'd52907, 16'd64932, 16'd40815, 16'd11812, 16'd5052, 16'd46714, 16'd16452, 16'd12875, 16'd38994, 16'd20217, 16'd6837, 16'd63146, 16'd62116, 16'd60959, 16'd47806, 16'd49834, 16'd23142, 16'd23153, 16'd29095, 16'd28885, 16'd31667, 16'd36161, 16'd33710});
	test_expansion(128'hdf610ccce2f095464cd28becac3efbc1, {16'd3719, 16'd3948, 16'd45382, 16'd11890, 16'd50174, 16'd29093, 16'd4495, 16'd58183, 16'd55946, 16'd23794, 16'd59869, 16'd50143, 16'd62368, 16'd5255, 16'd15283, 16'd54252, 16'd65193, 16'd22925, 16'd31500, 16'd7516, 16'd51085, 16'd47414, 16'd43172, 16'd21277, 16'd60764, 16'd56433});
	test_expansion(128'h622039ab32e91c022b5d624e07445341, {16'd29234, 16'd47378, 16'd62583, 16'd60678, 16'd53469, 16'd9226, 16'd5442, 16'd34556, 16'd26481, 16'd14865, 16'd51659, 16'd40591, 16'd65062, 16'd2385, 16'd11350, 16'd11563, 16'd36413, 16'd1041, 16'd60254, 16'd24230, 16'd38627, 16'd63351, 16'd31411, 16'd17223, 16'd4508, 16'd41330});
	test_expansion(128'h16e8eeef7a7656cff3ede2385260722a, {16'd12259, 16'd2214, 16'd4998, 16'd53567, 16'd14595, 16'd62364, 16'd39287, 16'd16687, 16'd44186, 16'd53905, 16'd30062, 16'd21880, 16'd19410, 16'd54504, 16'd5275, 16'd22031, 16'd45247, 16'd20196, 16'd52996, 16'd44245, 16'd4017, 16'd46851, 16'd13384, 16'd23399, 16'd23804, 16'd19551});
	test_expansion(128'haac79f4e967beac7eb37a12fbe971249, {16'd13287, 16'd40856, 16'd5833, 16'd46689, 16'd28037, 16'd12452, 16'd35138, 16'd41265, 16'd38518, 16'd47513, 16'd9675, 16'd19726, 16'd21593, 16'd46037, 16'd17672, 16'd19978, 16'd50447, 16'd49382, 16'd63997, 16'd55794, 16'd14651, 16'd47886, 16'd62420, 16'd4295, 16'd43047, 16'd21238});
	test_expansion(128'h2d05632c4b4fd102049bedffa3f8543a, {16'd45901, 16'd11157, 16'd3051, 16'd4942, 16'd18894, 16'd49762, 16'd5355, 16'd57855, 16'd32731, 16'd44165, 16'd52752, 16'd29228, 16'd21020, 16'd12759, 16'd59636, 16'd11932, 16'd59513, 16'd30537, 16'd29961, 16'd54730, 16'd6139, 16'd3588, 16'd45717, 16'd64658, 16'd34196, 16'd13944});
	test_expansion(128'h6fd38028eeb1083149979a3e8c1d8310, {16'd23594, 16'd61372, 16'd11717, 16'd52500, 16'd6369, 16'd32342, 16'd24386, 16'd31887, 16'd17432, 16'd3977, 16'd63792, 16'd22513, 16'd1562, 16'd27247, 16'd58394, 16'd30561, 16'd26075, 16'd50002, 16'd64079, 16'd28444, 16'd19189, 16'd8136, 16'd28578, 16'd6764, 16'd39458, 16'd49324});
	test_expansion(128'h308091c6ac024b23043d2857b9045548, {16'd29625, 16'd39158, 16'd50692, 16'd4262, 16'd29720, 16'd44540, 16'd39821, 16'd48580, 16'd32889, 16'd53530, 16'd34812, 16'd63231, 16'd50067, 16'd60284, 16'd13458, 16'd42187, 16'd40023, 16'd31634, 16'd52517, 16'd61645, 16'd56978, 16'd55698, 16'd47170, 16'd42549, 16'd31954, 16'd36232});
	test_expansion(128'hf95bc6dd4b0df23a231c337ac991dc4a, {16'd18556, 16'd5657, 16'd64331, 16'd24116, 16'd34098, 16'd19411, 16'd6799, 16'd8917, 16'd31202, 16'd21233, 16'd24338, 16'd40894, 16'd41872, 16'd60524, 16'd132, 16'd9492, 16'd37003, 16'd27503, 16'd36686, 16'd37617, 16'd21648, 16'd39846, 16'd20802, 16'd60353, 16'd45218, 16'd53813});
	test_expansion(128'h9a5b1ef8ae7437fac61124160c6e419b, {16'd32750, 16'd12679, 16'd33827, 16'd52982, 16'd31932, 16'd45179, 16'd2179, 16'd15666, 16'd43454, 16'd12644, 16'd41074, 16'd19869, 16'd6638, 16'd49023, 16'd63249, 16'd60933, 16'd41198, 16'd16441, 16'd46754, 16'd38114, 16'd15185, 16'd9596, 16'd148, 16'd31144, 16'd58057, 16'd29652});
	test_expansion(128'h817059d5552364d46ce7260746ce2d2a, {16'd16675, 16'd16898, 16'd46477, 16'd32182, 16'd62225, 16'd3341, 16'd6902, 16'd51776, 16'd63026, 16'd10411, 16'd43997, 16'd1299, 16'd7095, 16'd37718, 16'd4892, 16'd47271, 16'd15082, 16'd54929, 16'd12867, 16'd37965, 16'd18432, 16'd14099, 16'd58197, 16'd41512, 16'd36804, 16'd46417});
	test_expansion(128'hf6ca2df9f348e3e38ab23a1ce982a445, {16'd12980, 16'd29942, 16'd52318, 16'd49514, 16'd56144, 16'd11812, 16'd37990, 16'd45821, 16'd31950, 16'd50631, 16'd54508, 16'd32641, 16'd47643, 16'd2694, 16'd3217, 16'd58171, 16'd52615, 16'd56823, 16'd43585, 16'd9026, 16'd63766, 16'd42008, 16'd54892, 16'd61036, 16'd7928, 16'd60640});
	test_expansion(128'hd35010cf14da9e3d1f0000af4a66e9c0, {16'd7868, 16'd34299, 16'd37698, 16'd28492, 16'd52261, 16'd63235, 16'd35632, 16'd60599, 16'd59868, 16'd5982, 16'd60611, 16'd5366, 16'd6892, 16'd48349, 16'd44086, 16'd49937, 16'd39567, 16'd26681, 16'd40072, 16'd35977, 16'd53604, 16'd4994, 16'd10747, 16'd10734, 16'd31248, 16'd50059});
	test_expansion(128'h54039f306a7a271dc7233ebdc21e0a11, {16'd7102, 16'd6257, 16'd34896, 16'd34689, 16'd33064, 16'd11281, 16'd44609, 16'd15153, 16'd57626, 16'd49626, 16'd17537, 16'd7600, 16'd42855, 16'd24761, 16'd4360, 16'd51281, 16'd10275, 16'd13055, 16'd56740, 16'd43068, 16'd16551, 16'd63465, 16'd42326, 16'd54227, 16'd34219, 16'd50618});
	test_expansion(128'hffaf557de072ed679576c7f728fd203b, {16'd36773, 16'd52048, 16'd7189, 16'd58295, 16'd64216, 16'd23508, 16'd51915, 16'd56589, 16'd45970, 16'd50336, 16'd1138, 16'd18609, 16'd30877, 16'd65214, 16'd32247, 16'd33491, 16'd53515, 16'd21339, 16'd26722, 16'd24945, 16'd64124, 16'd8394, 16'd25231, 16'd16141, 16'd56377, 16'd20287});
	test_expansion(128'hb3feb2e31a8fd32fe38096790e3274ac, {16'd48193, 16'd8812, 16'd8314, 16'd36805, 16'd3401, 16'd56724, 16'd64559, 16'd32960, 16'd9523, 16'd47690, 16'd51703, 16'd49785, 16'd25935, 16'd60559, 16'd29443, 16'd16221, 16'd44071, 16'd63950, 16'd17008, 16'd27733, 16'd55003, 16'd44787, 16'd43357, 16'd18907, 16'd56524, 16'd263});
	test_expansion(128'h61cc3ae0f7b8613cd950fc48186cb625, {16'd33636, 16'd22933, 16'd47353, 16'd44983, 16'd23070, 16'd47649, 16'd54481, 16'd27239, 16'd46212, 16'd24335, 16'd18132, 16'd23510, 16'd18087, 16'd604, 16'd1481, 16'd1549, 16'd10218, 16'd52019, 16'd63346, 16'd54835, 16'd40915, 16'd61601, 16'd17411, 16'd3767, 16'd24826, 16'd15141});
	test_expansion(128'hcf9d3ab27e2e4c249603610959d11fb8, {16'd46998, 16'd17921, 16'd15954, 16'd58464, 16'd47559, 16'd2098, 16'd63808, 16'd12637, 16'd34813, 16'd37724, 16'd19468, 16'd15920, 16'd20707, 16'd64925, 16'd51775, 16'd48978, 16'd43378, 16'd47343, 16'd10672, 16'd53811, 16'd51687, 16'd40489, 16'd48584, 16'd10626, 16'd27724, 16'd63674});
	test_expansion(128'haf6575d9a88507f127aeb3d7d4bedc97, {16'd22400, 16'd47845, 16'd60072, 16'd59821, 16'd57881, 16'd59288, 16'd5916, 16'd8184, 16'd55771, 16'd51092, 16'd62806, 16'd47350, 16'd21479, 16'd20678, 16'd4398, 16'd43018, 16'd61460, 16'd16104, 16'd62655, 16'd39699, 16'd61011, 16'd45803, 16'd8367, 16'd32112, 16'd37322, 16'd58450});
	test_expansion(128'h40e46da2e4fadc99211a8807901a87c4, {16'd31016, 16'd64554, 16'd16889, 16'd33627, 16'd14868, 16'd47899, 16'd1459, 16'd30143, 16'd31352, 16'd49031, 16'd51298, 16'd34869, 16'd45035, 16'd44618, 16'd41976, 16'd51945, 16'd40619, 16'd22351, 16'd11550, 16'd13940, 16'd49283, 16'd57720, 16'd57784, 16'd2184, 16'd44521, 16'd1269});
	test_expansion(128'h8ae28b145967587bb082cd9c545702cd, {16'd23633, 16'd35195, 16'd21173, 16'd58847, 16'd19721, 16'd41963, 16'd32883, 16'd43292, 16'd12156, 16'd34885, 16'd51912, 16'd25868, 16'd3841, 16'd44330, 16'd29271, 16'd5814, 16'd56807, 16'd52463, 16'd15572, 16'd55769, 16'd33929, 16'd40436, 16'd62700, 16'd39205, 16'd63508, 16'd50915});
	test_expansion(128'h3566e77a61b860544cd278f52a98b991, {16'd29063, 16'd30077, 16'd53243, 16'd5362, 16'd43600, 16'd55960, 16'd7240, 16'd274, 16'd53511, 16'd55473, 16'd58458, 16'd7400, 16'd32024, 16'd24870, 16'd35302, 16'd46036, 16'd28274, 16'd7970, 16'd13712, 16'd39718, 16'd2701, 16'd7946, 16'd4133, 16'd39167, 16'd1806, 16'd14292});
	test_expansion(128'hf5bdd7bc37b520524445c5af06a7f7bc, {16'd54317, 16'd15883, 16'd7301, 16'd24596, 16'd43315, 16'd62064, 16'd15334, 16'd25647, 16'd40596, 16'd11624, 16'd44485, 16'd35139, 16'd28076, 16'd16893, 16'd34265, 16'd19388, 16'd36302, 16'd37169, 16'd57297, 16'd4352, 16'd52690, 16'd41440, 16'd53324, 16'd5196, 16'd8593, 16'd27076});
	test_expansion(128'h3812634da37573c9d79655979f2b6204, {16'd18286, 16'd14801, 16'd24707, 16'd8867, 16'd22393, 16'd20189, 16'd7544, 16'd14154, 16'd33663, 16'd26004, 16'd40188, 16'd6206, 16'd37954, 16'd61976, 16'd9093, 16'd23491, 16'd61861, 16'd15545, 16'd15503, 16'd61114, 16'd27162, 16'd35288, 16'd32958, 16'd30321, 16'd3547, 16'd27328});
	test_expansion(128'hb6a57655ebd1889eb964ec8d10f605f0, {16'd64491, 16'd14018, 16'd16064, 16'd55909, 16'd64585, 16'd58226, 16'd58562, 16'd1075, 16'd55565, 16'd46899, 16'd38114, 16'd48136, 16'd49146, 16'd49790, 16'd18157, 16'd6576, 16'd4296, 16'd58094, 16'd65301, 16'd49079, 16'd7187, 16'd9739, 16'd64044, 16'd60615, 16'd8106, 16'd6638});
	test_expansion(128'h647fdba97f2dadfbb4b15f8bc93b8099, {16'd3987, 16'd63090, 16'd33413, 16'd14318, 16'd49740, 16'd56889, 16'd51853, 16'd63194, 16'd38487, 16'd54036, 16'd44015, 16'd3972, 16'd7576, 16'd29439, 16'd60895, 16'd31258, 16'd31851, 16'd57769, 16'd4945, 16'd36487, 16'd12261, 16'd60910, 16'd30621, 16'd6011, 16'd28227, 16'd43084});
	test_expansion(128'hd5ef3175868dbad1c54dec0947d7ad6e, {16'd53186, 16'd62768, 16'd34677, 16'd23394, 16'd47890, 16'd13954, 16'd49196, 16'd32035, 16'd28988, 16'd24249, 16'd25721, 16'd14739, 16'd30256, 16'd34237, 16'd33922, 16'd26371, 16'd22030, 16'd48516, 16'd2988, 16'd7216, 16'd50734, 16'd11559, 16'd53198, 16'd20045, 16'd45576, 16'd33373});
	test_expansion(128'h270255ac444691d0b3c4c1ab2239a6c1, {16'd20801, 16'd29335, 16'd22213, 16'd37220, 16'd4755, 16'd7886, 16'd1469, 16'd41813, 16'd63814, 16'd60598, 16'd4688, 16'd34298, 16'd38070, 16'd15842, 16'd13592, 16'd3368, 16'd13154, 16'd7267, 16'd46961, 16'd86, 16'd19799, 16'd16672, 16'd63207, 16'd6896, 16'd20199, 16'd42055});
	test_expansion(128'h79da6c9a9a212e2a3d97cf8dfaeb2727, {16'd30402, 16'd45687, 16'd19675, 16'd18296, 16'd3367, 16'd63874, 16'd49869, 16'd28612, 16'd60191, 16'd23255, 16'd37940, 16'd4082, 16'd51644, 16'd42284, 16'd46143, 16'd57202, 16'd22010, 16'd52588, 16'd47314, 16'd60825, 16'd22754, 16'd49556, 16'd13090, 16'd45785, 16'd29105, 16'd38821});
	test_expansion(128'h3af37a9646e9caa86a2e71434c4cb7c1, {16'd58845, 16'd2484, 16'd46146, 16'd48916, 16'd19126, 16'd3210, 16'd46476, 16'd5568, 16'd799, 16'd52333, 16'd46159, 16'd4037, 16'd64972, 16'd3205, 16'd8003, 16'd43143, 16'd44453, 16'd24486, 16'd62259, 16'd26364, 16'd58294, 16'd35334, 16'd57534, 16'd59519, 16'd42992, 16'd51689});
	test_expansion(128'h84bf87671d200e238e76a624ca8cb90a, {16'd12974, 16'd28223, 16'd51093, 16'd65530, 16'd15404, 16'd22619, 16'd17866, 16'd3740, 16'd13328, 16'd11340, 16'd48069, 16'd21218, 16'd64044, 16'd12485, 16'd51690, 16'd1624, 16'd18404, 16'd46990, 16'd42515, 16'd41401, 16'd12693, 16'd25734, 16'd65317, 16'd933, 16'd3907, 16'd4367});
	test_expansion(128'hd3fac970b33211d47cc4d404b8ff6b1e, {16'd1579, 16'd44298, 16'd50096, 16'd62901, 16'd6550, 16'd25180, 16'd32897, 16'd52286, 16'd37818, 16'd64442, 16'd64205, 16'd22833, 16'd23862, 16'd42085, 16'd882, 16'd44953, 16'd29893, 16'd16831, 16'd22022, 16'd46690, 16'd24854, 16'd40647, 16'd49163, 16'd46116, 16'd47344, 16'd61434});
	test_expansion(128'h311b44fb47b6169f22569cf9d32271eb, {16'd53823, 16'd45690, 16'd46914, 16'd54279, 16'd47693, 16'd17089, 16'd48362, 16'd54478, 16'd52902, 16'd1628, 16'd31226, 16'd52345, 16'd30681, 16'd41293, 16'd19523, 16'd45278, 16'd21071, 16'd55774, 16'd30676, 16'd35424, 16'd7099, 16'd53956, 16'd33513, 16'd51565, 16'd22728, 16'd4604});
	test_expansion(128'hb348760e354040f7c43a4411861404eb, {16'd5870, 16'd13303, 16'd14408, 16'd14267, 16'd9406, 16'd8260, 16'd7475, 16'd35204, 16'd42408, 16'd36218, 16'd23801, 16'd23663, 16'd64209, 16'd5957, 16'd14726, 16'd32409, 16'd10250, 16'd51413, 16'd34536, 16'd63992, 16'd39009, 16'd19789, 16'd3316, 16'd44938, 16'd26, 16'd30730});
	test_expansion(128'hd38cf8798bf4181150f33f3def06725f, {16'd47954, 16'd12552, 16'd53163, 16'd14055, 16'd11835, 16'd30391, 16'd26836, 16'd40362, 16'd27808, 16'd12395, 16'd10634, 16'd30659, 16'd4561, 16'd44479, 16'd12355, 16'd3120, 16'd3092, 16'd4354, 16'd62414, 16'd47258, 16'd49406, 16'd38278, 16'd64893, 16'd11478, 16'd53143, 16'd50995});
	test_expansion(128'h3bea2af64a634129530d70bf7e7f29c7, {16'd21265, 16'd49832, 16'd40911, 16'd49830, 16'd47961, 16'd12345, 16'd62330, 16'd44348, 16'd5470, 16'd7197, 16'd40493, 16'd46347, 16'd20752, 16'd16498, 16'd26552, 16'd48614, 16'd5501, 16'd62345, 16'd40195, 16'd22541, 16'd48661, 16'd28848, 16'd24641, 16'd51194, 16'd64872, 16'd61851});
	test_expansion(128'hd5b8fe4a51d1a2e6e1743585cf8e338f, {16'd2956, 16'd64550, 16'd24804, 16'd23544, 16'd23993, 16'd30807, 16'd16675, 16'd24740, 16'd42351, 16'd16813, 16'd305, 16'd19952, 16'd56043, 16'd42916, 16'd8270, 16'd50772, 16'd5698, 16'd15958, 16'd49130, 16'd37966, 16'd43008, 16'd21066, 16'd28229, 16'd18512, 16'd28823, 16'd57131});
	test_expansion(128'heebaa55a6762e5fb7693c2e76c5166ab, {16'd53919, 16'd25882, 16'd1930, 16'd6124, 16'd33928, 16'd58170, 16'd30010, 16'd51596, 16'd15740, 16'd55442, 16'd37918, 16'd51286, 16'd26665, 16'd9825, 16'd47703, 16'd20731, 16'd33586, 16'd11099, 16'd18186, 16'd50431, 16'd16776, 16'd10758, 16'd5901, 16'd2986, 16'd44380, 16'd47745});
	test_expansion(128'h94270b4b2540ec88d85ff93a1ca5c874, {16'd45523, 16'd57633, 16'd43750, 16'd44920, 16'd57780, 16'd41232, 16'd25291, 16'd45568, 16'd46938, 16'd7400, 16'd38186, 16'd61091, 16'd24239, 16'd35264, 16'd40907, 16'd6336, 16'd29679, 16'd48258, 16'd26068, 16'd33958, 16'd35969, 16'd13723, 16'd60049, 16'd24884, 16'd53961, 16'd48469});
	test_expansion(128'h95fd610735841e23ceebd1a6c49f32f1, {16'd10609, 16'd8939, 16'd17065, 16'd51997, 16'd3384, 16'd26063, 16'd49248, 16'd42731, 16'd11193, 16'd43778, 16'd48808, 16'd34531, 16'd40088, 16'd48879, 16'd33360, 16'd4128, 16'd1220, 16'd37650, 16'd47654, 16'd57951, 16'd27293, 16'd1042, 16'd59883, 16'd55422, 16'd39235, 16'd7074});
	test_expansion(128'h85e5b69247065ea749aa89762e0419a8, {16'd43704, 16'd55136, 16'd4186, 16'd53371, 16'd63880, 16'd33557, 16'd55237, 16'd17479, 16'd54605, 16'd24658, 16'd50633, 16'd23255, 16'd59697, 16'd33255, 16'd9876, 16'd35589, 16'd42883, 16'd59678, 16'd222, 16'd63016, 16'd9934, 16'd31561, 16'd7563, 16'd55325, 16'd18608, 16'd11761});
	test_expansion(128'hcccd32a2f0908e693fe55a4b8f3d4213, {16'd26974, 16'd26116, 16'd60131, 16'd24298, 16'd33782, 16'd54858, 16'd14940, 16'd14932, 16'd3569, 16'd24738, 16'd40277, 16'd13543, 16'd18549, 16'd39185, 16'd14014, 16'd60742, 16'd9866, 16'd41631, 16'd58564, 16'd16830, 16'd33101, 16'd19305, 16'd8542, 16'd1416, 16'd20765, 16'd48852});
	test_expansion(128'h8c0e825fc2e200497654ce9cdd403090, {16'd43311, 16'd23448, 16'd10980, 16'd927, 16'd30933, 16'd19093, 16'd46286, 16'd52233, 16'd34265, 16'd59921, 16'd37746, 16'd58278, 16'd16092, 16'd16240, 16'd44031, 16'd17299, 16'd24534, 16'd48816, 16'd38034, 16'd9933, 16'd45422, 16'd30256, 16'd20566, 16'd55185, 16'd41997, 16'd64861});
	test_expansion(128'h8ab445502640e0a17b9ebc8aa5a0a5b4, {16'd32950, 16'd10863, 16'd51645, 16'd12959, 16'd10545, 16'd28302, 16'd44027, 16'd26464, 16'd9904, 16'd58730, 16'd35214, 16'd28506, 16'd38538, 16'd382, 16'd1132, 16'd42667, 16'd35204, 16'd65489, 16'd23420, 16'd46529, 16'd2613, 16'd19035, 16'd15517, 16'd65103, 16'd60681, 16'd10001});
	test_expansion(128'hd62ae8822236bb48ff57ca57125522e2, {16'd29652, 16'd59148, 16'd24358, 16'd28960, 16'd25175, 16'd15320, 16'd20311, 16'd29880, 16'd26070, 16'd49510, 16'd14176, 16'd65089, 16'd45420, 16'd58502, 16'd51877, 16'd42737, 16'd57589, 16'd53292, 16'd46859, 16'd43153, 16'd62413, 16'd33907, 16'd35465, 16'd24627, 16'd661, 16'd62489});
	test_expansion(128'h698905cf88b9cf2e918a1f4dd30da0ce, {16'd41483, 16'd31664, 16'd56461, 16'd50423, 16'd45327, 16'd55702, 16'd25844, 16'd23398, 16'd10177, 16'd24799, 16'd11257, 16'd24696, 16'd33553, 16'd1456, 16'd38542, 16'd47145, 16'd57083, 16'd50668, 16'd9853, 16'd28067, 16'd32634, 16'd20951, 16'd49903, 16'd18265, 16'd15483, 16'd39415});
	test_expansion(128'h6a811d6ba14cd29c06f39a9c45034c74, {16'd7116, 16'd18923, 16'd58653, 16'd378, 16'd40229, 16'd58921, 16'd16416, 16'd65002, 16'd64975, 16'd8267, 16'd28560, 16'd31253, 16'd8938, 16'd31122, 16'd49311, 16'd51125, 16'd62458, 16'd11834, 16'd47570, 16'd45706, 16'd49738, 16'd8385, 16'd34999, 16'd44590, 16'd62947, 16'd8411});
	test_expansion(128'h5a282bc39b19e70b6f5b1bf651d4ff45, {16'd47285, 16'd13623, 16'd28920, 16'd11435, 16'd19825, 16'd908, 16'd32979, 16'd56255, 16'd15957, 16'd40475, 16'd36114, 16'd21964, 16'd55917, 16'd9589, 16'd58344, 16'd15747, 16'd30570, 16'd29663, 16'd13748, 16'd753, 16'd16552, 16'd19752, 16'd9852, 16'd60407, 16'd6426, 16'd22419});
	test_expansion(128'h36fe32ea7d122cd4e7836b145cc284c8, {16'd52735, 16'd9654, 16'd65257, 16'd64897, 16'd36797, 16'd58211, 16'd64536, 16'd13096, 16'd27168, 16'd1121, 16'd15419, 16'd63716, 16'd23507, 16'd29901, 16'd55457, 16'd48361, 16'd37461, 16'd9063, 16'd1910, 16'd30531, 16'd48344, 16'd62853, 16'd26469, 16'd46659, 16'd29044, 16'd20595});
	test_expansion(128'heca47cfbaf29807a0af8e6f8dd7768eb, {16'd3780, 16'd48752, 16'd59355, 16'd16596, 16'd26990, 16'd27392, 16'd33086, 16'd13240, 16'd45894, 16'd32234, 16'd63901, 16'd38712, 16'd17721, 16'd53559, 16'd45128, 16'd43559, 16'd50476, 16'd48334, 16'd41271, 16'd52520, 16'd24257, 16'd55133, 16'd41710, 16'd23930, 16'd27651, 16'd15206});
	test_expansion(128'h923424f431e62f33358c7ae5c8dea8e2, {16'd34916, 16'd24387, 16'd14183, 16'd46532, 16'd57718, 16'd32868, 16'd34607, 16'd33708, 16'd5302, 16'd34072, 16'd45859, 16'd7909, 16'd21043, 16'd46897, 16'd64557, 16'd51946, 16'd62773, 16'd43930, 16'd51687, 16'd33403, 16'd7800, 16'd32105, 16'd22591, 16'd46205, 16'd1253, 16'd11705});
	test_expansion(128'h6564044a8d36f1242fd7f00b0b6f5a46, {16'd64892, 16'd58132, 16'd7280, 16'd44756, 16'd23514, 16'd46620, 16'd10507, 16'd3083, 16'd43687, 16'd65046, 16'd54140, 16'd35866, 16'd6929, 16'd35776, 16'd21407, 16'd43709, 16'd30826, 16'd39754, 16'd43226, 16'd37671, 16'd41361, 16'd25429, 16'd60946, 16'd15441, 16'd12447, 16'd22810});
	test_expansion(128'hcbfbe635ffa43e1d9059566e593fc0bf, {16'd45579, 16'd33694, 16'd9002, 16'd14976, 16'd2061, 16'd41776, 16'd65063, 16'd27860, 16'd2125, 16'd42752, 16'd37803, 16'd5740, 16'd40734, 16'd10560, 16'd60925, 16'd37629, 16'd32591, 16'd39123, 16'd59932, 16'd39619, 16'd56158, 16'd62548, 16'd46988, 16'd2633, 16'd34070, 16'd64559});
	test_expansion(128'hd0f6ddacd4cec0739811bf1b56dbe8b2, {16'd45241, 16'd46840, 16'd57129, 16'd59528, 16'd37649, 16'd40650, 16'd10529, 16'd2208, 16'd6982, 16'd56269, 16'd65049, 16'd54978, 16'd25578, 16'd56589, 16'd58455, 16'd50850, 16'd44563, 16'd49380, 16'd36261, 16'd10814, 16'd4155, 16'd25825, 16'd8661, 16'd12705, 16'd63503, 16'd10760});
	test_expansion(128'hef704e845106aff269ab33ea7c471c33, {16'd44187, 16'd45885, 16'd9603, 16'd44416, 16'd44698, 16'd35116, 16'd26372, 16'd38808, 16'd62960, 16'd27503, 16'd18313, 16'd11470, 16'd39207, 16'd12371, 16'd38879, 16'd13103, 16'd45904, 16'd28008, 16'd50806, 16'd63011, 16'd7766, 16'd18759, 16'd57631, 16'd62610, 16'd46916, 16'd9715});
	test_expansion(128'hb419be5c230799775c5d592f2051ba04, {16'd62745, 16'd62840, 16'd49788, 16'd11500, 16'd2863, 16'd14474, 16'd35034, 16'd58429, 16'd44842, 16'd52960, 16'd13866, 16'd35147, 16'd55620, 16'd65238, 16'd57837, 16'd21837, 16'd52628, 16'd12042, 16'd7648, 16'd37041, 16'd5277, 16'd60667, 16'd17972, 16'd58163, 16'd31130, 16'd17560});
	test_expansion(128'h9c0bb5d4c01a156b8fb2fe5754a9e1cb, {16'd32851, 16'd55202, 16'd58866, 16'd36526, 16'd33991, 16'd29882, 16'd2088, 16'd13859, 16'd4173, 16'd59761, 16'd539, 16'd34811, 16'd37168, 16'd19942, 16'd42019, 16'd44980, 16'd9767, 16'd35661, 16'd16271, 16'd45996, 16'd58223, 16'd29501, 16'd26366, 16'd64415, 16'd61626, 16'd23776});
	test_expansion(128'h6880f2d68ae8801e67b7b41c63a5fd0b, {16'd60222, 16'd55427, 16'd51811, 16'd416, 16'd61209, 16'd41965, 16'd10276, 16'd56692, 16'd44050, 16'd41631, 16'd44036, 16'd9071, 16'd43374, 16'd43746, 16'd54818, 16'd35820, 16'd29672, 16'd42520, 16'd5483, 16'd30244, 16'd62697, 16'd22761, 16'd29916, 16'd21904, 16'd54980, 16'd10625});
	test_expansion(128'h9a27affc438a2cf79a1ca2078399ef70, {16'd36196, 16'd44328, 16'd48971, 16'd58705, 16'd11754, 16'd15497, 16'd14370, 16'd48350, 16'd15062, 16'd18918, 16'd51294, 16'd29655, 16'd55189, 16'd23143, 16'd2265, 16'd63223, 16'd48397, 16'd19758, 16'd7821, 16'd36105, 16'd42755, 16'd50422, 16'd50330, 16'd41506, 16'd34521, 16'd56331});
	test_expansion(128'ha1f1e6cc7b14d3bf33a6432dfa9e30a4, {16'd6318, 16'd8347, 16'd38470, 16'd49315, 16'd23160, 16'd39861, 16'd3639, 16'd34027, 16'd38346, 16'd55037, 16'd61396, 16'd6366, 16'd47745, 16'd22641, 16'd8760, 16'd24042, 16'd49399, 16'd27507, 16'd10885, 16'd48807, 16'd36648, 16'd22426, 16'd48484, 16'd52863, 16'd6342, 16'd4974});
	test_expansion(128'h1c9bed8e0ff06fbbee128aac892eff2a, {16'd27998, 16'd26106, 16'd11075, 16'd2395, 16'd59980, 16'd26441, 16'd49136, 16'd32198, 16'd51585, 16'd65, 16'd54971, 16'd42237, 16'd38900, 16'd13748, 16'd65447, 16'd49890, 16'd49510, 16'd12500, 16'd60853, 16'd54922, 16'd50425, 16'd49969, 16'd55088, 16'd21119, 16'd37809, 16'd26499});
	test_expansion(128'h819c8f31c9069d2d2fc601b5cede620e, {16'd31859, 16'd41143, 16'd58949, 16'd64266, 16'd28101, 16'd43211, 16'd51026, 16'd20844, 16'd33115, 16'd33529, 16'd30257, 16'd21447, 16'd7164, 16'd26464, 16'd56997, 16'd8016, 16'd41084, 16'd28147, 16'd5640, 16'd27885, 16'd17831, 16'd45784, 16'd45675, 16'd34586, 16'd11730, 16'd1214});
	test_expansion(128'h10b632100910b5cfa4e8f7205c674e7c, {16'd50864, 16'd45674, 16'd6358, 16'd19828, 16'd11722, 16'd17705, 16'd34081, 16'd55668, 16'd4804, 16'd17254, 16'd43036, 16'd17812, 16'd51299, 16'd13756, 16'd34817, 16'd39639, 16'd5111, 16'd3616, 16'd12512, 16'd6546, 16'd46601, 16'd18561, 16'd43662, 16'd52331, 16'd46546, 16'd16751});
	test_expansion(128'h27dff77268e89415bcf1462c31af3fe5, {16'd47510, 16'd53526, 16'd45160, 16'd63140, 16'd42390, 16'd7711, 16'd36467, 16'd62880, 16'd2125, 16'd24842, 16'd22062, 16'd45482, 16'd35736, 16'd32774, 16'd17429, 16'd335, 16'd7780, 16'd9072, 16'd41980, 16'd13492, 16'd36343, 16'd65513, 16'd51726, 16'd48398, 16'd15814, 16'd33484});
	test_expansion(128'ha5e31edbdcf6b667573ce47c5fbcb787, {16'd65154, 16'd42774, 16'd11608, 16'd28401, 16'd13987, 16'd15666, 16'd49996, 16'd21806, 16'd18710, 16'd19662, 16'd1668, 16'd139, 16'd12495, 16'd43338, 16'd35504, 16'd62627, 16'd59821, 16'd49015, 16'd9002, 16'd85, 16'd30343, 16'd267, 16'd36194, 16'd18329, 16'd31637, 16'd12077});
	test_expansion(128'hc1a033374bd7f0fbdad29bec2410a5cf, {16'd46770, 16'd62795, 16'd31975, 16'd14335, 16'd39671, 16'd57226, 16'd6392, 16'd1158, 16'd50726, 16'd42936, 16'd65164, 16'd63428, 16'd29922, 16'd26903, 16'd21925, 16'd32932, 16'd13901, 16'd20927, 16'd1563, 16'd43925, 16'd26074, 16'd43147, 16'd33321, 16'd28018, 16'd11706, 16'd63753});
	test_expansion(128'h72afbdd75f527cae9c5dc65511048921, {16'd47149, 16'd8291, 16'd41453, 16'd32989, 16'd7212, 16'd27928, 16'd37723, 16'd28445, 16'd62204, 16'd45301, 16'd15995, 16'd10781, 16'd41798, 16'd61741, 16'd43650, 16'd2162, 16'd55121, 16'd18665, 16'd44491, 16'd28091, 16'd6208, 16'd37258, 16'd3290, 16'd37310, 16'd50070, 16'd59539});
	test_expansion(128'hb87c3f220a1d56749ae7a212bf467e2f, {16'd4756, 16'd48437, 16'd59763, 16'd31968, 16'd136, 16'd25290, 16'd40791, 16'd28528, 16'd58343, 16'd63009, 16'd57309, 16'd41487, 16'd58882, 16'd46983, 16'd61571, 16'd16933, 16'd62409, 16'd46916, 16'd52160, 16'd525, 16'd62285, 16'd63563, 16'd4321, 16'd13733, 16'd19041, 16'd58713});
	test_expansion(128'h428ba8a28525897e3fa179dabdc2dce9, {16'd26072, 16'd62802, 16'd62349, 16'd10776, 16'd44881, 16'd19850, 16'd36024, 16'd46360, 16'd42011, 16'd18506, 16'd15434, 16'd22354, 16'd30088, 16'd30779, 16'd34128, 16'd34650, 16'd3168, 16'd55205, 16'd45171, 16'd37898, 16'd17228, 16'd15567, 16'd20894, 16'd29614, 16'd35054, 16'd34635});
	test_expansion(128'heff29fd12095f6eb38042ef45d43b955, {16'd7923, 16'd63954, 16'd12623, 16'd56827, 16'd12691, 16'd35058, 16'd49610, 16'd43686, 16'd4712, 16'd53921, 16'd2105, 16'd54248, 16'd16851, 16'd727, 16'd18731, 16'd54896, 16'd10176, 16'd1979, 16'd6692, 16'd16683, 16'd19534, 16'd2254, 16'd40383, 16'd970, 16'd45985, 16'd11635});
	test_expansion(128'hde335be8c83d896ab3d4635340e80b2e, {16'd50323, 16'd38927, 16'd42119, 16'd40183, 16'd46883, 16'd18852, 16'd32585, 16'd36953, 16'd46531, 16'd15796, 16'd11334, 16'd55496, 16'd50649, 16'd15128, 16'd59185, 16'd47386, 16'd56813, 16'd7964, 16'd54228, 16'd29616, 16'd54183, 16'd57312, 16'd57725, 16'd4673, 16'd41197, 16'd18672});
	test_expansion(128'h376a071e1e3fb11a8aabcbf2e71cf78f, {16'd10847, 16'd33491, 16'd11593, 16'd33579, 16'd38151, 16'd4274, 16'd45957, 16'd28160, 16'd59450, 16'd12420, 16'd24635, 16'd35399, 16'd2909, 16'd12830, 16'd46249, 16'd49034, 16'd56960, 16'd4507, 16'd13388, 16'd13420, 16'd42336, 16'd15832, 16'd22991, 16'd7594, 16'd65218, 16'd28492});
	test_expansion(128'h9a60aa295ede6d0b273303a98a19fc2a, {16'd53730, 16'd26213, 16'd11009, 16'd51070, 16'd22471, 16'd8852, 16'd29880, 16'd29697, 16'd26987, 16'd22883, 16'd20301, 16'd29750, 16'd63257, 16'd51235, 16'd51601, 16'd17417, 16'd24522, 16'd15886, 16'd36981, 16'd60749, 16'd5994, 16'd36653, 16'd58773, 16'd41979, 16'd49075, 16'd11567});
	test_expansion(128'h0be6fb5007002bb652af4b61b130e73d, {16'd16860, 16'd3307, 16'd57243, 16'd64914, 16'd3072, 16'd14912, 16'd63513, 16'd26378, 16'd53397, 16'd45287, 16'd27629, 16'd62593, 16'd2910, 16'd26752, 16'd4370, 16'd18700, 16'd53562, 16'd41470, 16'd42291, 16'd51512, 16'd4548, 16'd50416, 16'd38013, 16'd59748, 16'd41713, 16'd52066});
	test_expansion(128'h14bac838d7eff08e9038477bcd486787, {16'd35349, 16'd23355, 16'd3866, 16'd55300, 16'd32846, 16'd18056, 16'd28025, 16'd48079, 16'd3161, 16'd19047, 16'd10491, 16'd7888, 16'd22754, 16'd36717, 16'd44902, 16'd60382, 16'd28165, 16'd64588, 16'd46321, 16'd17300, 16'd25536, 16'd24596, 16'd1853, 16'd55548, 16'd21889, 16'd11775});
	test_expansion(128'hec02d4a47f7976623480d4da16e9413b, {16'd46083, 16'd32876, 16'd55669, 16'd21185, 16'd34944, 16'd7774, 16'd4391, 16'd32028, 16'd52678, 16'd47879, 16'd11945, 16'd16500, 16'd58660, 16'd55466, 16'd53496, 16'd33153, 16'd48146, 16'd43235, 16'd11564, 16'd5910, 16'd36135, 16'd3930, 16'd15326, 16'd52554, 16'd23408, 16'd22393});
	test_expansion(128'h49bb0a5a67575b648f9afe8b969b285d, {16'd6545, 16'd2536, 16'd61552, 16'd19078, 16'd40362, 16'd569, 16'd25471, 16'd40221, 16'd8832, 16'd28868, 16'd42015, 16'd48858, 16'd11262, 16'd55172, 16'd35561, 16'd10187, 16'd63824, 16'd27625, 16'd2646, 16'd8651, 16'd46889, 16'd9207, 16'd24234, 16'd59473, 16'd42049, 16'd12180});
	test_expansion(128'h77a41a7cf9248403d0bbdc5ea29a5582, {16'd58382, 16'd4586, 16'd11427, 16'd57932, 16'd4988, 16'd46213, 16'd59351, 16'd50603, 16'd23401, 16'd22767, 16'd7750, 16'd29755, 16'd42506, 16'd46812, 16'd63324, 16'd52321, 16'd53949, 16'd55640, 16'd64952, 16'd32915, 16'd26140, 16'd37658, 16'd62425, 16'd36024, 16'd9245, 16'd9310});
	test_expansion(128'h7fde34fc0f4b52c1857914e5b3f10b54, {16'd43273, 16'd31516, 16'd32871, 16'd56281, 16'd42082, 16'd21560, 16'd4999, 16'd43329, 16'd19525, 16'd39573, 16'd63761, 16'd42545, 16'd35192, 16'd32625, 16'd13968, 16'd42982, 16'd30239, 16'd3974, 16'd19492, 16'd13710, 16'd23161, 16'd1965, 16'd59589, 16'd4051, 16'd7195, 16'd31394});
	test_expansion(128'h89319c63237571b3a9e0c2d009d9151c, {16'd18085, 16'd57421, 16'd62209, 16'd13499, 16'd10636, 16'd18319, 16'd33021, 16'd392, 16'd64607, 16'd19798, 16'd9847, 16'd43473, 16'd45910, 16'd59830, 16'd52567, 16'd4414, 16'd44577, 16'd21255, 16'd47326, 16'd34205, 16'd16482, 16'd18305, 16'd21909, 16'd21656, 16'd10517, 16'd44720});
	test_expansion(128'h2e814d3bed347c16af5ac23e22fc901f, {16'd52805, 16'd20033, 16'd57531, 16'd56421, 16'd52191, 16'd24086, 16'd16821, 16'd25964, 16'd11527, 16'd37315, 16'd51811, 16'd45664, 16'd24987, 16'd45142, 16'd23231, 16'd9612, 16'd26874, 16'd34561, 16'd62640, 16'd45427, 16'd4063, 16'd31057, 16'd20561, 16'd58193, 16'd61716, 16'd36115});
	test_expansion(128'hec7b24c743468329c3f48ea179fa4cb9, {16'd3981, 16'd31967, 16'd61623, 16'd5516, 16'd26032, 16'd23247, 16'd38089, 16'd44138, 16'd57212, 16'd48595, 16'd39662, 16'd27411, 16'd9487, 16'd32655, 16'd1179, 16'd12952, 16'd42246, 16'd32627, 16'd58300, 16'd15318, 16'd63366, 16'd65090, 16'd21047, 16'd44739, 16'd32402, 16'd35289});
	test_expansion(128'h0dabdacd64d256598c8c38086135a122, {16'd15225, 16'd64311, 16'd25132, 16'd58134, 16'd5913, 16'd40640, 16'd34527, 16'd7708, 16'd64054, 16'd21959, 16'd35051, 16'd32861, 16'd27811, 16'd65133, 16'd44266, 16'd17448, 16'd36458, 16'd53589, 16'd3667, 16'd19388, 16'd6205, 16'd17430, 16'd24997, 16'd31218, 16'd63687, 16'd63024});
	test_expansion(128'h44b53f7e7a5b9786394a4bc5ceff74df, {16'd12188, 16'd9769, 16'd47399, 16'd46902, 16'd40470, 16'd17986, 16'd7497, 16'd3637, 16'd39259, 16'd11134, 16'd8970, 16'd4889, 16'd18488, 16'd33012, 16'd42097, 16'd35057, 16'd35334, 16'd54471, 16'd20162, 16'd51522, 16'd40451, 16'd12206, 16'd20184, 16'd36677, 16'd22314, 16'd37078});
	test_expansion(128'h50e2e081d534e85c66b829eeefa22082, {16'd17958, 16'd61836, 16'd41679, 16'd34950, 16'd57004, 16'd60926, 16'd57030, 16'd25199, 16'd42866, 16'd14975, 16'd50070, 16'd37702, 16'd32773, 16'd2203, 16'd19375, 16'd27321, 16'd6653, 16'd43315, 16'd17624, 16'd34779, 16'd4873, 16'd30948, 16'd41045, 16'd21633, 16'd27090, 16'd20509});
	test_expansion(128'hea6142176c95a7f8592beec21455fd40, {16'd17617, 16'd47879, 16'd52705, 16'd15622, 16'd3923, 16'd9282, 16'd8237, 16'd12291, 16'd55307, 16'd3359, 16'd8761, 16'd34096, 16'd14188, 16'd25266, 16'd33879, 16'd15591, 16'd58107, 16'd63244, 16'd35977, 16'd16481, 16'd25928, 16'd43836, 16'd52121, 16'd61849, 16'd40152, 16'd62291});
	test_expansion(128'h69c2f172dc057987a3e99a94dfbc0262, {16'd62242, 16'd42477, 16'd44654, 16'd890, 16'd60334, 16'd15678, 16'd36532, 16'd8709, 16'd64451, 16'd51298, 16'd38877, 16'd45438, 16'd10962, 16'd32936, 16'd54297, 16'd57370, 16'd19153, 16'd3716, 16'd51763, 16'd63748, 16'd62169, 16'd39433, 16'd20674, 16'd25182, 16'd41720, 16'd46348});
	test_expansion(128'hba5827c858982935c109635c2e418955, {16'd21300, 16'd22834, 16'd49749, 16'd35623, 16'd6897, 16'd24076, 16'd44937, 16'd27424, 16'd50744, 16'd63747, 16'd47637, 16'd14002, 16'd19594, 16'd36045, 16'd39430, 16'd22986, 16'd20547, 16'd44232, 16'd50286, 16'd16838, 16'd64407, 16'd2125, 16'd52530, 16'd25998, 16'd64893, 16'd1305});
	test_expansion(128'hc95e90cd0566ef92ee05edff7b94ab15, {16'd9835, 16'd45148, 16'd56200, 16'd6974, 16'd63186, 16'd59396, 16'd7199, 16'd33037, 16'd9235, 16'd40313, 16'd60581, 16'd4194, 16'd41833, 16'd5148, 16'd46546, 16'd60984, 16'd23589, 16'd59815, 16'd24535, 16'd31426, 16'd45058, 16'd2081, 16'd64331, 16'd30580, 16'd55518, 16'd40972});
	test_expansion(128'hebd6520aa7b05c37f125b80d3caf0cef, {16'd59486, 16'd14074, 16'd53940, 16'd12441, 16'd45971, 16'd24186, 16'd63422, 16'd20364, 16'd53835, 16'd47239, 16'd25013, 16'd24529, 16'd22190, 16'd19579, 16'd5590, 16'd5527, 16'd43617, 16'd2608, 16'd37005, 16'd5509, 16'd46243, 16'd33896, 16'd11671, 16'd32519, 16'd47946, 16'd45988});
	test_expansion(128'h65fc4df3497a45b3848a907e6f91bd3e, {16'd55308, 16'd1847, 16'd24656, 16'd8346, 16'd46108, 16'd52258, 16'd19229, 16'd14994, 16'd59537, 16'd11726, 16'd18872, 16'd11422, 16'd4925, 16'd37373, 16'd50243, 16'd30246, 16'd62500, 16'd33646, 16'd57961, 16'd31929, 16'd58780, 16'd17440, 16'd18352, 16'd43678, 16'd24190, 16'd37953});
	test_expansion(128'h9c7173f16928903605b7a0aaa7f9a6b1, {16'd10700, 16'd55625, 16'd58025, 16'd298, 16'd44570, 16'd63303, 16'd51975, 16'd17259, 16'd63992, 16'd25490, 16'd2989, 16'd43453, 16'd35244, 16'd59549, 16'd16492, 16'd42467, 16'd30873, 16'd58164, 16'd61389, 16'd26000, 16'd52662, 16'd48852, 16'd16665, 16'd7139, 16'd46474, 16'd27547});
	test_expansion(128'hc1467c9ba10263e9714ed48873dde406, {16'd9651, 16'd8799, 16'd34816, 16'd21342, 16'd27063, 16'd2361, 16'd35185, 16'd1506, 16'd56604, 16'd52041, 16'd45677, 16'd20141, 16'd12254, 16'd43078, 16'd63172, 16'd45130, 16'd32192, 16'd18202, 16'd55478, 16'd30758, 16'd16831, 16'd55647, 16'd50135, 16'd27385, 16'd62410, 16'd39521});
	test_expansion(128'h96c38990026d35b371acc7267baee8c4, {16'd27920, 16'd3299, 16'd44634, 16'd37270, 16'd26577, 16'd1274, 16'd51622, 16'd15060, 16'd32540, 16'd63302, 16'd1759, 16'd41761, 16'd43110, 16'd38380, 16'd22974, 16'd20512, 16'd44908, 16'd26928, 16'd59746, 16'd15064, 16'd14202, 16'd46642, 16'd54197, 16'd19299, 16'd64679, 16'd18334});
	test_expansion(128'ha49cec1af54b0fa8a724ce550ea020bd, {16'd1806, 16'd39046, 16'd39940, 16'd36466, 16'd12169, 16'd41439, 16'd11456, 16'd3508, 16'd35997, 16'd41717, 16'd53386, 16'd640, 16'd6426, 16'd30315, 16'd43067, 16'd11833, 16'd62418, 16'd24851, 16'd7359, 16'd21242, 16'd20200, 16'd22094, 16'd24004, 16'd41837, 16'd29788, 16'd14129});
	test_expansion(128'h5654515112018493e9330ebbc5a4f965, {16'd57764, 16'd45048, 16'd35609, 16'd65486, 16'd17757, 16'd22848, 16'd27655, 16'd44254, 16'd26193, 16'd33394, 16'd21660, 16'd3032, 16'd52019, 16'd18677, 16'd37431, 16'd10336, 16'd1040, 16'd26976, 16'd34612, 16'd38475, 16'd38063, 16'd51284, 16'd41902, 16'd18629, 16'd64644, 16'd1281});
	test_expansion(128'h6ef042d9a826d54e1aa99fecc99d766d, {16'd62419, 16'd31688, 16'd61525, 16'd17781, 16'd5973, 16'd22703, 16'd16409, 16'd12095, 16'd61867, 16'd3387, 16'd34933, 16'd17218, 16'd13148, 16'd61113, 16'd38608, 16'd10088, 16'd54180, 16'd19261, 16'd14153, 16'd47073, 16'd2540, 16'd52787, 16'd4594, 16'd19892, 16'd40917, 16'd64536});
	test_expansion(128'h8cf8e8463fe9930e3e6a52f487970d59, {16'd30663, 16'd62054, 16'd34937, 16'd51050, 16'd5884, 16'd45534, 16'd52618, 16'd34471, 16'd42648, 16'd58412, 16'd28961, 16'd44313, 16'd41634, 16'd49390, 16'd45635, 16'd2985, 16'd56642, 16'd3405, 16'd47241, 16'd27167, 16'd13693, 16'd43482, 16'd58358, 16'd50278, 16'd24939, 16'd10030});
	test_expansion(128'h676418decf382815ae7483799a3a4ecf, {16'd23769, 16'd61703, 16'd62969, 16'd27161, 16'd53590, 16'd45917, 16'd34122, 16'd55923, 16'd15099, 16'd12391, 16'd1155, 16'd30388, 16'd44765, 16'd47306, 16'd58245, 16'd62978, 16'd42348, 16'd46044, 16'd17844, 16'd48308, 16'd58283, 16'd1711, 16'd32251, 16'd21819, 16'd61050, 16'd32926});
	test_expansion(128'hf4302cac362a520f71d9d31b596c0673, {16'd43801, 16'd24286, 16'd44419, 16'd52354, 16'd50785, 16'd24717, 16'd55516, 16'd43916, 16'd7724, 16'd13356, 16'd7412, 16'd57609, 16'd45560, 16'd19386, 16'd56766, 16'd57074, 16'd30902, 16'd3032, 16'd30277, 16'd23681, 16'd13799, 16'd997, 16'd15040, 16'd4559, 16'd13655, 16'd45435});
	test_expansion(128'h5e9eac2ed9fc75f8c5fec0ca5ce43a68, {16'd26393, 16'd11210, 16'd23236, 16'd29127, 16'd49572, 16'd37498, 16'd41353, 16'd18748, 16'd50785, 16'd54992, 16'd38908, 16'd27317, 16'd17222, 16'd4992, 16'd253, 16'd22897, 16'd21489, 16'd4982, 16'd31162, 16'd24372, 16'd62905, 16'd62343, 16'd23961, 16'd40885, 16'd8085, 16'd39973});
	test_expansion(128'h7d47907232244972f827ce067c6287c8, {16'd45042, 16'd42811, 16'd55690, 16'd22208, 16'd10974, 16'd20722, 16'd19653, 16'd65338, 16'd51463, 16'd60108, 16'd41827, 16'd27430, 16'd5987, 16'd12043, 16'd6517, 16'd10137, 16'd21715, 16'd57596, 16'd29503, 16'd47720, 16'd39520, 16'd47218, 16'd32989, 16'd5946, 16'd7565, 16'd35088});
	test_expansion(128'hb574678bd1eb1fb57251d69669ebecb7, {16'd64386, 16'd36351, 16'd62009, 16'd20134, 16'd18090, 16'd6498, 16'd43756, 16'd39420, 16'd9483, 16'd1854, 16'd43531, 16'd10441, 16'd33599, 16'd27079, 16'd5084, 16'd55118, 16'd64478, 16'd5689, 16'd26869, 16'd58126, 16'd14805, 16'd1061, 16'd34650, 16'd40568, 16'd17896, 16'd51236});
	test_expansion(128'h612e76e08c778c04973a84b7779b3ee3, {16'd53760, 16'd49902, 16'd20960, 16'd9315, 16'd8034, 16'd29762, 16'd31973, 16'd38803, 16'd60096, 16'd10670, 16'd62895, 16'd43562, 16'd59625, 16'd27944, 16'd46127, 16'd46089, 16'd8833, 16'd9092, 16'd12837, 16'd33813, 16'd56827, 16'd24905, 16'd37045, 16'd53982, 16'd32280, 16'd36582});
	test_expansion(128'h7df3cbaa4eb851ca6cb2e1b8e8743816, {16'd22700, 16'd39702, 16'd24076, 16'd19244, 16'd40835, 16'd27037, 16'd28331, 16'd22289, 16'd1203, 16'd31453, 16'd45124, 16'd58744, 16'd61630, 16'd54430, 16'd46180, 16'd11037, 16'd49437, 16'd18348, 16'd13736, 16'd36536, 16'd29015, 16'd28138, 16'd61333, 16'd32264, 16'd20314, 16'd19838});
	test_expansion(128'hca6ce43f7c87867383d1397130e67bd4, {16'd45953, 16'd33330, 16'd53782, 16'd51584, 16'd18893, 16'd45894, 16'd55248, 16'd33800, 16'd3836, 16'd36095, 16'd63919, 16'd30727, 16'd40847, 16'd45205, 16'd58157, 16'd18469, 16'd46788, 16'd51906, 16'd58347, 16'd62191, 16'd56984, 16'd42736, 16'd41056, 16'd8489, 16'd27963, 16'd38053});
	test_expansion(128'h10a31b52c9de775b42e5917c05e70f6e, {16'd58268, 16'd49032, 16'd604, 16'd22004, 16'd48182, 16'd42396, 16'd58613, 16'd24812, 16'd18619, 16'd40683, 16'd35715, 16'd20873, 16'd37816, 16'd31729, 16'd44679, 16'd30112, 16'd31860, 16'd47145, 16'd33865, 16'd51249, 16'd5733, 16'd43706, 16'd9810, 16'd45263, 16'd58472, 16'd25931});
	test_expansion(128'hb98bbbb605048b663e8c9c7d833540c4, {16'd23919, 16'd93, 16'd11582, 16'd40155, 16'd53152, 16'd11936, 16'd50118, 16'd59059, 16'd47892, 16'd24387, 16'd47159, 16'd64754, 16'd37216, 16'd19860, 16'd16310, 16'd38724, 16'd29029, 16'd19140, 16'd9608, 16'd14615, 16'd52019, 16'd3044, 16'd23755, 16'd9265, 16'd59039, 16'd48016});
	test_expansion(128'hf0b9d37d95b840eb66dc241eea6e4987, {16'd34746, 16'd60248, 16'd57116, 16'd25595, 16'd28005, 16'd11038, 16'd29737, 16'd31397, 16'd18831, 16'd11747, 16'd60775, 16'd19296, 16'd51152, 16'd48736, 16'd36212, 16'd20922, 16'd7203, 16'd42732, 16'd13262, 16'd31385, 16'd20277, 16'd57169, 16'd16621, 16'd6613, 16'd52801, 16'd21439});
	test_expansion(128'h105b44da1ae33eec6a841c04f3fb8b70, {16'd15641, 16'd27081, 16'd24469, 16'd45949, 16'd21208, 16'd20143, 16'd2848, 16'd7728, 16'd63668, 16'd31966, 16'd5239, 16'd11881, 16'd6391, 16'd30372, 16'd7327, 16'd31514, 16'd29809, 16'd53784, 16'd17528, 16'd13272, 16'd52951, 16'd43531, 16'd14985, 16'd47815, 16'd50157, 16'd24938});
	test_expansion(128'h247988718b91408ab1a76ba8eeaa269d, {16'd61443, 16'd60202, 16'd15494, 16'd17088, 16'd32105, 16'd58154, 16'd59227, 16'd57245, 16'd42595, 16'd63421, 16'd17341, 16'd57161, 16'd20037, 16'd38765, 16'd2129, 16'd58526, 16'd15448, 16'd34988, 16'd48527, 16'd52769, 16'd5154, 16'd34997, 16'd60509, 16'd31885, 16'd425, 16'd50573});
	test_expansion(128'hdcca4586892623dff6058da97578995f, {16'd6980, 16'd50103, 16'd10401, 16'd2157, 16'd59014, 16'd44068, 16'd9360, 16'd22852, 16'd51415, 16'd46498, 16'd43402, 16'd49368, 16'd4678, 16'd10648, 16'd27005, 16'd11361, 16'd9912, 16'd9334, 16'd28833, 16'd4437, 16'd49834, 16'd6422, 16'd25419, 16'd46174, 16'd17148, 16'd26817});
	test_expansion(128'h58a351433fb5251c363b5d9b72cd064a, {16'd11544, 16'd1392, 16'd44231, 16'd8498, 16'd17198, 16'd41463, 16'd33413, 16'd51050, 16'd9915, 16'd55242, 16'd62145, 16'd15047, 16'd22958, 16'd35103, 16'd17560, 16'd30043, 16'd59750, 16'd60674, 16'd22288, 16'd44673, 16'd52351, 16'd35831, 16'd55568, 16'd23805, 16'd55776, 16'd35330});
	test_expansion(128'ha7e426f093b03002ac9295b0437b85a1, {16'd47906, 16'd25848, 16'd51137, 16'd11927, 16'd61340, 16'd17230, 16'd48614, 16'd54856, 16'd40784, 16'd4232, 16'd37609, 16'd41170, 16'd25861, 16'd17435, 16'd57678, 16'd56569, 16'd17354, 16'd4231, 16'd18803, 16'd14745, 16'd32664, 16'd9333, 16'd17693, 16'd23021, 16'd3635, 16'd8188});
	test_expansion(128'hbba709058de92a04f88a494067963eeb, {16'd7745, 16'd61646, 16'd51739, 16'd22435, 16'd59637, 16'd56037, 16'd7138, 16'd33844, 16'd4710, 16'd50684, 16'd60037, 16'd21685, 16'd55896, 16'd64079, 16'd42246, 16'd12114, 16'd50845, 16'd52877, 16'd43442, 16'd53598, 16'd5266, 16'd40486, 16'd7256, 16'd27293, 16'd17580, 16'd33683});
	test_expansion(128'he18a0da19babbb371c38ce6c0b7c0db2, {16'd28079, 16'd7376, 16'd7588, 16'd38552, 16'd27320, 16'd488, 16'd26578, 16'd19687, 16'd55299, 16'd59295, 16'd17463, 16'd18113, 16'd13037, 16'd1629, 16'd21840, 16'd29539, 16'd37565, 16'd16755, 16'd22963, 16'd46099, 16'd59349, 16'd24270, 16'd36419, 16'd19489, 16'd26074, 16'd52046});
	test_expansion(128'h7559ce55f7a4c20eb7b595185192a588, {16'd21239, 16'd1111, 16'd9623, 16'd56728, 16'd26610, 16'd38807, 16'd14872, 16'd65388, 16'd27198, 16'd49874, 16'd3130, 16'd44865, 16'd59174, 16'd16564, 16'd60238, 16'd31943, 16'd12826, 16'd23960, 16'd28473, 16'd49428, 16'd8166, 16'd12351, 16'd39343, 16'd19950, 16'd25584, 16'd28523});
	test_expansion(128'h34f9dc06e547a052cdc36b49003b7885, {16'd11286, 16'd21986, 16'd44991, 16'd29670, 16'd17876, 16'd17166, 16'd46205, 16'd15407, 16'd7774, 16'd49785, 16'd27671, 16'd29504, 16'd21823, 16'd53249, 16'd37827, 16'd24835, 16'd51491, 16'd12339, 16'd61097, 16'd10762, 16'd61187, 16'd6896, 16'd48011, 16'd64986, 16'd14955, 16'd21957});
	test_expansion(128'h5fa42f4441efecd90abe79d59632d6d7, {16'd6530, 16'd56983, 16'd16083, 16'd33791, 16'd24016, 16'd5622, 16'd25226, 16'd8979, 16'd30711, 16'd27689, 16'd36100, 16'd46375, 16'd38419, 16'd22322, 16'd16099, 16'd54312, 16'd9747, 16'd14641, 16'd22115, 16'd10159, 16'd22531, 16'd62506, 16'd5789, 16'd59819, 16'd4344, 16'd39924});
	test_expansion(128'h180debce164be8ac79e4db9425636952, {16'd62010, 16'd4860, 16'd11838, 16'd64247, 16'd1895, 16'd31765, 16'd52199, 16'd31809, 16'd31545, 16'd31384, 16'd33057, 16'd46544, 16'd23754, 16'd63343, 16'd59835, 16'd28044, 16'd59343, 16'd63739, 16'd2315, 16'd45058, 16'd41991, 16'd10770, 16'd38613, 16'd52941, 16'd41243, 16'd3942});
	test_expansion(128'hd39a6bc2ccd81154b34bdcca9aa2803b, {16'd29316, 16'd21229, 16'd52631, 16'd9598, 16'd11138, 16'd31807, 16'd45973, 16'd9401, 16'd31987, 16'd15749, 16'd19296, 16'd25480, 16'd13153, 16'd60401, 16'd8553, 16'd49169, 16'd42925, 16'd12288, 16'd4571, 16'd25002, 16'd48739, 16'd46388, 16'd60163, 16'd24318, 16'd19074, 16'd63286});
	test_expansion(128'had38d04a3dd467e29d0e66131b380b7c, {16'd31796, 16'd5262, 16'd26589, 16'd23860, 16'd4284, 16'd25872, 16'd40198, 16'd58911, 16'd64144, 16'd3366, 16'd5087, 16'd43808, 16'd36808, 16'd61103, 16'd59065, 16'd41219, 16'd57340, 16'd31822, 16'd63364, 16'd20542, 16'd56223, 16'd48436, 16'd40724, 16'd28315, 16'd40845, 16'd40598});
	test_expansion(128'h3424861ad989bb00ae37bc9198d8a064, {16'd42834, 16'd36475, 16'd63153, 16'd7856, 16'd30838, 16'd60833, 16'd61125, 16'd32744, 16'd50937, 16'd19538, 16'd65321, 16'd50954, 16'd19355, 16'd9849, 16'd53456, 16'd6625, 16'd62400, 16'd40479, 16'd33344, 16'd53406, 16'd8179, 16'd56660, 16'd64327, 16'd43214, 16'd49309, 16'd46665});
	test_expansion(128'he8d963e79d27f3d02ef80b4b8ee5f81d, {16'd18265, 16'd5749, 16'd41950, 16'd37942, 16'd8361, 16'd47476, 16'd1659, 16'd35727, 16'd52936, 16'd41736, 16'd33985, 16'd4559, 16'd61476, 16'd8126, 16'd63730, 16'd59775, 16'd52057, 16'd54705, 16'd63151, 16'd57995, 16'd20366, 16'd31650, 16'd65243, 16'd20478, 16'd36409, 16'd23879});
	test_expansion(128'h7f890249d6832ee74e9c7985b38f32c3, {16'd20550, 16'd9363, 16'd22609, 16'd22760, 16'd24803, 16'd4481, 16'd53078, 16'd30413, 16'd24555, 16'd2102, 16'd15197, 16'd40439, 16'd47592, 16'd19014, 16'd11465, 16'd8046, 16'd37115, 16'd52940, 16'd23058, 16'd1593, 16'd51702, 16'd20323, 16'd26637, 16'd1136, 16'd48313, 16'd15802});
	test_expansion(128'h997d79ea8656a1ba6dd05055eb69e0fe, {16'd24151, 16'd54519, 16'd41714, 16'd27392, 16'd22028, 16'd32557, 16'd1089, 16'd28904, 16'd15269, 16'd38646, 16'd29162, 16'd27236, 16'd7871, 16'd49004, 16'd45234, 16'd32183, 16'd21742, 16'd30402, 16'd33428, 16'd61028, 16'd55123, 16'd40083, 16'd39871, 16'd31929, 16'd15074, 16'd3777});
	test_expansion(128'h5bc4885265400d6b67b7baf726f28b38, {16'd45144, 16'd25708, 16'd7576, 16'd3846, 16'd57165, 16'd4816, 16'd37780, 16'd60061, 16'd15007, 16'd21405, 16'd10259, 16'd10152, 16'd61440, 16'd44650, 16'd63659, 16'd28591, 16'd27291, 16'd55089, 16'd60227, 16'd30782, 16'd32775, 16'd64877, 16'd63565, 16'd12406, 16'd42427, 16'd18645});
	test_expansion(128'hfc8ad915e2ec5d0677c24e03183f0867, {16'd17746, 16'd51926, 16'd57769, 16'd8147, 16'd10451, 16'd55044, 16'd8240, 16'd48717, 16'd41186, 16'd30898, 16'd46103, 16'd7050, 16'd16152, 16'd49358, 16'd62957, 16'd44304, 16'd44379, 16'd57297, 16'd3466, 16'd29890, 16'd14140, 16'd741, 16'd1512, 16'd52883, 16'd27260, 16'd55749});
	test_expansion(128'h93c08f63641fd7105a9a633b499ca36f, {16'd43211, 16'd33021, 16'd64959, 16'd44546, 16'd64626, 16'd4770, 16'd15790, 16'd8924, 16'd30291, 16'd38245, 16'd40435, 16'd38325, 16'd64488, 16'd44061, 16'd4380, 16'd18802, 16'd913, 16'd23712, 16'd3897, 16'd8040, 16'd15029, 16'd35385, 16'd62849, 16'd50765, 16'd18132, 16'd14021});
	test_expansion(128'h1e6c005c59fd1a1da0e9a258a6ff3e28, {16'd14906, 16'd6600, 16'd27508, 16'd45712, 16'd41747, 16'd21650, 16'd43273, 16'd15086, 16'd25435, 16'd54911, 16'd16773, 16'd54729, 16'd53321, 16'd63890, 16'd49283, 16'd18658, 16'd11001, 16'd48118, 16'd29190, 16'd40638, 16'd20150, 16'd40309, 16'd20541, 16'd42117, 16'd14064, 16'd43375});
	test_expansion(128'h41a9165c6b1f2c7e151321737b018ff8, {16'd5339, 16'd58145, 16'd13922, 16'd58760, 16'd44053, 16'd717, 16'd33577, 16'd7777, 16'd43709, 16'd12133, 16'd41439, 16'd35788, 16'd37987, 16'd26840, 16'd42726, 16'd7846, 16'd19605, 16'd20996, 16'd20463, 16'd62428, 16'd12856, 16'd3160, 16'd22814, 16'd48750, 16'd62260, 16'd1180});
	test_expansion(128'h9467f78fc2f3404fd5c7148a020a4118, {16'd20723, 16'd11129, 16'd38609, 16'd4457, 16'd2424, 16'd40206, 16'd22344, 16'd52176, 16'd27280, 16'd48461, 16'd20553, 16'd48066, 16'd4028, 16'd31399, 16'd62438, 16'd29224, 16'd13497, 16'd19001, 16'd56975, 16'd27016, 16'd59412, 16'd35682, 16'd36752, 16'd49043, 16'd62953, 16'd17705});
	test_expansion(128'hc8dcea1a782771b4a69ff977d3c666c4, {16'd51065, 16'd62887, 16'd30197, 16'd34756, 16'd31054, 16'd56482, 16'd37820, 16'd56496, 16'd23026, 16'd32664, 16'd61070, 16'd16706, 16'd60108, 16'd9668, 16'd51872, 16'd26527, 16'd9325, 16'd52722, 16'd62027, 16'd61607, 16'd61231, 16'd46128, 16'd14490, 16'd39719, 16'd4420, 16'd29821});
	test_expansion(128'hb6f3edc616c35cb2afe643a7ae3653a9, {16'd21959, 16'd60934, 16'd17148, 16'd49132, 16'd6774, 16'd45118, 16'd49490, 16'd60890, 16'd19431, 16'd12325, 16'd22893, 16'd8952, 16'd50235, 16'd17004, 16'd16815, 16'd53241, 16'd45609, 16'd16487, 16'd6220, 16'd45185, 16'd4567, 16'd3428, 16'd27757, 16'd6737, 16'd7931, 16'd24866});
	test_expansion(128'hf8ccc03079535ddc60e1acec7162a124, {16'd29310, 16'd29230, 16'd1231, 16'd53159, 16'd35961, 16'd36091, 16'd28200, 16'd47383, 16'd19428, 16'd9522, 16'd40253, 16'd29676, 16'd3985, 16'd61929, 16'd2977, 16'd37289, 16'd36842, 16'd3047, 16'd932, 16'd3397, 16'd15732, 16'd16622, 16'd11224, 16'd38811, 16'd35348, 16'd19051});
	test_expansion(128'h6420686aca0f42fd580e962a551471be, {16'd31046, 16'd65433, 16'd42298, 16'd9925, 16'd9230, 16'd16411, 16'd20454, 16'd16707, 16'd42553, 16'd20135, 16'd25892, 16'd62047, 16'd10392, 16'd53955, 16'd53555, 16'd45936, 16'd58040, 16'd40934, 16'd39871, 16'd33070, 16'd52488, 16'd40365, 16'd51436, 16'd11445, 16'd42690, 16'd46895});
	test_expansion(128'ha27ab6ac656b9c46c30b80eedf423af9, {16'd57690, 16'd30345, 16'd16653, 16'd1598, 16'd3400, 16'd13400, 16'd27245, 16'd9772, 16'd33102, 16'd18573, 16'd26413, 16'd22689, 16'd40928, 16'd30512, 16'd46989, 16'd5911, 16'd23952, 16'd13832, 16'd64084, 16'd12997, 16'd41966, 16'd1441, 16'd41378, 16'd18139, 16'd31262, 16'd14770});
	test_expansion(128'h96bb04488196ca738a9b8a3c1ad03d24, {16'd19021, 16'd22043, 16'd32092, 16'd55437, 16'd40699, 16'd43368, 16'd6567, 16'd53599, 16'd57897, 16'd241, 16'd53328, 16'd3120, 16'd52477, 16'd46730, 16'd42978, 16'd30015, 16'd8905, 16'd62205, 16'd20725, 16'd50635, 16'd1337, 16'd35059, 16'd6051, 16'd17446, 16'd16881, 16'd30860});
	test_expansion(128'h6e6e8ab6f7c682cc4a5aecc2fd215bda, {16'd13935, 16'd5238, 16'd38297, 16'd46032, 16'd27318, 16'd18090, 16'd1569, 16'd32161, 16'd59020, 16'd30568, 16'd59698, 16'd61684, 16'd21784, 16'd50825, 16'd16513, 16'd34580, 16'd48622, 16'd35420, 16'd59386, 16'd45308, 16'd11598, 16'd58276, 16'd14321, 16'd41362, 16'd53786, 16'd60321});
	test_expansion(128'ha5a0dc0130424ac7358d0b803f528611, {16'd27604, 16'd61068, 16'd52602, 16'd4359, 16'd5746, 16'd14582, 16'd48598, 16'd42263, 16'd13602, 16'd54757, 16'd17680, 16'd42650, 16'd4217, 16'd42242, 16'd23285, 16'd22135, 16'd237, 16'd55419, 16'd47852, 16'd28573, 16'd48419, 16'd33775, 16'd30859, 16'd29317, 16'd50560, 16'd21255});
	test_expansion(128'h90df4687e2442f992bd075649a7ab8c3, {16'd25575, 16'd52459, 16'd21285, 16'd29441, 16'd56388, 16'd45601, 16'd14089, 16'd18095, 16'd12269, 16'd30734, 16'd19564, 16'd47953, 16'd18574, 16'd43628, 16'd41916, 16'd60581, 16'd12164, 16'd7469, 16'd46498, 16'd58826, 16'd9296, 16'd3135, 16'd14144, 16'd44932, 16'd31230, 16'd967});
	test_expansion(128'h86b313753b8dd6e251227de83545e706, {16'd48669, 16'd4363, 16'd24902, 16'd57957, 16'd2815, 16'd19350, 16'd39265, 16'd33589, 16'd40885, 16'd21710, 16'd30942, 16'd45566, 16'd28293, 16'd27539, 16'd11692, 16'd43409, 16'd28802, 16'd34522, 16'd1159, 16'd38672, 16'd242, 16'd63215, 16'd44810, 16'd56182, 16'd6891, 16'd6575});
	test_expansion(128'h189183a8e854f90b58a47e75e71c04ce, {16'd10971, 16'd6060, 16'd57593, 16'd13854, 16'd45731, 16'd61861, 16'd12030, 16'd3842, 16'd37720, 16'd347, 16'd90, 16'd47396, 16'd25962, 16'd13555, 16'd12007, 16'd22655, 16'd18736, 16'd5688, 16'd28894, 16'd24425, 16'd47553, 16'd54622, 16'd13649, 16'd9126, 16'd55784, 16'd3195});
	test_expansion(128'hfa514a4b7c8e3de0f91758d54e3d3092, {16'd5852, 16'd16882, 16'd50666, 16'd32253, 16'd6653, 16'd11219, 16'd40304, 16'd50355, 16'd49466, 16'd1611, 16'd55646, 16'd49528, 16'd12094, 16'd53835, 16'd43561, 16'd48836, 16'd4872, 16'd44725, 16'd48603, 16'd24397, 16'd60504, 16'd34138, 16'd8223, 16'd24575, 16'd35305, 16'd18357});
	test_expansion(128'hceb2572607c0a643ad6f73442c770326, {16'd29513, 16'd1498, 16'd54333, 16'd27303, 16'd35026, 16'd5294, 16'd63502, 16'd40304, 16'd39591, 16'd18460, 16'd57246, 16'd52327, 16'd52542, 16'd54767, 16'd55411, 16'd59833, 16'd5389, 16'd18383, 16'd16730, 16'd58592, 16'd43781, 16'd49261, 16'd50820, 16'd60638, 16'd54608, 16'd29988});
	test_expansion(128'hc9dec53213ecf16636af541891b5aa33, {16'd3928, 16'd40195, 16'd6312, 16'd35481, 16'd51673, 16'd65364, 16'd39224, 16'd59700, 16'd20688, 16'd3517, 16'd51255, 16'd46644, 16'd29410, 16'd16330, 16'd15970, 16'd60643, 16'd31110, 16'd44291, 16'd54493, 16'd21478, 16'd16269, 16'd19003, 16'd55340, 16'd64829, 16'd40673, 16'd61288});
	test_expansion(128'h19da4dea1b655ec3dd9f678e7f698f52, {16'd18432, 16'd8024, 16'd39505, 16'd42559, 16'd25402, 16'd27089, 16'd1092, 16'd38122, 16'd52970, 16'd38221, 16'd62475, 16'd34341, 16'd55120, 16'd46254, 16'd5015, 16'd57430, 16'd57489, 16'd25174, 16'd35145, 16'd57235, 16'd58520, 16'd58429, 16'd10777, 16'd49687, 16'd46246, 16'd59453});
	test_expansion(128'hc997d5677f0fbed45ceb3246419ddf26, {16'd41784, 16'd32937, 16'd57606, 16'd6364, 16'd1335, 16'd42979, 16'd30950, 16'd38400, 16'd48855, 16'd46072, 16'd59229, 16'd8939, 16'd15713, 16'd62565, 16'd7269, 16'd13097, 16'd2146, 16'd24478, 16'd63294, 16'd5532, 16'd2232, 16'd39840, 16'd2991, 16'd33538, 16'd46373, 16'd24121});
	test_expansion(128'h3fe4a5258116062b4acf3feb1ad00739, {16'd63977, 16'd45495, 16'd64106, 16'd44114, 16'd14852, 16'd57566, 16'd45796, 16'd14627, 16'd19076, 16'd40824, 16'd39646, 16'd64286, 16'd21505, 16'd10090, 16'd37478, 16'd5478, 16'd35541, 16'd18017, 16'd362, 16'd26815, 16'd58498, 16'd59529, 16'd50295, 16'd351, 16'd40363, 16'd62345});
	test_expansion(128'h256b1062363e882b8cf6e68a23728d0d, {16'd528, 16'd7853, 16'd953, 16'd37747, 16'd51205, 16'd60754, 16'd17437, 16'd27538, 16'd47844, 16'd16452, 16'd17924, 16'd57996, 16'd17635, 16'd23969, 16'd2811, 16'd23422, 16'd25922, 16'd15988, 16'd23328, 16'd39935, 16'd11112, 16'd38339, 16'd50907, 16'd65113, 16'd33217, 16'd51612});
	test_expansion(128'hb4601aa1883f3ee3b2c96f8a47644d06, {16'd7530, 16'd11133, 16'd23371, 16'd40305, 16'd41637, 16'd37286, 16'd39739, 16'd2636, 16'd44423, 16'd31119, 16'd17489, 16'd51477, 16'd17155, 16'd55066, 16'd10673, 16'd45762, 16'd12753, 16'd51708, 16'd4742, 16'd60650, 16'd22658, 16'd35626, 16'd10552, 16'd62838, 16'd13318, 16'd61025});
	test_expansion(128'h1d7ab113099dbeba98038c5b572b5f98, {16'd63212, 16'd20799, 16'd33004, 16'd44900, 16'd38618, 16'd54128, 16'd37473, 16'd19021, 16'd10829, 16'd40169, 16'd36038, 16'd19120, 16'd14557, 16'd30117, 16'd59129, 16'd21587, 16'd28284, 16'd19284, 16'd20880, 16'd19653, 16'd16327, 16'd59404, 16'd56810, 16'd18880, 16'd26079, 16'd41202});
	test_expansion(128'haa77dca962e4d136ecc026b69c75cd3f, {16'd24739, 16'd50965, 16'd19040, 16'd37238, 16'd51378, 16'd40422, 16'd60516, 16'd13212, 16'd27400, 16'd15636, 16'd20592, 16'd59777, 16'd22569, 16'd1492, 16'd27692, 16'd42729, 16'd15039, 16'd30180, 16'd57509, 16'd41905, 16'd62781, 16'd7488, 16'd2884, 16'd10454, 16'd20017, 16'd12853});
	test_expansion(128'h9c8b32f5cb95f79e6593bc77ecd685b9, {16'd53000, 16'd25460, 16'd31382, 16'd62605, 16'd13076, 16'd27601, 16'd58042, 16'd57498, 16'd19769, 16'd7178, 16'd64561, 16'd57430, 16'd59773, 16'd18804, 16'd26219, 16'd61892, 16'd14177, 16'd21864, 16'd27633, 16'd6639, 16'd51214, 16'd23455, 16'd13142, 16'd59434, 16'd8150, 16'd17127});
	test_expansion(128'h3975df4f2ced6d07d3dcddf924080c7b, {16'd23789, 16'd53779, 16'd26676, 16'd21546, 16'd35735, 16'd62784, 16'd52763, 16'd15110, 16'd27780, 16'd45353, 16'd49926, 16'd10684, 16'd4184, 16'd39313, 16'd29237, 16'd36027, 16'd17292, 16'd14639, 16'd37940, 16'd45563, 16'd37525, 16'd7484, 16'd25002, 16'd4033, 16'd63164, 16'd5751});
	test_expansion(128'h94686038967274814326ed04c935f8f0, {16'd64628, 16'd55301, 16'd531, 16'd43407, 16'd7112, 16'd3881, 16'd24719, 16'd25964, 16'd32956, 16'd59907, 16'd16182, 16'd53505, 16'd24052, 16'd30611, 16'd64442, 16'd7403, 16'd12433, 16'd19527, 16'd12633, 16'd54387, 16'd40387, 16'd37434, 16'd35696, 16'd28392, 16'd9811, 16'd24252});
	test_expansion(128'h9f53e26ab4f7023b9c832c03475bea5c, {16'd5717, 16'd46142, 16'd35463, 16'd59076, 16'd20495, 16'd39861, 16'd28927, 16'd42218, 16'd7620, 16'd62515, 16'd36165, 16'd32017, 16'd11204, 16'd44347, 16'd3462, 16'd56056, 16'd64740, 16'd62857, 16'd33710, 16'd51231, 16'd9267, 16'd51176, 16'd35674, 16'd58829, 16'd9053, 16'd63654});
	test_expansion(128'h100d7c5b1be297cb1be936753a1bb4bc, {16'd30322, 16'd32492, 16'd57999, 16'd15510, 16'd29618, 16'd51642, 16'd59319, 16'd21636, 16'd48614, 16'd44974, 16'd31914, 16'd33438, 16'd29747, 16'd17846, 16'd31052, 16'd30579, 16'd7216, 16'd61299, 16'd11365, 16'd58192, 16'd3149, 16'd28744, 16'd52842, 16'd4716, 16'd49835, 16'd11862});
	test_expansion(128'h879e2b821dc42e0ee659ad7babd36361, {16'd35182, 16'd9146, 16'd51575, 16'd63110, 16'd10745, 16'd47767, 16'd26871, 16'd59809, 16'd46878, 16'd27623, 16'd14033, 16'd13133, 16'd62751, 16'd43834, 16'd62217, 16'd39924, 16'd43322, 16'd42901, 16'd52340, 16'd11508, 16'd20398, 16'd63356, 16'd5283, 16'd59167, 16'd31059, 16'd37922});
	test_expansion(128'he60419db474379d2917c15ff44de2793, {16'd19860, 16'd15571, 16'd20664, 16'd44729, 16'd34416, 16'd23562, 16'd55489, 16'd13705, 16'd38754, 16'd40668, 16'd5982, 16'd38767, 16'd11707, 16'd35911, 16'd51752, 16'd3603, 16'd17178, 16'd1410, 16'd60639, 16'd47045, 16'd49005, 16'd6643, 16'd42442, 16'd49205, 16'd61344, 16'd5589});
	test_expansion(128'h785cce10a1a9fd4ddce3608023f45d77, {16'd5874, 16'd51699, 16'd34636, 16'd46275, 16'd8311, 16'd18759, 16'd29545, 16'd18351, 16'd21517, 16'd20675, 16'd63521, 16'd39596, 16'd59991, 16'd5265, 16'd8973, 16'd41481, 16'd53744, 16'd61597, 16'd47313, 16'd7399, 16'd30278, 16'd22801, 16'd18625, 16'd52047, 16'd47662, 16'd13277});
	test_expansion(128'h109d230d55bfbc0fedc514e6c61c5a8d, {16'd63356, 16'd26770, 16'd44789, 16'd62248, 16'd36860, 16'd58973, 16'd14196, 16'd63785, 16'd10084, 16'd1277, 16'd53154, 16'd57444, 16'd50234, 16'd21133, 16'd8078, 16'd3212, 16'd359, 16'd37915, 16'd64888, 16'd58965, 16'd53840, 16'd4364, 16'd64256, 16'd27875, 16'd62777, 16'd56036});
	test_expansion(128'h7f57926dca76560e64bb80a20635becd, {16'd3809, 16'd65289, 16'd36054, 16'd59249, 16'd41918, 16'd11881, 16'd44521, 16'd15847, 16'd17659, 16'd51315, 16'd11921, 16'd42236, 16'd42838, 16'd56490, 16'd61661, 16'd47888, 16'd49296, 16'd22076, 16'd41819, 16'd47574, 16'd57046, 16'd50732, 16'd25573, 16'd10553, 16'd54737, 16'd4752});
	test_expansion(128'hda5fc426d27034667149debb0d05aa4f, {16'd52128, 16'd7432, 16'd53447, 16'd14255, 16'd11882, 16'd34740, 16'd18298, 16'd3813, 16'd64404, 16'd37686, 16'd28825, 16'd34258, 16'd5783, 16'd11170, 16'd58993, 16'd9541, 16'd47384, 16'd42517, 16'd28337, 16'd44474, 16'd12618, 16'd47788, 16'd35881, 16'd54722, 16'd33259, 16'd33660});
	test_expansion(128'hf903388382cef4497f0217e0c3c73493, {16'd51876, 16'd52583, 16'd35410, 16'd57496, 16'd46289, 16'd64506, 16'd50227, 16'd20746, 16'd38308, 16'd47056, 16'd45954, 16'd21318, 16'd57974, 16'd51532, 16'd6771, 16'd59840, 16'd41511, 16'd27953, 16'd26930, 16'd55629, 16'd27077, 16'd23419, 16'd5233, 16'd36062, 16'd55968, 16'd40821});
	test_expansion(128'h3198ae21ce9e0d9670e69245ea9d6591, {16'd14940, 16'd35763, 16'd4482, 16'd14005, 16'd41210, 16'd24666, 16'd57829, 16'd4496, 16'd34868, 16'd41831, 16'd3760, 16'd12856, 16'd62974, 16'd40016, 16'd31011, 16'd58628, 16'd18187, 16'd25225, 16'd19813, 16'd19598, 16'd58917, 16'd41079, 16'd39655, 16'd59785, 16'd46743, 16'd36315});
	test_expansion(128'h71f20c50488ae0c164359f8c8c75612e, {16'd42139, 16'd11633, 16'd17164, 16'd8379, 16'd5755, 16'd51063, 16'd47366, 16'd45874, 16'd41679, 16'd6336, 16'd38971, 16'd25418, 16'd63731, 16'd11829, 16'd59373, 16'd23669, 16'd25385, 16'd52620, 16'd19461, 16'd37929, 16'd53481, 16'd35884, 16'd20235, 16'd4656, 16'd60271, 16'd31972});
	test_expansion(128'h279c9fe102cbe0ec4485844090ef87ef, {16'd3074, 16'd13358, 16'd64831, 16'd65038, 16'd1427, 16'd29218, 16'd52206, 16'd38965, 16'd5909, 16'd18677, 16'd56450, 16'd39294, 16'd60623, 16'd53667, 16'd24478, 16'd46359, 16'd30977, 16'd54205, 16'd18830, 16'd51045, 16'd36779, 16'd32875, 16'd903, 16'd26476, 16'd64705, 16'd56785});
	test_expansion(128'h9c36e41fdc92f369056021fe7717257a, {16'd50070, 16'd43027, 16'd51802, 16'd8016, 16'd6576, 16'd11052, 16'd48751, 16'd12246, 16'd52252, 16'd33865, 16'd35436, 16'd31210, 16'd3340, 16'd14787, 16'd11513, 16'd1969, 16'd37636, 16'd22551, 16'd27921, 16'd65169, 16'd56019, 16'd10037, 16'd10107, 16'd56397, 16'd24297, 16'd19695});
	test_expansion(128'hf285828705dd4eb77b14cc19a5ad88f5, {16'd27580, 16'd35623, 16'd58134, 16'd17032, 16'd24289, 16'd63900, 16'd23002, 16'd27439, 16'd49075, 16'd2084, 16'd19232, 16'd51914, 16'd50291, 16'd43254, 16'd26579, 16'd22407, 16'd51521, 16'd32958, 16'd20307, 16'd21730, 16'd42010, 16'd58608, 16'd16291, 16'd34247, 16'd46888, 16'd20145});
	test_expansion(128'hf24b930b6a0dd4ffb708b348e4f2e0b0, {16'd40669, 16'd55050, 16'd31951, 16'd15087, 16'd59589, 16'd6359, 16'd31409, 16'd31222, 16'd60639, 16'd35190, 16'd6866, 16'd20681, 16'd18402, 16'd11445, 16'd17443, 16'd20923, 16'd21256, 16'd16703, 16'd10117, 16'd22839, 16'd44609, 16'd50499, 16'd21582, 16'd21039, 16'd41471, 16'd15365});
	test_expansion(128'h36344501a57f71a6c9633759a05b9151, {16'd19680, 16'd64887, 16'd29384, 16'd46012, 16'd45343, 16'd12622, 16'd32013, 16'd64221, 16'd9809, 16'd29009, 16'd49385, 16'd46578, 16'd36482, 16'd64076, 16'd51217, 16'd52946, 16'd41317, 16'd58172, 16'd15056, 16'd10246, 16'd16420, 16'd25041, 16'd5217, 16'd7267, 16'd10072, 16'd4813});
	test_expansion(128'h9f1078cb7f78dced77087531a6670bbc, {16'd57565, 16'd62846, 16'd9896, 16'd45861, 16'd5492, 16'd42123, 16'd18551, 16'd39700, 16'd14914, 16'd5364, 16'd32760, 16'd34355, 16'd31372, 16'd38972, 16'd36851, 16'd52402, 16'd3251, 16'd15772, 16'd10853, 16'd60077, 16'd27153, 16'd21227, 16'd60335, 16'd55636, 16'd15844, 16'd11889});
	test_expansion(128'heb7b618a9c55272407b79e4fbe48d5cb, {16'd61065, 16'd48650, 16'd42109, 16'd8670, 16'd4606, 16'd14397, 16'd5292, 16'd59928, 16'd34264, 16'd4942, 16'd23725, 16'd51080, 16'd47526, 16'd27514, 16'd23140, 16'd27179, 16'd13160, 16'd62705, 16'd30414, 16'd5315, 16'd35500, 16'd20342, 16'd35486, 16'd40255, 16'd14661, 16'd16131});
	test_expansion(128'hf4ca9a5a5d0927fa98b24e33fb628018, {16'd51991, 16'd25842, 16'd36706, 16'd23949, 16'd62126, 16'd4155, 16'd64833, 16'd34641, 16'd23415, 16'd19231, 16'd63194, 16'd57772, 16'd32389, 16'd35507, 16'd60153, 16'd3650, 16'd63629, 16'd19629, 16'd44172, 16'd2633, 16'd64624, 16'd38524, 16'd29780, 16'd11457, 16'd64012, 16'd18621});
	test_expansion(128'hc3b5d33abbe550895f412988bf073fdb, {16'd65347, 16'd17899, 16'd5994, 16'd31187, 16'd20117, 16'd7229, 16'd3001, 16'd6100, 16'd39518, 16'd4617, 16'd47653, 16'd7889, 16'd44803, 16'd2393, 16'd34168, 16'd13750, 16'd17651, 16'd37248, 16'd53429, 16'd44759, 16'd40950, 16'd13532, 16'd13438, 16'd41309, 16'd31841, 16'd62338});
	test_expansion(128'hf3b27c31e8ad29fdbc4560f8a56255a2, {16'd12258, 16'd52048, 16'd26107, 16'd15280, 16'd27726, 16'd46124, 16'd15042, 16'd9853, 16'd49955, 16'd5156, 16'd45173, 16'd38883, 16'd53870, 16'd37228, 16'd32200, 16'd10446, 16'd49508, 16'd31976, 16'd43378, 16'd2080, 16'd38357, 16'd60215, 16'd64471, 16'd5997, 16'd46660, 16'd53921});
	test_expansion(128'hecbb9e326dbffaaf19c4aad5b2c540a6, {16'd21921, 16'd42271, 16'd8633, 16'd3930, 16'd44123, 16'd48925, 16'd35241, 16'd31257, 16'd52029, 16'd35781, 16'd11278, 16'd5716, 16'd8382, 16'd63628, 16'd20287, 16'd2174, 16'd13475, 16'd33358, 16'd2683, 16'd25327, 16'd40659, 16'd40053, 16'd9252, 16'd50912, 16'd57055, 16'd34986});
	test_expansion(128'hf908a02f32948ad274646b7483624ab5, {16'd20211, 16'd20373, 16'd13322, 16'd36108, 16'd8285, 16'd30756, 16'd15813, 16'd63401, 16'd44225, 16'd26185, 16'd43734, 16'd24953, 16'd50442, 16'd6146, 16'd53114, 16'd53439, 16'd38578, 16'd28195, 16'd1090, 16'd57859, 16'd21287, 16'd48662, 16'd61101, 16'd17632, 16'd18627, 16'd21974});
	test_expansion(128'h02dd6fc011b5e3f3fedd63d67888699d, {16'd29831, 16'd53675, 16'd61139, 16'd44055, 16'd34879, 16'd10920, 16'd39695, 16'd58334, 16'd9854, 16'd42879, 16'd9581, 16'd56928, 16'd21250, 16'd30859, 16'd64139, 16'd58745, 16'd7925, 16'd15966, 16'd57568, 16'd14088, 16'd9967, 16'd45913, 16'd61129, 16'd35095, 16'd6477, 16'd33703});
	test_expansion(128'h8f66b9cf9d415e2d1ee10b6bf6b07321, {16'd49614, 16'd1046, 16'd110, 16'd64309, 16'd26995, 16'd269, 16'd40056, 16'd3955, 16'd60365, 16'd24110, 16'd50793, 16'd44413, 16'd16919, 16'd45799, 16'd61007, 16'd48696, 16'd56696, 16'd3850, 16'd29082, 16'd26712, 16'd31985, 16'd24271, 16'd59522, 16'd3517, 16'd48325, 16'd31417});
	test_expansion(128'h41fb8aa70f24af2d1170c02f9ecc0c7e, {16'd30154, 16'd29253, 16'd35074, 16'd3086, 16'd17893, 16'd37029, 16'd51934, 16'd29328, 16'd13323, 16'd53001, 16'd35301, 16'd61283, 16'd52761, 16'd17168, 16'd9009, 16'd57374, 16'd38950, 16'd33409, 16'd34488, 16'd1951, 16'd57906, 16'd56358, 16'd4486, 16'd39633, 16'd40583, 16'd3280});
	test_expansion(128'h45f841e07204722e315e3b7d56cdf26d, {16'd16357, 16'd36111, 16'd13593, 16'd65091, 16'd8118, 16'd15733, 16'd34444, 16'd58046, 16'd53959, 16'd45070, 16'd20409, 16'd15627, 16'd64699, 16'd23783, 16'd42104, 16'd32631, 16'd26101, 16'd45231, 16'd5264, 16'd31065, 16'd46644, 16'd50641, 16'd44428, 16'd45286, 16'd30830, 16'd48331});
	test_expansion(128'h8e5909be538f0ab281ca6c98ade974c3, {16'd852, 16'd16924, 16'd38822, 16'd54012, 16'd13526, 16'd27445, 16'd31286, 16'd50674, 16'd18028, 16'd56673, 16'd28508, 16'd31316, 16'd10772, 16'd4074, 16'd48586, 16'd63027, 16'd13541, 16'd35589, 16'd56025, 16'd36465, 16'd60412, 16'd18748, 16'd40595, 16'd45037, 16'd40507, 16'd64434});
	test_expansion(128'h03dbbab4640c064d9cf7a837d7bbcce5, {16'd28575, 16'd46263, 16'd9144, 16'd41048, 16'd58452, 16'd56167, 16'd38250, 16'd24261, 16'd140, 16'd43368, 16'd11565, 16'd50849, 16'd53110, 16'd65169, 16'd43243, 16'd43093, 16'd25627, 16'd57548, 16'd49841, 16'd13232, 16'd17652, 16'd42755, 16'd10584, 16'd14126, 16'd708, 16'd34329});
	test_expansion(128'h4d4faa4c2b8ad96dfa3ef70ebcae1f66, {16'd38437, 16'd59254, 16'd50533, 16'd16994, 16'd5173, 16'd60480, 16'd1155, 16'd27385, 16'd57172, 16'd17623, 16'd39956, 16'd27951, 16'd40107, 16'd46987, 16'd29793, 16'd13535, 16'd27226, 16'd47167, 16'd21631, 16'd10355, 16'd52226, 16'd30670, 16'd26528, 16'd14993, 16'd55073, 16'd53500});
	test_expansion(128'h46db3f53c03010a22a3d24b766e0fabe, {16'd37175, 16'd27515, 16'd50316, 16'd30859, 16'd31913, 16'd8425, 16'd4094, 16'd1356, 16'd54656, 16'd45563, 16'd7621, 16'd50665, 16'd49217, 16'd42551, 16'd19307, 16'd38974, 16'd26881, 16'd9120, 16'd10413, 16'd64816, 16'd35528, 16'd629, 16'd1390, 16'd35066, 16'd55057, 16'd29253});
	test_expansion(128'hc5683567ac9b3f5afe0952cdfd2f2159, {16'd26672, 16'd15430, 16'd64502, 16'd36375, 16'd40821, 16'd12060, 16'd1332, 16'd28484, 16'd41957, 16'd7448, 16'd34483, 16'd19242, 16'd24945, 16'd41857, 16'd44076, 16'd20599, 16'd36263, 16'd21766, 16'd52956, 16'd36974, 16'd13081, 16'd46982, 16'd25056, 16'd56822, 16'd22006, 16'd13264});
	test_expansion(128'ha697cfabeecd7fe288d492156c18966f, {16'd34604, 16'd10086, 16'd64085, 16'd45883, 16'd17628, 16'd32707, 16'd60426, 16'd41738, 16'd1661, 16'd49741, 16'd48715, 16'd31987, 16'd63279, 16'd33821, 16'd37675, 16'd52044, 16'd63287, 16'd48047, 16'd6836, 16'd32098, 16'd40838, 16'd13853, 16'd48420, 16'd14241, 16'd49708, 16'd3296});
	test_expansion(128'h8295face35e6175ead045d35279eb35f, {16'd25914, 16'd19945, 16'd17069, 16'd26038, 16'd51252, 16'd56991, 16'd14841, 16'd61210, 16'd2183, 16'd23424, 16'd30478, 16'd34585, 16'd34827, 16'd39671, 16'd8237, 16'd47956, 16'd2984, 16'd55900, 16'd30748, 16'd64675, 16'd42659, 16'd51667, 16'd197, 16'd61264, 16'd43789, 16'd37122});
	test_expansion(128'h0953b5727b53004701a54a4c5ed7f7da, {16'd33110, 16'd26344, 16'd29902, 16'd28874, 16'd51193, 16'd10953, 16'd47320, 16'd33855, 16'd35430, 16'd20967, 16'd40613, 16'd30356, 16'd29277, 16'd16527, 16'd41403, 16'd43777, 16'd21931, 16'd26348, 16'd64502, 16'd11636, 16'd64101, 16'd48004, 16'd4008, 16'd50358, 16'd62756, 16'd549});
	test_expansion(128'h496bab014cbecaaa05c0c1f8594756c8, {16'd52571, 16'd30838, 16'd13349, 16'd12405, 16'd39589, 16'd60217, 16'd56634, 16'd2979, 16'd43204, 16'd27243, 16'd45652, 16'd52874, 16'd11367, 16'd15083, 16'd44576, 16'd62719, 16'd37008, 16'd56133, 16'd61326, 16'd11507, 16'd28607, 16'd31915, 16'd32554, 16'd32886, 16'd13355, 16'd63212});
	test_expansion(128'h35152d3fd3385a267508130ba29798b5, {16'd46074, 16'd10532, 16'd38622, 16'd13673, 16'd47541, 16'd5943, 16'd64687, 16'd21122, 16'd58136, 16'd24731, 16'd36947, 16'd2657, 16'd65369, 16'd17359, 16'd11429, 16'd11039, 16'd30723, 16'd63421, 16'd63017, 16'd56264, 16'd41042, 16'd14166, 16'd60394, 16'd4809, 16'd43539, 16'd20809});
	test_expansion(128'h8f2ff023da31dd8b091e0fb9ac7fe6cf, {16'd43508, 16'd55075, 16'd21679, 16'd47326, 16'd61939, 16'd26512, 16'd18418, 16'd25339, 16'd65116, 16'd35714, 16'd49370, 16'd26487, 16'd1867, 16'd26064, 16'd22592, 16'd41515, 16'd13316, 16'd51744, 16'd53021, 16'd20571, 16'd39582, 16'd2336, 16'd42132, 16'd45223, 16'd23696, 16'd43741});
	test_expansion(128'ha965295c1a64d400c5a0a776092fdbb0, {16'd336, 16'd38056, 16'd13368, 16'd31869, 16'd32127, 16'd1215, 16'd26068, 16'd35740, 16'd35382, 16'd16746, 16'd31616, 16'd29740, 16'd64481, 16'd2048, 16'd38648, 16'd56546, 16'd43402, 16'd50016, 16'd25049, 16'd65259, 16'd23879, 16'd56002, 16'd16442, 16'd1096, 16'd11162, 16'd14698});
	test_expansion(128'h0f3057ce1f33bc94d4bfd93ea4efafb6, {16'd20069, 16'd7259, 16'd47437, 16'd30791, 16'd40922, 16'd25092, 16'd51475, 16'd56567, 16'd48079, 16'd22016, 16'd12462, 16'd21421, 16'd47661, 16'd8969, 16'd26735, 16'd63466, 16'd20313, 16'd4678, 16'd63093, 16'd28638, 16'd41232, 16'd15352, 16'd9949, 16'd41765, 16'd4469, 16'd50175});
	test_expansion(128'h9e0d69f22c4a7e8c3d9e42439a7aa3ab, {16'd20548, 16'd32263, 16'd20499, 16'd4841, 16'd33737, 16'd42240, 16'd20104, 16'd33798, 16'd27281, 16'd55717, 16'd20008, 16'd5024, 16'd62935, 16'd59285, 16'd3377, 16'd22942, 16'd29148, 16'd1584, 16'd24940, 16'd34321, 16'd20039, 16'd33386, 16'd44418, 16'd14685, 16'd51605, 16'd63203});
	test_expansion(128'h4feca371e46d082b8c6eeb1103e4994c, {16'd46415, 16'd40586, 16'd55460, 16'd6193, 16'd11858, 16'd31621, 16'd58473, 16'd30555, 16'd806, 16'd51875, 16'd46209, 16'd36516, 16'd37788, 16'd64323, 16'd15164, 16'd12962, 16'd26147, 16'd28053, 16'd48019, 16'd1767, 16'd55306, 16'd50295, 16'd3098, 16'd12768, 16'd16355, 16'd58239});
	test_expansion(128'h4c8698fdc9618726bce963bd82b74f1a, {16'd35163, 16'd63108, 16'd3829, 16'd23243, 16'd6981, 16'd35922, 16'd4776, 16'd29954, 16'd15868, 16'd28175, 16'd18277, 16'd20713, 16'd17003, 16'd54457, 16'd43009, 16'd31925, 16'd14749, 16'd51626, 16'd63027, 16'd20657, 16'd15411, 16'd39891, 16'd24092, 16'd30615, 16'd62625, 16'd39513});
	test_expansion(128'h0262c68f1081833d52e68f25c647ffc1, {16'd2819, 16'd13570, 16'd43289, 16'd1340, 16'd52361, 16'd59050, 16'd911, 16'd37341, 16'd63231, 16'd65276, 16'd48111, 16'd28307, 16'd21630, 16'd7099, 16'd17317, 16'd42508, 16'd29589, 16'd22119, 16'd29788, 16'd46102, 16'd10223, 16'd63040, 16'd62624, 16'd1665, 16'd54305, 16'd34602});
	test_expansion(128'heee508ee43573dd55414373f2b5d6ca0, {16'd7025, 16'd63398, 16'd20897, 16'd17482, 16'd31453, 16'd10247, 16'd25984, 16'd58300, 16'd18441, 16'd36336, 16'd60151, 16'd28998, 16'd60322, 16'd24805, 16'd32667, 16'd7414, 16'd30158, 16'd62662, 16'd48621, 16'd53078, 16'd44968, 16'd23114, 16'd34643, 16'd20719, 16'd49320, 16'd12555});
	test_expansion(128'hdf06dc845d946833c197e9943c5b1719, {16'd8669, 16'd44725, 16'd12738, 16'd54364, 16'd51969, 16'd51105, 16'd25997, 16'd7659, 16'd299, 16'd22467, 16'd64336, 16'd874, 16'd55000, 16'd33094, 16'd7468, 16'd36716, 16'd43007, 16'd64662, 16'd30853, 16'd16586, 16'd49220, 16'd10380, 16'd58825, 16'd47669, 16'd26495, 16'd50058});
	test_expansion(128'h3f913fb1cc907478b66ae408f18a19ce, {16'd26457, 16'd64695, 16'd2803, 16'd64994, 16'd46232, 16'd58338, 16'd50234, 16'd37112, 16'd47274, 16'd57697, 16'd47106, 16'd34192, 16'd31403, 16'd44573, 16'd28835, 16'd20445, 16'd41311, 16'd14970, 16'd39217, 16'd41907, 16'd44684, 16'd976, 16'd15822, 16'd1390, 16'd16907, 16'd15851});
	test_expansion(128'hd34b3f9b2cbf2381b5180d1ea1c005ed, {16'd35469, 16'd41624, 16'd26706, 16'd6842, 16'd8789, 16'd24807, 16'd27518, 16'd8798, 16'd43928, 16'd38868, 16'd11776, 16'd981, 16'd17298, 16'd53394, 16'd8092, 16'd53240, 16'd13206, 16'd24419, 16'd18784, 16'd51961, 16'd33081, 16'd23893, 16'd18878, 16'd20916, 16'd20897, 16'd27096});
	test_expansion(128'h367b14c851b4aa2c5764c37c473ec6d5, {16'd8426, 16'd13523, 16'd36882, 16'd64796, 16'd5936, 16'd39582, 16'd48336, 16'd34862, 16'd24272, 16'd259, 16'd1649, 16'd52859, 16'd51462, 16'd33959, 16'd41905, 16'd21026, 16'd61298, 16'd6775, 16'd63015, 16'd36351, 16'd39059, 16'd44582, 16'd40291, 16'd14385, 16'd28919, 16'd40678});
	test_expansion(128'hf89b210db0c0e2b167f004edadfd2631, {16'd64317, 16'd8701, 16'd24152, 16'd63697, 16'd18859, 16'd261, 16'd48043, 16'd65196, 16'd25520, 16'd13232, 16'd9012, 16'd55366, 16'd36910, 16'd1461, 16'd26841, 16'd33254, 16'd12053, 16'd12007, 16'd29115, 16'd37685, 16'd56288, 16'd4236, 16'd37523, 16'd15735, 16'd44946, 16'd60573});
	test_expansion(128'h2d3c20ba5a0ae4d35fdda35e3bf82ab7, {16'd50881, 16'd17046, 16'd23087, 16'd7288, 16'd32582, 16'd65144, 16'd17982, 16'd6402, 16'd45222, 16'd3695, 16'd21183, 16'd52275, 16'd27191, 16'd38457, 16'd14069, 16'd61897, 16'd27992, 16'd1832, 16'd53539, 16'd57901, 16'd46583, 16'd7848, 16'd9299, 16'd24647, 16'd60449, 16'd14345});
	test_expansion(128'h9e40f44c6d8eba3ed433df5787a3538a, {16'd12313, 16'd47735, 16'd64957, 16'd42968, 16'd37104, 16'd44603, 16'd24636, 16'd11609, 16'd16770, 16'd17659, 16'd46696, 16'd40959, 16'd46925, 16'd13365, 16'd56663, 16'd46005, 16'd45239, 16'd55670, 16'd62396, 16'd29960, 16'd22818, 16'd5666, 16'd4768, 16'd28544, 16'd21132, 16'd31035});
	test_expansion(128'h5d20f77fa0788f4fe7abc94cd59228e6, {16'd39570, 16'd9089, 16'd1911, 16'd39795, 16'd6973, 16'd21252, 16'd1489, 16'd23005, 16'd52036, 16'd60616, 16'd49068, 16'd32442, 16'd26897, 16'd43851, 16'd39676, 16'd55453, 16'd8161, 16'd6979, 16'd58548, 16'd62749, 16'd64636, 16'd12095, 16'd17157, 16'd35759, 16'd7127, 16'd38655});
	test_expansion(128'h267567d1a8df3d4b326d4a5d4e2d474a, {16'd25281, 16'd30645, 16'd25148, 16'd2028, 16'd9730, 16'd45714, 16'd57753, 16'd45671, 16'd15271, 16'd63503, 16'd14910, 16'd42920, 16'd10251, 16'd22093, 16'd11618, 16'd20016, 16'd8697, 16'd18847, 16'd22315, 16'd9425, 16'd63948, 16'd50699, 16'd27043, 16'd14231, 16'd48617, 16'd27176});
	test_expansion(128'h94c3008c2f624089ea63ada638530f1b, {16'd21428, 16'd44908, 16'd15311, 16'd31916, 16'd61460, 16'd36300, 16'd9886, 16'd31373, 16'd14981, 16'd33062, 16'd9858, 16'd52136, 16'd35005, 16'd64461, 16'd52447, 16'd30724, 16'd16046, 16'd64190, 16'd17814, 16'd39277, 16'd46487, 16'd49959, 16'd11976, 16'd22122, 16'd2673, 16'd6581});
	test_expansion(128'h6aa8ac7527288ce7acd8159b7bd827a2, {16'd28448, 16'd57389, 16'd22311, 16'd64908, 16'd43068, 16'd30465, 16'd23580, 16'd35545, 16'd56662, 16'd32445, 16'd12719, 16'd17236, 16'd54114, 16'd40493, 16'd17842, 16'd47272, 16'd9172, 16'd41414, 16'd16667, 16'd32369, 16'd62146, 16'd21543, 16'd55646, 16'd44799, 16'd5867, 16'd14023});
	test_expansion(128'hcc422de5906454621e1ee53a20b2a33b, {16'd45321, 16'd18408, 16'd45743, 16'd2583, 16'd48355, 16'd32140, 16'd11429, 16'd47277, 16'd35057, 16'd50334, 16'd17810, 16'd26607, 16'd45063, 16'd12919, 16'd24968, 16'd32474, 16'd21315, 16'd37169, 16'd14441, 16'd3501, 16'd8862, 16'd19407, 16'd38531, 16'd42456, 16'd49843, 16'd19646});
	test_expansion(128'h4e7034c7ea319269325e2cbfdd5ce236, {16'd17477, 16'd2770, 16'd1411, 16'd12986, 16'd21051, 16'd33105, 16'd56571, 16'd7528, 16'd62982, 16'd738, 16'd3160, 16'd31174, 16'd25998, 16'd62594, 16'd9713, 16'd20414, 16'd41166, 16'd63794, 16'd21188, 16'd10032, 16'd19573, 16'd60144, 16'd61353, 16'd41198, 16'd39001, 16'd38951});
	test_expansion(128'h4fb4b6b7ac8e5286075e8348beccb3d7, {16'd54278, 16'd8327, 16'd8971, 16'd49102, 16'd48171, 16'd18801, 16'd16104, 16'd58621, 16'd61237, 16'd26661, 16'd43469, 16'd16077, 16'd60858, 16'd27426, 16'd22996, 16'd36714, 16'd47783, 16'd15020, 16'd57727, 16'd31146, 16'd37852, 16'd14870, 16'd28524, 16'd10659, 16'd2663, 16'd5250});
	test_expansion(128'h620183f3e2d1b3181faf1dfce181aba6, {16'd52829, 16'd3588, 16'd43274, 16'd20498, 16'd14578, 16'd58235, 16'd27001, 16'd2308, 16'd51463, 16'd10216, 16'd51739, 16'd41531, 16'd8558, 16'd31555, 16'd41046, 16'd34497, 16'd1002, 16'd24317, 16'd48223, 16'd17853, 16'd45771, 16'd44793, 16'd11716, 16'd7886, 16'd58992, 16'd22314});
	test_expansion(128'h9a8f2e25f390241bcd7b2082e83eae1a, {16'd17715, 16'd30291, 16'd10523, 16'd41057, 16'd40037, 16'd14669, 16'd50436, 16'd39414, 16'd52451, 16'd1990, 16'd18749, 16'd30646, 16'd23375, 16'd13919, 16'd27564, 16'd26104, 16'd17848, 16'd22228, 16'd36814, 16'd64999, 16'd37273, 16'd56852, 16'd7782, 16'd13651, 16'd27155, 16'd189});
	test_expansion(128'h9feab3c4fdd1ab5a145f170f16dd3ebc, {16'd55672, 16'd62369, 16'd41508, 16'd30657, 16'd4490, 16'd50715, 16'd18520, 16'd944, 16'd33856, 16'd15808, 16'd12478, 16'd23664, 16'd51495, 16'd25740, 16'd54237, 16'd32705, 16'd4552, 16'd47896, 16'd49258, 16'd6058, 16'd41433, 16'd45763, 16'd43201, 16'd2475, 16'd12549, 16'd19971});
	test_expansion(128'h20fdf802a0693469abcb10cf55705b8f, {16'd33426, 16'd4094, 16'd34237, 16'd24436, 16'd2974, 16'd22792, 16'd45913, 16'd9138, 16'd2369, 16'd34, 16'd56254, 16'd31371, 16'd10100, 16'd24500, 16'd40458, 16'd65208, 16'd11020, 16'd43500, 16'd5623, 16'd14750, 16'd8974, 16'd5489, 16'd28141, 16'd1487, 16'd58581, 16'd44894});
	test_expansion(128'h42260c16d96dc8b5e0c8e0d9e5fea762, {16'd22236, 16'd48260, 16'd51731, 16'd60981, 16'd2234, 16'd62467, 16'd12406, 16'd1305, 16'd37609, 16'd51293, 16'd31318, 16'd58302, 16'd7608, 16'd21439, 16'd24437, 16'd54123, 16'd29605, 16'd19185, 16'd15062, 16'd41403, 16'd35135, 16'd40892, 16'd36757, 16'd56186, 16'd14411, 16'd61349});
	test_expansion(128'he4496e3f0d1239ae14acd323d195e6a7, {16'd12646, 16'd52113, 16'd26468, 16'd63789, 16'd28214, 16'd42874, 16'd22242, 16'd1772, 16'd19432, 16'd23852, 16'd44152, 16'd7275, 16'd11954, 16'd24706, 16'd54428, 16'd25161, 16'd63865, 16'd6582, 16'd63936, 16'd14422, 16'd8859, 16'd4549, 16'd27591, 16'd35386, 16'd55604, 16'd25780});
	test_expansion(128'h9af902d02a8434207048cd8b31eb81be, {16'd62121, 16'd8387, 16'd26643, 16'd1873, 16'd31074, 16'd7206, 16'd7734, 16'd13303, 16'd11116, 16'd36895, 16'd24263, 16'd35832, 16'd25843, 16'd53708, 16'd323, 16'd48466, 16'd21722, 16'd34139, 16'd48049, 16'd2537, 16'd28844, 16'd20635, 16'd25857, 16'd64339, 16'd21034, 16'd3067});
	test_expansion(128'hb9571e96b72ae7f33270f1a1ca428ee6, {16'd623, 16'd64379, 16'd49623, 16'd43960, 16'd38019, 16'd58002, 16'd32025, 16'd20162, 16'd18527, 16'd7968, 16'd12816, 16'd9751, 16'd24299, 16'd42802, 16'd26106, 16'd24801, 16'd12949, 16'd64193, 16'd25146, 16'd60992, 16'd24123, 16'd37989, 16'd43106, 16'd43204, 16'd36943, 16'd20714});
	test_expansion(128'h4dcbd2190aec5b091cbd85d184900eae, {16'd7170, 16'd3749, 16'd16308, 16'd3043, 16'd5459, 16'd27764, 16'd24160, 16'd36023, 16'd29448, 16'd26188, 16'd48331, 16'd4932, 16'd61477, 16'd52793, 16'd55796, 16'd41641, 16'd14998, 16'd31274, 16'd58966, 16'd1646, 16'd64405, 16'd1235, 16'd26089, 16'd16123, 16'd10372, 16'd29196});
	test_expansion(128'ha0bb27a5ed7efcc0513a419f81dd2621, {16'd2582, 16'd55022, 16'd29514, 16'd686, 16'd32242, 16'd4982, 16'd32016, 16'd28490, 16'd55700, 16'd57440, 16'd21454, 16'd60625, 16'd49032, 16'd56394, 16'd36348, 16'd39236, 16'd27425, 16'd4535, 16'd59926, 16'd3855, 16'd32705, 16'd5200, 16'd18271, 16'd3752, 16'd54673, 16'd3102});
	test_expansion(128'h2aa0b52933bcd45a5bed6cbd40183a04, {16'd7345, 16'd27700, 16'd39605, 16'd14875, 16'd39238, 16'd48684, 16'd37962, 16'd57792, 16'd5865, 16'd53649, 16'd60519, 16'd45302, 16'd7227, 16'd27649, 16'd31319, 16'd46137, 16'd31152, 16'd56282, 16'd48691, 16'd1794, 16'd41410, 16'd3144, 16'd13738, 16'd10308, 16'd9538, 16'd25422});
	test_expansion(128'hc0fcbef50ea6ecdd5b14b65fdaef1970, {16'd7027, 16'd33544, 16'd28358, 16'd61791, 16'd46757, 16'd56870, 16'd64055, 16'd13807, 16'd44406, 16'd48875, 16'd17609, 16'd53119, 16'd19360, 16'd38824, 16'd29520, 16'd36225, 16'd53259, 16'd31331, 16'd37063, 16'd61541, 16'd33111, 16'd44602, 16'd56821, 16'd38667, 16'd11542, 16'd59530});
	test_expansion(128'h7f397c999e431a7afd87d2e2633cb136, {16'd50476, 16'd27266, 16'd22201, 16'd29901, 16'd49932, 16'd36549, 16'd6599, 16'd20930, 16'd61629, 16'd29223, 16'd57678, 16'd48305, 16'd37459, 16'd62729, 16'd6056, 16'd55206, 16'd19438, 16'd16622, 16'd40280, 16'd41557, 16'd16415, 16'd63915, 16'd28155, 16'd42286, 16'd42391, 16'd64490});
	test_expansion(128'h9354619758d156e9b11d852a73072b9f, {16'd30970, 16'd53057, 16'd36699, 16'd43722, 16'd22795, 16'd31661, 16'd40518, 16'd42479, 16'd6719, 16'd7859, 16'd36179, 16'd7505, 16'd8754, 16'd60668, 16'd42100, 16'd15898, 16'd63130, 16'd37063, 16'd10254, 16'd52633, 16'd9169, 16'd52691, 16'd51013, 16'd47266, 16'd19684, 16'd61851});
	test_expansion(128'h9bb2ed977ec2f96f3578ad94d898aa07, {16'd18554, 16'd33501, 16'd8360, 16'd8111, 16'd13268, 16'd40127, 16'd38368, 16'd19673, 16'd48101, 16'd14673, 16'd3392, 16'd1757, 16'd53409, 16'd25960, 16'd48961, 16'd62492, 16'd44608, 16'd28791, 16'd63057, 16'd27621, 16'd54975, 16'd2648, 16'd54623, 16'd50881, 16'd9204, 16'd28588});
	test_expansion(128'h365b02b3c95e3efb809da64c0bacc115, {16'd47838, 16'd27751, 16'd39187, 16'd52538, 16'd16983, 16'd48938, 16'd35547, 16'd5132, 16'd36447, 16'd8194, 16'd33436, 16'd22452, 16'd22885, 16'd63991, 16'd230, 16'd44058, 16'd47473, 16'd12889, 16'd28211, 16'd59540, 16'd53079, 16'd53088, 16'd57094, 16'd9463, 16'd6209, 16'd13867});
	test_expansion(128'hb14d99fb03610e36a84b388914cbd136, {16'd42962, 16'd32940, 16'd58407, 16'd41887, 16'd7471, 16'd55150, 16'd44193, 16'd40615, 16'd27725, 16'd49571, 16'd14381, 16'd32937, 16'd33100, 16'd16127, 16'd45235, 16'd32149, 16'd64715, 16'd8411, 16'd58919, 16'd594, 16'd52068, 16'd51626, 16'd62358, 16'd45038, 16'd64402, 16'd1909});
	test_expansion(128'h11dc773e513b08d4264147cc828edb51, {16'd17125, 16'd54012, 16'd13207, 16'd38978, 16'd45406, 16'd37053, 16'd13476, 16'd4776, 16'd16794, 16'd56547, 16'd40834, 16'd5580, 16'd38291, 16'd14394, 16'd44781, 16'd41272, 16'd2006, 16'd24352, 16'd8649, 16'd42074, 16'd5858, 16'd29581, 16'd54834, 16'd33331, 16'd4120, 16'd15193});
	test_expansion(128'h7cad93553997679e145eeb701935e73c, {16'd6946, 16'd24671, 16'd35465, 16'd63297, 16'd24982, 16'd57155, 16'd43395, 16'd30443, 16'd61841, 16'd53095, 16'd19653, 16'd17824, 16'd50112, 16'd56873, 16'd19044, 16'd26828, 16'd47022, 16'd1678, 16'd17607, 16'd54072, 16'd51964, 16'd45378, 16'd30397, 16'd23562, 16'd41856, 16'd49070});
	test_expansion(128'hd019f8d07882a56b81ee1b25103a8ca1, {16'd10434, 16'd45232, 16'd39098, 16'd44527, 16'd62066, 16'd52989, 16'd6779, 16'd40768, 16'd30637, 16'd50651, 16'd60356, 16'd25677, 16'd22371, 16'd49022, 16'd6270, 16'd62075, 16'd18555, 16'd5290, 16'd18020, 16'd51934, 16'd27411, 16'd52812, 16'd27459, 16'd39514, 16'd43609, 16'd46807});
	test_expansion(128'hf0df3a46e9b2057345a9f1d288e4e32f, {16'd61868, 16'd45665, 16'd3739, 16'd22610, 16'd51346, 16'd6979, 16'd65440, 16'd54825, 16'd41111, 16'd31408, 16'd20210, 16'd29607, 16'd23270, 16'd20813, 16'd56381, 16'd48094, 16'd31147, 16'd60401, 16'd52166, 16'd50907, 16'd29683, 16'd21424, 16'd22343, 16'd5339, 16'd65413, 16'd21923});
	test_expansion(128'hf5a4711d0002b4de5d1114442c6265b0, {16'd31493, 16'd13324, 16'd23019, 16'd37993, 16'd25178, 16'd34920, 16'd217, 16'd17424, 16'd13896, 16'd34031, 16'd25807, 16'd20953, 16'd7072, 16'd53114, 16'd21912, 16'd14318, 16'd51513, 16'd30390, 16'd63845, 16'd47345, 16'd49204, 16'd41999, 16'd25918, 16'd51491, 16'd49201, 16'd34874});
	test_expansion(128'h4df573d2ec20a71f3593f2ee8d66a7ba, {16'd35445, 16'd64313, 16'd61759, 16'd26577, 16'd16775, 16'd17721, 16'd41642, 16'd63220, 16'd34978, 16'd2873, 16'd54588, 16'd34624, 16'd4860, 16'd21131, 16'd3651, 16'd18773, 16'd16834, 16'd50662, 16'd25867, 16'd59860, 16'd18057, 16'd17815, 16'd7691, 16'd8845, 16'd63413, 16'd25982});
	test_expansion(128'h5dc5cd4faa9ac37f7f3e72ee07d5a0cd, {16'd5071, 16'd41817, 16'd18178, 16'd4700, 16'd8476, 16'd61983, 16'd30601, 16'd26448, 16'd40279, 16'd40211, 16'd52177, 16'd38246, 16'd57192, 16'd39608, 16'd34032, 16'd35397, 16'd58205, 16'd33845, 16'd39796, 16'd37407, 16'd26477, 16'd53874, 16'd45238, 16'd38703, 16'd2657, 16'd49078});
	test_expansion(128'h52ca3e0415ff27d9f6582640bc0e7577, {16'd56963, 16'd27752, 16'd28146, 16'd9615, 16'd44546, 16'd52275, 16'd6876, 16'd4410, 16'd49751, 16'd17497, 16'd14018, 16'd27491, 16'd29894, 16'd8686, 16'd20705, 16'd55618, 16'd36339, 16'd50143, 16'd22092, 16'd21395, 16'd4182, 16'd18740, 16'd44713, 16'd65179, 16'd49646, 16'd4941});
	test_expansion(128'hba7eaaf8a2ecb80f9b17c7010e2b937a, {16'd34240, 16'd43654, 16'd17306, 16'd4077, 16'd31376, 16'd18141, 16'd38945, 16'd40149, 16'd59948, 16'd46719, 16'd38528, 16'd50389, 16'd24776, 16'd17960, 16'd63302, 16'd39155, 16'd20865, 16'd3590, 16'd57007, 16'd51658, 16'd519, 16'd36714, 16'd7015, 16'd56891, 16'd1853, 16'd34023});
	test_expansion(128'h27ce13944c3b24059cde536832a1e158, {16'd52104, 16'd11687, 16'd59347, 16'd37059, 16'd17380, 16'd38069, 16'd34833, 16'd1998, 16'd62599, 16'd60672, 16'd25671, 16'd16380, 16'd48453, 16'd18790, 16'd15611, 16'd20061, 16'd46670, 16'd9115, 16'd45470, 16'd11081, 16'd8578, 16'd63810, 16'd51448, 16'd17129, 16'd47499, 16'd22271});
	test_expansion(128'h3b3cb0a29f0fe4a3360cd84e3f16c18e, {16'd39416, 16'd14028, 16'd65411, 16'd20469, 16'd24883, 16'd14552, 16'd53046, 16'd30530, 16'd40995, 16'd1921, 16'd27044, 16'd37606, 16'd59411, 16'd5550, 16'd65106, 16'd42612, 16'd9336, 16'd6906, 16'd44430, 16'd52921, 16'd34839, 16'd7392, 16'd26667, 16'd99, 16'd21878, 16'd2066});
	test_expansion(128'h840172a3b7eb934f3662231beb05b7ae, {16'd34998, 16'd32839, 16'd34800, 16'd35311, 16'd50408, 16'd21978, 16'd55649, 16'd25039, 16'd412, 16'd24249, 16'd7343, 16'd30433, 16'd10677, 16'd57917, 16'd59, 16'd18563, 16'd26952, 16'd26332, 16'd24514, 16'd4764, 16'd27251, 16'd44911, 16'd48757, 16'd28997, 16'd22287, 16'd19994});
	test_expansion(128'h900883f6352f959985825bb146b200b7, {16'd32109, 16'd47758, 16'd29470, 16'd26226, 16'd46056, 16'd30058, 16'd16745, 16'd59365, 16'd48806, 16'd60494, 16'd59891, 16'd22012, 16'd56307, 16'd48988, 16'd17225, 16'd52274, 16'd12748, 16'd11236, 16'd27918, 16'd44649, 16'd28820, 16'd3763, 16'd45155, 16'd250, 16'd5233, 16'd10246});
	test_expansion(128'hc0b24b6eb01c68fa994e9ff982c07ac3, {16'd59220, 16'd27245, 16'd10033, 16'd56790, 16'd31657, 16'd4804, 16'd44784, 16'd8849, 16'd32744, 16'd539, 16'd15174, 16'd50276, 16'd2659, 16'd11735, 16'd36559, 16'd63295, 16'd8638, 16'd41763, 16'd37818, 16'd33348, 16'd1671, 16'd21802, 16'd41468, 16'd39423, 16'd13018, 16'd23141});
	test_expansion(128'h1377ae2ce62455145d9306a7d36ae5c2, {16'd39926, 16'd1442, 16'd4096, 16'd1903, 16'd63987, 16'd50186, 16'd29708, 16'd10649, 16'd14040, 16'd40145, 16'd52613, 16'd20358, 16'd52825, 16'd55222, 16'd60498, 16'd13340, 16'd35205, 16'd8533, 16'd49688, 16'd17828, 16'd4831, 16'd54884, 16'd59835, 16'd30078, 16'd21022, 16'd28087});
	test_expansion(128'h2665751cdc07d1dfd9807b94e1b91d5b, {16'd604, 16'd9703, 16'd40001, 16'd14035, 16'd64472, 16'd62207, 16'd37024, 16'd10001, 16'd30283, 16'd54752, 16'd57106, 16'd17233, 16'd17417, 16'd47133, 16'd56238, 16'd55602, 16'd48868, 16'd52893, 16'd1490, 16'd31836, 16'd57062, 16'd62199, 16'd999, 16'd30766, 16'd65261, 16'd29721});
	test_expansion(128'h06c0e6c8fce2a8e8516de15d003ecc48, {16'd58927, 16'd41160, 16'd23346, 16'd12730, 16'd10664, 16'd15938, 16'd57095, 16'd44028, 16'd56762, 16'd4264, 16'd5152, 16'd37859, 16'd1321, 16'd4003, 16'd24686, 16'd44781, 16'd11212, 16'd47041, 16'd15761, 16'd62622, 16'd42815, 16'd35396, 16'd47247, 16'd9098, 16'd53123, 16'd17800});
	test_expansion(128'h72993e5fd8656460072cf53d38d5c39d, {16'd32547, 16'd38538, 16'd29183, 16'd10509, 16'd2416, 16'd61966, 16'd12655, 16'd12836, 16'd47693, 16'd42900, 16'd32095, 16'd8260, 16'd24594, 16'd25799, 16'd47672, 16'd59599, 16'd62911, 16'd34181, 16'd19504, 16'd52617, 16'd40582, 16'd56840, 16'd60778, 16'd7620, 16'd53472, 16'd21058});
	test_expansion(128'h917364cf6bbb202a8a606f519fabbc5f, {16'd24661, 16'd21854, 16'd54178, 16'd62652, 16'd34785, 16'd59257, 16'd60056, 16'd54270, 16'd55593, 16'd34166, 16'd2879, 16'd48916, 16'd4297, 16'd16143, 16'd49592, 16'd6554, 16'd31210, 16'd19658, 16'd54165, 16'd2595, 16'd31785, 16'd55011, 16'd44278, 16'd53570, 16'd44473, 16'd40014});
	test_expansion(128'he229ab9b3d89695d27efe6aebcc9a6cb, {16'd17466, 16'd36209, 16'd33603, 16'd30493, 16'd6408, 16'd30278, 16'd32650, 16'd37629, 16'd47885, 16'd26663, 16'd19678, 16'd19416, 16'd41654, 16'd9129, 16'd28716, 16'd53752, 16'd32608, 16'd65001, 16'd32456, 16'd6168, 16'd61476, 16'd33265, 16'd14562, 16'd63144, 16'd3473, 16'd14369});
	test_expansion(128'h011f1ad6f48aae8cf4017d336e15b884, {16'd23132, 16'd38167, 16'd41500, 16'd42391, 16'd39573, 16'd50820, 16'd52459, 16'd27715, 16'd12130, 16'd20839, 16'd40132, 16'd64358, 16'd4086, 16'd27662, 16'd45659, 16'd61988, 16'd39534, 16'd1120, 16'd50937, 16'd37987, 16'd55033, 16'd65047, 16'd20315, 16'd39563, 16'd55493, 16'd46584});
	test_expansion(128'h920ebe5fa97406a34c1ba31031b14a8b, {16'd24645, 16'd11702, 16'd49818, 16'd667, 16'd5671, 16'd8315, 16'd13951, 16'd45661, 16'd30700, 16'd37788, 16'd32025, 16'd64464, 16'd5447, 16'd57351, 16'd12316, 16'd22676, 16'd36524, 16'd5246, 16'd27560, 16'd46989, 16'd35187, 16'd2100, 16'd949, 16'd49269, 16'd46669, 16'd53353});
	test_expansion(128'hee304d725f5b7e6251b947c218c30590, {16'd62604, 16'd11082, 16'd43943, 16'd32301, 16'd40448, 16'd61975, 16'd45724, 16'd53432, 16'd58288, 16'd21605, 16'd2831, 16'd49965, 16'd50587, 16'd38655, 16'd5618, 16'd20150, 16'd4563, 16'd32221, 16'd56931, 16'd16341, 16'd35752, 16'd44043, 16'd19012, 16'd38188, 16'd53449, 16'd9489});
	test_expansion(128'hcf0f5555062bf2097b6dbd584dab37d9, {16'd38456, 16'd22309, 16'd6583, 16'd9776, 16'd49778, 16'd11410, 16'd60451, 16'd54347, 16'd5165, 16'd49594, 16'd40633, 16'd28988, 16'd59463, 16'd2203, 16'd55353, 16'd11049, 16'd12626, 16'd57288, 16'd20702, 16'd9518, 16'd50295, 16'd31607, 16'd41721, 16'd60898, 16'd33531, 16'd22673});
	test_expansion(128'h5bda799c50571d6d4a3badb3f3a926fb, {16'd46429, 16'd60899, 16'd23119, 16'd45284, 16'd6372, 16'd18635, 16'd44893, 16'd35152, 16'd32948, 16'd1392, 16'd10950, 16'd60160, 16'd60949, 16'd59589, 16'd43195, 16'd57376, 16'd2349, 16'd48264, 16'd60471, 16'd62757, 16'd59104, 16'd11425, 16'd20722, 16'd38429, 16'd11332, 16'd2002});
	test_expansion(128'h120c4e6fafcf6f75437d3b5aba451a98, {16'd2852, 16'd1124, 16'd32428, 16'd5860, 16'd56456, 16'd28545, 16'd49816, 16'd30175, 16'd18429, 16'd43412, 16'd11002, 16'd19809, 16'd48190, 16'd33550, 16'd57515, 16'd43106, 16'd63230, 16'd51480, 16'd44828, 16'd33534, 16'd17190, 16'd39082, 16'd34832, 16'd11749, 16'd44427, 16'd44084});
	test_expansion(128'hab501f7d1283b8f7528d214086ba542f, {16'd56734, 16'd45598, 16'd52278, 16'd11817, 16'd15968, 16'd4720, 16'd36857, 16'd26898, 16'd62796, 16'd3512, 16'd40666, 16'd5614, 16'd56152, 16'd34666, 16'd21831, 16'd12378, 16'd28525, 16'd7992, 16'd18212, 16'd35236, 16'd49148, 16'd17416, 16'd17870, 16'd29907, 16'd50713, 16'd61542});
	test_expansion(128'h4c590122a39764606d87e2d18f4c2c7c, {16'd51941, 16'd48658, 16'd30236, 16'd59784, 16'd33264, 16'd45875, 16'd992, 16'd11157, 16'd39260, 16'd65403, 16'd64967, 16'd9728, 16'd9968, 16'd51505, 16'd44821, 16'd36728, 16'd2595, 16'd9322, 16'd59645, 16'd53145, 16'd19105, 16'd13218, 16'd17114, 16'd60309, 16'd23611, 16'd23038});
	test_expansion(128'h8d1f445eeedcfb42ec28da8e55862424, {16'd8717, 16'd17221, 16'd25760, 16'd14627, 16'd30441, 16'd46680, 16'd30314, 16'd12716, 16'd53511, 16'd47700, 16'd37889, 16'd49611, 16'd36933, 16'd24879, 16'd43985, 16'd21383, 16'd11042, 16'd38783, 16'd47452, 16'd1279, 16'd8101, 16'd41420, 16'd50310, 16'd53360, 16'd30997, 16'd35625});
	test_expansion(128'h3b5d77c6efe89573f8ff480c52f45f40, {16'd19050, 16'd36717, 16'd33524, 16'd30431, 16'd15961, 16'd39361, 16'd59903, 16'd30103, 16'd11593, 16'd46519, 16'd15538, 16'd9021, 16'd50869, 16'd45223, 16'd59558, 16'd41829, 16'd34011, 16'd28653, 16'd44901, 16'd5495, 16'd22010, 16'd22283, 16'd30929, 16'd45490, 16'd51707, 16'd2048});
	test_expansion(128'hfd51247c0dd295038646f90abc7e1ae5, {16'd3647, 16'd22678, 16'd19043, 16'd51435, 16'd27973, 16'd42009, 16'd59936, 16'd44738, 16'd6219, 16'd48236, 16'd43129, 16'd15480, 16'd7580, 16'd61231, 16'd9264, 16'd29102, 16'd35230, 16'd54043, 16'd27969, 16'd10699, 16'd33756, 16'd50061, 16'd30131, 16'd58680, 16'd9712, 16'd6090});
	test_expansion(128'ha262cd2a34836ff45b71245070ca6bf1, {16'd46073, 16'd13750, 16'd1719, 16'd17338, 16'd1558, 16'd15542, 16'd20509, 16'd20969, 16'd48975, 16'd37384, 16'd59411, 16'd13396, 16'd12943, 16'd32698, 16'd29222, 16'd31745, 16'd43265, 16'd20208, 16'd20617, 16'd34369, 16'd11847, 16'd23574, 16'd4225, 16'd42393, 16'd10101, 16'd63316});
	test_expansion(128'h7caa7253ae9edf9dfbd252af6d68ec51, {16'd64280, 16'd21430, 16'd57156, 16'd64703, 16'd27500, 16'd58765, 16'd32223, 16'd544, 16'd62376, 16'd14265, 16'd285, 16'd56220, 16'd56014, 16'd25729, 16'd65444, 16'd18204, 16'd48161, 16'd40369, 16'd1439, 16'd40215, 16'd4017, 16'd37782, 16'd8090, 16'd36211, 16'd25348, 16'd177});
	test_expansion(128'hbaa97005ef2721895593468f6e2e4eea, {16'd48099, 16'd44494, 16'd28851, 16'd46327, 16'd7144, 16'd39855, 16'd1829, 16'd30888, 16'd14500, 16'd34705, 16'd62284, 16'd62216, 16'd8978, 16'd53798, 16'd13933, 16'd57308, 16'd11518, 16'd23996, 16'd55280, 16'd30317, 16'd42193, 16'd50647, 16'd32335, 16'd24837, 16'd12694, 16'd46364});
	test_expansion(128'h7e0217885f211744815e1bbdd053e985, {16'd60638, 16'd4671, 16'd35676, 16'd34468, 16'd62414, 16'd62115, 16'd41424, 16'd32294, 16'd1459, 16'd61158, 16'd65306, 16'd18672, 16'd18049, 16'd4993, 16'd37634, 16'd40282, 16'd11272, 16'd58942, 16'd10779, 16'd41425, 16'd28140, 16'd24512, 16'd20304, 16'd2600, 16'd61514, 16'd54891});
	test_expansion(128'hd790f075aa60dbaaab9f7bca84f6c187, {16'd48257, 16'd55425, 16'd38656, 16'd34641, 16'd23623, 16'd350, 16'd36435, 16'd35018, 16'd45090, 16'd8213, 16'd6737, 16'd44600, 16'd19556, 16'd38008, 16'd54626, 16'd44968, 16'd57859, 16'd55871, 16'd55173, 16'd47748, 16'd34149, 16'd21714, 16'd53452, 16'd55631, 16'd32551, 16'd21547});
	test_expansion(128'h6db77d48a540c0a84dcfdf5960075c5d, {16'd8389, 16'd36343, 16'd54206, 16'd26865, 16'd37724, 16'd49662, 16'd11661, 16'd47273, 16'd10993, 16'd19349, 16'd46751, 16'd38397, 16'd32483, 16'd33735, 16'd26585, 16'd44437, 16'd20335, 16'd58634, 16'd60144, 16'd42928, 16'd7409, 16'd61834, 16'd28163, 16'd32607, 16'd24171, 16'd54854});
	test_expansion(128'heeedadf1349494466bd8437f66ef433f, {16'd65513, 16'd4810, 16'd3602, 16'd59138, 16'd29034, 16'd43927, 16'd41999, 16'd46535, 16'd9105, 16'd36816, 16'd18992, 16'd50718, 16'd61836, 16'd49787, 16'd15604, 16'd27040, 16'd26594, 16'd48522, 16'd59679, 16'd4236, 16'd27578, 16'd17068, 16'd52745, 16'd53960, 16'd64260, 16'd41165});
	test_expansion(128'h374ad536c92969d0666c6e980756db5e, {16'd42566, 16'd3371, 16'd5865, 16'd49361, 16'd23940, 16'd56010, 16'd61127, 16'd47954, 16'd63860, 16'd39834, 16'd60474, 16'd44859, 16'd41618, 16'd54580, 16'd19485, 16'd62341, 16'd11993, 16'd41119, 16'd21058, 16'd42105, 16'd46160, 16'd53346, 16'd35641, 16'd16531, 16'd5490, 16'd7621});
	test_expansion(128'h0992eda84b926f1ba62d5b6ede35741c, {16'd60627, 16'd27249, 16'd54879, 16'd42428, 16'd57564, 16'd1651, 16'd49711, 16'd6976, 16'd62775, 16'd58622, 16'd64456, 16'd8171, 16'd142, 16'd19092, 16'd2109, 16'd35188, 16'd31376, 16'd20607, 16'd32618, 16'd7998, 16'd14138, 16'd136, 16'd32021, 16'd38959, 16'd33754, 16'd7644});
	test_expansion(128'h8151c6769dd537ae32f240734b19bc83, {16'd37908, 16'd36010, 16'd55612, 16'd56364, 16'd24005, 16'd30814, 16'd14661, 16'd15445, 16'd24219, 16'd41236, 16'd25702, 16'd14599, 16'd52768, 16'd36054, 16'd53247, 16'd55053, 16'd63095, 16'd32972, 16'd8770, 16'd7876, 16'd22463, 16'd56287, 16'd23785, 16'd57431, 16'd29448, 16'd42031});
	test_expansion(128'h3a9e75b32c2e7d07beb2851eb652338b, {16'd54277, 16'd39546, 16'd21968, 16'd12173, 16'd7025, 16'd7900, 16'd23644, 16'd26544, 16'd50421, 16'd5457, 16'd18964, 16'd45926, 16'd23958, 16'd22097, 16'd6408, 16'd61801, 16'd42156, 16'd3179, 16'd63376, 16'd3615, 16'd18104, 16'd36984, 16'd45520, 16'd12182, 16'd48390, 16'd15171});
	test_expansion(128'h2c18c635d2f29e2a1ef5a490f1fa9117, {16'd60362, 16'd49013, 16'd62908, 16'd11354, 16'd58530, 16'd2712, 16'd33224, 16'd35166, 16'd63548, 16'd46789, 16'd51010, 16'd40839, 16'd10818, 16'd23064, 16'd4960, 16'd25725, 16'd60965, 16'd25894, 16'd12963, 16'd12005, 16'd17145, 16'd61713, 16'd10534, 16'd32213, 16'd8442, 16'd52823});
	test_expansion(128'h3ffe3f5b8efea5a7f644a083f2acbf58, {16'd52275, 16'd42404, 16'd9698, 16'd11646, 16'd31635, 16'd47350, 16'd44091, 16'd57270, 16'd27744, 16'd23879, 16'd48330, 16'd41199, 16'd17935, 16'd10655, 16'd40422, 16'd24331, 16'd41216, 16'd57730, 16'd40632, 16'd16144, 16'd11543, 16'd32359, 16'd33772, 16'd19774, 16'd16434, 16'd23105});
	test_expansion(128'ha15b9bfa61b8ddeee6c7965280a42529, {16'd52824, 16'd32182, 16'd27626, 16'd42953, 16'd46255, 16'd39542, 16'd5237, 16'd37101, 16'd36265, 16'd21258, 16'd28638, 16'd42836, 16'd19396, 16'd63591, 16'd58375, 16'd2229, 16'd35770, 16'd1727, 16'd1881, 16'd65062, 16'd49179, 16'd42138, 16'd32844, 16'd46094, 16'd9600, 16'd58583});
	test_expansion(128'h4d38d8fea75aa22912499d535d39313d, {16'd18357, 16'd60204, 16'd36352, 16'd55899, 16'd54172, 16'd42558, 16'd47609, 16'd63275, 16'd45858, 16'd9544, 16'd42586, 16'd55173, 16'd63281, 16'd23735, 16'd32076, 16'd27268, 16'd40565, 16'd1333, 16'd4185, 16'd49020, 16'd25082, 16'd32098, 16'd54755, 16'd25140, 16'd27549, 16'd64952});
	test_expansion(128'h7561f59de8d2b758cf21eb79f2ffa7b9, {16'd9969, 16'd36485, 16'd46405, 16'd61822, 16'd2177, 16'd33163, 16'd41962, 16'd19065, 16'd36730, 16'd1518, 16'd37435, 16'd62017, 16'd21386, 16'd27090, 16'd16129, 16'd52823, 16'd25708, 16'd40152, 16'd40431, 16'd42756, 16'd37898, 16'd63309, 16'd15323, 16'd29448, 16'd26037, 16'd7182});
	test_expansion(128'h169b5af2af43ba91860bc2f8afc6beb3, {16'd52302, 16'd28796, 16'd49994, 16'd59689, 16'd22309, 16'd14019, 16'd60943, 16'd56066, 16'd26491, 16'd46756, 16'd25976, 16'd19671, 16'd61850, 16'd34746, 16'd31121, 16'd61107, 16'd25548, 16'd26238, 16'd64583, 16'd48260, 16'd60422, 16'd10068, 16'd63083, 16'd33765, 16'd53451, 16'd26584});
	test_expansion(128'ha9e7603d6644973b36ee09bfc5c4db17, {16'd55439, 16'd14461, 16'd15579, 16'd59602, 16'd20107, 16'd59621, 16'd5496, 16'd24347, 16'd2812, 16'd37246, 16'd7175, 16'd58137, 16'd64721, 16'd33457, 16'd15146, 16'd9619, 16'd42111, 16'd55622, 16'd16007, 16'd9529, 16'd10214, 16'd18523, 16'd25479, 16'd53908, 16'd23790, 16'd6959});
	test_expansion(128'h2eb808c4ee144650d91d50aa841a3723, {16'd17556, 16'd11388, 16'd5111, 16'd22297, 16'd17275, 16'd39626, 16'd20428, 16'd39902, 16'd39007, 16'd4458, 16'd21499, 16'd8041, 16'd51175, 16'd49455, 16'd37473, 16'd17145, 16'd30463, 16'd45870, 16'd36576, 16'd2216, 16'd22349, 16'd28957, 16'd46918, 16'd54869, 16'd41857, 16'd55168});
	test_expansion(128'h7f28bac79519a60ca714376ef515d226, {16'd39299, 16'd31619, 16'd49890, 16'd35355, 16'd28302, 16'd26359, 16'd16951, 16'd64298, 16'd44812, 16'd24134, 16'd19546, 16'd5198, 16'd50053, 16'd48080, 16'd55430, 16'd16030, 16'd59140, 16'd9171, 16'd23528, 16'd44876, 16'd2238, 16'd34131, 16'd22889, 16'd29258, 16'd23634, 16'd50559});
	test_expansion(128'h9219d91fa3a77e7fc9b52f1b1f882805, {16'd18514, 16'd59285, 16'd41797, 16'd45571, 16'd7690, 16'd43335, 16'd39662, 16'd13747, 16'd36519, 16'd51133, 16'd60689, 16'd6839, 16'd25831, 16'd48082, 16'd12284, 16'd41168, 16'd64134, 16'd45421, 16'd43233, 16'd19535, 16'd2645, 16'd54535, 16'd50063, 16'd43127, 16'd24182, 16'd63452});
	test_expansion(128'he9042a01f5a8131882fe610c17ca01e6, {16'd25258, 16'd58884, 16'd57413, 16'd3476, 16'd17771, 16'd53715, 16'd16877, 16'd19735, 16'd57621, 16'd28015, 16'd37783, 16'd25808, 16'd57399, 16'd14459, 16'd52667, 16'd65407, 16'd64698, 16'd61622, 16'd8452, 16'd31645, 16'd19411, 16'd19328, 16'd32637, 16'd37476, 16'd56836, 16'd29218});
	test_expansion(128'h74a59fc63e15b7018ebb54dfe9077782, {16'd38140, 16'd33678, 16'd40325, 16'd15357, 16'd26735, 16'd31552, 16'd64390, 16'd24778, 16'd52235, 16'd24340, 16'd59412, 16'd8821, 16'd42169, 16'd15037, 16'd29025, 16'd10929, 16'd63642, 16'd23720, 16'd31304, 16'd61061, 16'd36949, 16'd36257, 16'd44648, 16'd12909, 16'd46047, 16'd12027});
	test_expansion(128'ha0638c02849596acd51ce811059ccf24, {16'd52755, 16'd57408, 16'd50664, 16'd46866, 16'd48779, 16'd13836, 16'd44784, 16'd56588, 16'd57482, 16'd13737, 16'd25866, 16'd35138, 16'd13983, 16'd48368, 16'd34599, 16'd31226, 16'd388, 16'd51722, 16'd40365, 16'd32398, 16'd49498, 16'd13495, 16'd47105, 16'd33340, 16'd34195, 16'd64931});
	test_expansion(128'h4a885f81aaeec2eda3202e1c590a21ee, {16'd60019, 16'd7981, 16'd65000, 16'd46477, 16'd33459, 16'd31224, 16'd3669, 16'd39691, 16'd15154, 16'd64437, 16'd48826, 16'd28351, 16'd65200, 16'd9931, 16'd45956, 16'd42883, 16'd62538, 16'd32020, 16'd9265, 16'd28918, 16'd54449, 16'd44323, 16'd23968, 16'd8538, 16'd31909, 16'd14241});
	test_expansion(128'hb0b9cfcd76468a32f668c9f7a5fa3a6e, {16'd49641, 16'd26631, 16'd23178, 16'd61954, 16'd49083, 16'd50976, 16'd55157, 16'd57429, 16'd15729, 16'd18001, 16'd43326, 16'd29142, 16'd7296, 16'd59282, 16'd56970, 16'd7860, 16'd41995, 16'd25007, 16'd40774, 16'd6195, 16'd14291, 16'd9872, 16'd56576, 16'd22242, 16'd24299, 16'd61084});
	test_expansion(128'hc0ebc5a93e9591710126e133b0825085, {16'd18456, 16'd38978, 16'd25993, 16'd36404, 16'd27756, 16'd24249, 16'd40591, 16'd36428, 16'd51065, 16'd14121, 16'd36847, 16'd51169, 16'd33889, 16'd245, 16'd65455, 16'd31211, 16'd789, 16'd20336, 16'd21745, 16'd55162, 16'd63850, 16'd25241, 16'd50004, 16'd12698, 16'd64015, 16'd15290});
	test_expansion(128'hb1889701a9d145181f8a16dddac981fa, {16'd19341, 16'd19046, 16'd27954, 16'd25027, 16'd11555, 16'd38355, 16'd48654, 16'd55395, 16'd5277, 16'd26817, 16'd35929, 16'd59406, 16'd64378, 16'd52591, 16'd35625, 16'd61861, 16'd22019, 16'd15482, 16'd9148, 16'd38501, 16'd35299, 16'd62389, 16'd60626, 16'd24153, 16'd61208, 16'd16571});
	test_expansion(128'h1673e626c949c3617612c91fe5480129, {16'd16733, 16'd1745, 16'd27318, 16'd45801, 16'd7450, 16'd36742, 16'd18535, 16'd17314, 16'd20962, 16'd15901, 16'd33355, 16'd55439, 16'd17823, 16'd53352, 16'd27191, 16'd52796, 16'd23371, 16'd60741, 16'd46169, 16'd46793, 16'd64560, 16'd42350, 16'd1809, 16'd58505, 16'd16884, 16'd9683});
	test_expansion(128'h76d1d7509574bab9771d768870226407, {16'd4424, 16'd29594, 16'd12031, 16'd61227, 16'd5280, 16'd53242, 16'd20938, 16'd49495, 16'd10137, 16'd20250, 16'd39588, 16'd29753, 16'd7728, 16'd21022, 16'd47481, 16'd46597, 16'd32136, 16'd4837, 16'd3021, 16'd16009, 16'd12433, 16'd29319, 16'd39458, 16'd24728, 16'd24741, 16'd38417});
	test_expansion(128'h1748e899f8e096f41912c18cf4ca6e16, {16'd47228, 16'd59792, 16'd55648, 16'd48010, 16'd48082, 16'd3265, 16'd11706, 16'd18434, 16'd14243, 16'd7538, 16'd50332, 16'd225, 16'd19987, 16'd52770, 16'd54138, 16'd1054, 16'd61261, 16'd28208, 16'd9397, 16'd29748, 16'd65383, 16'd32371, 16'd14153, 16'd1363, 16'd63957, 16'd46216});
	test_expansion(128'hbe11d020c09b6871208b60103cb06be7, {16'd30127, 16'd13337, 16'd61642, 16'd23080, 16'd65383, 16'd61252, 16'd8038, 16'd59396, 16'd22368, 16'd36363, 16'd19757, 16'd23677, 16'd63338, 16'd49950, 16'd28385, 16'd51793, 16'd59871, 16'd11176, 16'd42845, 16'd42582, 16'd34521, 16'd40396, 16'd58290, 16'd58021, 16'd19274, 16'd48923});
	test_expansion(128'hc13445ce92929866acb36549d0d14b1c, {16'd6176, 16'd43454, 16'd15139, 16'd956, 16'd62166, 16'd53509, 16'd41794, 16'd11680, 16'd52716, 16'd19674, 16'd47195, 16'd50050, 16'd9147, 16'd20515, 16'd64863, 16'd55759, 16'd42312, 16'd26957, 16'd11104, 16'd46037, 16'd48057, 16'd45882, 16'd50117, 16'd49413, 16'd31501, 16'd52836});
	test_expansion(128'h8b18910375fab27240ce7a319701fbb8, {16'd50402, 16'd1830, 16'd40330, 16'd15408, 16'd57206, 16'd45903, 16'd41193, 16'd24748, 16'd49962, 16'd46739, 16'd32064, 16'd34704, 16'd20133, 16'd7006, 16'd48879, 16'd13669, 16'd20824, 16'd7458, 16'd5130, 16'd29392, 16'd15340, 16'd34733, 16'd21099, 16'd16623, 16'd28403, 16'd57769});
	test_expansion(128'h8dbfbdcb980e4daf65daf251e38b63c5, {16'd46775, 16'd6148, 16'd62975, 16'd42588, 16'd63844, 16'd56768, 16'd268, 16'd56091, 16'd62675, 16'd62476, 16'd20226, 16'd4977, 16'd21511, 16'd9549, 16'd53710, 16'd59946, 16'd29940, 16'd34150, 16'd59549, 16'd23685, 16'd558, 16'd8949, 16'd54768, 16'd27628, 16'd31524, 16'd61740});
	test_expansion(128'h05dedde0b18dc213ea6b8383570a21d9, {16'd26585, 16'd39414, 16'd44383, 16'd30339, 16'd11337, 16'd10216, 16'd39802, 16'd9836, 16'd14362, 16'd31907, 16'd16114, 16'd31615, 16'd1642, 16'd34158, 16'd31646, 16'd4085, 16'd24404, 16'd25041, 16'd4259, 16'd3108, 16'd27746, 16'd28206, 16'd18669, 16'd23705, 16'd35916, 16'd33242});
	test_expansion(128'h7e482e62d03f0b24dde98ec144d53832, {16'd24885, 16'd274, 16'd4690, 16'd15315, 16'd52147, 16'd24048, 16'd44073, 16'd59474, 16'd54603, 16'd49536, 16'd45800, 16'd42811, 16'd49794, 16'd8194, 16'd58513, 16'd40519, 16'd35671, 16'd56889, 16'd19361, 16'd4077, 16'd18503, 16'd62260, 16'd54400, 16'd43190, 16'd38336, 16'd2386});
	test_expansion(128'hfd73aff453d61983f6f7d3c81efbf470, {16'd28179, 16'd14120, 16'd19739, 16'd60183, 16'd53395, 16'd35647, 16'd64648, 16'd11215, 16'd55627, 16'd54222, 16'd18864, 16'd15778, 16'd35111, 16'd38860, 16'd41271, 16'd61453, 16'd61461, 16'd42044, 16'd11491, 16'd64011, 16'd14242, 16'd62429, 16'd64500, 16'd19824, 16'd17765, 16'd14322});
	test_expansion(128'h80f4f534109a0c1fb1f55d2e799fc3b0, {16'd19108, 16'd3118, 16'd21776, 16'd55284, 16'd9087, 16'd57874, 16'd43802, 16'd18793, 16'd24202, 16'd60202, 16'd6606, 16'd30009, 16'd64793, 16'd36698, 16'd13542, 16'd21601, 16'd28190, 16'd16709, 16'd21623, 16'd23128, 16'd34649, 16'd32553, 16'd21488, 16'd21281, 16'd3618, 16'd13742});
	test_expansion(128'hfd75f9ce06073d2c67c26207fd97298f, {16'd9667, 16'd13882, 16'd40384, 16'd54502, 16'd47210, 16'd32443, 16'd46913, 16'd25826, 16'd62407, 16'd7559, 16'd33462, 16'd44309, 16'd41216, 16'd51737, 16'd31249, 16'd52775, 16'd25237, 16'd55992, 16'd56142, 16'd61162, 16'd29965, 16'd24631, 16'd28896, 16'd54901, 16'd46688, 16'd11873});
	test_expansion(128'h9e80847e06c88c3a5fbd1be093c2fea8, {16'd55036, 16'd57259, 16'd7599, 16'd43521, 16'd40907, 16'd4599, 16'd40926, 16'd28366, 16'd55009, 16'd53892, 16'd22890, 16'd55466, 16'd31885, 16'd2154, 16'd60587, 16'd1203, 16'd3967, 16'd52106, 16'd57402, 16'd15032, 16'd63560, 16'd40822, 16'd50977, 16'd58549, 16'd3471, 16'd9001});
	test_expansion(128'h4423a034ac9abc30442b2baf07fb7856, {16'd30664, 16'd3913, 16'd21464, 16'd56822, 16'd49503, 16'd63532, 16'd60777, 16'd6613, 16'd59153, 16'd41252, 16'd37919, 16'd6671, 16'd27015, 16'd14714, 16'd54356, 16'd6575, 16'd57152, 16'd54708, 16'd64102, 16'd27197, 16'd17093, 16'd429, 16'd19647, 16'd7454, 16'd14006, 16'd18504});
	test_expansion(128'hbaf64ccb1a1b98348d8f417e9481c377, {16'd5103, 16'd1591, 16'd9959, 16'd34887, 16'd46575, 16'd44613, 16'd54854, 16'd44933, 16'd17709, 16'd30770, 16'd37311, 16'd1747, 16'd17480, 16'd3352, 16'd2902, 16'd52859, 16'd23751, 16'd56649, 16'd23269, 16'd48996, 16'd38601, 16'd26891, 16'd7663, 16'd27643, 16'd21962, 16'd33623});
	test_expansion(128'hbfc6a774c608504147043800959dd459, {16'd26732, 16'd49167, 16'd7809, 16'd7538, 16'd35741, 16'd10298, 16'd44070, 16'd16183, 16'd60492, 16'd30854, 16'd49349, 16'd58573, 16'd55955, 16'd34071, 16'd28897, 16'd47283, 16'd62254, 16'd30455, 16'd62850, 16'd54033, 16'd27026, 16'd54273, 16'd54918, 16'd43493, 16'd3607, 16'd40700});
	test_expansion(128'h732dadc5e8ab35884915a8dc089f0512, {16'd37064, 16'd10660, 16'd35535, 16'd29335, 16'd15602, 16'd40305, 16'd45851, 16'd48677, 16'd15661, 16'd27481, 16'd5791, 16'd64353, 16'd1590, 16'd60118, 16'd55089, 16'd16907, 16'd114, 16'd16429, 16'd6392, 16'd48098, 16'd28626, 16'd57965, 16'd10843, 16'd61094, 16'd19624, 16'd23150});
	test_expansion(128'h2ea1a9f90887d0f74002c82115a99db5, {16'd32353, 16'd1781, 16'd28313, 16'd5412, 16'd48245, 16'd30802, 16'd40069, 16'd26605, 16'd49914, 16'd9536, 16'd31433, 16'd31061, 16'd23227, 16'd27621, 16'd49929, 16'd53547, 16'd50093, 16'd15251, 16'd25524, 16'd63659, 16'd1866, 16'd44280, 16'd54196, 16'd3422, 16'd22368, 16'd23148});
	test_expansion(128'ha571b690686754de515f91d922abeb9b, {16'd920, 16'd7297, 16'd45744, 16'd54274, 16'd44209, 16'd11200, 16'd33790, 16'd16308, 16'd11377, 16'd48900, 16'd64301, 16'd44779, 16'd6487, 16'd8635, 16'd6958, 16'd44558, 16'd46885, 16'd37721, 16'd20949, 16'd52265, 16'd10987, 16'd55754, 16'd45187, 16'd13525, 16'd49400, 16'd35663});
	test_expansion(128'h577cf32db8efda51793e60e016a54a2f, {16'd27566, 16'd46241, 16'd25515, 16'd2129, 16'd38124, 16'd42707, 16'd1399, 16'd33480, 16'd7495, 16'd33500, 16'd23022, 16'd13747, 16'd47925, 16'd60363, 16'd48558, 16'd1772, 16'd16091, 16'd39103, 16'd52425, 16'd55041, 16'd53753, 16'd18084, 16'd42584, 16'd22154, 16'd21258, 16'd40684});
	test_expansion(128'hebe8df6f1de7124559adfd87342b7acf, {16'd23040, 16'd27043, 16'd46245, 16'd27722, 16'd40682, 16'd39341, 16'd15768, 16'd32874, 16'd20367, 16'd52666, 16'd28074, 16'd6153, 16'd46678, 16'd58832, 16'd34699, 16'd58307, 16'd62489, 16'd1110, 16'd7511, 16'd10112, 16'd3192, 16'd739, 16'd55247, 16'd63663, 16'd48407, 16'd22139});
	test_expansion(128'hc52a3ece695b34413338a5d9107cf15a, {16'd41633, 16'd10354, 16'd42005, 16'd64487, 16'd36289, 16'd31694, 16'd62068, 16'd21493, 16'd8193, 16'd32660, 16'd52242, 16'd22416, 16'd49753, 16'd30820, 16'd19618, 16'd50470, 16'd49411, 16'd5554, 16'd42970, 16'd50239, 16'd60988, 16'd29095, 16'd24190, 16'd63077, 16'd8006, 16'd9290});
	test_expansion(128'h9f34f9a0cf3e545751b01fee71871f01, {16'd22118, 16'd63492, 16'd38410, 16'd30112, 16'd11828, 16'd58559, 16'd19157, 16'd9032, 16'd22742, 16'd37323, 16'd37945, 16'd40149, 16'd28305, 16'd32296, 16'd7016, 16'd26315, 16'd50799, 16'd39394, 16'd40327, 16'd42311, 16'd38020, 16'd50438, 16'd20673, 16'd21749, 16'd37567, 16'd56216});
	test_expansion(128'ha75d3cf3fe88fd32d64c88f679aff08e, {16'd58125, 16'd4037, 16'd32797, 16'd9872, 16'd15209, 16'd40382, 16'd27841, 16'd56216, 16'd25050, 16'd51573, 16'd24444, 16'd57887, 16'd6491, 16'd48823, 16'd52800, 16'd8272, 16'd44298, 16'd31757, 16'd9464, 16'd3786, 16'd60313, 16'd7542, 16'd3915, 16'd50225, 16'd49039, 16'd16296});
	test_expansion(128'hcfd279d02cae262399b770b2efe56d15, {16'd17475, 16'd16873, 16'd9137, 16'd56061, 16'd55880, 16'd43382, 16'd39310, 16'd52211, 16'd16373, 16'd43493, 16'd11208, 16'd41739, 16'd64900, 16'd63772, 16'd59211, 16'd45678, 16'd26686, 16'd31985, 16'd65037, 16'd51348, 16'd37259, 16'd57871, 16'd9024, 16'd18790, 16'd12695, 16'd37818});
	test_expansion(128'h50b95353ee9afcf481356958216e7a2b, {16'd44320, 16'd12121, 16'd2359, 16'd61426, 16'd46845, 16'd47668, 16'd63856, 16'd25674, 16'd39946, 16'd50381, 16'd31665, 16'd27846, 16'd15956, 16'd42953, 16'd1274, 16'd59078, 16'd57327, 16'd51140, 16'd32763, 16'd58961, 16'd11986, 16'd55014, 16'd33915, 16'd24324, 16'd30765, 16'd11511});
	test_expansion(128'hd03b18e31e821dd90d315fc1f79c385d, {16'd19932, 16'd31602, 16'd15689, 16'd2993, 16'd51906, 16'd23059, 16'd20035, 16'd65528, 16'd46914, 16'd9121, 16'd55388, 16'd58487, 16'd63847, 16'd55681, 16'd43032, 16'd7105, 16'd7962, 16'd24772, 16'd54429, 16'd3111, 16'd5173, 16'd210, 16'd38534, 16'd42827, 16'd30931, 16'd61873});
	test_expansion(128'h280828f77e48b8f4f470f2192713b521, {16'd22619, 16'd937, 16'd2545, 16'd16284, 16'd33820, 16'd55994, 16'd33202, 16'd6453, 16'd56824, 16'd34367, 16'd56432, 16'd27149, 16'd39789, 16'd37935, 16'd45571, 16'd1788, 16'd62948, 16'd41249, 16'd11539, 16'd29323, 16'd23429, 16'd51969, 16'd2912, 16'd27206, 16'd9002, 16'd17549});
	test_expansion(128'hccdc0a2f2e0e5b20a7bdbe399f5a975d, {16'd32590, 16'd26589, 16'd57141, 16'd13325, 16'd56285, 16'd17255, 16'd48994, 16'd28074, 16'd4600, 16'd31617, 16'd3174, 16'd58717, 16'd35360, 16'd33835, 16'd25662, 16'd65194, 16'd40697, 16'd38258, 16'd8657, 16'd206, 16'd46323, 16'd1121, 16'd17587, 16'd34040, 16'd4155, 16'd52735});
	test_expansion(128'hb7b7f184364e0afa52f3706d60127c05, {16'd12519, 16'd29980, 16'd36397, 16'd1270, 16'd36452, 16'd21622, 16'd13031, 16'd500, 16'd53997, 16'd56867, 16'd22493, 16'd59163, 16'd1119, 16'd36513, 16'd56471, 16'd36286, 16'd2846, 16'd55970, 16'd13678, 16'd33116, 16'd13512, 16'd55906, 16'd50000, 16'd46276, 16'd43821, 16'd52586});
	test_expansion(128'h16c4cd9668980bc218cec65259e37ea1, {16'd30948, 16'd23021, 16'd17654, 16'd27892, 16'd54639, 16'd808, 16'd18258, 16'd6726, 16'd55301, 16'd63113, 16'd30576, 16'd10370, 16'd64421, 16'd22795, 16'd39661, 16'd46067, 16'd59093, 16'd25586, 16'd36668, 16'd25712, 16'd62664, 16'd12111, 16'd48856, 16'd23046, 16'd54083, 16'd41448});
	test_expansion(128'hce4288ffa4d745a912e4406635bc7bc4, {16'd45220, 16'd56412, 16'd27491, 16'd18107, 16'd6884, 16'd39968, 16'd45821, 16'd63595, 16'd31717, 16'd17941, 16'd10639, 16'd25806, 16'd42405, 16'd32553, 16'd41193, 16'd8224, 16'd64235, 16'd20569, 16'd62121, 16'd40068, 16'd30823, 16'd60652, 16'd10533, 16'd2650, 16'd28668, 16'd23730});
	test_expansion(128'h010fc851cdd8d0ccf4df893fe463fa4b, {16'd8223, 16'd36512, 16'd26237, 16'd39666, 16'd10164, 16'd51575, 16'd39078, 16'd32928, 16'd11880, 16'd17023, 16'd54064, 16'd518, 16'd54555, 16'd19346, 16'd30592, 16'd10985, 16'd34446, 16'd58404, 16'd29385, 16'd3465, 16'd33416, 16'd55476, 16'd54421, 16'd22474, 16'd752, 16'd26499});
	test_expansion(128'h87774a2138974e01b482102a6aa1cc05, {16'd7916, 16'd63674, 16'd23868, 16'd5641, 16'd45462, 16'd17648, 16'd14786, 16'd63363, 16'd7971, 16'd44560, 16'd28924, 16'd30970, 16'd33201, 16'd30788, 16'd44147, 16'd33281, 16'd12308, 16'd15669, 16'd23925, 16'd8997, 16'd403, 16'd63606, 16'd305, 16'd40367, 16'd60040, 16'd15835});
	test_expansion(128'h1edf1d5174c17d89b63d44f0cb441c4f, {16'd59084, 16'd45335, 16'd6458, 16'd7203, 16'd28527, 16'd28038, 16'd56282, 16'd533, 16'd19463, 16'd53997, 16'd14679, 16'd22630, 16'd63125, 16'd31182, 16'd9446, 16'd31989, 16'd42332, 16'd8754, 16'd52471, 16'd10557, 16'd38413, 16'd23347, 16'd60349, 16'd45272, 16'd41308, 16'd24423});
	test_expansion(128'h84599c8b3deee336d0d721f9b04e754a, {16'd5634, 16'd23622, 16'd56373, 16'd59947, 16'd49452, 16'd514, 16'd52017, 16'd24670, 16'd65165, 16'd51933, 16'd60174, 16'd14508, 16'd30310, 16'd14215, 16'd34877, 16'd5356, 16'd38313, 16'd36137, 16'd32819, 16'd13468, 16'd50625, 16'd1118, 16'd10059, 16'd52094, 16'd41617, 16'd53647});
	test_expansion(128'h2eb884adfa3463c187edb172027f1d0b, {16'd28442, 16'd13237, 16'd42912, 16'd62214, 16'd21456, 16'd799, 16'd221, 16'd6420, 16'd43179, 16'd55317, 16'd29232, 16'd38045, 16'd8886, 16'd52091, 16'd62306, 16'd64721, 16'd12974, 16'd30106, 16'd61142, 16'd27297, 16'd18468, 16'd47435, 16'd16421, 16'd26213, 16'd59230, 16'd15704});
	test_expansion(128'h4c5802de02cd5d6fcd3a15b846eba1f5, {16'd18670, 16'd30553, 16'd45149, 16'd56, 16'd38037, 16'd10030, 16'd64661, 16'd61125, 16'd27207, 16'd54421, 16'd23238, 16'd10992, 16'd48289, 16'd65129, 16'd37513, 16'd51847, 16'd34816, 16'd21215, 16'd26660, 16'd38240, 16'd33756, 16'd28259, 16'd37103, 16'd30380, 16'd38837, 16'd8793});
	test_expansion(128'he4f71c9bfe762bb9e19fee9c5fb0c436, {16'd44112, 16'd6848, 16'd26561, 16'd16040, 16'd35367, 16'd22924, 16'd59470, 16'd33867, 16'd51627, 16'd33189, 16'd47966, 16'd60818, 16'd4140, 16'd12652, 16'd20863, 16'd37914, 16'd34965, 16'd29042, 16'd54087, 16'd6177, 16'd56251, 16'd13924, 16'd35904, 16'd20232, 16'd13573, 16'd39599});
	test_expansion(128'hdc633bfd29bcfa6fca8060abdfd017ea, {16'd59690, 16'd13240, 16'd550, 16'd44624, 16'd37481, 16'd42077, 16'd39967, 16'd31630, 16'd25343, 16'd44810, 16'd704, 16'd48041, 16'd30150, 16'd12326, 16'd21680, 16'd21887, 16'd1806, 16'd62743, 16'd41537, 16'd46616, 16'd23815, 16'd26715, 16'd1930, 16'd61920, 16'd20137, 16'd7931});
	test_expansion(128'h606da19fa25932ea8c7a574447719b5b, {16'd44323, 16'd14086, 16'd3911, 16'd7500, 16'd47758, 16'd25485, 16'd17621, 16'd18785, 16'd52076, 16'd7764, 16'd33413, 16'd60255, 16'd24713, 16'd59061, 16'd58504, 16'd34651, 16'd46747, 16'd27335, 16'd11756, 16'd29216, 16'd8040, 16'd46511, 16'd53614, 16'd28833, 16'd65151, 16'd33451});
	test_expansion(128'h9a3e4c58f765e3898392bf376a94094d, {16'd9412, 16'd58372, 16'd57816, 16'd61891, 16'd7117, 16'd41784, 16'd1441, 16'd13590, 16'd24984, 16'd64828, 16'd46928, 16'd12245, 16'd5284, 16'd43056, 16'd34857, 16'd35037, 16'd8204, 16'd39177, 16'd63139, 16'd29728, 16'd31358, 16'd20367, 16'd1297, 16'd30016, 16'd31250, 16'd36442});
	test_expansion(128'h08bbb49046cddd583a6fc9141efcf705, {16'd52766, 16'd55426, 16'd15788, 16'd21671, 16'd48859, 16'd30859, 16'd57795, 16'd50578, 16'd704, 16'd30671, 16'd15920, 16'd46837, 16'd58020, 16'd9984, 16'd5712, 16'd59983, 16'd61514, 16'd25273, 16'd64558, 16'd52448, 16'd23394, 16'd27103, 16'd62445, 16'd44313, 16'd61628, 16'd10616});
	test_expansion(128'h2dc2dee37102a873888ce694daac39e2, {16'd2496, 16'd8203, 16'd51496, 16'd51084, 16'd47717, 16'd55791, 16'd12102, 16'd15618, 16'd63590, 16'd1319, 16'd28077, 16'd22577, 16'd27257, 16'd39445, 16'd31162, 16'd19623, 16'd59922, 16'd36700, 16'd30205, 16'd64853, 16'd29500, 16'd6270, 16'd46304, 16'd16299, 16'd43902, 16'd55697});
	test_expansion(128'h075dd44cf9795cec874c21081b51ad43, {16'd6312, 16'd63814, 16'd55236, 16'd32152, 16'd21970, 16'd41969, 16'd52999, 16'd63355, 16'd40800, 16'd63671, 16'd30352, 16'd4102, 16'd61511, 16'd32401, 16'd14500, 16'd20157, 16'd25375, 16'd49270, 16'd1771, 16'd9241, 16'd9081, 16'd29787, 16'd25430, 16'd29231, 16'd36500, 16'd24860});
	test_expansion(128'h312f512318329e88c5e6c204d73fa8a7, {16'd10906, 16'd15885, 16'd25514, 16'd38532, 16'd4956, 16'd33116, 16'd35978, 16'd60873, 16'd47712, 16'd20013, 16'd51511, 16'd8870, 16'd50674, 16'd42302, 16'd40965, 16'd36183, 16'd29004, 16'd3501, 16'd13466, 16'd18821, 16'd40136, 16'd5456, 16'd56228, 16'd42094, 16'd51176, 16'd2629});
	test_expansion(128'h9affb62844f7c6910aa11dc29d183589, {16'd61304, 16'd7510, 16'd8768, 16'd62623, 16'd27235, 16'd18270, 16'd8839, 16'd65215, 16'd50874, 16'd40404, 16'd28500, 16'd25374, 16'd52237, 16'd24083, 16'd25650, 16'd23435, 16'd56700, 16'd21361, 16'd37817, 16'd59567, 16'd65262, 16'd29550, 16'd40452, 16'd12173, 16'd33352, 16'd50064});
	test_expansion(128'he834efb7055c3ab3bac5a2772c45a30c, {16'd2418, 16'd14691, 16'd28291, 16'd24497, 16'd58192, 16'd15503, 16'd21297, 16'd56906, 16'd36464, 16'd43144, 16'd36296, 16'd53538, 16'd39855, 16'd25515, 16'd28632, 16'd6605, 16'd49604, 16'd44758, 16'd53244, 16'd65224, 16'd19846, 16'd8665, 16'd51598, 16'd14629, 16'd27153, 16'd49554});
	test_expansion(128'h6e153171536794e01e4f38cd311f7e2a, {16'd54400, 16'd63828, 16'd59048, 16'd51432, 16'd13840, 16'd57744, 16'd44483, 16'd8499, 16'd33514, 16'd40075, 16'd17924, 16'd44300, 16'd34481, 16'd1199, 16'd59508, 16'd43012, 16'd43358, 16'd16723, 16'd57402, 16'd5429, 16'd46401, 16'd6458, 16'd7654, 16'd19942, 16'd42431, 16'd27323});
	test_expansion(128'h640a60ac22cb864651e84ca887d8d30d, {16'd41497, 16'd13289, 16'd32084, 16'd46947, 16'd12953, 16'd18818, 16'd7767, 16'd36350, 16'd19348, 16'd51748, 16'd58089, 16'd21309, 16'd55691, 16'd4482, 16'd6582, 16'd58898, 16'd48902, 16'd58831, 16'd49326, 16'd46732, 16'd28158, 16'd33880, 16'd24695, 16'd47278, 16'd29553, 16'd65227});
	test_expansion(128'h58053fb01e5935df85e73baa49f8656f, {16'd2159, 16'd54670, 16'd37773, 16'd36774, 16'd55517, 16'd51620, 16'd60045, 16'd14911, 16'd59252, 16'd10986, 16'd21651, 16'd52264, 16'd57578, 16'd7425, 16'd1933, 16'd55155, 16'd29561, 16'd12866, 16'd22059, 16'd25474, 16'd25613, 16'd22102, 16'd50095, 16'd65105, 16'd48754, 16'd25790});
	test_expansion(128'hb2ca4044de2a9d5eebb9aeac04ee99cb, {16'd11696, 16'd9834, 16'd15969, 16'd1883, 16'd8232, 16'd9376, 16'd274, 16'd36052, 16'd53279, 16'd12807, 16'd8695, 16'd47322, 16'd57286, 16'd7931, 16'd34887, 16'd47583, 16'd1120, 16'd58377, 16'd60774, 16'd7267, 16'd11, 16'd22070, 16'd42659, 16'd42272, 16'd31982, 16'd32723});
	test_expansion(128'h40c3fecaafdfa79a01db064c6a692340, {16'd36638, 16'd15145, 16'd53866, 16'd29907, 16'd49612, 16'd62534, 16'd18356, 16'd50734, 16'd37089, 16'd28844, 16'd64555, 16'd14426, 16'd20856, 16'd22252, 16'd31767, 16'd5313, 16'd10916, 16'd52380, 16'd61107, 16'd64937, 16'd58041, 16'd64250, 16'd49615, 16'd63798, 16'd49335, 16'd3512});
	test_expansion(128'h4116ba1396cce5f7ba0d6414433dad0f, {16'd40426, 16'd17443, 16'd24569, 16'd78, 16'd44954, 16'd64171, 16'd17958, 16'd54762, 16'd22586, 16'd37549, 16'd46488, 16'd51882, 16'd36182, 16'd25866, 16'd49072, 16'd6240, 16'd43041, 16'd59904, 16'd35294, 16'd52104, 16'd20920, 16'd50775, 16'd30623, 16'd62723, 16'd32681, 16'd27913});
	test_expansion(128'hdd9720a6fae2257d4b4cc5ef3ef2d9b6, {16'd24148, 16'd35019, 16'd35593, 16'd53531, 16'd40382, 16'd43511, 16'd22815, 16'd14846, 16'd29601, 16'd18269, 16'd54877, 16'd15550, 16'd45841, 16'd19485, 16'd9894, 16'd38046, 16'd12059, 16'd37854, 16'd35816, 16'd9194, 16'd47137, 16'd34773, 16'd15877, 16'd38781, 16'd12348, 16'd42810});
	test_expansion(128'h4ae2c79a767766edc047d36c8af2ae10, {16'd50019, 16'd62187, 16'd5372, 16'd59822, 16'd3617, 16'd34364, 16'd22141, 16'd60064, 16'd14527, 16'd14251, 16'd6275, 16'd38477, 16'd2287, 16'd20317, 16'd21074, 16'd24485, 16'd27987, 16'd63033, 16'd17367, 16'd47225, 16'd61363, 16'd60532, 16'd25579, 16'd45905, 16'd17773, 16'd35145});
	test_expansion(128'h7c0064df891f1a52f8d0adaf4b1ef89a, {16'd61021, 16'd50888, 16'd43469, 16'd37203, 16'd26482, 16'd63835, 16'd4164, 16'd40895, 16'd37878, 16'd31363, 16'd25792, 16'd38817, 16'd23553, 16'd27092, 16'd2628, 16'd37813, 16'd13049, 16'd3163, 16'd511, 16'd15737, 16'd17862, 16'd61600, 16'd34978, 16'd36062, 16'd34503, 16'd57516});
	test_expansion(128'h9be1293d6b4447c927a5741d6f73012e, {16'd34971, 16'd33629, 16'd43106, 16'd34022, 16'd14723, 16'd20145, 16'd57453, 16'd2304, 16'd13822, 16'd23052, 16'd30927, 16'd47088, 16'd43609, 16'd38220, 16'd20616, 16'd61005, 16'd18334, 16'd48002, 16'd43846, 16'd38851, 16'd32806, 16'd50407, 16'd26447, 16'd26956, 16'd62539, 16'd12508});
	test_expansion(128'hf0016323ccb7ad4e2bbce33ed1f2caf0, {16'd58882, 16'd8283, 16'd42430, 16'd46418, 16'd22730, 16'd5521, 16'd33877, 16'd10850, 16'd11760, 16'd31953, 16'd65010, 16'd10382, 16'd50792, 16'd51238, 16'd58328, 16'd30122, 16'd59898, 16'd61386, 16'd11294, 16'd9335, 16'd41155, 16'd13714, 16'd57402, 16'd3948, 16'd25652, 16'd36193});
	test_expansion(128'h0dd0f1810fa7aec3c101a7af07b20aaf, {16'd58310, 16'd17639, 16'd20340, 16'd52289, 16'd37100, 16'd12249, 16'd30157, 16'd26523, 16'd501, 16'd63698, 16'd60433, 16'd58825, 16'd35850, 16'd35237, 16'd33929, 16'd54285, 16'd56886, 16'd2830, 16'd7953, 16'd63599, 16'd56576, 16'd50534, 16'd63450, 16'd9784, 16'd61956, 16'd1426});
	test_expansion(128'hdb1cc6c77772124599f56e49713e6691, {16'd41463, 16'd18445, 16'd55279, 16'd5086, 16'd20982, 16'd34413, 16'd47396, 16'd30357, 16'd43178, 16'd36423, 16'd7059, 16'd11332, 16'd36486, 16'd8725, 16'd20191, 16'd48006, 16'd7260, 16'd57138, 16'd59455, 16'd35040, 16'd63209, 16'd61136, 16'd11246, 16'd28949, 16'd19054, 16'd47573});
	test_expansion(128'hca15c6cecc61ad28df9de28d3008beb8, {16'd48856, 16'd57951, 16'd64650, 16'd619, 16'd62853, 16'd37347, 16'd45646, 16'd45080, 16'd24739, 16'd45928, 16'd61529, 16'd9677, 16'd64697, 16'd38627, 16'd51796, 16'd60158, 16'd29042, 16'd4572, 16'd21139, 16'd32161, 16'd57512, 16'd23910, 16'd64060, 16'd8370, 16'd35637, 16'd45914});
	test_expansion(128'h8bbebba534e6193d33e4b133a0362e63, {16'd1136, 16'd30786, 16'd35209, 16'd47083, 16'd56752, 16'd22299, 16'd33549, 16'd23437, 16'd44205, 16'd32438, 16'd36289, 16'd65334, 16'd17944, 16'd22988, 16'd49233, 16'd1378, 16'd42985, 16'd48672, 16'd60994, 16'd57401, 16'd12458, 16'd9241, 16'd45164, 16'd14806, 16'd45118, 16'd55181});
	test_expansion(128'h03f5d893210f6e0d3959958064ff208f, {16'd50718, 16'd46402, 16'd51064, 16'd43022, 16'd8751, 16'd28839, 16'd44958, 16'd33274, 16'd11072, 16'd1981, 16'd45981, 16'd61266, 16'd61850, 16'd58376, 16'd62356, 16'd49398, 16'd19455, 16'd21325, 16'd4770, 16'd13148, 16'd23079, 16'd24110, 16'd62140, 16'd14435, 16'd64521, 16'd37182});
	test_expansion(128'ha0f4c609ce2bc856d6b31d01460564c9, {16'd31177, 16'd45562, 16'd54268, 16'd3032, 16'd10583, 16'd10937, 16'd48872, 16'd34027, 16'd40757, 16'd63956, 16'd60600, 16'd218, 16'd25836, 16'd42453, 16'd4979, 16'd61139, 16'd29268, 16'd39200, 16'd26515, 16'd64953, 16'd59891, 16'd11414, 16'd65528, 16'd45468, 16'd62443, 16'd18567});
	test_expansion(128'h3beb6cdf8dd3d14210115dfe8bb5f430, {16'd46118, 16'd39188, 16'd23506, 16'd52934, 16'd2320, 16'd37804, 16'd63488, 16'd19588, 16'd62841, 16'd49771, 16'd14650, 16'd7577, 16'd1409, 16'd61177, 16'd14890, 16'd6054, 16'd55508, 16'd40775, 16'd45152, 16'd60031, 16'd56890, 16'd56187, 16'd49387, 16'd48026, 16'd58599, 16'd16639});
	test_expansion(128'h1b5196efab5e7fe3e1417d6ebb3f8d33, {16'd52022, 16'd43985, 16'd1882, 16'd57553, 16'd47864, 16'd32484, 16'd30935, 16'd40531, 16'd49344, 16'd43586, 16'd45060, 16'd6143, 16'd23687, 16'd24239, 16'd52766, 16'd47674, 16'd14587, 16'd52076, 16'd12245, 16'd15942, 16'd4716, 16'd13534, 16'd5226, 16'd12269, 16'd10150, 16'd26243});
	test_expansion(128'h58740dbe7b1068050c28050dac9e2772, {16'd32841, 16'd50329, 16'd6071, 16'd64276, 16'd55007, 16'd61595, 16'd48390, 16'd25112, 16'd38529, 16'd33744, 16'd4232, 16'd13353, 16'd32909, 16'd48636, 16'd1417, 16'd3871, 16'd9697, 16'd34702, 16'd39084, 16'd41890, 16'd47789, 16'd37347, 16'd54174, 16'd42413, 16'd17096, 16'd9197});
	test_expansion(128'he93a00ec4f7f1a05332264f63ffb38d4, {16'd38068, 16'd55681, 16'd60976, 16'd20620, 16'd45845, 16'd14232, 16'd42842, 16'd49893, 16'd63957, 16'd38342, 16'd57639, 16'd8854, 16'd23306, 16'd39641, 16'd35335, 16'd59955, 16'd49554, 16'd5589, 16'd57816, 16'd68, 16'd54939, 16'd34913, 16'd39387, 16'd54172, 16'd33321, 16'd32714});
	test_expansion(128'h99632b03ac8e10cb1a9359bcd4fd662e, {16'd54400, 16'd37831, 16'd18946, 16'd38720, 16'd10905, 16'd54005, 16'd1826, 16'd11115, 16'd55544, 16'd56862, 16'd13670, 16'd2390, 16'd46372, 16'd324, 16'd48859, 16'd15930, 16'd15855, 16'd10484, 16'd55383, 16'd40096, 16'd27496, 16'd2215, 16'd64683, 16'd39341, 16'd1161, 16'd4089});
	test_expansion(128'h34767e322d27c85093acba1af4cecd6f, {16'd7306, 16'd38997, 16'd58552, 16'd44479, 16'd36274, 16'd559, 16'd10057, 16'd60349, 16'd6443, 16'd65413, 16'd17940, 16'd28268, 16'd42068, 16'd2871, 16'd4702, 16'd14071, 16'd44669, 16'd35628, 16'd5170, 16'd35309, 16'd51488, 16'd21858, 16'd38208, 16'd12582, 16'd7647, 16'd62511});
	test_expansion(128'hf249aa81e684f3fbac654f1e1b62755c, {16'd33129, 16'd64799, 16'd62597, 16'd38625, 16'd3792, 16'd39299, 16'd2008, 16'd42531, 16'd33661, 16'd16997, 16'd48799, 16'd42615, 16'd28098, 16'd38346, 16'd27024, 16'd5209, 16'd14360, 16'd43292, 16'd60588, 16'd55306, 16'd61710, 16'd56515, 16'd25509, 16'd63572, 16'd9672, 16'd49319});
	test_expansion(128'h3d4c7e61e64c02b449ba84fa8268bd3c, {16'd58967, 16'd39908, 16'd63893, 16'd33484, 16'd5462, 16'd51994, 16'd18404, 16'd45845, 16'd64391, 16'd50367, 16'd44379, 16'd42239, 16'd45088, 16'd25478, 16'd25432, 16'd29675, 16'd20076, 16'd9467, 16'd49452, 16'd53225, 16'd57932, 16'd41984, 16'd25610, 16'd13032, 16'd2477, 16'd14349});
	test_expansion(128'h2fa344175611ee0fb9729e8ad09b0464, {16'd53459, 16'd13610, 16'd59556, 16'd2272, 16'd20597, 16'd63442, 16'd18259, 16'd45210, 16'd24879, 16'd40860, 16'd28366, 16'd53005, 16'd61003, 16'd61592, 16'd20429, 16'd5568, 16'd8133, 16'd49766, 16'd4037, 16'd44927, 16'd19464, 16'd26113, 16'd35401, 16'd27928, 16'd50325, 16'd32409});
	test_expansion(128'h31fdcf4c0373535d0c7498c6ad3bfe48, {16'd1929, 16'd23928, 16'd41937, 16'd28059, 16'd44486, 16'd33881, 16'd52637, 16'd45607, 16'd56154, 16'd33035, 16'd11187, 16'd19909, 16'd34639, 16'd33807, 16'd40099, 16'd35830, 16'd4731, 16'd21684, 16'd13293, 16'd7741, 16'd4423, 16'd48577, 16'd25174, 16'd46324, 16'd46416, 16'd15211});
	test_expansion(128'hed2ddb289a0d7ee3074fed90c7f491b9, {16'd25993, 16'd57025, 16'd43265, 16'd58895, 16'd15742, 16'd9517, 16'd43755, 16'd26092, 16'd31271, 16'd63434, 16'd51148, 16'd31011, 16'd64108, 16'd7872, 16'd42420, 16'd8880, 16'd20275, 16'd25922, 16'd41078, 16'd16985, 16'd44982, 16'd16261, 16'd20036, 16'd58131, 16'd43299, 16'd2800});
	test_expansion(128'h7957fb85820894ba53c90e43485675bd, {16'd4667, 16'd46501, 16'd64169, 16'd10288, 16'd3293, 16'd4324, 16'd38512, 16'd55814, 16'd64124, 16'd20505, 16'd21434, 16'd9379, 16'd17158, 16'd59625, 16'd2117, 16'd34676, 16'd44789, 16'd14582, 16'd48770, 16'd1105, 16'd55049, 16'd40828, 16'd59141, 16'd28965, 16'd3196, 16'd43646});
	test_expansion(128'h7c09bea7688451266ba0418a25a6ea09, {16'd18192, 16'd25079, 16'd56405, 16'd40804, 16'd52388, 16'd48315, 16'd63869, 16'd17831, 16'd65487, 16'd53065, 16'd40933, 16'd54577, 16'd63584, 16'd45178, 16'd9477, 16'd14082, 16'd30737, 16'd51950, 16'd49399, 16'd29017, 16'd15813, 16'd6513, 16'd27121, 16'd49506, 16'd12185, 16'd20385});
	test_expansion(128'h3af5871087271c7e8f33a6433b564715, {16'd17344, 16'd24228, 16'd60134, 16'd3512, 16'd61585, 16'd31384, 16'd14755, 16'd42319, 16'd23601, 16'd51215, 16'd22366, 16'd4516, 16'd22812, 16'd34408, 16'd24527, 16'd64673, 16'd51481, 16'd24569, 16'd19261, 16'd54669, 16'd23033, 16'd43108, 16'd58036, 16'd8649, 16'd23573, 16'd25163});
	test_expansion(128'hc22131d66f49f95e438db7b2e9575c92, {16'd33170, 16'd26504, 16'd22941, 16'd32387, 16'd8930, 16'd41261, 16'd3596, 16'd35384, 16'd10080, 16'd9430, 16'd11750, 16'd47474, 16'd51083, 16'd41370, 16'd42018, 16'd5589, 16'd42503, 16'd11116, 16'd59631, 16'd15445, 16'd62646, 16'd53812, 16'd53202, 16'd10572, 16'd19102, 16'd54511});
	test_expansion(128'hc8cdad5da07acc7521887286387ba97c, {16'd48334, 16'd23251, 16'd22850, 16'd674, 16'd22471, 16'd43048, 16'd6170, 16'd45036, 16'd2237, 16'd16504, 16'd12631, 16'd13902, 16'd58432, 16'd5764, 16'd45934, 16'd11926, 16'd40927, 16'd28414, 16'd31061, 16'd10809, 16'd54466, 16'd13284, 16'd8152, 16'd41891, 16'd1651, 16'd14289});
	test_expansion(128'h183d4ce25e6c1cbf5b8b15af49ed822f, {16'd35061, 16'd10961, 16'd27444, 16'd55875, 16'd49028, 16'd7562, 16'd38358, 16'd50412, 16'd49815, 16'd9621, 16'd50839, 16'd9030, 16'd31502, 16'd5907, 16'd29064, 16'd2134, 16'd14150, 16'd26399, 16'd57847, 16'd34724, 16'd45120, 16'd2739, 16'd37858, 16'd51569, 16'd21064, 16'd46063});
	test_expansion(128'h998b367a9b4e7c63b251e4ee4bfcee38, {16'd21457, 16'd41950, 16'd55011, 16'd54935, 16'd59219, 16'd35187, 16'd8182, 16'd38181, 16'd41789, 16'd47572, 16'd19172, 16'd13676, 16'd45126, 16'd53539, 16'd51056, 16'd10355, 16'd39940, 16'd11174, 16'd24801, 16'd24993, 16'd24298, 16'd6210, 16'd45419, 16'd18815, 16'd31115, 16'd16365});
	test_expansion(128'h61b13efe1cfb8c3b407c594d9660469c, {16'd59539, 16'd42404, 16'd29477, 16'd36050, 16'd11752, 16'd3740, 16'd60327, 16'd51816, 16'd41539, 16'd13482, 16'd63280, 16'd35921, 16'd5738, 16'd29865, 16'd37910, 16'd39247, 16'd31395, 16'd54976, 16'd34388, 16'd4468, 16'd50453, 16'd39080, 16'd29852, 16'd23150, 16'd7010, 16'd46774});
	test_expansion(128'h86cb10c12be414d68c9c138964906b0e, {16'd56682, 16'd22219, 16'd32366, 16'd31729, 16'd24046, 16'd62998, 16'd40943, 16'd61308, 16'd37505, 16'd28680, 16'd24034, 16'd29656, 16'd28455, 16'd59464, 16'd45145, 16'd57314, 16'd35370, 16'd49422, 16'd49086, 16'd476, 16'd38400, 16'd16068, 16'd12018, 16'd41628, 16'd58014, 16'd13842});
	test_expansion(128'h2e818cf21fc53f22f3829223721d1dab, {16'd30836, 16'd51479, 16'd44117, 16'd56092, 16'd28200, 16'd11208, 16'd44436, 16'd40102, 16'd61119, 16'd22172, 16'd26670, 16'd54884, 16'd11421, 16'd65449, 16'd22115, 16'd45410, 16'd13335, 16'd49981, 16'd54825, 16'd58134, 16'd15835, 16'd27132, 16'd21807, 16'd38778, 16'd40817, 16'd54279});
	test_expansion(128'hf87f6a7905afbb9733f582522a0a32bd, {16'd56641, 16'd31471, 16'd16443, 16'd30977, 16'd24328, 16'd19706, 16'd1946, 16'd24108, 16'd48141, 16'd12909, 16'd1370, 16'd58356, 16'd23911, 16'd21804, 16'd40484, 16'd17965, 16'd28355, 16'd23419, 16'd20906, 16'd38021, 16'd38828, 16'd5856, 16'd17181, 16'd32962, 16'd3816, 16'd29897});
	test_expansion(128'h6e8674b0ab7e8436d00ac7dc66cd1fa8, {16'd11300, 16'd57089, 16'd17804, 16'd24580, 16'd3631, 16'd34660, 16'd36595, 16'd56965, 16'd40710, 16'd52957, 16'd36176, 16'd44656, 16'd23618, 16'd5688, 16'd60187, 16'd39523, 16'd63559, 16'd37861, 16'd63599, 16'd2044, 16'd65153, 16'd42989, 16'd38004, 16'd21921, 16'd3436, 16'd55027});
	test_expansion(128'hcf8130ad339e205f57e6e727a8974ac9, {16'd61174, 16'd32706, 16'd46242, 16'd11211, 16'd39565, 16'd19292, 16'd26950, 16'd62217, 16'd2896, 16'd36301, 16'd10139, 16'd31434, 16'd12632, 16'd55962, 16'd15504, 16'd47555, 16'd39013, 16'd51434, 16'd53260, 16'd16886, 16'd58361, 16'd28963, 16'd61200, 16'd24722, 16'd13657, 16'd30255});
	test_expansion(128'hfbcd765a12398e7951ef2c30f7af1c7e, {16'd23984, 16'd20894, 16'd55361, 16'd1859, 16'd12390, 16'd26837, 16'd39480, 16'd60819, 16'd46524, 16'd63695, 16'd45424, 16'd25187, 16'd37118, 16'd27102, 16'd12234, 16'd56147, 16'd18544, 16'd16571, 16'd26575, 16'd13200, 16'd32366, 16'd53259, 16'd11122, 16'd58491, 16'd56829, 16'd5081});
	test_expansion(128'h80cf9e2bd47e20988a934308adc5c277, {16'd27680, 16'd28248, 16'd11466, 16'd3396, 16'd62972, 16'd58407, 16'd10844, 16'd25270, 16'd21681, 16'd62966, 16'd34991, 16'd986, 16'd25571, 16'd60406, 16'd64289, 16'd32127, 16'd29090, 16'd61755, 16'd45798, 16'd55705, 16'd62232, 16'd575, 16'd32042, 16'd7973, 16'd61137, 16'd29776});
	test_expansion(128'hfcb8091a3206be1226394037a7100294, {16'd46576, 16'd13727, 16'd59299, 16'd24599, 16'd37858, 16'd1346, 16'd34790, 16'd55115, 16'd48003, 16'd42967, 16'd56434, 16'd22432, 16'd813, 16'd15807, 16'd48456, 16'd14648, 16'd33261, 16'd22584, 16'd30615, 16'd19952, 16'd37130, 16'd63478, 16'd3014, 16'd65163, 16'd2643, 16'd2538});
	test_expansion(128'ha1d51c6ad9d03e2c2e223ddcaccf3a64, {16'd64395, 16'd48819, 16'd3770, 16'd58049, 16'd26167, 16'd31289, 16'd919, 16'd17822, 16'd30185, 16'd7180, 16'd27496, 16'd52089, 16'd11776, 16'd31455, 16'd48950, 16'd49133, 16'd31859, 16'd34841, 16'd31776, 16'd55433, 16'd12329, 16'd20150, 16'd45442, 16'd46431, 16'd57024, 16'd9913});
	test_expansion(128'h09b8fc0979b8736975316203363e300c, {16'd21797, 16'd6504, 16'd64712, 16'd29216, 16'd26103, 16'd7181, 16'd58477, 16'd35631, 16'd26637, 16'd39258, 16'd39798, 16'd28904, 16'd41968, 16'd28135, 16'd54868, 16'd23713, 16'd24679, 16'd8128, 16'd59013, 16'd56243, 16'd7137, 16'd51857, 16'd26811, 16'd25015, 16'd23130, 16'd55766});
	test_expansion(128'hec111aac9798d880540dc409157966ab, {16'd60550, 16'd14885, 16'd15960, 16'd10966, 16'd38307, 16'd62716, 16'd14690, 16'd4135, 16'd3268, 16'd34611, 16'd45353, 16'd40949, 16'd4, 16'd34301, 16'd26902, 16'd65332, 16'd56577, 16'd58635, 16'd32774, 16'd32149, 16'd40424, 16'd43848, 16'd48443, 16'd26939, 16'd24876, 16'd33965});
	test_expansion(128'hd99c55b9bc02af7cb3f78ae1d4f68016, {16'd63718, 16'd64672, 16'd47613, 16'd32624, 16'd18193, 16'd13466, 16'd32259, 16'd10434, 16'd20134, 16'd59041, 16'd49575, 16'd35249, 16'd37107, 16'd58580, 16'd31103, 16'd23974, 16'd42814, 16'd29933, 16'd38778, 16'd53474, 16'd1215, 16'd24420, 16'd269, 16'd8727, 16'd58027, 16'd28573});
	test_expansion(128'hccd5c9adc0681aaabcdfa154d236ed98, {16'd34763, 16'd55826, 16'd11837, 16'd14626, 16'd6293, 16'd37571, 16'd43182, 16'd45768, 16'd5517, 16'd2696, 16'd43909, 16'd38485, 16'd4886, 16'd37814, 16'd58775, 16'd53008, 16'd35440, 16'd61565, 16'd35918, 16'd17224, 16'd60525, 16'd9455, 16'd24843, 16'd49021, 16'd61563, 16'd6777});
	test_expansion(128'hfb9cd392801029bdaca6b0bef20864b0, {16'd44111, 16'd36506, 16'd54260, 16'd65012, 16'd60894, 16'd37812, 16'd45219, 16'd55771, 16'd4659, 16'd14310, 16'd45946, 16'd60297, 16'd3241, 16'd42022, 16'd21399, 16'd18993, 16'd3712, 16'd26588, 16'd52606, 16'd58385, 16'd33421, 16'd38071, 16'd10384, 16'd25721, 16'd34696, 16'd58984});
	test_expansion(128'h6ee5036fbf3c496a7fb3717d0e1d8e02, {16'd1097, 16'd9024, 16'd33976, 16'd60331, 16'd8658, 16'd49219, 16'd42016, 16'd9787, 16'd13502, 16'd58951, 16'd9578, 16'd50337, 16'd233, 16'd46208, 16'd36516, 16'd32183, 16'd63344, 16'd29889, 16'd54888, 16'd60491, 16'd54497, 16'd7804, 16'd52603, 16'd38499, 16'd9524, 16'd31567});
	test_expansion(128'h35ef5136af0b3c82461c29eaf7230542, {16'd64220, 16'd26225, 16'd51932, 16'd10650, 16'd11799, 16'd59605, 16'd54047, 16'd26268, 16'd142, 16'd46572, 16'd29720, 16'd2383, 16'd26705, 16'd40587, 16'd38556, 16'd43845, 16'd36952, 16'd218, 16'd16914, 16'd18517, 16'd45518, 16'd64009, 16'd34465, 16'd65111, 16'd24825, 16'd32872});
	test_expansion(128'hde2480b790010209f83c1a78ba8affb8, {16'd24195, 16'd18063, 16'd10764, 16'd1331, 16'd46601, 16'd27033, 16'd55636, 16'd52475, 16'd10951, 16'd50899, 16'd61864, 16'd8401, 16'd21726, 16'd62648, 16'd36725, 16'd29360, 16'd29359, 16'd8406, 16'd17280, 16'd27571, 16'd36260, 16'd19422, 16'd35553, 16'd55468, 16'd16854, 16'd64892});
	test_expansion(128'h999f2e9ce4df60899aff04a7c5d82592, {16'd53131, 16'd64608, 16'd65249, 16'd10464, 16'd55552, 16'd58137, 16'd31586, 16'd3582, 16'd27398, 16'd8336, 16'd8787, 16'd43399, 16'd3373, 16'd13844, 16'd44339, 16'd16640, 16'd25015, 16'd54966, 16'd745, 16'd23785, 16'd4370, 16'd23805, 16'd10300, 16'd50602, 16'd22564, 16'd39115});
	test_expansion(128'ha7c9f766076dbc6cb60da18d0d2791b1, {16'd958, 16'd10308, 16'd25453, 16'd24503, 16'd53576, 16'd27022, 16'd45980, 16'd42903, 16'd56974, 16'd15868, 16'd49548, 16'd5287, 16'd24860, 16'd61913, 16'd19138, 16'd43796, 16'd40410, 16'd28077, 16'd9240, 16'd32377, 16'd54534, 16'd60216, 16'd4193, 16'd26338, 16'd30856, 16'd2250});
	test_expansion(128'hc68832bb0220174068978feb0848a14a, {16'd17633, 16'd7602, 16'd53229, 16'd47606, 16'd5012, 16'd5550, 16'd22368, 16'd53905, 16'd20386, 16'd40275, 16'd756, 16'd39727, 16'd36138, 16'd61848, 16'd24699, 16'd61047, 16'd53143, 16'd5750, 16'd4615, 16'd65397, 16'd49386, 16'd60263, 16'd18651, 16'd22710, 16'd10725, 16'd29925});
	test_expansion(128'he520d2a7947fc4486b2d481fb5e92458, {16'd57168, 16'd35776, 16'd17921, 16'd57735, 16'd64417, 16'd6883, 16'd11321, 16'd14905, 16'd46536, 16'd54547, 16'd40462, 16'd32106, 16'd63508, 16'd58174, 16'd53616, 16'd55834, 16'd37879, 16'd3645, 16'd58978, 16'd60980, 16'd55611, 16'd51155, 16'd13722, 16'd5185, 16'd36689, 16'd60209});
	test_expansion(128'h3194c1a4f188259d56d6d5e7d4233923, {16'd12969, 16'd60035, 16'd32971, 16'd43832, 16'd36994, 16'd46211, 16'd18472, 16'd896, 16'd37238, 16'd43007, 16'd60152, 16'd52995, 16'd20312, 16'd27888, 16'd29589, 16'd224, 16'd42433, 16'd29395, 16'd5331, 16'd7227, 16'd27523, 16'd27250, 16'd59895, 16'd4469, 16'd1067, 16'd51315});
	test_expansion(128'h9d863b1047b9bd0c7694f653e163d2bd, {16'd33844, 16'd8202, 16'd2611, 16'd4674, 16'd43057, 16'd57357, 16'd49726, 16'd39077, 16'd5551, 16'd54098, 16'd49940, 16'd13370, 16'd45655, 16'd29496, 16'd33123, 16'd22021, 16'd55946, 16'd31864, 16'd25806, 16'd11696, 16'd20467, 16'd61395, 16'd5844, 16'd6953, 16'd18095, 16'd54611});
	test_expansion(128'h5979c6c394f3c6b24b39efe5854d9ec8, {16'd22255, 16'd31204, 16'd2190, 16'd53437, 16'd6063, 16'd56620, 16'd15710, 16'd51567, 16'd20102, 16'd30726, 16'd23730, 16'd55251, 16'd18865, 16'd40381, 16'd18486, 16'd2991, 16'd48449, 16'd478, 16'd41896, 16'd37009, 16'd65161, 16'd42837, 16'd17924, 16'd52921, 16'd31745, 16'd46019});
	test_expansion(128'hbe95bbe2873eee08fef8414d09d2eb86, {16'd43060, 16'd31141, 16'd60947, 16'd38206, 16'd4974, 16'd37674, 16'd36867, 16'd41701, 16'd32750, 16'd43127, 16'd50660, 16'd57766, 16'd36670, 16'd25287, 16'd30707, 16'd24760, 16'd50427, 16'd36713, 16'd62260, 16'd44704, 16'd27508, 16'd38652, 16'd60537, 16'd44733, 16'd56701, 16'd54559});
	test_expansion(128'h88c965a4ce1b9da562f9b599d94e89fd, {16'd53899, 16'd44081, 16'd48995, 16'd13843, 16'd54159, 16'd12308, 16'd44335, 16'd9388, 16'd8719, 16'd14825, 16'd59803, 16'd62048, 16'd56764, 16'd54162, 16'd17837, 16'd18655, 16'd41334, 16'd54820, 16'd18137, 16'd57323, 16'd52552, 16'd10723, 16'd37600, 16'd25379, 16'd38484, 16'd33825});
	test_expansion(128'h145243841720320c852ae2381423b476, {16'd2049, 16'd1701, 16'd15980, 16'd50333, 16'd7105, 16'd64098, 16'd6532, 16'd31547, 16'd51370, 16'd52797, 16'd34835, 16'd2368, 16'd37821, 16'd59373, 16'd51482, 16'd26738, 16'd63004, 16'd15758, 16'd59949, 16'd49684, 16'd44500, 16'd53987, 16'd61531, 16'd61217, 16'd57502, 16'd47196});
	test_expansion(128'h4c876c7f6a44feff7b3f456739edffcb, {16'd3793, 16'd10888, 16'd53707, 16'd10384, 16'd58612, 16'd62755, 16'd56811, 16'd23695, 16'd22944, 16'd47308, 16'd52632, 16'd39727, 16'd29625, 16'd51475, 16'd26264, 16'd16524, 16'd63922, 16'd20610, 16'd33143, 16'd43405, 16'd3888, 16'd35531, 16'd37727, 16'd31506, 16'd14776, 16'd27881});
	test_expansion(128'hbff43fe8f7f80b52b5c1ba44caa852de, {16'd46839, 16'd44257, 16'd19132, 16'd45375, 16'd42150, 16'd13783, 16'd5479, 16'd1729, 16'd32350, 16'd9965, 16'd40421, 16'd31973, 16'd35289, 16'd9574, 16'd64522, 16'd64343, 16'd65447, 16'd19623, 16'd32566, 16'd51504, 16'd47480, 16'd42232, 16'd16163, 16'd58981, 16'd1894, 16'd43121});
	test_expansion(128'h5a8cee8cb45cc55c3dbc034bf9e28c0c, {16'd14411, 16'd13000, 16'd37823, 16'd31513, 16'd49678, 16'd13348, 16'd22440, 16'd34800, 16'd25622, 16'd47607, 16'd25596, 16'd58194, 16'd64098, 16'd65157, 16'd15524, 16'd26569, 16'd22905, 16'd29247, 16'd47970, 16'd23744, 16'd32682, 16'd18774, 16'd55776, 16'd30797, 16'd9702, 16'd47732});
	test_expansion(128'h6abedc296387eeda7a4819c66a6a659e, {16'd57931, 16'd11628, 16'd38998, 16'd17786, 16'd55911, 16'd20391, 16'd59724, 16'd18162, 16'd40994, 16'd36577, 16'd45606, 16'd42716, 16'd58499, 16'd62720, 16'd48332, 16'd59602, 16'd7992, 16'd50385, 16'd54407, 16'd36146, 16'd8865, 16'd13322, 16'd26924, 16'd53856, 16'd65303, 16'd45647});
	test_expansion(128'h0aba83695484a8ba770790a590863f84, {16'd42235, 16'd10006, 16'd55052, 16'd11095, 16'd14542, 16'd24801, 16'd62807, 16'd25617, 16'd34921, 16'd41056, 16'd60802, 16'd11526, 16'd61783, 16'd40837, 16'd48166, 16'd18483, 16'd54229, 16'd36465, 16'd63690, 16'd34563, 16'd34164, 16'd48592, 16'd55253, 16'd63803, 16'd50140, 16'd32107});
	test_expansion(128'h5b855b4eaeb8ea6e7e74ee5c930a268c, {16'd22092, 16'd61155, 16'd45046, 16'd65256, 16'd33428, 16'd55905, 16'd50123, 16'd21363, 16'd23258, 16'd64322, 16'd49061, 16'd41284, 16'd23102, 16'd58219, 16'd35591, 16'd51143, 16'd8490, 16'd38826, 16'd7134, 16'd44541, 16'd29668, 16'd41254, 16'd64384, 16'd65031, 16'd55862, 16'd54114});
	test_expansion(128'h99fee199cd2eb242a96ddbcd65e5581e, {16'd37715, 16'd13268, 16'd38646, 16'd7659, 16'd13244, 16'd40206, 16'd20724, 16'd41721, 16'd37383, 16'd15064, 16'd62903, 16'd17867, 16'd7707, 16'd36787, 16'd38890, 16'd51129, 16'd6908, 16'd37103, 16'd21207, 16'd39625, 16'd53135, 16'd27091, 16'd21774, 16'd53766, 16'd2863, 16'd6936});
	test_expansion(128'h2340535d63ec2f0d1b8eeb2a7a469a4c, {16'd8012, 16'd42879, 16'd57037, 16'd33794, 16'd54941, 16'd58408, 16'd34585, 16'd39028, 16'd59298, 16'd56663, 16'd56536, 16'd52690, 16'd21067, 16'd65402, 16'd35324, 16'd15632, 16'd18400, 16'd64721, 16'd42446, 16'd54858, 16'd31154, 16'd3072, 16'd7103, 16'd58615, 16'd15113, 16'd29965});
	test_expansion(128'hf7287f9948e098c80e3f27d4066a6538, {16'd43724, 16'd46187, 16'd65197, 16'd10066, 16'd46398, 16'd3336, 16'd25091, 16'd19279, 16'd43391, 16'd26377, 16'd48237, 16'd4606, 16'd45354, 16'd24612, 16'd4982, 16'd18064, 16'd53493, 16'd36137, 16'd60448, 16'd35720, 16'd40267, 16'd8326, 16'd40783, 16'd9953, 16'd40405, 16'd40497});
	test_expansion(128'h3977af374edea2610130408660511c91, {16'd13682, 16'd47188, 16'd53922, 16'd47394, 16'd18905, 16'd47004, 16'd38870, 16'd13529, 16'd29773, 16'd13508, 16'd65525, 16'd44301, 16'd18381, 16'd21872, 16'd30961, 16'd23609, 16'd5884, 16'd24195, 16'd54885, 16'd26288, 16'd59649, 16'd2471, 16'd4656, 16'd44444, 16'd41488, 16'd54273});
	test_expansion(128'hcd2d8329a542fe76720592578c1ec3fc, {16'd14523, 16'd16177, 16'd18611, 16'd27047, 16'd13953, 16'd28336, 16'd65110, 16'd36097, 16'd49086, 16'd5565, 16'd18030, 16'd7734, 16'd45060, 16'd47864, 16'd23438, 16'd25724, 16'd21279, 16'd48632, 16'd54031, 16'd18411, 16'd15295, 16'd44691, 16'd4540, 16'd45060, 16'd12614, 16'd23366});
	test_expansion(128'h97597d1f98133baef5c2d053b15da935, {16'd36450, 16'd18234, 16'd53114, 16'd49011, 16'd22675, 16'd7368, 16'd13924, 16'd42000, 16'd24820, 16'd53302, 16'd63327, 16'd32012, 16'd1885, 16'd21589, 16'd62101, 16'd5702, 16'd28761, 16'd28484, 16'd40237, 16'd63631, 16'd50975, 16'd1370, 16'd29452, 16'd13530, 16'd31379, 16'd26521});
	test_expansion(128'h38709bdd09545bfcf68af7bf2fa17d52, {16'd50655, 16'd61208, 16'd54347, 16'd46597, 16'd51356, 16'd12049, 16'd51339, 16'd3429, 16'd8311, 16'd26788, 16'd11206, 16'd39943, 16'd42561, 16'd28638, 16'd15943, 16'd3624, 16'd31047, 16'd5844, 16'd3483, 16'd16798, 16'd12664, 16'd14570, 16'd8588, 16'd6122, 16'd21069, 16'd16612});
	test_expansion(128'h4221d2ee164074817c23c8cd7aea2295, {16'd19546, 16'd43238, 16'd58511, 16'd65437, 16'd59320, 16'd34247, 16'd44192, 16'd31351, 16'd7098, 16'd65409, 16'd32125, 16'd56463, 16'd58455, 16'd32662, 16'd54915, 16'd16520, 16'd31647, 16'd31827, 16'd61073, 16'd20417, 16'd59915, 16'd52682, 16'd17080, 16'd17893, 16'd47137, 16'd38882});
	test_expansion(128'hc76a530ed423e40832467902f0a7f926, {16'd44423, 16'd11084, 16'd50827, 16'd24719, 16'd2724, 16'd43990, 16'd13632, 16'd58885, 16'd15204, 16'd12209, 16'd45440, 16'd18187, 16'd4016, 16'd11853, 16'd37781, 16'd1005, 16'd698, 16'd9817, 16'd52202, 16'd59199, 16'd15049, 16'd23470, 16'd23030, 16'd25214, 16'd21224, 16'd26449});
	test_expansion(128'h1ca6064a3f5f106d0c2ac079251b0a26, {16'd7754, 16'd25341, 16'd40167, 16'd24270, 16'd19307, 16'd42251, 16'd43471, 16'd64208, 16'd64973, 16'd42184, 16'd42714, 16'd16184, 16'd57252, 16'd52746, 16'd63988, 16'd47539, 16'd13261, 16'd57138, 16'd59542, 16'd47038, 16'd31064, 16'd38091, 16'd33505, 16'd8976, 16'd53992, 16'd54500});
	test_expansion(128'h94eb11692c6fecb441cf08c85e51b6c4, {16'd50627, 16'd16179, 16'd46553, 16'd2336, 16'd9644, 16'd12803, 16'd61715, 16'd44503, 16'd47406, 16'd861, 16'd59860, 16'd41966, 16'd52259, 16'd3426, 16'd23208, 16'd344, 16'd20674, 16'd34224, 16'd29509, 16'd24767, 16'd24705, 16'd49753, 16'd48302, 16'd33851, 16'd58628, 16'd20390});
	test_expansion(128'h5fb54864dc589a9b5cd7beb37d637f69, {16'd3127, 16'd24636, 16'd31507, 16'd14983, 16'd21280, 16'd2731, 16'd57766, 16'd48732, 16'd8413, 16'd24140, 16'd24316, 16'd58296, 16'd8475, 16'd18701, 16'd27496, 16'd2137, 16'd32353, 16'd12235, 16'd60380, 16'd49460, 16'd535, 16'd3188, 16'd7343, 16'd23349, 16'd10847, 16'd25138});
	test_expansion(128'h249075a90dd217189026c2f3bee067ac, {16'd57786, 16'd63715, 16'd40571, 16'd46229, 16'd518, 16'd64977, 16'd62809, 16'd45852, 16'd18310, 16'd52366, 16'd27170, 16'd55006, 16'd31276, 16'd62603, 16'd64593, 16'd43074, 16'd24106, 16'd38251, 16'd18784, 16'd4379, 16'd49107, 16'd47764, 16'd48152, 16'd16930, 16'd1936, 16'd41387});
	test_expansion(128'hc86b45869679f03cbdf9fddd96a98807, {16'd54730, 16'd10187, 16'd59158, 16'd15651, 16'd12415, 16'd56916, 16'd51359, 16'd10131, 16'd45413, 16'd5991, 16'd7470, 16'd6705, 16'd26070, 16'd53546, 16'd30331, 16'd26931, 16'd8183, 16'd53742, 16'd31797, 16'd42053, 16'd12945, 16'd16182, 16'd18258, 16'd58857, 16'd45018, 16'd12556});
	test_expansion(128'h28a33e930c0873b072f50c07f68771c2, {16'd726, 16'd37556, 16'd32649, 16'd50446, 16'd47488, 16'd40771, 16'd15662, 16'd31914, 16'd27712, 16'd20673, 16'd30136, 16'd38131, 16'd55046, 16'd33416, 16'd51465, 16'd49592, 16'd63994, 16'd37540, 16'd25705, 16'd18052, 16'd21293, 16'd60312, 16'd42540, 16'd51517, 16'd22212, 16'd48954});
	test_expansion(128'h8e84081652673a7dcdc063f701c1ecb3, {16'd11779, 16'd2493, 16'd36705, 16'd25409, 16'd9129, 16'd41749, 16'd52674, 16'd1748, 16'd52624, 16'd50055, 16'd56858, 16'd27757, 16'd35704, 16'd15284, 16'd55112, 16'd40217, 16'd36727, 16'd12677, 16'd32197, 16'd54507, 16'd43039, 16'd60099, 16'd38766, 16'd49772, 16'd40015, 16'd63900});
	test_expansion(128'hb5f2ea39b92d2ba0183f927ac098808a, {16'd45637, 16'd22146, 16'd54827, 16'd44778, 16'd10420, 16'd22754, 16'd46282, 16'd40052, 16'd14438, 16'd48200, 16'd56975, 16'd2724, 16'd12089, 16'd11909, 16'd49973, 16'd54262, 16'd38086, 16'd22831, 16'd45173, 16'd37729, 16'd14879, 16'd8846, 16'd671, 16'd12544, 16'd18932, 16'd47860});
	test_expansion(128'hb97225b536144b114ba384741c3ca369, {16'd57321, 16'd12961, 16'd27796, 16'd259, 16'd39411, 16'd23756, 16'd11656, 16'd39451, 16'd37263, 16'd33129, 16'd21100, 16'd32130, 16'd59928, 16'd44474, 16'd15730, 16'd36424, 16'd35859, 16'd4501, 16'd36281, 16'd37311, 16'd33632, 16'd52292, 16'd2897, 16'd37347, 16'd58158, 16'd35706});
	test_expansion(128'h3c3cea044cdbcb34978d3d1500dfb1da, {16'd16423, 16'd17479, 16'd19700, 16'd41249, 16'd36452, 16'd64677, 16'd54736, 16'd42345, 16'd57637, 16'd17000, 16'd63652, 16'd26564, 16'd20369, 16'd24913, 16'd9619, 16'd48313, 16'd46167, 16'd13078, 16'd39526, 16'd2080, 16'd38049, 16'd40600, 16'd14126, 16'd65009, 16'd45373, 16'd33062});
	test_expansion(128'h9decaa6beb6df89ca3a3c638b1436e80, {16'd34144, 16'd36123, 16'd43675, 16'd21184, 16'd17044, 16'd13691, 16'd35832, 16'd14823, 16'd12761, 16'd34239, 16'd49802, 16'd32889, 16'd44051, 16'd15682, 16'd10766, 16'd44527, 16'd42333, 16'd3359, 16'd49274, 16'd18843, 16'd36272, 16'd13586, 16'd36234, 16'd64229, 16'd62308, 16'd5500});
	test_expansion(128'h5bd6dce42cf1988fde474b64b8fa1993, {16'd45172, 16'd57731, 16'd7522, 16'd40322, 16'd5950, 16'd27109, 16'd53847, 16'd56242, 16'd36241, 16'd49940, 16'd48156, 16'd34199, 16'd32356, 16'd4004, 16'd23645, 16'd48277, 16'd51249, 16'd48562, 16'd49304, 16'd2062, 16'd28351, 16'd60965, 16'd50231, 16'd32328, 16'd24122, 16'd43064});
	test_expansion(128'h0a9de0c452b181168563185bda520fce, {16'd36206, 16'd22624, 16'd60725, 16'd4492, 16'd56948, 16'd59653, 16'd42084, 16'd31367, 16'd2524, 16'd52391, 16'd41892, 16'd22199, 16'd43999, 16'd32488, 16'd65088, 16'd20695, 16'd38419, 16'd13564, 16'd39117, 16'd6781, 16'd44402, 16'd61587, 16'd42929, 16'd5414, 16'd54351, 16'd49662});
	test_expansion(128'hc56466ce4de6d6d0c33ffd65a87e9d60, {16'd25175, 16'd49413, 16'd25175, 16'd29060, 16'd27743, 16'd52297, 16'd7342, 16'd22873, 16'd59970, 16'd40944, 16'd42373, 16'd19880, 16'd22402, 16'd1634, 16'd48364, 16'd53355, 16'd29560, 16'd1431, 16'd30034, 16'd61074, 16'd28217, 16'd31496, 16'd28370, 16'd6505, 16'd61034, 16'd53652});
	test_expansion(128'h174e99ddee443043ab5b2db4e3b2a9b1, {16'd37544, 16'd28965, 16'd4558, 16'd24467, 16'd36826, 16'd10158, 16'd29544, 16'd9261, 16'd58197, 16'd5420, 16'd53545, 16'd21841, 16'd31721, 16'd56148, 16'd31230, 16'd28267, 16'd65043, 16'd56889, 16'd30308, 16'd39369, 16'd46847, 16'd61447, 16'd23551, 16'd18976, 16'd23574, 16'd5144});
	test_expansion(128'hf17e5eb5983752aac369b4d10d73abab, {16'd56833, 16'd6033, 16'd4437, 16'd39013, 16'd10850, 16'd51697, 16'd32261, 16'd60574, 16'd21143, 16'd27040, 16'd19467, 16'd40280, 16'd52782, 16'd32412, 16'd30262, 16'd3172, 16'd48825, 16'd12871, 16'd17010, 16'd25162, 16'd41641, 16'd33750, 16'd37336, 16'd15530, 16'd57832, 16'd41670});
	test_expansion(128'hdc0b173dfc30b7fd06a9e583ce4424dd, {16'd59785, 16'd58799, 16'd14821, 16'd60864, 16'd18931, 16'd54308, 16'd8057, 16'd19928, 16'd52894, 16'd31855, 16'd44665, 16'd29883, 16'd8931, 16'd55749, 16'd1965, 16'd9749, 16'd55484, 16'd20975, 16'd38219, 16'd65067, 16'd41890, 16'd51588, 16'd45609, 16'd24652, 16'd27954, 16'd22981});
	test_expansion(128'hdf6a207d590a20257a8867c7f5415152, {16'd34813, 16'd51841, 16'd16991, 16'd21657, 16'd47459, 16'd65025, 16'd42820, 16'd27414, 16'd59999, 16'd34292, 16'd63527, 16'd60199, 16'd10678, 16'd30420, 16'd1338, 16'd14499, 16'd24353, 16'd63585, 16'd11488, 16'd46826, 16'd12187, 16'd7239, 16'd25364, 16'd27675, 16'd47040, 16'd49423});
	test_expansion(128'h03d5a30c9d899e37545ed3c33e4b13b5, {16'd59040, 16'd59713, 16'd2277, 16'd8093, 16'd6167, 16'd33531, 16'd61878, 16'd25569, 16'd22279, 16'd38233, 16'd49306, 16'd48803, 16'd24364, 16'd1471, 16'd1537, 16'd18945, 16'd10218, 16'd2190, 16'd65007, 16'd1675, 16'd50262, 16'd40930, 16'd27081, 16'd1543, 16'd44576, 16'd47610});
	test_expansion(128'hb98a864a65430cc81d4bde5099e5b54d, {16'd60253, 16'd14532, 16'd52357, 16'd1744, 16'd44376, 16'd9132, 16'd35046, 16'd33697, 16'd28870, 16'd56047, 16'd44083, 16'd46866, 16'd18578, 16'd5051, 16'd3464, 16'd48404, 16'd21118, 16'd8832, 16'd57044, 16'd10317, 16'd54348, 16'd60393, 16'd55411, 16'd54888, 16'd35258, 16'd63043});
	test_expansion(128'hf3ebaeabb95a912e4b3529306ac80854, {16'd51223, 16'd43109, 16'd4146, 16'd23680, 16'd2084, 16'd32986, 16'd44153, 16'd62792, 16'd40698, 16'd64661, 16'd22009, 16'd63971, 16'd34833, 16'd53742, 16'd20765, 16'd57510, 16'd668, 16'd55426, 16'd49605, 16'd57209, 16'd49933, 16'd64872, 16'd32753, 16'd59863, 16'd32848, 16'd60679});
	test_expansion(128'h84696e99087f073d07fa730832bc0777, {16'd15477, 16'd55356, 16'd37388, 16'd30734, 16'd63691, 16'd28271, 16'd39348, 16'd26606, 16'd40815, 16'd43786, 16'd56049, 16'd40498, 16'd16030, 16'd18243, 16'd33493, 16'd18286, 16'd48691, 16'd12580, 16'd45495, 16'd21086, 16'd42965, 16'd64357, 16'd42584, 16'd56386, 16'd17836, 16'd21459});
	test_expansion(128'h320ccccd84b992b490926b7526994611, {16'd25017, 16'd33181, 16'd32036, 16'd42102, 16'd11938, 16'd14552, 16'd29106, 16'd28103, 16'd21563, 16'd5352, 16'd37027, 16'd1037, 16'd56653, 16'd48575, 16'd46621, 16'd47495, 16'd60006, 16'd27480, 16'd8279, 16'd46523, 16'd24235, 16'd4386, 16'd53397, 16'd22096, 16'd5356, 16'd57607});
	test_expansion(128'h95c928b492a6e9791f2145fa2fc1823b, {16'd46196, 16'd32718, 16'd11772, 16'd34906, 16'd10306, 16'd34917, 16'd1140, 16'd42610, 16'd9179, 16'd25356, 16'd26363, 16'd19928, 16'd31009, 16'd9766, 16'd12134, 16'd14536, 16'd58213, 16'd379, 16'd43758, 16'd42500, 16'd45258, 16'd58730, 16'd29350, 16'd61788, 16'd65301, 16'd20329});
	test_expansion(128'h30c64f6a33471f2ed3a9213073722bc3, {16'd12785, 16'd30202, 16'd28266, 16'd34819, 16'd15876, 16'd34489, 16'd2377, 16'd48195, 16'd17030, 16'd64353, 16'd21923, 16'd214, 16'd30996, 16'd41314, 16'd39264, 16'd48214, 16'd29666, 16'd5452, 16'd36213, 16'd2871, 16'd54282, 16'd12093, 16'd19226, 16'd39604, 16'd29124, 16'd9421});
	test_expansion(128'h44a7fb206d7f30c358226bef7aafeabb, {16'd64072, 16'd60745, 16'd2798, 16'd38726, 16'd54130, 16'd19718, 16'd29809, 16'd36650, 16'd14286, 16'd33106, 16'd15112, 16'd59755, 16'd40388, 16'd12593, 16'd41536, 16'd11249, 16'd45986, 16'd49846, 16'd16132, 16'd34916, 16'd14200, 16'd32058, 16'd61232, 16'd6312, 16'd48377, 16'd26823});
	test_expansion(128'h6b29de706043e0c070cb63830089ce22, {16'd13833, 16'd30793, 16'd53176, 16'd38826, 16'd62698, 16'd715, 16'd52360, 16'd55250, 16'd13172, 16'd17169, 16'd5411, 16'd7125, 16'd48592, 16'd38439, 16'd20737, 16'd9010, 16'd57201, 16'd27215, 16'd18854, 16'd38254, 16'd698, 16'd43650, 16'd46309, 16'd11295, 16'd31977, 16'd20479});
	test_expansion(128'hc525895d247579856dce9c2be216618d, {16'd46763, 16'd18767, 16'd241, 16'd62820, 16'd40598, 16'd24222, 16'd60788, 16'd32214, 16'd42245, 16'd49804, 16'd31086, 16'd53854, 16'd32686, 16'd31482, 16'd31372, 16'd49497, 16'd54152, 16'd62361, 16'd11896, 16'd47130, 16'd55659, 16'd24262, 16'd8377, 16'd63283, 16'd52160, 16'd51063});
	test_expansion(128'hf878e8455eacfe5ab60afd9f3924bcc7, {16'd40172, 16'd38679, 16'd6495, 16'd56340, 16'd60885, 16'd16384, 16'd36849, 16'd64103, 16'd32304, 16'd65408, 16'd56960, 16'd16055, 16'd37692, 16'd31029, 16'd59583, 16'd44816, 16'd122, 16'd46982, 16'd42400, 16'd64535, 16'd18755, 16'd63668, 16'd21747, 16'd64869, 16'd47722, 16'd37368});
	test_expansion(128'hc40146c2b8184acf4799846b6b14c063, {16'd44548, 16'd3130, 16'd55287, 16'd46756, 16'd21069, 16'd33843, 16'd61540, 16'd18057, 16'd10322, 16'd21904, 16'd22675, 16'd62564, 16'd22381, 16'd1235, 16'd11466, 16'd57470, 16'd39551, 16'd31019, 16'd57873, 16'd5690, 16'd32964, 16'd60015, 16'd36240, 16'd30140, 16'd55715, 16'd45289});
	test_expansion(128'hb0f68deed69773961ac6422ecf5e1481, {16'd48171, 16'd63912, 16'd21906, 16'd53200, 16'd31105, 16'd4660, 16'd22243, 16'd1147, 16'd27498, 16'd54030, 16'd52009, 16'd39662, 16'd49493, 16'd1514, 16'd41756, 16'd24276, 16'd27651, 16'd3233, 16'd26891, 16'd9432, 16'd38269, 16'd52229, 16'd9785, 16'd28375, 16'd34829, 16'd21251});
	test_expansion(128'h0ddccd6d450bbfd0bd1144d47b03834a, {16'd32545, 16'd54403, 16'd48642, 16'd13941, 16'd52949, 16'd26923, 16'd6217, 16'd4888, 16'd53711, 16'd36111, 16'd18035, 16'd1487, 16'd3041, 16'd1971, 16'd45324, 16'd34118, 16'd19632, 16'd61015, 16'd63396, 16'd30879, 16'd49815, 16'd13160, 16'd20118, 16'd38761, 16'd50392, 16'd47889});
	test_expansion(128'he8dd71f9ad3bf871173cc95cf5afafb8, {16'd37311, 16'd5233, 16'd26850, 16'd25762, 16'd2301, 16'd29608, 16'd25189, 16'd22452, 16'd7099, 16'd51244, 16'd7147, 16'd7029, 16'd27227, 16'd43553, 16'd35720, 16'd30797, 16'd42801, 16'd47502, 16'd40988, 16'd19121, 16'd17613, 16'd32353, 16'd48641, 16'd33423, 16'd24954, 16'd10305});
	test_expansion(128'hac7bd40f9b64a4c735515297d8dfa4bc, {16'd56136, 16'd20814, 16'd11065, 16'd37590, 16'd19627, 16'd47250, 16'd47378, 16'd1666, 16'd30461, 16'd24687, 16'd31885, 16'd49667, 16'd31219, 16'd28554, 16'd43450, 16'd6922, 16'd56078, 16'd61778, 16'd1458, 16'd59344, 16'd47235, 16'd446, 16'd24887, 16'd13533, 16'd9749, 16'd59412});
	test_expansion(128'hd2636a27e1dd529ab49194b4ec24bc1a, {16'd32986, 16'd31713, 16'd13806, 16'd19153, 16'd30339, 16'd47736, 16'd25362, 16'd27630, 16'd17539, 16'd35617, 16'd45331, 16'd29227, 16'd23287, 16'd15393, 16'd19468, 16'd62859, 16'd34550, 16'd31234, 16'd7883, 16'd7017, 16'd52483, 16'd61435, 16'd53968, 16'd22394, 16'd37113, 16'd26599});
	test_expansion(128'hf9ac70d913ee076fa8a94ca095fdae44, {16'd52676, 16'd19265, 16'd61434, 16'd54724, 16'd25984, 16'd17942, 16'd55375, 16'd40395, 16'd19331, 16'd25513, 16'd26342, 16'd9828, 16'd24198, 16'd26331, 16'd38974, 16'd18267, 16'd28788, 16'd59217, 16'd22292, 16'd29203, 16'd39586, 16'd28472, 16'd52987, 16'd7078, 16'd36258, 16'd14889});
	test_expansion(128'h777a0a66e2c9dc598c9c5f38fada0a5f, {16'd44600, 16'd30694, 16'd38470, 16'd7789, 16'd6379, 16'd36192, 16'd20263, 16'd38005, 16'd888, 16'd58416, 16'd29095, 16'd22419, 16'd47723, 16'd41062, 16'd21117, 16'd38567, 16'd15346, 16'd40284, 16'd15605, 16'd57291, 16'd37062, 16'd32605, 16'd31399, 16'd41815, 16'd62870, 16'd62023});
	test_expansion(128'h8e5cd28c8823bc70eed4faae3e5bc985, {16'd30304, 16'd65419, 16'd5628, 16'd35374, 16'd2651, 16'd40407, 16'd61747, 16'd6778, 16'd24255, 16'd315, 16'd9212, 16'd40444, 16'd25510, 16'd23570, 16'd33986, 16'd31315, 16'd43005, 16'd6810, 16'd9269, 16'd53129, 16'd7333, 16'd2961, 16'd33073, 16'd24302, 16'd20490, 16'd15894});
	test_expansion(128'h98db4b25454f85b4b14cac1477160a43, {16'd20828, 16'd41474, 16'd29133, 16'd51968, 16'd61276, 16'd30627, 16'd8786, 16'd63031, 16'd8552, 16'd62970, 16'd64023, 16'd63963, 16'd61634, 16'd41275, 16'd32344, 16'd14574, 16'd23318, 16'd4247, 16'd64221, 16'd43442, 16'd2939, 16'd40065, 16'd26279, 16'd15922, 16'd34543, 16'd20467});
	test_expansion(128'h24d349fa88afd27d6c97bcb765dc5212, {16'd48390, 16'd49128, 16'd46753, 16'd20422, 16'd1519, 16'd9489, 16'd19273, 16'd33705, 16'd13581, 16'd23626, 16'd44237, 16'd15995, 16'd40408, 16'd10784, 16'd45774, 16'd515, 16'd14970, 16'd9278, 16'd33789, 16'd5728, 16'd43085, 16'd5929, 16'd23873, 16'd48332, 16'd29203, 16'd28066});
	test_expansion(128'h949554921ef2310f33b6cb4b2b942793, {16'd12073, 16'd11304, 16'd51121, 16'd55647, 16'd46447, 16'd30990, 16'd41431, 16'd50259, 16'd24082, 16'd48585, 16'd28474, 16'd5056, 16'd31319, 16'd16146, 16'd51211, 16'd26122, 16'd53316, 16'd7376, 16'd33856, 16'd12634, 16'd26123, 16'd45009, 16'd22043, 16'd39434, 16'd3711, 16'd59267});
	test_expansion(128'hc3060655534efd19e3677dbd245828f4, {16'd16507, 16'd61698, 16'd49596, 16'd51533, 16'd15985, 16'd17764, 16'd38868, 16'd29830, 16'd39201, 16'd16726, 16'd6966, 16'd19177, 16'd20171, 16'd42093, 16'd1306, 16'd35900, 16'd35992, 16'd33428, 16'd29608, 16'd24516, 16'd13480, 16'd55328, 16'd47905, 16'd35169, 16'd61671, 16'd42578});
	test_expansion(128'h20df4e0afcb71bd92a66c15578ba9f1c, {16'd43442, 16'd16862, 16'd33886, 16'd42667, 16'd46785, 16'd49789, 16'd45553, 16'd62689, 16'd60192, 16'd65411, 16'd19344, 16'd9340, 16'd55530, 16'd22257, 16'd63782, 16'd35388, 16'd54370, 16'd50108, 16'd2274, 16'd60078, 16'd10238, 16'd17831, 16'd4583, 16'd43573, 16'd22254, 16'd28012});
	test_expansion(128'hb8426ffa18a55fea19439c6175870bd2, {16'd10635, 16'd54619, 16'd26649, 16'd40388, 16'd16538, 16'd44685, 16'd54412, 16'd46842, 16'd44562, 16'd41429, 16'd23869, 16'd2145, 16'd13995, 16'd47209, 16'd8341, 16'd12549, 16'd34721, 16'd50004, 16'd19445, 16'd31047, 16'd65355, 16'd18547, 16'd46637, 16'd14128, 16'd45049, 16'd15474});
	test_expansion(128'h629fd80ca00e5906be00fd41927df6b6, {16'd15345, 16'd64535, 16'd55085, 16'd128, 16'd44788, 16'd60046, 16'd45212, 16'd37402, 16'd2552, 16'd62331, 16'd1603, 16'd31875, 16'd41023, 16'd19255, 16'd17585, 16'd6795, 16'd23022, 16'd41141, 16'd52627, 16'd2940, 16'd28037, 16'd17484, 16'd16052, 16'd53056, 16'd42469, 16'd17201});
	test_expansion(128'haa1e3a3bc7ea5c0c5e0264012e69eeb9, {16'd69, 16'd30189, 16'd207, 16'd2597, 16'd30445, 16'd15851, 16'd14085, 16'd26762, 16'd18660, 16'd53191, 16'd16882, 16'd15394, 16'd39671, 16'd12924, 16'd19550, 16'd1094, 16'd7714, 16'd35191, 16'd19364, 16'd63090, 16'd6214, 16'd8337, 16'd7935, 16'd53981, 16'd44122, 16'd22333});
	test_expansion(128'h90abece967ee890aa2947fe6ac02a6e1, {16'd30924, 16'd52066, 16'd21687, 16'd2479, 16'd12370, 16'd60899, 16'd41509, 16'd26630, 16'd39352, 16'd2125, 16'd33674, 16'd36328, 16'd35262, 16'd51280, 16'd43874, 16'd21830, 16'd55910, 16'd40265, 16'd47036, 16'd10293, 16'd687, 16'd46217, 16'd49392, 16'd57173, 16'd53571, 16'd36181});
	test_expansion(128'h4b649c9a2660290f3ff961f31419ce35, {16'd31098, 16'd63447, 16'd1487, 16'd26756, 16'd62567, 16'd10159, 16'd5220, 16'd60914, 16'd7495, 16'd41772, 16'd29709, 16'd32506, 16'd53006, 16'd21259, 16'd44927, 16'd25212, 16'd13243, 16'd56418, 16'd57364, 16'd5867, 16'd63275, 16'd41329, 16'd47947, 16'd20538, 16'd1150, 16'd55106});
	test_expansion(128'h97a6024327b8ea9df78509ddd775b848, {16'd45346, 16'd49040, 16'd4073, 16'd54818, 16'd51447, 16'd21136, 16'd17304, 16'd34742, 16'd40412, 16'd58997, 16'd54789, 16'd2684, 16'd32165, 16'd48619, 16'd4114, 16'd23974, 16'd3104, 16'd10819, 16'd63729, 16'd55011, 16'd53050, 16'd28998, 16'd50085, 16'd60655, 16'd37408, 16'd17550});
	test_expansion(128'h9f65e2c70fb41dd8db47ca745428d191, {16'd57830, 16'd16115, 16'd34308, 16'd32156, 16'd12616, 16'd218, 16'd57816, 16'd3885, 16'd12206, 16'd48766, 16'd65321, 16'd14786, 16'd19809, 16'd37368, 16'd65324, 16'd10049, 16'd35329, 16'd48846, 16'd18861, 16'd7070, 16'd17701, 16'd1380, 16'd42306, 16'd34544, 16'd53611, 16'd42069});
	test_expansion(128'h8662848b71f2ab5dcc27a0f22666fe7e, {16'd24003, 16'd40061, 16'd54887, 16'd62327, 16'd58993, 16'd58534, 16'd37208, 16'd55530, 16'd16454, 16'd32156, 16'd27675, 16'd36309, 16'd18202, 16'd64655, 16'd38994, 16'd60268, 16'd26066, 16'd1268, 16'd56986, 16'd35327, 16'd60597, 16'd52439, 16'd47760, 16'd2574, 16'd62355, 16'd44580});
	test_expansion(128'hec4f9fcc9c708b9c8d6e912b62060b32, {16'd35508, 16'd60427, 16'd13436, 16'd62145, 16'd69, 16'd36628, 16'd39042, 16'd8418, 16'd57088, 16'd43313, 16'd42279, 16'd64847, 16'd48491, 16'd64816, 16'd43261, 16'd15061, 16'd6514, 16'd58727, 16'd53324, 16'd50458, 16'd41060, 16'd49227, 16'd65300, 16'd58426, 16'd34002, 16'd19206});
	test_expansion(128'hb0cd4f51eb9bc4a418dd1be20e960811, {16'd11047, 16'd35629, 16'd61597, 16'd10601, 16'd11357, 16'd2570, 16'd58469, 16'd2782, 16'd29432, 16'd46677, 16'd15831, 16'd8334, 16'd25002, 16'd1295, 16'd57860, 16'd25176, 16'd44919, 16'd34766, 16'd31628, 16'd52948, 16'd21890, 16'd49798, 16'd57488, 16'd27900, 16'd9814, 16'd13926});
	test_expansion(128'h7bc003512ef08a8e070e4aef2abb97c7, {16'd40511, 16'd12833, 16'd47128, 16'd24053, 16'd16865, 16'd14286, 16'd55280, 16'd23793, 16'd54086, 16'd36245, 16'd25248, 16'd44669, 16'd11117, 16'd45734, 16'd7700, 16'd49333, 16'd32649, 16'd40947, 16'd49272, 16'd42898, 16'd3237, 16'd29457, 16'd5850, 16'd58086, 16'd25740, 16'd33425});
	test_expansion(128'h9b22da8a81990f8aaa55ae04e08b2ad2, {16'd38567, 16'd21002, 16'd62782, 16'd29595, 16'd7797, 16'd34689, 16'd61007, 16'd64966, 16'd51384, 16'd54922, 16'd58752, 16'd24167, 16'd60353, 16'd17201, 16'd6545, 16'd25542, 16'd13822, 16'd54748, 16'd21020, 16'd38853, 16'd27300, 16'd31855, 16'd5207, 16'd50601, 16'd13104, 16'd41317});
	test_expansion(128'h16e3544a85537a5ae993af2f7d2fa05b, {16'd29716, 16'd12345, 16'd65090, 16'd17549, 16'd5761, 16'd27919, 16'd536, 16'd37798, 16'd54023, 16'd46418, 16'd18684, 16'd22387, 16'd17465, 16'd63464, 16'd36167, 16'd52335, 16'd44062, 16'd31108, 16'd28898, 16'd20512, 16'd5680, 16'd34920, 16'd47166, 16'd45036, 16'd34753, 16'd12106});
	test_expansion(128'h3d04eb0d6943b3258664d9ae57bea2fb, {16'd25646, 16'd38190, 16'd58130, 16'd1561, 16'd61334, 16'd30009, 16'd6318, 16'd50296, 16'd42477, 16'd29618, 16'd11611, 16'd16401, 16'd16046, 16'd43156, 16'd60569, 16'd47520, 16'd49073, 16'd17638, 16'd28143, 16'd17602, 16'd39578, 16'd5474, 16'd13699, 16'd44987, 16'd55790, 16'd62248});
	test_expansion(128'h676099a5b3b4e3778dbfb04ea22afaca, {16'd11887, 16'd17867, 16'd19579, 16'd21438, 16'd31059, 16'd45681, 16'd25767, 16'd33826, 16'd61402, 16'd64222, 16'd6141, 16'd22671, 16'd40216, 16'd39647, 16'd48651, 16'd46880, 16'd7783, 16'd16315, 16'd10486, 16'd21024, 16'd30920, 16'd10687, 16'd63351, 16'd25424, 16'd61217, 16'd3594});
	test_expansion(128'h13e22dab8eac8e22787262873e6baf72, {16'd6283, 16'd25724, 16'd41931, 16'd33832, 16'd57560, 16'd2851, 16'd56482, 16'd34969, 16'd13103, 16'd5400, 16'd11330, 16'd2566, 16'd52040, 16'd5144, 16'd1060, 16'd1585, 16'd38524, 16'd50953, 16'd52655, 16'd40314, 16'd56740, 16'd35934, 16'd10913, 16'd42967, 16'd38043, 16'd37591});
	test_expansion(128'h1993ebddda511a4147df15f9a2a9e260, {16'd51627, 16'd41336, 16'd56569, 16'd63795, 16'd52546, 16'd6018, 16'd14661, 16'd8368, 16'd4697, 16'd55117, 16'd15668, 16'd36976, 16'd11244, 16'd6179, 16'd25359, 16'd10178, 16'd37264, 16'd53417, 16'd38104, 16'd56511, 16'd17016, 16'd2492, 16'd18164, 16'd51709, 16'd28450, 16'd55922});
	test_expansion(128'h83d518bf61b7545dd029955cf23fe081, {16'd58828, 16'd33135, 16'd12176, 16'd23921, 16'd57951, 16'd15501, 16'd63892, 16'd62122, 16'd31543, 16'd58843, 16'd26865, 16'd39679, 16'd51533, 16'd58075, 16'd45583, 16'd8034, 16'd54839, 16'd40978, 16'd1399, 16'd58420, 16'd4218, 16'd12655, 16'd48154, 16'd9257, 16'd62212, 16'd59043});
	test_expansion(128'h69f4dd685ff38dc391b4d4beecc3e55e, {16'd12699, 16'd52734, 16'd29786, 16'd33261, 16'd41653, 16'd4422, 16'd55061, 16'd2695, 16'd30129, 16'd29571, 16'd37288, 16'd40135, 16'd60387, 16'd25259, 16'd37873, 16'd22272, 16'd57418, 16'd49837, 16'd47956, 16'd25604, 16'd43441, 16'd24791, 16'd48776, 16'd44673, 16'd9718, 16'd13514});
	test_expansion(128'h6f0bbc6afacf1bee44c4fa3794abb270, {16'd48855, 16'd11921, 16'd60139, 16'd56524, 16'd47227, 16'd52118, 16'd35412, 16'd32251, 16'd41719, 16'd8619, 16'd13558, 16'd6116, 16'd33862, 16'd35242, 16'd64518, 16'd13783, 16'd29976, 16'd40693, 16'd7507, 16'd6470, 16'd39347, 16'd4729, 16'd53790, 16'd40565, 16'd38227, 16'd47421});
	test_expansion(128'h7b33ba938ae6d0796fd313ab8d83f5a2, {16'd34623, 16'd50734, 16'd62656, 16'd15961, 16'd54968, 16'd41221, 16'd7366, 16'd9841, 16'd23766, 16'd63273, 16'd40079, 16'd20430, 16'd30024, 16'd19375, 16'd34004, 16'd4538, 16'd12191, 16'd52766, 16'd46911, 16'd31380, 16'd53457, 16'd12024, 16'd7669, 16'd1974, 16'd37860, 16'd31133});
	test_expansion(128'h1b1816276382f4bfb55901d42efa74bc, {16'd38132, 16'd29909, 16'd30537, 16'd43938, 16'd37742, 16'd19711, 16'd17981, 16'd50217, 16'd42870, 16'd50476, 16'd55075, 16'd32497, 16'd59151, 16'd4046, 16'd15269, 16'd59545, 16'd17625, 16'd53509, 16'd58881, 16'd62974, 16'd33563, 16'd16572, 16'd27492, 16'd4364, 16'd21801, 16'd47730});
	test_expansion(128'h1d9be146fc6a26cd329fdd3d3c6a8871, {16'd44337, 16'd44703, 16'd387, 16'd19750, 16'd5635, 16'd31492, 16'd12005, 16'd30407, 16'd62755, 16'd6630, 16'd17593, 16'd39279, 16'd5217, 16'd11566, 16'd45159, 16'd59730, 16'd47060, 16'd47082, 16'd38673, 16'd11235, 16'd32655, 16'd5443, 16'd30757, 16'd3599, 16'd29403, 16'd64842});
	test_expansion(128'h3cb7cbf5809704ca906100e4ed360574, {16'd6342, 16'd31682, 16'd64603, 16'd10094, 16'd36466, 16'd21036, 16'd9607, 16'd18603, 16'd39127, 16'd2911, 16'd58560, 16'd34284, 16'd55963, 16'd14404, 16'd42562, 16'd25889, 16'd45722, 16'd9496, 16'd14678, 16'd61438, 16'd21493, 16'd33863, 16'd28284, 16'd26733, 16'd35932, 16'd57489});
	test_expansion(128'h5576d6b1e8f187d3301d8b24514827d3, {16'd4508, 16'd526, 16'd7760, 16'd58348, 16'd21032, 16'd4641, 16'd15324, 16'd28950, 16'd1133, 16'd58416, 16'd59814, 16'd62019, 16'd46977, 16'd26625, 16'd57304, 16'd13458, 16'd16109, 16'd30524, 16'd21039, 16'd42300, 16'd25774, 16'd59338, 16'd15190, 16'd38927, 16'd43428, 16'd42607});
	test_expansion(128'h55c517f58461a2b2459bc8caa9e70639, {16'd48378, 16'd34553, 16'd9150, 16'd7448, 16'd6636, 16'd24738, 16'd56437, 16'd16650, 16'd45512, 16'd55174, 16'd7982, 16'd59635, 16'd12057, 16'd7728, 16'd65258, 16'd13611, 16'd13793, 16'd37205, 16'd64030, 16'd5784, 16'd10094, 16'd12679, 16'd16834, 16'd14741, 16'd12777, 16'd16445});
	test_expansion(128'hb1ef96f7c48600dbe1d421a96c2b4834, {16'd13504, 16'd65266, 16'd34106, 16'd64931, 16'd63102, 16'd38490, 16'd23436, 16'd32522, 16'd19272, 16'd6929, 16'd18426, 16'd49834, 16'd21444, 16'd1705, 16'd34375, 16'd20801, 16'd20044, 16'd52116, 16'd2183, 16'd60870, 16'd19157, 16'd28683, 16'd14922, 16'd3642, 16'd44771, 16'd15900});
	test_expansion(128'h797284b7a291563228330917a00b5fdd, {16'd5670, 16'd17676, 16'd9140, 16'd50384, 16'd5826, 16'd63478, 16'd2095, 16'd52645, 16'd50936, 16'd64053, 16'd24058, 16'd7987, 16'd10371, 16'd7764, 16'd63581, 16'd48711, 16'd39871, 16'd53397, 16'd32297, 16'd33181, 16'd17457, 16'd29829, 16'd55456, 16'd50832, 16'd32235, 16'd63458});
	test_expansion(128'h35cf2ee3bb0c4892caf88cc7260423a6, {16'd23153, 16'd17263, 16'd56017, 16'd51491, 16'd19390, 16'd55847, 16'd34982, 16'd35104, 16'd29605, 16'd61508, 16'd56891, 16'd55198, 16'd4425, 16'd23839, 16'd29523, 16'd27717, 16'd64476, 16'd53188, 16'd63864, 16'd12769, 16'd4250, 16'd21181, 16'd38808, 16'd53376, 16'd4975, 16'd23372});
	test_expansion(128'h34c206443c8548ac0f50aa4fa19226a1, {16'd24653, 16'd12657, 16'd38841, 16'd7392, 16'd30890, 16'd31199, 16'd1353, 16'd58610, 16'd19209, 16'd22215, 16'd58193, 16'd62224, 16'd29359, 16'd13153, 16'd52803, 16'd39895, 16'd19927, 16'd8360, 16'd38931, 16'd56385, 16'd5086, 16'd28841, 16'd26397, 16'd42134, 16'd9352, 16'd34795});
	test_expansion(128'h464134516b3e74b72b794fdcd77c96f0, {16'd29682, 16'd58553, 16'd47573, 16'd8656, 16'd12205, 16'd30479, 16'd25574, 16'd17333, 16'd37992, 16'd26703, 16'd29621, 16'd22907, 16'd11934, 16'd36208, 16'd37074, 16'd10349, 16'd47327, 16'd54295, 16'd17432, 16'd47995, 16'd36806, 16'd27298, 16'd41068, 16'd40472, 16'd17458, 16'd52240});
	test_expansion(128'hd08b0e121384057441e59c9d1dee7f55, {16'd41645, 16'd52369, 16'd52404, 16'd50313, 16'd53080, 16'd39302, 16'd31470, 16'd23790, 16'd49656, 16'd40128, 16'd33574, 16'd15694, 16'd24391, 16'd19556, 16'd31236, 16'd44602, 16'd14757, 16'd43601, 16'd63189, 16'd25558, 16'd46875, 16'd54083, 16'd18827, 16'd34749, 16'd59142, 16'd29722});
	test_expansion(128'h0fc56a972ef1746cf6b57772ad603fb2, {16'd17327, 16'd44561, 16'd4628, 16'd38937, 16'd35984, 16'd14193, 16'd43116, 16'd9599, 16'd48557, 16'd39545, 16'd45119, 16'd24455, 16'd12467, 16'd16033, 16'd30758, 16'd16900, 16'd32193, 16'd39948, 16'd5005, 16'd45652, 16'd12494, 16'd46436, 16'd60654, 16'd2356, 16'd38273, 16'd7448});
	test_expansion(128'ha60820c44879035087624e7a7145ee9c, {16'd48807, 16'd6148, 16'd61145, 16'd29346, 16'd64248, 16'd56182, 16'd40993, 16'd15174, 16'd44353, 16'd21641, 16'd22259, 16'd45909, 16'd7630, 16'd24903, 16'd6748, 16'd40158, 16'd238, 16'd23500, 16'd43333, 16'd30887, 16'd34819, 16'd37444, 16'd29628, 16'd47089, 16'd12807, 16'd32916});
	test_expansion(128'he25040dedf1a09a61d28fcecb8e0bc7f, {16'd54885, 16'd50228, 16'd51144, 16'd61207, 16'd24702, 16'd12807, 16'd6185, 16'd3785, 16'd43885, 16'd8118, 16'd59535, 16'd53596, 16'd57382, 16'd11062, 16'd39059, 16'd50165, 16'd14800, 16'd30724, 16'd15030, 16'd64098, 16'd43640, 16'd19640, 16'd509, 16'd579, 16'd21456, 16'd39427});
	test_expansion(128'hd3d21508d126b871ae7a2859d704b566, {16'd23215, 16'd16323, 16'd1326, 16'd3356, 16'd57233, 16'd17400, 16'd19847, 16'd22009, 16'd37844, 16'd36342, 16'd36800, 16'd30536, 16'd33816, 16'd25731, 16'd8327, 16'd2857, 16'd6331, 16'd16834, 16'd11688, 16'd33278, 16'd43548, 16'd13428, 16'd53529, 16'd34079, 16'd47885, 16'd24267});
	test_expansion(128'h15ff464a22de2012bec803e23e574106, {16'd8933, 16'd6942, 16'd17083, 16'd63747, 16'd57275, 16'd15834, 16'd15693, 16'd52430, 16'd26301, 16'd42796, 16'd32722, 16'd20720, 16'd15031, 16'd25725, 16'd2925, 16'd60647, 16'd11720, 16'd52142, 16'd35833, 16'd58134, 16'd35542, 16'd7455, 16'd63707, 16'd26547, 16'd61300, 16'd12234});
	test_expansion(128'hcdfdb486746adf3b756b5473a2e8830d, {16'd17773, 16'd59331, 16'd51310, 16'd7996, 16'd47686, 16'd31667, 16'd55353, 16'd9710, 16'd61205, 16'd31274, 16'd12423, 16'd16367, 16'd17158, 16'd31036, 16'd14746, 16'd12006, 16'd37555, 16'd6898, 16'd52198, 16'd35926, 16'd15429, 16'd35805, 16'd28200, 16'd36432, 16'd36736, 16'd22244});
	test_expansion(128'h3f4fc3bd374d1f2f58360c69793ae0f1, {16'd52256, 16'd1988, 16'd26836, 16'd2751, 16'd63652, 16'd19483, 16'd7835, 16'd51755, 16'd42509, 16'd24010, 16'd33844, 16'd35608, 16'd46407, 16'd8752, 16'd59299, 16'd48143, 16'd50581, 16'd39607, 16'd58772, 16'd4299, 16'd16443, 16'd56954, 16'd13635, 16'd34086, 16'd15921, 16'd21571});
	test_expansion(128'hcff496bc3f5293900f13577bd165cf7a, {16'd18424, 16'd59261, 16'd49605, 16'd61594, 16'd36798, 16'd50043, 16'd41634, 16'd40546, 16'd23069, 16'd2944, 16'd19628, 16'd22229, 16'd51230, 16'd38337, 16'd39450, 16'd42323, 16'd32453, 16'd42872, 16'd33606, 16'd39724, 16'd54110, 16'd13342, 16'd5442, 16'd35083, 16'd28827, 16'd24892});
	test_expansion(128'ha70dcf8dcd1c0c4c7c4ce0d9464fc126, {16'd4724, 16'd48114, 16'd55473, 16'd4545, 16'd58473, 16'd57367, 16'd62447, 16'd20988, 16'd49370, 16'd14155, 16'd13454, 16'd19037, 16'd3110, 16'd35213, 16'd12509, 16'd39080, 16'd62372, 16'd49528, 16'd63780, 16'd38107, 16'd14334, 16'd53465, 16'd22391, 16'd23020, 16'd42912, 16'd16303});
	test_expansion(128'h2574988d7f1f736b998f7d38349bb30c, {16'd31356, 16'd1657, 16'd23426, 16'd20072, 16'd12571, 16'd22429, 16'd59509, 16'd24090, 16'd17719, 16'd36219, 16'd5174, 16'd62276, 16'd52355, 16'd63292, 16'd3122, 16'd21666, 16'd24181, 16'd62712, 16'd5208, 16'd42784, 16'd40337, 16'd20957, 16'd27549, 16'd7133, 16'd47721, 16'd41877});
	test_expansion(128'h52cb645ef180ad85ba87c41194eea91d, {16'd37222, 16'd52761, 16'd6912, 16'd55085, 16'd21506, 16'd58398, 16'd53777, 16'd19133, 16'd55710, 16'd19626, 16'd56345, 16'd2807, 16'd26289, 16'd1863, 16'd37007, 16'd57909, 16'd62050, 16'd37354, 16'd37838, 16'd47888, 16'd38619, 16'd14548, 16'd50524, 16'd21901, 16'd34706, 16'd30009});
	test_expansion(128'h8fd6d18473cabe1652aa39feba740d76, {16'd37841, 16'd8009, 16'd16326, 16'd35752, 16'd20322, 16'd62827, 16'd35882, 16'd47658, 16'd53654, 16'd22514, 16'd38052, 16'd51014, 16'd42715, 16'd58178, 16'd8957, 16'd34538, 16'd54459, 16'd6146, 16'd62225, 16'd43513, 16'd23828, 16'd31804, 16'd45632, 16'd32093, 16'd766, 16'd32291});
	test_expansion(128'h728cb93d1251274280a8c85c182f4f35, {16'd36614, 16'd50739, 16'd21134, 16'd49955, 16'd4392, 16'd20249, 16'd12982, 16'd59290, 16'd1638, 16'd63551, 16'd22601, 16'd23209, 16'd8527, 16'd54743, 16'd64375, 16'd63465, 16'd18747, 16'd38656, 16'd55531, 16'd62528, 16'd21018, 16'd5467, 16'd45619, 16'd22596, 16'd49317, 16'd25483});
	test_expansion(128'h0279b4b35a45b1290f46e46559307fa2, {16'd8435, 16'd41473, 16'd57442, 16'd31889, 16'd6814, 16'd28367, 16'd20094, 16'd17489, 16'd49555, 16'd40976, 16'd3002, 16'd36535, 16'd35429, 16'd28454, 16'd12135, 16'd54858, 16'd55400, 16'd33618, 16'd63028, 16'd27296, 16'd29026, 16'd13880, 16'd14517, 16'd17252, 16'd51910, 16'd58152});
	test_expansion(128'h9df8f05ecd9e3a2036d6a9971a18cd75, {16'd52079, 16'd45773, 16'd26, 16'd1422, 16'd51200, 16'd56965, 16'd28014, 16'd34464, 16'd564, 16'd42032, 16'd60583, 16'd18306, 16'd61044, 16'd32850, 16'd12916, 16'd29928, 16'd40747, 16'd48360, 16'd62208, 16'd11966, 16'd14090, 16'd41672, 16'd59897, 16'd38056, 16'd62076, 16'd31926});
	test_expansion(128'he57e3ce38dc9d026c92f619585c4fd9f, {16'd54009, 16'd23061, 16'd30145, 16'd61723, 16'd7920, 16'd16439, 16'd23074, 16'd11867, 16'd4933, 16'd4761, 16'd28995, 16'd31722, 16'd43882, 16'd5603, 16'd6508, 16'd48731, 16'd30583, 16'd51960, 16'd40051, 16'd25451, 16'd55032, 16'd64245, 16'd12667, 16'd55417, 16'd4520, 16'd3781});
	test_expansion(128'h8a952a8a5b2161e4f9c38b3ec5c4729e, {16'd56313, 16'd21542, 16'd47315, 16'd24558, 16'd57691, 16'd48119, 16'd8166, 16'd45826, 16'd46360, 16'd20511, 16'd44322, 16'd6303, 16'd50080, 16'd31630, 16'd8663, 16'd54986, 16'd34529, 16'd55718, 16'd19466, 16'd64819, 16'd28708, 16'd37504, 16'd12464, 16'd62874, 16'd64253, 16'd41578});
	test_expansion(128'h033fa4edda099e0f1a833423a957a869, {16'd23400, 16'd45098, 16'd51292, 16'd16576, 16'd63924, 16'd54651, 16'd21404, 16'd46215, 16'd64975, 16'd30680, 16'd20854, 16'd33537, 16'd39748, 16'd17269, 16'd29070, 16'd9613, 16'd6805, 16'd62717, 16'd5143, 16'd42598, 16'd50327, 16'd5168, 16'd24042, 16'd48239, 16'd14028, 16'd24054});
	test_expansion(128'h280e9785f3640241743acb0284a987d8, {16'd35062, 16'd38918, 16'd64899, 16'd30977, 16'd53404, 16'd12425, 16'd33599, 16'd44277, 16'd6984, 16'd23680, 16'd26682, 16'd10055, 16'd7733, 16'd2895, 16'd17719, 16'd22425, 16'd9721, 16'd42803, 16'd50205, 16'd21649, 16'd34472, 16'd51212, 16'd25398, 16'd18112, 16'd2908, 16'd40654});
	test_expansion(128'h542686241b01ae4be1499ec8e5eee43b, {16'd21586, 16'd51257, 16'd42951, 16'd41053, 16'd54052, 16'd6073, 16'd28311, 16'd46065, 16'd8949, 16'd24455, 16'd58893, 16'd35567, 16'd25571, 16'd55883, 16'd33723, 16'd10450, 16'd31795, 16'd22748, 16'd58111, 16'd25268, 16'd25323, 16'd45153, 16'd16906, 16'd45724, 16'd23113, 16'd28527});
	test_expansion(128'h7abd6dcefea3336573ccf860e75b483c, {16'd61195, 16'd7933, 16'd2014, 16'd52174, 16'd16117, 16'd16468, 16'd54537, 16'd62441, 16'd51654, 16'd21131, 16'd22428, 16'd26312, 16'd55629, 16'd26189, 16'd13896, 16'd38273, 16'd28835, 16'd27461, 16'd3059, 16'd27026, 16'd16588, 16'd27796, 16'd39924, 16'd20122, 16'd6390, 16'd26945});
	test_expansion(128'hedebf78e4836cd9def3ab96f4e9e2313, {16'd57966, 16'd31920, 16'd33670, 16'd4744, 16'd58533, 16'd50198, 16'd29992, 16'd35923, 16'd2760, 16'd23859, 16'd49004, 16'd18883, 16'd35560, 16'd38403, 16'd28340, 16'd10069, 16'd39969, 16'd13182, 16'd26358, 16'd1148, 16'd3613, 16'd130, 16'd48814, 16'd50416, 16'd11640, 16'd14498});
	test_expansion(128'h4d7bdd0b9458f348ad53f27604028257, {16'd51471, 16'd15219, 16'd25999, 16'd46034, 16'd25620, 16'd48057, 16'd34548, 16'd21849, 16'd22963, 16'd25530, 16'd14010, 16'd9531, 16'd35734, 16'd50038, 16'd37096, 16'd50595, 16'd55648, 16'd54700, 16'd13851, 16'd65324, 16'd19120, 16'd56101, 16'd13383, 16'd37579, 16'd15569, 16'd15211});
	test_expansion(128'h0ac3d183189ca0fabeaf94c2a72ebe55, {16'd11706, 16'd39046, 16'd13798, 16'd54855, 16'd11274, 16'd50552, 16'd30325, 16'd34719, 16'd48877, 16'd24722, 16'd10103, 16'd52637, 16'd64479, 16'd62524, 16'd980, 16'd44489, 16'd36308, 16'd58184, 16'd8966, 16'd27516, 16'd27472, 16'd14004, 16'd40547, 16'd20766, 16'd43812, 16'd13278});
	test_expansion(128'h0ab2e5fb0925fdd431e480f46681324a, {16'd60593, 16'd27006, 16'd31830, 16'd9300, 16'd58683, 16'd24709, 16'd60688, 16'd22393, 16'd25802, 16'd63004, 16'd9722, 16'd34091, 16'd62756, 16'd5568, 16'd22815, 16'd54746, 16'd39053, 16'd8443, 16'd33542, 16'd848, 16'd42337, 16'd36965, 16'd49878, 16'd9400, 16'd14358, 16'd4366});
	test_expansion(128'h9dce575dc5c9d957ca54e1bdfe690f41, {16'd60149, 16'd61197, 16'd14681, 16'd47435, 16'd64353, 16'd57935, 16'd42464, 16'd56947, 16'd22856, 16'd8357, 16'd61611, 16'd13667, 16'd65286, 16'd29914, 16'd1214, 16'd28691, 16'd52052, 16'd31484, 16'd63173, 16'd63601, 16'd1031, 16'd37942, 16'd26494, 16'd42928, 16'd29402, 16'd38536});
	test_expansion(128'h803404b9cedf5882ed38df024289ec2a, {16'd53562, 16'd52771, 16'd16734, 16'd63518, 16'd17384, 16'd61313, 16'd51724, 16'd36557, 16'd22935, 16'd8512, 16'd10379, 16'd40076, 16'd37631, 16'd42246, 16'd50490, 16'd42820, 16'd62432, 16'd28439, 16'd763, 16'd23553, 16'd64222, 16'd57282, 16'd19746, 16'd32877, 16'd33315, 16'd58530});
	test_expansion(128'h0558f51fff00e09e4a08ebad06bf3ccc, {16'd49966, 16'd4949, 16'd28857, 16'd26190, 16'd57022, 16'd6276, 16'd23398, 16'd64072, 16'd43253, 16'd21579, 16'd63577, 16'd31468, 16'd43700, 16'd52081, 16'd23859, 16'd18387, 16'd42329, 16'd18051, 16'd8352, 16'd22671, 16'd35137, 16'd15889, 16'd64782, 16'd33509, 16'd62135, 16'd19120});
	test_expansion(128'hc22cdb1dbe1dc1aa2304b317e0934653, {16'd32685, 16'd40450, 16'd13006, 16'd17097, 16'd15996, 16'd59630, 16'd50640, 16'd197, 16'd47034, 16'd64565, 16'd34379, 16'd31749, 16'd36047, 16'd13292, 16'd5827, 16'd38187, 16'd1343, 16'd48733, 16'd29355, 16'd55223, 16'd2335, 16'd2297, 16'd35989, 16'd65010, 16'd53686, 16'd18567});
	test_expansion(128'h497ef8c7621808d49ded0ba475b2252d, {16'd46171, 16'd46207, 16'd37475, 16'd64089, 16'd56332, 16'd11586, 16'd5622, 16'd48097, 16'd57139, 16'd58677, 16'd9825, 16'd13942, 16'd15487, 16'd35257, 16'd6562, 16'd49286, 16'd42020, 16'd34946, 16'd41046, 16'd50937, 16'd61730, 16'd53058, 16'd61339, 16'd16044, 16'd32569, 16'd35519});
	test_expansion(128'he08368847c5107a44341a834fa22abaa, {16'd26738, 16'd62443, 16'd50152, 16'd43425, 16'd42554, 16'd51788, 16'd23254, 16'd22267, 16'd5347, 16'd519, 16'd16654, 16'd43708, 16'd39003, 16'd16378, 16'd56613, 16'd40538, 16'd30177, 16'd36257, 16'd21252, 16'd31807, 16'd44762, 16'd32988, 16'd38494, 16'd22289, 16'd40480, 16'd58601});
	test_expansion(128'hcca540c570c5cc7522ee576bf35dc335, {16'd33177, 16'd41263, 16'd18065, 16'd38798, 16'd26239, 16'd50408, 16'd20503, 16'd21034, 16'd63647, 16'd40956, 16'd55827, 16'd42749, 16'd6074, 16'd34829, 16'd45695, 16'd56824, 16'd23695, 16'd33948, 16'd23767, 16'd7092, 16'd37137, 16'd33230, 16'd41099, 16'd63999, 16'd59020, 16'd32717});
	test_expansion(128'h2839bab6c9d077163b6455b8b1f2ba43, {16'd21938, 16'd1271, 16'd41434, 16'd49564, 16'd15592, 16'd65284, 16'd44920, 16'd20037, 16'd54922, 16'd36167, 16'd37070, 16'd41107, 16'd29519, 16'd19051, 16'd25512, 16'd31862, 16'd15314, 16'd11033, 16'd36742, 16'd31490, 16'd6015, 16'd5172, 16'd60364, 16'd10145, 16'd16290, 16'd29006});
	test_expansion(128'h4fc95d7a82532ca2d7d67c47fae60855, {16'd47839, 16'd58480, 16'd16453, 16'd12797, 16'd15279, 16'd27565, 16'd8746, 16'd46785, 16'd13703, 16'd9455, 16'd50869, 16'd29876, 16'd53239, 16'd43259, 16'd60451, 16'd42606, 16'd19874, 16'd11809, 16'd64632, 16'd46730, 16'd61015, 16'd9158, 16'd14404, 16'd14398, 16'd40940, 16'd27801});
	test_expansion(128'hdba23519655d999249a388eed81b8178, {16'd26587, 16'd28468, 16'd7290, 16'd35375, 16'd17715, 16'd13588, 16'd53657, 16'd23155, 16'd26786, 16'd61134, 16'd63563, 16'd27585, 16'd2816, 16'd54672, 16'd37886, 16'd27428, 16'd19929, 16'd26071, 16'd38521, 16'd38805, 16'd60400, 16'd5249, 16'd64508, 16'd14222, 16'd60502, 16'd49679});
	test_expansion(128'h163efe111e1678156fda446b466c1a02, {16'd25987, 16'd59668, 16'd45476, 16'd57846, 16'd42124, 16'd16331, 16'd18851, 16'd7962, 16'd15655, 16'd5429, 16'd47018, 16'd24870, 16'd38480, 16'd21876, 16'd51269, 16'd17328, 16'd21487, 16'd31472, 16'd41058, 16'd57958, 16'd28204, 16'd43460, 16'd36958, 16'd25947, 16'd61055, 16'd48582});
	test_expansion(128'hfb0e919cab8d59da6ae3151a5175b533, {16'd55074, 16'd49997, 16'd53625, 16'd12307, 16'd52605, 16'd44903, 16'd28464, 16'd48349, 16'd8214, 16'd39053, 16'd16019, 16'd37178, 16'd3453, 16'd6895, 16'd43671, 16'd29840, 16'd5447, 16'd6839, 16'd11481, 16'd37182, 16'd21884, 16'd38128, 16'd5044, 16'd35612, 16'd8304, 16'd41463});
	test_expansion(128'hf15228a76d5fb876bb164ffb6516d72e, {16'd13825, 16'd52468, 16'd42137, 16'd63089, 16'd17492, 16'd65472, 16'd43799, 16'd60291, 16'd33593, 16'd21704, 16'd6325, 16'd55881, 16'd52227, 16'd28142, 16'd47030, 16'd12172, 16'd4958, 16'd44043, 16'd27383, 16'd49241, 16'd4883, 16'd64096, 16'd14268, 16'd53300, 16'd42994, 16'd24537});
	test_expansion(128'h8f3750d58ba6a723f2edad625651af76, {16'd25647, 16'd18896, 16'd15077, 16'd32975, 16'd26, 16'd40994, 16'd22420, 16'd28111, 16'd43942, 16'd28936, 16'd64002, 16'd64839, 16'd43503, 16'd48261, 16'd17973, 16'd32582, 16'd27652, 16'd12417, 16'd10867, 16'd19791, 16'd4723, 16'd21552, 16'd6355, 16'd44515, 16'd47261, 16'd56276});
	test_expansion(128'h697edf5c551b6ea82f6958a724ccec2d, {16'd28732, 16'd25386, 16'd40487, 16'd36990, 16'd42313, 16'd24959, 16'd56736, 16'd47044, 16'd23637, 16'd61742, 16'd53279, 16'd15494, 16'd53757, 16'd41333, 16'd322, 16'd45553, 16'd41932, 16'd51704, 16'd5655, 16'd11855, 16'd38944, 16'd6951, 16'd6083, 16'd36416, 16'd49712, 16'd14383});
	test_expansion(128'h84440384fcaf5d76b71a75cdbcfa9e93, {16'd24042, 16'd21717, 16'd62649, 16'd53182, 16'd8211, 16'd6971, 16'd60702, 16'd62518, 16'd44799, 16'd45184, 16'd47644, 16'd38695, 16'd25272, 16'd28835, 16'd18273, 16'd7302, 16'd35355, 16'd58688, 16'd14494, 16'd51462, 16'd1358, 16'd33722, 16'd5417, 16'd62632, 16'd45737, 16'd63856});
	test_expansion(128'h813b6e790fe91d017d7a8ab593a273b0, {16'd11315, 16'd33457, 16'd65124, 16'd12023, 16'd30714, 16'd19098, 16'd15667, 16'd17961, 16'd1221, 16'd42579, 16'd42653, 16'd22887, 16'd64947, 16'd22770, 16'd47230, 16'd25907, 16'd30590, 16'd22330, 16'd2952, 16'd15827, 16'd8356, 16'd61222, 16'd45504, 16'd51333, 16'd16061, 16'd59093});
	test_expansion(128'hd84eaf97b393981aee54676d5213ad01, {16'd19161, 16'd39212, 16'd17143, 16'd35256, 16'd7765, 16'd50269, 16'd35638, 16'd48353, 16'd30610, 16'd19467, 16'd55311, 16'd47627, 16'd7324, 16'd33403, 16'd27044, 16'd14938, 16'd33201, 16'd59385, 16'd46880, 16'd54873, 16'd41014, 16'd4592, 16'd30174, 16'd46884, 16'd47539, 16'd16920});
	test_expansion(128'hdfdf0e0d63e350999c7fb02acbc8f298, {16'd40345, 16'd25125, 16'd16581, 16'd20358, 16'd50750, 16'd10391, 16'd51424, 16'd14684, 16'd53188, 16'd44509, 16'd22731, 16'd45116, 16'd40681, 16'd24300, 16'd59412, 16'd10069, 16'd1574, 16'd10966, 16'd13983, 16'd11098, 16'd2488, 16'd12830, 16'd27976, 16'd49392, 16'd45202, 16'd54407});
	test_expansion(128'h969f04d84fbeb91fe2f810052a40d9c7, {16'd44572, 16'd48965, 16'd14996, 16'd16805, 16'd39374, 16'd31455, 16'd19523, 16'd4480, 16'd20383, 16'd29672, 16'd43751, 16'd38086, 16'd15502, 16'd57454, 16'd54429, 16'd24629, 16'd24117, 16'd27460, 16'd33354, 16'd63663, 16'd30556, 16'd27266, 16'd9427, 16'd63479, 16'd21005, 16'd57373});
	test_expansion(128'ha154c2568059b8b94a8d681bf57617fc, {16'd54118, 16'd10509, 16'd29507, 16'd2707, 16'd29389, 16'd39344, 16'd52376, 16'd44517, 16'd2731, 16'd7932, 16'd17696, 16'd13736, 16'd51263, 16'd51648, 16'd59995, 16'd35285, 16'd20519, 16'd3153, 16'd38221, 16'd54873, 16'd23633, 16'd57393, 16'd53819, 16'd27346, 16'd5048, 16'd12776});
	test_expansion(128'h73bffcd7061c2d0a6fdddeae1b67690a, {16'd40260, 16'd10906, 16'd41832, 16'd12353, 16'd9621, 16'd28638, 16'd41011, 16'd48565, 16'd45521, 16'd3243, 16'd8497, 16'd35357, 16'd23613, 16'd25264, 16'd64169, 16'd16716, 16'd37968, 16'd17908, 16'd40148, 16'd64051, 16'd44371, 16'd32450, 16'd16091, 16'd13774, 16'd19999, 16'd20994});
	test_expansion(128'h38d96f900d48ba53c7edaf91ace46420, {16'd2877, 16'd18510, 16'd6947, 16'd46531, 16'd42134, 16'd3119, 16'd46906, 16'd15302, 16'd22316, 16'd35073, 16'd13523, 16'd8824, 16'd47392, 16'd21647, 16'd20275, 16'd24790, 16'd32267, 16'd36594, 16'd25830, 16'd20949, 16'd46820, 16'd15193, 16'd34167, 16'd17927, 16'd15031, 16'd39385});
	test_expansion(128'hb6b6a253f54ef7ec0129f4211cf8705a, {16'd34549, 16'd53250, 16'd63929, 16'd49626, 16'd1123, 16'd26920, 16'd11889, 16'd45644, 16'd3016, 16'd59985, 16'd25089, 16'd25708, 16'd6252, 16'd10476, 16'd55176, 16'd16374, 16'd61362, 16'd45293, 16'd34831, 16'd64022, 16'd25126, 16'd42029, 16'd10730, 16'd30505, 16'd4028, 16'd26288});
	test_expansion(128'hf347a94452e71628c38fd85bc2c0c813, {16'd22844, 16'd8561, 16'd59883, 16'd39097, 16'd26497, 16'd6338, 16'd47194, 16'd45134, 16'd29655, 16'd43341, 16'd17217, 16'd50269, 16'd30716, 16'd19369, 16'd12735, 16'd44284, 16'd15359, 16'd12112, 16'd15550, 16'd55673, 16'd53768, 16'd47009, 16'd28182, 16'd50193, 16'd33317, 16'd64944});
	test_expansion(128'h31a15c7bfe399fbdfc82a1b81cbb7a94, {16'd61156, 16'd44081, 16'd3568, 16'd41471, 16'd51482, 16'd56897, 16'd51661, 16'd35759, 16'd59623, 16'd55668, 16'd39146, 16'd58916, 16'd60296, 16'd17446, 16'd22956, 16'd1064, 16'd36909, 16'd45437, 16'd14551, 16'd18398, 16'd16046, 16'd50406, 16'd49100, 16'd39284, 16'd51434, 16'd62763});
	test_expansion(128'hdad4278c4f3aa88b4b070250ef7f1c04, {16'd29374, 16'd31204, 16'd61152, 16'd10008, 16'd35772, 16'd61917, 16'd13455, 16'd12442, 16'd53019, 16'd25073, 16'd47763, 16'd22704, 16'd48525, 16'd53145, 16'd46997, 16'd63273, 16'd28474, 16'd53052, 16'd54595, 16'd45846, 16'd1418, 16'd49210, 16'd6695, 16'd11138, 16'd33445, 16'd19977});
	test_expansion(128'h7e1549323d34c563c7b35bba615d5fd0, {16'd49869, 16'd61568, 16'd43499, 16'd21327, 16'd24410, 16'd64411, 16'd62122, 16'd4861, 16'd25341, 16'd58163, 16'd51765, 16'd8893, 16'd2799, 16'd3536, 16'd16718, 16'd16797, 16'd29335, 16'd63855, 16'd2926, 16'd58877, 16'd23129, 16'd21532, 16'd6908, 16'd312, 16'd45389, 16'd65430});
	test_expansion(128'h9791f88f5801adeb2388e9d285d10718, {16'd28869, 16'd14437, 16'd47849, 16'd55912, 16'd38224, 16'd24964, 16'd62088, 16'd48858, 16'd50542, 16'd36578, 16'd50886, 16'd998, 16'd27361, 16'd63388, 16'd32753, 16'd62485, 16'd364, 16'd40314, 16'd27868, 16'd23650, 16'd49866, 16'd3328, 16'd42394, 16'd47696, 16'd2264, 16'd64848});
	test_expansion(128'h9c3089783691163dff0df7cb2bda229c, {16'd31162, 16'd59870, 16'd23173, 16'd61595, 16'd56558, 16'd10900, 16'd29266, 16'd52181, 16'd47594, 16'd19887, 16'd12265, 16'd14345, 16'd24196, 16'd48928, 16'd51901, 16'd15837, 16'd38704, 16'd32782, 16'd20566, 16'd27376, 16'd47489, 16'd59973, 16'd12411, 16'd26355, 16'd48938, 16'd2139});
	test_expansion(128'h246d0cd76151d2fcda19012b270240e5, {16'd28318, 16'd30953, 16'd3699, 16'd57133, 16'd10359, 16'd12036, 16'd63699, 16'd62742, 16'd52573, 16'd52162, 16'd57064, 16'd17328, 16'd42957, 16'd36072, 16'd51558, 16'd59981, 16'd30539, 16'd43875, 16'd12892, 16'd55238, 16'd55182, 16'd55500, 16'd13402, 16'd47390, 16'd20098, 16'd50419});
	test_expansion(128'h3106fdb6c8be3a2580920d06a1c82b2b, {16'd2667, 16'd12433, 16'd53084, 16'd62620, 16'd7346, 16'd44334, 16'd13624, 16'd21497, 16'd16900, 16'd11115, 16'd39490, 16'd2043, 16'd19183, 16'd14636, 16'd21093, 16'd5704, 16'd25492, 16'd14635, 16'd45127, 16'd40341, 16'd51304, 16'd21414, 16'd17355, 16'd44792, 16'd6114, 16'd45391});
	test_expansion(128'ha2dc2870a752f0d41f7b61294700f1de, {16'd62838, 16'd31674, 16'd55119, 16'd6369, 16'd27005, 16'd5074, 16'd2374, 16'd62396, 16'd47347, 16'd59678, 16'd43142, 16'd13540, 16'd25709, 16'd51071, 16'd47009, 16'd40257, 16'd28723, 16'd11, 16'd14568, 16'd46228, 16'd41187, 16'd11310, 16'd31991, 16'd31857, 16'd57406, 16'd1064});
	test_expansion(128'he10d8efc689d7b1c17e8ebd8dc941507, {16'd20571, 16'd55692, 16'd20264, 16'd58537, 16'd64531, 16'd43178, 16'd50157, 16'd5272, 16'd5826, 16'd44670, 16'd13753, 16'd60305, 16'd25950, 16'd55621, 16'd33574, 16'd62701, 16'd18199, 16'd12661, 16'd52569, 16'd46270, 16'd31284, 16'd7620, 16'd34355, 16'd2149, 16'd18166, 16'd6675});
	test_expansion(128'h217ad3957302385290df1a0d590065de, {16'd3105, 16'd22129, 16'd45005, 16'd36313, 16'd18099, 16'd31845, 16'd17628, 16'd12859, 16'd46847, 16'd20665, 16'd47399, 16'd42835, 16'd36018, 16'd11291, 16'd55999, 16'd33214, 16'd63408, 16'd18896, 16'd32221, 16'd17062, 16'd65271, 16'd33908, 16'd60496, 16'd1035, 16'd22888, 16'd31203});
	test_expansion(128'h34e75cc8b6ab0e114ad4d8375c31ecf7, {16'd4800, 16'd51238, 16'd61035, 16'd6398, 16'd26095, 16'd39112, 16'd51836, 16'd2053, 16'd29958, 16'd35344, 16'd42048, 16'd1287, 16'd48631, 16'd9388, 16'd29837, 16'd36375, 16'd47489, 16'd15612, 16'd17395, 16'd60260, 16'd3776, 16'd58385, 16'd17606, 16'd10636, 16'd65287, 16'd3562});
	test_expansion(128'hb31791224d5fc9944bb680abeda77bc5, {16'd56565, 16'd47064, 16'd65322, 16'd55333, 16'd25364, 16'd54505, 16'd22317, 16'd4846, 16'd43560, 16'd51205, 16'd38583, 16'd6839, 16'd7823, 16'd4365, 16'd33283, 16'd24854, 16'd44962, 16'd18890, 16'd14033, 16'd30025, 16'd28800, 16'd2726, 16'd36798, 16'd39999, 16'd58711, 16'd19607});
	test_expansion(128'hcaf978a4ab9c5957dd340aa986fcb209, {16'd41827, 16'd57992, 16'd7048, 16'd46626, 16'd101, 16'd38306, 16'd36217, 16'd6986, 16'd37818, 16'd21616, 16'd38606, 16'd53124, 16'd1528, 16'd31195, 16'd4596, 16'd23689, 16'd11344, 16'd44569, 16'd19088, 16'd19465, 16'd10857, 16'd19816, 16'd62951, 16'd51095, 16'd64031, 16'd56228});
	test_expansion(128'h7c501699dd1d0873eb471d9d8cbc1640, {16'd26471, 16'd59472, 16'd19189, 16'd17319, 16'd38, 16'd53006, 16'd16638, 16'd11891, 16'd41144, 16'd58741, 16'd54907, 16'd34338, 16'd45212, 16'd60520, 16'd46099, 16'd44436, 16'd1026, 16'd31072, 16'd17446, 16'd59440, 16'd13930, 16'd20804, 16'd29375, 16'd2230, 16'd13061, 16'd40242});
	test_expansion(128'h3b39bd8c4575cda69d4fd7de4d947cb5, {16'd28999, 16'd4734, 16'd62983, 16'd33315, 16'd11652, 16'd11727, 16'd13047, 16'd17573, 16'd42750, 16'd29212, 16'd3889, 16'd9938, 16'd20910, 16'd62185, 16'd40259, 16'd46740, 16'd17882, 16'd38283, 16'd47196, 16'd5901, 16'd13573, 16'd50788, 16'd60994, 16'd34428, 16'd56719, 16'd53621});
	test_expansion(128'h040aa3125b585d5730d7448a3590739d, {16'd8934, 16'd14675, 16'd10316, 16'd1556, 16'd42203, 16'd63849, 16'd48546, 16'd49701, 16'd28948, 16'd27326, 16'd35915, 16'd44887, 16'd7090, 16'd32247, 16'd57040, 16'd38123, 16'd42435, 16'd20231, 16'd58247, 16'd43826, 16'd14124, 16'd2795, 16'd28236, 16'd41609, 16'd9323, 16'd60078});
	test_expansion(128'hb9ec991823b83cd64f0abef140c0c56d, {16'd31261, 16'd26743, 16'd30558, 16'd40090, 16'd47636, 16'd37588, 16'd33416, 16'd51434, 16'd45612, 16'd23233, 16'd31070, 16'd48661, 16'd58486, 16'd4542, 16'd56286, 16'd950, 16'd38694, 16'd53015, 16'd7275, 16'd13229, 16'd40611, 16'd25780, 16'd42800, 16'd44078, 16'd60481, 16'd22646});
	test_expansion(128'h67eaf29c3da62c3de546e87d80137b81, {16'd48263, 16'd2682, 16'd45030, 16'd58623, 16'd56246, 16'd52034, 16'd47688, 16'd4943, 16'd44354, 16'd31205, 16'd10791, 16'd37861, 16'd30733, 16'd4732, 16'd45981, 16'd3880, 16'd46565, 16'd45144, 16'd30149, 16'd57253, 16'd35230, 16'd32082, 16'd24967, 16'd38052, 16'd36195, 16'd22493});
	test_expansion(128'h749c4cb81721b78d6492aa9ebed01712, {16'd15708, 16'd6297, 16'd26464, 16'd14887, 16'd60738, 16'd61700, 16'd28757, 16'd22387, 16'd22647, 16'd41104, 16'd12115, 16'd46047, 16'd6939, 16'd33058, 16'd25781, 16'd34955, 16'd65293, 16'd31133, 16'd28973, 16'd25121, 16'd6504, 16'd8433, 16'd26761, 16'd114, 16'd48790, 16'd57686});
	test_expansion(128'h0b80faab30149fe8682c8f59ad3de3ae, {16'd4197, 16'd62565, 16'd24609, 16'd28879, 16'd3159, 16'd43506, 16'd41627, 16'd30738, 16'd63746, 16'd38359, 16'd61628, 16'd56818, 16'd23958, 16'd35243, 16'd45195, 16'd40170, 16'd20525, 16'd14295, 16'd7937, 16'd52727, 16'd42199, 16'd27313, 16'd1124, 16'd16435, 16'd48043, 16'd51429});
	test_expansion(128'hb81679f3b002edecd6d2e16fefc00304, {16'd29525, 16'd60143, 16'd1860, 16'd51284, 16'd27047, 16'd24858, 16'd23313, 16'd24038, 16'd9534, 16'd26417, 16'd18854, 16'd11733, 16'd20432, 16'd40980, 16'd32595, 16'd59306, 16'd4876, 16'd61512, 16'd18752, 16'd39296, 16'd60342, 16'd50279, 16'd23362, 16'd33237, 16'd19393, 16'd6903});
	test_expansion(128'hc0da6402e96cc010ff3675e1addd8b94, {16'd13759, 16'd59787, 16'd32203, 16'd60793, 16'd10780, 16'd5227, 16'd26221, 16'd4175, 16'd33868, 16'd54710, 16'd61831, 16'd17987, 16'd62536, 16'd13356, 16'd43410, 16'd64898, 16'd13100, 16'd43844, 16'd56306, 16'd7564, 16'd34070, 16'd3942, 16'd21839, 16'd26080, 16'd25784, 16'd55808});
	test_expansion(128'hb0e8d75ddb60017779b16308bbd6d0e7, {16'd29759, 16'd55616, 16'd1372, 16'd43295, 16'd16628, 16'd60102, 16'd54054, 16'd57408, 16'd61509, 16'd57822, 16'd48805, 16'd59746, 16'd22901, 16'd62577, 16'd35258, 16'd62069, 16'd44394, 16'd2659, 16'd44828, 16'd45847, 16'd44251, 16'd36448, 16'd1451, 16'd31807, 16'd55636, 16'd39147});
	test_expansion(128'ha1aaf41dabec5ebfe93ccb7f2673228e, {16'd33476, 16'd30807, 16'd3786, 16'd22688, 16'd59036, 16'd4553, 16'd49378, 16'd2156, 16'd12643, 16'd96, 16'd26558, 16'd30987, 16'd44862, 16'd7942, 16'd21139, 16'd57618, 16'd57662, 16'd61958, 16'd46690, 16'd19932, 16'd566, 16'd52527, 16'd65489, 16'd20515, 16'd30639, 16'd4326});
	test_expansion(128'h90a01181182adc039fd00fe0818bbd33, {16'd20853, 16'd52164, 16'd15633, 16'd13368, 16'd54246, 16'd46828, 16'd63992, 16'd57026, 16'd60394, 16'd53610, 16'd30618, 16'd42127, 16'd17049, 16'd39054, 16'd8776, 16'd26492, 16'd14916, 16'd29090, 16'd47541, 16'd26563, 16'd19003, 16'd10389, 16'd61910, 16'd44334, 16'd44067, 16'd42274});
	test_expansion(128'h2bc05fff8439e96c9a9e5c4282a3d819, {16'd6628, 16'd40595, 16'd56658, 16'd27915, 16'd33561, 16'd31482, 16'd56087, 16'd36377, 16'd55380, 16'd9860, 16'd26420, 16'd64658, 16'd52617, 16'd17739, 16'd21386, 16'd49552, 16'd12926, 16'd57191, 16'd43228, 16'd26408, 16'd37696, 16'd36720, 16'd29915, 16'd60132, 16'd25193, 16'd52624});
	test_expansion(128'h094af4454d8eb8497c5559b41fe01296, {16'd60027, 16'd16372, 16'd44055, 16'd54907, 16'd34452, 16'd2864, 16'd7756, 16'd11570, 16'd57185, 16'd7365, 16'd4242, 16'd14919, 16'd4047, 16'd29941, 16'd21885, 16'd43216, 16'd59833, 16'd4170, 16'd10878, 16'd40960, 16'd6056, 16'd39296, 16'd9291, 16'd7174, 16'd52738, 16'd16507});
	test_expansion(128'hec890dfa89cd5bc72ea74891c1279c63, {16'd61095, 16'd25476, 16'd1093, 16'd43083, 16'd11333, 16'd48954, 16'd17715, 16'd1776, 16'd37814, 16'd20550, 16'd43177, 16'd60609, 16'd24616, 16'd43810, 16'd64508, 16'd38880, 16'd20400, 16'd45082, 16'd12763, 16'd26807, 16'd5389, 16'd56179, 16'd44031, 16'd27968, 16'd54630, 16'd38860});
	test_expansion(128'h4149cdf9cc0c80a5592662c2a263554d, {16'd21903, 16'd43751, 16'd23433, 16'd5225, 16'd3393, 16'd11651, 16'd44881, 16'd14515, 16'd53896, 16'd4113, 16'd39163, 16'd33805, 16'd57579, 16'd33615, 16'd15962, 16'd49147, 16'd12683, 16'd21911, 16'd14639, 16'd56119, 16'd2335, 16'd37650, 16'd37349, 16'd32864, 16'd15144, 16'd44441});
	test_expansion(128'hf889f2b648c76070037198adde5c6a4f, {16'd31175, 16'd38389, 16'd11459, 16'd62076, 16'd8764, 16'd8174, 16'd40318, 16'd49671, 16'd61904, 16'd35360, 16'd28397, 16'd52244, 16'd42077, 16'd50377, 16'd33983, 16'd37509, 16'd9521, 16'd47008, 16'd25903, 16'd40226, 16'd5792, 16'd60914, 16'd63182, 16'd24967, 16'd41553, 16'd29235});
	test_expansion(128'h1b1f62b1841c44ead98d235bfc02082f, {16'd8755, 16'd23591, 16'd12200, 16'd19665, 16'd10080, 16'd4636, 16'd23814, 16'd51292, 16'd45245, 16'd58825, 16'd62418, 16'd59351, 16'd3438, 16'd41034, 16'd30791, 16'd38636, 16'd5045, 16'd2755, 16'd63551, 16'd4455, 16'd42593, 16'd46781, 16'd13262, 16'd25700, 16'd59805, 16'd53172});
	test_expansion(128'hc3a10b6e9ab1658b267781e1556d2ac1, {16'd14787, 16'd33749, 16'd23304, 16'd27250, 16'd11100, 16'd24663, 16'd7665, 16'd57312, 16'd47242, 16'd20314, 16'd59380, 16'd56243, 16'd29103, 16'd48802, 16'd18144, 16'd21601, 16'd40203, 16'd41829, 16'd26030, 16'd63058, 16'd12051, 16'd51700, 16'd48772, 16'd48675, 16'd3914, 16'd23912});
	test_expansion(128'hba81e9d4296e017953a371f323ee3a94, {16'd48801, 16'd16493, 16'd32940, 16'd10763, 16'd5900, 16'd16509, 16'd34840, 16'd23384, 16'd14459, 16'd21455, 16'd22869, 16'd43215, 16'd52966, 16'd55714, 16'd20137, 16'd63229, 16'd7474, 16'd14598, 16'd43023, 16'd48187, 16'd51206, 16'd56650, 16'd26110, 16'd54941, 16'd38266, 16'd28409});
	test_expansion(128'hc300b0003b5f3e48ccd2ba9a96561319, {16'd2608, 16'd4532, 16'd42916, 16'd26798, 16'd21449, 16'd36913, 16'd63264, 16'd51184, 16'd48322, 16'd12010, 16'd41525, 16'd33175, 16'd30321, 16'd64550, 16'd16193, 16'd53504, 16'd32369, 16'd63344, 16'd38762, 16'd12038, 16'd35684, 16'd60334, 16'd30841, 16'd43468, 16'd28271, 16'd37024});
	test_expansion(128'h632eddf48f17a75d26c22b663e851df6, {16'd9410, 16'd11034, 16'd65293, 16'd64114, 16'd51434, 16'd15626, 16'd58469, 16'd46593, 16'd21631, 16'd65507, 16'd40676, 16'd34285, 16'd49733, 16'd53592, 16'd32440, 16'd50569, 16'd44632, 16'd36410, 16'd47345, 16'd32423, 16'd63331, 16'd38918, 16'd28860, 16'd37207, 16'd1608, 16'd1822});
	test_expansion(128'h332b028b095d8a7b0796efdb2b8bd5c4, {16'd50840, 16'd59662, 16'd32533, 16'd32188, 16'd60715, 16'd5804, 16'd2273, 16'd8933, 16'd9351, 16'd13610, 16'd13183, 16'd15757, 16'd50096, 16'd13031, 16'd59621, 16'd8721, 16'd11151, 16'd51933, 16'd12511, 16'd47809, 16'd25650, 16'd64871, 16'd34992, 16'd54835, 16'd9554, 16'd32304});
	test_expansion(128'h0737a5ac82705137c77f24faf8f49833, {16'd25614, 16'd16036, 16'd27179, 16'd63761, 16'd40881, 16'd43611, 16'd27182, 16'd44129, 16'd12366, 16'd36820, 16'd35012, 16'd9619, 16'd29841, 16'd35922, 16'd5284, 16'd33619, 16'd17137, 16'd49211, 16'd28735, 16'd44023, 16'd470, 16'd11524, 16'd26348, 16'd13755, 16'd9554, 16'd15303});
	test_expansion(128'h0f85042affe4eb5ff6e41179455dde33, {16'd15090, 16'd36138, 16'd29677, 16'd53022, 16'd23876, 16'd29220, 16'd49583, 16'd42922, 16'd53865, 16'd57298, 16'd50174, 16'd49715, 16'd14861, 16'd30260, 16'd9591, 16'd2187, 16'd41289, 16'd15685, 16'd44117, 16'd9937, 16'd32255, 16'd46830, 16'd55124, 16'd14207, 16'd11138, 16'd48258});
	test_expansion(128'hf471aa02acd2d13a0f5e1104e9e84b54, {16'd4742, 16'd29915, 16'd18484, 16'd9046, 16'd15221, 16'd62895, 16'd49849, 16'd43038, 16'd19611, 16'd31062, 16'd1359, 16'd20809, 16'd29208, 16'd60852, 16'd46944, 16'd54906, 16'd47509, 16'd17397, 16'd29507, 16'd25090, 16'd39946, 16'd35789, 16'd61839, 16'd17072, 16'd40177, 16'd30654});
	test_expansion(128'h2cf1fc76c75a787db8bbda576eb6d9c9, {16'd50238, 16'd20494, 16'd12415, 16'd62715, 16'd19175, 16'd42720, 16'd18540, 16'd14811, 16'd50772, 16'd686, 16'd51656, 16'd31416, 16'd29043, 16'd56373, 16'd62747, 16'd39478, 16'd28210, 16'd40729, 16'd35085, 16'd20979, 16'd12300, 16'd4355, 16'd17958, 16'd39420, 16'd56759, 16'd13097});
	test_expansion(128'hbc91e986776b0a28c3a3106fefd7db62, {16'd21431, 16'd4317, 16'd45386, 16'd13930, 16'd8281, 16'd28803, 16'd41609, 16'd65279, 16'd46222, 16'd31876, 16'd47846, 16'd18582, 16'd27479, 16'd54508, 16'd51189, 16'd35467, 16'd18632, 16'd23946, 16'd6887, 16'd54093, 16'd64950, 16'd5328, 16'd4972, 16'd28583, 16'd48138, 16'd36780});
	test_expansion(128'h4414ec7bc8a93a3af3dcf8606cd2689d, {16'd62422, 16'd63174, 16'd34816, 16'd2949, 16'd29882, 16'd65381, 16'd65163, 16'd26285, 16'd14816, 16'd11351, 16'd60818, 16'd4341, 16'd42522, 16'd31108, 16'd56061, 16'd5754, 16'd34289, 16'd58074, 16'd9916, 16'd39265, 16'd522, 16'd12672, 16'd22026, 16'd14406, 16'd38737, 16'd45778});
	test_expansion(128'h57d447913d18c5ae1ba017eaa0a1274d, {16'd45962, 16'd44473, 16'd25252, 16'd45826, 16'd44573, 16'd21670, 16'd35873, 16'd45309, 16'd22920, 16'd2608, 16'd41519, 16'd1735, 16'd58198, 16'd22781, 16'd44269, 16'd26951, 16'd16402, 16'd56312, 16'd183, 16'd31444, 16'd35550, 16'd4362, 16'd17290, 16'd20830, 16'd55804, 16'd40037});
	test_expansion(128'h26de326cf16486570d05ade3c8b2ed5a, {16'd63054, 16'd31008, 16'd33443, 16'd40717, 16'd9302, 16'd16092, 16'd24534, 16'd18558, 16'd28257, 16'd20966, 16'd56709, 16'd45072, 16'd52779, 16'd58728, 16'd34347, 16'd60931, 16'd22603, 16'd3730, 16'd46202, 16'd27255, 16'd14728, 16'd46607, 16'd53589, 16'd54157, 16'd6158, 16'd40175});
	test_expansion(128'hb8bd437518b5b9a33507bc799743f21c, {16'd27286, 16'd14848, 16'd13552, 16'd19056, 16'd4135, 16'd55088, 16'd59548, 16'd24018, 16'd63346, 16'd37722, 16'd27920, 16'd38234, 16'd56757, 16'd59936, 16'd42636, 16'd52198, 16'd5932, 16'd8080, 16'd11321, 16'd29771, 16'd50968, 16'd54030, 16'd34889, 16'd26834, 16'd20529, 16'd45024});
	test_expansion(128'h4c9e8754adf294d719f7bf93c0c9540c, {16'd6079, 16'd26638, 16'd34966, 16'd42941, 16'd38180, 16'd50415, 16'd42211, 16'd38817, 16'd16152, 16'd53627, 16'd30458, 16'd4202, 16'd36909, 16'd13850, 16'd3393, 16'd47005, 16'd64596, 16'd46638, 16'd49453, 16'd10878, 16'd49066, 16'd1869, 16'd52555, 16'd16637, 16'd44287, 16'd20345});
	test_expansion(128'hc99e4bbe55f07f20d1020586eea3381a, {16'd42475, 16'd39606, 16'd32848, 16'd235, 16'd60561, 16'd23640, 16'd26095, 16'd15022, 16'd17812, 16'd9110, 16'd8017, 16'd53536, 16'd4427, 16'd634, 16'd2649, 16'd59150, 16'd44706, 16'd43766, 16'd35271, 16'd21189, 16'd29825, 16'd62175, 16'd454, 16'd5339, 16'd5293, 16'd59579});
	test_expansion(128'hc21ff8aa1bec6b881d55a93d6a66324f, {16'd62280, 16'd20141, 16'd1060, 16'd6195, 16'd8725, 16'd61312, 16'd22189, 16'd24323, 16'd51634, 16'd48481, 16'd41816, 16'd25303, 16'd6977, 16'd47165, 16'd61578, 16'd62939, 16'd47248, 16'd11813, 16'd43485, 16'd13341, 16'd56879, 16'd61142, 16'd37249, 16'd31117, 16'd14121, 16'd8023});
	test_expansion(128'h5f0388680d1e7650321a265b8baca78d, {16'd34664, 16'd13511, 16'd12834, 16'd12640, 16'd47095, 16'd49984, 16'd60966, 16'd1639, 16'd38934, 16'd31433, 16'd54558, 16'd27359, 16'd54311, 16'd49291, 16'd31263, 16'd48552, 16'd34639, 16'd51617, 16'd60164, 16'd43428, 16'd30816, 16'd33319, 16'd33644, 16'd2801, 16'd15038, 16'd53499});
	test_expansion(128'h2941d6488f9f2abd72fc88f74eac1215, {16'd4248, 16'd32804, 16'd11654, 16'd22963, 16'd30127, 16'd28418, 16'd29130, 16'd25132, 16'd8014, 16'd5888, 16'd35404, 16'd58767, 16'd26000, 16'd57572, 16'd55666, 16'd15512, 16'd57215, 16'd4893, 16'd57541, 16'd361, 16'd46073, 16'd64721, 16'd33013, 16'd43373, 16'd806, 16'd26514});
	test_expansion(128'h0e38227b3434395d80682d149e399499, {16'd3004, 16'd29245, 16'd53090, 16'd41147, 16'd1927, 16'd7350, 16'd18338, 16'd42196, 16'd61184, 16'd57053, 16'd59508, 16'd39147, 16'd56380, 16'd22579, 16'd56716, 16'd26144, 16'd64068, 16'd33927, 16'd8537, 16'd20422, 16'd6082, 16'd34484, 16'd17503, 16'd18443, 16'd1255, 16'd63866});
	test_expansion(128'h979cb1e9e1ea1d635508d2ad6217e1ef, {16'd59843, 16'd2304, 16'd37635, 16'd10595, 16'd35557, 16'd1955, 16'd12981, 16'd56272, 16'd21190, 16'd8878, 16'd16736, 16'd29614, 16'd47402, 16'd58566, 16'd45896, 16'd63744, 16'd25437, 16'd56941, 16'd16793, 16'd39515, 16'd65050, 16'd48944, 16'd5392, 16'd8101, 16'd56220, 16'd2231});
	test_expansion(128'hb8825116ee7936f695516835366e8622, {16'd47061, 16'd13405, 16'd54722, 16'd51134, 16'd17074, 16'd2361, 16'd28739, 16'd15192, 16'd30285, 16'd4041, 16'd45452, 16'd36366, 16'd49952, 16'd44056, 16'd39174, 16'd60452, 16'd39748, 16'd60899, 16'd50458, 16'd51045, 16'd29105, 16'd15244, 16'd783, 16'd15999, 16'd57603, 16'd38628});
	test_expansion(128'h8f3066224bdbed3946ee4fca8eec389f, {16'd6343, 16'd24197, 16'd13870, 16'd6220, 16'd11522, 16'd9401, 16'd29466, 16'd55789, 16'd15634, 16'd34453, 16'd42806, 16'd12970, 16'd12028, 16'd61082, 16'd65329, 16'd3796, 16'd9493, 16'd46414, 16'd8358, 16'd56692, 16'd41173, 16'd28332, 16'd3211, 16'd12992, 16'd17124, 16'd43951});
	test_expansion(128'h13e7cb0122c93294ac61b30e4c24751f, {16'd61434, 16'd23700, 16'd45808, 16'd52249, 16'd19363, 16'd8289, 16'd55396, 16'd12730, 16'd19725, 16'd34439, 16'd65531, 16'd50086, 16'd44487, 16'd12834, 16'd30535, 16'd37915, 16'd59010, 16'd16462, 16'd28882, 16'd55410, 16'd22402, 16'd35368, 16'd44578, 16'd44931, 16'd53359, 16'd56140});
	test_expansion(128'h6cf0c7dd40e1bb332c63a0f7241b82dd, {16'd51511, 16'd25122, 16'd27972, 16'd34270, 16'd64735, 16'd58498, 16'd42144, 16'd46657, 16'd26659, 16'd63158, 16'd64305, 16'd56010, 16'd8744, 16'd56557, 16'd26575, 16'd27311, 16'd30279, 16'd26808, 16'd8836, 16'd59304, 16'd63019, 16'd50065, 16'd14292, 16'd65085, 16'd29092, 16'd25321});
	test_expansion(128'hb02c8424560be6d4df761382507c2af3, {16'd33254, 16'd57358, 16'd63881, 16'd26080, 16'd60202, 16'd38177, 16'd16596, 16'd57090, 16'd44146, 16'd28974, 16'd34845, 16'd10646, 16'd7614, 16'd7230, 16'd47667, 16'd28413, 16'd15903, 16'd1297, 16'd12215, 16'd57359, 16'd43853, 16'd64153, 16'd32222, 16'd41056, 16'd46977, 16'd38428});
	test_expansion(128'h50e6a95613347017af25bcf6cbdd1c7e, {16'd22281, 16'd13128, 16'd21452, 16'd33507, 16'd47309, 16'd64837, 16'd8502, 16'd63215, 16'd6020, 16'd33359, 16'd37814, 16'd5542, 16'd16264, 16'd8488, 16'd1405, 16'd44357, 16'd15631, 16'd56944, 16'd7327, 16'd58150, 16'd42103, 16'd64088, 16'd9783, 16'd22246, 16'd41771, 16'd43679});
	test_expansion(128'he65c281e892def3e440dcc0070a35fb1, {16'd31550, 16'd45927, 16'd30792, 16'd23249, 16'd50728, 16'd49944, 16'd63346, 16'd64854, 16'd49473, 16'd44169, 16'd38129, 16'd53540, 16'd18736, 16'd6725, 16'd17814, 16'd57176, 16'd30818, 16'd2737, 16'd32213, 16'd61570, 16'd7041, 16'd15990, 16'd21099, 16'd3747, 16'd37803, 16'd44401});
	test_expansion(128'h699b9d2da45f5e7d790522fad9dc6750, {16'd35617, 16'd54125, 16'd16640, 16'd56897, 16'd23319, 16'd20084, 16'd9233, 16'd52892, 16'd3641, 16'd52264, 16'd56434, 16'd833, 16'd7570, 16'd30925, 16'd24874, 16'd23046, 16'd34800, 16'd4683, 16'd53311, 16'd4109, 16'd43506, 16'd59786, 16'd40819, 16'd44215, 16'd34201, 16'd9259});
	test_expansion(128'h3ba9efe444eda4ed73947c171683ca2f, {16'd2240, 16'd61984, 16'd36744, 16'd23134, 16'd8356, 16'd5869, 16'd20368, 16'd28405, 16'd6433, 16'd3269, 16'd5857, 16'd11107, 16'd26404, 16'd55876, 16'd63065, 16'd1463, 16'd15709, 16'd37030, 16'd48934, 16'd18478, 16'd62501, 16'd29237, 16'd46342, 16'd21750, 16'd54102, 16'd24971});
	test_expansion(128'h83ff994ead3b3309c7f5fc487417ce2c, {16'd53059, 16'd55491, 16'd9232, 16'd29782, 16'd46243, 16'd9329, 16'd49111, 16'd61779, 16'd27764, 16'd60749, 16'd24314, 16'd13105, 16'd50399, 16'd44832, 16'd43964, 16'd26368, 16'd35813, 16'd49290, 16'd53963, 16'd6525, 16'd48026, 16'd54857, 16'd17306, 16'd21868, 16'd57711, 16'd59323});
	test_expansion(128'h9d9cdeb162a85aa269b4e4ad4025186f, {16'd35025, 16'd37004, 16'd27097, 16'd56215, 16'd17603, 16'd65165, 16'd28825, 16'd9385, 16'd17363, 16'd55999, 16'd7616, 16'd53363, 16'd9323, 16'd46856, 16'd51407, 16'd34687, 16'd50035, 16'd52139, 16'd57972, 16'd6483, 16'd36779, 16'd6467, 16'd49071, 16'd14622, 16'd29025, 16'd45367});
	test_expansion(128'hf095f5ca56bb35a6914199ee08683016, {16'd12396, 16'd51357, 16'd30943, 16'd58874, 16'd56032, 16'd32199, 16'd24955, 16'd61290, 16'd58974, 16'd53210, 16'd28373, 16'd39366, 16'd48282, 16'd63424, 16'd36166, 16'd46406, 16'd64249, 16'd3881, 16'd46217, 16'd32336, 16'd28546, 16'd19075, 16'd13611, 16'd43094, 16'd37931, 16'd33522});
	test_expansion(128'h966307cafbbe7c83e71ed751d35101a7, {16'd31715, 16'd62774, 16'd63117, 16'd13979, 16'd45962, 16'd25136, 16'd34120, 16'd55545, 16'd59087, 16'd46782, 16'd12740, 16'd21488, 16'd40055, 16'd49719, 16'd22030, 16'd25586, 16'd9399, 16'd33331, 16'd46983, 16'd36978, 16'd60589, 16'd6093, 16'd4627, 16'd64056, 16'd26034, 16'd19248});
	test_expansion(128'he78a438b09a005441cdff9baa8b8e40a, {16'd31995, 16'd61343, 16'd38091, 16'd28941, 16'd31854, 16'd39814, 16'd57575, 16'd40585, 16'd20799, 16'd8882, 16'd61787, 16'd11696, 16'd11433, 16'd52766, 16'd37997, 16'd7968, 16'd42613, 16'd46034, 16'd7523, 16'd11640, 16'd63698, 16'd31312, 16'd61792, 16'd34134, 16'd51029, 16'd32112});
	test_expansion(128'h80100759551672d60ea4ea9761a3df92, {16'd58087, 16'd37168, 16'd50850, 16'd45575, 16'd19490, 16'd23446, 16'd12602, 16'd9948, 16'd63435, 16'd16639, 16'd26444, 16'd2724, 16'd30926, 16'd37509, 16'd21969, 16'd14778, 16'd57229, 16'd960, 16'd23831, 16'd18370, 16'd49396, 16'd3689, 16'd20080, 16'd44682, 16'd5240, 16'd65382});
	test_expansion(128'hc90e7d356d5e23b6c8420adaf857ee93, {16'd52306, 16'd42830, 16'd39263, 16'd12157, 16'd46661, 16'd35868, 16'd44056, 16'd51845, 16'd43460, 16'd7716, 16'd4671, 16'd40487, 16'd33207, 16'd25803, 16'd9659, 16'd59566, 16'd55953, 16'd23319, 16'd53906, 16'd50946, 16'd43299, 16'd56819, 16'd21082, 16'd31186, 16'd17975, 16'd24507});
	test_expansion(128'h14c1aab19aecdeb647d1d146fe6c472d, {16'd6635, 16'd52849, 16'd1426, 16'd44430, 16'd10656, 16'd10298, 16'd19432, 16'd17635, 16'd64772, 16'd6384, 16'd37224, 16'd61085, 16'd28449, 16'd23571, 16'd41275, 16'd10962, 16'd57580, 16'd32764, 16'd23920, 16'd23422, 16'd9781, 16'd15273, 16'd1467, 16'd16805, 16'd23121, 16'd144});
	test_expansion(128'h2d6b5e3b0f11c33a26d331385ffd05eb, {16'd40303, 16'd42100, 16'd12877, 16'd57667, 16'd7515, 16'd4881, 16'd43196, 16'd46272, 16'd8304, 16'd615, 16'd16807, 16'd42226, 16'd4694, 16'd60563, 16'd13892, 16'd23751, 16'd48840, 16'd8352, 16'd10037, 16'd56435, 16'd55777, 16'd43795, 16'd38344, 16'd4843, 16'd4526, 16'd24576});
	test_expansion(128'hd95be9ca44be0acc4f2af4dd811c15f4, {16'd56111, 16'd9089, 16'd61507, 16'd41090, 16'd56898, 16'd44997, 16'd18063, 16'd30165, 16'd16701, 16'd64940, 16'd45409, 16'd34617, 16'd59122, 16'd3759, 16'd22244, 16'd61769, 16'd25163, 16'd48524, 16'd55973, 16'd4064, 16'd40640, 16'd38241, 16'd33717, 16'd61242, 16'd27807, 16'd20762});
	test_expansion(128'h6934180a782bd79aa2b72f0c593de0f3, {16'd51399, 16'd20069, 16'd19172, 16'd58448, 16'd25043, 16'd57142, 16'd53966, 16'd23135, 16'd22302, 16'd12789, 16'd39712, 16'd8914, 16'd39010, 16'd59853, 16'd38084, 16'd58897, 16'd41188, 16'd65158, 16'd59708, 16'd50568, 16'd6175, 16'd40035, 16'd45167, 16'd8683, 16'd34269, 16'd28802});
	test_expansion(128'h8eb63a46101128977df21e03084f3398, {16'd10552, 16'd35358, 16'd45705, 16'd1176, 16'd28189, 16'd21502, 16'd17455, 16'd40310, 16'd45749, 16'd46073, 16'd47214, 16'd1461, 16'd28623, 16'd50491, 16'd40317, 16'd24047, 16'd32378, 16'd43341, 16'd13637, 16'd33784, 16'd50542, 16'd58249, 16'd28520, 16'd49298, 16'd64110, 16'd27068});
	test_expansion(128'hadc7e125dba5f65553488a2c7305559f, {16'd8874, 16'd36263, 16'd22952, 16'd28155, 16'd17630, 16'd20823, 16'd17333, 16'd21660, 16'd48421, 16'd58295, 16'd12252, 16'd36044, 16'd6578, 16'd34837, 16'd45682, 16'd57864, 16'd31834, 16'd1468, 16'd47973, 16'd6377, 16'd35659, 16'd12293, 16'd58919, 16'd59585, 16'd59176, 16'd34096});
	test_expansion(128'hc406bff5a06cbe9a0f021e8b21a2c107, {16'd10351, 16'd35303, 16'd52950, 16'd38026, 16'd25824, 16'd37886, 16'd21037, 16'd24340, 16'd8417, 16'd58940, 16'd53972, 16'd35579, 16'd23188, 16'd98, 16'd29466, 16'd44410, 16'd17986, 16'd35261, 16'd33473, 16'd10740, 16'd5616, 16'd21514, 16'd53914, 16'd10620, 16'd17974, 16'd46825});
	test_expansion(128'h61cbaeb89eafc4b1936d01a1bbb74b0d, {16'd29376, 16'd51777, 16'd52687, 16'd1369, 16'd26228, 16'd36718, 16'd51069, 16'd41371, 16'd26311, 16'd46628, 16'd12392, 16'd8710, 16'd61905, 16'd12080, 16'd23883, 16'd30045, 16'd35087, 16'd26692, 16'd8112, 16'd50976, 16'd19799, 16'd31695, 16'd46363, 16'd35095, 16'd45892, 16'd16180});
	test_expansion(128'h6cac006716752d09f183dbc30f3ec35f, {16'd7257, 16'd62055, 16'd28394, 16'd64183, 16'd33860, 16'd18669, 16'd51277, 16'd13417, 16'd5901, 16'd10208, 16'd17194, 16'd23711, 16'd26780, 16'd15250, 16'd60208, 16'd51470, 16'd52906, 16'd30567, 16'd12452, 16'd50474, 16'd14656, 16'd5372, 16'd16333, 16'd35837, 16'd58241, 16'd15479});
	test_expansion(128'hcf5914fa0fa7cf9339fa254278ec2b37, {16'd54894, 16'd2689, 16'd53965, 16'd58227, 16'd9649, 16'd50779, 16'd23248, 16'd37292, 16'd8291, 16'd39376, 16'd18770, 16'd36273, 16'd40485, 16'd7506, 16'd51865, 16'd36040, 16'd59222, 16'd44972, 16'd27834, 16'd24949, 16'd9880, 16'd58654, 16'd27595, 16'd1478, 16'd29925, 16'd11265});
	test_expansion(128'he326c71e556e637f9e868e98608a84f2, {16'd50876, 16'd28111, 16'd16991, 16'd51284, 16'd48774, 16'd1628, 16'd29927, 16'd44361, 16'd60176, 16'd48451, 16'd40983, 16'd33151, 16'd34436, 16'd61038, 16'd30008, 16'd36304, 16'd9443, 16'd20605, 16'd59021, 16'd35277, 16'd2467, 16'd58367, 16'd13863, 16'd32370, 16'd52463, 16'd33546});
	test_expansion(128'h189ae12402507b83fbf77b417299c753, {16'd17502, 16'd43153, 16'd48856, 16'd36392, 16'd10345, 16'd22805, 16'd62390, 16'd11835, 16'd63354, 16'd18124, 16'd48044, 16'd5938, 16'd56456, 16'd11868, 16'd44777, 16'd64583, 16'd29134, 16'd58171, 16'd35492, 16'd17833, 16'd29623, 16'd45607, 16'd36164, 16'd405, 16'd41317, 16'd49277});
	test_expansion(128'h937476eb432349e3ece36b09ff56f8dd, {16'd28880, 16'd42443, 16'd8422, 16'd43614, 16'd33361, 16'd9126, 16'd49830, 16'd40650, 16'd37716, 16'd31418, 16'd12913, 16'd15865, 16'd7378, 16'd17956, 16'd63170, 16'd29165, 16'd19578, 16'd28752, 16'd43718, 16'd32482, 16'd30, 16'd14642, 16'd56281, 16'd43449, 16'd5196, 16'd39462});
	test_expansion(128'hc44e318b7901038d14dd72a8c6aeea7a, {16'd5596, 16'd39078, 16'd63336, 16'd6404, 16'd51632, 16'd50086, 16'd2586, 16'd12338, 16'd51953, 16'd46397, 16'd25358, 16'd23692, 16'd40409, 16'd8633, 16'd244, 16'd17430, 16'd43154, 16'd31313, 16'd54281, 16'd65159, 16'd38315, 16'd7254, 16'd53883, 16'd51347, 16'd24658, 16'd59859});
	test_expansion(128'h5ec423f5b40de4e85e0730c2489440f0, {16'd8190, 16'd33288, 16'd56223, 16'd36767, 16'd48423, 16'd29779, 16'd51458, 16'd42313, 16'd7427, 16'd61608, 16'd19251, 16'd57707, 16'd2297, 16'd33220, 16'd65445, 16'd4636, 16'd63840, 16'd34465, 16'd45650, 16'd41793, 16'd41040, 16'd38025, 16'd22016, 16'd19804, 16'd27701, 16'd58065});
	test_expansion(128'hd48375d3e85bbcdf0588a19734e05937, {16'd55618, 16'd1487, 16'd60936, 16'd60771, 16'd43934, 16'd7128, 16'd18418, 16'd45057, 16'd34376, 16'd39903, 16'd49341, 16'd64937, 16'd38882, 16'd4554, 16'd60533, 16'd890, 16'd38222, 16'd49025, 16'd9806, 16'd31544, 16'd3608, 16'd25084, 16'd41201, 16'd37680, 16'd52702, 16'd22967});
	test_expansion(128'hdad2fe9e25c333a2590bf5aef8d14f6b, {16'd28543, 16'd259, 16'd64040, 16'd37375, 16'd35681, 16'd18567, 16'd22461, 16'd35641, 16'd12085, 16'd43756, 16'd385, 16'd36527, 16'd61175, 16'd4238, 16'd31597, 16'd27260, 16'd18973, 16'd37558, 16'd45956, 16'd20705, 16'd33354, 16'd36811, 16'd53547, 16'd57785, 16'd1830, 16'd6802});
	test_expansion(128'h1a77ce5bb327923f7545b89d4767346b, {16'd16280, 16'd29145, 16'd61581, 16'd52253, 16'd39313, 16'd32976, 16'd9551, 16'd16697, 16'd43730, 16'd29147, 16'd7328, 16'd38246, 16'd22309, 16'd43639, 16'd11006, 16'd46388, 16'd12076, 16'd38415, 16'd59378, 16'd15060, 16'd30688, 16'd48962, 16'd26911, 16'd45487, 16'd16807, 16'd50086});
	test_expansion(128'h123a84262c172c41443afe5c11fdc282, {16'd33738, 16'd47249, 16'd14312, 16'd4374, 16'd22427, 16'd4333, 16'd10542, 16'd13083, 16'd35147, 16'd63926, 16'd40339, 16'd48523, 16'd59973, 16'd43620, 16'd41683, 16'd30266, 16'd55087, 16'd53336, 16'd26567, 16'd39768, 16'd33222, 16'd56834, 16'd57703, 16'd47966, 16'd64616, 16'd24039});
	test_expansion(128'h4bc53487d551446a507413981f157295, {16'd40377, 16'd827, 16'd42659, 16'd53444, 16'd12704, 16'd48963, 16'd27614, 16'd47416, 16'd39606, 16'd47065, 16'd65203, 16'd3268, 16'd59050, 16'd12097, 16'd45278, 16'd17767, 16'd41216, 16'd57580, 16'd26675, 16'd12031, 16'd17719, 16'd58652, 16'd40749, 16'd56733, 16'd52241, 16'd34082});
	test_expansion(128'hef1d4b248d29e57eb444fa560ceaa9ab, {16'd51955, 16'd62668, 16'd13442, 16'd27219, 16'd4015, 16'd46286, 16'd21069, 16'd12273, 16'd57073, 16'd13003, 16'd59461, 16'd13679, 16'd47624, 16'd41072, 16'd62700, 16'd26191, 16'd18361, 16'd25340, 16'd3929, 16'd17285, 16'd36707, 16'd48847, 16'd22637, 16'd22330, 16'd62849, 16'd16185});
	test_expansion(128'ha2f889122659e1bdd6af61432c4ce2a7, {16'd52102, 16'd65020, 16'd18414, 16'd35329, 16'd2727, 16'd5849, 16'd53023, 16'd55093, 16'd14266, 16'd26044, 16'd5025, 16'd45887, 16'd47592, 16'd23810, 16'd16500, 16'd4147, 16'd19969, 16'd46453, 16'd45870, 16'd59221, 16'd1201, 16'd2514, 16'd26645, 16'd33801, 16'd64832, 16'd31456});
	test_expansion(128'hd6e53366db42bfc5d13ddaa8b45c48d3, {16'd60699, 16'd41482, 16'd41176, 16'd2176, 16'd28682, 16'd56507, 16'd2086, 16'd31615, 16'd48850, 16'd48307, 16'd23654, 16'd45329, 16'd10983, 16'd63055, 16'd47355, 16'd8461, 16'd30740, 16'd1130, 16'd54053, 16'd24256, 16'd19218, 16'd55389, 16'd59367, 16'd58939, 16'd50837, 16'd7582});
	test_expansion(128'hd93f104d359e37bc1750a9bb6dac5992, {16'd8644, 16'd10443, 16'd58147, 16'd59039, 16'd5745, 16'd10282, 16'd31788, 16'd30859, 16'd8522, 16'd55698, 16'd32053, 16'd56640, 16'd49965, 16'd9742, 16'd21091, 16'd30452, 16'd57069, 16'd19580, 16'd5770, 16'd30260, 16'd52, 16'd28420, 16'd30546, 16'd45115, 16'd43888, 16'd37940});
	test_expansion(128'h552ec654d7d9be72895c0a22cd268ca5, {16'd30357, 16'd9651, 16'd9673, 16'd29254, 16'd47109, 16'd935, 16'd28952, 16'd42619, 16'd15991, 16'd40672, 16'd25909, 16'd32824, 16'd9580, 16'd55821, 16'd13649, 16'd50317, 16'd763, 16'd23315, 16'd31859, 16'd62952, 16'd5784, 16'd2465, 16'd32154, 16'd34945, 16'd3557, 16'd29087});
	test_expansion(128'h479ced42c1e1321fa516243147ac695c, {16'd31331, 16'd49062, 16'd44175, 16'd44249, 16'd26852, 16'd2104, 16'd56048, 16'd19082, 16'd46727, 16'd42302, 16'd45528, 16'd38619, 16'd49514, 16'd45854, 16'd41227, 16'd62941, 16'd36284, 16'd13990, 16'd1352, 16'd47993, 16'd53989, 16'd45211, 16'd53817, 16'd5731, 16'd17563, 16'd20225});
	test_expansion(128'hb91d7fdc6b10c378a0690ca3537a527f, {16'd2842, 16'd17805, 16'd12722, 16'd38272, 16'd37772, 16'd41649, 16'd65345, 16'd18373, 16'd26305, 16'd49026, 16'd35899, 16'd30153, 16'd39763, 16'd15079, 16'd50127, 16'd35114, 16'd34944, 16'd50891, 16'd14545, 16'd51240, 16'd31350, 16'd2261, 16'd43426, 16'd35009, 16'd52152, 16'd37179});
	test_expansion(128'h8cf920a9aefd2c7be04d18c7d5c1854f, {16'd13245, 16'd12851, 16'd60576, 16'd48366, 16'd18710, 16'd50658, 16'd34322, 16'd11088, 16'd37375, 16'd50474, 16'd12372, 16'd8093, 16'd25250, 16'd13301, 16'd57968, 16'd679, 16'd5764, 16'd32782, 16'd22979, 16'd49670, 16'd18799, 16'd37349, 16'd26084, 16'd53731, 16'd22595, 16'd9618});
	test_expansion(128'ha2e0e0d7ec8d9db6968aac7bbff2e4bc, {16'd16944, 16'd31957, 16'd60016, 16'd23485, 16'd29756, 16'd21024, 16'd48149, 16'd62304, 16'd63623, 16'd8191, 16'd39497, 16'd10125, 16'd15732, 16'd53143, 16'd13692, 16'd50530, 16'd58776, 16'd37097, 16'd49851, 16'd56051, 16'd16538, 16'd60809, 16'd7367, 16'd60586, 16'd36209, 16'd50717});
	test_expansion(128'h2dc130341892c98da720f2cb28b38590, {16'd22649, 16'd17432, 16'd58933, 16'd61710, 16'd50415, 16'd41141, 16'd37777, 16'd2819, 16'd42900, 16'd47872, 16'd63551, 16'd8373, 16'd55039, 16'd63464, 16'd6028, 16'd29564, 16'd37617, 16'd39888, 16'd45489, 16'd3357, 16'd59259, 16'd21511, 16'd34204, 16'd43381, 16'd25614, 16'd39096});
	test_expansion(128'h53aa1bf6d6e32622faff3f4959c71013, {16'd40591, 16'd12108, 16'd40248, 16'd34231, 16'd25415, 16'd45455, 16'd6514, 16'd19035, 16'd64146, 16'd44512, 16'd2347, 16'd41060, 16'd3849, 16'd41634, 16'd41505, 16'd24383, 16'd22524, 16'd52882, 16'd13459, 16'd44383, 16'd32803, 16'd52412, 16'd13793, 16'd48928, 16'd56716, 16'd53261});
	test_expansion(128'h12cd1ff3f389bed9cb188eb5655e84c3, {16'd55445, 16'd56190, 16'd17530, 16'd32323, 16'd50623, 16'd43050, 16'd13210, 16'd38664, 16'd13462, 16'd583, 16'd8644, 16'd35944, 16'd50641, 16'd41450, 16'd25104, 16'd11513, 16'd36543, 16'd64529, 16'd61780, 16'd60459, 16'd58728, 16'd22927, 16'd38610, 16'd57635, 16'd11659, 16'd26338});
	test_expansion(128'hb811f6b38d05307211c913cc6ec7136a, {16'd34244, 16'd5031, 16'd29201, 16'd21712, 16'd57473, 16'd7702, 16'd53065, 16'd10839, 16'd54310, 16'd8357, 16'd6159, 16'd60309, 16'd55157, 16'd44597, 16'd19968, 16'd20500, 16'd616, 16'd18591, 16'd54971, 16'd38217, 16'd22195, 16'd3955, 16'd23065, 16'd64800, 16'd45119, 16'd61708});
	test_expansion(128'h654058e032864597f694ad129b0f0b04, {16'd57909, 16'd27172, 16'd1189, 16'd33625, 16'd34039, 16'd60399, 16'd43989, 16'd48616, 16'd46999, 16'd57326, 16'd52077, 16'd22808, 16'd49308, 16'd33330, 16'd11180, 16'd45520, 16'd25184, 16'd29491, 16'd22322, 16'd34012, 16'd59990, 16'd29688, 16'd36905, 16'd7521, 16'd18353, 16'd11943});
	test_expansion(128'hb52216945bcf795035d3215a4ff68d0c, {16'd53273, 16'd40997, 16'd58957, 16'd30801, 16'd36700, 16'd23098, 16'd46344, 16'd14270, 16'd23983, 16'd48573, 16'd29754, 16'd17442, 16'd15988, 16'd30391, 16'd55373, 16'd58648, 16'd19298, 16'd48593, 16'd33937, 16'd50086, 16'd35525, 16'd40078, 16'd34630, 16'd31670, 16'd53671, 16'd21929});
	test_expansion(128'h5e61df75d901cf6b1ed36083f9004b0f, {16'd32298, 16'd38819, 16'd59887, 16'd15519, 16'd61704, 16'd37964, 16'd37408, 16'd24573, 16'd32851, 16'd41569, 16'd21201, 16'd11427, 16'd22551, 16'd52196, 16'd13442, 16'd20730, 16'd2774, 16'd5682, 16'd50315, 16'd10017, 16'd29277, 16'd39885, 16'd53148, 16'd17297, 16'd35107, 16'd53576});
	test_expansion(128'h2add1f7fde01205684ecc816e53250bf, {16'd48120, 16'd6774, 16'd3924, 16'd37124, 16'd51112, 16'd11211, 16'd38098, 16'd35922, 16'd39603, 16'd35221, 16'd64528, 16'd32284, 16'd60501, 16'd19614, 16'd60963, 16'd33065, 16'd33660, 16'd18664, 16'd12576, 16'd60264, 16'd6196, 16'd57432, 16'd36126, 16'd21460, 16'd10571, 16'd7110});
	test_expansion(128'h90c76ee6f5f5a7511e4522c12da7a034, {16'd29737, 16'd26286, 16'd9260, 16'd3784, 16'd40986, 16'd25131, 16'd33673, 16'd13586, 16'd38919, 16'd39589, 16'd24332, 16'd45465, 16'd19060, 16'd29103, 16'd28268, 16'd59887, 16'd31582, 16'd44407, 16'd3661, 16'd62463, 16'd38881, 16'd44983, 16'd9167, 16'd59, 16'd3040, 16'd47839});
	test_expansion(128'h1a14c23577313904a87f759928a1f75b, {16'd6690, 16'd28987, 16'd21825, 16'd24106, 16'd28299, 16'd50159, 16'd7252, 16'd15544, 16'd29265, 16'd41849, 16'd41335, 16'd7499, 16'd6775, 16'd62749, 16'd24758, 16'd554, 16'd57395, 16'd48108, 16'd29226, 16'd12085, 16'd44941, 16'd56271, 16'd50102, 16'd58562, 16'd65024, 16'd61370});
	test_expansion(128'hae17a4ce5ab969b4bfb9de5cc6810605, {16'd4350, 16'd23550, 16'd11830, 16'd17552, 16'd20191, 16'd45050, 16'd64328, 16'd20259, 16'd40158, 16'd1373, 16'd11511, 16'd28103, 16'd17599, 16'd29496, 16'd8539, 16'd1514, 16'd4252, 16'd8357, 16'd6569, 16'd1498, 16'd60365, 16'd2556, 16'd27633, 16'd4514, 16'd17733, 16'd34284});
	test_expansion(128'h53481bee07b86185cc10a2ebb8056da9, {16'd45048, 16'd13490, 16'd1807, 16'd24680, 16'd22207, 16'd21446, 16'd7716, 16'd62500, 16'd53468, 16'd35369, 16'd34150, 16'd61199, 16'd29959, 16'd38646, 16'd58343, 16'd8934, 16'd28788, 16'd7633, 16'd65060, 16'd59737, 16'd15937, 16'd13742, 16'd48968, 16'd55314, 16'd28117, 16'd25738});
	test_expansion(128'h32fd60e8c2f885347c5975b3faace1aa, {16'd9593, 16'd3838, 16'd40290, 16'd44538, 16'd40935, 16'd23454, 16'd32752, 16'd38843, 16'd34832, 16'd15232, 16'd28571, 16'd39585, 16'd63160, 16'd1249, 16'd38836, 16'd28314, 16'd18065, 16'd34507, 16'd24858, 16'd39959, 16'd4344, 16'd16094, 16'd10563, 16'd63960, 16'd64855, 16'd5950});
	test_expansion(128'he72e83ff435ac7f072b99afafd16d096, {16'd19882, 16'd36721, 16'd29648, 16'd39652, 16'd61144, 16'd51304, 16'd56539, 16'd9350, 16'd10987, 16'd11085, 16'd951, 16'd33099, 16'd15966, 16'd16220, 16'd54899, 16'd1704, 16'd33636, 16'd1207, 16'd42954, 16'd40293, 16'd4495, 16'd41328, 16'd56716, 16'd32622, 16'd4192, 16'd30789});
	test_expansion(128'ha71d0d021f2b5cd7c1c035cced21ef22, {16'd23656, 16'd3234, 16'd20123, 16'd41138, 16'd51616, 16'd2938, 16'd23053, 16'd3292, 16'd47971, 16'd26864, 16'd61627, 16'd57841, 16'd29517, 16'd18127, 16'd8876, 16'd39960, 16'd47905, 16'd14870, 16'd47146, 16'd60428, 16'd6658, 16'd49223, 16'd43754, 16'd7690, 16'd37993, 16'd51346});
	test_expansion(128'h84441764d7d63beb1ea5146eedce6b94, {16'd36999, 16'd18200, 16'd53581, 16'd42325, 16'd44902, 16'd13733, 16'd31347, 16'd32237, 16'd52610, 16'd53940, 16'd11747, 16'd24819, 16'd65022, 16'd43224, 16'd35813, 16'd30308, 16'd61903, 16'd22938, 16'd59921, 16'd4550, 16'd54696, 16'd32453, 16'd64533, 16'd25653, 16'd19887, 16'd27572});
	test_expansion(128'h10f8645bd4a9f1e5021d1b03d829707c, {16'd63267, 16'd32149, 16'd35623, 16'd6023, 16'd4869, 16'd30798, 16'd4616, 16'd10719, 16'd29553, 16'd29870, 16'd49625, 16'd34468, 16'd18285, 16'd16004, 16'd24791, 16'd35290, 16'd28853, 16'd49353, 16'd39445, 16'd16485, 16'd7559, 16'd25544, 16'd37543, 16'd47704, 16'd5931, 16'd9411});
	test_expansion(128'hba75a56f38eea6e0d5207746272b74c4, {16'd10088, 16'd59218, 16'd16858, 16'd45836, 16'd4625, 16'd27858, 16'd41034, 16'd25640, 16'd13172, 16'd50864, 16'd7335, 16'd27361, 16'd47805, 16'd12472, 16'd11145, 16'd28215, 16'd31182, 16'd62572, 16'd45358, 16'd36753, 16'd42520, 16'd56877, 16'd45402, 16'd34534, 16'd56300, 16'd271});
	test_expansion(128'hcfbe9d428c9cc1f6056efab310b34544, {16'd7621, 16'd13092, 16'd53673, 16'd7792, 16'd49651, 16'd39473, 16'd16554, 16'd5615, 16'd9217, 16'd64152, 16'd1791, 16'd1242, 16'd40175, 16'd61993, 16'd10528, 16'd25790, 16'd3046, 16'd11110, 16'd18641, 16'd2562, 16'd58309, 16'd914, 16'd7660, 16'd44446, 16'd32940, 16'd41048});
	test_expansion(128'h5a92e69b008aa8a6ad02ee9608b550bb, {16'd35700, 16'd15106, 16'd29876, 16'd31694, 16'd18820, 16'd48797, 16'd60082, 16'd53571, 16'd30044, 16'd48331, 16'd54946, 16'd34374, 16'd17563, 16'd32530, 16'd43124, 16'd44063, 16'd44479, 16'd33741, 16'd30620, 16'd31199, 16'd62320, 16'd50502, 16'd47840, 16'd59325, 16'd6102, 16'd51413});
	test_expansion(128'h7a5e6fcbbb010537cf697c15eb256a38, {16'd61965, 16'd49262, 16'd51471, 16'd53184, 16'd40759, 16'd31157, 16'd16192, 16'd25338, 16'd47809, 16'd28421, 16'd30331, 16'd52580, 16'd33102, 16'd17748, 16'd54256, 16'd4150, 16'd58029, 16'd19577, 16'd13420, 16'd5426, 16'd36588, 16'd34608, 16'd27350, 16'd24386, 16'd62443, 16'd48981});
	test_expansion(128'h0210b13e628e79d88c26db562f4be760, {16'd51964, 16'd41473, 16'd10134, 16'd55300, 16'd25321, 16'd48648, 16'd1773, 16'd29447, 16'd57648, 16'd7945, 16'd23143, 16'd53378, 16'd11599, 16'd60932, 16'd33427, 16'd20359, 16'd20856, 16'd58835, 16'd14198, 16'd7661, 16'd57190, 16'd2769, 16'd36970, 16'd40397, 16'd108, 16'd35772});
	test_expansion(128'h7948cd84afd2ac85b1a42307669e430e, {16'd17054, 16'd64774, 16'd22043, 16'd22205, 16'd55314, 16'd28607, 16'd62148, 16'd12458, 16'd63708, 16'd941, 16'd11926, 16'd59866, 16'd13313, 16'd54579, 16'd19084, 16'd2502, 16'd55737, 16'd33322, 16'd41161, 16'd38204, 16'd2352, 16'd7394, 16'd9473, 16'd56429, 16'd20011, 16'd18955});
	test_expansion(128'h2941f3641fd25619814ad4bb09a56f73, {16'd4171, 16'd8519, 16'd47045, 16'd42950, 16'd43666, 16'd32062, 16'd42243, 16'd38104, 16'd58337, 16'd18872, 16'd13122, 16'd48315, 16'd5193, 16'd6437, 16'd7104, 16'd44289, 16'd55162, 16'd56606, 16'd38674, 16'd2376, 16'd61862, 16'd37490, 16'd59386, 16'd2635, 16'd57574, 16'd9988});
	test_expansion(128'h54182dbff3d3f7b3d5de6ec6cd0e22ab, {16'd28483, 16'd46122, 16'd13575, 16'd48054, 16'd20579, 16'd40169, 16'd12062, 16'd3736, 16'd56726, 16'd16571, 16'd13968, 16'd34941, 16'd15550, 16'd31392, 16'd46123, 16'd36883, 16'd23240, 16'd63540, 16'd29599, 16'd33567, 16'd3661, 16'd18634, 16'd10744, 16'd5199, 16'd26801, 16'd58711});
	test_expansion(128'hd845de9c3d9c9aaac0a189636f90432b, {16'd49710, 16'd40063, 16'd32050, 16'd10664, 16'd30467, 16'd41530, 16'd17666, 16'd31550, 16'd47149, 16'd30583, 16'd15591, 16'd33022, 16'd13378, 16'd18593, 16'd11711, 16'd46799, 16'd12603, 16'd28506, 16'd3197, 16'd62526, 16'd29360, 16'd50694, 16'd37957, 16'd53508, 16'd64189, 16'd40381});
	test_expansion(128'h5d74cc3555c4e983e0bf46d64b07f9db, {16'd40395, 16'd17269, 16'd8275, 16'd19565, 16'd17295, 16'd47928, 16'd8604, 16'd8619, 16'd44959, 16'd11014, 16'd62821, 16'd21726, 16'd36382, 16'd26670, 16'd23854, 16'd37780, 16'd40238, 16'd30400, 16'd5728, 16'd25929, 16'd5446, 16'd18873, 16'd39243, 16'd55032, 16'd5924, 16'd50594});
	test_expansion(128'h0dcf27e88694850e8e47674ca729a5b4, {16'd62755, 16'd6265, 16'd62686, 16'd43069, 16'd313, 16'd35007, 16'd59068, 16'd51460, 16'd35956, 16'd6792, 16'd36221, 16'd31674, 16'd11762, 16'd33261, 16'd62587, 16'd29278, 16'd37473, 16'd51751, 16'd8124, 16'd788, 16'd64077, 16'd45051, 16'd52322, 16'd58049, 16'd28865, 16'd60110});
	test_expansion(128'h340856e9f59502db6274ffbb3e180387, {16'd13457, 16'd2155, 16'd7257, 16'd62365, 16'd13996, 16'd8341, 16'd59096, 16'd3032, 16'd45675, 16'd35364, 16'd15763, 16'd21876, 16'd43012, 16'd19485, 16'd38848, 16'd37784, 16'd50020, 16'd36901, 16'd47040, 16'd2025, 16'd7702, 16'd30494, 16'd55195, 16'd7516, 16'd45612, 16'd3833});
	test_expansion(128'ha2d80f03676deabcddad6a3b7cdfc4db, {16'd27142, 16'd1030, 16'd63613, 16'd58088, 16'd51608, 16'd21523, 16'd46930, 16'd20298, 16'd36384, 16'd14654, 16'd62437, 16'd20746, 16'd47201, 16'd14970, 16'd9814, 16'd30457, 16'd38962, 16'd18613, 16'd11816, 16'd50807, 16'd16102, 16'd50803, 16'd5270, 16'd31084, 16'd63593, 16'd50963});
	test_expansion(128'hdbb3ad7c9e7e923864d881cdfbd220be, {16'd55076, 16'd29981, 16'd20756, 16'd32604, 16'd32634, 16'd10517, 16'd8825, 16'd44243, 16'd35931, 16'd8628, 16'd3912, 16'd49266, 16'd15101, 16'd54908, 16'd7219, 16'd33724, 16'd1965, 16'd30764, 16'd13839, 16'd36201, 16'd56515, 16'd58542, 16'd38102, 16'd10832, 16'd1879, 16'd40397});
	test_expansion(128'hbc7d2718ddb2c9b99c9982954d2ba8da, {16'd48299, 16'd31497, 16'd15341, 16'd63276, 16'd42244, 16'd29686, 16'd63517, 16'd51853, 16'd28343, 16'd16327, 16'd28681, 16'd11086, 16'd22135, 16'd42942, 16'd10082, 16'd28957, 16'd22325, 16'd33856, 16'd65330, 16'd58704, 16'd57496, 16'd54980, 16'd6758, 16'd28441, 16'd8596, 16'd60044});
	test_expansion(128'heafbf893acd8aeb5ea43055a66b5a327, {16'd5206, 16'd18701, 16'd33591, 16'd26236, 16'd32559, 16'd56361, 16'd33744, 16'd8759, 16'd60059, 16'd57471, 16'd57566, 16'd11731, 16'd62470, 16'd8440, 16'd28877, 16'd4485, 16'd21344, 16'd5444, 16'd63570, 16'd21602, 16'd7126, 16'd21260, 16'd49192, 16'd12584, 16'd6296, 16'd65101});
	test_expansion(128'he4d82f698c1dbcae9f8650c580d5479a, {16'd50386, 16'd56151, 16'd15004, 16'd59092, 16'd27279, 16'd27290, 16'd57810, 16'd32666, 16'd37988, 16'd42830, 16'd61826, 16'd11172, 16'd23966, 16'd48392, 16'd64742, 16'd26380, 16'd18104, 16'd31463, 16'd51345, 16'd33782, 16'd39965, 16'd55060, 16'd64333, 16'd24854, 16'd60913, 16'd17000});
	test_expansion(128'h24b27efaf6d78cb5488d34855965b91e, {16'd35523, 16'd28390, 16'd37897, 16'd35787, 16'd16510, 16'd50629, 16'd30674, 16'd30409, 16'd42789, 16'd3578, 16'd50801, 16'd37266, 16'd40629, 16'd39756, 16'd28755, 16'd62603, 16'd62426, 16'd61002, 16'd47413, 16'd59642, 16'd12143, 16'd36888, 16'd6332, 16'd60137, 16'd47461, 16'd52433});
	test_expansion(128'h9b4b9be0616aeaf1f7f4952c8412369d, {16'd20819, 16'd18417, 16'd31273, 16'd8240, 16'd36514, 16'd13230, 16'd35009, 16'd37631, 16'd25125, 16'd52304, 16'd47354, 16'd47221, 16'd41503, 16'd31263, 16'd27827, 16'd22673, 16'd44477, 16'd2287, 16'd40764, 16'd27394, 16'd40619, 16'd59930, 16'd20856, 16'd50262, 16'd11235, 16'd60257});
	test_expansion(128'h19fc77173b29c351d581feb4f7747c2f, {16'd20690, 16'd47624, 16'd21542, 16'd53392, 16'd13750, 16'd35868, 16'd24579, 16'd36584, 16'd24076, 16'd38234, 16'd16815, 16'd28683, 16'd61615, 16'd13076, 16'd55521, 16'd48667, 16'd60988, 16'd42356, 16'd20314, 16'd28072, 16'd7941, 16'd15976, 16'd52197, 16'd2249, 16'd60815, 16'd31743});
	test_expansion(128'ha81b6ce640969f2b60df88958059d7eb, {16'd20218, 16'd48586, 16'd19947, 16'd32125, 16'd7079, 16'd23456, 16'd8279, 16'd54230, 16'd48269, 16'd29505, 16'd6814, 16'd29497, 16'd1478, 16'd3423, 16'd55437, 16'd32902, 16'd33372, 16'd38470, 16'd60472, 16'd42537, 16'd34025, 16'd32698, 16'd63242, 16'd47351, 16'd210, 16'd22819});
	test_expansion(128'h0ff421afdae8a79ffd18af9573dca156, {16'd41754, 16'd32231, 16'd21377, 16'd41922, 16'd10480, 16'd38333, 16'd52615, 16'd51841, 16'd64624, 16'd27360, 16'd31616, 16'd12397, 16'd15687, 16'd41306, 16'd3679, 16'd25460, 16'd37374, 16'd2868, 16'd32349, 16'd18341, 16'd63692, 16'd50593, 16'd45494, 16'd42889, 16'd59446, 16'd21418});
	test_expansion(128'hbf00edea8972afcb45106ada3196941e, {16'd26508, 16'd46451, 16'd12288, 16'd27126, 16'd46719, 16'd27887, 16'd49941, 16'd41285, 16'd65368, 16'd12848, 16'd31430, 16'd64633, 16'd6741, 16'd31406, 16'd63872, 16'd5251, 16'd64039, 16'd11054, 16'd52528, 16'd51080, 16'd44318, 16'd35284, 16'd16173, 16'd52409, 16'd49088, 16'd38415});
	test_expansion(128'h10cc9842affa1b300804f7145a082c00, {16'd40343, 16'd38321, 16'd52519, 16'd28287, 16'd56607, 16'd20620, 16'd17931, 16'd32008, 16'd50775, 16'd29701, 16'd12917, 16'd27801, 16'd63515, 16'd3073, 16'd49821, 16'd2634, 16'd5192, 16'd29924, 16'd54636, 16'd56229, 16'd10612, 16'd62520, 16'd4927, 16'd28944, 16'd54237, 16'd3853});
	test_expansion(128'h6e3abc208e683dddf219a7734af36624, {16'd46754, 16'd21322, 16'd50021, 16'd61485, 16'd59677, 16'd39017, 16'd286, 16'd30699, 16'd37133, 16'd26027, 16'd37661, 16'd54883, 16'd28103, 16'd29670, 16'd63458, 16'd24189, 16'd31140, 16'd20633, 16'd17861, 16'd9106, 16'd34846, 16'd31555, 16'd31998, 16'd44250, 16'd31936, 16'd41911});
	test_expansion(128'hee9014267dca1944545032a95e581b39, {16'd38886, 16'd15390, 16'd7587, 16'd5206, 16'd8483, 16'd17527, 16'd59565, 16'd26104, 16'd24699, 16'd18658, 16'd57235, 16'd58116, 16'd60495, 16'd28163, 16'd15403, 16'd19129, 16'd33920, 16'd50192, 16'd38893, 16'd35060, 16'd11130, 16'd62965, 16'd52666, 16'd24177, 16'd19238, 16'd47055});
	test_expansion(128'h7a5c985618af74ac07e8e9ab8f9c3f85, {16'd3058, 16'd20922, 16'd10156, 16'd24667, 16'd25050, 16'd42074, 16'd18227, 16'd15645, 16'd6414, 16'd27096, 16'd922, 16'd18399, 16'd15187, 16'd35563, 16'd44329, 16'd36073, 16'd61293, 16'd44857, 16'd52662, 16'd45751, 16'd44944, 16'd3924, 16'd44500, 16'd58433, 16'd8539, 16'd47500});
	test_expansion(128'h110e075401d48a1f74b9f55466eb8437, {16'd32291, 16'd28488, 16'd39002, 16'd21453, 16'd7155, 16'd10476, 16'd40869, 16'd17140, 16'd59904, 16'd3603, 16'd57420, 16'd27192, 16'd25029, 16'd52546, 16'd42815, 16'd25862, 16'd3621, 16'd12603, 16'd29639, 16'd56223, 16'd1285, 16'd16595, 16'd7470, 16'd51419, 16'd10197, 16'd26182});
	test_expansion(128'h7ea6c4b3b4afd5e617339490031f66a9, {16'd4788, 16'd15362, 16'd42997, 16'd10177, 16'd51113, 16'd8664, 16'd38357, 16'd39476, 16'd24318, 16'd51572, 16'd30232, 16'd35, 16'd53701, 16'd65410, 16'd10344, 16'd25995, 16'd12613, 16'd30660, 16'd22597, 16'd58747, 16'd59794, 16'd40493, 16'd52819, 16'd64218, 16'd28097, 16'd40395});
	test_expansion(128'hccca1b81a8e8bb96a2bb755c358f4609, {16'd23242, 16'd63755, 16'd6758, 16'd52806, 16'd32793, 16'd37476, 16'd61535, 16'd61452, 16'd10814, 16'd4629, 16'd36710, 16'd63, 16'd8096, 16'd51282, 16'd27102, 16'd51807, 16'd1693, 16'd22131, 16'd4047, 16'd50174, 16'd54728, 16'd4499, 16'd1256, 16'd47729, 16'd40781, 16'd47056});
	test_expansion(128'hfbe545c1ae5afd6c0e88fd5458930827, {16'd30663, 16'd50755, 16'd16713, 16'd36975, 16'd51089, 16'd16655, 16'd52060, 16'd31957, 16'd51834, 16'd7578, 16'd10394, 16'd50963, 16'd65239, 16'd22485, 16'd47449, 16'd21493, 16'd34651, 16'd48316, 16'd21943, 16'd12763, 16'd55983, 16'd3473, 16'd36251, 16'd29178, 16'd59056, 16'd60284});
	test_expansion(128'h114f75bdbd12df5f861ff873d7e74d03, {16'd51103, 16'd50461, 16'd49605, 16'd22377, 16'd64046, 16'd47153, 16'd27295, 16'd39785, 16'd42505, 16'd8285, 16'd48215, 16'd8504, 16'd34274, 16'd3482, 16'd58870, 16'd60405, 16'd10528, 16'd53773, 16'd27765, 16'd16957, 16'd10943, 16'd16076, 16'd28254, 16'd61695, 16'd50212, 16'd46884});
	test_expansion(128'h1f8cfed1d19713c750c9779132311bd4, {16'd2833, 16'd26978, 16'd14736, 16'd61932, 16'd14367, 16'd18501, 16'd11787, 16'd10816, 16'd53439, 16'd45105, 16'd56245, 16'd62814, 16'd39416, 16'd63665, 16'd35168, 16'd22203, 16'd38523, 16'd21256, 16'd38814, 16'd16267, 16'd42149, 16'd58856, 16'd26272, 16'd48476, 16'd54613, 16'd3897});
	test_expansion(128'ha079b1255038b759b8c51a9a2c9b21fe, {16'd9107, 16'd48095, 16'd15560, 16'd32651, 16'd19799, 16'd25934, 16'd47041, 16'd6621, 16'd19611, 16'd62358, 16'd57270, 16'd27510, 16'd40103, 16'd50283, 16'd7588, 16'd12828, 16'd33671, 16'd51570, 16'd57509, 16'd34733, 16'd34729, 16'd42892, 16'd22833, 16'd3055, 16'd41949, 16'd57411});
	test_expansion(128'h6396173d673b33ea975c29efa56bc216, {16'd29130, 16'd17040, 16'd52587, 16'd29371, 16'd63280, 16'd14348, 16'd63980, 16'd56756, 16'd51174, 16'd56557, 16'd56534, 16'd57712, 16'd32352, 16'd64230, 16'd6580, 16'd64063, 16'd3719, 16'd40522, 16'd41259, 16'd22294, 16'd24383, 16'd6858, 16'd47865, 16'd18151, 16'd49424, 16'd36457});
	test_expansion(128'h54016a802fd9cb0c78c231471a903535, {16'd43211, 16'd15766, 16'd37290, 16'd26045, 16'd22057, 16'd18858, 16'd26373, 16'd42244, 16'd55771, 16'd58104, 16'd26090, 16'd26555, 16'd51951, 16'd31310, 16'd61346, 16'd23985, 16'd16765, 16'd64678, 16'd62926, 16'd57037, 16'd22112, 16'd16826, 16'd49827, 16'd36044, 16'd4086, 16'd63695});
	test_expansion(128'h8ea8dbc52a74e02665df277917c18037, {16'd15913, 16'd6621, 16'd21928, 16'd9759, 16'd33467, 16'd47733, 16'd86, 16'd63691, 16'd27740, 16'd6484, 16'd42899, 16'd14693, 16'd4703, 16'd8668, 16'd23384, 16'd12714, 16'd30280, 16'd11786, 16'd20211, 16'd50437, 16'd4260, 16'd56941, 16'd45246, 16'd47645, 16'd25193, 16'd8689});
	test_expansion(128'h91e717438d169ca59b39cc9b6eb75973, {16'd26020, 16'd1268, 16'd20292, 16'd16338, 16'd23588, 16'd16393, 16'd40354, 16'd64321, 16'd30296, 16'd5443, 16'd58761, 16'd55614, 16'd8289, 16'd8387, 16'd31399, 16'd25784, 16'd24188, 16'd27643, 16'd52011, 16'd35524, 16'd42965, 16'd45601, 16'd6443, 16'd56679, 16'd29611, 16'd9357});
	test_expansion(128'h8e66214e0ddfe2f5617a75fad2183951, {16'd59079, 16'd1770, 16'd34903, 16'd52391, 16'd38418, 16'd36192, 16'd60500, 16'd25332, 16'd38191, 16'd27236, 16'd1390, 16'd30002, 16'd55584, 16'd25176, 16'd64611, 16'd36296, 16'd40861, 16'd39429, 16'd62782, 16'd31291, 16'd23541, 16'd43451, 16'd42261, 16'd25568, 16'd36561, 16'd14086});
	test_expansion(128'hbce0b70d5b26171d2d08e6c656d8c58e, {16'd40588, 16'd43169, 16'd20512, 16'd45164, 16'd47430, 16'd41447, 16'd34858, 16'd44137, 16'd27827, 16'd24926, 16'd38437, 16'd18027, 16'd2185, 16'd11992, 16'd4958, 16'd30052, 16'd2576, 16'd10074, 16'd58273, 16'd8485, 16'd23197, 16'd20561, 16'd1619, 16'd3264, 16'd7806, 16'd48055});
	test_expansion(128'h774548f44bd05e168fad0d94cb762ab6, {16'd41212, 16'd49902, 16'd52303, 16'd24284, 16'd57104, 16'd51083, 16'd15223, 16'd4588, 16'd49193, 16'd15893, 16'd10332, 16'd50597, 16'd56747, 16'd4534, 16'd28745, 16'd37081, 16'd57419, 16'd32761, 16'd46442, 16'd37234, 16'd44029, 16'd65170, 16'd48014, 16'd7626, 16'd26729, 16'd58387});
	test_expansion(128'h53efe8d92d412e5ae0da155791d84db5, {16'd15445, 16'd21675, 16'd38464, 16'd18074, 16'd25492, 16'd46661, 16'd17974, 16'd6565, 16'd20587, 16'd14387, 16'd62331, 16'd6459, 16'd35622, 16'd33121, 16'd53489, 16'd11525, 16'd29574, 16'd34860, 16'd56588, 16'd54038, 16'd52644, 16'd4957, 16'd12211, 16'd27587, 16'd37625, 16'd34039});
	test_expansion(128'hf004d1ad427a46c14050bd4a13453bac, {16'd59981, 16'd19908, 16'd36055, 16'd43420, 16'd49123, 16'd38383, 16'd62697, 16'd43193, 16'd20073, 16'd9603, 16'd23715, 16'd7662, 16'd20984, 16'd50018, 16'd50303, 16'd65298, 16'd32675, 16'd42047, 16'd58723, 16'd40847, 16'd34897, 16'd28733, 16'd64191, 16'd36305, 16'd55872, 16'd51716});
	test_expansion(128'hd153b46d7c6df6b9144c133dfb91eff0, {16'd32626, 16'd64903, 16'd28568, 16'd7816, 16'd27377, 16'd33071, 16'd20008, 16'd48084, 16'd17415, 16'd61126, 16'd28750, 16'd18942, 16'd14930, 16'd59531, 16'd25589, 16'd48012, 16'd15854, 16'd57160, 16'd22639, 16'd62410, 16'd37315, 16'd4404, 16'd16932, 16'd2545, 16'd58586, 16'd39387});
	test_expansion(128'h13a7cceb0afabcb4d60e7ce38dcb813b, {16'd2508, 16'd53887, 16'd16560, 16'd11031, 16'd11243, 16'd57452, 16'd27905, 16'd61194, 16'd9176, 16'd42236, 16'd21908, 16'd35601, 16'd20812, 16'd40265, 16'd12544, 16'd29385, 16'd26285, 16'd919, 16'd30902, 16'd3797, 16'd44077, 16'd11811, 16'd3481, 16'd60654, 16'd52814, 16'd10742});
	test_expansion(128'h5240259ac63ecc8ace2c48eaf5f7e2b2, {16'd28472, 16'd47093, 16'd8881, 16'd59126, 16'd53042, 16'd32805, 16'd36147, 16'd45830, 16'd65056, 16'd19902, 16'd42567, 16'd23079, 16'd4467, 16'd8786, 16'd41314, 16'd13426, 16'd9098, 16'd15443, 16'd16939, 16'd14544, 16'd33016, 16'd18195, 16'd3601, 16'd60033, 16'd22045, 16'd39391});
	test_expansion(128'h40d4edbb212af4b9f1beecf7282e2a38, {16'd53729, 16'd55963, 16'd20845, 16'd11295, 16'd47546, 16'd11586, 16'd40395, 16'd56033, 16'd3282, 16'd55298, 16'd63389, 16'd31168, 16'd12778, 16'd22422, 16'd29831, 16'd31099, 16'd17298, 16'd41240, 16'd21607, 16'd44409, 16'd20591, 16'd16558, 16'd61200, 16'd6034, 16'd17974, 16'd31393});
	test_expansion(128'h44c880f408fa5f2cc642900afcd2e564, {16'd54617, 16'd43946, 16'd56086, 16'd24537, 16'd20918, 16'd36773, 16'd3386, 16'd22631, 16'd27115, 16'd27642, 16'd48409, 16'd18053, 16'd8156, 16'd10537, 16'd15003, 16'd63805, 16'd40272, 16'd31048, 16'd10149, 16'd53353, 16'd55616, 16'd377, 16'd53612, 16'd36309, 16'd32309, 16'd1827});
	test_expansion(128'hde2533081082cc6f752977d0bcf18f9f, {16'd35707, 16'd18079, 16'd1718, 16'd2379, 16'd28380, 16'd62021, 16'd46187, 16'd53345, 16'd56217, 16'd56099, 16'd33681, 16'd49696, 16'd11779, 16'd57829, 16'd18128, 16'd7625, 16'd22162, 16'd63653, 16'd40848, 16'd31893, 16'd63325, 16'd49399, 16'd27810, 16'd49951, 16'd39310, 16'd43421});
	test_expansion(128'h6b29b80e43ffd48ba42d47c55b41f14d, {16'd14617, 16'd26577, 16'd39510, 16'd32166, 16'd22379, 16'd5536, 16'd47428, 16'd61387, 16'd30182, 16'd21971, 16'd26032, 16'd42347, 16'd39200, 16'd36762, 16'd41481, 16'd25676, 16'd11481, 16'd3544, 16'd39756, 16'd37040, 16'd11256, 16'd42336, 16'd35244, 16'd56060, 16'd59624, 16'd34004});
	test_expansion(128'h04323375bc9442af0c68fc7bd1b47fb3, {16'd28890, 16'd18008, 16'd20782, 16'd18046, 16'd43741, 16'd2703, 16'd21009, 16'd14720, 16'd41986, 16'd9767, 16'd16569, 16'd39748, 16'd59222, 16'd27828, 16'd28553, 16'd46018, 16'd3314, 16'd2940, 16'd547, 16'd9684, 16'd40208, 16'd17970, 16'd12573, 16'd50816, 16'd20049, 16'd10846});
	test_expansion(128'hb15f9390a60b85a20b199301f503739a, {16'd42579, 16'd50475, 16'd32548, 16'd35227, 16'd34691, 16'd55744, 16'd54671, 16'd12579, 16'd21966, 16'd18998, 16'd6265, 16'd36773, 16'd24297, 16'd55983, 16'd57676, 16'd58973, 16'd44131, 16'd24217, 16'd49030, 16'd28188, 16'd56665, 16'd15857, 16'd14508, 16'd60956, 16'd18552, 16'd51746});
	test_expansion(128'h7b245d174045975646890ab3100e4380, {16'd21367, 16'd53940, 16'd33547, 16'd33679, 16'd5758, 16'd44459, 16'd25671, 16'd16621, 16'd25560, 16'd29795, 16'd59744, 16'd2145, 16'd19503, 16'd50314, 16'd704, 16'd45789, 16'd20832, 16'd19519, 16'd1989, 16'd56983, 16'd23583, 16'd32496, 16'd49035, 16'd6139, 16'd36857, 16'd2779});
	test_expansion(128'hf715f874068b579ee2717bdd89cf083b, {16'd58137, 16'd33630, 16'd41819, 16'd45844, 16'd42815, 16'd15950, 16'd19729, 16'd6948, 16'd13971, 16'd58557, 16'd43306, 16'd52972, 16'd20169, 16'd54047, 16'd61754, 16'd64032, 16'd14764, 16'd63, 16'd40072, 16'd14279, 16'd14677, 16'd25110, 16'd15322, 16'd20052, 16'd14055, 16'd11719});
	test_expansion(128'hd0c2c0561e16ac411b15b22d9056d83e, {16'd24694, 16'd42037, 16'd29015, 16'd7161, 16'd51926, 16'd60071, 16'd47753, 16'd5096, 16'd38557, 16'd62130, 16'd8853, 16'd2438, 16'd36821, 16'd23435, 16'd21899, 16'd6981, 16'd43170, 16'd11541, 16'd38734, 16'd22437, 16'd18556, 16'd44207, 16'd36586, 16'd11464, 16'd39282, 16'd43470});
	test_expansion(128'h141dceeee656d8766892757c33bb1b3f, {16'd9142, 16'd42175, 16'd2259, 16'd20845, 16'd62228, 16'd27184, 16'd12343, 16'd54877, 16'd62209, 16'd7372, 16'd48854, 16'd23454, 16'd14841, 16'd54108, 16'd59471, 16'd41234, 16'd45308, 16'd35466, 16'd1334, 16'd12073, 16'd29091, 16'd64687, 16'd22838, 16'd22621, 16'd25759, 16'd23640});
	test_expansion(128'h485a0a1a09d70c05a706cdcb37872135, {16'd34788, 16'd18824, 16'd10008, 16'd49471, 16'd19392, 16'd65139, 16'd39407, 16'd31174, 16'd25252, 16'd50780, 16'd7972, 16'd58280, 16'd52797, 16'd64407, 16'd57905, 16'd34539, 16'd43250, 16'd44171, 16'd62033, 16'd14921, 16'd44675, 16'd26989, 16'd36523, 16'd59417, 16'd5856, 16'd54889});
	test_expansion(128'h6292fb8285195c408826290a4dcf0fb7, {16'd24771, 16'd7848, 16'd23009, 16'd30818, 16'd60911, 16'd3915, 16'd48534, 16'd47162, 16'd13840, 16'd9843, 16'd42968, 16'd31797, 16'd17285, 16'd61869, 16'd64698, 16'd13592, 16'd30222, 16'd57847, 16'd696, 16'd29947, 16'd62014, 16'd2491, 16'd55628, 16'd10631, 16'd40222, 16'd54125});
	test_expansion(128'hcbd0c05e1a86dfa2d9ec9edc9734809a, {16'd52977, 16'd1498, 16'd14334, 16'd9802, 16'd29792, 16'd25178, 16'd43916, 16'd57503, 16'd62602, 16'd55199, 16'd64220, 16'd63654, 16'd46675, 16'd33008, 16'd62318, 16'd23152, 16'd13795, 16'd38183, 16'd18933, 16'd62627, 16'd36879, 16'd28609, 16'd29762, 16'd18387, 16'd18819, 16'd25331});
	test_expansion(128'h4540ed860e55fee6a5645cfada563e53, {16'd17937, 16'd8334, 16'd61493, 16'd43684, 16'd25390, 16'd60729, 16'd57045, 16'd34580, 16'd22930, 16'd39703, 16'd8479, 16'd9473, 16'd61954, 16'd62161, 16'd45797, 16'd4078, 16'd37537, 16'd615, 16'd57382, 16'd63620, 16'd40717, 16'd59205, 16'd47809, 16'd22275, 16'd50697, 16'd14228});
	test_expansion(128'hda6e349429505a533361d1722ffdd970, {16'd49351, 16'd51609, 16'd18309, 16'd52826, 16'd49388, 16'd39330, 16'd55349, 16'd25733, 16'd36583, 16'd55353, 16'd50856, 16'd8245, 16'd14795, 16'd9750, 16'd63669, 16'd33912, 16'd24903, 16'd40884, 16'd19948, 16'd11823, 16'd31861, 16'd51661, 16'd41839, 16'd12560, 16'd36210, 16'd47328});
	test_expansion(128'h5b6ef5d855a089e9923f926868c335b2, {16'd38628, 16'd9897, 16'd14663, 16'd22143, 16'd16388, 16'd40000, 16'd60539, 16'd58255, 16'd36371, 16'd7943, 16'd53183, 16'd16694, 16'd30584, 16'd36246, 16'd32688, 16'd713, 16'd10372, 16'd54445, 16'd46445, 16'd10835, 16'd34188, 16'd52570, 16'd30149, 16'd31297, 16'd30001, 16'd26154});
	test_expansion(128'h628a0b0adafb68f090cb1cb657fc667c, {16'd39468, 16'd2661, 16'd26983, 16'd35789, 16'd10701, 16'd8420, 16'd24201, 16'd58313, 16'd44716, 16'd38468, 16'd47359, 16'd12311, 16'd29263, 16'd45536, 16'd14098, 16'd24181, 16'd33480, 16'd21476, 16'd29315, 16'd3273, 16'd45400, 16'd40765, 16'd17955, 16'd30712, 16'd46208, 16'd3803});
	test_expansion(128'h5b15b9b65386fe5f75fafcbf09f77691, {16'd54795, 16'd15359, 16'd58576, 16'd62682, 16'd8693, 16'd50329, 16'd24882, 16'd21368, 16'd1914, 16'd33352, 16'd10604, 16'd17993, 16'd39640, 16'd20607, 16'd48694, 16'd40824, 16'd52779, 16'd54104, 16'd41559, 16'd57665, 16'd8438, 16'd25244, 16'd39056, 16'd50660, 16'd40365, 16'd3892});
	test_expansion(128'h0cec8c30291e4dbbfce33c481e3da03e, {16'd50379, 16'd55514, 16'd22196, 16'd16489, 16'd52136, 16'd4192, 16'd41554, 16'd46043, 16'd53512, 16'd63144, 16'd45843, 16'd7814, 16'd57722, 16'd41845, 16'd63984, 16'd30318, 16'd44785, 16'd64538, 16'd62720, 16'd3824, 16'd5439, 16'd7076, 16'd51461, 16'd44744, 16'd56932, 16'd1647});
	test_expansion(128'h9c28a1968698142b946620f6b99c1761, {16'd3779, 16'd34228, 16'd63431, 16'd53568, 16'd17352, 16'd46823, 16'd10318, 16'd3574, 16'd33620, 16'd28840, 16'd54308, 16'd41472, 16'd8668, 16'd46839, 16'd60292, 16'd25392, 16'd45823, 16'd63407, 16'd54160, 16'd1794, 16'd36255, 16'd40669, 16'd13695, 16'd57226, 16'd57690, 16'd28428});
	test_expansion(128'hb316f90560f665c94d3461d1c87f018f, {16'd59077, 16'd54859, 16'd44639, 16'd21662, 16'd4862, 16'd15988, 16'd53342, 16'd21177, 16'd1517, 16'd11596, 16'd62272, 16'd58498, 16'd48653, 16'd22695, 16'd21943, 16'd42730, 16'd12478, 16'd15162, 16'd63169, 16'd63470, 16'd61426, 16'd37853, 16'd53122, 16'd48414, 16'd26707, 16'd16610});
	test_expansion(128'h922fb3d49030127fb385b5ce9ec9115e, {16'd11833, 16'd53201, 16'd63707, 16'd37351, 16'd16069, 16'd3313, 16'd57432, 16'd65198, 16'd41447, 16'd35895, 16'd18533, 16'd42958, 16'd50316, 16'd30944, 16'd61533, 16'd11651, 16'd13828, 16'd59555, 16'd2733, 16'd14819, 16'd4, 16'd10257, 16'd37394, 16'd44720, 16'd1693, 16'd32519});
	test_expansion(128'hf42da3ad6947025d06f3c202040be3ac, {16'd47980, 16'd29488, 16'd56703, 16'd19918, 16'd28217, 16'd50982, 16'd184, 16'd55709, 16'd62707, 16'd55065, 16'd31476, 16'd50334, 16'd58086, 16'd48239, 16'd12156, 16'd53113, 16'd17604, 16'd44402, 16'd26527, 16'd12268, 16'd55234, 16'd719, 16'd39516, 16'd45813, 16'd10408, 16'd16219});
	test_expansion(128'h91bef60796e9592e2dd29457057811d9, {16'd42024, 16'd19347, 16'd44045, 16'd61812, 16'd30690, 16'd21320, 16'd45703, 16'd5112, 16'd8060, 16'd55538, 16'd25555, 16'd33591, 16'd39372, 16'd8957, 16'd4274, 16'd7954, 16'd40430, 16'd54534, 16'd56433, 16'd57115, 16'd17087, 16'd48571, 16'd33929, 16'd15573, 16'd47590, 16'd63207});
	test_expansion(128'h12fc46f4e3d372142184b8ceec1f171f, {16'd18631, 16'd54182, 16'd32485, 16'd42163, 16'd20623, 16'd54640, 16'd23640, 16'd20610, 16'd37991, 16'd26060, 16'd64764, 16'd59896, 16'd12701, 16'd41404, 16'd12400, 16'd53285, 16'd51250, 16'd27196, 16'd26896, 16'd46353, 16'd39916, 16'd43911, 16'd2732, 16'd10783, 16'd45851, 16'd40799});
	test_expansion(128'hf503a7861d38ed2b48eaddb544e276fb, {16'd1439, 16'd1828, 16'd3879, 16'd29943, 16'd4056, 16'd5639, 16'd20675, 16'd39935, 16'd50343, 16'd34676, 16'd41808, 16'd51042, 16'd10962, 16'd53404, 16'd20106, 16'd44576, 16'd41755, 16'd22067, 16'd6688, 16'd63013, 16'd3215, 16'd11204, 16'd51472, 16'd54590, 16'd36956, 16'd15621});
	test_expansion(128'h407e18be564eb0788b01e890d1c87605, {16'd1506, 16'd65283, 16'd59125, 16'd32251, 16'd18972, 16'd58139, 16'd62097, 16'd61657, 16'd654, 16'd57047, 16'd52012, 16'd43794, 16'd4479, 16'd9751, 16'd64499, 16'd46532, 16'd35777, 16'd5717, 16'd11877, 16'd12414, 16'd47015, 16'd39352, 16'd16728, 16'd37380, 16'd23847, 16'd12895});
	test_expansion(128'h14831d0e371eda45de5cbeb33935327b, {16'd33673, 16'd25142, 16'd36527, 16'd28502, 16'd48880, 16'd24714, 16'd12386, 16'd38434, 16'd37729, 16'd274, 16'd41663, 16'd4783, 16'd60935, 16'd37274, 16'd54597, 16'd58075, 16'd49274, 16'd63706, 16'd27474, 16'd4167, 16'd27266, 16'd55954, 16'd29520, 16'd47292, 16'd20511, 16'd40345});
	test_expansion(128'hf34eca05e654feeeca2a3f34276e2100, {16'd55410, 16'd60184, 16'd57270, 16'd43387, 16'd16186, 16'd15959, 16'd37819, 16'd54034, 16'd35572, 16'd19031, 16'd1476, 16'd8674, 16'd13335, 16'd45728, 16'd60552, 16'd41335, 16'd23048, 16'd12109, 16'd15126, 16'd8259, 16'd49901, 16'd52661, 16'd64592, 16'd31829, 16'd13667, 16'd22434});
	test_expansion(128'h85d96f788b301e65d06ee6606ebe26ec, {16'd72, 16'd48898, 16'd27063, 16'd60441, 16'd6835, 16'd14410, 16'd27090, 16'd337, 16'd41138, 16'd19127, 16'd12636, 16'd21395, 16'd7095, 16'd19290, 16'd37998, 16'd40153, 16'd56449, 16'd47569, 16'd16482, 16'd65139, 16'd23771, 16'd43139, 16'd11480, 16'd37558, 16'd57661, 16'd3303});
	test_expansion(128'hbd006718b377656b235dbf6571af8748, {16'd62405, 16'd26501, 16'd56042, 16'd46936, 16'd2652, 16'd45921, 16'd61787, 16'd58162, 16'd50868, 16'd38422, 16'd55565, 16'd27527, 16'd16720, 16'd45957, 16'd56664, 16'd31940, 16'd54336, 16'd61357, 16'd50050, 16'd45575, 16'd35894, 16'd19743, 16'd54401, 16'd63067, 16'd1293, 16'd64180});
	test_expansion(128'h885f7831fd2d27e4738811ef06f41ebc, {16'd44049, 16'd8295, 16'd59961, 16'd50818, 16'd13298, 16'd35240, 16'd26414, 16'd24920, 16'd33821, 16'd50889, 16'd56939, 16'd30037, 16'd11109, 16'd23271, 16'd54668, 16'd4335, 16'd39634, 16'd11668, 16'd21366, 16'd21659, 16'd61969, 16'd48048, 16'd49123, 16'd13393, 16'd50960, 16'd34211});
	test_expansion(128'h97af5a222d2cf32c65c3c96007dec5b2, {16'd8346, 16'd29225, 16'd60179, 16'd16844, 16'd45241, 16'd50466, 16'd30377, 16'd43260, 16'd25876, 16'd13077, 16'd43559, 16'd43986, 16'd35036, 16'd47546, 16'd16577, 16'd52981, 16'd65279, 16'd29617, 16'd30720, 16'd8579, 16'd52535, 16'd2396, 16'd33854, 16'd51726, 16'd9152, 16'd15685});
	test_expansion(128'ha9c30dc526da0f08e50f45ba8a9b8df5, {16'd24385, 16'd51271, 16'd54336, 16'd27583, 16'd9287, 16'd3583, 16'd3848, 16'd24419, 16'd48905, 16'd12080, 16'd6202, 16'd30761, 16'd15072, 16'd16033, 16'd3957, 16'd65238, 16'd28601, 16'd3251, 16'd7533, 16'd229, 16'd7673, 16'd50512, 16'd54386, 16'd6273, 16'd26400, 16'd49888});
	test_expansion(128'h2400aec876d89ea14c2d7d984d1748c9, {16'd7148, 16'd37340, 16'd31644, 16'd64859, 16'd17384, 16'd57727, 16'd58564, 16'd26797, 16'd30378, 16'd52183, 16'd43185, 16'd5366, 16'd18313, 16'd35376, 16'd3043, 16'd42019, 16'd57628, 16'd56424, 16'd20684, 16'd11486, 16'd16918, 16'd62990, 16'd7566, 16'd42941, 16'd27486, 16'd64798});
	test_expansion(128'h962c8992bfe36d93a8a7977413a88f83, {16'd39723, 16'd39980, 16'd22844, 16'd37526, 16'd40042, 16'd54317, 16'd55422, 16'd33665, 16'd56403, 16'd51082, 16'd42867, 16'd51041, 16'd6060, 16'd28811, 16'd2062, 16'd45595, 16'd58879, 16'd18700, 16'd52505, 16'd44846, 16'd17890, 16'd33712, 16'd43095, 16'd45195, 16'd3309, 16'd28769});
	test_expansion(128'he0ab521f2364253bf7b2ca566dcc5324, {16'd63054, 16'd55265, 16'd1956, 16'd53919, 16'd43632, 16'd52500, 16'd37735, 16'd32004, 16'd30947, 16'd34183, 16'd21148, 16'd52487, 16'd46335, 16'd14998, 16'd48360, 16'd7777, 16'd53831, 16'd64636, 16'd9869, 16'd51000, 16'd42449, 16'd46638, 16'd48967, 16'd37412, 16'd49177, 16'd37925});
	test_expansion(128'hff08ab97e9a347343170c6a72298cfdd, {16'd24559, 16'd46437, 16'd6026, 16'd31368, 16'd62315, 16'd877, 16'd32415, 16'd18996, 16'd52042, 16'd31924, 16'd42045, 16'd57463, 16'd48951, 16'd19938, 16'd55709, 16'd51724, 16'd17519, 16'd59570, 16'd54788, 16'd55420, 16'd17347, 16'd61682, 16'd1231, 16'd11643, 16'd27559, 16'd809});
	test_expansion(128'hb40ec9e45d210727ac3699735f35433e, {16'd26079, 16'd56365, 16'd50956, 16'd33859, 16'd63894, 16'd10896, 16'd5227, 16'd58686, 16'd32164, 16'd56580, 16'd42252, 16'd32606, 16'd13032, 16'd15033, 16'd35172, 16'd38549, 16'd37257, 16'd25270, 16'd63957, 16'd48859, 16'd2447, 16'd13167, 16'd16241, 16'd46379, 16'd50987, 16'd27953});
	test_expansion(128'h2e7f32c0b4bb18c58a312db2f9f9181b, {16'd45181, 16'd58253, 16'd24341, 16'd41912, 16'd63953, 16'd63927, 16'd64958, 16'd57386, 16'd31845, 16'd12975, 16'd9247, 16'd25982, 16'd14566, 16'd47987, 16'd23486, 16'd133, 16'd65297, 16'd57365, 16'd10167, 16'd29725, 16'd43547, 16'd20046, 16'd19069, 16'd36529, 16'd55306, 16'd9398});
	test_expansion(128'heb712b1f8ae9d741472c0d4b52b54375, {16'd3907, 16'd9055, 16'd17584, 16'd29397, 16'd14946, 16'd21520, 16'd32444, 16'd40613, 16'd5855, 16'd32931, 16'd26905, 16'd27733, 16'd64871, 16'd37755, 16'd13815, 16'd60905, 16'd14555, 16'd52994, 16'd6495, 16'd362, 16'd24920, 16'd45844, 16'd62085, 16'd15585, 16'd10028, 16'd59602});
	test_expansion(128'h0671e52e395abf71b841f9a2a5a776e7, {16'd21413, 16'd64233, 16'd36521, 16'd44126, 16'd63490, 16'd51279, 16'd20417, 16'd27270, 16'd41456, 16'd42815, 16'd50910, 16'd25841, 16'd56283, 16'd8551, 16'd33737, 16'd65122, 16'd15139, 16'd48334, 16'd23531, 16'd35680, 16'd15073, 16'd15181, 16'd63129, 16'd9736, 16'd52172, 16'd40847});
	test_expansion(128'h69391d7c83737a81559dc7f321992733, {16'd14552, 16'd42727, 16'd32305, 16'd61369, 16'd61686, 16'd33069, 16'd3550, 16'd13758, 16'd32507, 16'd57027, 16'd30665, 16'd21951, 16'd4134, 16'd50163, 16'd5810, 16'd1813, 16'd46991, 16'd38848, 16'd20791, 16'd56487, 16'd63284, 16'd25347, 16'd6248, 16'd65142, 16'd60949, 16'd26129});
	test_expansion(128'h90db63c5525dde189e6c725074b1c613, {16'd37738, 16'd12616, 16'd4063, 16'd58700, 16'd57358, 16'd54952, 16'd4161, 16'd15120, 16'd51827, 16'd13892, 16'd43086, 16'd37958, 16'd57879, 16'd17372, 16'd29969, 16'd50647, 16'd45178, 16'd7001, 16'd23531, 16'd53561, 16'd43787, 16'd27595, 16'd41363, 16'd50174, 16'd38581, 16'd57760});
	test_expansion(128'h835117e19de1943641629536c1ca3f80, {16'd63422, 16'd35723, 16'd35998, 16'd56190, 16'd5259, 16'd45199, 16'd17882, 16'd25105, 16'd22283, 16'd41065, 16'd64465, 16'd49686, 16'd24600, 16'd55490, 16'd20972, 16'd38594, 16'd14722, 16'd63452, 16'd51625, 16'd884, 16'd43770, 16'd61373, 16'd26983, 16'd41296, 16'd19475, 16'd9445});
	test_expansion(128'h7107efaa454a35649094d5e89428e018, {16'd60011, 16'd329, 16'd37243, 16'd2005, 16'd57037, 16'd11881, 16'd62323, 16'd48358, 16'd57401, 16'd16586, 16'd27702, 16'd41214, 16'd47231, 16'd6880, 16'd30552, 16'd34279, 16'd64951, 16'd11384, 16'd59215, 16'd52820, 16'd18405, 16'd64465, 16'd44695, 16'd55025, 16'd27234, 16'd21459});
	test_expansion(128'h76fab402c5b4767f4d4d733a6f94ba85, {16'd25951, 16'd30071, 16'd38527, 16'd19342, 16'd58041, 16'd21200, 16'd58461, 16'd32889, 16'd42451, 16'd27428, 16'd45204, 16'd51461, 16'd8801, 16'd17678, 16'd3300, 16'd52656, 16'd48543, 16'd567, 16'd40529, 16'd21720, 16'd39846, 16'd18456, 16'd39240, 16'd3477, 16'd56345, 16'd38631});
	test_expansion(128'h447ae4758050545da92b6b4c8f838e5d, {16'd12633, 16'd15505, 16'd48384, 16'd33922, 16'd51265, 16'd5516, 16'd10641, 16'd49450, 16'd38652, 16'd59631, 16'd9994, 16'd49922, 16'd57553, 16'd45937, 16'd1168, 16'd61680, 16'd50515, 16'd64176, 16'd57857, 16'd33661, 16'd1749, 16'd10634, 16'd51842, 16'd9723, 16'd23721, 16'd44515});
	test_expansion(128'h3d79568cdb5ae64330167c20552f7489, {16'd37167, 16'd33037, 16'd21049, 16'd11238, 16'd36997, 16'd609, 16'd57559, 16'd42383, 16'd25442, 16'd59079, 16'd20735, 16'd15935, 16'd65011, 16'd53074, 16'd8771, 16'd63459, 16'd46147, 16'd37793, 16'd61273, 16'd57003, 16'd36613, 16'd26226, 16'd54866, 16'd54301, 16'd13457, 16'd56647});
	test_expansion(128'hb03ad70d65f4f79a8930004534e2daf9, {16'd22413, 16'd44133, 16'd54080, 16'd63031, 16'd63722, 16'd39770, 16'd62915, 16'd58834, 16'd35707, 16'd18363, 16'd20980, 16'd26500, 16'd60929, 16'd60376, 16'd7965, 16'd5251, 16'd4445, 16'd43938, 16'd55114, 16'd51285, 16'd12640, 16'd1224, 16'd25832, 16'd19513, 16'd9513, 16'd33803});
	test_expansion(128'hf214a325e4eef3083e54be2b3fe50a6e, {16'd7002, 16'd28978, 16'd34968, 16'd42614, 16'd31402, 16'd3319, 16'd65344, 16'd471, 16'd13425, 16'd5764, 16'd29419, 16'd46390, 16'd9845, 16'd60774, 16'd35803, 16'd45755, 16'd64576, 16'd5585, 16'd45074, 16'd47265, 16'd36123, 16'd26439, 16'd61942, 16'd48606, 16'd28790, 16'd11275});
	test_expansion(128'h834ef9f893a36c5011ee6002104f889c, {16'd8697, 16'd55715, 16'd34433, 16'd34651, 16'd59230, 16'd65136, 16'd22133, 16'd40025, 16'd11948, 16'd16852, 16'd16345, 16'd39394, 16'd50815, 16'd47837, 16'd58717, 16'd9220, 16'd20522, 16'd43789, 16'd61414, 16'd32024, 16'd12099, 16'd59732, 16'd32683, 16'd31601, 16'd26698, 16'd42503});
	test_expansion(128'h4773ba44e9ee3598b8ae8b45bc9cba68, {16'd48629, 16'd58478, 16'd27510, 16'd57462, 16'd48666, 16'd17820, 16'd38316, 16'd41549, 16'd64737, 16'd56096, 16'd12338, 16'd17474, 16'd29830, 16'd30990, 16'd12894, 16'd43512, 16'd25609, 16'd18636, 16'd44321, 16'd21913, 16'd19952, 16'd49974, 16'd29515, 16'd43073, 16'd16091, 16'd8297});
	test_expansion(128'h5abc9d73dd9abc14a7690f29f25750ff, {16'd34258, 16'd5981, 16'd38455, 16'd55785, 16'd57897, 16'd34018, 16'd55864, 16'd29406, 16'd57903, 16'd1842, 16'd47512, 16'd48411, 16'd28111, 16'd8556, 16'd34690, 16'd8894, 16'd26807, 16'd22518, 16'd58763, 16'd54226, 16'd61403, 16'd51283, 16'd33489, 16'd16863, 16'd64608, 16'd21175});
	test_expansion(128'h8d24e13b622511c37a6ba2698bbf5452, {16'd15234, 16'd27976, 16'd9427, 16'd14225, 16'd59893, 16'd6237, 16'd28556, 16'd11725, 16'd13162, 16'd29097, 16'd32788, 16'd14613, 16'd59568, 16'd37545, 16'd47180, 16'd31711, 16'd50344, 16'd60056, 16'd11110, 16'd30720, 16'd1187, 16'd43525, 16'd45401, 16'd438, 16'd932, 16'd45673});
	test_expansion(128'h4d5abae0200cf05eecd6ff8847a31b8b, {16'd51137, 16'd42689, 16'd63982, 16'd25464, 16'd2140, 16'd59496, 16'd29649, 16'd54707, 16'd43378, 16'd39179, 16'd47922, 16'd21719, 16'd34363, 16'd23796, 16'd5246, 16'd41158, 16'd52525, 16'd4126, 16'd48134, 16'd12227, 16'd57313, 16'd23464, 16'd59874, 16'd5657, 16'd25122, 16'd55993});
	test_expansion(128'h5bf9b5e364270113ca8fdf81949d4568, {16'd55635, 16'd34845, 16'd57513, 16'd35886, 16'd21339, 16'd27165, 16'd2213, 16'd47766, 16'd29726, 16'd52011, 16'd11664, 16'd27668, 16'd55588, 16'd17410, 16'd39470, 16'd13285, 16'd19308, 16'd48852, 16'd14152, 16'd55311, 16'd2071, 16'd35064, 16'd39270, 16'd4122, 16'd16995, 16'd3744});
	test_expansion(128'h3b29e7e1dc65508ac3f7c57a27e10a01, {16'd26584, 16'd43751, 16'd13000, 16'd40259, 16'd1351, 16'd42440, 16'd16973, 16'd15370, 16'd33241, 16'd48597, 16'd40357, 16'd27640, 16'd26646, 16'd9211, 16'd7215, 16'd61490, 16'd61719, 16'd23763, 16'd10488, 16'd22952, 16'd32077, 16'd47956, 16'd19298, 16'd64458, 16'd26296, 16'd7670});
	test_expansion(128'hbe900c4ce8c830650851df8712a19485, {16'd2558, 16'd856, 16'd57313, 16'd51372, 16'd58621, 16'd12519, 16'd58912, 16'd28921, 16'd36374, 16'd26618, 16'd36510, 16'd64243, 16'd21320, 16'd15630, 16'd52631, 16'd119, 16'd22093, 16'd14835, 16'd10855, 16'd23290, 16'd25312, 16'd63583, 16'd24725, 16'd29173, 16'd3501, 16'd27434});
	test_expansion(128'hec7410c20783677b025e00bc8ed1ec8d, {16'd5954, 16'd50770, 16'd25867, 16'd8645, 16'd57133, 16'd26853, 16'd28253, 16'd58876, 16'd39517, 16'd2685, 16'd45783, 16'd33040, 16'd27071, 16'd65340, 16'd12010, 16'd62596, 16'd30539, 16'd6401, 16'd35745, 16'd58614, 16'd9149, 16'd51637, 16'd57273, 16'd3759, 16'd11544, 16'd34305});
	test_expansion(128'h7b09e829dde33950a75abf72a96352bf, {16'd30406, 16'd8168, 16'd31099, 16'd47673, 16'd44375, 16'd46652, 16'd54341, 16'd11446, 16'd5602, 16'd31456, 16'd41783, 16'd63041, 16'd50831, 16'd50947, 16'd8410, 16'd55931, 16'd22557, 16'd34591, 16'd3592, 16'd30165, 16'd19976, 16'd53367, 16'd48360, 16'd45619, 16'd63132, 16'd53275});
	test_expansion(128'h80b13bf8bba7bbee1c6ff491fafe596c, {16'd12843, 16'd51903, 16'd54580, 16'd7007, 16'd503, 16'd9613, 16'd31060, 16'd9221, 16'd25049, 16'd29683, 16'd61488, 16'd62489, 16'd45540, 16'd31853, 16'd49699, 16'd35021, 16'd16608, 16'd28204, 16'd27865, 16'd3313, 16'd22151, 16'd32731, 16'd28551, 16'd10532, 16'd43443, 16'd20033});
	test_expansion(128'h1f6eab21d1823202f17468391dcbf073, {16'd35099, 16'd60012, 16'd41194, 16'd11112, 16'd3052, 16'd20046, 16'd8604, 16'd8999, 16'd16474, 16'd49038, 16'd25882, 16'd8417, 16'd41745, 16'd30445, 16'd2874, 16'd12745, 16'd41754, 16'd30600, 16'd60561, 16'd57463, 16'd44873, 16'd38740, 16'd46709, 16'd31040, 16'd4368, 16'd7443});
	test_expansion(128'he225b82ee1c5594cf53d2265331412aa, {16'd27228, 16'd53511, 16'd45414, 16'd38435, 16'd32380, 16'd60807, 16'd29529, 16'd13186, 16'd7639, 16'd40485, 16'd22077, 16'd13071, 16'd64001, 16'd55723, 16'd40679, 16'd30006, 16'd29757, 16'd43545, 16'd28661, 16'd47524, 16'd45513, 16'd12904, 16'd38280, 16'd13133, 16'd14557, 16'd31181});
	test_expansion(128'h51aa305a2e43b5cc7f9dcdf075853cd3, {16'd21097, 16'd34791, 16'd55406, 16'd60336, 16'd51220, 16'd9494, 16'd3576, 16'd7969, 16'd42856, 16'd4725, 16'd60332, 16'd48826, 16'd52835, 16'd46454, 16'd26751, 16'd56214, 16'd6529, 16'd46696, 16'd14982, 16'd19084, 16'd837, 16'd30467, 16'd20160, 16'd63917, 16'd9865, 16'd164});
	test_expansion(128'hd5cec66e5db535a42d110f7134c0f851, {16'd56086, 16'd54789, 16'd63634, 16'd54156, 16'd59653, 16'd50055, 16'd36127, 16'd27676, 16'd61848, 16'd10535, 16'd65400, 16'd62433, 16'd63033, 16'd5544, 16'd29278, 16'd19859, 16'd20206, 16'd54415, 16'd1383, 16'd36107, 16'd58247, 16'd40010, 16'd46776, 16'd22938, 16'd32599, 16'd27220});
	test_expansion(128'hf59c357d7bca8dbf0a26751129822d9f, {16'd14966, 16'd38696, 16'd56872, 16'd56038, 16'd46696, 16'd61991, 16'd14117, 16'd45884, 16'd20168, 16'd45476, 16'd18070, 16'd22662, 16'd14712, 16'd19673, 16'd38130, 16'd24249, 16'd11580, 16'd64600, 16'd64633, 16'd20161, 16'd46576, 16'd42522, 16'd11824, 16'd19606, 16'd4662, 16'd60314});
	test_expansion(128'ha792085e9034425e14cbfc1b749f037e, {16'd41303, 16'd4752, 16'd30362, 16'd27073, 16'd58398, 16'd45818, 16'd63490, 16'd48385, 16'd28414, 16'd35331, 16'd45516, 16'd58939, 16'd50245, 16'd49042, 16'd22944, 16'd56204, 16'd56619, 16'd33547, 16'd28131, 16'd27196, 16'd57827, 16'd29871, 16'd2133, 16'd35870, 16'd47257, 16'd29574});
	test_expansion(128'hf875fa5e07adc4b5eb44898ba1f1e813, {16'd19479, 16'd2880, 16'd33772, 16'd62530, 16'd46639, 16'd222, 16'd41289, 16'd7383, 16'd3392, 16'd1586, 16'd2392, 16'd30953, 16'd7064, 16'd52559, 16'd26067, 16'd36705, 16'd6677, 16'd28364, 16'd23326, 16'd33161, 16'd23102, 16'd19798, 16'd59672, 16'd33406, 16'd34257, 16'd30502});
	test_expansion(128'h317e2d085246ac246b9837f2dabf200e, {16'd49357, 16'd24998, 16'd33014, 16'd9199, 16'd24797, 16'd45720, 16'd828, 16'd30376, 16'd14326, 16'd59350, 16'd34939, 16'd61390, 16'd26794, 16'd9159, 16'd31371, 16'd45773, 16'd23974, 16'd663, 16'd18121, 16'd31340, 16'd49122, 16'd56923, 16'd48984, 16'd17789, 16'd867, 16'd51076});
	test_expansion(128'h228c21090fd180967a92b4295e68505b, {16'd42654, 16'd26142, 16'd30078, 16'd50986, 16'd48959, 16'd19373, 16'd17621, 16'd13635, 16'd31593, 16'd23197, 16'd29506, 16'd49733, 16'd8296, 16'd11954, 16'd39629, 16'd34772, 16'd64019, 16'd3135, 16'd38614, 16'd50228, 16'd51857, 16'd46215, 16'd42615, 16'd63275, 16'd36338, 16'd48197});
	test_expansion(128'hb990aff68cebd440f1689da2175e0513, {16'd54042, 16'd44852, 16'd9602, 16'd13525, 16'd32194, 16'd54364, 16'd37668, 16'd16, 16'd31069, 16'd29365, 16'd58909, 16'd63848, 16'd56746, 16'd26097, 16'd34609, 16'd12555, 16'd21858, 16'd56330, 16'd23462, 16'd63209, 16'd64460, 16'd20646, 16'd48231, 16'd29959, 16'd59643, 16'd33275});
	test_expansion(128'h17695e7d96222c53c4b3f843920f5251, {16'd13136, 16'd29336, 16'd11, 16'd35439, 16'd57379, 16'd7181, 16'd35476, 16'd17707, 16'd15543, 16'd39885, 16'd58289, 16'd32469, 16'd50977, 16'd42291, 16'd49882, 16'd9601, 16'd47736, 16'd2281, 16'd43115, 16'd10058, 16'd27760, 16'd58468, 16'd2853, 16'd320, 16'd48983, 16'd36589});
	test_expansion(128'h40fd98fae838f70e40286b8e111b8894, {16'd42678, 16'd46711, 16'd46240, 16'd36402, 16'd30885, 16'd40826, 16'd55486, 16'd25538, 16'd29896, 16'd53573, 16'd54107, 16'd59814, 16'd62815, 16'd62032, 16'd15926, 16'd5478, 16'd28517, 16'd36081, 16'd51578, 16'd32458, 16'd8870, 16'd42362, 16'd3889, 16'd22734, 16'd13793, 16'd13216});
	test_expansion(128'h8cd27af9f1563d109d59d8c6ee40b707, {16'd43860, 16'd49792, 16'd23500, 16'd11291, 16'd36136, 16'd33289, 16'd1225, 16'd23457, 16'd23387, 16'd32585, 16'd42538, 16'd41842, 16'd20741, 16'd12162, 16'd37243, 16'd32023, 16'd21623, 16'd47873, 16'd44358, 16'd18663, 16'd27071, 16'd42570, 16'd26958, 16'd382, 16'd15429, 16'd30803});
	test_expansion(128'h3b6084a3b0fb7d57693a197d713e5001, {16'd63831, 16'd56692, 16'd19242, 16'd30454, 16'd23182, 16'd63910, 16'd65033, 16'd3231, 16'd26087, 16'd12642, 16'd45112, 16'd30515, 16'd57512, 16'd58534, 16'd328, 16'd55071, 16'd27330, 16'd46173, 16'd25170, 16'd11891, 16'd57645, 16'd54958, 16'd38021, 16'd35015, 16'd17646, 16'd27570});
	test_expansion(128'h04233f79ca6dd643d6e63ab549189238, {16'd1294, 16'd50621, 16'd62827, 16'd6249, 16'd22505, 16'd34847, 16'd17119, 16'd40166, 16'd36103, 16'd9632, 16'd51403, 16'd22131, 16'd58126, 16'd51306, 16'd26773, 16'd59235, 16'd59128, 16'd63162, 16'd29028, 16'd1342, 16'd27210, 16'd9570, 16'd26934, 16'd60, 16'd60114, 16'd57430});
	test_expansion(128'hd3e643a380b240e38db35147ad77a519, {16'd37267, 16'd41717, 16'd32446, 16'd9136, 16'd26361, 16'd3765, 16'd9571, 16'd4010, 16'd60797, 16'd46958, 16'd6276, 16'd57768, 16'd57420, 16'd32861, 16'd58431, 16'd6587, 16'd32594, 16'd42625, 16'd40955, 16'd33207, 16'd62857, 16'd14191, 16'd31248, 16'd18940, 16'd23630, 16'd63319});
	test_expansion(128'hbe3ef6be8be07896856b6e49930c276c, {16'd28714, 16'd63194, 16'd23488, 16'd13592, 16'd28548, 16'd14274, 16'd53677, 16'd10535, 16'd19708, 16'd50860, 16'd9694, 16'd48370, 16'd12447, 16'd44081, 16'd22048, 16'd7331, 16'd61149, 16'd21639, 16'd558, 16'd57419, 16'd32858, 16'd3865, 16'd11615, 16'd64869, 16'd25998, 16'd34742});
	test_expansion(128'he0657a2a88a03a3d962e93be00c8693f, {16'd49546, 16'd42934, 16'd1579, 16'd24612, 16'd3938, 16'd22511, 16'd12425, 16'd42793, 16'd51538, 16'd57475, 16'd38194, 16'd47934, 16'd28448, 16'd42745, 16'd2510, 16'd57776, 16'd21913, 16'd39437, 16'd29405, 16'd10829, 16'd30973, 16'd44771, 16'd52995, 16'd7508, 16'd62722, 16'd40341});
	test_expansion(128'ha4deaa2e7388d0ad0d1b5bc63cca7191, {16'd36878, 16'd21412, 16'd15502, 16'd61450, 16'd15795, 16'd59884, 16'd34620, 16'd62901, 16'd12453, 16'd52286, 16'd16327, 16'd45670, 16'd17535, 16'd50977, 16'd1400, 16'd3082, 16'd28011, 16'd55547, 16'd27147, 16'd47196, 16'd984, 16'd40902, 16'd22292, 16'd50438, 16'd24062, 16'd31333});
	test_expansion(128'h1acc873eeb3899226599623b9b2d5b58, {16'd41486, 16'd20591, 16'd8656, 16'd54606, 16'd29527, 16'd13426, 16'd20720, 16'd41579, 16'd46071, 16'd37524, 16'd4187, 16'd6541, 16'd43023, 16'd49577, 16'd943, 16'd50350, 16'd19122, 16'd56659, 16'd51476, 16'd53618, 16'd56024, 16'd18006, 16'd20975, 16'd20895, 16'd30358, 16'd61453});
	test_expansion(128'h7a0cc6961bfa84db02c94e6fb84ddd85, {16'd11712, 16'd6530, 16'd60541, 16'd35381, 16'd25243, 16'd36824, 16'd18032, 16'd62224, 16'd36188, 16'd3845, 16'd50642, 16'd56004, 16'd44208, 16'd64535, 16'd14965, 16'd20547, 16'd49169, 16'd2857, 16'd22398, 16'd46435, 16'd54834, 16'd46437, 16'd16173, 16'd23957, 16'd13305, 16'd27589});
	test_expansion(128'h4c2133f0840f676fb82d4505bfa54301, {16'd30318, 16'd49283, 16'd58918, 16'd43714, 16'd6420, 16'd8954, 16'd41864, 16'd29716, 16'd62562, 16'd19811, 16'd40803, 16'd29812, 16'd60239, 16'd38220, 16'd474, 16'd6755, 16'd25277, 16'd58370, 16'd40207, 16'd32993, 16'd60563, 16'd20438, 16'd37094, 16'd65258, 16'd7617, 16'd41987});
	test_expansion(128'ha7ae461be738b646233cd3b6e5f0c2e5, {16'd25337, 16'd30229, 16'd63588, 16'd60433, 16'd43527, 16'd19146, 16'd5107, 16'd40905, 16'd36338, 16'd12513, 16'd37827, 16'd11428, 16'd63946, 16'd11281, 16'd22752, 16'd10238, 16'd37855, 16'd7983, 16'd45724, 16'd22024, 16'd57871, 16'd9231, 16'd19269, 16'd64015, 16'd9244, 16'd32912});
	test_expansion(128'h87c1fb7167cb4c09ca2cf00f207a5f56, {16'd25933, 16'd36616, 16'd28609, 16'd34535, 16'd49248, 16'd50433, 16'd63083, 16'd37264, 16'd11429, 16'd52458, 16'd36667, 16'd30236, 16'd12241, 16'd27479, 16'd47159, 16'd14494, 16'd6524, 16'd50673, 16'd41285, 16'd20224, 16'd13160, 16'd33778, 16'd34999, 16'd33170, 16'd36296, 16'd51554});
	test_expansion(128'h496fcfd01c1ea76f878db8d76c9d2f36, {16'd7083, 16'd25458, 16'd50320, 16'd41033, 16'd55855, 16'd30025, 16'd29404, 16'd11900, 16'd53600, 16'd8690, 16'd25335, 16'd60981, 16'd16394, 16'd2119, 16'd15263, 16'd24869, 16'd14738, 16'd34803, 16'd31966, 16'd55072, 16'd37794, 16'd56844, 16'd770, 16'd4700, 16'd39303, 16'd18337});
	test_expansion(128'h883334f52dc1c971ec7cf898beb5a4e3, {16'd24903, 16'd61312, 16'd24746, 16'd44522, 16'd59400, 16'd55830, 16'd40877, 16'd7893, 16'd28329, 16'd20447, 16'd50186, 16'd64339, 16'd38232, 16'd49446, 16'd19634, 16'd47563, 16'd53981, 16'd23131, 16'd51887, 16'd60777, 16'd39493, 16'd56804, 16'd44907, 16'd19999, 16'd1970, 16'd13335});
	test_expansion(128'hd735b735d9dc3b27223a1d606477a44a, {16'd6230, 16'd1945, 16'd28021, 16'd23361, 16'd36596, 16'd63300, 16'd28667, 16'd14132, 16'd8000, 16'd46784, 16'd38082, 16'd63257, 16'd2366, 16'd19562, 16'd62944, 16'd58662, 16'd59516, 16'd62969, 16'd64326, 16'd31574, 16'd45314, 16'd13185, 16'd29713, 16'd62947, 16'd10958, 16'd37382});
	test_expansion(128'haac26931437a605b43680ef16b90ce75, {16'd30183, 16'd24475, 16'd38254, 16'd46604, 16'd63996, 16'd29483, 16'd27130, 16'd37093, 16'd64836, 16'd14037, 16'd51640, 16'd3129, 16'd62499, 16'd9107, 16'd3464, 16'd18321, 16'd15694, 16'd43602, 16'd40288, 16'd38239, 16'd22523, 16'd36111, 16'd18008, 16'd60385, 16'd19480, 16'd39501});
	test_expansion(128'hedb8976a2be7f5ad8de6dab9c0d893a2, {16'd3743, 16'd13949, 16'd56041, 16'd7230, 16'd5050, 16'd59910, 16'd11225, 16'd46513, 16'd23549, 16'd47488, 16'd39190, 16'd50577, 16'd34509, 16'd35672, 16'd12969, 16'd26251, 16'd61006, 16'd36264, 16'd44528, 16'd9648, 16'd18688, 16'd61238, 16'd23993, 16'd3131, 16'd40204, 16'd12979});
	test_expansion(128'h6db4cae0c116700995f4bdda25d85913, {16'd55760, 16'd52143, 16'd13812, 16'd19234, 16'd15935, 16'd38869, 16'd17265, 16'd15134, 16'd15924, 16'd58395, 16'd47513, 16'd35674, 16'd1237, 16'd23937, 16'd31362, 16'd63340, 16'd31328, 16'd6588, 16'd16107, 16'd64943, 16'd9552, 16'd30241, 16'd50635, 16'd36417, 16'd38182, 16'd8595});
	test_expansion(128'h5132291781b498ab2ef12c0c58419dbb, {16'd42576, 16'd52502, 16'd59953, 16'd64027, 16'd14123, 16'd37718, 16'd23414, 16'd17286, 16'd50570, 16'd48954, 16'd54501, 16'd37335, 16'd26381, 16'd39500, 16'd60298, 16'd6444, 16'd27296, 16'd61004, 16'd20708, 16'd21272, 16'd4108, 16'd55185, 16'd4616, 16'd3934, 16'd16708, 16'd18765});
	test_expansion(128'hd2d4738c3b9375be910c88b58ab32e51, {16'd38645, 16'd19745, 16'd36826, 16'd19391, 16'd30119, 16'd24613, 16'd47372, 16'd1904, 16'd13943, 16'd32561, 16'd44483, 16'd24508, 16'd32504, 16'd40860, 16'd37974, 16'd29839, 16'd51292, 16'd45927, 16'd6668, 16'd42787, 16'd49111, 16'd5767, 16'd36846, 16'd41486, 16'd35242, 16'd51041});
	test_expansion(128'hf4b11b0bd4ca707a112033054897b4f1, {16'd61460, 16'd8968, 16'd60849, 16'd38796, 16'd57810, 16'd37645, 16'd16038, 16'd60692, 16'd49778, 16'd10289, 16'd6080, 16'd41563, 16'd43020, 16'd776, 16'd34737, 16'd10058, 16'd28846, 16'd43794, 16'd35453, 16'd44169, 16'd10283, 16'd40688, 16'd2760, 16'd42039, 16'd8000, 16'd46530});
	test_expansion(128'h4bed8f55ab434436838877e8dcb77034, {16'd37838, 16'd36203, 16'd11110, 16'd13876, 16'd24887, 16'd9290, 16'd57367, 16'd4868, 16'd31956, 16'd20748, 16'd65139, 16'd6803, 16'd55057, 16'd45777, 16'd39787, 16'd54526, 16'd11632, 16'd32669, 16'd35489, 16'd27514, 16'd11192, 16'd59581, 16'd27616, 16'd23642, 16'd21835, 16'd16720});
	test_expansion(128'hc261ce2645210dfeb1bb7584c227a0b7, {16'd18900, 16'd52916, 16'd56319, 16'd16781, 16'd9520, 16'd40824, 16'd61053, 16'd11221, 16'd37926, 16'd60547, 16'd49362, 16'd57069, 16'd14799, 16'd9096, 16'd23662, 16'd14307, 16'd33380, 16'd34383, 16'd9753, 16'd6379, 16'd14708, 16'd23996, 16'd32404, 16'd62512, 16'd40750, 16'd25631});
	test_expansion(128'h7dfa974e390a75a981abb144684be22d, {16'd26106, 16'd10602, 16'd23659, 16'd38174, 16'd32917, 16'd386, 16'd34922, 16'd26613, 16'd30868, 16'd40932, 16'd1781, 16'd42414, 16'd644, 16'd49800, 16'd50671, 16'd51361, 16'd39054, 16'd61190, 16'd35592, 16'd321, 16'd55765, 16'd13604, 16'd19701, 16'd52569, 16'd11503, 16'd62475});
	test_expansion(128'hab9d15dc06dc3777afbcc60633a455f6, {16'd57797, 16'd40238, 16'd18967, 16'd42624, 16'd64577, 16'd8326, 16'd50331, 16'd11134, 16'd25857, 16'd31094, 16'd48955, 16'd4034, 16'd13111, 16'd28576, 16'd64187, 16'd54654, 16'd47041, 16'd8705, 16'd3449, 16'd60707, 16'd18922, 16'd7887, 16'd9013, 16'd37853, 16'd63563, 16'd48944});
	test_expansion(128'hf6e6fe830e671df942fde75f8a0f32ea, {16'd6583, 16'd14710, 16'd15464, 16'd22300, 16'd43076, 16'd44262, 16'd47055, 16'd34622, 16'd59952, 16'd48453, 16'd31590, 16'd4938, 16'd36533, 16'd56367, 16'd29134, 16'd2310, 16'd11947, 16'd20725, 16'd51699, 16'd46970, 16'd44934, 16'd2802, 16'd51670, 16'd9561, 16'd9582, 16'd48414});
	test_expansion(128'hd2d3e7b8451f3528e5221545d686c3b8, {16'd14654, 16'd13152, 16'd59497, 16'd51115, 16'd33783, 16'd9240, 16'd38291, 16'd12549, 16'd43732, 16'd8411, 16'd35236, 16'd36702, 16'd63383, 16'd20769, 16'd8349, 16'd11176, 16'd50465, 16'd35236, 16'd1537, 16'd5748, 16'd21245, 16'd63012, 16'd53267, 16'd40413, 16'd34171, 16'd42796});
	test_expansion(128'h9629b4b2e5e6e004db39e3ff16b17d7c, {16'd17842, 16'd1845, 16'd23954, 16'd45380, 16'd23259, 16'd46228, 16'd64121, 16'd21551, 16'd41617, 16'd48749, 16'd49164, 16'd14390, 16'd30134, 16'd36293, 16'd30651, 16'd53944, 16'd18538, 16'd50666, 16'd53375, 16'd23623, 16'd33015, 16'd464, 16'd14059, 16'd65175, 16'd62379, 16'd3592});
	test_expansion(128'ha02384f98a0a30d56a94cee6511053cd, {16'd15236, 16'd13540, 16'd215, 16'd15069, 16'd57540, 16'd25517, 16'd59590, 16'd26107, 16'd52117, 16'd2001, 16'd35466, 16'd35569, 16'd3628, 16'd17038, 16'd51745, 16'd35884, 16'd20600, 16'd25801, 16'd22932, 16'd34619, 16'd21844, 16'd22050, 16'd26563, 16'd55186, 16'd49650, 16'd57615});
	test_expansion(128'he3550c9978e8206098b5a83295ea8cf1, {16'd50940, 16'd9060, 16'd9148, 16'd47615, 16'd9260, 16'd19924, 16'd11875, 16'd30742, 16'd29619, 16'd32758, 16'd19143, 16'd38137, 16'd18385, 16'd13052, 16'd49058, 16'd42711, 16'd41050, 16'd40320, 16'd15918, 16'd39565, 16'd112, 16'd4115, 16'd32567, 16'd42938, 16'd41565, 16'd49012});
	test_expansion(128'h050a23491af0c2d794c9b6c7c04e8c90, {16'd5834, 16'd25988, 16'd29905, 16'd53798, 16'd44167, 16'd22863, 16'd50146, 16'd18469, 16'd55729, 16'd64078, 16'd17367, 16'd17126, 16'd38363, 16'd55277, 16'd26786, 16'd60833, 16'd12143, 16'd27660, 16'd45951, 16'd27946, 16'd39103, 16'd46973, 16'd55153, 16'd32094, 16'd45014, 16'd61882});
	test_expansion(128'h6a21d1e3bdc77e3c5fd44b213b742d82, {16'd34507, 16'd52255, 16'd44990, 16'd37938, 16'd51155, 16'd31359, 16'd37484, 16'd42621, 16'd64049, 16'd58737, 16'd2714, 16'd55501, 16'd29469, 16'd61805, 16'd35317, 16'd25333, 16'd52977, 16'd48335, 16'd49651, 16'd58497, 16'd28670, 16'd25555, 16'd49146, 16'd27172, 16'd54221, 16'd44629});
	test_expansion(128'hbf424164c7917f91c04bf8362567e6c1, {16'd897, 16'd27375, 16'd29431, 16'd6133, 16'd9431, 16'd59967, 16'd64140, 16'd29757, 16'd32294, 16'd46374, 16'd18506, 16'd50201, 16'd53621, 16'd28708, 16'd14730, 16'd45275, 16'd55829, 16'd34490, 16'd6072, 16'd27545, 16'd13432, 16'd17091, 16'd46205, 16'd64549, 16'd41865, 16'd54083});
	test_expansion(128'h71206efdbed917e7e956d83bb7290c20, {16'd36867, 16'd26420, 16'd51030, 16'd38760, 16'd44572, 16'd55842, 16'd56307, 16'd16792, 16'd20789, 16'd64448, 16'd10698, 16'd24384, 16'd5735, 16'd16370, 16'd25315, 16'd40561, 16'd2940, 16'd9841, 16'd60813, 16'd3352, 16'd52798, 16'd43721, 16'd43631, 16'd31787, 16'd53423, 16'd31897});
	test_expansion(128'h0b593e40de2e7d901025e377e85e0a16, {16'd58985, 16'd48975, 16'd23944, 16'd42963, 16'd20734, 16'd64385, 16'd4437, 16'd8201, 16'd44107, 16'd2876, 16'd29333, 16'd45448, 16'd20561, 16'd36666, 16'd7712, 16'd39580, 16'd22580, 16'd16231, 16'd18528, 16'd33732, 16'd44667, 16'd16605, 16'd49739, 16'd2753, 16'd64420, 16'd21336});
	test_expansion(128'h23defd4d8e3b7b1c132f817ce6c07754, {16'd36756, 16'd42446, 16'd36343, 16'd58597, 16'd27369, 16'd8895, 16'd56333, 16'd46136, 16'd10144, 16'd15638, 16'd39644, 16'd20517, 16'd44286, 16'd8192, 16'd27921, 16'd19550, 16'd49396, 16'd30641, 16'd7018, 16'd20495, 16'd34012, 16'd43064, 16'd4916, 16'd63520, 16'd535, 16'd7227});
	test_expansion(128'hd8fd2961dcbffe8e3e79dc96fd783f2b, {16'd21604, 16'd61527, 16'd3014, 16'd42523, 16'd39559, 16'd28668, 16'd36945, 16'd44372, 16'd34229, 16'd7884, 16'd37580, 16'd32943, 16'd33831, 16'd22627, 16'd19960, 16'd50727, 16'd44500, 16'd8717, 16'd53932, 16'd1781, 16'd27057, 16'd12510, 16'd33463, 16'd4639, 16'd48846, 16'd24484});
	test_expansion(128'h861289afdc1f8f5b904862d1eff4e9ce, {16'd34343, 16'd25238, 16'd36102, 16'd41928, 16'd27815, 16'd14355, 16'd7922, 16'd42915, 16'd25161, 16'd4238, 16'd51895, 16'd65374, 16'd15107, 16'd54567, 16'd59850, 16'd35826, 16'd24147, 16'd48646, 16'd20196, 16'd42636, 16'd57808, 16'd14880, 16'd55370, 16'd40176, 16'd7279, 16'd758});
	test_expansion(128'hbb08953ad44221c371960f470dc14f68, {16'd48747, 16'd18134, 16'd52548, 16'd42818, 16'd47507, 16'd51496, 16'd7213, 16'd30491, 16'd52202, 16'd27665, 16'd39728, 16'd29763, 16'd29408, 16'd60459, 16'd32028, 16'd51732, 16'd50121, 16'd64974, 16'd2932, 16'd3416, 16'd17780, 16'd1305, 16'd56328, 16'd24810, 16'd15457, 16'd51899});
	test_expansion(128'h8674067d6abe8a294e60e8a0400233b1, {16'd51325, 16'd14622, 16'd60931, 16'd26469, 16'd34072, 16'd55684, 16'd26984, 16'd51842, 16'd48566, 16'd24295, 16'd50986, 16'd3894, 16'd46558, 16'd24710, 16'd36073, 16'd53417, 16'd37478, 16'd17407, 16'd39812, 16'd41582, 16'd51500, 16'd26074, 16'd9083, 16'd56169, 16'd60257, 16'd19273});
	test_expansion(128'h293f113355cba4a39d75d2e31b7e96a8, {16'd26353, 16'd39429, 16'd57272, 16'd59562, 16'd11869, 16'd48248, 16'd46882, 16'd43256, 16'd2750, 16'd43277, 16'd6497, 16'd17361, 16'd35986, 16'd65341, 16'd17862, 16'd49702, 16'd2342, 16'd58473, 16'd53191, 16'd47625, 16'd30996, 16'd55566, 16'd61356, 16'd24997, 16'd17561, 16'd169});
	test_expansion(128'heab0b095ec919d4e11cda77d75264333, {16'd22410, 16'd49727, 16'd43291, 16'd61095, 16'd49009, 16'd36093, 16'd38864, 16'd1913, 16'd44644, 16'd37877, 16'd21774, 16'd12382, 16'd47711, 16'd56872, 16'd12008, 16'd5932, 16'd29185, 16'd31233, 16'd26390, 16'd11383, 16'd6932, 16'd15425, 16'd1838, 16'd50423, 16'd3161, 16'd25219});
	test_expansion(128'h129b63f7c3641f369ba0b1b5229d4c9a, {16'd7376, 16'd2355, 16'd62265, 16'd37734, 16'd59939, 16'd20185, 16'd7664, 16'd40248, 16'd16930, 16'd5028, 16'd46662, 16'd4043, 16'd10791, 16'd64818, 16'd3724, 16'd52893, 16'd60801, 16'd45041, 16'd50275, 16'd21863, 16'd55523, 16'd2834, 16'd44621, 16'd59263, 16'd64838, 16'd60147});
	test_expansion(128'h1c244cbe373812712629f9260c3f3b82, {16'd4636, 16'd19485, 16'd46670, 16'd23564, 16'd32183, 16'd12867, 16'd8195, 16'd30716, 16'd53699, 16'd8705, 16'd35848, 16'd16996, 16'd54751, 16'd26401, 16'd41039, 16'd37744, 16'd57724, 16'd47594, 16'd44833, 16'd41817, 16'd25503, 16'd19840, 16'd5367, 16'd210, 16'd25499, 16'd13238});
	test_expansion(128'hc0d050cceb2ad3a86ba322b7dd0e80c3, {16'd65460, 16'd64788, 16'd8996, 16'd21345, 16'd12961, 16'd29102, 16'd21472, 16'd40624, 16'd3345, 16'd593, 16'd13722, 16'd31626, 16'd59639, 16'd2268, 16'd3789, 16'd27287, 16'd62309, 16'd2022, 16'd32722, 16'd47529, 16'd60717, 16'd39663, 16'd19251, 16'd38750, 16'd60241, 16'd13588});
	test_expansion(128'h3b0b492f36fd8a192d6184763e796bd4, {16'd28832, 16'd45612, 16'd21871, 16'd58574, 16'd37136, 16'd10158, 16'd61586, 16'd58397, 16'd42922, 16'd65092, 16'd56294, 16'd30720, 16'd17263, 16'd35624, 16'd25207, 16'd30603, 16'd9934, 16'd5954, 16'd9877, 16'd62519, 16'd50985, 16'd16695, 16'd60212, 16'd23824, 16'd5922, 16'd63565});
	test_expansion(128'h0f25f83294d7e3e14bb94e12be48dfd6, {16'd3248, 16'd52635, 16'd40688, 16'd52390, 16'd23561, 16'd60466, 16'd63672, 16'd21187, 16'd57782, 16'd12084, 16'd59125, 16'd36372, 16'd52841, 16'd42779, 16'd45552, 16'd8427, 16'd1623, 16'd60779, 16'd21424, 16'd19462, 16'd25912, 16'd33548, 16'd56999, 16'd18322, 16'd61646, 16'd21284});
	test_expansion(128'h37562b111b7bab1b591f39a1fda4d0dd, {16'd45050, 16'd15912, 16'd21903, 16'd26133, 16'd44513, 16'd9891, 16'd58617, 16'd11786, 16'd56899, 16'd33693, 16'd15499, 16'd26932, 16'd7337, 16'd8744, 16'd40170, 16'd49979, 16'd61714, 16'd38311, 16'd45869, 16'd42094, 16'd25154, 16'd31562, 16'd7825, 16'd26426, 16'd63862, 16'd40664});
	test_expansion(128'h2160119937df29f5d505f24ab44fe645, {16'd36211, 16'd56095, 16'd54587, 16'd5587, 16'd57256, 16'd21872, 16'd34983, 16'd58693, 16'd22775, 16'd19861, 16'd4622, 16'd42766, 16'd17545, 16'd40870, 16'd46827, 16'd57445, 16'd51126, 16'd64743, 16'd13357, 16'd63059, 16'd33538, 16'd54038, 16'd32639, 16'd9149, 16'd13860, 16'd9208});
	test_expansion(128'hda008f8604be7fb5c08c2d80371d8a53, {16'd5837, 16'd64764, 16'd44044, 16'd55595, 16'd17593, 16'd19958, 16'd35571, 16'd24545, 16'd47425, 16'd57782, 16'd22193, 16'd13302, 16'd51602, 16'd21761, 16'd62413, 16'd3282, 16'd46067, 16'd16517, 16'd338, 16'd63731, 16'd30570, 16'd41361, 16'd3207, 16'd30189, 16'd41712, 16'd1347});
	test_expansion(128'h29ffa55bb4decdc0598646267a693340, {16'd25418, 16'd36428, 16'd24690, 16'd2003, 16'd9563, 16'd64465, 16'd39612, 16'd14735, 16'd24154, 16'd57154, 16'd25858, 16'd32262, 16'd57693, 16'd35991, 16'd42977, 16'd63944, 16'd35186, 16'd16129, 16'd43168, 16'd40754, 16'd56003, 16'd41668, 16'd33648, 16'd14175, 16'd61522, 16'd43437});
	test_expansion(128'ha43ad0bbf43777a5c680eb1628a83144, {16'd34794, 16'd52595, 16'd28788, 16'd6137, 16'd2522, 16'd37149, 16'd18241, 16'd50667, 16'd39834, 16'd26759, 16'd40959, 16'd38331, 16'd54262, 16'd47263, 16'd58989, 16'd49550, 16'd36430, 16'd1588, 16'd22193, 16'd43204, 16'd39919, 16'd2612, 16'd17275, 16'd31211, 16'd60615, 16'd29451});
	test_expansion(128'h4aef900280120df79bfcd28fa2c791ea, {16'd8422, 16'd59432, 16'd17376, 16'd38774, 16'd27681, 16'd59402, 16'd13882, 16'd36256, 16'd50561, 16'd58703, 16'd44291, 16'd50632, 16'd15533, 16'd62308, 16'd12912, 16'd56766, 16'd53350, 16'd58476, 16'd33604, 16'd50752, 16'd726, 16'd51093, 16'd35301, 16'd3469, 16'd9640, 16'd17726});
	test_expansion(128'ha3b6733a1703b1ee3db1a7ef197964e5, {16'd16581, 16'd42620, 16'd27956, 16'd9239, 16'd18726, 16'd45741, 16'd63596, 16'd46661, 16'd9990, 16'd15379, 16'd52996, 16'd61143, 16'd54302, 16'd24678, 16'd6321, 16'd52616, 16'd1211, 16'd15031, 16'd17112, 16'd23101, 16'd7683, 16'd14474, 16'd4672, 16'd21138, 16'd29577, 16'd5244});
	test_expansion(128'h62e031047daac42379edf0b6323582ef, {16'd63781, 16'd28540, 16'd12008, 16'd51498, 16'd40285, 16'd3406, 16'd44203, 16'd60852, 16'd64274, 16'd44468, 16'd38616, 16'd12202, 16'd25934, 16'd11161, 16'd52880, 16'd869, 16'd27838, 16'd41737, 16'd45897, 16'd63966, 16'd52317, 16'd47556, 16'd21809, 16'd27701, 16'd19627, 16'd13296});
	test_expansion(128'h32841f4782c8207115a291901063202f, {16'd14654, 16'd14584, 16'd8818, 16'd29187, 16'd20401, 16'd22780, 16'd58368, 16'd37533, 16'd50246, 16'd2070, 16'd13283, 16'd47042, 16'd27197, 16'd49520, 16'd12420, 16'd18768, 16'd21314, 16'd6202, 16'd3922, 16'd12785, 16'd37666, 16'd32122, 16'd13723, 16'd51844, 16'd46250, 16'd21454});
	test_expansion(128'hb6bf427a238d1dc9ffec683a75bac926, {16'd27609, 16'd15651, 16'd36446, 16'd33766, 16'd8450, 16'd5446, 16'd61357, 16'd20147, 16'd14583, 16'd56430, 16'd58770, 16'd54560, 16'd12076, 16'd12174, 16'd42410, 16'd35023, 16'd619, 16'd24404, 16'd49391, 16'd5803, 16'd47455, 16'd36452, 16'd55245, 16'd47657, 16'd19774, 16'd19503});
	test_expansion(128'h5ced88a1c5fb8f69b24cb0adc15a8b33, {16'd21370, 16'd23472, 16'd2456, 16'd50675, 16'd6084, 16'd60832, 16'd62073, 16'd39783, 16'd11410, 16'd35519, 16'd19933, 16'd23404, 16'd24914, 16'd1936, 16'd62900, 16'd5307, 16'd55586, 16'd60043, 16'd11315, 16'd24465, 16'd47492, 16'd4108, 16'd5862, 16'd6925, 16'd19223, 16'd22259});
	test_expansion(128'he7340793e03429366f09df38cce0e406, {16'd16352, 16'd63399, 16'd61963, 16'd29616, 16'd63911, 16'd12118, 16'd59074, 16'd42733, 16'd36292, 16'd23233, 16'd28958, 16'd46060, 16'd48390, 16'd19544, 16'd23668, 16'd26455, 16'd40052, 16'd19656, 16'd52475, 16'd29989, 16'd37618, 16'd52857, 16'd35952, 16'd53702, 16'd129, 16'd43223});
	test_expansion(128'h6422bb814bad3fdc42b112e6aab2bf4e, {16'd16356, 16'd36930, 16'd49929, 16'd18155, 16'd58146, 16'd55418, 16'd58180, 16'd33446, 16'd63626, 16'd47319, 16'd26279, 16'd31742, 16'd43940, 16'd9759, 16'd43240, 16'd40524, 16'd49595, 16'd41453, 16'd13968, 16'd15732, 16'd21121, 16'd28006, 16'd51816, 16'd17205, 16'd43684, 16'd15115});
	test_expansion(128'h9f97113aee19203af3178303eff52219, {16'd28711, 16'd13381, 16'd41188, 16'd56883, 16'd54410, 16'd40321, 16'd57902, 16'd25555, 16'd1013, 16'd51824, 16'd19928, 16'd63367, 16'd34883, 16'd60806, 16'd15217, 16'd895, 16'd1923, 16'd9714, 16'd39104, 16'd2583, 16'd47495, 16'd60540, 16'd16258, 16'd58907, 16'd44595, 16'd63792});
	test_expansion(128'hf6437041a27a8b9692e77de821692bc1, {16'd50959, 16'd63666, 16'd62297, 16'd26863, 16'd52389, 16'd26885, 16'd33453, 16'd9824, 16'd20877, 16'd47689, 16'd36311, 16'd57124, 16'd15801, 16'd38977, 16'd46709, 16'd7687, 16'd37282, 16'd12724, 16'd51565, 16'd62284, 16'd56835, 16'd1430, 16'd33804, 16'd672, 16'd1618, 16'd33457});
	test_expansion(128'h16581c17c2073512b7e82729259bdebb, {16'd48173, 16'd774, 16'd42791, 16'd7818, 16'd46341, 16'd65050, 16'd43935, 16'd58952, 16'd28269, 16'd14591, 16'd10779, 16'd5736, 16'd54681, 16'd9106, 16'd28381, 16'd52809, 16'd46881, 16'd893, 16'd40326, 16'd31174, 16'd49690, 16'd25509, 16'd36420, 16'd13801, 16'd12345, 16'd10632});
	test_expansion(128'h5d96d7f6a39fa20676c7cf93df53e5a1, {16'd52036, 16'd4147, 16'd6780, 16'd31382, 16'd51334, 16'd9917, 16'd1477, 16'd58371, 16'd60435, 16'd14894, 16'd24354, 16'd57263, 16'd13083, 16'd15957, 16'd5148, 16'd52066, 16'd53733, 16'd19615, 16'd38764, 16'd58490, 16'd21870, 16'd64359, 16'd35683, 16'd64752, 16'd26240, 16'd16342});
	test_expansion(128'h9950cec8fc8a3677349a0414c40da2d9, {16'd23180, 16'd38521, 16'd28665, 16'd24570, 16'd31568, 16'd49795, 16'd12302, 16'd10565, 16'd37584, 16'd15847, 16'd53415, 16'd20923, 16'd55197, 16'd16387, 16'd47368, 16'd37636, 16'd31126, 16'd40546, 16'd10260, 16'd52345, 16'd57987, 16'd10002, 16'd54148, 16'd20929, 16'd57878, 16'd19658});
	test_expansion(128'h807c79cf94657d2321767e6478e3fce3, {16'd7880, 16'd27791, 16'd57749, 16'd65206, 16'd35951, 16'd16437, 16'd54108, 16'd42225, 16'd33347, 16'd32545, 16'd55182, 16'd58800, 16'd27294, 16'd30619, 16'd19109, 16'd27346, 16'd60635, 16'd10674, 16'd1532, 16'd62862, 16'd3445, 16'd62679, 16'd59694, 16'd11337, 16'd21782, 16'd45308});
	test_expansion(128'h7e152423ef191d90104ea2d3c03f6363, {16'd19373, 16'd23584, 16'd28762, 16'd718, 16'd54612, 16'd15142, 16'd52721, 16'd29156, 16'd30302, 16'd29613, 16'd8989, 16'd47751, 16'd23125, 16'd52566, 16'd31192, 16'd12392, 16'd26231, 16'd3419, 16'd64267, 16'd19273, 16'd54800, 16'd17981, 16'd17075, 16'd3900, 16'd23889, 16'd21261});
	test_expansion(128'h76597204579ce983e423baf115340460, {16'd5512, 16'd53131, 16'd19154, 16'd1131, 16'd31663, 16'd24169, 16'd23566, 16'd26606, 16'd3994, 16'd143, 16'd46135, 16'd40715, 16'd6144, 16'd37142, 16'd43246, 16'd17982, 16'd55559, 16'd61432, 16'd44752, 16'd45245, 16'd30543, 16'd53858, 16'd16910, 16'd26015, 16'd17158, 16'd8859});
	test_expansion(128'h9017f23a6936b1b1a8e0e65688911d73, {16'd16459, 16'd43502, 16'd50673, 16'd21188, 16'd19321, 16'd25473, 16'd32987, 16'd39578, 16'd15728, 16'd48042, 16'd45805, 16'd65181, 16'd58371, 16'd51439, 16'd64322, 16'd42559, 16'd22498, 16'd64160, 16'd29835, 16'd22876, 16'd47428, 16'd55766, 16'd30357, 16'd9392, 16'd59421, 16'd21870});
	test_expansion(128'h7e5cd700c8dfb3a9fe0caec78946fd75, {16'd2661, 16'd32637, 16'd53623, 16'd8590, 16'd43102, 16'd63833, 16'd46423, 16'd12955, 16'd1893, 16'd38169, 16'd40289, 16'd17305, 16'd24298, 16'd20434, 16'd13841, 16'd16767, 16'd50824, 16'd37736, 16'd40382, 16'd49832, 16'd57494, 16'd45587, 16'd12986, 16'd50810, 16'd36830, 16'd41352});
	test_expansion(128'hbaef23e89e1121582fb63a3b71dcbcfa, {16'd9415, 16'd37418, 16'd3994, 16'd26941, 16'd56942, 16'd53489, 16'd65369, 16'd10375, 16'd40950, 16'd14617, 16'd15981, 16'd30902, 16'd13566, 16'd48012, 16'd4746, 16'd17803, 16'd40678, 16'd49591, 16'd24282, 16'd61828, 16'd48716, 16'd18321, 16'd59868, 16'd55032, 16'd37118, 16'd44205});
	test_expansion(128'hdbb643206e1cdd1eb910c8daca7d4373, {16'd11829, 16'd279, 16'd38095, 16'd47838, 16'd49782, 16'd18539, 16'd27529, 16'd34149, 16'd28930, 16'd42508, 16'd56541, 16'd2844, 16'd33283, 16'd7861, 16'd44996, 16'd44683, 16'd56559, 16'd53747, 16'd2536, 16'd64552, 16'd24675, 16'd15431, 16'd50222, 16'd31142, 16'd20111, 16'd49892});
	test_expansion(128'ha13f1003cebbd611bd191daff3d62541, {16'd25333, 16'd4711, 16'd15105, 16'd6408, 16'd55084, 16'd24404, 16'd39591, 16'd60250, 16'd21364, 16'd31577, 16'd27331, 16'd60395, 16'd39034, 16'd23915, 16'd18561, 16'd35970, 16'd3508, 16'd44902, 16'd28934, 16'd48655, 16'd9839, 16'd25208, 16'd4364, 16'd3557, 16'd56290, 16'd7583});
	test_expansion(128'h396723f2507467a5d52df70e47f0aea3, {16'd48891, 16'd57373, 16'd42144, 16'd23785, 16'd50857, 16'd25571, 16'd11569, 16'd21948, 16'd458, 16'd2334, 16'd2701, 16'd7916, 16'd12788, 16'd27647, 16'd56546, 16'd631, 16'd18753, 16'd22954, 16'd54967, 16'd54044, 16'd64311, 16'd63731, 16'd37934, 16'd2953, 16'd49697, 16'd62869});
	test_expansion(128'h5058be1fcccaeb8c42c2eb4744553dc1, {16'd49715, 16'd6771, 16'd45577, 16'd28494, 16'd60088, 16'd28600, 16'd40493, 16'd53611, 16'd44914, 16'd17937, 16'd34257, 16'd17268, 16'd7436, 16'd27540, 16'd32830, 16'd8468, 16'd38659, 16'd19653, 16'd29367, 16'd54846, 16'd50062, 16'd39333, 16'd40927, 16'd44178, 16'd43557, 16'd25112});
	test_expansion(128'h2a70421c0adf9f4cf5ff24f278af5e54, {16'd16154, 16'd31322, 16'd50693, 16'd51622, 16'd38272, 16'd61589, 16'd60493, 16'd19516, 16'd60309, 16'd35836, 16'd62610, 16'd38291, 16'd5554, 16'd52136, 16'd48294, 16'd37850, 16'd10639, 16'd14937, 16'd30387, 16'd1146, 16'd62096, 16'd52629, 16'd10320, 16'd13993, 16'd56276, 16'd54187});
	test_expansion(128'hb8b8b2e347d1b0e58f95218e3bd6c8ae, {16'd6602, 16'd6636, 16'd4041, 16'd23399, 16'd27595, 16'd1445, 16'd47925, 16'd22591, 16'd19102, 16'd44753, 16'd37080, 16'd39224, 16'd5306, 16'd29648, 16'd21046, 16'd59164, 16'd28519, 16'd34764, 16'd20639, 16'd50089, 16'd43691, 16'd62224, 16'd30063, 16'd6816, 16'd18173, 16'd1928});
	test_expansion(128'h447fd0c4ff38f217b0a4042880a9e3a5, {16'd32984, 16'd18258, 16'd45492, 16'd37164, 16'd36293, 16'd30112, 16'd33681, 16'd29424, 16'd22286, 16'd19569, 16'd29607, 16'd64437, 16'd20619, 16'd36711, 16'd63959, 16'd59144, 16'd7958, 16'd27761, 16'd61412, 16'd20178, 16'd40073, 16'd56481, 16'd33503, 16'd18291, 16'd50073, 16'd33107});
	test_expansion(128'hbca9f2e33dbe05b7317cf5bd1698aa6d, {16'd65434, 16'd48534, 16'd19588, 16'd857, 16'd8526, 16'd46779, 16'd55401, 16'd54427, 16'd29366, 16'd35920, 16'd35182, 16'd55770, 16'd47359, 16'd12086, 16'd61680, 16'd43616, 16'd13658, 16'd24310, 16'd57884, 16'd63384, 16'd31786, 16'd61385, 16'd12893, 16'd57155, 16'd2283, 16'd25429});
	test_expansion(128'h4816cc1135a9746cc6ec9fb8f4d59f9d, {16'd1216, 16'd19943, 16'd40654, 16'd33261, 16'd54500, 16'd32816, 16'd46442, 16'd53737, 16'd39869, 16'd45580, 16'd57788, 16'd39481, 16'd64819, 16'd9499, 16'd38512, 16'd19409, 16'd21193, 16'd34514, 16'd30036, 16'd4019, 16'd8880, 16'd49841, 16'd42122, 16'd65455, 16'd49805, 16'd32878});
	test_expansion(128'h9701485d4e9f3aa61dae2fee01eb3443, {16'd59921, 16'd22381, 16'd2707, 16'd29574, 16'd1463, 16'd56075, 16'd12208, 16'd39738, 16'd8677, 16'd32003, 16'd35866, 16'd54751, 16'd3305, 16'd23933, 16'd4575, 16'd979, 16'd257, 16'd38699, 16'd7366, 16'd51052, 16'd49934, 16'd49210, 16'd15468, 16'd56808, 16'd18468, 16'd37628});
	test_expansion(128'he69957d51072fa252efb4a38fd19a107, {16'd31545, 16'd53647, 16'd27400, 16'd46555, 16'd30539, 16'd12066, 16'd43329, 16'd19681, 16'd53856, 16'd41234, 16'd1970, 16'd8057, 16'd6199, 16'd22276, 16'd21742, 16'd11618, 16'd1828, 16'd11854, 16'd24857, 16'd16774, 16'd65049, 16'd46834, 16'd16478, 16'd29507, 16'd39439, 16'd14355});
	test_expansion(128'he67f22abc8d9da49a6a635090745aa28, {16'd58706, 16'd6109, 16'd35151, 16'd16542, 16'd51648, 16'd587, 16'd33770, 16'd27646, 16'd15010, 16'd45383, 16'd58400, 16'd1337, 16'd50338, 16'd27225, 16'd5045, 16'd23105, 16'd11125, 16'd47188, 16'd19755, 16'd14218, 16'd58092, 16'd20472, 16'd35400, 16'd13450, 16'd17443, 16'd1993});
	test_expansion(128'h5b6b82dd19f1911f305ae4ccae21ba15, {16'd23338, 16'd22598, 16'd5028, 16'd2068, 16'd22324, 16'd63059, 16'd48681, 16'd47595, 16'd21122, 16'd48781, 16'd40980, 16'd6398, 16'd41905, 16'd3915, 16'd38241, 16'd49589, 16'd13298, 16'd52726, 16'd56565, 16'd20017, 16'd51001, 16'd28703, 16'd62907, 16'd12183, 16'd30556, 16'd32926});
	test_expansion(128'h820cf437613be3460e986ec0bfff9605, {16'd39701, 16'd33482, 16'd13008, 16'd22528, 16'd41500, 16'd63069, 16'd44278, 16'd58416, 16'd29762, 16'd34584, 16'd22779, 16'd19565, 16'd35586, 16'd13026, 16'd44091, 16'd18141, 16'd21762, 16'd18232, 16'd12274, 16'd47892, 16'd9382, 16'd52606, 16'd28442, 16'd6819, 16'd31046, 16'd34515});
	test_expansion(128'h413a8cc77ece23d5490f9f3e6d9095f7, {16'd5124, 16'd54797, 16'd8971, 16'd27120, 16'd44422, 16'd61949, 16'd43222, 16'd47867, 16'd14626, 16'd61888, 16'd44614, 16'd41169, 16'd8204, 16'd64508, 16'd27249, 16'd471, 16'd58819, 16'd1846, 16'd4597, 16'd49672, 16'd39981, 16'd16023, 16'd55199, 16'd23920, 16'd30041, 16'd42527});
	test_expansion(128'ha5983109404a4cf318029ed9cc9d510c, {16'd18637, 16'd50508, 16'd3203, 16'd2242, 16'd50938, 16'd28615, 16'd7380, 16'd36075, 16'd25025, 16'd16760, 16'd10906, 16'd37139, 16'd2577, 16'd40076, 16'd48189, 16'd7016, 16'd14414, 16'd37006, 16'd18553, 16'd49882, 16'd28032, 16'd46878, 16'd18359, 16'd65240, 16'd30729, 16'd62398});
	test_expansion(128'hcb44ce1f904dccc2f32c5a2fba70546a, {16'd55537, 16'd23825, 16'd23022, 16'd58798, 16'd58387, 16'd15194, 16'd21015, 16'd22282, 16'd47567, 16'd36874, 16'd58084, 16'd13191, 16'd51078, 16'd1849, 16'd37897, 16'd18005, 16'd26438, 16'd39045, 16'd20781, 16'd24599, 16'd19147, 16'd18928, 16'd8245, 16'd28649, 16'd51067, 16'd38957});
	test_expansion(128'he653af7f6cea7ad699a50f4aab79b401, {16'd34266, 16'd60903, 16'd9945, 16'd6057, 16'd869, 16'd42166, 16'd5453, 16'd18947, 16'd30306, 16'd47220, 16'd660, 16'd46173, 16'd60389, 16'd52499, 16'd10608, 16'd45754, 16'd8227, 16'd45113, 16'd19138, 16'd65319, 16'd24857, 16'd58654, 16'd52098, 16'd9091, 16'd9913, 16'd63736});
	test_expansion(128'h6fd8bd3671ef48977e6edd2e1b9e9682, {16'd35068, 16'd30015, 16'd11445, 16'd50573, 16'd30903, 16'd23575, 16'd51270, 16'd51272, 16'd18152, 16'd15207, 16'd28150, 16'd26963, 16'd17178, 16'd59784, 16'd48020, 16'd9131, 16'd45014, 16'd63399, 16'd10185, 16'd58845, 16'd32987, 16'd44619, 16'd23368, 16'd27774, 16'd24351, 16'd7063});
	test_expansion(128'hcd78cc86c43fad5734011c1d74707c02, {16'd3799, 16'd61068, 16'd25849, 16'd38898, 16'd29553, 16'd64648, 16'd36075, 16'd7101, 16'd24402, 16'd19497, 16'd59644, 16'd62863, 16'd56783, 16'd29536, 16'd28758, 16'd28858, 16'd18485, 16'd4768, 16'd20748, 16'd55490, 16'd43754, 16'd8823, 16'd38517, 16'd525, 16'd28117, 16'd4500});
	test_expansion(128'h19712e58f34a3a7a47efc4e7fcf96c20, {16'd65400, 16'd51016, 16'd47005, 16'd12713, 16'd39234, 16'd61511, 16'd43284, 16'd48286, 16'd63598, 16'd23345, 16'd16876, 16'd9565, 16'd16872, 16'd9625, 16'd20227, 16'd26430, 16'd54665, 16'd11328, 16'd8632, 16'd52639, 16'd16651, 16'd6141, 16'd42867, 16'd10731, 16'd18190, 16'd63476});
	test_expansion(128'h09358105fb75c3ce1098423f4317465f, {16'd23751, 16'd11787, 16'd13688, 16'd20164, 16'd1012, 16'd2417, 16'd42526, 16'd24723, 16'd6162, 16'd64475, 16'd21219, 16'd27759, 16'd41125, 16'd61418, 16'd44557, 16'd20893, 16'd13629, 16'd5882, 16'd7501, 16'd63338, 16'd55909, 16'd1187, 16'd40111, 16'd1381, 16'd35670, 16'd47611});
	test_expansion(128'h5c48c6f98d71eb007a6197fba97c9b06, {16'd18086, 16'd30821, 16'd46640, 16'd29892, 16'd33039, 16'd60829, 16'd11543, 16'd52453, 16'd28091, 16'd34559, 16'd34266, 16'd11983, 16'd36856, 16'd50701, 16'd26880, 16'd31505, 16'd25553, 16'd25696, 16'd15476, 16'd7486, 16'd59866, 16'd45289, 16'd25008, 16'd17371, 16'd40257, 16'd56224});
	test_expansion(128'h28dc8de35fbddb6ddb48bf3f9491c6ea, {16'd11146, 16'd4520, 16'd39678, 16'd3104, 16'd34533, 16'd6040, 16'd42154, 16'd59978, 16'd25413, 16'd32160, 16'd38945, 16'd15510, 16'd58923, 16'd4805, 16'd38978, 16'd60507, 16'd5767, 16'd28236, 16'd55059, 16'd55725, 16'd55386, 16'd44595, 16'd36460, 16'd16286, 16'd53819, 16'd62394});
	test_expansion(128'hdf6d5af2942f0026ba7612613c72cfbd, {16'd26542, 16'd8463, 16'd12721, 16'd62168, 16'd31275, 16'd14376, 16'd16086, 16'd60145, 16'd60676, 16'd47666, 16'd44864, 16'd61840, 16'd38270, 16'd34471, 16'd58605, 16'd31366, 16'd3640, 16'd59907, 16'd9003, 16'd59319, 16'd28014, 16'd43506, 16'd30796, 16'd44707, 16'd37968, 16'd40306});
	test_expansion(128'h115fd1a24d919358b7bbd5d59485a2bc, {16'd20389, 16'd55031, 16'd49736, 16'd62055, 16'd30788, 16'd46273, 16'd23920, 16'd57741, 16'd35233, 16'd44521, 16'd44101, 16'd55227, 16'd5534, 16'd56134, 16'd39092, 16'd29784, 16'd19855, 16'd7494, 16'd37105, 16'd41357, 16'd36895, 16'd10622, 16'd46947, 16'd16467, 16'd26135, 16'd9546});
	test_expansion(128'hd1de4183a429499b5c24455d06dfbc76, {16'd1982, 16'd34022, 16'd35987, 16'd63259, 16'd42509, 16'd52786, 16'd61145, 16'd41841, 16'd25228, 16'd10924, 16'd11650, 16'd15948, 16'd31603, 16'd3847, 16'd49439, 16'd13197, 16'd12669, 16'd62636, 16'd5272, 16'd44740, 16'd44112, 16'd61018, 16'd43088, 16'd30608, 16'd27001, 16'd34654});
	test_expansion(128'h43494a08afd49e283523d2a22032d3eb, {16'd31082, 16'd27421, 16'd10867, 16'd36635, 16'd27721, 16'd34107, 16'd39004, 16'd10158, 16'd37335, 16'd34980, 16'd50800, 16'd23106, 16'd37268, 16'd56287, 16'd46895, 16'd9997, 16'd51603, 16'd15855, 16'd56792, 16'd46334, 16'd60120, 16'd60106, 16'd51786, 16'd47427, 16'd49482, 16'd44242});
	test_expansion(128'hce29fe594f6b1f66560bb63206865fa1, {16'd44801, 16'd37730, 16'd8424, 16'd63524, 16'd55117, 16'd47786, 16'd45900, 16'd48224, 16'd44629, 16'd8944, 16'd10502, 16'd26581, 16'd48811, 16'd28967, 16'd58317, 16'd1820, 16'd5746, 16'd17069, 16'd13593, 16'd12909, 16'd43633, 16'd35913, 16'd7219, 16'd52155, 16'd52792, 16'd37321});
	test_expansion(128'h17636e65f66ce8e09da1a3b762c89990, {16'd32540, 16'd47851, 16'd46687, 16'd61168, 16'd49007, 16'd37370, 16'd32364, 16'd26103, 16'd56654, 16'd3215, 16'd57413, 16'd56982, 16'd62080, 16'd15387, 16'd21706, 16'd46355, 16'd34595, 16'd36971, 16'd55028, 16'd28575, 16'd28832, 16'd59533, 16'd35605, 16'd41459, 16'd47258, 16'd33485});
	test_expansion(128'h1622336216935236bb535e272e7cfaeb, {16'd62589, 16'd21460, 16'd38075, 16'd30386, 16'd6738, 16'd34257, 16'd65093, 16'd7549, 16'd30481, 16'd11494, 16'd13379, 16'd44933, 16'd40096, 16'd55127, 16'd46811, 16'd6236, 16'd62748, 16'd5890, 16'd33007, 16'd9041, 16'd32661, 16'd49512, 16'd50110, 16'd62853, 16'd3714, 16'd63128});
	test_expansion(128'ha7f60eb62362dd16525012454d2130ef, {16'd22585, 16'd33475, 16'd1897, 16'd37014, 16'd13725, 16'd23008, 16'd40454, 16'd2629, 16'd57213, 16'd28441, 16'd6345, 16'd48020, 16'd9875, 16'd62410, 16'd60166, 16'd63110, 16'd48983, 16'd25395, 16'd37600, 16'd9580, 16'd47620, 16'd8336, 16'd14784, 16'd53041, 16'd51387, 16'd60690});
	test_expansion(128'h56db1c2c37441c0cf478d608127c3391, {16'd55645, 16'd37166, 16'd18583, 16'd25914, 16'd41408, 16'd2018, 16'd7682, 16'd15817, 16'd15738, 16'd10754, 16'd48415, 16'd13999, 16'd50664, 16'd62030, 16'd43916, 16'd15084, 16'd27585, 16'd53351, 16'd37316, 16'd15701, 16'd21975, 16'd14986, 16'd46888, 16'd55765, 16'd34251, 16'd28618});
	test_expansion(128'h2048e1fcb93bd622a291b90028da7788, {16'd38230, 16'd5329, 16'd10718, 16'd27909, 16'd58189, 16'd41847, 16'd9370, 16'd20495, 16'd42586, 16'd52303, 16'd46166, 16'd44767, 16'd17025, 16'd63194, 16'd41450, 16'd61648, 16'd10293, 16'd65282, 16'd51488, 16'd51689, 16'd44900, 16'd25868, 16'd2979, 16'd50548, 16'd10592, 16'd4166});
	test_expansion(128'hc670f4ababffaf45d473bbb63667a7f6, {16'd50244, 16'd44349, 16'd35672, 16'd25596, 16'd25349, 16'd23368, 16'd9073, 16'd39494, 16'd35727, 16'd21196, 16'd37013, 16'd38113, 16'd11214, 16'd40155, 16'd42241, 16'd57762, 16'd51030, 16'd18409, 16'd57471, 16'd28125, 16'd55406, 16'd12033, 16'd14728, 16'd18948, 16'd50730, 16'd53439});
	test_expansion(128'h1be88f04371a620eaf478bf45e21fb26, {16'd9639, 16'd49222, 16'd19204, 16'd7420, 16'd18224, 16'd37042, 16'd4896, 16'd47357, 16'd50863, 16'd49749, 16'd32572, 16'd27051, 16'd24627, 16'd9571, 16'd15662, 16'd5871, 16'd53161, 16'd40286, 16'd45739, 16'd36363, 16'd52035, 16'd4413, 16'd21020, 16'd2923, 16'd169, 16'd45688});
	test_expansion(128'hb35119b7ce351374dcd36e096dc3feb0, {16'd32561, 16'd4405, 16'd9419, 16'd63096, 16'd25232, 16'd58453, 16'd51104, 16'd60524, 16'd35628, 16'd33308, 16'd18630, 16'd51673, 16'd50873, 16'd53976, 16'd12747, 16'd33614, 16'd12494, 16'd37704, 16'd49838, 16'd20301, 16'd38469, 16'd3393, 16'd57045, 16'd11849, 16'd35965, 16'd48279});
	test_expansion(128'hcdadf4c62bc25b55f5ae4a751a6f451d, {16'd51642, 16'd31504, 16'd23823, 16'd16345, 16'd47950, 16'd50953, 16'd30776, 16'd5569, 16'd39144, 16'd5197, 16'd6806, 16'd15823, 16'd21259, 16'd18614, 16'd15383, 16'd16929, 16'd17270, 16'd63781, 16'd44441, 16'd2200, 16'd60233, 16'd42127, 16'd36079, 16'd27710, 16'd34663, 16'd35406});
	test_expansion(128'h28d41c31b3a239f1f6df361c30795b7d, {16'd54305, 16'd36033, 16'd58935, 16'd13927, 16'd50674, 16'd65465, 16'd37550, 16'd27923, 16'd44285, 16'd23880, 16'd9659, 16'd61983, 16'd19084, 16'd63039, 16'd35063, 16'd44901, 16'd59977, 16'd32832, 16'd22430, 16'd57139, 16'd14063, 16'd20819, 16'd61019, 16'd57260, 16'd24672, 16'd9520});
	test_expansion(128'hbcc69a72618170f406c4c65ee0e73a4b, {16'd4226, 16'd60723, 16'd50305, 16'd16424, 16'd29089, 16'd22074, 16'd31801, 16'd33572, 16'd56881, 16'd3374, 16'd25620, 16'd25769, 16'd43523, 16'd1771, 16'd21615, 16'd21509, 16'd13826, 16'd27103, 16'd16434, 16'd35149, 16'd26551, 16'd48464, 16'd31877, 16'd6212, 16'd58989, 16'd57021});
	test_expansion(128'hff490984628b72f6d3c0c24ea83fa00e, {16'd48742, 16'd54600, 16'd44118, 16'd3325, 16'd5833, 16'd49790, 16'd40255, 16'd2075, 16'd2166, 16'd56047, 16'd5977, 16'd65011, 16'd5744, 16'd18668, 16'd797, 16'd37696, 16'd52643, 16'd65237, 16'd23507, 16'd37034, 16'd50301, 16'd37138, 16'd31351, 16'd61900, 16'd53512, 16'd53223});
	test_expansion(128'h3e244ba890cdc2ba7cd3c3e895eac55f, {16'd57462, 16'd52131, 16'd57937, 16'd30866, 16'd35011, 16'd15682, 16'd12898, 16'd20820, 16'd51341, 16'd57483, 16'd2973, 16'd10800, 16'd28910, 16'd14377, 16'd50139, 16'd38322, 16'd28728, 16'd37828, 16'd64941, 16'd12855, 16'd63645, 16'd51884, 16'd3181, 16'd35740, 16'd54313, 16'd5809});
	test_expansion(128'h69e0a16b3039aa6e286951418e90fbbd, {16'd53970, 16'd29897, 16'd23569, 16'd18396, 16'd59989, 16'd42009, 16'd8079, 16'd45067, 16'd49841, 16'd61684, 16'd57845, 16'd54788, 16'd2185, 16'd26548, 16'd8018, 16'd24271, 16'd49851, 16'd9858, 16'd36928, 16'd28676, 16'd64382, 16'd57949, 16'd52912, 16'd61803, 16'd13096, 16'd26055});
	test_expansion(128'hf52fe407b133abc9833c16c02a764bbe, {16'd55047, 16'd14231, 16'd35362, 16'd696, 16'd12434, 16'd26770, 16'd23997, 16'd9856, 16'd32011, 16'd55898, 16'd9500, 16'd19110, 16'd65397, 16'd38260, 16'd50898, 16'd1570, 16'd9999, 16'd37466, 16'd14974, 16'd13646, 16'd32239, 16'd36416, 16'd40731, 16'd24652, 16'd3742, 16'd22432});
	test_expansion(128'h6fdc4387e0ba7fc33209d6098d851cf5, {16'd38068, 16'd18634, 16'd37108, 16'd36333, 16'd13220, 16'd6836, 16'd65481, 16'd6574, 16'd64479, 16'd40914, 16'd7812, 16'd33934, 16'd58418, 16'd45914, 16'd32097, 16'd9627, 16'd46243, 16'd5449, 16'd48424, 16'd47671, 16'd10167, 16'd50892, 16'd5420, 16'd35620, 16'd57930, 16'd51890});
	test_expansion(128'h24072c67259a81020ca142bb8acf00a2, {16'd65384, 16'd22053, 16'd30956, 16'd47995, 16'd58492, 16'd38052, 16'd5747, 16'd59387, 16'd54954, 16'd36750, 16'd37934, 16'd57860, 16'd13388, 16'd7326, 16'd64532, 16'd3272, 16'd9434, 16'd30479, 16'd10766, 16'd615, 16'd34965, 16'd6290, 16'd2545, 16'd59118, 16'd48704, 16'd26458});
	test_expansion(128'h3078258680e3e5f7de56f67851e9e59e, {16'd20201, 16'd163, 16'd14604, 16'd9826, 16'd32291, 16'd46470, 16'd56527, 16'd32894, 16'd24900, 16'd60640, 16'd19021, 16'd54537, 16'd7155, 16'd38325, 16'd62145, 16'd5346, 16'd33080, 16'd28258, 16'd17653, 16'd27831, 16'd50729, 16'd40857, 16'd60107, 16'd47518, 16'd13576, 16'd19464});
	test_expansion(128'h733401623319d01b91a93628ee75c4d3, {16'd37250, 16'd32668, 16'd49944, 16'd11603, 16'd54886, 16'd49890, 16'd5932, 16'd5499, 16'd50584, 16'd57988, 16'd37579, 16'd34160, 16'd60185, 16'd12118, 16'd33730, 16'd18453, 16'd56310, 16'd15144, 16'd4210, 16'd24460, 16'd32290, 16'd25166, 16'd23332, 16'd685, 16'd18651, 16'd59387});
	test_expansion(128'h7cdbbe80f86438be05607fc1d05c0607, {16'd34672, 16'd41020, 16'd62320, 16'd22085, 16'd10689, 16'd21442, 16'd41432, 16'd6354, 16'd35963, 16'd25733, 16'd48634, 16'd46171, 16'd634, 16'd28698, 16'd4897, 16'd27825, 16'd7625, 16'd36165, 16'd50604, 16'd11432, 16'd1722, 16'd43726, 16'd53074, 16'd50967, 16'd58796, 16'd63336});
	test_expansion(128'h71b79f478ae1e020ad5afcf5799e90fa, {16'd9762, 16'd24470, 16'd55839, 16'd46946, 16'd51357, 16'd40073, 16'd30425, 16'd64902, 16'd49256, 16'd23227, 16'd586, 16'd41488, 16'd14155, 16'd7484, 16'd47974, 16'd65486, 16'd33115, 16'd539, 16'd36672, 16'd52022, 16'd44366, 16'd8350, 16'd50549, 16'd38609, 16'd44672, 16'd43131});
	test_expansion(128'ha69d4839e5f3e2ed5852a0b3212fcb59, {16'd33975, 16'd5363, 16'd23064, 16'd56471, 16'd7162, 16'd54804, 16'd7506, 16'd11945, 16'd20440, 16'd39002, 16'd33018, 16'd36304, 16'd36469, 16'd26922, 16'd9870, 16'd21019, 16'd45997, 16'd58394, 16'd59405, 16'd3437, 16'd819, 16'd35686, 16'd793, 16'd42161, 16'd15648, 16'd11671});
	test_expansion(128'h9efdd90983618bf47cbd8f8b7952682e, {16'd30346, 16'd40139, 16'd32754, 16'd28902, 16'd9737, 16'd25120, 16'd18049, 16'd10591, 16'd925, 16'd28693, 16'd31335, 16'd5321, 16'd55974, 16'd44753, 16'd1002, 16'd1787, 16'd27645, 16'd4339, 16'd58203, 16'd15950, 16'd6579, 16'd27068, 16'd17850, 16'd42714, 16'd14042, 16'd18870});
	test_expansion(128'h657c292f0424eb1ddaab0a4adaa9b21f, {16'd32126, 16'd57775, 16'd60159, 16'd11951, 16'd463, 16'd21895, 16'd5341, 16'd34212, 16'd18661, 16'd17626, 16'd4330, 16'd19073, 16'd34921, 16'd17266, 16'd55801, 16'd7575, 16'd28396, 16'd7133, 16'd3633, 16'd27057, 16'd35902, 16'd43276, 16'd43823, 16'd41072, 16'd44048, 16'd19405});
	test_expansion(128'h2e9ae4a3845220258df70e2a7ba050b8, {16'd57355, 16'd29924, 16'd44587, 16'd11118, 16'd58716, 16'd27620, 16'd51349, 16'd431, 16'd5703, 16'd42476, 16'd19517, 16'd2059, 16'd14111, 16'd23149, 16'd60719, 16'd15901, 16'd47635, 16'd34916, 16'd45363, 16'd54397, 16'd61776, 16'd51611, 16'd59443, 16'd48787, 16'd57176, 16'd44166});
	test_expansion(128'h6635f850b9d6b87d0214f4575366d930, {16'd29846, 16'd11027, 16'd1454, 16'd40402, 16'd61087, 16'd12868, 16'd42501, 16'd6506, 16'd31664, 16'd10655, 16'd56542, 16'd26261, 16'd36074, 16'd56498, 16'd44974, 16'd1083, 16'd29036, 16'd12244, 16'd61161, 16'd10309, 16'd50328, 16'd18834, 16'd5439, 16'd45505, 16'd34676, 16'd54768});
	test_expansion(128'hc19cf9403d015301fcd4e5bb1cb160c6, {16'd47206, 16'd2307, 16'd45390, 16'd16588, 16'd13197, 16'd11666, 16'd35035, 16'd26374, 16'd22717, 16'd26339, 16'd46967, 16'd48648, 16'd9573, 16'd34197, 16'd11027, 16'd38498, 16'd6737, 16'd2185, 16'd7258, 16'd49763, 16'd37434, 16'd48712, 16'd36643, 16'd1262, 16'd58031, 16'd43086});
	test_expansion(128'h422a12d8daec5f5e728d5860bca679c8, {16'd8891, 16'd19664, 16'd60269, 16'd55114, 16'd25546, 16'd64338, 16'd43590, 16'd16905, 16'd50446, 16'd11047, 16'd15035, 16'd14002, 16'd28779, 16'd43816, 16'd41009, 16'd4225, 16'd64565, 16'd53052, 16'd32029, 16'd11189, 16'd38819, 16'd20836, 16'd6426, 16'd58969, 16'd36240, 16'd57248});
	test_expansion(128'h63d059a7057c0f9fc4db274a9e5a5930, {16'd18083, 16'd16984, 16'd30217, 16'd58630, 16'd11290, 16'd36416, 16'd64436, 16'd34502, 16'd42868, 16'd3990, 16'd46123, 16'd44564, 16'd57035, 16'd32950, 16'd25933, 16'd18981, 16'd56934, 16'd31952, 16'd27541, 16'd52368, 16'd17703, 16'd46131, 16'd12830, 16'd51375, 16'd55959, 16'd22161});
	test_expansion(128'h82d26b3359e1e1d70732e11f161938fd, {16'd30680, 16'd3183, 16'd8734, 16'd44253, 16'd17147, 16'd53117, 16'd39081, 16'd11513, 16'd18329, 16'd59064, 16'd50075, 16'd19866, 16'd19176, 16'd42142, 16'd53047, 16'd44660, 16'd45080, 16'd17093, 16'd54651, 16'd42116, 16'd40411, 16'd43704, 16'd30590, 16'd56380, 16'd31794, 16'd49423});
	test_expansion(128'h8be4fa0e865e5a61ef1be243319542a7, {16'd50283, 16'd40739, 16'd63490, 16'd19275, 16'd29214, 16'd42695, 16'd23660, 16'd20737, 16'd19271, 16'd36841, 16'd28722, 16'd7481, 16'd25406, 16'd8206, 16'd55997, 16'd56404, 16'd20161, 16'd58872, 16'd57960, 16'd30458, 16'd2929, 16'd55521, 16'd8024, 16'd26201, 16'd37072, 16'd31551});
	test_expansion(128'hdcbfd3e4730324552b54ce390b046e0b, {16'd42373, 16'd12353, 16'd48051, 16'd21740, 16'd55251, 16'd21994, 16'd54374, 16'd26817, 16'd36339, 16'd5063, 16'd7002, 16'd50394, 16'd37752, 16'd35676, 16'd29016, 16'd38234, 16'd64194, 16'd21870, 16'd8130, 16'd64571, 16'd27208, 16'd27570, 16'd9711, 16'd64427, 16'd40107, 16'd34657});
	test_expansion(128'hfcdbb95383adc732a508ada43e82851f, {16'd41244, 16'd26043, 16'd27304, 16'd28221, 16'd25797, 16'd11757, 16'd55189, 16'd25800, 16'd22311, 16'd41440, 16'd50366, 16'd45614, 16'd50778, 16'd23891, 16'd23829, 16'd37645, 16'd9431, 16'd30182, 16'd38553, 16'd39304, 16'd24551, 16'd14899, 16'd23092, 16'd17530, 16'd41119, 16'd48364});
	test_expansion(128'h937e2f233614a43db439d96d09b448d2, {16'd8358, 16'd4870, 16'd51248, 16'd52034, 16'd35716, 16'd12141, 16'd53568, 16'd48579, 16'd21018, 16'd9373, 16'd42179, 16'd64559, 16'd24900, 16'd29192, 16'd63025, 16'd14307, 16'd32865, 16'd12025, 16'd52433, 16'd43311, 16'd618, 16'd57928, 16'd49604, 16'd8274, 16'd19931, 16'd33626});
	test_expansion(128'h957752dcc70e74f65a830e96ace095e0, {16'd13410, 16'd38914, 16'd57135, 16'd613, 16'd2644, 16'd13120, 16'd37020, 16'd45504, 16'd64700, 16'd17722, 16'd21802, 16'd31706, 16'd39735, 16'd14315, 16'd34622, 16'd22431, 16'd32300, 16'd12661, 16'd32287, 16'd53054, 16'd38314, 16'd22752, 16'd41004, 16'd63694, 16'd44083, 16'd40072});
	test_expansion(128'h6111ac5af3256213f1833956f0478d69, {16'd52334, 16'd34301, 16'd58560, 16'd62087, 16'd49972, 16'd15179, 16'd3084, 16'd60107, 16'd50171, 16'd48539, 16'd61998, 16'd18892, 16'd25358, 16'd60355, 16'd64306, 16'd11761, 16'd12316, 16'd51497, 16'd3004, 16'd23979, 16'd16147, 16'd3930, 16'd35759, 16'd31549, 16'd11357, 16'd41220});
	test_expansion(128'hbcfdcafa9f4966a005b0c5778d0db402, {16'd2507, 16'd63647, 16'd64848, 16'd48261, 16'd47943, 16'd16484, 16'd11272, 16'd60718, 16'd52787, 16'd50747, 16'd58218, 16'd19456, 16'd45319, 16'd36989, 16'd43895, 16'd54929, 16'd56752, 16'd60679, 16'd9728, 16'd40217, 16'd17505, 16'd63480, 16'd6127, 16'd26043, 16'd38453, 16'd51539});
	test_expansion(128'h6ca3f052a136ec42711df718c8dd14a7, {16'd56356, 16'd8197, 16'd53014, 16'd43862, 16'd21379, 16'd16674, 16'd44117, 16'd25801, 16'd12571, 16'd32446, 16'd39789, 16'd13767, 16'd30677, 16'd64193, 16'd32909, 16'd21070, 16'd23541, 16'd13317, 16'd60180, 16'd35738, 16'd46714, 16'd58112, 16'd59814, 16'd56260, 16'd9, 16'd20478});
	test_expansion(128'he820737b1a1ca2f9ff28ad15d6b856a8, {16'd37002, 16'd43790, 16'd212, 16'd8940, 16'd29163, 16'd61896, 16'd30269, 16'd56455, 16'd8243, 16'd60199, 16'd34766, 16'd54760, 16'd34365, 16'd9178, 16'd13411, 16'd50978, 16'd4117, 16'd11836, 16'd7863, 16'd37088, 16'd62550, 16'd39784, 16'd32930, 16'd7852, 16'd26633, 16'd7613});
	test_expansion(128'h6e769c43b495c0a28a6cb18c60c0c88e, {16'd56827, 16'd21737, 16'd40540, 16'd48782, 16'd46767, 16'd3020, 16'd64993, 16'd38598, 16'd47135, 16'd54290, 16'd15511, 16'd49550, 16'd54928, 16'd31246, 16'd18363, 16'd46812, 16'd49943, 16'd23415, 16'd33903, 16'd35596, 16'd11041, 16'd7664, 16'd60857, 16'd37044, 16'd41539, 16'd44155});
	test_expansion(128'h98e9ac692178e440200889ebdc836e9f, {16'd17544, 16'd23481, 16'd44418, 16'd38983, 16'd36635, 16'd4704, 16'd60318, 16'd44829, 16'd62617, 16'd14881, 16'd57645, 16'd46716, 16'd20086, 16'd21952, 16'd48848, 16'd36428, 16'd33599, 16'd62054, 16'd15762, 16'd61434, 16'd50909, 16'd8431, 16'd64504, 16'd61228, 16'd37427, 16'd17751});
	test_expansion(128'h2f99b8eaa7a70cdb50adc471dd21d436, {16'd5956, 16'd25990, 16'd8200, 16'd63755, 16'd18126, 16'd1944, 16'd43779, 16'd10034, 16'd25411, 16'd59076, 16'd44173, 16'd62283, 16'd28711, 16'd23255, 16'd26784, 16'd24889, 16'd9071, 16'd22972, 16'd23537, 16'd909, 16'd42440, 16'd4789, 16'd64115, 16'd46367, 16'd15540, 16'd51412});
	test_expansion(128'hf30e193dfc68d9613aa14d2f93de22d8, {16'd27297, 16'd12242, 16'd14973, 16'd20218, 16'd45204, 16'd60573, 16'd10419, 16'd43026, 16'd41226, 16'd26041, 16'd36880, 16'd27393, 16'd14868, 16'd2377, 16'd20650, 16'd2414, 16'd58323, 16'd62611, 16'd11013, 16'd63831, 16'd48107, 16'd59145, 16'd37429, 16'd65206, 16'd24988, 16'd10511});
	test_expansion(128'hbc274bcd107d18cb7cf8794aa01e7331, {16'd47361, 16'd60242, 16'd65431, 16'd61327, 16'd65089, 16'd35227, 16'd39720, 16'd23717, 16'd35018, 16'd7316, 16'd47714, 16'd58541, 16'd4894, 16'd9488, 16'd9969, 16'd34421, 16'd56842, 16'd46436, 16'd56668, 16'd35270, 16'd689, 16'd29369, 16'd32488, 16'd29756, 16'd18680, 16'd52733});
	test_expansion(128'h1454a14e8ba58baa29c0525873a22608, {16'd61112, 16'd55269, 16'd41297, 16'd60915, 16'd48724, 16'd14616, 16'd3452, 16'd59470, 16'd20820, 16'd45975, 16'd39658, 16'd53976, 16'd46418, 16'd32177, 16'd14478, 16'd62068, 16'd49314, 16'd61154, 16'd16704, 16'd63368, 16'd18632, 16'd48452, 16'd45994, 16'd40188, 16'd46121, 16'd42046});
	test_expansion(128'hb8895fc2cb026e275e094c4ac9e11481, {16'd59193, 16'd46369, 16'd45483, 16'd28460, 16'd15340, 16'd34349, 16'd61766, 16'd51173, 16'd35725, 16'd63125, 16'd10529, 16'd47129, 16'd7409, 16'd17373, 16'd9619, 16'd65332, 16'd56650, 16'd13544, 16'd47584, 16'd53282, 16'd43978, 16'd7064, 16'd37875, 16'd50849, 16'd13918, 16'd64836});
	test_expansion(128'hb0c2f7c4310c966976858d8050855b8f, {16'd56731, 16'd38450, 16'd61550, 16'd61852, 16'd31639, 16'd15421, 16'd59147, 16'd62059, 16'd39686, 16'd25198, 16'd42399, 16'd37954, 16'd23508, 16'd27487, 16'd20948, 16'd38318, 16'd42526, 16'd4464, 16'd18288, 16'd39225, 16'd19610, 16'd11280, 16'd62417, 16'd53463, 16'd8603, 16'd40940});
	test_expansion(128'hac031fd636a97e507283901fb09b8dfd, {16'd8335, 16'd30484, 16'd61302, 16'd17704, 16'd54758, 16'd12614, 16'd62420, 16'd35989, 16'd23422, 16'd63442, 16'd33879, 16'd18674, 16'd25935, 16'd61286, 16'd43886, 16'd7229, 16'd38873, 16'd33570, 16'd3501, 16'd28991, 16'd45048, 16'd32535, 16'd38716, 16'd19286, 16'd57472, 16'd36827});
	test_expansion(128'h7a8abdee380ba56334fb6cc45212df87, {16'd57258, 16'd48100, 16'd27934, 16'd242, 16'd20149, 16'd32889, 16'd64692, 16'd37508, 16'd50405, 16'd12312, 16'd42702, 16'd23124, 16'd63783, 16'd47472, 16'd37518, 16'd1370, 16'd52322, 16'd34507, 16'd47231, 16'd47507, 16'd32809, 16'd59337, 16'd14544, 16'd7093, 16'd20934, 16'd40893});
	test_expansion(128'hfda0744388a38a0a4fda9e68a359ebbf, {16'd56412, 16'd26714, 16'd4860, 16'd17846, 16'd55841, 16'd50996, 16'd33056, 16'd28747, 16'd42751, 16'd47139, 16'd57960, 16'd30671, 16'd42334, 16'd29686, 16'd7929, 16'd15146, 16'd46699, 16'd3196, 16'd9124, 16'd60027, 16'd37858, 16'd46514, 16'd13959, 16'd58197, 16'd16438, 16'd54577});
	test_expansion(128'h2c78299e4dad3f946a91608e2eb6c0b5, {16'd59837, 16'd48991, 16'd18661, 16'd19505, 16'd45996, 16'd8960, 16'd19642, 16'd27185, 16'd48590, 16'd9423, 16'd3416, 16'd10781, 16'd15032, 16'd16840, 16'd26173, 16'd45673, 16'd22493, 16'd38716, 16'd56655, 16'd6859, 16'd46956, 16'd14203, 16'd65092, 16'd63745, 16'd39338, 16'd15061});
	test_expansion(128'he6ba894de6705d56d3e6b75661ef7ed8, {16'd42059, 16'd31220, 16'd6713, 16'd30077, 16'd58078, 16'd1397, 16'd30426, 16'd18735, 16'd29772, 16'd64175, 16'd12813, 16'd12584, 16'd28448, 16'd20664, 16'd1484, 16'd2237, 16'd38670, 16'd26408, 16'd27128, 16'd11032, 16'd650, 16'd613, 16'd22186, 16'd16226, 16'd45486, 16'd55703});
	test_expansion(128'h08400fbe5cd33b3be4877d60daf2230c, {16'd17089, 16'd53758, 16'd61150, 16'd29704, 16'd10816, 16'd21748, 16'd58394, 16'd23974, 16'd5432, 16'd4918, 16'd55092, 16'd50169, 16'd39829, 16'd31606, 16'd48697, 16'd28637, 16'd2711, 16'd33806, 16'd11136, 16'd59094, 16'd54084, 16'd15502, 16'd61, 16'd39942, 16'd41957, 16'd18500});
	test_expansion(128'hacd1c03f67ce9eaca7eff44d8cfdb5ed, {16'd40620, 16'd40359, 16'd29146, 16'd19461, 16'd13115, 16'd49197, 16'd54726, 16'd51653, 16'd57675, 16'd64739, 16'd32116, 16'd44508, 16'd42145, 16'd29082, 16'd60667, 16'd8835, 16'd40838, 16'd58202, 16'd40063, 16'd63131, 16'd36531, 16'd22170, 16'd18227, 16'd1115, 16'd234, 16'd13501});
	test_expansion(128'h838b09dc144c921e4c6ec6c544a2f15a, {16'd52049, 16'd43908, 16'd20816, 16'd38167, 16'd35659, 16'd21993, 16'd29340, 16'd144, 16'd17039, 16'd48171, 16'd39058, 16'd1484, 16'd18718, 16'd42787, 16'd8938, 16'd4155, 16'd28246, 16'd65194, 16'd58010, 16'd23417, 16'd51156, 16'd65512, 16'd56852, 16'd44422, 16'd430, 16'd7219});
	test_expansion(128'h77a7f0d0ae33f3fa3d28199cc81ee341, {16'd11044, 16'd11531, 16'd63240, 16'd40095, 16'd26281, 16'd6697, 16'd43659, 16'd21007, 16'd47915, 16'd62027, 16'd51305, 16'd48630, 16'd46974, 16'd31331, 16'd57314, 16'd47405, 16'd10950, 16'd42760, 16'd42872, 16'd13557, 16'd33907, 16'd57451, 16'd32523, 16'd19007, 16'd51047, 16'd14550});
	test_expansion(128'h4fede245091cbb4c3093ea9968451245, {16'd12697, 16'd57700, 16'd47583, 16'd14473, 16'd52121, 16'd63154, 16'd57040, 16'd56993, 16'd59790, 16'd13956, 16'd56763, 16'd14829, 16'd18506, 16'd17837, 16'd14623, 16'd26940, 16'd21496, 16'd16478, 16'd46305, 16'd16914, 16'd15214, 16'd5138, 16'd12000, 16'd8213, 16'd38508, 16'd30308});
	test_expansion(128'h646472c455e1c94828549ac175265360, {16'd7761, 16'd6168, 16'd47392, 16'd48932, 16'd34287, 16'd28888, 16'd9420, 16'd16969, 16'd37373, 16'd39872, 16'd24534, 16'd57404, 16'd15754, 16'd3402, 16'd5506, 16'd30533, 16'd56512, 16'd20485, 16'd20109, 16'd18571, 16'd30786, 16'd25697, 16'd46079, 16'd64485, 16'd11604, 16'd17910});
	test_expansion(128'h6dd845fe1c5b6c3d89a2d5e5bb69a44d, {16'd9076, 16'd57327, 16'd38041, 16'd63991, 16'd14165, 16'd49668, 16'd20918, 16'd38707, 16'd23272, 16'd46902, 16'd11737, 16'd29278, 16'd20597, 16'd23319, 16'd61714, 16'd9192, 16'd34102, 16'd24423, 16'd11323, 16'd11244, 16'd3889, 16'd15179, 16'd58450, 16'd57892, 16'd52580, 16'd20543});
	test_expansion(128'hfac9d1b523f8b2985ff112560f381b77, {16'd9285, 16'd58704, 16'd50874, 16'd47536, 16'd18087, 16'd24610, 16'd4616, 16'd3459, 16'd10184, 16'd2246, 16'd35471, 16'd26392, 16'd15133, 16'd35084, 16'd27175, 16'd34039, 16'd17363, 16'd49310, 16'd44258, 16'd54691, 16'd5719, 16'd44176, 16'd6100, 16'd14960, 16'd16106, 16'd36693});
	test_expansion(128'h92e9d6642098ee2a266e8b9079b6aa27, {16'd19255, 16'd39048, 16'd40470, 16'd40160, 16'd17775, 16'd46403, 16'd38006, 16'd59409, 16'd22082, 16'd46394, 16'd13936, 16'd1092, 16'd54368, 16'd39370, 16'd57877, 16'd5564, 16'd28878, 16'd36593, 16'd40767, 16'd14625, 16'd42458, 16'd17503, 16'd15484, 16'd45089, 16'd19173, 16'd55786});
	test_expansion(128'h20e07c20645f1bcdad7306c906c68314, {16'd4741, 16'd61565, 16'd27908, 16'd13527, 16'd24641, 16'd25946, 16'd17847, 16'd5479, 16'd10782, 16'd28673, 16'd38375, 16'd34063, 16'd58460, 16'd35392, 16'd34469, 16'd52053, 16'd63570, 16'd18045, 16'd26927, 16'd17584, 16'd49416, 16'd43621, 16'd993, 16'd16418, 16'd15069, 16'd60789});
	test_expansion(128'h6eaaca11bdc9863232da0463d623d2fb, {16'd18295, 16'd65228, 16'd30019, 16'd18132, 16'd28594, 16'd23928, 16'd3852, 16'd58177, 16'd17109, 16'd63546, 16'd42297, 16'd6122, 16'd60981, 16'd45599, 16'd60524, 16'd10024, 16'd31078, 16'd47019, 16'd25570, 16'd12985, 16'd29091, 16'd40872, 16'd52434, 16'd60659, 16'd13089, 16'd2727});
	test_expansion(128'h10938bbd2ad6f4a413ab439296558faa, {16'd12798, 16'd49563, 16'd722, 16'd35772, 16'd24095, 16'd60084, 16'd35077, 16'd54744, 16'd11867, 16'd28954, 16'd20699, 16'd41910, 16'd2842, 16'd29870, 16'd52640, 16'd22227, 16'd46997, 16'd45901, 16'd58570, 16'd39972, 16'd14950, 16'd62548, 16'd14954, 16'd18720, 16'd1376, 16'd32597});
	test_expansion(128'h81294362e830f8303f4e9388762808fd, {16'd16849, 16'd41996, 16'd46434, 16'd30075, 16'd24755, 16'd62500, 16'd1592, 16'd48156, 16'd46023, 16'd21746, 16'd57399, 16'd10740, 16'd38640, 16'd1129, 16'd15685, 16'd36069, 16'd31671, 16'd37924, 16'd29763, 16'd35240, 16'd45158, 16'd14237, 16'd12163, 16'd51704, 16'd59406, 16'd30341});
	test_expansion(128'ha45387170418aa2ca4af4de1e826f515, {16'd22424, 16'd23411, 16'd62274, 16'd8325, 16'd34976, 16'd8870, 16'd54379, 16'd51171, 16'd35268, 16'd47144, 16'd15421, 16'd12093, 16'd32869, 16'd40632, 16'd22618, 16'd50993, 16'd49759, 16'd42850, 16'd19961, 16'd24698, 16'd34526, 16'd33987, 16'd6092, 16'd5467, 16'd38368, 16'd33946});
	test_expansion(128'h9e4883fd7eb042d6763f97c11079c347, {16'd64274, 16'd60323, 16'd46442, 16'd19365, 16'd58851, 16'd34097, 16'd4820, 16'd58591, 16'd44889, 16'd44022, 16'd8597, 16'd59937, 16'd60711, 16'd15566, 16'd44839, 16'd27280, 16'd40938, 16'd14364, 16'd21909, 16'd58740, 16'd64266, 16'd35456, 16'd11855, 16'd31391, 16'd58626, 16'd61652});
	test_expansion(128'h5a6303c600841f5b9a749cb1605d40ae, {16'd32985, 16'd44795, 16'd64565, 16'd23003, 16'd35708, 16'd19230, 16'd30250, 16'd57090, 16'd30196, 16'd57868, 16'd27893, 16'd39445, 16'd52948, 16'd52209, 16'd50043, 16'd6270, 16'd9400, 16'd1680, 16'd60974, 16'd18893, 16'd18983, 16'd2635, 16'd45730, 16'd17023, 16'd51674, 16'd51493});
	test_expansion(128'hdbbc997a55c1a961d1cb8a9611cc254c, {16'd55767, 16'd20450, 16'd23884, 16'd6088, 16'd35164, 16'd25941, 16'd13382, 16'd1130, 16'd7491, 16'd30816, 16'd54431, 16'd33765, 16'd2948, 16'd63661, 16'd8221, 16'd45738, 16'd55029, 16'd47743, 16'd26415, 16'd36936, 16'd15283, 16'd34862, 16'd30971, 16'd33879, 16'd3150, 16'd8148});
	test_expansion(128'h4927bb25646dcfc3c2bcd24619c70261, {16'd42513, 16'd37147, 16'd38952, 16'd26163, 16'd24914, 16'd57952, 16'd47930, 16'd42002, 16'd23079, 16'd34666, 16'd29533, 16'd40130, 16'd31838, 16'd59772, 16'd26357, 16'd7340, 16'd14525, 16'd26773, 16'd22556, 16'd53007, 16'd20323, 16'd55785, 16'd10627, 16'd7566, 16'd29452, 16'd18033});
	test_expansion(128'h4a4ec721b3c5824737de93420f8204b0, {16'd24002, 16'd13950, 16'd40412, 16'd6491, 16'd25888, 16'd21663, 16'd26475, 16'd18598, 16'd52625, 16'd30582, 16'd21089, 16'd29771, 16'd61491, 16'd50238, 16'd6647, 16'd65254, 16'd37808, 16'd44176, 16'd54284, 16'd5621, 16'd1352, 16'd61998, 16'd40025, 16'd54594, 16'd35571, 16'd37592});
	test_expansion(128'h5c33f080ebdb16e27fe5c7cab4f61786, {16'd916, 16'd29814, 16'd28311, 16'd38802, 16'd39649, 16'd51839, 16'd55193, 16'd44281, 16'd37713, 16'd63237, 16'd63754, 16'd5917, 16'd22236, 16'd833, 16'd45560, 16'd28405, 16'd39206, 16'd35801, 16'd7147, 16'd54506, 16'd50462, 16'd58267, 16'd41943, 16'd33978, 16'd39890, 16'd43439});
	test_expansion(128'hb4e8a2a061308a6d375ef8befdf6b8e8, {16'd17945, 16'd26121, 16'd62138, 16'd5126, 16'd20479, 16'd36012, 16'd47656, 16'd1647, 16'd35792, 16'd17967, 16'd31013, 16'd46923, 16'd49986, 16'd35642, 16'd56385, 16'd37327, 16'd6863, 16'd53753, 16'd14256, 16'd12741, 16'd25203, 16'd59639, 16'd48567, 16'd16921, 16'd39440, 16'd11561});
	test_expansion(128'h298c7ca0b9ad8dea45931761c6ccbcc3, {16'd59955, 16'd55521, 16'd22551, 16'd51909, 16'd49122, 16'd55130, 16'd43802, 16'd19027, 16'd9619, 16'd41111, 16'd37971, 16'd13154, 16'd18207, 16'd48331, 16'd54262, 16'd32631, 16'd19867, 16'd54242, 16'd56753, 16'd14017, 16'd31473, 16'd7392, 16'd35291, 16'd29396, 16'd7156, 16'd2909});
	test_expansion(128'hb1aeac4c279038e10ad14adf00d8ed03, {16'd39229, 16'd49037, 16'd42070, 16'd20563, 16'd44287, 16'd7716, 16'd49943, 16'd2023, 16'd313, 16'd30554, 16'd58405, 16'd19679, 16'd22813, 16'd17048, 16'd3680, 16'd57760, 16'd40631, 16'd34540, 16'd5190, 16'd14632, 16'd30764, 16'd16281, 16'd64781, 16'd10596, 16'd14264, 16'd21931});
	test_expansion(128'h7d7952c9f112ba23d462973bebffff8d, {16'd43899, 16'd54809, 16'd19466, 16'd7485, 16'd61782, 16'd57026, 16'd55052, 16'd42378, 16'd14910, 16'd12188, 16'd29796, 16'd40296, 16'd15881, 16'd41297, 16'd12905, 16'd21572, 16'd65067, 16'd60472, 16'd10155, 16'd32454, 16'd51240, 16'd26575, 16'd54908, 16'd37824, 16'd7829, 16'd62724});
	test_expansion(128'h8857111c177e768833bf270682cb8586, {16'd25923, 16'd43180, 16'd59223, 16'd28744, 16'd58710, 16'd56066, 16'd53771, 16'd60362, 16'd7423, 16'd32044, 16'd63900, 16'd16001, 16'd35425, 16'd14160, 16'd64249, 16'd51022, 16'd32931, 16'd17996, 16'd2949, 16'd36265, 16'd20009, 16'd26378, 16'd57538, 16'd2812, 16'd8575, 16'd14097});
	test_expansion(128'hfd83c625421b9f92286c4ce9a7c0d69c, {16'd57899, 16'd26651, 16'd22789, 16'd12406, 16'd4689, 16'd21098, 16'd20058, 16'd1413, 16'd55812, 16'd38840, 16'd45246, 16'd57127, 16'd30960, 16'd23274, 16'd18758, 16'd30862, 16'd16188, 16'd9310, 16'd31691, 16'd55521, 16'd4127, 16'd40201, 16'd63386, 16'd14892, 16'd54744, 16'd5545});
	test_expansion(128'hbbc0678b9e7fa820837e844021a9c31f, {16'd51702, 16'd47400, 16'd41136, 16'd48655, 16'd35271, 16'd44579, 16'd63847, 16'd41447, 16'd22512, 16'd51104, 16'd3209, 16'd59409, 16'd58529, 16'd52006, 16'd3282, 16'd51775, 16'd7113, 16'd33185, 16'd21464, 16'd36654, 16'd4787, 16'd43605, 16'd53587, 16'd46196, 16'd37090, 16'd50662});
	test_expansion(128'hecbcac8db1e0363eaf594c6213dab12c, {16'd33516, 16'd19501, 16'd37432, 16'd56826, 16'd22031, 16'd30109, 16'd6206, 16'd65277, 16'd45841, 16'd419, 16'd20454, 16'd4216, 16'd47263, 16'd18609, 16'd61390, 16'd56770, 16'd18446, 16'd5740, 16'd18380, 16'd49385, 16'd54206, 16'd41882, 16'd61333, 16'd11542, 16'd32429, 16'd55632});
	test_expansion(128'hb4fc4844ee9326900f560e1f45b566ae, {16'd56867, 16'd56990, 16'd29599, 16'd27612, 16'd46385, 16'd5756, 16'd23546, 16'd29047, 16'd30625, 16'd40302, 16'd52262, 16'd14517, 16'd24258, 16'd3525, 16'd29676, 16'd55556, 16'd61111, 16'd43084, 16'd27124, 16'd61404, 16'd63656, 16'd41659, 16'd42939, 16'd29915, 16'd52370, 16'd4021});
	test_expansion(128'hacba0a12956092d798cdedcdd4f6c0d3, {16'd11148, 16'd10317, 16'd61466, 16'd35014, 16'd29754, 16'd65392, 16'd8753, 16'd11982, 16'd14439, 16'd38208, 16'd42480, 16'd1720, 16'd32227, 16'd53898, 16'd54600, 16'd54664, 16'd4401, 16'd22095, 16'd22025, 16'd9073, 16'd15558, 16'd37878, 16'd41027, 16'd17222, 16'd14296, 16'd5365});
	test_expansion(128'h88e7635b347d9fb639af3372c947bd4c, {16'd48984, 16'd47325, 16'd62835, 16'd14445, 16'd46466, 16'd5852, 16'd35, 16'd54019, 16'd40548, 16'd42936, 16'd32408, 16'd43915, 16'd33143, 16'd1065, 16'd26658, 16'd15114, 16'd14472, 16'd15301, 16'd32431, 16'd20427, 16'd11814, 16'd10567, 16'd56095, 16'd37702, 16'd823, 16'd34924});
	test_expansion(128'h83ecc1b38745a62e1a970ea33eb121bb, {16'd28524, 16'd57539, 16'd36245, 16'd7200, 16'd6577, 16'd57500, 16'd19148, 16'd11684, 16'd41981, 16'd61050, 16'd21426, 16'd28432, 16'd52694, 16'd32776, 16'd26271, 16'd41454, 16'd51818, 16'd42293, 16'd9631, 16'd2677, 16'd63392, 16'd58945, 16'd12501, 16'd23168, 16'd48074, 16'd28884});
	test_expansion(128'h6a2b42c88644cf47d9bcb292591e6ee4, {16'd48750, 16'd48263, 16'd26678, 16'd27976, 16'd59824, 16'd55462, 16'd23943, 16'd57555, 16'd45435, 16'd31607, 16'd25946, 16'd31464, 16'd27006, 16'd3196, 16'd33044, 16'd21801, 16'd60129, 16'd44990, 16'd63091, 16'd53740, 16'd27166, 16'd8269, 16'd54821, 16'd16881, 16'd38529, 16'd63035});
	test_expansion(128'h921f8583b291360a50b51143e6bed6e5, {16'd43331, 16'd49252, 16'd5011, 16'd21070, 16'd35691, 16'd57668, 16'd31452, 16'd39673, 16'd61561, 16'd50402, 16'd8416, 16'd38276, 16'd50582, 16'd56475, 16'd61516, 16'd23399, 16'd49736, 16'd1860, 16'd56613, 16'd2470, 16'd28041, 16'd32988, 16'd1562, 16'd1127, 16'd7946, 16'd47541});
	test_expansion(128'hee8bea7b1df28b65020e2dd3b245fe48, {16'd7895, 16'd65149, 16'd20938, 16'd16223, 16'd25331, 16'd48327, 16'd9607, 16'd58274, 16'd30783, 16'd36082, 16'd21631, 16'd46638, 16'd53644, 16'd3762, 16'd44503, 16'd1374, 16'd57953, 16'd53797, 16'd29576, 16'd51865, 16'd58958, 16'd11462, 16'd4138, 16'd43770, 16'd58150, 16'd41436});
	test_expansion(128'hcc7de9ec1e63dcfb47e5fceb5389ba32, {16'd25490, 16'd57437, 16'd58613, 16'd48150, 16'd12037, 16'd6298, 16'd51091, 16'd23950, 16'd1437, 16'd21807, 16'd7159, 16'd49444, 16'd36523, 16'd62069, 16'd16269, 16'd3450, 16'd7430, 16'd62092, 16'd50260, 16'd49584, 16'd55561, 16'd7855, 16'd53826, 16'd24320, 16'd62574, 16'd26349});
	test_expansion(128'h724a2da070320a2ac0f02f043660ac8d, {16'd43501, 16'd20951, 16'd61506, 16'd14241, 16'd28494, 16'd3876, 16'd53876, 16'd56507, 16'd4316, 16'd38364, 16'd14827, 16'd33738, 16'd9286, 16'd33044, 16'd57448, 16'd50890, 16'd59817, 16'd717, 16'd34200, 16'd24289, 16'd14951, 16'd31729, 16'd21789, 16'd12325, 16'd554, 16'd37610});
	test_expansion(128'h2f69be1de5a102f4261fe647a1b2357e, {16'd28671, 16'd5679, 16'd27937, 16'd64938, 16'd51601, 16'd64637, 16'd10010, 16'd33970, 16'd2451, 16'd64212, 16'd39372, 16'd31670, 16'd19239, 16'd30905, 16'd30768, 16'd63884, 16'd21641, 16'd60490, 16'd31781, 16'd55817, 16'd21936, 16'd32665, 16'd28800, 16'd38051, 16'd47460, 16'd61337});
	test_expansion(128'ha75802b04a09e2ba74fbb56c1f8ac130, {16'd26596, 16'd7234, 16'd51255, 16'd37163, 16'd13036, 16'd8204, 16'd50233, 16'd36649, 16'd58173, 16'd5466, 16'd36365, 16'd6103, 16'd23122, 16'd50068, 16'd46504, 16'd15123, 16'd14694, 16'd16234, 16'd59278, 16'd12851, 16'd31901, 16'd9611, 16'd28717, 16'd7740, 16'd4945, 16'd40284});
	test_expansion(128'hd4946a35708e9ac7add8cf767a3b5df5, {16'd43025, 16'd29458, 16'd7470, 16'd24800, 16'd38508, 16'd46647, 16'd40273, 16'd49202, 16'd5584, 16'd20404, 16'd44687, 16'd56889, 16'd25175, 16'd36491, 16'd39769, 16'd32774, 16'd4058, 16'd60558, 16'd31225, 16'd22610, 16'd43409, 16'd26970, 16'd19190, 16'd4121, 16'd63942, 16'd61303});
	test_expansion(128'he4beb48e197f30846141cdec0ffc6bcf, {16'd46606, 16'd17485, 16'd26844, 16'd44860, 16'd53666, 16'd9647, 16'd23980, 16'd40595, 16'd56069, 16'd25401, 16'd40207, 16'd9463, 16'd55080, 16'd10618, 16'd34189, 16'd46236, 16'd11573, 16'd59529, 16'd14482, 16'd19182, 16'd5262, 16'd37850, 16'd44660, 16'd49397, 16'd26562, 16'd26606});
	test_expansion(128'h0cc414e0a145e33d8f7bef2f03ae5cda, {16'd9279, 16'd29863, 16'd58163, 16'd31822, 16'd31870, 16'd5403, 16'd30672, 16'd38252, 16'd535, 16'd28671, 16'd24146, 16'd14613, 16'd38762, 16'd47797, 16'd48091, 16'd17022, 16'd2107, 16'd61980, 16'd51957, 16'd56001, 16'd8497, 16'd43575, 16'd34366, 16'd36458, 16'd21302, 16'd11945});
	test_expansion(128'hd543c0c12ddca97f02ed740f3f35cd34, {16'd59372, 16'd60034, 16'd16139, 16'd28979, 16'd42119, 16'd65038, 16'd20989, 16'd5788, 16'd18194, 16'd45418, 16'd47859, 16'd13780, 16'd33473, 16'd52413, 16'd29144, 16'd58176, 16'd49733, 16'd47320, 16'd49462, 16'd29230, 16'd45118, 16'd55327, 16'd706, 16'd54547, 16'd20540, 16'd64654});
	test_expansion(128'hb6b4b20b78dfd56204e30c1171d856a6, {16'd30695, 16'd18514, 16'd17269, 16'd16757, 16'd23861, 16'd26407, 16'd20691, 16'd23400, 16'd51878, 16'd39555, 16'd6316, 16'd5691, 16'd47499, 16'd11241, 16'd36065, 16'd53545, 16'd50932, 16'd48680, 16'd65121, 16'd737, 16'd7234, 16'd22265, 16'd56759, 16'd46695, 16'd32013, 16'd43816});
	test_expansion(128'h3bfbf1a3507d4398e4532a1d774fca99, {16'd37927, 16'd15949, 16'd32760, 16'd24846, 16'd16001, 16'd23380, 16'd17823, 16'd45863, 16'd23285, 16'd4588, 16'd12455, 16'd17617, 16'd53599, 16'd60559, 16'd42508, 16'd14256, 16'd45787, 16'd63148, 16'd36767, 16'd11191, 16'd8144, 16'd57344, 16'd36704, 16'd37118, 16'd17627, 16'd13175});
	test_expansion(128'h297cd44bb08f4a3ea3e3d30b90f83bae, {16'd7510, 16'd38371, 16'd8263, 16'd50158, 16'd34501, 16'd9922, 16'd42577, 16'd26210, 16'd23839, 16'd42497, 16'd16835, 16'd37065, 16'd62895, 16'd38041, 16'd31549, 16'd15616, 16'd50838, 16'd5428, 16'd13897, 16'd47197, 16'd14300, 16'd51062, 16'd20947, 16'd35548, 16'd55602, 16'd16723});
	test_expansion(128'h87e11c3c46d55866b4487e4766dfd0a6, {16'd42476, 16'd22750, 16'd47065, 16'd3765, 16'd23817, 16'd62346, 16'd6012, 16'd38704, 16'd5228, 16'd62526, 16'd17907, 16'd12146, 16'd18474, 16'd8134, 16'd7987, 16'd64294, 16'd38150, 16'd26931, 16'd398, 16'd10576, 16'd32204, 16'd10970, 16'd58132, 16'd1666, 16'd57827, 16'd17480});
	test_expansion(128'hb54bb990081dd2b3e47d11ea3efd7ac4, {16'd53656, 16'd20640, 16'd4152, 16'd59299, 16'd57732, 16'd23431, 16'd28382, 16'd46744, 16'd63027, 16'd28939, 16'd61019, 16'd49547, 16'd43666, 16'd61217, 16'd50739, 16'd27360, 16'd27523, 16'd58083, 16'd43844, 16'd54951, 16'd35844, 16'd23514, 16'd53423, 16'd8589, 16'd53801, 16'd37135});
	test_expansion(128'h370a6777d9b623fa2705ac67f6a58ca7, {16'd42125, 16'd12827, 16'd17954, 16'd18825, 16'd51490, 16'd24669, 16'd62358, 16'd4906, 16'd36841, 16'd9362, 16'd38634, 16'd3657, 16'd55007, 16'd61057, 16'd7958, 16'd36175, 16'd18098, 16'd53097, 16'd34097, 16'd33784, 16'd26461, 16'd40512, 16'd3703, 16'd19381, 16'd53931, 16'd54654});
	test_expansion(128'h983c972fed44f0ebd9522bff092703f6, {16'd61575, 16'd60243, 16'd36765, 16'd55369, 16'd25298, 16'd17213, 16'd49784, 16'd65382, 16'd35609, 16'd7845, 16'd33240, 16'd47979, 16'd37975, 16'd51438, 16'd8199, 16'd51734, 16'd37846, 16'd33793, 16'd47025, 16'd32761, 16'd27859, 16'd50790, 16'd52875, 16'd9825, 16'd40909, 16'd10329});
	test_expansion(128'h2bbc52f69ad17966bbed9567cbadb233, {16'd30780, 16'd55262, 16'd19894, 16'd54394, 16'd13039, 16'd54493, 16'd47275, 16'd35546, 16'd56967, 16'd2647, 16'd44776, 16'd36759, 16'd22969, 16'd31861, 16'd18070, 16'd53116, 16'd53795, 16'd52191, 16'd23287, 16'd34568, 16'd42479, 16'd9830, 16'd6973, 16'd7042, 16'd51599, 16'd30397});
	test_expansion(128'h60e2a02358054bef1c3adc17d7738929, {16'd51276, 16'd9123, 16'd26944, 16'd28618, 16'd17168, 16'd17586, 16'd63123, 16'd728, 16'd47828, 16'd32623, 16'd37316, 16'd15521, 16'd60905, 16'd53563, 16'd23040, 16'd48600, 16'd63321, 16'd19733, 16'd11862, 16'd5602, 16'd41695, 16'd13720, 16'd48927, 16'd6546, 16'd13635, 16'd50087});
	test_expansion(128'h4b6cd5a6003671aa53155862a0bfd662, {16'd53648, 16'd29852, 16'd30732, 16'd16559, 16'd33884, 16'd18150, 16'd5520, 16'd55388, 16'd10716, 16'd30935, 16'd14400, 16'd4711, 16'd18089, 16'd10166, 16'd55834, 16'd36157, 16'd6512, 16'd3657, 16'd51487, 16'd52842, 16'd12561, 16'd53144, 16'd3470, 16'd51900, 16'd20576, 16'd38355});
	test_expansion(128'hacf164f626b986b779e3da962ede04a2, {16'd62811, 16'd8734, 16'd58701, 16'd22034, 16'd21, 16'd15688, 16'd38732, 16'd897, 16'd52860, 16'd1974, 16'd23560, 16'd20962, 16'd28555, 16'd58253, 16'd44811, 16'd38425, 16'd20172, 16'd25802, 16'd65057, 16'd47167, 16'd24916, 16'd19248, 16'd30278, 16'd21252, 16'd29019, 16'd34298});
	test_expansion(128'ha5208db1245cfb90129f9dd092f8098c, {16'd59100, 16'd1418, 16'd45521, 16'd25347, 16'd52795, 16'd13295, 16'd61825, 16'd9674, 16'd33820, 16'd49875, 16'd15916, 16'd34145, 16'd64815, 16'd12429, 16'd23381, 16'd26705, 16'd53104, 16'd62994, 16'd28257, 16'd50081, 16'd21590, 16'd33284, 16'd2300, 16'd22177, 16'd34352, 16'd21168});
	test_expansion(128'hb183da65c070370afa47fcc80c378ff5, {16'd39477, 16'd55170, 16'd42531, 16'd4265, 16'd31000, 16'd58166, 16'd56310, 16'd20658, 16'd45481, 16'd26852, 16'd65494, 16'd32213, 16'd12243, 16'd19049, 16'd45995, 16'd30912, 16'd16517, 16'd59553, 16'd10504, 16'd41467, 16'd44857, 16'd44950, 16'd56922, 16'd24293, 16'd27863, 16'd18800});
	test_expansion(128'h9fbbaa41bdddd0757d7b5e29488d15df, {16'd29686, 16'd1839, 16'd86, 16'd12509, 16'd56440, 16'd10011, 16'd57305, 16'd15344, 16'd26100, 16'd2765, 16'd1374, 16'd2865, 16'd29004, 16'd46410, 16'd17172, 16'd18149, 16'd55646, 16'd15526, 16'd33558, 16'd18685, 16'd21029, 16'd19260, 16'd33902, 16'd12860, 16'd54453, 16'd4271});
	test_expansion(128'hab5fd7cccf860089ced15136fe3c2515, {16'd12208, 16'd24360, 16'd52944, 16'd63171, 16'd18840, 16'd34667, 16'd59763, 16'd20194, 16'd6969, 16'd60599, 16'd8752, 16'd4123, 16'd29223, 16'd40399, 16'd38129, 16'd44669, 16'd15533, 16'd6893, 16'd48666, 16'd17134, 16'd44125, 16'd60250, 16'd43116, 16'd62559, 16'd54490, 16'd39805});
	test_expansion(128'h7fde9be6a0b409fa441c0aa9710620e9, {16'd6348, 16'd15026, 16'd31991, 16'd59126, 16'd4948, 16'd5221, 16'd21950, 16'd37511, 16'd23151, 16'd19991, 16'd37977, 16'd28343, 16'd7094, 16'd35692, 16'd53005, 16'd35977, 16'd28798, 16'd61492, 16'd64583, 16'd3969, 16'd20191, 16'd6249, 16'd21146, 16'd31030, 16'd39957, 16'd15816});
	test_expansion(128'hf3e207f6d094a9852a574e3524bb5298, {16'd26204, 16'd36384, 16'd25714, 16'd26550, 16'd15133, 16'd57517, 16'd41257, 16'd47244, 16'd9189, 16'd6295, 16'd31625, 16'd22468, 16'd4087, 16'd41641, 16'd16964, 16'd21456, 16'd25090, 16'd11194, 16'd21371, 16'd38377, 16'd27374, 16'd58818, 16'd26256, 16'd29293, 16'd49963, 16'd48794});
	test_expansion(128'ha2283cee200b2356bb5b9789717580ce, {16'd59988, 16'd21437, 16'd45547, 16'd5978, 16'd30172, 16'd62782, 16'd4123, 16'd23462, 16'd1248, 16'd35398, 16'd20728, 16'd49589, 16'd54552, 16'd14052, 16'd28262, 16'd62404, 16'd65, 16'd33411, 16'd22777, 16'd4337, 16'd15805, 16'd55156, 16'd30990, 16'd23838, 16'd39473, 16'd58630});
	test_expansion(128'h041732f03ab273e42075c963cb906ee9, {16'd48932, 16'd56824, 16'd4338, 16'd41326, 16'd21483, 16'd27216, 16'd13999, 16'd42946, 16'd61116, 16'd39646, 16'd2627, 16'd44784, 16'd56087, 16'd20177, 16'd14687, 16'd52349, 16'd39155, 16'd5985, 16'd41514, 16'd28651, 16'd54742, 16'd57352, 16'd46962, 16'd47655, 16'd31958, 16'd4094});
	test_expansion(128'h47287041f6f22034a8ab839b608fa01e, {16'd23758, 16'd17820, 16'd11063, 16'd17022, 16'd42804, 16'd63694, 16'd43157, 16'd54977, 16'd1657, 16'd1173, 16'd38432, 16'd38274, 16'd54245, 16'd18672, 16'd47772, 16'd57055, 16'd45750, 16'd39358, 16'd20954, 16'd39013, 16'd9322, 16'd5983, 16'd47669, 16'd30100, 16'd32544, 16'd864});
	test_expansion(128'ha3e74c5422e4fd4058f6f1b4f3fbd3f3, {16'd59634, 16'd15945, 16'd47647, 16'd46583, 16'd12020, 16'd41887, 16'd13094, 16'd30539, 16'd14977, 16'd61421, 16'd42352, 16'd54726, 16'd14628, 16'd46669, 16'd23713, 16'd41076, 16'd6698, 16'd19940, 16'd54221, 16'd19409, 16'd5327, 16'd1611, 16'd51766, 16'd7850, 16'd7994, 16'd32173});
	test_expansion(128'h5dd3db7612ce4d0a9eb295160e8923aa, {16'd64989, 16'd34815, 16'd1997, 16'd3607, 16'd11499, 16'd20648, 16'd45221, 16'd27385, 16'd47479, 16'd35327, 16'd37961, 16'd54966, 16'd9293, 16'd25665, 16'd26881, 16'd25291, 16'd35449, 16'd42805, 16'd54926, 16'd60751, 16'd17733, 16'd14635, 16'd45577, 16'd15065, 16'd28595, 16'd57059});
	test_expansion(128'h2c4e2691779e6c20e3f50fd6997124b3, {16'd57267, 16'd65413, 16'd61798, 16'd12612, 16'd38069, 16'd2335, 16'd55169, 16'd13220, 16'd59769, 16'd44794, 16'd41385, 16'd36820, 16'd4683, 16'd58196, 16'd25143, 16'd61971, 16'd65455, 16'd64939, 16'd62773, 16'd1755, 16'd19645, 16'd29765, 16'd40432, 16'd41470, 16'd37039, 16'd12334});
	test_expansion(128'h5267264579874b3b48c805fdfe5cbfe8, {16'd17195, 16'd43210, 16'd29146, 16'd37955, 16'd11292, 16'd16868, 16'd17969, 16'd58753, 16'd23828, 16'd50155, 16'd17509, 16'd65180, 16'd46351, 16'd55303, 16'd39965, 16'd30372, 16'd13940, 16'd64516, 16'd47815, 16'd42583, 16'd45692, 16'd39704, 16'd5572, 16'd33259, 16'd249, 16'd29070});
	test_expansion(128'h32dc6479c08615af0e3e5a1db2dd3ed0, {16'd64184, 16'd23642, 16'd36998, 16'd31625, 16'd31359, 16'd36738, 16'd48930, 16'd36880, 16'd33215, 16'd51421, 16'd34735, 16'd36527, 16'd3742, 16'd60811, 16'd49706, 16'd20793, 16'd53870, 16'd29511, 16'd27645, 16'd5321, 16'd36086, 16'd40823, 16'd13402, 16'd58473, 16'd17067, 16'd56223});
	test_expansion(128'h60e3eb86b6817ecac52f7a501c76f4df, {16'd16589, 16'd2053, 16'd35263, 16'd58692, 16'd2193, 16'd5046, 16'd59528, 16'd55086, 16'd16380, 16'd57804, 16'd16475, 16'd27770, 16'd49718, 16'd47752, 16'd16498, 16'd14562, 16'd47734, 16'd19423, 16'd47066, 16'd4152, 16'd5750, 16'd61640, 16'd12898, 16'd64565, 16'd38559, 16'd34078});
	test_expansion(128'hc4d299bc42b91230c3735df9eb6fc974, {16'd26491, 16'd22924, 16'd48085, 16'd5707, 16'd2907, 16'd8100, 16'd59463, 16'd25784, 16'd41828, 16'd13484, 16'd63931, 16'd3862, 16'd2181, 16'd18302, 16'd1348, 16'd45197, 16'd11801, 16'd26229, 16'd7444, 16'd12197, 16'd33755, 16'd24746, 16'd60646, 16'd16787, 16'd42463, 16'd42372});
	test_expansion(128'hbf8f1b7426df49a97660c922c989da23, {16'd37207, 16'd23626, 16'd52650, 16'd45449, 16'd39252, 16'd27221, 16'd16147, 16'd51790, 16'd4797, 16'd2941, 16'd49112, 16'd7808, 16'd8131, 16'd7559, 16'd7518, 16'd64246, 16'd29944, 16'd45894, 16'd30406, 16'd33646, 16'd24199, 16'd10560, 16'd49415, 16'd30256, 16'd30665, 16'd43929});
	test_expansion(128'h6f156c58dc1ccf36339395dfaf55e244, {16'd13096, 16'd50315, 16'd21534, 16'd47570, 16'd38599, 16'd24731, 16'd50755, 16'd14561, 16'd30909, 16'd34622, 16'd43224, 16'd9213, 16'd30950, 16'd13748, 16'd31744, 16'd20290, 16'd30581, 16'd11763, 16'd11431, 16'd40185, 16'd55162, 16'd61859, 16'd59727, 16'd3656, 16'd22279, 16'd17289});
	test_expansion(128'h9e7e792fb38976262019c2764a4167f7, {16'd40627, 16'd22928, 16'd55184, 16'd62994, 16'd28256, 16'd14622, 16'd27074, 16'd30760, 16'd50644, 16'd23563, 16'd61962, 16'd59841, 16'd56044, 16'd65214, 16'd12125, 16'd39214, 16'd61639, 16'd50120, 16'd12821, 16'd21403, 16'd40301, 16'd31132, 16'd28378, 16'd57885, 16'd64501, 16'd49141});
	test_expansion(128'h2c346abc6080733d3c84f71cdfd52719, {16'd7925, 16'd5186, 16'd15165, 16'd12917, 16'd56206, 16'd4115, 16'd52180, 16'd55489, 16'd11628, 16'd16992, 16'd10268, 16'd63223, 16'd45027, 16'd64970, 16'd58195, 16'd867, 16'd31219, 16'd9500, 16'd11626, 16'd26609, 16'd14870, 16'd15546, 16'd56967, 16'd5864, 16'd16118, 16'd13254});
	test_expansion(128'h50e7a06a05cbd0e9c0f06daba5936d64, {16'd36549, 16'd38537, 16'd41585, 16'd8345, 16'd54384, 16'd16300, 16'd18525, 16'd62958, 16'd8303, 16'd48459, 16'd54160, 16'd56240, 16'd13534, 16'd3159, 16'd61502, 16'd23251, 16'd17646, 16'd7215, 16'd28230, 16'd30471, 16'd41936, 16'd37552, 16'd58458, 16'd34038, 16'd18406, 16'd43960});
	test_expansion(128'h1f45c80d0f74854d937b4153e1b7d874, {16'd19974, 16'd12388, 16'd39643, 16'd33202, 16'd42181, 16'd63148, 16'd32849, 16'd35245, 16'd13979, 16'd44266, 16'd38512, 16'd12946, 16'd12077, 16'd51387, 16'd64382, 16'd64129, 16'd51858, 16'd5069, 16'd52749, 16'd24994, 16'd49708, 16'd37638, 16'd42001, 16'd28079, 16'd33647, 16'd57215});
	test_expansion(128'hf88dacf5247870eab03478aa41250786, {16'd32835, 16'd9978, 16'd16414, 16'd61205, 16'd46856, 16'd63225, 16'd40061, 16'd54451, 16'd22403, 16'd33008, 16'd39158, 16'd22909, 16'd33928, 16'd62971, 16'd41413, 16'd7110, 16'd29553, 16'd52287, 16'd49378, 16'd24179, 16'd12719, 16'd13988, 16'd48918, 16'd5049, 16'd38091, 16'd22615});
	test_expansion(128'h3d1006a4b2a94f04bd7fd4f55956c08f, {16'd46877, 16'd3392, 16'd3650, 16'd65135, 16'd56728, 16'd11355, 16'd53373, 16'd55008, 16'd61907, 16'd63097, 16'd15310, 16'd38697, 16'd64731, 16'd43586, 16'd32264, 16'd54244, 16'd20898, 16'd15209, 16'd22572, 16'd44794, 16'd5299, 16'd23710, 16'd61762, 16'd12983, 16'd35088, 16'd38846});
	test_expansion(128'hd25ffecfa51ec2413ecc2d8f6b80dcec, {16'd7977, 16'd65051, 16'd16322, 16'd57551, 16'd14579, 16'd15434, 16'd44741, 16'd7184, 16'd19342, 16'd54697, 16'd5139, 16'd18687, 16'd29645, 16'd1667, 16'd50089, 16'd47532, 16'd21999, 16'd40203, 16'd28795, 16'd62434, 16'd5681, 16'd56908, 16'd8422, 16'd39899, 16'd632, 16'd43406});
	test_expansion(128'h51a6d5f0e593b6c1e9c5e119ce7b7640, {16'd18350, 16'd45546, 16'd64435, 16'd14991, 16'd29137, 16'd46478, 16'd29932, 16'd41294, 16'd12203, 16'd54228, 16'd37854, 16'd41884, 16'd2324, 16'd6392, 16'd37016, 16'd38166, 16'd21797, 16'd8729, 16'd360, 16'd10760, 16'd16577, 16'd5763, 16'd36957, 16'd65285, 16'd37417, 16'd37055});
	test_expansion(128'hf3dbb4093ff57f147d7e3e328cc8f721, {16'd64925, 16'd31429, 16'd28063, 16'd18653, 16'd24505, 16'd13239, 16'd33708, 16'd40852, 16'd25352, 16'd53412, 16'd8608, 16'd9547, 16'd36132, 16'd10793, 16'd8124, 16'd57887, 16'd29943, 16'd9095, 16'd62788, 16'd59010, 16'd61744, 16'd64618, 16'd60022, 16'd50466, 16'd41031, 16'd20994});
	test_expansion(128'hf42129beb8e643f6c629a5d71958b463, {16'd53703, 16'd7030, 16'd37636, 16'd28268, 16'd39772, 16'd4033, 16'd9287, 16'd30872, 16'd1392, 16'd21851, 16'd3297, 16'd55072, 16'd35182, 16'd23471, 16'd46901, 16'd27196, 16'd6935, 16'd35020, 16'd33882, 16'd34868, 16'd61791, 16'd38763, 16'd14097, 16'd58607, 16'd2015, 16'd50525});
	test_expansion(128'hd075a8fa837859760f5f48fbaed9a86a, {16'd53113, 16'd19472, 16'd57623, 16'd61469, 16'd19429, 16'd4673, 16'd48541, 16'd50694, 16'd17291, 16'd2613, 16'd31865, 16'd61663, 16'd5258, 16'd49102, 16'd50861, 16'd54214, 16'd32319, 16'd50247, 16'd64195, 16'd37765, 16'd59014, 16'd4862, 16'd34047, 16'd280, 16'd42846, 16'd16725});
	test_expansion(128'h830705514e5b8ff7cd299d74dd176577, {16'd60849, 16'd24237, 16'd15656, 16'd28143, 16'd39865, 16'd37249, 16'd56945, 16'd49912, 16'd59535, 16'd13565, 16'd2657, 16'd42720, 16'd6006, 16'd60393, 16'd33710, 16'd31279, 16'd14531, 16'd58249, 16'd64898, 16'd22153, 16'd5453, 16'd50342, 16'd39543, 16'd1856, 16'd41856, 16'd18485});
	test_expansion(128'hd396f15869fc87074609ed7e2d578005, {16'd54481, 16'd40583, 16'd858, 16'd37255, 16'd40696, 16'd25505, 16'd39580, 16'd14349, 16'd10641, 16'd36775, 16'd24142, 16'd65266, 16'd21782, 16'd7689, 16'd11541, 16'd48240, 16'd60281, 16'd56723, 16'd46302, 16'd38753, 16'd18872, 16'd51407, 16'd2816, 16'd16706, 16'd64938, 16'd5042});
	test_expansion(128'h258b4dcb7123cfc345eddc394acaca75, {16'd19785, 16'd11866, 16'd62203, 16'd30626, 16'd53016, 16'd60229, 16'd32359, 16'd30604, 16'd42968, 16'd26549, 16'd7102, 16'd45162, 16'd14801, 16'd21082, 16'd19468, 16'd28941, 16'd11147, 16'd64805, 16'd56532, 16'd16903, 16'd46329, 16'd45617, 16'd20879, 16'd33793, 16'd54286, 16'd34482});
	test_expansion(128'hb8202d40e3bec06d1c1270cf337bc49c, {16'd11559, 16'd2628, 16'd60470, 16'd37855, 16'd45166, 16'd18165, 16'd61943, 16'd25645, 16'd46930, 16'd1113, 16'd19574, 16'd46069, 16'd10059, 16'd25840, 16'd59691, 16'd47863, 16'd37090, 16'd22338, 16'd55538, 16'd46851, 16'd53201, 16'd18559, 16'd29082, 16'd10276, 16'd63158, 16'd27861});
	test_expansion(128'h43991b17e05cde53813f1ba0990c49cb, {16'd58058, 16'd50493, 16'd44921, 16'd51019, 16'd31551, 16'd12805, 16'd28551, 16'd51830, 16'd3938, 16'd38438, 16'd31709, 16'd47688, 16'd33841, 16'd57004, 16'd2257, 16'd11569, 16'd7998, 16'd20200, 16'd56045, 16'd61619, 16'd53038, 16'd27974, 16'd20392, 16'd1548, 16'd31077, 16'd21093});
	test_expansion(128'h9ee8bfa76e7ec238b47215d427ea083c, {16'd22800, 16'd59160, 16'd22427, 16'd36469, 16'd46664, 16'd15058, 16'd8112, 16'd29816, 16'd3988, 16'd17594, 16'd63346, 16'd64399, 16'd46672, 16'd53491, 16'd60684, 16'd50339, 16'd38341, 16'd2229, 16'd36248, 16'd3714, 16'd18068, 16'd8676, 16'd41317, 16'd19254, 16'd48956, 16'd61348});
	test_expansion(128'h4d149a6f231b66eeec0b651330d5ceb9, {16'd12381, 16'd1322, 16'd21031, 16'd34722, 16'd24486, 16'd17096, 16'd60556, 16'd24473, 16'd34651, 16'd14509, 16'd33843, 16'd49647, 16'd46441, 16'd61461, 16'd13114, 16'd52982, 16'd63769, 16'd52165, 16'd55329, 16'd58778, 16'd58424, 16'd9214, 16'd38670, 16'd34328, 16'd64704, 16'd30217});
	test_expansion(128'hab5df2c5f4daf37f21a413a5fb5ce249, {16'd37824, 16'd5632, 16'd42978, 16'd44553, 16'd2478, 16'd5486, 16'd63226, 16'd15362, 16'd10803, 16'd40435, 16'd47591, 16'd52399, 16'd38275, 16'd38659, 16'd22781, 16'd29373, 16'd30851, 16'd22394, 16'd7862, 16'd9919, 16'd34562, 16'd1126, 16'd1997, 16'd51879, 16'd18056, 16'd13183});
	test_expansion(128'h2fc60464325f6cec0b40b520ea27cbe0, {16'd61210, 16'd3738, 16'd12230, 16'd11435, 16'd21221, 16'd58541, 16'd9083, 16'd38224, 16'd24298, 16'd13810, 16'd58125, 16'd59938, 16'd45353, 16'd63623, 16'd14325, 16'd57199, 16'd47193, 16'd10909, 16'd62668, 16'd12120, 16'd11286, 16'd11636, 16'd9908, 16'd51793, 16'd61180, 16'd3177});
	test_expansion(128'hee125bdb44581e6ea385024ec1d20dd2, {16'd14030, 16'd30686, 16'd10127, 16'd4121, 16'd27583, 16'd55520, 16'd20641, 16'd1999, 16'd6768, 16'd52419, 16'd11658, 16'd30836, 16'd60223, 16'd16246, 16'd41566, 16'd12034, 16'd32226, 16'd17755, 16'd28851, 16'd37601, 16'd50853, 16'd14602, 16'd36632, 16'd50604, 16'd21442, 16'd58204});
	test_expansion(128'hafa4719dfd1dbb988ae602beef0919aa, {16'd63584, 16'd52079, 16'd19394, 16'd12295, 16'd20070, 16'd56864, 16'd55905, 16'd26450, 16'd13129, 16'd38412, 16'd24791, 16'd21445, 16'd21149, 16'd21337, 16'd43619, 16'd20270, 16'd40304, 16'd21714, 16'd16864, 16'd37868, 16'd15725, 16'd2897, 16'd48020, 16'd4434, 16'd30202, 16'd30615});
	test_expansion(128'hd39415ef67df6dc7d3e783128f999503, {16'd53310, 16'd44300, 16'd6830, 16'd2833, 16'd1772, 16'd60032, 16'd9111, 16'd45839, 16'd51070, 16'd65406, 16'd33442, 16'd44432, 16'd28811, 16'd53031, 16'd17015, 16'd54893, 16'd61751, 16'd39699, 16'd56706, 16'd12402, 16'd32941, 16'd39297, 16'd6560, 16'd45879, 16'd50531, 16'd36576});
	test_expansion(128'h6a8788bea0070e98b1a966fc19cc3cf7, {16'd7919, 16'd56763, 16'd10802, 16'd60773, 16'd6218, 16'd30520, 16'd38169, 16'd5821, 16'd61184, 16'd1548, 16'd54262, 16'd19799, 16'd52230, 16'd39245, 16'd45779, 16'd9982, 16'd4082, 16'd24448, 16'd19881, 16'd63426, 16'd45077, 16'd36305, 16'd50408, 16'd15295, 16'd22861, 16'd21069});
	test_expansion(128'hb498d97ce5c8090e36e49c742cad635b, {16'd47227, 16'd39016, 16'd42704, 16'd26241, 16'd57416, 16'd24760, 16'd45344, 16'd11573, 16'd61749, 16'd28275, 16'd9347, 16'd31744, 16'd20544, 16'd58605, 16'd42093, 16'd5169, 16'd50558, 16'd58100, 16'd13585, 16'd42409, 16'd41633, 16'd34922, 16'd29348, 16'd22242, 16'd57299, 16'd9775});
	test_expansion(128'h36603d6159e45055693c97deb6aaf533, {16'd29705, 16'd10845, 16'd17994, 16'd7698, 16'd61979, 16'd3958, 16'd21399, 16'd20677, 16'd27565, 16'd58460, 16'd934, 16'd56384, 16'd27197, 16'd24897, 16'd50476, 16'd31361, 16'd16437, 16'd20784, 16'd54051, 16'd26197, 16'd46765, 16'd3010, 16'd5874, 16'd55245, 16'd24012, 16'd46674});
	test_expansion(128'h63952b5f855d3268e85c6c02face6cfe, {16'd36192, 16'd5948, 16'd26241, 16'd62974, 16'd46526, 16'd55156, 16'd14936, 16'd23122, 16'd52805, 16'd64324, 16'd36547, 16'd25469, 16'd42486, 16'd17738, 16'd8442, 16'd11505, 16'd43383, 16'd62113, 16'd47020, 16'd29221, 16'd9122, 16'd51892, 16'd33390, 16'd54784, 16'd20594, 16'd35020});
	test_expansion(128'h9da819b38b51727456f0a6d6d18dee99, {16'd42355, 16'd13245, 16'd64258, 16'd48595, 16'd44659, 16'd19599, 16'd26023, 16'd40538, 16'd62160, 16'd12425, 16'd34048, 16'd64900, 16'd19387, 16'd15837, 16'd11904, 16'd36658, 16'd38756, 16'd33423, 16'd39106, 16'd57535, 16'd40353, 16'd36512, 16'd32653, 16'd44385, 16'd29264, 16'd11682});
	test_expansion(128'hd46bd9d3de3681042b2f07315717dfee, {16'd18940, 16'd5688, 16'd788, 16'd31525, 16'd42933, 16'd54377, 16'd65184, 16'd24844, 16'd64764, 16'd59762, 16'd54077, 16'd56050, 16'd45537, 16'd54245, 16'd10928, 16'd42497, 16'd34540, 16'd25527, 16'd25991, 16'd4362, 16'd13246, 16'd60257, 16'd40640, 16'd45417, 16'd7050, 16'd25875});
	test_expansion(128'h39f51a6d734b6c36f68559fbbc553032, {16'd60799, 16'd49973, 16'd62664, 16'd41822, 16'd32178, 16'd13280, 16'd14702, 16'd51765, 16'd33731, 16'd53319, 16'd11992, 16'd61331, 16'd73, 16'd7626, 16'd49392, 16'd51130, 16'd8783, 16'd24951, 16'd62403, 16'd9663, 16'd55410, 16'd49505, 16'd12989, 16'd32738, 16'd47854, 16'd45221});
	test_expansion(128'hebb7b92bb35a6d016f6583f7767077f3, {16'd35277, 16'd7252, 16'd48823, 16'd60017, 16'd50797, 16'd59624, 16'd62720, 16'd54570, 16'd24301, 16'd24507, 16'd45257, 16'd16409, 16'd7959, 16'd37359, 16'd41688, 16'd29155, 16'd46949, 16'd20817, 16'd3812, 16'd58431, 16'd8841, 16'd44089, 16'd10094, 16'd38025, 16'd47806, 16'd61197});
	test_expansion(128'h14237b49cf652d3d264f1c01eb9ae898, {16'd766, 16'd19136, 16'd5314, 16'd28609, 16'd6098, 16'd32381, 16'd31689, 16'd64812, 16'd56196, 16'd47350, 16'd37197, 16'd53170, 16'd12073, 16'd33732, 16'd38700, 16'd20650, 16'd61073, 16'd32511, 16'd63023, 16'd42414, 16'd62124, 16'd56945, 16'd41925, 16'd40970, 16'd21258, 16'd58515});
	test_expansion(128'h22b228006611de3aad7a0dc90e1455b3, {16'd39454, 16'd2352, 16'd14798, 16'd64214, 16'd18214, 16'd17038, 16'd47825, 16'd25873, 16'd2327, 16'd56368, 16'd11395, 16'd24086, 16'd5612, 16'd20114, 16'd46194, 16'd26852, 16'd12274, 16'd54317, 16'd18466, 16'd3881, 16'd17721, 16'd10354, 16'd15699, 16'd41723, 16'd54456, 16'd16432});
	test_expansion(128'h752efb35493717330c084e2ef42b499b, {16'd10922, 16'd62755, 16'd42497, 16'd9630, 16'd15910, 16'd25527, 16'd13533, 16'd32816, 16'd31894, 16'd3533, 16'd6160, 16'd26477, 16'd51608, 16'd57756, 16'd27544, 16'd29720, 16'd11818, 16'd9129, 16'd16313, 16'd29443, 16'd3876, 16'd5172, 16'd201, 16'd24643, 16'd55636, 16'd5579});
	test_expansion(128'hb4c6b076c31bea43f37e4e942518cbfd, {16'd6900, 16'd279, 16'd24425, 16'd47225, 16'd37971, 16'd1067, 16'd23644, 16'd26414, 16'd7436, 16'd12418, 16'd8480, 16'd6196, 16'd51888, 16'd54632, 16'd56266, 16'd7683, 16'd54865, 16'd20614, 16'd27673, 16'd63522, 16'd41982, 16'd27059, 16'd47753, 16'd59277, 16'd64226, 16'd28445});
	test_expansion(128'hdbc49166ba927661506e6e85bf51cc14, {16'd44039, 16'd37495, 16'd50464, 16'd24409, 16'd54452, 16'd38212, 16'd39123, 16'd15092, 16'd35023, 16'd48086, 16'd2463, 16'd18244, 16'd40880, 16'd53459, 16'd518, 16'd3803, 16'd10885, 16'd57509, 16'd56204, 16'd50270, 16'd10087, 16'd45157, 16'd52194, 16'd22119, 16'd26046, 16'd29492});
	test_expansion(128'hf8d60c3675425f59244cd018fb7bd6f9, {16'd16174, 16'd13791, 16'd19238, 16'd43192, 16'd19830, 16'd40005, 16'd19591, 16'd39320, 16'd61782, 16'd21536, 16'd51194, 16'd44854, 16'd22135, 16'd29710, 16'd59079, 16'd57853, 16'd60901, 16'd18277, 16'd50895, 16'd23573, 16'd9915, 16'd6218, 16'd6963, 16'd19875, 16'd58421, 16'd60357});
	test_expansion(128'h08edb1be6ef29ba955a1ed61cc554f18, {16'd38712, 16'd546, 16'd22835, 16'd63368, 16'd25845, 16'd31158, 16'd21951, 16'd52857, 16'd39423, 16'd61907, 16'd56827, 16'd57213, 16'd49846, 16'd17243, 16'd19301, 16'd23604, 16'd34578, 16'd44898, 16'd29807, 16'd33958, 16'd55702, 16'd64196, 16'd25010, 16'd38411, 16'd13159, 16'd12522});
	test_expansion(128'h106fcabe9566ed423baec78a52f4187e, {16'd27466, 16'd2334, 16'd46755, 16'd44675, 16'd16974, 16'd18314, 16'd22090, 16'd47, 16'd533, 16'd57779, 16'd34396, 16'd28605, 16'd63724, 16'd21967, 16'd32421, 16'd34714, 16'd39682, 16'd65469, 16'd5351, 16'd41853, 16'd19898, 16'd44164, 16'd3529, 16'd21863, 16'd23756, 16'd17167});
	test_expansion(128'h02ffab7e1ddfe9df78a241ccc9aec320, {16'd17491, 16'd63108, 16'd14002, 16'd39713, 16'd25325, 16'd24792, 16'd7861, 16'd21464, 16'd30940, 16'd13580, 16'd13381, 16'd59805, 16'd9764, 16'd51210, 16'd40389, 16'd26818, 16'd50733, 16'd27820, 16'd50047, 16'd31828, 16'd59712, 16'd26585, 16'd41194, 16'd57591, 16'd4705, 16'd21227});
	test_expansion(128'hfa4f1639da042afe7f2b93cd2af750e7, {16'd24655, 16'd6782, 16'd57460, 16'd11283, 16'd47460, 16'd30536, 16'd58260, 16'd10555, 16'd63275, 16'd32446, 16'd13400, 16'd27798, 16'd13344, 16'd37154, 16'd40908, 16'd37175, 16'd22683, 16'd34196, 16'd50885, 16'd27217, 16'd15216, 16'd981, 16'd49978, 16'd56223, 16'd17800, 16'd23487});
	test_expansion(128'hede66a46a9fe49341f81099c5087ebf0, {16'd6523, 16'd10677, 16'd8593, 16'd32013, 16'd39387, 16'd19278, 16'd53647, 16'd26611, 16'd46086, 16'd4780, 16'd21220, 16'd59710, 16'd61206, 16'd39227, 16'd4320, 16'd5022, 16'd32024, 16'd22149, 16'd26951, 16'd46166, 16'd34683, 16'd10967, 16'd7444, 16'd24985, 16'd51146, 16'd28520});
	test_expansion(128'hc6e1638e05ec135e0a5dc5a99540652e, {16'd45205, 16'd21628, 16'd1413, 16'd122, 16'd45823, 16'd63483, 16'd61318, 16'd11622, 16'd9698, 16'd35930, 16'd43124, 16'd45617, 16'd5274, 16'd16183, 16'd57028, 16'd61863, 16'd21946, 16'd34646, 16'd26321, 16'd1264, 16'd43468, 16'd65362, 16'd42148, 16'd19494, 16'd44233, 16'd63817});
	test_expansion(128'ha282c54bc871842a2c5c92a7cc17dd48, {16'd39075, 16'd37141, 16'd37273, 16'd54281, 16'd48014, 16'd60704, 16'd31476, 16'd26222, 16'd18227, 16'd48941, 16'd2694, 16'd29230, 16'd49816, 16'd52086, 16'd33417, 16'd57779, 16'd43705, 16'd25370, 16'd3764, 16'd30093, 16'd24361, 16'd60705, 16'd63664, 16'd16679, 16'd35550, 16'd52673});
	test_expansion(128'h57238a48b1bc4c86eb05444da75969ea, {16'd12858, 16'd20267, 16'd35719, 16'd13113, 16'd21125, 16'd8594, 16'd10169, 16'd29961, 16'd56353, 16'd32808, 16'd49307, 16'd18816, 16'd45097, 16'd38372, 16'd39189, 16'd36334, 16'd5869, 16'd16127, 16'd54527, 16'd48492, 16'd7897, 16'd17475, 16'd589, 16'd43579, 16'd19216, 16'd51405});
	test_expansion(128'h2ef54d0f492a356b608b74d6fcf7017b, {16'd52001, 16'd22559, 16'd9771, 16'd42581, 16'd12901, 16'd6529, 16'd62401, 16'd38363, 16'd20069, 16'd12403, 16'd63347, 16'd6456, 16'd63794, 16'd6281, 16'd43106, 16'd46694, 16'd47869, 16'd16643, 16'd31677, 16'd3664, 16'd49291, 16'd63902, 16'd59828, 16'd28322, 16'd13972, 16'd64567});
	test_expansion(128'h745caff577a6bbec6600b874d2dadd01, {16'd54220, 16'd45387, 16'd3146, 16'd19728, 16'd44436, 16'd21441, 16'd35937, 16'd11314, 16'd19218, 16'd31016, 16'd47676, 16'd57572, 16'd62991, 16'd54989, 16'd9461, 16'd57375, 16'd22641, 16'd27838, 16'd41102, 16'd30314, 16'd61298, 16'd31981, 16'd53344, 16'd5878, 16'd40705, 16'd60722});
	test_expansion(128'he4f6a9e0ae97e518fb613ce1af2b5540, {16'd13594, 16'd43106, 16'd13104, 16'd52985, 16'd8832, 16'd40697, 16'd1632, 16'd22643, 16'd29729, 16'd46990, 16'd5535, 16'd10315, 16'd51824, 16'd39609, 16'd2451, 16'd43610, 16'd51724, 16'd26961, 16'd51076, 16'd6518, 16'd65303, 16'd32733, 16'd46621, 16'd41331, 16'd59918, 16'd57399});
	test_expansion(128'hebf7812c71fe1812c1e2d4b24a278174, {16'd12936, 16'd39662, 16'd25594, 16'd48531, 16'd62540, 16'd60601, 16'd51349, 16'd47292, 16'd7805, 16'd41697, 16'd13921, 16'd57912, 16'd24883, 16'd54357, 16'd37942, 16'd18704, 16'd46103, 16'd22856, 16'd23461, 16'd25095, 16'd34851, 16'd55205, 16'd1533, 16'd32169, 16'd54813, 16'd9472});
	test_expansion(128'h6316bd59df200f2e9953993efa9a3f0b, {16'd56917, 16'd47810, 16'd55260, 16'd27346, 16'd44358, 16'd20917, 16'd53698, 16'd55071, 16'd54234, 16'd59778, 16'd16439, 16'd31486, 16'd46081, 16'd62321, 16'd51566, 16'd58935, 16'd52129, 16'd48984, 16'd59639, 16'd57862, 16'd56161, 16'd50029, 16'd57034, 16'd44850, 16'd2848, 16'd63431});
	test_expansion(128'h4c41eb8f320a908bc7c3f417427cfd3b, {16'd54407, 16'd65082, 16'd64219, 16'd33362, 16'd36684, 16'd45514, 16'd49134, 16'd26370, 16'd14159, 16'd6756, 16'd41531, 16'd21712, 16'd7088, 16'd32908, 16'd63293, 16'd62348, 16'd11453, 16'd51928, 16'd2648, 16'd24118, 16'd10686, 16'd26380, 16'd48228, 16'd65072, 16'd43990, 16'd22374});
	test_expansion(128'hd49e7ba9c4dca0d987a42f5668f2bb4f, {16'd4030, 16'd26831, 16'd53604, 16'd43433, 16'd2361, 16'd65082, 16'd22776, 16'd32810, 16'd14729, 16'd63988, 16'd50447, 16'd17399, 16'd654, 16'd1956, 16'd33868, 16'd42259, 16'd48317, 16'd12286, 16'd4034, 16'd51753, 16'd38367, 16'd35801, 16'd46638, 16'd37173, 16'd20440, 16'd43677});
	test_expansion(128'h1d43b5c1c674d138cad435e309921709, {16'd23268, 16'd35365, 16'd33460, 16'd61611, 16'd26435, 16'd50582, 16'd53882, 16'd14309, 16'd19816, 16'd41875, 16'd60622, 16'd3142, 16'd38501, 16'd12925, 16'd24620, 16'd32507, 16'd60256, 16'd62606, 16'd3787, 16'd8183, 16'd7461, 16'd4066, 16'd39611, 16'd5757, 16'd55032, 16'd55636});
	test_expansion(128'haaf871d953c8baaa3b211fab3064560d, {16'd27160, 16'd47225, 16'd41372, 16'd4550, 16'd46298, 16'd11684, 16'd38751, 16'd25158, 16'd22718, 16'd28287, 16'd12177, 16'd15495, 16'd64037, 16'd54529, 16'd44654, 16'd38022, 16'd38444, 16'd34823, 16'd63551, 16'd27412, 16'd16623, 16'd4021, 16'd59260, 16'd29382, 16'd8509, 16'd18896});
	test_expansion(128'h5d5026cc67ff3c2cd85ffb7283df008b, {16'd4366, 16'd18729, 16'd10694, 16'd59236, 16'd24453, 16'd57892, 16'd35160, 16'd50296, 16'd8936, 16'd53232, 16'd51571, 16'd55929, 16'd22572, 16'd24479, 16'd4220, 16'd57585, 16'd27982, 16'd51381, 16'd51438, 16'd62043, 16'd1834, 16'd41607, 16'd51593, 16'd54267, 16'd23212, 16'd34722});
	test_expansion(128'hcab36421bb226ad0f4ff5ae165b13196, {16'd51055, 16'd41842, 16'd4867, 16'd58948, 16'd12000, 16'd21330, 16'd28322, 16'd58138, 16'd30484, 16'd32917, 16'd24368, 16'd27752, 16'd55447, 16'd62481, 16'd34149, 16'd48634, 16'd38369, 16'd2049, 16'd52314, 16'd3220, 16'd22759, 16'd23635, 16'd1135, 16'd56844, 16'd22158, 16'd63532});
	test_expansion(128'h4a680bfbeb05c26970b8c23f757a573c, {16'd51494, 16'd41098, 16'd64793, 16'd38233, 16'd9059, 16'd35263, 16'd37336, 16'd46367, 16'd11118, 16'd48885, 16'd27651, 16'd55628, 16'd39266, 16'd12105, 16'd56711, 16'd36873, 16'd23305, 16'd43921, 16'd56709, 16'd53167, 16'd63925, 16'd30031, 16'd685, 16'd53240, 16'd37930, 16'd25002});
	test_expansion(128'hab14951100fb3276b4d7d4e2564b642e, {16'd1155, 16'd45569, 16'd65105, 16'd18713, 16'd45157, 16'd10491, 16'd13152, 16'd19017, 16'd30275, 16'd18666, 16'd20962, 16'd5787, 16'd62647, 16'd36222, 16'd52802, 16'd38940, 16'd36755, 16'd20281, 16'd5890, 16'd39885, 16'd32299, 16'd37845, 16'd25912, 16'd52776, 16'd28076, 16'd50764});
	test_expansion(128'h67e67ec0df259729e49313343b8125a3, {16'd42778, 16'd26976, 16'd58878, 16'd51299, 16'd15916, 16'd4244, 16'd19773, 16'd47773, 16'd21220, 16'd28714, 16'd19155, 16'd45601, 16'd39985, 16'd14098, 16'd45324, 16'd20008, 16'd12311, 16'd620, 16'd13025, 16'd46496, 16'd15434, 16'd35010, 16'd19405, 16'd44087, 16'd54908, 16'd53621});
	test_expansion(128'h0f5a7ee87eb8a004ea5f345c3e09ae95, {16'd29170, 16'd47490, 16'd34594, 16'd15989, 16'd31211, 16'd11656, 16'd41071, 16'd6146, 16'd33935, 16'd2878, 16'd47671, 16'd54699, 16'd32735, 16'd9412, 16'd20761, 16'd30634, 16'd23163, 16'd5030, 16'd15330, 16'd64069, 16'd30856, 16'd34057, 16'd36598, 16'd55541, 16'd18153, 16'd2731});
	test_expansion(128'h5b658f91e43238266f8039b716781e2d, {16'd33147, 16'd44158, 16'd29643, 16'd21409, 16'd57927, 16'd39239, 16'd25621, 16'd22007, 16'd20913, 16'd61886, 16'd19317, 16'd65272, 16'd22886, 16'd43709, 16'd60476, 16'd38272, 16'd35853, 16'd42540, 16'd62808, 16'd50245, 16'd46260, 16'd10125, 16'd17847, 16'd42680, 16'd44278, 16'd36800});
	test_expansion(128'h5769cff45f7c62e984292b26b6c6c1c7, {16'd41942, 16'd43164, 16'd36550, 16'd41696, 16'd63578, 16'd15545, 16'd9384, 16'd56871, 16'd51733, 16'd50216, 16'd28575, 16'd64151, 16'd37050, 16'd28329, 16'd49282, 16'd8464, 16'd8236, 16'd51596, 16'd32964, 16'd43441, 16'd5273, 16'd19796, 16'd65145, 16'd44304, 16'd17688, 16'd55010});
	test_expansion(128'hfc3b0ecab3c8b598eade83b604993e77, {16'd20488, 16'd40915, 16'd43501, 16'd52853, 16'd16931, 16'd52715, 16'd10521, 16'd43371, 16'd11344, 16'd11288, 16'd37505, 16'd44297, 16'd26030, 16'd35776, 16'd56988, 16'd13877, 16'd44770, 16'd12402, 16'd53955, 16'd43976, 16'd17928, 16'd28899, 16'd2745, 16'd4237, 16'd887, 16'd1553});
	test_expansion(128'h55fe7da0a0890e8b75972365ae1b7909, {16'd20904, 16'd43936, 16'd11657, 16'd41200, 16'd20448, 16'd12159, 16'd5644, 16'd51101, 16'd22056, 16'd32071, 16'd12580, 16'd31814, 16'd32097, 16'd6032, 16'd42273, 16'd32721, 16'd36701, 16'd57798, 16'd29988, 16'd11571, 16'd1843, 16'd33878, 16'd4057, 16'd18594, 16'd2107, 16'd32696});
	test_expansion(128'hbce94ac2315fb3dde096a15c526bdfce, {16'd24741, 16'd16056, 16'd13146, 16'd15217, 16'd40658, 16'd25870, 16'd41268, 16'd32671, 16'd30827, 16'd34201, 16'd56166, 16'd1918, 16'd19317, 16'd24294, 16'd24966, 16'd13649, 16'd59552, 16'd52483, 16'd24844, 16'd14059, 16'd272, 16'd19309, 16'd10543, 16'd58423, 16'd5276, 16'd41179});
	test_expansion(128'hb0ee3f5e069000406da40d5277faf3f2, {16'd49772, 16'd47202, 16'd58262, 16'd6331, 16'd39175, 16'd52930, 16'd3206, 16'd9047, 16'd50234, 16'd46939, 16'd62113, 16'd36694, 16'd18992, 16'd26608, 16'd62107, 16'd53375, 16'd58710, 16'd3375, 16'd55899, 16'd20303, 16'd62800, 16'd50689, 16'd17648, 16'd32968, 16'd2457, 16'd9438});
	test_expansion(128'hb2151a314a56dd9b10a00b386e3d7e4f, {16'd34990, 16'd25507, 16'd17226, 16'd54338, 16'd43840, 16'd56467, 16'd26178, 16'd37950, 16'd9092, 16'd6696, 16'd46423, 16'd49611, 16'd39887, 16'd41985, 16'd34435, 16'd61458, 16'd57931, 16'd18635, 16'd40302, 16'd60138, 16'd55690, 16'd48904, 16'd14305, 16'd16576, 16'd17648, 16'd42696});
	test_expansion(128'h0f5729558de6ecc4a1abf3e73be92d6c, {16'd29977, 16'd16621, 16'd62038, 16'd44602, 16'd4259, 16'd46208, 16'd60635, 16'd10777, 16'd37964, 16'd1248, 16'd52476, 16'd30181, 16'd43167, 16'd60796, 16'd38003, 16'd21194, 16'd64757, 16'd61954, 16'd59095, 16'd63367, 16'd7556, 16'd17997, 16'd13043, 16'd3156, 16'd14385, 16'd10206});
	test_expansion(128'hbe395b5a85c418fd85185fa934a3a484, {16'd47152, 16'd62500, 16'd27526, 16'd36222, 16'd9948, 16'd45160, 16'd39638, 16'd27839, 16'd28318, 16'd2271, 16'd37548, 16'd56993, 16'd6579, 16'd5394, 16'd37802, 16'd30319, 16'd2912, 16'd64263, 16'd24147, 16'd38163, 16'd63129, 16'd8760, 16'd63230, 16'd62018, 16'd30898, 16'd36040});
	test_expansion(128'h70b93a7dea90455f0e50caa74360d102, {16'd27476, 16'd15952, 16'd40764, 16'd4393, 16'd36093, 16'd44704, 16'd46414, 16'd25807, 16'd45738, 16'd23977, 16'd42359, 16'd50277, 16'd33455, 16'd46852, 16'd20057, 16'd13339, 16'd15958, 16'd36422, 16'd51850, 16'd7855, 16'd35392, 16'd1068, 16'd31817, 16'd40990, 16'd6355, 16'd26191});
	test_expansion(128'h0ecf2bac89aac9efbf2f6389ea3b71c1, {16'd10282, 16'd12848, 16'd17125, 16'd13404, 16'd56174, 16'd14065, 16'd6821, 16'd62697, 16'd4797, 16'd62329, 16'd20134, 16'd3991, 16'd30802, 16'd33141, 16'd39456, 16'd48316, 16'd61653, 16'd44732, 16'd58611, 16'd26023, 16'd61853, 16'd34633, 16'd14209, 16'd54434, 16'd1700, 16'd27585});
	test_expansion(128'h7074c52f21d0567ead8b220734ba33e7, {16'd57499, 16'd52031, 16'd17890, 16'd1654, 16'd65242, 16'd64506, 16'd62397, 16'd15470, 16'd18472, 16'd58983, 16'd41821, 16'd33175, 16'd10330, 16'd35706, 16'd10427, 16'd58942, 16'd17990, 16'd54444, 16'd6393, 16'd60623, 16'd6243, 16'd53947, 16'd11466, 16'd54391, 16'd39872, 16'd621});
	test_expansion(128'hf71a564c6f075ed75515cbce81d481be, {16'd49170, 16'd22403, 16'd47788, 16'd17614, 16'd9115, 16'd9369, 16'd2168, 16'd46979, 16'd26174, 16'd25900, 16'd38340, 16'd17791, 16'd37111, 16'd37810, 16'd61991, 16'd49181, 16'd65097, 16'd18928, 16'd52415, 16'd55155, 16'd14652, 16'd18474, 16'd21054, 16'd64210, 16'd47202, 16'd56689});
	test_expansion(128'hea8a64cd16373381fcb3d61280c3d555, {16'd52478, 16'd9941, 16'd1152, 16'd28302, 16'd56889, 16'd23305, 16'd51512, 16'd7240, 16'd13329, 16'd45834, 16'd23721, 16'd30094, 16'd49903, 16'd36093, 16'd31723, 16'd1134, 16'd63932, 16'd55227, 16'd21832, 16'd21893, 16'd61887, 16'd6879, 16'd53807, 16'd27396, 16'd4251, 16'd8605});
	test_expansion(128'h0a20e88eee71b2f16ef73e130a7f8a84, {16'd10752, 16'd62630, 16'd9067, 16'd5958, 16'd2581, 16'd14118, 16'd61702, 16'd42052, 16'd59506, 16'd58514, 16'd19654, 16'd17382, 16'd28441, 16'd749, 16'd33952, 16'd40578, 16'd59203, 16'd5842, 16'd58039, 16'd3250, 16'd26896, 16'd47468, 16'd6485, 16'd13611, 16'd45287, 16'd10444});
	test_expansion(128'h1ca6a5802f28c27ab119137ed023aca3, {16'd49666, 16'd56749, 16'd62054, 16'd63185, 16'd28212, 16'd41447, 16'd58778, 16'd50244, 16'd1536, 16'd16468, 16'd7213, 16'd58004, 16'd17358, 16'd29505, 16'd63391, 16'd28500, 16'd60644, 16'd65427, 16'd20441, 16'd50342, 16'd18017, 16'd28045, 16'd4155, 16'd31190, 16'd242, 16'd494});
	test_expansion(128'hf0c84e3c93d3b3542bc608557990f891, {16'd63282, 16'd8782, 16'd60903, 16'd17880, 16'd38827, 16'd55064, 16'd48284, 16'd59722, 16'd39465, 16'd25819, 16'd14595, 16'd50781, 16'd6962, 16'd19846, 16'd8415, 16'd61483, 16'd4519, 16'd36017, 16'd50450, 16'd48446, 16'd17668, 16'd27334, 16'd30141, 16'd18460, 16'd55079, 16'd35863});
	test_expansion(128'h411232729c25515745c940bae42f104c, {16'd53452, 16'd2572, 16'd55684, 16'd30913, 16'd42485, 16'd43821, 16'd27721, 16'd44993, 16'd30347, 16'd18202, 16'd55914, 16'd55750, 16'd39776, 16'd5061, 16'd52381, 16'd11614, 16'd2893, 16'd32039, 16'd4256, 16'd48602, 16'd52829, 16'd40339, 16'd37667, 16'd58536, 16'd40138, 16'd31159});
	test_expansion(128'h83b6b83418698383e25d064f365748c9, {16'd14876, 16'd37971, 16'd11750, 16'd63311, 16'd44313, 16'd8925, 16'd59760, 16'd4932, 16'd15691, 16'd38023, 16'd39930, 16'd52201, 16'd2994, 16'd4056, 16'd25814, 16'd8004, 16'd63000, 16'd19840, 16'd4160, 16'd59665, 16'd54848, 16'd62616, 16'd50991, 16'd7899, 16'd9614, 16'd58907});
	test_expansion(128'ha605a9b9093221f7934060a674ac893b, {16'd24539, 16'd50964, 16'd13950, 16'd8675, 16'd55691, 16'd14469, 16'd27876, 16'd29980, 16'd5434, 16'd43184, 16'd41929, 16'd41806, 16'd60921, 16'd28381, 16'd41086, 16'd58871, 16'd56554, 16'd8083, 16'd25825, 16'd43840, 16'd15532, 16'd57279, 16'd47495, 16'd44067, 16'd34566, 16'd52252});
	test_expansion(128'h2a07ba3e491ed0a4a5bebfd090599baa, {16'd61070, 16'd59940, 16'd48629, 16'd49829, 16'd39650, 16'd59519, 16'd18197, 16'd61897, 16'd14296, 16'd37367, 16'd62187, 16'd32374, 16'd41170, 16'd4105, 16'd37618, 16'd48834, 16'd50766, 16'd43904, 16'd25276, 16'd54612, 16'd1, 16'd36384, 16'd13400, 16'd1124, 16'd15920, 16'd45988});
	test_expansion(128'hfb3373a5415c05df49f1e57207323056, {16'd60087, 16'd48351, 16'd58913, 16'd54044, 16'd20435, 16'd6796, 16'd34520, 16'd50025, 16'd64364, 16'd54909, 16'd56901, 16'd35367, 16'd21795, 16'd16900, 16'd25246, 16'd61746, 16'd60636, 16'd19195, 16'd57806, 16'd45604, 16'd9661, 16'd10253, 16'd51187, 16'd59967, 16'd56464, 16'd9262});
	test_expansion(128'h80463514ccb59d58c7dc0190ceb06ca6, {16'd52074, 16'd39980, 16'd35644, 16'd31409, 16'd28470, 16'd60107, 16'd16097, 16'd59595, 16'd46912, 16'd8212, 16'd5725, 16'd32738, 16'd56916, 16'd47521, 16'd55603, 16'd2874, 16'd33964, 16'd34554, 16'd34510, 16'd47153, 16'd25112, 16'd60499, 16'd9686, 16'd6762, 16'd34878, 16'd42059});
	test_expansion(128'h31c45c16a7c1a931471f119a44efd4e5, {16'd46131, 16'd42544, 16'd6899, 16'd3786, 16'd27063, 16'd2393, 16'd60996, 16'd18779, 16'd64400, 16'd41692, 16'd36862, 16'd21313, 16'd63404, 16'd20474, 16'd1408, 16'd12814, 16'd6197, 16'd14380, 16'd36576, 16'd4956, 16'd62888, 16'd11448, 16'd58091, 16'd9522, 16'd30304, 16'd13607});
	test_expansion(128'h690eb455d1534bd5cae149a43af47240, {16'd7654, 16'd6311, 16'd30748, 16'd9527, 16'd26482, 16'd17524, 16'd17809, 16'd64806, 16'd65057, 16'd16605, 16'd40287, 16'd25399, 16'd20132, 16'd1337, 16'd9836, 16'd25542, 16'd21634, 16'd30392, 16'd11923, 16'd15087, 16'd9798, 16'd39049, 16'd54518, 16'd11573, 16'd57329, 16'd36350});
	test_expansion(128'h38956a37568badbc1f604a5263afdbd0, {16'd33511, 16'd58981, 16'd7537, 16'd36273, 16'd51910, 16'd57055, 16'd17463, 16'd33403, 16'd63872, 16'd57309, 16'd60513, 16'd7420, 16'd33390, 16'd21398, 16'd7093, 16'd41282, 16'd44454, 16'd43424, 16'd48590, 16'd25721, 16'd51297, 16'd9124, 16'd48358, 16'd64630, 16'd62323, 16'd19045});
	test_expansion(128'h29bd289b1b61a946981c31fa752ccfa4, {16'd5063, 16'd29294, 16'd43673, 16'd33566, 16'd43837, 16'd48377, 16'd20644, 16'd17579, 16'd10928, 16'd55758, 16'd28721, 16'd19679, 16'd20081, 16'd30972, 16'd47713, 16'd59190, 16'd61386, 16'd13849, 16'd23026, 16'd5528, 16'd43699, 16'd4496, 16'd8323, 16'd59982, 16'd64440, 16'd18697});
	test_expansion(128'h316f2a9d00ff50f37a18f06eeca2cd85, {16'd27788, 16'd22908, 16'd50590, 16'd55336, 16'd39580, 16'd7733, 16'd7354, 16'd15408, 16'd41873, 16'd57156, 16'd3881, 16'd61230, 16'd8102, 16'd1673, 16'd25118, 16'd53587, 16'd29059, 16'd4939, 16'd62755, 16'd8146, 16'd6328, 16'd15294, 16'd39514, 16'd48767, 16'd25038, 16'd53753});
	test_expansion(128'h6375d91758f2515c8971f2cd486f8d8d, {16'd40674, 16'd5466, 16'd20340, 16'd22313, 16'd23869, 16'd36992, 16'd28397, 16'd7607, 16'd20917, 16'd10890, 16'd20070, 16'd65028, 16'd39389, 16'd7655, 16'd62995, 16'd36951, 16'd38182, 16'd11037, 16'd12125, 16'd153, 16'd63245, 16'd34589, 16'd34917, 16'd8796, 16'd4926, 16'd62059});
	test_expansion(128'h007aab6dfa0f414d7b6b224608c85aee, {16'd47550, 16'd47295, 16'd10826, 16'd33287, 16'd59641, 16'd25450, 16'd4184, 16'd49898, 16'd50683, 16'd2237, 16'd30340, 16'd57151, 16'd19045, 16'd63722, 16'd51410, 16'd27177, 16'd24699, 16'd35070, 16'd44588, 16'd21702, 16'd11839, 16'd54790, 16'd17528, 16'd5695, 16'd23451, 16'd2262});
	test_expansion(128'h85f2e667c25391034a999d2ca3897b6e, {16'd34413, 16'd35225, 16'd1632, 16'd37005, 16'd63304, 16'd21573, 16'd26006, 16'd33336, 16'd43647, 16'd28592, 16'd51397, 16'd62467, 16'd29061, 16'd25262, 16'd41090, 16'd51600, 16'd31529, 16'd32061, 16'd9105, 16'd27850, 16'd31305, 16'd1151, 16'd1033, 16'd20787, 16'd25286, 16'd45626});
	test_expansion(128'h6156967aaed8f7445b997dd345744d58, {16'd43792, 16'd14339, 16'd21509, 16'd62198, 16'd34590, 16'd36331, 16'd2186, 16'd23888, 16'd3208, 16'd430, 16'd2477, 16'd55561, 16'd45219, 16'd8218, 16'd15874, 16'd21611, 16'd34233, 16'd38938, 16'd1471, 16'd45611, 16'd39087, 16'd61682, 16'd56249, 16'd28068, 16'd47659, 16'd60761});
	test_expansion(128'h795df76f9826140f942593bb27063702, {16'd40299, 16'd7470, 16'd12471, 16'd12290, 16'd13639, 16'd33400, 16'd2467, 16'd36652, 16'd1009, 16'd49903, 16'd39927, 16'd42731, 16'd34315, 16'd25299, 16'd6245, 16'd32044, 16'd45280, 16'd16728, 16'd48205, 16'd58896, 16'd63497, 16'd65036, 16'd41588, 16'd44814, 16'd6640, 16'd35127});
	test_expansion(128'h0b36ff75e73eb3ae061eec403e29fb10, {16'd56394, 16'd16757, 16'd52060, 16'd6534, 16'd44846, 16'd54072, 16'd40311, 16'd44988, 16'd33555, 16'd51383, 16'd18673, 16'd10969, 16'd62973, 16'd64620, 16'd10535, 16'd35757, 16'd44681, 16'd63156, 16'd50226, 16'd45260, 16'd2067, 16'd16934, 16'd54189, 16'd2016, 16'd29847, 16'd25030});
	test_expansion(128'h209a9f788edd48111cebdd194d394f16, {16'd6876, 16'd38954, 16'd47979, 16'd52096, 16'd59535, 16'd26407, 16'd42627, 16'd9646, 16'd60297, 16'd28424, 16'd57780, 16'd9443, 16'd17894, 16'd47199, 16'd34479, 16'd53056, 16'd35808, 16'd17193, 16'd64923, 16'd44730, 16'd1722, 16'd16207, 16'd52485, 16'd43363, 16'd21337, 16'd50620});
	test_expansion(128'h8a892c0cc258c57822df4ada95d75b0d, {16'd21664, 16'd2131, 16'd54530, 16'd3509, 16'd61982, 16'd33207, 16'd48167, 16'd36285, 16'd11350, 16'd55063, 16'd17017, 16'd17075, 16'd50817, 16'd39157, 16'd36373, 16'd37455, 16'd3839, 16'd51049, 16'd14888, 16'd26583, 16'd42209, 16'd11426, 16'd997, 16'd13274, 16'd402, 16'd2985});
	test_expansion(128'h4992c9513d6a01c2663c9d9f84f900f2, {16'd24257, 16'd5011, 16'd52126, 16'd4718, 16'd46370, 16'd15491, 16'd15210, 16'd15381, 16'd28328, 16'd58710, 16'd61397, 16'd33235, 16'd22388, 16'd53013, 16'd63280, 16'd32990, 16'd59443, 16'd61384, 16'd40204, 16'd4860, 16'd39387, 16'd35581, 16'd13838, 16'd40408, 16'd63292, 16'd48119});
	test_expansion(128'ha6e49ebd3b92810f4a2d1fbdb8d80ae0, {16'd8697, 16'd60249, 16'd24232, 16'd25379, 16'd17340, 16'd44772, 16'd14512, 16'd41489, 16'd49064, 16'd59113, 16'd20120, 16'd58085, 16'd52659, 16'd25711, 16'd10283, 16'd17533, 16'd62633, 16'd46356, 16'd55949, 16'd49808, 16'd52785, 16'd55473, 16'd60085, 16'd12204, 16'd33854, 16'd65431});
	test_expansion(128'h9848c12ad0751b9bbae4470eae609e13, {16'd22370, 16'd15278, 16'd34533, 16'd16891, 16'd51252, 16'd47797, 16'd959, 16'd38149, 16'd21263, 16'd14264, 16'd25758, 16'd50160, 16'd3946, 16'd61167, 16'd7527, 16'd43354, 16'd17456, 16'd27733, 16'd55585, 16'd8932, 16'd18801, 16'd28017, 16'd46985, 16'd34284, 16'd53071, 16'd51940});
	test_expansion(128'h5cb1c04fe176b442c72d484e8effccb0, {16'd37480, 16'd4038, 16'd65344, 16'd35570, 16'd34442, 16'd19502, 16'd37292, 16'd33936, 16'd12666, 16'd14200, 16'd23805, 16'd14811, 16'd14295, 16'd26557, 16'd28665, 16'd55356, 16'd62540, 16'd48727, 16'd413, 16'd53757, 16'd23485, 16'd38198, 16'd27234, 16'd21107, 16'd43667, 16'd28972});
	test_expansion(128'h6dae479e2527bf3ddadd57dec85cbaf9, {16'd37614, 16'd36523, 16'd44642, 16'd19295, 16'd60839, 16'd60389, 16'd30785, 16'd64385, 16'd31115, 16'd39545, 16'd56556, 16'd46554, 16'd14809, 16'd5427, 16'd34837, 16'd44291, 16'd46961, 16'd23008, 16'd7409, 16'd4555, 16'd16238, 16'd2478, 16'd27838, 16'd19259, 16'd51261, 16'd10530});
	test_expansion(128'h8b7e0a29f88c4f3e06307587a84020fc, {16'd56572, 16'd33825, 16'd1177, 16'd64395, 16'd770, 16'd16993, 16'd60780, 16'd10512, 16'd65175, 16'd47055, 16'd43715, 16'd42702, 16'd43944, 16'd2961, 16'd24113, 16'd20399, 16'd44973, 16'd55693, 16'd56177, 16'd17000, 16'd59138, 16'd49930, 16'd22983, 16'd10622, 16'd58629, 16'd39490});
	test_expansion(128'hd71588a0b1e7261604202c9f448ded0e, {16'd45127, 16'd26447, 16'd27054, 16'd42066, 16'd40481, 16'd36887, 16'd45749, 16'd65309, 16'd22474, 16'd43251, 16'd38187, 16'd54250, 16'd14755, 16'd33449, 16'd58161, 16'd18440, 16'd15177, 16'd22449, 16'd22010, 16'd54057, 16'd64262, 16'd33108, 16'd11126, 16'd35307, 16'd22877, 16'd50508});
	test_expansion(128'h814cb570e3c1cddf31a7c9659d08718d, {16'd30775, 16'd56692, 16'd41751, 16'd34015, 16'd28807, 16'd53633, 16'd17537, 16'd32320, 16'd51682, 16'd11477, 16'd17852, 16'd35546, 16'd64980, 16'd54363, 16'd56900, 16'd64019, 16'd10415, 16'd34579, 16'd18880, 16'd5019, 16'd13523, 16'd225, 16'd7360, 16'd65289, 16'd64459, 16'd33760});
	test_expansion(128'h788d10da036c89246afab78e386d0fb6, {16'd25209, 16'd33337, 16'd7727, 16'd16757, 16'd63769, 16'd19594, 16'd9866, 16'd277, 16'd41818, 16'd12935, 16'd11521, 16'd63093, 16'd24629, 16'd47663, 16'd61733, 16'd717, 16'd29122, 16'd6870, 16'd7721, 16'd14788, 16'd38684, 16'd22442, 16'd39284, 16'd37869, 16'd44810, 16'd51463});
	test_expansion(128'h661d2ef94df9e173f98ae3109422b180, {16'd12054, 16'd43113, 16'd40435, 16'd64351, 16'd52887, 16'd51336, 16'd3338, 16'd9884, 16'd55841, 16'd55070, 16'd4233, 16'd55646, 16'd14184, 16'd14130, 16'd26081, 16'd31324, 16'd30232, 16'd32818, 16'd36493, 16'd45708, 16'd31654, 16'd16288, 16'd5111, 16'd40103, 16'd13074, 16'd12736});
	test_expansion(128'h3cde6d453544b0609cf22ed435516bd4, {16'd59893, 16'd22415, 16'd7998, 16'd52819, 16'd40352, 16'd43096, 16'd54445, 16'd44831, 16'd46698, 16'd53190, 16'd27215, 16'd20024, 16'd56408, 16'd43777, 16'd35740, 16'd45283, 16'd12978, 16'd40029, 16'd35849, 16'd52305, 16'd6262, 16'd22549, 16'd20834, 16'd25019, 16'd57787, 16'd20486});
	test_expansion(128'h268d9cf804517ef5ab247fc3d1aae819, {16'd20591, 16'd6465, 16'd33605, 16'd1198, 16'd39770, 16'd11797, 16'd26505, 16'd56859, 16'd21676, 16'd15184, 16'd20206, 16'd48043, 16'd31855, 16'd41351, 16'd10739, 16'd60141, 16'd8059, 16'd17777, 16'd27197, 16'd34466, 16'd39522, 16'd17994, 16'd38300, 16'd20973, 16'd62181, 16'd40516});
	test_expansion(128'hdf1764a85cdcc560cbb1679274cd5af7, {16'd35871, 16'd13506, 16'd41538, 16'd34569, 16'd25429, 16'd30005, 16'd7980, 16'd8525, 16'd58736, 16'd47690, 16'd62785, 16'd55007, 16'd6650, 16'd52310, 16'd40347, 16'd35175, 16'd56921, 16'd43821, 16'd20173, 16'd30570, 16'd30554, 16'd31148, 16'd3415, 16'd47954, 16'd11069, 16'd58467});
	test_expansion(128'h974fbd04c5de4135e10e9fe568e39d84, {16'd62890, 16'd3732, 16'd25449, 16'd316, 16'd19708, 16'd32724, 16'd7078, 16'd56335, 16'd27698, 16'd28479, 16'd9679, 16'd25060, 16'd6923, 16'd10446, 16'd8344, 16'd21472, 16'd55782, 16'd2865, 16'd1450, 16'd64193, 16'd57866, 16'd44512, 16'd28783, 16'd57045, 16'd3803, 16'd13942});
	test_expansion(128'h4bd7349b6b8e89e87237fc7ed12cbb0f, {16'd46990, 16'd27625, 16'd25495, 16'd11370, 16'd34122, 16'd18215, 16'd59730, 16'd65336, 16'd61815, 16'd35647, 16'd18220, 16'd55993, 16'd54186, 16'd61300, 16'd7316, 16'd10854, 16'd1183, 16'd51139, 16'd4156, 16'd29240, 16'd35748, 16'd52215, 16'd22764, 16'd22981, 16'd16366, 16'd55595});
	test_expansion(128'h0d3326d7203e3d563191c67a11af74ca, {16'd57873, 16'd22001, 16'd56694, 16'd57318, 16'd26597, 16'd44689, 16'd41455, 16'd48556, 16'd44488, 16'd39594, 16'd27078, 16'd31876, 16'd722, 16'd4498, 16'd11650, 16'd15426, 16'd58610, 16'd25259, 16'd2940, 16'd45501, 16'd30547, 16'd4965, 16'd34098, 16'd20111, 16'd2836, 16'd51984});
	test_expansion(128'h3211e0095afbe2667021a3314d6b4382, {16'd9030, 16'd25077, 16'd33629, 16'd57069, 16'd2880, 16'd61585, 16'd30760, 16'd14255, 16'd12428, 16'd13693, 16'd28780, 16'd23283, 16'd59663, 16'd17870, 16'd63794, 16'd60136, 16'd59702, 16'd47664, 16'd62142, 16'd24752, 16'd59322, 16'd57855, 16'd62253, 16'd27611, 16'd54444, 16'd53720});
	test_expansion(128'h79f676800ba193ae2df6388043730aec, {16'd44385, 16'd62849, 16'd16002, 16'd23156, 16'd49722, 16'd49120, 16'd5009, 16'd7206, 16'd30383, 16'd51181, 16'd40632, 16'd23256, 16'd24126, 16'd31062, 16'd29090, 16'd21770, 16'd23048, 16'd5771, 16'd35408, 16'd28782, 16'd46077, 16'd13671, 16'd44648, 16'd61746, 16'd46495, 16'd53283});
	test_expansion(128'h39826fe48a42d086fa45d0fabc849e6b, {16'd40560, 16'd48817, 16'd43671, 16'd64967, 16'd41575, 16'd17577, 16'd49975, 16'd17179, 16'd57724, 16'd42968, 16'd64962, 16'd37823, 16'd42562, 16'd61214, 16'd61512, 16'd2838, 16'd15058, 16'd64207, 16'd11659, 16'd6718, 16'd35254, 16'd3742, 16'd14739, 16'd53966, 16'd276, 16'd8906});
	test_expansion(128'h3a13715e076742a479a33229950d9275, {16'd41249, 16'd15722, 16'd12313, 16'd531, 16'd25787, 16'd25038, 16'd63533, 16'd48518, 16'd52212, 16'd49698, 16'd4676, 16'd32553, 16'd26795, 16'd63541, 16'd43549, 16'd31780, 16'd56080, 16'd44312, 16'd471, 16'd41738, 16'd25341, 16'd24261, 16'd44595, 16'd35666, 16'd42030, 16'd52766});
	test_expansion(128'h18dbe9c46c592b608c0b6973905937b6, {16'd8422, 16'd51314, 16'd19708, 16'd61496, 16'd1647, 16'd4582, 16'd63389, 16'd42843, 16'd30320, 16'd50174, 16'd43523, 16'd23517, 16'd49525, 16'd23021, 16'd50160, 16'd38554, 16'd62459, 16'd9383, 16'd62808, 16'd605, 16'd36125, 16'd44802, 16'd9474, 16'd11400, 16'd43333, 16'd49020});
	test_expansion(128'h97c2ec277bb82023eb6b0a52cd1df93e, {16'd7505, 16'd47895, 16'd36844, 16'd11836, 16'd42242, 16'd40342, 16'd54787, 16'd59458, 16'd52570, 16'd27133, 16'd11445, 16'd55818, 16'd62990, 16'd56740, 16'd35796, 16'd29907, 16'd25427, 16'd62479, 16'd39051, 16'd55838, 16'd24315, 16'd58704, 16'd32767, 16'd40662, 16'd9517, 16'd42953});
	test_expansion(128'hd900adfe02d03f7e2ce4bf3ebcfde0fa, {16'd5977, 16'd3954, 16'd5808, 16'd25958, 16'd33039, 16'd53531, 16'd57064, 16'd36184, 16'd56989, 16'd54648, 16'd50239, 16'd25457, 16'd41925, 16'd61071, 16'd34248, 16'd32383, 16'd9461, 16'd28313, 16'd3986, 16'd7823, 16'd30113, 16'd64615, 16'd26299, 16'd27528, 16'd12730, 16'd3501});
	test_expansion(128'h99880850826b37ac9c232a45cde6c59e, {16'd25114, 16'd65472, 16'd5495, 16'd36620, 16'd37764, 16'd32894, 16'd990, 16'd28950, 16'd16163, 16'd57635, 16'd33044, 16'd46909, 16'd8269, 16'd23807, 16'd15104, 16'd7839, 16'd55161, 16'd5982, 16'd35971, 16'd51395, 16'd9579, 16'd49507, 16'd47351, 16'd11475, 16'd34090, 16'd58800});
	test_expansion(128'h51bc6610cea9d20db15cea841fbe6d61, {16'd3276, 16'd35570, 16'd54483, 16'd54548, 16'd30071, 16'd21812, 16'd53236, 16'd32992, 16'd63364, 16'd16244, 16'd53031, 16'd48393, 16'd33537, 16'd62674, 16'd23083, 16'd30533, 16'd57696, 16'd58054, 16'd30197, 16'd51193, 16'd27962, 16'd42514, 16'd37837, 16'd53971, 16'd5825, 16'd52031});
	test_expansion(128'h8b84850899f3cd4b7c89a71292170c65, {16'd15971, 16'd65179, 16'd6426, 16'd31887, 16'd23830, 16'd6073, 16'd22116, 16'd34480, 16'd45752, 16'd20993, 16'd19938, 16'd6540, 16'd57261, 16'd18979, 16'd23270, 16'd36105, 16'd16284, 16'd61591, 16'd33815, 16'd2283, 16'd6880, 16'd13212, 16'd57894, 16'd19333, 16'd42711, 16'd56439});
	test_expansion(128'hd9eadb642b3d748fbc76a69a6c3e5a17, {16'd53294, 16'd22908, 16'd26811, 16'd6270, 16'd64611, 16'd20103, 16'd12390, 16'd31159, 16'd19264, 16'd33483, 16'd32906, 16'd9792, 16'd14219, 16'd44256, 16'd53657, 16'd305, 16'd15665, 16'd47109, 16'd24038, 16'd8901, 16'd44450, 16'd52253, 16'd9048, 16'd3815, 16'd21460, 16'd37341});
	test_expansion(128'he735eb23fa9cb28144a8b9518d9306a1, {16'd17909, 16'd39910, 16'd58780, 16'd29445, 16'd252, 16'd48729, 16'd38280, 16'd25477, 16'd62024, 16'd30415, 16'd51959, 16'd17241, 16'd52997, 16'd50075, 16'd55142, 16'd35129, 16'd56171, 16'd2314, 16'd63953, 16'd43461, 16'd24671, 16'd49578, 16'd59967, 16'd11524, 16'd60186, 16'd1577});
	test_expansion(128'h632ffeaaa8cc35c900409af981655934, {16'd11098, 16'd18448, 16'd39711, 16'd27280, 16'd46130, 16'd2195, 16'd8148, 16'd57834, 16'd6283, 16'd62677, 16'd42998, 16'd36521, 16'd8171, 16'd37654, 16'd54336, 16'd41263, 16'd45230, 16'd9653, 16'd2219, 16'd49145, 16'd29647, 16'd13633, 16'd53751, 16'd62807, 16'd27365, 16'd64450});
	test_expansion(128'hacd4d8521a85a458e02bbd034612db19, {16'd59175, 16'd42046, 16'd24774, 16'd43221, 16'd64967, 16'd6388, 16'd33879, 16'd29219, 16'd19473, 16'd2773, 16'd19325, 16'd57072, 16'd10172, 16'd7275, 16'd40722, 16'd24586, 16'd44067, 16'd14255, 16'd11345, 16'd57885, 16'd25673, 16'd49223, 16'd12502, 16'd47961, 16'd36975, 16'd30242});
	test_expansion(128'h6f229c98b64866e2bda794f92f8e035b, {16'd30426, 16'd16225, 16'd38105, 16'd57461, 16'd56680, 16'd19449, 16'd8382, 16'd50522, 16'd33524, 16'd30235, 16'd20460, 16'd57466, 16'd22169, 16'd45000, 16'd27381, 16'd3469, 16'd55794, 16'd23597, 16'd59179, 16'd6863, 16'd43630, 16'd61108, 16'd55084, 16'd50549, 16'd46682, 16'd59214});
	test_expansion(128'h95214f1bcb11cd757dec27f0f075887c, {16'd9165, 16'd26709, 16'd3119, 16'd5309, 16'd13628, 16'd1977, 16'd33696, 16'd27951, 16'd34391, 16'd20445, 16'd53855, 16'd52070, 16'd36184, 16'd752, 16'd26301, 16'd18638, 16'd1383, 16'd22805, 16'd56221, 16'd31008, 16'd44244, 16'd44263, 16'd57341, 16'd13446, 16'd12368, 16'd14356});
	test_expansion(128'h8b770c8afc7fdeef2b1ba05b82f765a3, {16'd37809, 16'd5126, 16'd6091, 16'd50144, 16'd55297, 16'd36207, 16'd40487, 16'd60345, 16'd9234, 16'd46470, 16'd13025, 16'd63742, 16'd22993, 16'd31829, 16'd53384, 16'd4495, 16'd58967, 16'd28897, 16'd30850, 16'd28494, 16'd38297, 16'd30080, 16'd5604, 16'd17497, 16'd3499, 16'd52170});
	test_expansion(128'he3f06eb2f69424a0250050a6d0048034, {16'd22175, 16'd3652, 16'd33463, 16'd31232, 16'd44265, 16'd33647, 16'd45211, 16'd60257, 16'd65049, 16'd4217, 16'd27631, 16'd29944, 16'd53886, 16'd6574, 16'd4067, 16'd22363, 16'd13907, 16'd64765, 16'd22275, 16'd14474, 16'd24803, 16'd43483, 16'd22750, 16'd64257, 16'd64725, 16'd28793});
	test_expansion(128'hd5315cd0bef83fc82402155ffef4a59c, {16'd9949, 16'd23892, 16'd38903, 16'd50807, 16'd40399, 16'd27547, 16'd43544, 16'd44577, 16'd7665, 16'd62418, 16'd24951, 16'd32232, 16'd5567, 16'd23728, 16'd50569, 16'd5696, 16'd49964, 16'd32631, 16'd48649, 16'd10983, 16'd58378, 16'd51811, 16'd41408, 16'd23811, 16'd15055, 16'd17217});
	test_expansion(128'heb97777e18d4ae51025bbdfeedbc6de9, {16'd3901, 16'd38452, 16'd1677, 16'd2353, 16'd61677, 16'd58746, 16'd58552, 16'd7769, 16'd29826, 16'd2781, 16'd25899, 16'd24780, 16'd10433, 16'd20304, 16'd11040, 16'd39036, 16'd50849, 16'd10293, 16'd19893, 16'd31968, 16'd39943, 16'd54530, 16'd40801, 16'd38926, 16'd33939, 16'd20895});
	test_expansion(128'h6c53313af46c7b6ef765a356f6e35028, {16'd58517, 16'd33208, 16'd39457, 16'd54974, 16'd8612, 16'd10334, 16'd14450, 16'd28222, 16'd46388, 16'd15338, 16'd6089, 16'd6408, 16'd30124, 16'd33482, 16'd16316, 16'd44473, 16'd56076, 16'd42760, 16'd36454, 16'd41723, 16'd59171, 16'd19490, 16'd46873, 16'd45650, 16'd58193, 16'd35193});
	test_expansion(128'h50fa2f355a561650d48fef90ad9959f6, {16'd9230, 16'd41672, 16'd26251, 16'd22519, 16'd50431, 16'd27312, 16'd38675, 16'd9166, 16'd44373, 16'd4899, 16'd41318, 16'd37335, 16'd16862, 16'd7163, 16'd41878, 16'd29088, 16'd22494, 16'd26562, 16'd54493, 16'd5170, 16'd12460, 16'd32926, 16'd10296, 16'd5617, 16'd21955, 16'd16762});
	test_expansion(128'he61fcab130b8ab979501fea966e17600, {16'd52692, 16'd27468, 16'd38612, 16'd6494, 16'd19410, 16'd63234, 16'd61791, 16'd58363, 16'd15942, 16'd38279, 16'd57939, 16'd5402, 16'd63584, 16'd59399, 16'd46861, 16'd46424, 16'd10252, 16'd45024, 16'd23132, 16'd3861, 16'd52390, 16'd46161, 16'd60182, 16'd28174, 16'd44219, 16'd17606});
	test_expansion(128'h77c6e0208ac670b4b5e074613506a76f, {16'd14426, 16'd15058, 16'd51130, 16'd11349, 16'd11196, 16'd24830, 16'd37373, 16'd24216, 16'd61024, 16'd38457, 16'd42214, 16'd44803, 16'd8745, 16'd27144, 16'd29471, 16'd6708, 16'd45612, 16'd11142, 16'd43411, 16'd59157, 16'd62724, 16'd8, 16'd15702, 16'd16157, 16'd22525, 16'd21979});
	test_expansion(128'hcf40a88b9d95218ad1d617dc426ef9bc, {16'd7148, 16'd21436, 16'd6826, 16'd25875, 16'd56152, 16'd42825, 16'd7176, 16'd43926, 16'd56097, 16'd6155, 16'd55339, 16'd58434, 16'd54961, 16'd23169, 16'd19832, 16'd4952, 16'd7465, 16'd49206, 16'd47800, 16'd40232, 16'd23193, 16'd53373, 16'd60596, 16'd40318, 16'd25482, 16'd39128});
	test_expansion(128'hac9108452e61ebf740988047354b79f3, {16'd15171, 16'd11883, 16'd21148, 16'd58794, 16'd9267, 16'd7508, 16'd54763, 16'd36917, 16'd58226, 16'd55903, 16'd58863, 16'd8376, 16'd62463, 16'd61831, 16'd51002, 16'd16203, 16'd37181, 16'd33654, 16'd58485, 16'd49485, 16'd41755, 16'd7461, 16'd7985, 16'd52901, 16'd40972, 16'd52106});
	test_expansion(128'hf3896832d219d45b8fd9623212dce472, {16'd29376, 16'd58398, 16'd38045, 16'd6957, 16'd58181, 16'd27160, 16'd49233, 16'd5157, 16'd20854, 16'd32453, 16'd17798, 16'd24206, 16'd26503, 16'd53706, 16'd8274, 16'd5910, 16'd31271, 16'd25326, 16'd47625, 16'd56536, 16'd11657, 16'd22221, 16'd56820, 16'd39597, 16'd63047, 16'd25930});
	test_expansion(128'h4d7a355e61d4f1b907acbd9e0af5e0c4, {16'd3239, 16'd47558, 16'd59167, 16'd61939, 16'd31622, 16'd6204, 16'd39895, 16'd18643, 16'd43757, 16'd64108, 16'd64576, 16'd40434, 16'd40935, 16'd64019, 16'd65105, 16'd28012, 16'd21340, 16'd44790, 16'd63879, 16'd48794, 16'd25292, 16'd28183, 16'd17277, 16'd30946, 16'd22801, 16'd51363});
	test_expansion(128'h00df544afb30c3b79ae5906e361dc672, {16'd5970, 16'd58187, 16'd16394, 16'd8019, 16'd7053, 16'd52490, 16'd20021, 16'd47461, 16'd48314, 16'd34989, 16'd21387, 16'd15934, 16'd14155, 16'd63978, 16'd4394, 16'd30345, 16'd2717, 16'd20543, 16'd60495, 16'd51008, 16'd15562, 16'd39759, 16'd45357, 16'd42384, 16'd36920, 16'd38584});
	test_expansion(128'h934e67528382d79f0a96b5c82ed4afed, {16'd8024, 16'd17200, 16'd61927, 16'd64294, 16'd31082, 16'd62038, 16'd43293, 16'd59331, 16'd46087, 16'd32168, 16'd18038, 16'd45149, 16'd5789, 16'd18910, 16'd54230, 16'd40563, 16'd32516, 16'd12221, 16'd61355, 16'd20220, 16'd17272, 16'd10485, 16'd60670, 16'd17983, 16'd59811, 16'd56015});
	test_expansion(128'h872771e97de587929c23c663ba774c59, {16'd22463, 16'd59129, 16'd65398, 16'd15854, 16'd44358, 16'd48769, 16'd26689, 16'd10966, 16'd54924, 16'd18753, 16'd5471, 16'd30801, 16'd33258, 16'd57322, 16'd18214, 16'd60530, 16'd2522, 16'd50656, 16'd13603, 16'd460, 16'd30789, 16'd47820, 16'd17119, 16'd6418, 16'd22201, 16'd5437});
	test_expansion(128'h407b0dd690af3c06de6048374f22e045, {16'd64075, 16'd26272, 16'd32112, 16'd10838, 16'd50248, 16'd58073, 16'd60570, 16'd25399, 16'd21198, 16'd26881, 16'd18445, 16'd63141, 16'd61618, 16'd15931, 16'd51945, 16'd3025, 16'd14979, 16'd44134, 16'd42762, 16'd38345, 16'd45343, 16'd46733, 16'd19458, 16'd28744, 16'd19138, 16'd31104});
	test_expansion(128'h84b320db4237876aaf0df26ce4eab3c3, {16'd46937, 16'd8184, 16'd35825, 16'd43772, 16'd39274, 16'd17476, 16'd17271, 16'd53827, 16'd32127, 16'd27899, 16'd47710, 16'd4137, 16'd29227, 16'd36019, 16'd44563, 16'd11390, 16'd50674, 16'd56308, 16'd47334, 16'd28436, 16'd41515, 16'd35660, 16'd22288, 16'd14410, 16'd21416, 16'd38583});
	test_expansion(128'ha49ad7c0d83c1087ce838516efadf1ac, {16'd21728, 16'd58236, 16'd3340, 16'd11441, 16'd13355, 16'd48866, 16'd52998, 16'd35633, 16'd29544, 16'd62691, 16'd48701, 16'd38609, 16'd40280, 16'd27262, 16'd39887, 16'd1841, 16'd59563, 16'd22909, 16'd30917, 16'd58181, 16'd29417, 16'd31003, 16'd35295, 16'd12324, 16'd27672, 16'd6844});
	test_expansion(128'hd491e9176517d45e451ac84621230f33, {16'd10346, 16'd39624, 16'd40922, 16'd22189, 16'd41776, 16'd1027, 16'd33579, 16'd53423, 16'd13855, 16'd63194, 16'd2664, 16'd19709, 16'd18015, 16'd35057, 16'd55802, 16'd5628, 16'd23730, 16'd3687, 16'd52168, 16'd39368, 16'd54868, 16'd52, 16'd31043, 16'd45840, 16'd4548, 16'd9042});
	test_expansion(128'hacb4e13f55ab5c882128fcc2885b5225, {16'd44589, 16'd32040, 16'd62141, 16'd16273, 16'd13320, 16'd33107, 16'd51475, 16'd41292, 16'd35188, 16'd34726, 16'd60083, 16'd25068, 16'd56366, 16'd23075, 16'd65403, 16'd41600, 16'd1941, 16'd34664, 16'd28491, 16'd25616, 16'd41914, 16'd49951, 16'd36794, 16'd37316, 16'd43588, 16'd8767});
	test_expansion(128'ha90dc0e93cecc6a97563fce703729d0e, {16'd12181, 16'd27548, 16'd16025, 16'd65150, 16'd50460, 16'd47223, 16'd19303, 16'd10878, 16'd61011, 16'd37803, 16'd50736, 16'd33142, 16'd31358, 16'd6922, 16'd2980, 16'd11682, 16'd1678, 16'd50535, 16'd37331, 16'd38357, 16'd42985, 16'd30396, 16'd24857, 16'd45752, 16'd25380, 16'd22329});
	test_expansion(128'h9465a33d6b749fdfb08f16c9d44ec810, {16'd22903, 16'd25103, 16'd56273, 16'd53106, 16'd8090, 16'd2425, 16'd19296, 16'd56664, 16'd56214, 16'd47472, 16'd51543, 16'd65092, 16'd62201, 16'd41345, 16'd56391, 16'd20152, 16'd59129, 16'd55428, 16'd24370, 16'd9293, 16'd28018, 16'd12661, 16'd52718, 16'd52053, 16'd54914, 16'd9169});
	test_expansion(128'he78bb50f6ed4512b230784087774e7b8, {16'd14995, 16'd15425, 16'd40792, 16'd35028, 16'd7788, 16'd18471, 16'd4436, 16'd28453, 16'd48214, 16'd19435, 16'd59169, 16'd38012, 16'd17328, 16'd62881, 16'd20647, 16'd4069, 16'd2289, 16'd21644, 16'd22305, 16'd24742, 16'd13676, 16'd30294, 16'd16865, 16'd10427, 16'd53316, 16'd37436});
	test_expansion(128'h9748021f11a0d4c3c76971298bfba28e, {16'd42715, 16'd10040, 16'd15840, 16'd27558, 16'd60660, 16'd29477, 16'd41981, 16'd38376, 16'd32885, 16'd55169, 16'd56628, 16'd34799, 16'd22548, 16'd15244, 16'd44655, 16'd16265, 16'd55429, 16'd48021, 16'd25655, 16'd34623, 16'd56706, 16'd48175, 16'd50513, 16'd228, 16'd48816, 16'd41013});
	test_expansion(128'h6388157089f3d19bec4ba12ee9136bc4, {16'd9825, 16'd20859, 16'd60740, 16'd11783, 16'd37602, 16'd5165, 16'd1921, 16'd55619, 16'd63142, 16'd29945, 16'd59316, 16'd16651, 16'd16353, 16'd1467, 16'd42559, 16'd13137, 16'd6645, 16'd7274, 16'd54672, 16'd20370, 16'd23471, 16'd26725, 16'd54997, 16'd34434, 16'd26439, 16'd11898});
	test_expansion(128'h4b52f6b87fc4087f8d94112dfb884df4, {16'd54558, 16'd29221, 16'd29931, 16'd50978, 16'd56983, 16'd47474, 16'd63076, 16'd24960, 16'd47066, 16'd36201, 16'd11056, 16'd31606, 16'd51802, 16'd40581, 16'd28246, 16'd19824, 16'd28991, 16'd10298, 16'd2413, 16'd1874, 16'd54981, 16'd42832, 16'd44924, 16'd16271, 16'd47106, 16'd32002});
	test_expansion(128'hdbe06e2880e6bdb5937324ae8adfda96, {16'd24643, 16'd57922, 16'd41592, 16'd58738, 16'd55985, 16'd37795, 16'd12897, 16'd2331, 16'd64511, 16'd5822, 16'd59529, 16'd19211, 16'd62645, 16'd16854, 16'd23757, 16'd40482, 16'd32844, 16'd55316, 16'd59359, 16'd15632, 16'd26505, 16'd17368, 16'd6493, 16'd14588, 16'd31206, 16'd42165});
	test_expansion(128'h936507fc62eb6a11556d59aadbc80622, {16'd46710, 16'd59257, 16'd48023, 16'd58540, 16'd50450, 16'd2167, 16'd8997, 16'd47881, 16'd15350, 16'd24920, 16'd7323, 16'd39289, 16'd4635, 16'd16590, 16'd41032, 16'd44375, 16'd13880, 16'd2710, 16'd54952, 16'd43017, 16'd41262, 16'd59594, 16'd46760, 16'd43230, 16'd62203, 16'd3884});
	test_expansion(128'h5d5d17552f45805721e0050e9822a2f8, {16'd57801, 16'd35139, 16'd44490, 16'd62609, 16'd19641, 16'd61706, 16'd51012, 16'd51215, 16'd47046, 16'd61642, 16'd15177, 16'd30141, 16'd27540, 16'd6637, 16'd18372, 16'd937, 16'd3533, 16'd44393, 16'd23927, 16'd8679, 16'd56512, 16'd39909, 16'd54029, 16'd43906, 16'd41360, 16'd43447});
	test_expansion(128'hc1fa94be1da7630e5ea75b91abb977ea, {16'd48956, 16'd47698, 16'd37391, 16'd7494, 16'd48281, 16'd45289, 16'd55076, 16'd58247, 16'd60142, 16'd27629, 16'd21730, 16'd63763, 16'd13029, 16'd18819, 16'd9401, 16'd52511, 16'd42067, 16'd27643, 16'd37972, 16'd65352, 16'd33427, 16'd50008, 16'd51517, 16'd55836, 16'd59778, 16'd63950});
	test_expansion(128'h813c286a303eb7b9c57d9e1e15b7b830, {16'd20975, 16'd54972, 16'd41865, 16'd7805, 16'd32221, 16'd17938, 16'd48380, 16'd22193, 16'd48024, 16'd14651, 16'd2127, 16'd17906, 16'd641, 16'd45203, 16'd17370, 16'd9711, 16'd45078, 16'd42624, 16'd35457, 16'd53763, 16'd13486, 16'd56064, 16'd20273, 16'd56851, 16'd20522, 16'd21547});
	test_expansion(128'haf39e7829b2daab871bfc2e76671b18c, {16'd37836, 16'd18529, 16'd2718, 16'd4752, 16'd26414, 16'd64659, 16'd30451, 16'd51120, 16'd40830, 16'd48531, 16'd62414, 16'd63529, 16'd44852, 16'd40879, 16'd8737, 16'd32404, 16'd29171, 16'd5481, 16'd9067, 16'd14380, 16'd60592, 16'd48254, 16'd7686, 16'd45012, 16'd16976, 16'd11890});
	test_expansion(128'h60c6a0953a64efc34b12e7926237a682, {16'd58722, 16'd39005, 16'd48518, 16'd39183, 16'd9283, 16'd65186, 16'd23809, 16'd44872, 16'd61283, 16'd53870, 16'd4713, 16'd34949, 16'd5506, 16'd25333, 16'd49812, 16'd48382, 16'd40380, 16'd38683, 16'd3285, 16'd35989, 16'd46259, 16'd23190, 16'd8449, 16'd40123, 16'd16546, 16'd4468});
	test_expansion(128'h7d5f14b12516be82492b55591a2c8546, {16'd41188, 16'd57924, 16'd58208, 16'd64044, 16'd37711, 16'd43793, 16'd42143, 16'd43704, 16'd44013, 16'd15458, 16'd50433, 16'd20415, 16'd5803, 16'd57958, 16'd37830, 16'd57740, 16'd50807, 16'd19195, 16'd40812, 16'd43867, 16'd32535, 16'd49984, 16'd11564, 16'd2749, 16'd19503, 16'd28887});
	test_expansion(128'h25befb06260b5dd1ba68179b26eaf9e1, {16'd49036, 16'd21491, 16'd36480, 16'd14901, 16'd5041, 16'd28256, 16'd39090, 16'd50131, 16'd35475, 16'd5356, 16'd46290, 16'd3234, 16'd14849, 16'd35350, 16'd15983, 16'd31924, 16'd58906, 16'd10719, 16'd3373, 16'd33518, 16'd2875, 16'd35088, 16'd61388, 16'd41100, 16'd32514, 16'd11105});
	test_expansion(128'h934c40bb2ae289f1ee6d366c2fe79caf, {16'd11290, 16'd58683, 16'd48642, 16'd7933, 16'd7078, 16'd37224, 16'd1858, 16'd39473, 16'd13544, 16'd14746, 16'd51937, 16'd32144, 16'd41494, 16'd39885, 16'd40106, 16'd11289, 16'd2992, 16'd14917, 16'd5171, 16'd41610, 16'd64013, 16'd33182, 16'd51503, 16'd49133, 16'd18134, 16'd8095});
	test_expansion(128'hc8688ac51c171239124462fac3abadbb, {16'd24023, 16'd39364, 16'd41414, 16'd59868, 16'd2919, 16'd23215, 16'd57264, 16'd61898, 16'd18784, 16'd12624, 16'd32091, 16'd56916, 16'd33342, 16'd31419, 16'd48638, 16'd45461, 16'd34861, 16'd11611, 16'd15327, 16'd36445, 16'd24687, 16'd18089, 16'd43143, 16'd34827, 16'd62607, 16'd39060});
	test_expansion(128'ha4285d07426aa46702af63acd94d3eba, {16'd4628, 16'd65095, 16'd27492, 16'd20080, 16'd38694, 16'd49766, 16'd15932, 16'd27850, 16'd20573, 16'd7210, 16'd16455, 16'd5297, 16'd28120, 16'd61226, 16'd22522, 16'd15330, 16'd35358, 16'd58711, 16'd6799, 16'd63285, 16'd9265, 16'd16509, 16'd9445, 16'd19973, 16'd32543, 16'd21082});
	test_expansion(128'h0770dc1ce0f7143df1b2053ebb5c565a, {16'd57825, 16'd35427, 16'd29335, 16'd45535, 16'd21691, 16'd53092, 16'd41338, 16'd14545, 16'd59770, 16'd30226, 16'd60645, 16'd64868, 16'd20406, 16'd24893, 16'd29955, 16'd5144, 16'd46083, 16'd4034, 16'd30864, 16'd1394, 16'd44069, 16'd52800, 16'd16563, 16'd2365, 16'd24091, 16'd35842});
	test_expansion(128'hf3cc0d2232f4eb968343ebdee235416d, {16'd24905, 16'd60808, 16'd30717, 16'd58058, 16'd36764, 16'd12799, 16'd15674, 16'd39097, 16'd48502, 16'd49604, 16'd23667, 16'd37378, 16'd33683, 16'd48894, 16'd21726, 16'd28807, 16'd23601, 16'd58802, 16'd45979, 16'd16109, 16'd29057, 16'd15556, 16'd41088, 16'd10131, 16'd40375, 16'd54638});
	test_expansion(128'h068a3eabea6fecf59e85d265e3495cf3, {16'd31210, 16'd9308, 16'd64395, 16'd20922, 16'd45845, 16'd60710, 16'd38659, 16'd57137, 16'd54253, 16'd53262, 16'd20648, 16'd2734, 16'd42226, 16'd41225, 16'd10791, 16'd54317, 16'd10843, 16'd57220, 16'd1655, 16'd39643, 16'd9459, 16'd12433, 16'd1767, 16'd45248, 16'd53417, 16'd4324});
	test_expansion(128'h5a5c8f18ba501643d0d3856b21fdb83f, {16'd49015, 16'd62591, 16'd3685, 16'd15771, 16'd24620, 16'd14751, 16'd28829, 16'd51730, 16'd9196, 16'd22669, 16'd46870, 16'd51420, 16'd37675, 16'd37330, 16'd14131, 16'd26601, 16'd52513, 16'd6594, 16'd38544, 16'd57941, 16'd41240, 16'd42036, 16'd25558, 16'd10252, 16'd41031, 16'd63266});
	test_expansion(128'h32e7ba9903501b4d40023c7b2450ac0f, {16'd62697, 16'd41249, 16'd58702, 16'd24372, 16'd3471, 16'd4019, 16'd4973, 16'd10899, 16'd39434, 16'd17457, 16'd54776, 16'd51384, 16'd4170, 16'd62449, 16'd21032, 16'd57652, 16'd47218, 16'd55213, 16'd24183, 16'd5837, 16'd51007, 16'd11434, 16'd29884, 16'd7295, 16'd39574, 16'd65454});
	test_expansion(128'h3fc51e2e642eb594b4ae2b3e2914ef89, {16'd33897, 16'd19800, 16'd4475, 16'd46868, 16'd28909, 16'd36957, 16'd16566, 16'd50259, 16'd53276, 16'd57290, 16'd10139, 16'd50617, 16'd6288, 16'd7081, 16'd41285, 16'd45421, 16'd20630, 16'd42320, 16'd20764, 16'd56298, 16'd24579, 16'd59038, 16'd5247, 16'd61286, 16'd52801, 16'd26015});
	test_expansion(128'h37801165671c90130de8d4085e1ec020, {16'd37682, 16'd64808, 16'd37465, 16'd9127, 16'd57640, 16'd34516, 16'd39733, 16'd28895, 16'd27216, 16'd41988, 16'd55138, 16'd47940, 16'd47212, 16'd22793, 16'd35158, 16'd39487, 16'd48508, 16'd19210, 16'd45871, 16'd31841, 16'd64573, 16'd24404, 16'd34142, 16'd13234, 16'd55969, 16'd4181});
	test_expansion(128'h1a2958a3a4c24b0af33fee39fdf5c902, {16'd11915, 16'd61013, 16'd65176, 16'd56018, 16'd61213, 16'd389, 16'd58769, 16'd55219, 16'd32174, 16'd53424, 16'd17498, 16'd13141, 16'd29715, 16'd7515, 16'd65367, 16'd41640, 16'd44949, 16'd35091, 16'd50177, 16'd22528, 16'd34812, 16'd2665, 16'd47281, 16'd46803, 16'd51119, 16'd3363});
	test_expansion(128'h4a9510294be76e89353a82f55eb2828d, {16'd9148, 16'd35107, 16'd31663, 16'd51481, 16'd49925, 16'd971, 16'd20968, 16'd51203, 16'd13038, 16'd41169, 16'd51935, 16'd31099, 16'd37383, 16'd40816, 16'd57315, 16'd30956, 16'd13547, 16'd60284, 16'd20398, 16'd62560, 16'd41405, 16'd47047, 16'd20323, 16'd32040, 16'd13107, 16'd29254});
	test_expansion(128'h0c7812345c63a6baeb22b8e5a2dd0b3b, {16'd48009, 16'd53329, 16'd56638, 16'd23532, 16'd50260, 16'd42498, 16'd55469, 16'd3203, 16'd7960, 16'd7954, 16'd46919, 16'd18822, 16'd48640, 16'd10662, 16'd10230, 16'd50248, 16'd30366, 16'd31898, 16'd61428, 16'd1867, 16'd27376, 16'd62458, 16'd62114, 16'd46599, 16'd52693, 16'd11065});
	test_expansion(128'h5f3b7191890dcedd63c29eadbeafce92, {16'd40250, 16'd61010, 16'd21984, 16'd20589, 16'd41389, 16'd53484, 16'd25535, 16'd21131, 16'd19281, 16'd15193, 16'd18032, 16'd7856, 16'd49634, 16'd8545, 16'd56133, 16'd31008, 16'd49036, 16'd40132, 16'd51958, 16'd29822, 16'd63235, 16'd9029, 16'd32189, 16'd54513, 16'd32071, 16'd14278});
	test_expansion(128'hed05fc2de629b5b0536d9460617bd04c, {16'd48202, 16'd47876, 16'd22049, 16'd37283, 16'd36451, 16'd48409, 16'd3199, 16'd44777, 16'd44686, 16'd51604, 16'd56514, 16'd7721, 16'd32854, 16'd10716, 16'd18353, 16'd44652, 16'd24807, 16'd51134, 16'd7778, 16'd14036, 16'd21792, 16'd9917, 16'd41990, 16'd5776, 16'd32619, 16'd46552});
	test_expansion(128'hc73588bc32b9adab3626b958cad92ea8, {16'd21103, 16'd31211, 16'd34805, 16'd17199, 16'd15396, 16'd55597, 16'd35271, 16'd59108, 16'd54797, 16'd39463, 16'd2067, 16'd52761, 16'd63888, 16'd56217, 16'd26573, 16'd40489, 16'd30097, 16'd26835, 16'd6679, 16'd12135, 16'd9729, 16'd46609, 16'd8857, 16'd55523, 16'd44130, 16'd57227});
	test_expansion(128'hb385515b802ddf7765137610db2dd133, {16'd6611, 16'd13541, 16'd24286, 16'd28589, 16'd38007, 16'd4175, 16'd59591, 16'd5820, 16'd27114, 16'd38388, 16'd38841, 16'd5623, 16'd31063, 16'd44129, 16'd9415, 16'd64279, 16'd57552, 16'd947, 16'd3718, 16'd8501, 16'd15038, 16'd50090, 16'd35230, 16'd64086, 16'd598, 16'd49230});
	test_expansion(128'h6f8972722bcf0b081be7db0cc2b3f114, {16'd23580, 16'd42160, 16'd11907, 16'd64010, 16'd48855, 16'd6343, 16'd24436, 16'd24773, 16'd16234, 16'd8011, 16'd15039, 16'd42769, 16'd40949, 16'd40056, 16'd34735, 16'd15515, 16'd21728, 16'd34028, 16'd20140, 16'd35301, 16'd55290, 16'd35813, 16'd7586, 16'd55856, 16'd65105, 16'd38411});
	test_expansion(128'hf467ef50c374c984e0399b8f13a6f91b, {16'd11412, 16'd12812, 16'd36683, 16'd26728, 16'd7416, 16'd1076, 16'd15932, 16'd13300, 16'd22857, 16'd2089, 16'd58870, 16'd30374, 16'd34104, 16'd60726, 16'd46071, 16'd46751, 16'd21405, 16'd62193, 16'd32609, 16'd2389, 16'd26578, 16'd3190, 16'd49909, 16'd9284, 16'd65532, 16'd28049});
	test_expansion(128'hec414ff1fd3b58301e88ba4331bb462e, {16'd48527, 16'd28187, 16'd65077, 16'd11792, 16'd50458, 16'd60827, 16'd5279, 16'd4839, 16'd15160, 16'd61439, 16'd64036, 16'd55382, 16'd46739, 16'd22061, 16'd39942, 16'd62591, 16'd28800, 16'd33204, 16'd26854, 16'd10802, 16'd35657, 16'd35436, 16'd20346, 16'd43319, 16'd61859, 16'd48558});
	test_expansion(128'h0420cbbe53bd9e9a73b5f1640729e8a0, {16'd5717, 16'd44595, 16'd12128, 16'd65006, 16'd37908, 16'd40291, 16'd14910, 16'd40734, 16'd44269, 16'd47400, 16'd46717, 16'd52467, 16'd12397, 16'd22372, 16'd64488, 16'd63713, 16'd44551, 16'd33977, 16'd44034, 16'd61165, 16'd11880, 16'd1437, 16'd64067, 16'd57065, 16'd2538, 16'd27567});
	test_expansion(128'hd18f828491181f32e097264b7d508eb4, {16'd16629, 16'd4747, 16'd28436, 16'd45119, 16'd47816, 16'd57437, 16'd29215, 16'd37210, 16'd59251, 16'd52577, 16'd42526, 16'd54006, 16'd57427, 16'd53249, 16'd42664, 16'd58810, 16'd18674, 16'd18847, 16'd65049, 16'd15822, 16'd633, 16'd41784, 16'd852, 16'd19498, 16'd30342, 16'd15641});
	test_expansion(128'hee40cb70547d9d03cd201e1df5efa3e0, {16'd36557, 16'd613, 16'd20479, 16'd50055, 16'd21992, 16'd42414, 16'd32002, 16'd56865, 16'd12700, 16'd38891, 16'd56963, 16'd51076, 16'd14091, 16'd43650, 16'd28327, 16'd25881, 16'd32955, 16'd61323, 16'd47813, 16'd51995, 16'd35071, 16'd40386, 16'd4078, 16'd27572, 16'd60218, 16'd4128});
	test_expansion(128'he0b2c163d806a8cda75743c74a0ffbf4, {16'd54869, 16'd39648, 16'd45992, 16'd62714, 16'd9704, 16'd45645, 16'd43616, 16'd10921, 16'd51143, 16'd56759, 16'd40184, 16'd60276, 16'd33834, 16'd45218, 16'd25285, 16'd14167, 16'd58126, 16'd44618, 16'd46224, 16'd28449, 16'd19311, 16'd31487, 16'd53013, 16'd21685, 16'd23799, 16'd39252});
	test_expansion(128'h3fa45edc59dcfe5187e5da315d5c211f, {16'd49960, 16'd8032, 16'd55166, 16'd52878, 16'd4805, 16'd29197, 16'd25793, 16'd46522, 16'd38375, 16'd13054, 16'd57639, 16'd26325, 16'd15018, 16'd11638, 16'd30128, 16'd35183, 16'd33540, 16'd48547, 16'd32012, 16'd8815, 16'd38236, 16'd20634, 16'd25746, 16'd63973, 16'd65085, 16'd30171});
	test_expansion(128'h96f1bcd5799abb70d49078be1974d3fa, {16'd61730, 16'd7314, 16'd25637, 16'd52840, 16'd52173, 16'd27354, 16'd24576, 16'd36176, 16'd25116, 16'd44462, 16'd13505, 16'd27487, 16'd10496, 16'd37392, 16'd26842, 16'd49064, 16'd56817, 16'd44294, 16'd40803, 16'd4929, 16'd56276, 16'd27118, 16'd61290, 16'd26374, 16'd20876, 16'd63298});
	test_expansion(128'h1aa8ff099c6441de3f297348cfc38757, {16'd7833, 16'd41533, 16'd62503, 16'd548, 16'd33076, 16'd35469, 16'd54612, 16'd326, 16'd22368, 16'd27259, 16'd11537, 16'd2553, 16'd15003, 16'd5308, 16'd34094, 16'd12645, 16'd16167, 16'd59842, 16'd38839, 16'd5959, 16'd11789, 16'd27909, 16'd12260, 16'd11591, 16'd61829, 16'd5700});
	test_expansion(128'h8a62ffbfacab368a3e5e9d1136cb86f5, {16'd14411, 16'd58808, 16'd61497, 16'd29959, 16'd19170, 16'd7697, 16'd53195, 16'd4204, 16'd60916, 16'd33433, 16'd33762, 16'd34104, 16'd8393, 16'd23862, 16'd2030, 16'd767, 16'd55926, 16'd35853, 16'd49833, 16'd29511, 16'd38470, 16'd26793, 16'd63409, 16'd5952, 16'd5953, 16'd28067});
	test_expansion(128'h10214f9a1e8b7931805769e98e53f31a, {16'd6543, 16'd1629, 16'd44236, 16'd28717, 16'd7508, 16'd53936, 16'd59635, 16'd855, 16'd10927, 16'd19639, 16'd20984, 16'd11738, 16'd11001, 16'd41781, 16'd43741, 16'd48003, 16'd3016, 16'd47579, 16'd2204, 16'd64347, 16'd38231, 16'd13413, 16'd15272, 16'd42920, 16'd32850, 16'd42679});
	test_expansion(128'h7b09f30257d10feb44099fabcc97b4a3, {16'd6420, 16'd13994, 16'd31006, 16'd16856, 16'd17508, 16'd61334, 16'd2042, 16'd7321, 16'd22691, 16'd54735, 16'd13515, 16'd10707, 16'd54794, 16'd19762, 16'd21099, 16'd17058, 16'd11815, 16'd6015, 16'd49209, 16'd31909, 16'd61073, 16'd1068, 16'd22112, 16'd4595, 16'd38660, 16'd43373});
	test_expansion(128'ha7c681dceda800b5d4ad0ba431575183, {16'd37314, 16'd5594, 16'd13980, 16'd48703, 16'd66, 16'd12614, 16'd61084, 16'd23075, 16'd49525, 16'd65526, 16'd18999, 16'd64255, 16'd56536, 16'd27244, 16'd499, 16'd3028, 16'd49680, 16'd35617, 16'd14031, 16'd50664, 16'd58795, 16'd41949, 16'd30283, 16'd61522, 16'd59330, 16'd58605});
	test_expansion(128'h35cbce3cd8b7afc05fc00aa84c5176d7, {16'd54153, 16'd12876, 16'd39132, 16'd37557, 16'd44915, 16'd64912, 16'd60972, 16'd7542, 16'd27691, 16'd2259, 16'd50325, 16'd62602, 16'd25493, 16'd9162, 16'd52116, 16'd30537, 16'd26706, 16'd59706, 16'd49550, 16'd56158, 16'd15689, 16'd19035, 16'd54736, 16'd62664, 16'd20204, 16'd9261});
	test_expansion(128'hbf6435b55e4e3cd0cade8aca35004996, {16'd63089, 16'd14250, 16'd52454, 16'd8426, 16'd2699, 16'd32183, 16'd24422, 16'd1442, 16'd7852, 16'd30168, 16'd5285, 16'd23840, 16'd44385, 16'd36752, 16'd53636, 16'd45217, 16'd21347, 16'd19427, 16'd41978, 16'd2648, 16'd2024, 16'd13533, 16'd40974, 16'd9544, 16'd40528, 16'd40212});
	test_expansion(128'h00224f19000f602407680c38b840e7dd, {16'd1663, 16'd55344, 16'd45601, 16'd47280, 16'd22697, 16'd48543, 16'd56025, 16'd36079, 16'd8294, 16'd11315, 16'd49688, 16'd33818, 16'd38699, 16'd6028, 16'd7434, 16'd4010, 16'd3375, 16'd53896, 16'd9811, 16'd19058, 16'd1921, 16'd50293, 16'd37607, 16'd18200, 16'd28781, 16'd8978});
	test_expansion(128'h22509d3f6a61ce57b4ff7973f567a260, {16'd5064, 16'd5096, 16'd50787, 16'd44865, 16'd16542, 16'd29950, 16'd39593, 16'd60353, 16'd59138, 16'd6862, 16'd35411, 16'd43398, 16'd6698, 16'd36102, 16'd14711, 16'd20968, 16'd20557, 16'd64309, 16'd21594, 16'd65215, 16'd22273, 16'd23848, 16'd19559, 16'd35023, 16'd43357, 16'd6014});
	test_expansion(128'h311c5ab04de2270bc184782d6238b60f, {16'd46023, 16'd38096, 16'd26636, 16'd7078, 16'd44170, 16'd55852, 16'd7578, 16'd9337, 16'd21133, 16'd44429, 16'd1132, 16'd8679, 16'd48292, 16'd14381, 16'd42750, 16'd65216, 16'd23264, 16'd38876, 16'd31192, 16'd8303, 16'd13015, 16'd13886, 16'd854, 16'd18899, 16'd61669, 16'd46929});
	test_expansion(128'hadd5735831b7566c5d1c90829ad88fed, {16'd948, 16'd65427, 16'd58045, 16'd61169, 16'd19888, 16'd11263, 16'd30202, 16'd16994, 16'd44236, 16'd62851, 16'd30896, 16'd36479, 16'd26555, 16'd13054, 16'd47794, 16'd48720, 16'd35293, 16'd11501, 16'd32885, 16'd2118, 16'd44750, 16'd2531, 16'd49111, 16'd10629, 16'd36086, 16'd32694});
	test_expansion(128'h10ff9c40ce076b2713c3e8e6ef88d1fc, {16'd23198, 16'd5646, 16'd54338, 16'd41973, 16'd37076, 16'd31164, 16'd14844, 16'd33369, 16'd44576, 16'd29239, 16'd30470, 16'd29817, 16'd44559, 16'd51592, 16'd12446, 16'd26034, 16'd8289, 16'd27580, 16'd25138, 16'd25969, 16'd60801, 16'd56560, 16'd38561, 16'd2146, 16'd29060, 16'd49567});
	test_expansion(128'h1b4aa67acf893d3722e34e997431739f, {16'd23654, 16'd5770, 16'd18921, 16'd31367, 16'd46129, 16'd705, 16'd56541, 16'd28914, 16'd1501, 16'd39815, 16'd34775, 16'd31429, 16'd2983, 16'd24419, 16'd27654, 16'd3279, 16'd46369, 16'd8224, 16'd46008, 16'd55209, 16'd56068, 16'd14931, 16'd45398, 16'd12078, 16'd31556, 16'd51738});
	test_expansion(128'h828552deb872ef07541a7858023d4357, {16'd21102, 16'd24223, 16'd24807, 16'd26664, 16'd13462, 16'd52434, 16'd39394, 16'd61378, 16'd52730, 16'd45311, 16'd33921, 16'd24689, 16'd24808, 16'd62202, 16'd39700, 16'd57116, 16'd29601, 16'd25114, 16'd44351, 16'd2710, 16'd62086, 16'd47852, 16'd54310, 16'd43748, 16'd21889, 16'd51344});
	test_expansion(128'h0e86ab577c99b31caffe68059ac11ad7, {16'd64243, 16'd14485, 16'd58455, 16'd22612, 16'd47782, 16'd1249, 16'd53437, 16'd5962, 16'd49519, 16'd61506, 16'd9326, 16'd8609, 16'd18150, 16'd61163, 16'd30539, 16'd19253, 16'd60162, 16'd3979, 16'd18432, 16'd5089, 16'd61072, 16'd8527, 16'd38877, 16'd29848, 16'd3084, 16'd39169});
	test_expansion(128'hf671a4fec1a38191e421c2cbab2f84e6, {16'd4354, 16'd64465, 16'd44369, 16'd28879, 16'd4570, 16'd60882, 16'd45552, 16'd27357, 16'd38050, 16'd36572, 16'd1834, 16'd47962, 16'd34352, 16'd59856, 16'd63532, 16'd49372, 16'd6634, 16'd39131, 16'd52028, 16'd5105, 16'd28403, 16'd63973, 16'd24172, 16'd37553, 16'd56659, 16'd43177});
	test_expansion(128'hf169c1e74a10c9501b89e3bb6edfef3c, {16'd41723, 16'd20518, 16'd52155, 16'd59710, 16'd20719, 16'd34207, 16'd52013, 16'd34941, 16'd2037, 16'd49899, 16'd46972, 16'd24774, 16'd29568, 16'd24662, 16'd39498, 16'd42759, 16'd46786, 16'd11131, 16'd35974, 16'd58674, 16'd35096, 16'd4777, 16'd34853, 16'd46671, 16'd55836, 16'd65394});
	test_expansion(128'hbc14d0ff3d113e6df99aa16f70b758f5, {16'd46669, 16'd60688, 16'd58188, 16'd63750, 16'd29780, 16'd55744, 16'd19231, 16'd64721, 16'd59425, 16'd43018, 16'd61575, 16'd37438, 16'd574, 16'd63097, 16'd62078, 16'd2249, 16'd9473, 16'd42138, 16'd6750, 16'd57401, 16'd42061, 16'd62424, 16'd63629, 16'd1572, 16'd48424, 16'd49284});
	test_expansion(128'h590796331b60a8d0b665be610c283811, {16'd37778, 16'd63314, 16'd12841, 16'd15414, 16'd51793, 16'd44222, 16'd51987, 16'd2620, 16'd4697, 16'd27015, 16'd49901, 16'd3285, 16'd49472, 16'd32987, 16'd44828, 16'd16252, 16'd57706, 16'd15405, 16'd11688, 16'd31860, 16'd8178, 16'd13901, 16'd42439, 16'd7390, 16'd64309, 16'd20802});
	test_expansion(128'h1a1084810cd3519234343be31b9ec9f8, {16'd64267, 16'd27629, 16'd34724, 16'd7299, 16'd28980, 16'd7498, 16'd24117, 16'd41588, 16'd32465, 16'd32795, 16'd44620, 16'd28827, 16'd56841, 16'd4583, 16'd29698, 16'd59006, 16'd485, 16'd16994, 16'd52533, 16'd26013, 16'd39528, 16'd52979, 16'd20845, 16'd2371, 16'd58128, 16'd19980});
	test_expansion(128'h414510137fb723a51e3184455e49bcb2, {16'd31444, 16'd40657, 16'd39881, 16'd63355, 16'd27313, 16'd22377, 16'd60926, 16'd64006, 16'd4740, 16'd37893, 16'd37205, 16'd58814, 16'd32340, 16'd56242, 16'd16063, 16'd54698, 16'd17530, 16'd2706, 16'd58842, 16'd21085, 16'd42318, 16'd25514, 16'd25159, 16'd11163, 16'd59615, 16'd6796});
	test_expansion(128'hffd67945b84acdc09bc1ad03a7102c6f, {16'd17893, 16'd9631, 16'd60188, 16'd36601, 16'd2370, 16'd54824, 16'd55514, 16'd11085, 16'd4083, 16'd15309, 16'd21389, 16'd56926, 16'd647, 16'd51051, 16'd23156, 16'd61901, 16'd32387, 16'd43792, 16'd35131, 16'd39497, 16'd65003, 16'd50247, 16'd19959, 16'd40207, 16'd14583, 16'd47028});
	test_expansion(128'hc49fe17b391023ba93c2bada1d00379f, {16'd39911, 16'd60143, 16'd64155, 16'd21508, 16'd1586, 16'd25003, 16'd40485, 16'd36390, 16'd27874, 16'd58522, 16'd55222, 16'd54962, 16'd1334, 16'd47259, 16'd17354, 16'd53093, 16'd52717, 16'd46137, 16'd53245, 16'd8700, 16'd1583, 16'd6281, 16'd14222, 16'd15582, 16'd48010, 16'd934});
	test_expansion(128'h1c80d28ec9be964d09893dbada0760dc, {16'd57188, 16'd36604, 16'd33698, 16'd12449, 16'd13748, 16'd22978, 16'd45279, 16'd33170, 16'd46227, 16'd25821, 16'd33026, 16'd51035, 16'd36588, 16'd64109, 16'd21366, 16'd13426, 16'd11873, 16'd20876, 16'd29890, 16'd27924, 16'd5957, 16'd39077, 16'd31995, 16'd34544, 16'd662, 16'd36338});
	test_expansion(128'h06e76a511f9c4844c3d4ff9909002e25, {16'd5837, 16'd28353, 16'd19209, 16'd27675, 16'd35158, 16'd47265, 16'd14446, 16'd11303, 16'd3368, 16'd43646, 16'd17300, 16'd38771, 16'd34658, 16'd53424, 16'd33314, 16'd29702, 16'd31045, 16'd52322, 16'd27569, 16'd5255, 16'd42561, 16'd2099, 16'd17122, 16'd13380, 16'd3774, 16'd32081});
	test_expansion(128'hac4721a3e1aa97841b28210b8efc7edc, {16'd15752, 16'd41672, 16'd60947, 16'd62955, 16'd37388, 16'd36047, 16'd20991, 16'd2077, 16'd53229, 16'd10519, 16'd37728, 16'd13111, 16'd14311, 16'd61258, 16'd41019, 16'd46407, 16'd9167, 16'd63477, 16'd51298, 16'd20582, 16'd35415, 16'd27505, 16'd16956, 16'd27855, 16'd12053, 16'd19689});
	test_expansion(128'h5f516d6527353da9dfb9b03898f940c5, {16'd58977, 16'd56940, 16'd32442, 16'd1167, 16'd9551, 16'd60298, 16'd910, 16'd41225, 16'd36089, 16'd18974, 16'd50114, 16'd29705, 16'd58312, 16'd22354, 16'd556, 16'd54560, 16'd21667, 16'd38688, 16'd976, 16'd15377, 16'd18992, 16'd48568, 16'd32090, 16'd56969, 16'd9778, 16'd61886});
	test_expansion(128'h81a7bbfa6928dbb3e440f40a22f7df03, {16'd19391, 16'd53550, 16'd24008, 16'd63039, 16'd29696, 16'd41052, 16'd47954, 16'd8309, 16'd42415, 16'd16624, 16'd48145, 16'd61859, 16'd39773, 16'd11484, 16'd65290, 16'd26913, 16'd55393, 16'd32124, 16'd16058, 16'd52387, 16'd14368, 16'd49148, 16'd42403, 16'd43969, 16'd16847, 16'd13456});
	test_expansion(128'hbca7b6d15d4c7adb5ce870eaf6dd90c1, {16'd56620, 16'd35480, 16'd16670, 16'd32915, 16'd21976, 16'd11413, 16'd22736, 16'd11347, 16'd39247, 16'd34686, 16'd10647, 16'd34473, 16'd9773, 16'd61556, 16'd37790, 16'd412, 16'd36765, 16'd42221, 16'd18433, 16'd6070, 16'd19163, 16'd23851, 16'd36144, 16'd13733, 16'd19160, 16'd57508});
	test_expansion(128'hdae26a488aa0ad257942204c0b59d1c1, {16'd408, 16'd50870, 16'd22111, 16'd26171, 16'd21143, 16'd14947, 16'd42933, 16'd55240, 16'd16226, 16'd58075, 16'd36075, 16'd13321, 16'd62142, 16'd32283, 16'd58490, 16'd16032, 16'd61097, 16'd50831, 16'd48892, 16'd50450, 16'd63912, 16'd15627, 16'd38165, 16'd52319, 16'd30248, 16'd39051});
	test_expansion(128'h22cc293250156ab7a92ed61275d741e6, {16'd19584, 16'd38971, 16'd7896, 16'd3502, 16'd47209, 16'd1148, 16'd58266, 16'd50484, 16'd41948, 16'd38741, 16'd9209, 16'd62209, 16'd58663, 16'd54165, 16'd6625, 16'd58735, 16'd45905, 16'd25768, 16'd41603, 16'd34532, 16'd54846, 16'd34527, 16'd55877, 16'd50388, 16'd65008, 16'd7771});
	test_expansion(128'h07d13ab4148bec61b97da41ab18bfcfc, {16'd55533, 16'd18204, 16'd26544, 16'd29146, 16'd27596, 16'd49452, 16'd64230, 16'd10045, 16'd11861, 16'd7986, 16'd62059, 16'd19983, 16'd35595, 16'd57792, 16'd42829, 16'd26198, 16'd22250, 16'd33437, 16'd13887, 16'd50749, 16'd53579, 16'd41209, 16'd57283, 16'd54825, 16'd63136, 16'd30003});
	test_expansion(128'h070e7080623f98d00acc20f3000f5c49, {16'd26354, 16'd26851, 16'd24278, 16'd54259, 16'd18196, 16'd45022, 16'd2438, 16'd12292, 16'd32787, 16'd24729, 16'd6416, 16'd51794, 16'd3246, 16'd16937, 16'd32864, 16'd55155, 16'd41114, 16'd5689, 16'd7387, 16'd3114, 16'd61378, 16'd15840, 16'd13153, 16'd36624, 16'd15769, 16'd27923});
	test_expansion(128'h69395ccaea1f8cff6f45826ba618b182, {16'd23852, 16'd41974, 16'd53992, 16'd41933, 16'd47224, 16'd44413, 16'd21799, 16'd27012, 16'd32958, 16'd19727, 16'd4234, 16'd2667, 16'd50817, 16'd2159, 16'd22515, 16'd31387, 16'd47571, 16'd63962, 16'd46398, 16'd32073, 16'd6377, 16'd62393, 16'd40421, 16'd47064, 16'd30764, 16'd56948});
	test_expansion(128'h56a564598d2216ccb2e659cab330148f, {16'd17052, 16'd4616, 16'd32250, 16'd14558, 16'd64811, 16'd11721, 16'd30601, 16'd23169, 16'd56502, 16'd49392, 16'd30978, 16'd24406, 16'd33651, 16'd2732, 16'd56328, 16'd45115, 16'd4362, 16'd35911, 16'd45982, 16'd14840, 16'd84, 16'd49761, 16'd2870, 16'd63890, 16'd13540, 16'd12921});
	test_expansion(128'hd92d70b5c40200cb0b650aa079e4d6ae, {16'd12769, 16'd56049, 16'd51990, 16'd44540, 16'd15714, 16'd48118, 16'd9938, 16'd9709, 16'd28581, 16'd52705, 16'd12911, 16'd30598, 16'd21319, 16'd49404, 16'd32016, 16'd18716, 16'd61052, 16'd1180, 16'd48803, 16'd34580, 16'd10843, 16'd57333, 16'd50520, 16'd52524, 16'd11153, 16'd20011});
	test_expansion(128'he8cb6c3670af636c7315db296d097632, {16'd3026, 16'd14513, 16'd29177, 16'd59221, 16'd32436, 16'd3747, 16'd10663, 16'd61994, 16'd38274, 16'd59188, 16'd26625, 16'd37822, 16'd4747, 16'd25519, 16'd21606, 16'd48888, 16'd31227, 16'd62069, 16'd37570, 16'd42639, 16'd49685, 16'd48540, 16'd4624, 16'd35896, 16'd20261, 16'd122});
	test_expansion(128'h756e3ec613999375883a87c2c62e46fc, {16'd18845, 16'd30905, 16'd32511, 16'd44912, 16'd60021, 16'd12674, 16'd29219, 16'd26763, 16'd10179, 16'd25609, 16'd63680, 16'd32658, 16'd22117, 16'd54212, 16'd61993, 16'd43976, 16'd19511, 16'd44088, 16'd16804, 16'd63104, 16'd35682, 16'd36680, 16'd54123, 16'd10233, 16'd31080, 16'd40642});
	test_expansion(128'h9f5208e05a155086a8cfe63f3cb68daf, {16'd12319, 16'd4402, 16'd11383, 16'd29878, 16'd49850, 16'd38583, 16'd22702, 16'd16828, 16'd48279, 16'd53804, 16'd20886, 16'd55516, 16'd1668, 16'd51200, 16'd20752, 16'd45808, 16'd13060, 16'd29083, 16'd10759, 16'd21423, 16'd2690, 16'd22589, 16'd41136, 16'd54136, 16'd52075, 16'd51965});
	test_expansion(128'hb66280e853e06c89d030c2ce013f5a7a, {16'd5801, 16'd34538, 16'd40070, 16'd12434, 16'd6047, 16'd36064, 16'd21682, 16'd8487, 16'd2089, 16'd64702, 16'd18932, 16'd47925, 16'd56521, 16'd10239, 16'd13638, 16'd43474, 16'd6216, 16'd19387, 16'd31692, 16'd17149, 16'd39758, 16'd1155, 16'd30495, 16'd55930, 16'd54988, 16'd33073});
	test_expansion(128'h8b42ecfb4e3c146d521c01631beab3a5, {16'd56926, 16'd24857, 16'd6890, 16'd7253, 16'd27694, 16'd47282, 16'd22656, 16'd57347, 16'd59283, 16'd62751, 16'd32966, 16'd45873, 16'd20586, 16'd8981, 16'd51306, 16'd37603, 16'd4190, 16'd32440, 16'd22859, 16'd57958, 16'd5586, 16'd692, 16'd64815, 16'd23066, 16'd17162, 16'd27344});
	test_expansion(128'h25aac2caa184a73c408efe5759d2b758, {16'd41624, 16'd40641, 16'd47787, 16'd62483, 16'd40546, 16'd56454, 16'd42549, 16'd24912, 16'd65442, 16'd32813, 16'd19608, 16'd34814, 16'd19315, 16'd24877, 16'd56856, 16'd42274, 16'd41176, 16'd43856, 16'd63259, 16'd6714, 16'd24961, 16'd26753, 16'd8156, 16'd21088, 16'd65159, 16'd19358});
	test_expansion(128'hba7fa9ed88fe9f9f1e9ff4c1ed63569d, {16'd4921, 16'd59784, 16'd33645, 16'd47770, 16'd19544, 16'd46293, 16'd40629, 16'd1548, 16'd53917, 16'd61033, 16'd25819, 16'd40038, 16'd39731, 16'd28662, 16'd20932, 16'd33534, 16'd62446, 16'd33780, 16'd44635, 16'd36484, 16'd24907, 16'd34821, 16'd39889, 16'd13629, 16'd23384, 16'd64932});
	test_expansion(128'h42e0290f28caa57cf31b535206867160, {16'd24143, 16'd26209, 16'd12024, 16'd21281, 16'd52196, 16'd46944, 16'd24657, 16'd43703, 16'd29473, 16'd61311, 16'd35964, 16'd31248, 16'd27304, 16'd15434, 16'd61348, 16'd21464, 16'd49955, 16'd8357, 16'd39129, 16'd60255, 16'd13539, 16'd2342, 16'd42529, 16'd29980, 16'd14735, 16'd57750});
	test_expansion(128'h875506cf37bd5602a275e133c64eb7b6, {16'd23860, 16'd341, 16'd29755, 16'd17740, 16'd40704, 16'd23527, 16'd26760, 16'd20889, 16'd57393, 16'd10986, 16'd36810, 16'd9762, 16'd38417, 16'd53531, 16'd14306, 16'd22312, 16'd23808, 16'd36730, 16'd24416, 16'd46524, 16'd37895, 16'd37524, 16'd61868, 16'd4172, 16'd46753, 16'd62272});
	test_expansion(128'h72861c09936ae409e565ecf3286efc42, {16'd19696, 16'd58760, 16'd37750, 16'd63445, 16'd16555, 16'd64824, 16'd21258, 16'd3822, 16'd47935, 16'd54958, 16'd24183, 16'd11438, 16'd42682, 16'd16269, 16'd54446, 16'd16191, 16'd22423, 16'd55916, 16'd57612, 16'd8214, 16'd39242, 16'd53409, 16'd51692, 16'd8462, 16'd29316, 16'd63791});
	test_expansion(128'h670f8c5be6def12e6ae8f2ae81b728ea, {16'd33995, 16'd40132, 16'd60119, 16'd49989, 16'd25143, 16'd22557, 16'd4450, 16'd48078, 16'd63233, 16'd6076, 16'd62147, 16'd35442, 16'd57718, 16'd18517, 16'd36473, 16'd51789, 16'd42190, 16'd5473, 16'd65089, 16'd49315, 16'd65247, 16'd59251, 16'd63524, 16'd5591, 16'd8480, 16'd26473});
	test_expansion(128'h7dd49c389952cc475fac8ecb8232c04b, {16'd51313, 16'd54746, 16'd2146, 16'd27344, 16'd56824, 16'd6298, 16'd65211, 16'd28414, 16'd38373, 16'd34721, 16'd62929, 16'd60889, 16'd41387, 16'd63209, 16'd36135, 16'd36135, 16'd58566, 16'd53655, 16'd27934, 16'd13312, 16'd11969, 16'd7187, 16'd12416, 16'd34853, 16'd1904, 16'd25341});
	test_expansion(128'h9dd8f4c900876ff2ee907d759cfc9f37, {16'd16719, 16'd6094, 16'd35628, 16'd18493, 16'd4242, 16'd1447, 16'd44331, 16'd23650, 16'd47499, 16'd52368, 16'd33449, 16'd60567, 16'd15070, 16'd11650, 16'd10258, 16'd49867, 16'd36517, 16'd9426, 16'd37540, 16'd61331, 16'd14812, 16'd36558, 16'd4414, 16'd51154, 16'd29485, 16'd25928});
	test_expansion(128'h334189542c015cb48131b494845407e2, {16'd57622, 16'd56724, 16'd45118, 16'd6168, 16'd47142, 16'd53450, 16'd23122, 16'd36318, 16'd33426, 16'd42805, 16'd52088, 16'd52486, 16'd32906, 16'd19614, 16'd16527, 16'd58784, 16'd59738, 16'd10239, 16'd56308, 16'd27416, 16'd60638, 16'd27429, 16'd41344, 16'd61537, 16'd5730, 16'd24511});
	test_expansion(128'hea8c2d66371a3fe882e2a04a34a5bd0f, {16'd20380, 16'd39279, 16'd44540, 16'd2807, 16'd18998, 16'd55145, 16'd26274, 16'd42118, 16'd56388, 16'd63533, 16'd30596, 16'd2650, 16'd17347, 16'd65098, 16'd33100, 16'd4924, 16'd43960, 16'd62715, 16'd20775, 16'd36759, 16'd11652, 16'd52322, 16'd64147, 16'd32310, 16'd39889, 16'd65094});
	test_expansion(128'he239b8b42c32886a4f60776f33ee85b8, {16'd60340, 16'd49614, 16'd13669, 16'd23219, 16'd8598, 16'd61579, 16'd41478, 16'd62242, 16'd46075, 16'd1840, 16'd50726, 16'd52937, 16'd13855, 16'd13331, 16'd51642, 16'd37787, 16'd7364, 16'd51276, 16'd54941, 16'd54046, 16'd32682, 16'd60592, 16'd9391, 16'd28523, 16'd9826, 16'd28554});
	test_expansion(128'hfa3698ebcc467c0e92f3bb2d98a1c93d, {16'd45326, 16'd37726, 16'd51061, 16'd29238, 16'd11090, 16'd65163, 16'd46468, 16'd55444, 16'd27923, 16'd1351, 16'd35628, 16'd10582, 16'd64224, 16'd50545, 16'd8217, 16'd33456, 16'd27804, 16'd43828, 16'd1751, 16'd42337, 16'd47271, 16'd51441, 16'd48933, 16'd64, 16'd32419, 16'd62789});
	test_expansion(128'h2a1634b2c396adf956e69fd8292fff93, {16'd15575, 16'd35088, 16'd33159, 16'd12726, 16'd404, 16'd32263, 16'd41098, 16'd13232, 16'd62609, 16'd17280, 16'd61399, 16'd65459, 16'd19467, 16'd35311, 16'd27268, 16'd11311, 16'd34013, 16'd43721, 16'd9842, 16'd3588, 16'd49407, 16'd24170, 16'd9143, 16'd51852, 16'd43139, 16'd33147});
	test_expansion(128'hb583820794e8e8aa3010110537c921a6, {16'd64875, 16'd48506, 16'd54726, 16'd22028, 16'd48057, 16'd46012, 16'd30790, 16'd50433, 16'd8502, 16'd57591, 16'd8941, 16'd54817, 16'd5667, 16'd59222, 16'd36488, 16'd2913, 16'd31809, 16'd45952, 16'd13173, 16'd20448, 16'd28638, 16'd20407, 16'd24761, 16'd54837, 16'd31330, 16'd5227});
	test_expansion(128'hcf64712d449612b2721c8b344633f230, {16'd6507, 16'd30651, 16'd5410, 16'd6818, 16'd64520, 16'd15362, 16'd10817, 16'd42936, 16'd13519, 16'd10530, 16'd32715, 16'd55185, 16'd5156, 16'd8739, 16'd62014, 16'd55796, 16'd14572, 16'd37846, 16'd7856, 16'd40909, 16'd23504, 16'd37377, 16'd12662, 16'd10640, 16'd35486, 16'd4543});
	test_expansion(128'h2face4705ce2b2159948affe12078a7e, {16'd15737, 16'd57828, 16'd20370, 16'd15768, 16'd61285, 16'd45794, 16'd2764, 16'd58937, 16'd8330, 16'd35436, 16'd37431, 16'd20382, 16'd65333, 16'd24528, 16'd13438, 16'd7620, 16'd41970, 16'd64800, 16'd12277, 16'd54450, 16'd28472, 16'd34786, 16'd367, 16'd28691, 16'd58645, 16'd18460});
	test_expansion(128'h6041a1e90efbbff7ce58d7bf69922565, {16'd53639, 16'd61507, 16'd1764, 16'd29376, 16'd46251, 16'd31097, 16'd9206, 16'd42524, 16'd10261, 16'd10377, 16'd13638, 16'd58949, 16'd61552, 16'd20778, 16'd39809, 16'd6393, 16'd56687, 16'd30128, 16'd30824, 16'd40905, 16'd30341, 16'd48411, 16'd39808, 16'd50000, 16'd49633, 16'd9748});
	test_expansion(128'h468d1dce42502254f7abb1096809b8c2, {16'd44673, 16'd4120, 16'd44668, 16'd65225, 16'd40822, 16'd33029, 16'd48041, 16'd5274, 16'd47492, 16'd4570, 16'd49787, 16'd18728, 16'd22865, 16'd50484, 16'd51370, 16'd38476, 16'd47936, 16'd22573, 16'd23637, 16'd44015, 16'd5079, 16'd37021, 16'd37709, 16'd30429, 16'd1147, 16'd56169});
	test_expansion(128'hba723c667c52ba62607a81142d67be11, {16'd16850, 16'd18282, 16'd20881, 16'd38381, 16'd61503, 16'd36950, 16'd45525, 16'd20330, 16'd64340, 16'd38306, 16'd47258, 16'd29131, 16'd39691, 16'd60151, 16'd40720, 16'd13373, 16'd36545, 16'd22926, 16'd24339, 16'd14233, 16'd2477, 16'd6173, 16'd17694, 16'd19806, 16'd10501, 16'd54809});
	test_expansion(128'he6949ffc9a24694e3170fce3de4473fb, {16'd46272, 16'd47447, 16'd5775, 16'd46801, 16'd35534, 16'd48060, 16'd476, 16'd56848, 16'd32851, 16'd65460, 16'd52009, 16'd37925, 16'd17025, 16'd54045, 16'd30190, 16'd30634, 16'd52964, 16'd45879, 16'd32275, 16'd57293, 16'd11438, 16'd27939, 16'd49451, 16'd62359, 16'd37394, 16'd12296});
	test_expansion(128'ha7407a480fa5b774fd4780c6b756fecf, {16'd10632, 16'd33606, 16'd11035, 16'd22774, 16'd33923, 16'd18765, 16'd47973, 16'd24837, 16'd58055, 16'd62422, 16'd24255, 16'd23030, 16'd60619, 16'd34483, 16'd15923, 16'd42333, 16'd8797, 16'd16697, 16'd30961, 16'd37216, 16'd43837, 16'd43780, 16'd49808, 16'd13609, 16'd27770, 16'd32819});
	test_expansion(128'h6669803c7308a461d0f14a772bede6dc, {16'd29915, 16'd18816, 16'd36776, 16'd10501, 16'd35150, 16'd23655, 16'd55181, 16'd26214, 16'd60901, 16'd10180, 16'd53698, 16'd45635, 16'd42263, 16'd216, 16'd25890, 16'd25423, 16'd40411, 16'd5733, 16'd37320, 16'd29196, 16'd21554, 16'd16375, 16'd48744, 16'd19595, 16'd43856, 16'd14976});
	test_expansion(128'hb6184b7ccbe478b8df0641969729a63d, {16'd21041, 16'd17681, 16'd4107, 16'd42560, 16'd37613, 16'd1331, 16'd56541, 16'd60013, 16'd64632, 16'd8443, 16'd23354, 16'd2985, 16'd28239, 16'd31531, 16'd59488, 16'd5808, 16'd42958, 16'd30841, 16'd10993, 16'd44059, 16'd15197, 16'd27489, 16'd17994, 16'd53977, 16'd21011, 16'd8544});
	test_expansion(128'h0caafefe77a9fa98b4bd64ab191634e5, {16'd42808, 16'd51141, 16'd62329, 16'd38559, 16'd62540, 16'd5165, 16'd58501, 16'd9308, 16'd29383, 16'd16162, 16'd26836, 16'd20870, 16'd52811, 16'd41870, 16'd49704, 16'd62573, 16'd58137, 16'd57463, 16'd12584, 16'd21302, 16'd31613, 16'd24934, 16'd62573, 16'd28538, 16'd64831, 16'd23254});
	test_expansion(128'h36c41a96360ccc32ca20729e592f2cf9, {16'd9835, 16'd56227, 16'd53968, 16'd17909, 16'd35705, 16'd6099, 16'd52914, 16'd45054, 16'd28517, 16'd50952, 16'd41541, 16'd1720, 16'd62985, 16'd1780, 16'd16510, 16'd45348, 16'd3963, 16'd28315, 16'd43763, 16'd7941, 16'd3768, 16'd38918, 16'd3545, 16'd20700, 16'd45407, 16'd17093});
	test_expansion(128'hc110c491fda5c2a00c1df98cc269f713, {16'd38558, 16'd48462, 16'd18783, 16'd14989, 16'd17144, 16'd54459, 16'd465, 16'd41563, 16'd10728, 16'd19945, 16'd1575, 16'd37584, 16'd25575, 16'd45207, 16'd60357, 16'd64427, 16'd23161, 16'd101, 16'd64878, 16'd52934, 16'd20710, 16'd51976, 16'd12248, 16'd22297, 16'd25450, 16'd17905});
	test_expansion(128'hf5221e3af7520f5e777172137ae389f8, {16'd41189, 16'd51650, 16'd10916, 16'd20191, 16'd40061, 16'd41044, 16'd27051, 16'd63917, 16'd49939, 16'd7730, 16'd17858, 16'd1423, 16'd43573, 16'd49357, 16'd5078, 16'd60600, 16'd29140, 16'd38609, 16'd29131, 16'd48531, 16'd43135, 16'd8742, 16'd16351, 16'd13839, 16'd48798, 16'd57466});
	test_expansion(128'h72605d63498378d0f400449bc32f320f, {16'd50255, 16'd11221, 16'd31800, 16'd17807, 16'd35963, 16'd20433, 16'd33134, 16'd30666, 16'd61344, 16'd28690, 16'd7899, 16'd31350, 16'd23534, 16'd1928, 16'd23467, 16'd50389, 16'd14455, 16'd18397, 16'd61371, 16'd36873, 16'd11502, 16'd17682, 16'd31716, 16'd57816, 16'd11365, 16'd49682});
	test_expansion(128'hb8279b350ef86a6db67abbb11d4786dd, {16'd32554, 16'd27637, 16'd57931, 16'd51462, 16'd23478, 16'd10585, 16'd56738, 16'd28919, 16'd1237, 16'd4008, 16'd54936, 16'd12780, 16'd6300, 16'd39757, 16'd48036, 16'd57861, 16'd51796, 16'd32067, 16'd43378, 16'd38359, 16'd39534, 16'd36693, 16'd462, 16'd39081, 16'd42991, 16'd21547});
	test_expansion(128'h3ac3bd514292ed18fae21dfb5e48f64b, {16'd38643, 16'd20985, 16'd56431, 16'd24715, 16'd18259, 16'd460, 16'd8162, 16'd39022, 16'd62613, 16'd37136, 16'd46282, 16'd63917, 16'd3537, 16'd6154, 16'd28810, 16'd10515, 16'd33884, 16'd13990, 16'd6491, 16'd16932, 16'd12397, 16'd30329, 16'd40326, 16'd23931, 16'd26600, 16'd5718});
	test_expansion(128'h34d263741632815eaa4c80c3e4d8fa4e, {16'd25481, 16'd14862, 16'd28100, 16'd10750, 16'd26920, 16'd64460, 16'd21267, 16'd11006, 16'd31895, 16'd59415, 16'd55769, 16'd24496, 16'd58251, 16'd37765, 16'd42832, 16'd18473, 16'd48008, 16'd63906, 16'd47955, 16'd54769, 16'd12874, 16'd64721, 16'd7453, 16'd1796, 16'd14684, 16'd31665});
	test_expansion(128'h54d7b8184474ec8d881eb17992787282, {16'd14832, 16'd18176, 16'd58091, 16'd2548, 16'd1887, 16'd29910, 16'd271, 16'd23382, 16'd15550, 16'd33433, 16'd51486, 16'd867, 16'd22277, 16'd12233, 16'd38678, 16'd60089, 16'd26074, 16'd63701, 16'd4495, 16'd41782, 16'd40008, 16'd8631, 16'd19398, 16'd48699, 16'd479, 16'd41015});
	test_expansion(128'h94bd56c83faae559fe70bf46f3fb9b9c, {16'd12297, 16'd19115, 16'd25115, 16'd35699, 16'd8730, 16'd21438, 16'd24119, 16'd25912, 16'd25736, 16'd46129, 16'd14527, 16'd16309, 16'd57513, 16'd46965, 16'd4128, 16'd6552, 16'd2125, 16'd23956, 16'd42583, 16'd24685, 16'd9284, 16'd26709, 16'd63867, 16'd3026, 16'd11796, 16'd29256});
	test_expansion(128'h2c5721abb1f3650dfa3b5c0cb3065e03, {16'd42996, 16'd22884, 16'd8876, 16'd38843, 16'd10656, 16'd5477, 16'd5685, 16'd58952, 16'd842, 16'd31246, 16'd17534, 16'd301, 16'd51034, 16'd10325, 16'd18742, 16'd23402, 16'd11684, 16'd9606, 16'd29919, 16'd60629, 16'd31819, 16'd365, 16'd34505, 16'd26258, 16'd41804, 16'd48085});
	test_expansion(128'h8cfca0f976fbd2fa02d2fedf0585c3c1, {16'd59953, 16'd61134, 16'd50669, 16'd27378, 16'd12176, 16'd40003, 16'd21926, 16'd62292, 16'd32443, 16'd48239, 16'd36656, 16'd39165, 16'd4144, 16'd13496, 16'd45781, 16'd48162, 16'd11209, 16'd52683, 16'd52468, 16'd58795, 16'd48047, 16'd49984, 16'd65006, 16'd23274, 16'd14134, 16'd59601});
	test_expansion(128'h4d3ea92bf2200a19571bcaec65a9836c, {16'd11270, 16'd64495, 16'd55857, 16'd17440, 16'd21631, 16'd46143, 16'd12611, 16'd33411, 16'd7761, 16'd5819, 16'd7292, 16'd62318, 16'd20242, 16'd58069, 16'd64524, 16'd16141, 16'd43526, 16'd34110, 16'd49179, 16'd21470, 16'd54146, 16'd34027, 16'd17167, 16'd26039, 16'd56393, 16'd51215});
	test_expansion(128'h01fbfc146ce9e594f5731ad1a2edcb07, {16'd15236, 16'd39835, 16'd37339, 16'd5450, 16'd42963, 16'd34994, 16'd37641, 16'd7516, 16'd37134, 16'd3995, 16'd989, 16'd33175, 16'd19901, 16'd8179, 16'd28011, 16'd27844, 16'd10413, 16'd57383, 16'd59024, 16'd20217, 16'd13390, 16'd33369, 16'd64237, 16'd21298, 16'd47500, 16'd38627});
	test_expansion(128'h85928b9d4cdb14920ca1adc35beacc02, {16'd10504, 16'd21472, 16'd11868, 16'd52901, 16'd28736, 16'd35096, 16'd64649, 16'd9007, 16'd28973, 16'd50882, 16'd39235, 16'd32630, 16'd37427, 16'd21673, 16'd39586, 16'd55335, 16'd2840, 16'd7046, 16'd6225, 16'd14888, 16'd28402, 16'd32674, 16'd17975, 16'd16003, 16'd50690, 16'd44512});
	test_expansion(128'he46d0bd71016dfdfff2dc8e7567e0a4a, {16'd63425, 16'd39211, 16'd65447, 16'd32411, 16'd63433, 16'd43113, 16'd59023, 16'd34632, 16'd35273, 16'd62531, 16'd51558, 16'd18741, 16'd58464, 16'd42745, 16'd14797, 16'd51683, 16'd45816, 16'd54714, 16'd11330, 16'd61595, 16'd9220, 16'd20498, 16'd7561, 16'd55852, 16'd33330, 16'd31573});
	test_expansion(128'h859fa6c50254abacfb8ee103acc66ab4, {16'd57852, 16'd5822, 16'd28393, 16'd40691, 16'd12431, 16'd21362, 16'd39120, 16'd31265, 16'd11605, 16'd21466, 16'd6055, 16'd25467, 16'd39485, 16'd29772, 16'd53144, 16'd33930, 16'd15089, 16'd57848, 16'd18621, 16'd46040, 16'd6157, 16'd59032, 16'd62526, 16'd6167, 16'd1737, 16'd754});
	test_expansion(128'h3306aa4f4ce7b299506a262e7a74aea6, {16'd61221, 16'd22553, 16'd33395, 16'd38248, 16'd17108, 16'd8460, 16'd23607, 16'd36126, 16'd57758, 16'd17941, 16'd40216, 16'd22428, 16'd39680, 16'd64589, 16'd10220, 16'd18705, 16'd44264, 16'd60828, 16'd61076, 16'd7905, 16'd64006, 16'd61083, 16'd36009, 16'd16142, 16'd22406, 16'd48932});
	test_expansion(128'hec9f796360d7c717c192cdcb598d8fd4, {16'd57566, 16'd6336, 16'd19674, 16'd47099, 16'd60530, 16'd55296, 16'd5969, 16'd21667, 16'd62063, 16'd35626, 16'd63251, 16'd46254, 16'd59015, 16'd55301, 16'd22190, 16'd53346, 16'd17909, 16'd35761, 16'd58277, 16'd37122, 16'd29197, 16'd2222, 16'd17241, 16'd28024, 16'd42598, 16'd60826});
	test_expansion(128'h6298be542b14447ad427bc849be4c861, {16'd52880, 16'd23768, 16'd5019, 16'd11214, 16'd12858, 16'd52238, 16'd17169, 16'd61575, 16'd22824, 16'd59601, 16'd4765, 16'd40513, 16'd9917, 16'd26207, 16'd31322, 16'd20552, 16'd38357, 16'd40182, 16'd52049, 16'd36764, 16'd29753, 16'd2929, 16'd59578, 16'd37594, 16'd42436, 16'd57861});
	test_expansion(128'h607c0374d65d0beba04d38e0e2c9d2ab, {16'd38499, 16'd15973, 16'd48470, 16'd64966, 16'd44806, 16'd50759, 16'd54900, 16'd55893, 16'd55610, 16'd41690, 16'd50097, 16'd49864, 16'd36601, 16'd31296, 16'd61456, 16'd29412, 16'd33936, 16'd13820, 16'd36444, 16'd15097, 16'd41318, 16'd62173, 16'd6721, 16'd47083, 16'd49589, 16'd26290});
	test_expansion(128'h2b2eb385d94c2cc04dbb129ad9144f9a, {16'd65068, 16'd29525, 16'd6223, 16'd22922, 16'd34966, 16'd1626, 16'd50554, 16'd61323, 16'd6850, 16'd28271, 16'd13553, 16'd25403, 16'd18539, 16'd58924, 16'd55520, 16'd36604, 16'd17524, 16'd48573, 16'd64674, 16'd57607, 16'd1458, 16'd1842, 16'd2344, 16'd16639, 16'd40378, 16'd4268});
	test_expansion(128'h977246a37353ebb4e58c1110d70af609, {16'd27426, 16'd44587, 16'd20481, 16'd18537, 16'd2301, 16'd29749, 16'd51773, 16'd3642, 16'd32322, 16'd9655, 16'd61145, 16'd2120, 16'd22108, 16'd33690, 16'd41531, 16'd45635, 16'd54001, 16'd11703, 16'd43346, 16'd33693, 16'd22399, 16'd29015, 16'd11788, 16'd53885, 16'd49487, 16'd13639});
	test_expansion(128'h0069cd6ae6a7c1ede53863b3a13654f8, {16'd13228, 16'd34762, 16'd6024, 16'd50320, 16'd431, 16'd23948, 16'd40860, 16'd36888, 16'd48884, 16'd51174, 16'd41803, 16'd1674, 16'd53954, 16'd1230, 16'd32511, 16'd17142, 16'd31721, 16'd53238, 16'd25737, 16'd29849, 16'd41107, 16'd39768, 16'd19135, 16'd24277, 16'd38474, 16'd6802});
	test_expansion(128'h5bc49547e069a9c6b8e9df6b8c48d0e9, {16'd22779, 16'd38009, 16'd25964, 16'd8917, 16'd26899, 16'd63991, 16'd54322, 16'd6229, 16'd55983, 16'd24772, 16'd19238, 16'd19266, 16'd61642, 16'd56051, 16'd63097, 16'd19412, 16'd15181, 16'd44047, 16'd22369, 16'd45167, 16'd37088, 16'd30824, 16'd54649, 16'd5562, 16'd13364, 16'd25096});
	test_expansion(128'haaf02d322b99484e17a9cf2dde559486, {16'd47476, 16'd45839, 16'd19825, 16'd3723, 16'd47617, 16'd44846, 16'd10821, 16'd17204, 16'd48736, 16'd40437, 16'd28500, 16'd582, 16'd17658, 16'd23334, 16'd27288, 16'd28737, 16'd31937, 16'd59034, 16'd35377, 16'd13091, 16'd45078, 16'd27272, 16'd59156, 16'd39490, 16'd56351, 16'd23037});
	test_expansion(128'h29b41b9624cf799e09ac84eefb07a55e, {16'd10675, 16'd22130, 16'd32330, 16'd30952, 16'd35538, 16'd48263, 16'd58614, 16'd11984, 16'd60053, 16'd59932, 16'd32588, 16'd38760, 16'd13346, 16'd15495, 16'd62861, 16'd26043, 16'd29624, 16'd8467, 16'd37721, 16'd54716, 16'd12070, 16'd28253, 16'd63330, 16'd57009, 16'd14569, 16'd48922});
	test_expansion(128'h428daa5479efc2e820eabc64ee661f3b, {16'd65323, 16'd11152, 16'd25894, 16'd20820, 16'd35798, 16'd31377, 16'd7051, 16'd1020, 16'd10451, 16'd31628, 16'd33001, 16'd40915, 16'd27960, 16'd40008, 16'd19784, 16'd47726, 16'd8821, 16'd34001, 16'd54198, 16'd2601, 16'd47700, 16'd37009, 16'd29236, 16'd9564, 16'd56821, 16'd64348});
	test_expansion(128'h53515c5f3fe1c63d39dd1614da24ba5a, {16'd5194, 16'd46840, 16'd31938, 16'd19954, 16'd61310, 16'd32935, 16'd50330, 16'd62792, 16'd11187, 16'd53998, 16'd24841, 16'd63183, 16'd22649, 16'd53190, 16'd64516, 16'd58689, 16'd57077, 16'd31116, 16'd3352, 16'd10419, 16'd14235, 16'd24647, 16'd45991, 16'd6709, 16'd59057, 16'd11609});
	test_expansion(128'hb500cb7fb33d8a1b859400d75378c5e9, {16'd63671, 16'd58202, 16'd36064, 16'd36402, 16'd47548, 16'd13942, 16'd14494, 16'd19032, 16'd17890, 16'd37194, 16'd7500, 16'd53362, 16'd56968, 16'd64212, 16'd4161, 16'd8279, 16'd3181, 16'd31013, 16'd6275, 16'd42271, 16'd9098, 16'd64616, 16'd47881, 16'd8769, 16'd29394, 16'd11476});
	test_expansion(128'hec64b08db05943cc3cef8017861f17a0, {16'd8826, 16'd9824, 16'd60197, 16'd60406, 16'd25479, 16'd63483, 16'd51516, 16'd2484, 16'd30626, 16'd54387, 16'd17709, 16'd9163, 16'd57744, 16'd42751, 16'd53966, 16'd16434, 16'd60367, 16'd40572, 16'd25412, 16'd43695, 16'd3596, 16'd36334, 16'd48868, 16'd9915, 16'd61414, 16'd30757});
	test_expansion(128'h0e64b9b4450e558fd998289a40cc0301, {16'd31011, 16'd62858, 16'd53164, 16'd3644, 16'd45139, 16'd59254, 16'd19256, 16'd8569, 16'd58237, 16'd53883, 16'd60973, 16'd56228, 16'd62363, 16'd42045, 16'd24030, 16'd813, 16'd18376, 16'd6456, 16'd7394, 16'd22000, 16'd10885, 16'd64142, 16'd27937, 16'd5745, 16'd22190, 16'd34195});
	test_expansion(128'h71dc7003df8833ed2eb1b666c128cd1f, {16'd26612, 16'd5086, 16'd58954, 16'd57349, 16'd25876, 16'd19148, 16'd12071, 16'd156, 16'd60542, 16'd54847, 16'd2712, 16'd29893, 16'd62109, 16'd15962, 16'd49920, 16'd62397, 16'd51831, 16'd51456, 16'd64225, 16'd8204, 16'd49672, 16'd43984, 16'd40826, 16'd11989, 16'd57776, 16'd15716});
	test_expansion(128'h16d1742161a215aab3b0597f1851610f, {16'd28254, 16'd60282, 16'd27852, 16'd31969, 16'd22845, 16'd12229, 16'd57114, 16'd65448, 16'd35749, 16'd34727, 16'd2686, 16'd32021, 16'd6940, 16'd15501, 16'd50667, 16'd39842, 16'd48038, 16'd6237, 16'd47862, 16'd41961, 16'd26082, 16'd30789, 16'd10795, 16'd55569, 16'd49272, 16'd55334});
	test_expansion(128'h33a2986814471f69503f8ad57a8b36b1, {16'd36249, 16'd55707, 16'd44262, 16'd57070, 16'd34103, 16'd647, 16'd26627, 16'd64801, 16'd2474, 16'd52080, 16'd51867, 16'd27096, 16'd54057, 16'd32028, 16'd54935, 16'd17962, 16'd37257, 16'd26860, 16'd25996, 16'd10896, 16'd21304, 16'd16403, 16'd41710, 16'd15539, 16'd56384, 16'd33460});
	test_expansion(128'h7b68dd2ff088c3f493ca247aa2136d4a, {16'd61342, 16'd58391, 16'd31103, 16'd11342, 16'd48032, 16'd38440, 16'd17012, 16'd37150, 16'd60980, 16'd50676, 16'd5471, 16'd43991, 16'd40794, 16'd33893, 16'd24650, 16'd6281, 16'd9536, 16'd7474, 16'd38940, 16'd43884, 16'd32941, 16'd11396, 16'd63415, 16'd58433, 16'd41661, 16'd44217});
	test_expansion(128'h4ade8e9e94aac1e3536827544d181cb5, {16'd64334, 16'd28286, 16'd9718, 16'd63434, 16'd55213, 16'd58577, 16'd45979, 16'd2166, 16'd308, 16'd14543, 16'd54331, 16'd47409, 16'd46761, 16'd62859, 16'd20911, 16'd14062, 16'd11294, 16'd60692, 16'd39628, 16'd30166, 16'd14044, 16'd21459, 16'd33661, 16'd44731, 16'd14553, 16'd6643});
	test_expansion(128'hb5e99e6312a99e8bbf9f3eb8797fd7aa, {16'd59871, 16'd41017, 16'd50985, 16'd5086, 16'd47874, 16'd46189, 16'd53229, 16'd63145, 16'd46760, 16'd17263, 16'd54870, 16'd42582, 16'd30569, 16'd53513, 16'd41153, 16'd64834, 16'd30974, 16'd45661, 16'd62224, 16'd34045, 16'd17700, 16'd7738, 16'd17511, 16'd20952, 16'd30286, 16'd37231});
	test_expansion(128'hc62d19e9fe5ee61e9232399dfd08c3ec, {16'd6616, 16'd26024, 16'd14921, 16'd25542, 16'd57655, 16'd20144, 16'd5113, 16'd31502, 16'd20513, 16'd31065, 16'd5961, 16'd48352, 16'd32748, 16'd27728, 16'd5136, 16'd63701, 16'd32861, 16'd42676, 16'd53559, 16'd26855, 16'd49075, 16'd19486, 16'd33230, 16'd31858, 16'd60685, 16'd56205});
	test_expansion(128'h7efe401150f7966636e747ce20c8214b, {16'd61780, 16'd11377, 16'd65246, 16'd33699, 16'd28086, 16'd29798, 16'd52645, 16'd49776, 16'd38074, 16'd3248, 16'd53807, 16'd27808, 16'd25227, 16'd24358, 16'd23133, 16'd12290, 16'd43301, 16'd36639, 16'd31488, 16'd54151, 16'd44660, 16'd41389, 16'd47779, 16'd20969, 16'd58089, 16'd3247});
	test_expansion(128'h1b054e55c444258729d8aeef83c841e2, {16'd52878, 16'd54570, 16'd10633, 16'd19835, 16'd22100, 16'd2520, 16'd45357, 16'd47660, 16'd32461, 16'd34967, 16'd18545, 16'd8414, 16'd53480, 16'd17325, 16'd30407, 16'd49300, 16'd54177, 16'd1334, 16'd33806, 16'd64219, 16'd27444, 16'd28568, 16'd42316, 16'd33113, 16'd4691, 16'd59449});
	test_expansion(128'h42633854809c4707c4991d6e510181ae, {16'd9225, 16'd3523, 16'd51593, 16'd2350, 16'd17806, 16'd50423, 16'd15890, 16'd13750, 16'd6658, 16'd7906, 16'd11135, 16'd21267, 16'd64617, 16'd48409, 16'd3173, 16'd28623, 16'd2661, 16'd58711, 16'd49522, 16'd544, 16'd623, 16'd65335, 16'd5577, 16'd4882, 16'd38959, 16'd30018});
	test_expansion(128'hc19bcfbb4a36d5af5554d2e63a4880e5, {16'd7234, 16'd62798, 16'd44925, 16'd28740, 16'd25539, 16'd1300, 16'd61078, 16'd26084, 16'd38243, 16'd57002, 16'd17299, 16'd51805, 16'd55238, 16'd4902, 16'd8959, 16'd17037, 16'd35328, 16'd54110, 16'd2140, 16'd54159, 16'd59654, 16'd31296, 16'd61908, 16'd40084, 16'd38232, 16'd23213});
	test_expansion(128'hbb3a3dfbe79e7167cd743ee81bc0c89f, {16'd39508, 16'd41483, 16'd26586, 16'd63785, 16'd33227, 16'd43917, 16'd54311, 16'd26228, 16'd48739, 16'd42439, 16'd33463, 16'd2187, 16'd59874, 16'd59227, 16'd27260, 16'd50870, 16'd54436, 16'd15822, 16'd63696, 16'd20628, 16'd63180, 16'd9820, 16'd39851, 16'd63081, 16'd51284, 16'd45471});
	test_expansion(128'h88868713146abc05c0fbf285920d19db, {16'd47688, 16'd53224, 16'd36901, 16'd38611, 16'd58974, 16'd37758, 16'd44945, 16'd23148, 16'd62605, 16'd8535, 16'd40919, 16'd819, 16'd15413, 16'd57337, 16'd14125, 16'd50214, 16'd27507, 16'd41796, 16'd51295, 16'd24179, 16'd43886, 16'd17232, 16'd6092, 16'd41378, 16'd15712, 16'd18836});
	test_expansion(128'hdb6edefb2cfdbaebc06040bbd8b4910a, {16'd19164, 16'd28354, 16'd6737, 16'd1426, 16'd64285, 16'd42459, 16'd35188, 16'd6554, 16'd20633, 16'd56786, 16'd41705, 16'd15250, 16'd1683, 16'd26536, 16'd20028, 16'd51400, 16'd63944, 16'd63037, 16'd12361, 16'd33415, 16'd3146, 16'd44497, 16'd24309, 16'd42422, 16'd60729, 16'd64776});
	test_expansion(128'h2988f6181a23db3047ab1d63e21a0d2e, {16'd44888, 16'd22606, 16'd21135, 16'd55250, 16'd54346, 16'd42863, 16'd22453, 16'd24830, 16'd16451, 16'd35097, 16'd29570, 16'd15070, 16'd18069, 16'd36494, 16'd64610, 16'd665, 16'd12966, 16'd63782, 16'd30415, 16'd9764, 16'd27148, 16'd747, 16'd54160, 16'd3710, 16'd50987, 16'd45758});
	test_expansion(128'hbe4b8750b3a9cfef012c3afceff11024, {16'd45604, 16'd19463, 16'd14935, 16'd46188, 16'd40561, 16'd28696, 16'd59943, 16'd50112, 16'd6913, 16'd2890, 16'd45454, 16'd34855, 16'd3677, 16'd21833, 16'd13778, 16'd54076, 16'd64081, 16'd9174, 16'd56732, 16'd44846, 16'd63576, 16'd10449, 16'd32459, 16'd38749, 16'd2040, 16'd20742});
	test_expansion(128'h5d929d869e56c3f6de52b9c83136c80f, {16'd55979, 16'd44703, 16'd49332, 16'd31302, 16'd8195, 16'd33424, 16'd11455, 16'd49096, 16'd60028, 16'd58980, 16'd19357, 16'd4766, 16'd31456, 16'd7799, 16'd23339, 16'd15411, 16'd23786, 16'd21828, 16'd1357, 16'd47601, 16'd42506, 16'd33104, 16'd57584, 16'd19079, 16'd62296, 16'd62908});
	test_expansion(128'h1c8679cc84ca6ba14e6298662f3122ac, {16'd5796, 16'd36419, 16'd38341, 16'd19854, 16'd4094, 16'd49024, 16'd58773, 16'd1689, 16'd27982, 16'd21816, 16'd43377, 16'd18924, 16'd26881, 16'd40868, 16'd41679, 16'd15882, 16'd14860, 16'd13632, 16'd28381, 16'd56328, 16'd32512, 16'd33627, 16'd60193, 16'd22472, 16'd6299, 16'd10838});
	test_expansion(128'ha8b3f208321620d92b28ac815fc65216, {16'd34629, 16'd43619, 16'd6063, 16'd25613, 16'd38928, 16'd59270, 16'd60569, 16'd37836, 16'd5827, 16'd30967, 16'd40825, 16'd36947, 16'd20509, 16'd6467, 16'd20048, 16'd34212, 16'd52422, 16'd41590, 16'd27475, 16'd15114, 16'd56873, 16'd52905, 16'd47748, 16'd49026, 16'd16303, 16'd56013});
	test_expansion(128'h43579fa1f63e2b5574b75135771a4af1, {16'd23957, 16'd52837, 16'd1036, 16'd25653, 16'd6175, 16'd26991, 16'd44673, 16'd49052, 16'd23371, 16'd34733, 16'd47426, 16'd49051, 16'd30466, 16'd28428, 16'd53878, 16'd10029, 16'd32556, 16'd26886, 16'd9346, 16'd6374, 16'd24593, 16'd62004, 16'd2841, 16'd5544, 16'd65058, 16'd22770});
	test_expansion(128'hb2cefd677ca49250b7dbed48cb8c9e85, {16'd5212, 16'd43197, 16'd6055, 16'd32015, 16'd31887, 16'd12535, 16'd65048, 16'd43593, 16'd50620, 16'd250, 16'd45769, 16'd27024, 16'd52825, 16'd45810, 16'd45661, 16'd24095, 16'd60920, 16'd61210, 16'd2566, 16'd44100, 16'd51693, 16'd47143, 16'd56093, 16'd62062, 16'd760, 16'd41047});
	test_expansion(128'hebfc0facc2e27f6cfc1e824612dbeafa, {16'd2360, 16'd65277, 16'd17321, 16'd22289, 16'd40413, 16'd14948, 16'd17483, 16'd54732, 16'd49606, 16'd30408, 16'd17809, 16'd43830, 16'd53020, 16'd28350, 16'd2181, 16'd2987, 16'd33681, 16'd9135, 16'd28098, 16'd50165, 16'd44785, 16'd5115, 16'd5867, 16'd41849, 16'd22863, 16'd17420});
	test_expansion(128'h67269437d29d7c957c7f6b1ec5bac017, {16'd7843, 16'd55993, 16'd17854, 16'd18940, 16'd24111, 16'd10034, 16'd52851, 16'd7537, 16'd1558, 16'd64024, 16'd62074, 16'd46618, 16'd34076, 16'd12906, 16'd56692, 16'd55510, 16'd36455, 16'd31022, 16'd37950, 16'd3935, 16'd46296, 16'd18404, 16'd17721, 16'd26246, 16'd33380, 16'd32513});
	test_expansion(128'hfad3621d1b5202487b542e69934f839f, {16'd60796, 16'd2681, 16'd13580, 16'd6707, 16'd58654, 16'd21206, 16'd49027, 16'd13258, 16'd11008, 16'd61811, 16'd43463, 16'd28539, 16'd57134, 16'd10538, 16'd6677, 16'd32671, 16'd37840, 16'd7184, 16'd31397, 16'd8145, 16'd17460, 16'd38421, 16'd61185, 16'd57847, 16'd26678, 16'd7766});
	test_expansion(128'h1786b195d8a73cf81d396b99becc406a, {16'd7440, 16'd62297, 16'd14300, 16'd15219, 16'd13108, 16'd33945, 16'd38891, 16'd5645, 16'd35299, 16'd41368, 16'd12709, 16'd3782, 16'd7741, 16'd42552, 16'd17066, 16'd23889, 16'd47933, 16'd29457, 16'd54426, 16'd21561, 16'd39669, 16'd59117, 16'd7345, 16'd51453, 16'd16897, 16'd12240});
	test_expansion(128'h570000505751fb644dbbdacdfe985af3, {16'd43099, 16'd52260, 16'd12818, 16'd56220, 16'd14514, 16'd60376, 16'd43443, 16'd34451, 16'd15960, 16'd55169, 16'd38045, 16'd683, 16'd9861, 16'd36652, 16'd5162, 16'd41565, 16'd12091, 16'd64919, 16'd29280, 16'd56047, 16'd40264, 16'd61345, 16'd52094, 16'd3342, 16'd58695, 16'd59740});
	test_expansion(128'hd9836a1791d25529b7a80ff5b0b779e2, {16'd36931, 16'd7278, 16'd64393, 16'd63481, 16'd22973, 16'd7364, 16'd6579, 16'd16007, 16'd55002, 16'd47109, 16'd33771, 16'd43701, 16'd20626, 16'd46447, 16'd40004, 16'd10268, 16'd15076, 16'd30324, 16'd53974, 16'd28942, 16'd59985, 16'd58284, 16'd43772, 16'd11297, 16'd56645, 16'd57610});
	test_expansion(128'hd29b99aec25bd9f78923a156f418b817, {16'd699, 16'd30945, 16'd11277, 16'd53998, 16'd52421, 16'd13701, 16'd11304, 16'd29880, 16'd13982, 16'd29461, 16'd19944, 16'd50403, 16'd17794, 16'd41972, 16'd49198, 16'd62574, 16'd50156, 16'd55285, 16'd36221, 16'd48845, 16'd26283, 16'd65268, 16'd38058, 16'd61292, 16'd8279, 16'd32725});
	test_expansion(128'h6479fb9b967d31e8baac66737dcc165d, {16'd41989, 16'd40926, 16'd35896, 16'd49874, 16'd15783, 16'd5002, 16'd27330, 16'd41721, 16'd27989, 16'd45240, 16'd13461, 16'd15973, 16'd13030, 16'd24608, 16'd19464, 16'd65221, 16'd63485, 16'd8037, 16'd61878, 16'd3025, 16'd24172, 16'd22578, 16'd30133, 16'd425, 16'd55387, 16'd48069});
	test_expansion(128'h62fc6901af824c680b6b82ba05432eaa, {16'd12464, 16'd6242, 16'd55941, 16'd33561, 16'd49727, 16'd32688, 16'd12086, 16'd34683, 16'd46440, 16'd32103, 16'd15230, 16'd61666, 16'd45900, 16'd3313, 16'd38897, 16'd22306, 16'd44382, 16'd50624, 16'd52387, 16'd10662, 16'd23071, 16'd8279, 16'd36259, 16'd9547, 16'd7575, 16'd30900});
	test_expansion(128'h99ed4305740a29b6bac2d2ed2303b4f0, {16'd1838, 16'd27686, 16'd51499, 16'd53379, 16'd54343, 16'd12448, 16'd38871, 16'd5675, 16'd16952, 16'd36516, 16'd8589, 16'd43600, 16'd22262, 16'd41264, 16'd42479, 16'd22423, 16'd1211, 16'd23445, 16'd1571, 16'd43399, 16'd46870, 16'd711, 16'd31730, 16'd43167, 16'd31264, 16'd22947});
	test_expansion(128'he68c642e1513b55f8d72cb1b455ca8e6, {16'd11774, 16'd1707, 16'd30305, 16'd10360, 16'd27360, 16'd7388, 16'd24686, 16'd14508, 16'd44219, 16'd36009, 16'd45552, 16'd51154, 16'd9322, 16'd47266, 16'd46159, 16'd6416, 16'd25606, 16'd3124, 16'd46105, 16'd31406, 16'd7045, 16'd13000, 16'd62424, 16'd31088, 16'd11888, 16'd13981});
	test_expansion(128'h60fa7365ba2c854a13dac6838cd87b7a, {16'd54850, 16'd22071, 16'd13418, 16'd44451, 16'd5939, 16'd36015, 16'd61226, 16'd33703, 16'd26277, 16'd47296, 16'd43611, 16'd7011, 16'd2802, 16'd39392, 16'd23608, 16'd44815, 16'd64171, 16'd42750, 16'd759, 16'd11020, 16'd59936, 16'd55818, 16'd65311, 16'd31186, 16'd65229, 16'd57098});
	test_expansion(128'h53295b6a06e3f3ad31e9c421e0bb0544, {16'd9047, 16'd50181, 16'd30522, 16'd10588, 16'd3901, 16'd30692, 16'd60178, 16'd15262, 16'd10020, 16'd24394, 16'd27073, 16'd23070, 16'd30181, 16'd63064, 16'd28821, 16'd34771, 16'd36361, 16'd15110, 16'd53041, 16'd21803, 16'd33607, 16'd1133, 16'd41449, 16'd39642, 16'd3586, 16'd47895});
	test_expansion(128'h912548c6ff0f19dfd2604640123885a7, {16'd16425, 16'd57444, 16'd51900, 16'd14327, 16'd20845, 16'd22119, 16'd56893, 16'd22455, 16'd60045, 16'd39337, 16'd27090, 16'd12769, 16'd45554, 16'd18924, 16'd25895, 16'd16026, 16'd36819, 16'd15907, 16'd34889, 16'd32067, 16'd56856, 16'd20558, 16'd55331, 16'd41169, 16'd33744, 16'd59953});
	test_expansion(128'h285f3780b95f1d874e3f8a14a5a9b723, {16'd35586, 16'd28200, 16'd7166, 16'd31940, 16'd54159, 16'd9093, 16'd49895, 16'd19163, 16'd57360, 16'd57792, 16'd55341, 16'd8749, 16'd30201, 16'd15712, 16'd64958, 16'd47154, 16'd28895, 16'd12019, 16'd51546, 16'd5599, 16'd782, 16'd47640, 16'd6534, 16'd35135, 16'd46549, 16'd65390});
	test_expansion(128'h2723ef72c4dc946ed553a96fb72e2d07, {16'd53711, 16'd16506, 16'd22059, 16'd52936, 16'd9970, 16'd23217, 16'd5859, 16'd63418, 16'd12404, 16'd40447, 16'd18324, 16'd18531, 16'd16185, 16'd61562, 16'd37540, 16'd49358, 16'd48018, 16'd39103, 16'd46461, 16'd51064, 16'd14601, 16'd42045, 16'd33460, 16'd53657, 16'd50902, 16'd21101});
	test_expansion(128'h4e70af54dd0b31b20cb80223e110d4f2, {16'd11027, 16'd37585, 16'd855, 16'd64528, 16'd24809, 16'd37677, 16'd21605, 16'd32740, 16'd8295, 16'd972, 16'd38224, 16'd44298, 16'd44437, 16'd46711, 16'd49115, 16'd39660, 16'd27992, 16'd28642, 16'd38181, 16'd33584, 16'd27838, 16'd6527, 16'd62779, 16'd26918, 16'd32317, 16'd5175});
	test_expansion(128'hf508bf4ba0e110472242d4620a0515c9, {16'd32227, 16'd27051, 16'd12435, 16'd18045, 16'd8567, 16'd45987, 16'd787, 16'd22429, 16'd26141, 16'd62908, 16'd24749, 16'd57362, 16'd49595, 16'd17876, 16'd54602, 16'd28644, 16'd11318, 16'd30019, 16'd59939, 16'd58473, 16'd22201, 16'd22891, 16'd10412, 16'd49099, 16'd9364, 16'd1416});
	test_expansion(128'hb224089c7a92f37d1b39ad15a060831a, {16'd17097, 16'd3001, 16'd47330, 16'd37566, 16'd12561, 16'd7842, 16'd35624, 16'd51224, 16'd24753, 16'd961, 16'd39458, 16'd9513, 16'd58577, 16'd26129, 16'd140, 16'd60364, 16'd46944, 16'd19959, 16'd44975, 16'd20560, 16'd10442, 16'd35021, 16'd55082, 16'd13641, 16'd17018, 16'd7079});
	test_expansion(128'hf272a6a2dfbb63b141a121d2be2e6abe, {16'd10251, 16'd63653, 16'd29037, 16'd12257, 16'd18062, 16'd8352, 16'd60358, 16'd25970, 16'd53931, 16'd11863, 16'd21638, 16'd50998, 16'd57651, 16'd47515, 16'd5168, 16'd13828, 16'd27365, 16'd45760, 16'd8917, 16'd58214, 16'd36387, 16'd36111, 16'd28838, 16'd28986, 16'd17702, 16'd9424});
	test_expansion(128'h0f70c023ae85eb581925e3c5c552b779, {16'd49760, 16'd38429, 16'd2531, 16'd27840, 16'd30284, 16'd64953, 16'd19558, 16'd56985, 16'd1136, 16'd1732, 16'd47026, 16'd61786, 16'd32746, 16'd23966, 16'd29766, 16'd2286, 16'd33960, 16'd45111, 16'd63870, 16'd6757, 16'd4443, 16'd22678, 16'd20891, 16'd60970, 16'd23856, 16'd18725});
	test_expansion(128'had2dfd08333d729aa488211c2dcc08c1, {16'd57376, 16'd53384, 16'd29403, 16'd45710, 16'd47892, 16'd37339, 16'd48222, 16'd7125, 16'd63151, 16'd4031, 16'd46384, 16'd24688, 16'd1777, 16'd16157, 16'd26427, 16'd45052, 16'd46418, 16'd44222, 16'd59777, 16'd51134, 16'd31113, 16'd26963, 16'd12803, 16'd23170, 16'd16267, 16'd32851});
	test_expansion(128'h25741f5eb8919914f765817a753b392e, {16'd37259, 16'd10516, 16'd26399, 16'd34378, 16'd8195, 16'd42297, 16'd7770, 16'd11159, 16'd62647, 16'd34762, 16'd32321, 16'd32704, 16'd39012, 16'd11138, 16'd42282, 16'd59604, 16'd24344, 16'd60287, 16'd65330, 16'd22952, 16'd19848, 16'd25065, 16'd1797, 16'd63004, 16'd19854, 16'd3061});
	test_expansion(128'h331309ab322c6c9cc6216bea085bdcc5, {16'd54230, 16'd53754, 16'd15753, 16'd25595, 16'd54791, 16'd1035, 16'd10107, 16'd61546, 16'd10141, 16'd9646, 16'd23051, 16'd750, 16'd31174, 16'd4054, 16'd13405, 16'd46819, 16'd61289, 16'd51249, 16'd22487, 16'd41533, 16'd63861, 16'd37311, 16'd22601, 16'd58046, 16'd40661, 16'd31463});
	test_expansion(128'h6bb385858644ae0590fd162ec785ddec, {16'd25613, 16'd33296, 16'd24587, 16'd10783, 16'd21103, 16'd27596, 16'd44459, 16'd61139, 16'd55959, 16'd42783, 16'd26723, 16'd11299, 16'd20953, 16'd1324, 16'd42777, 16'd56840, 16'd25168, 16'd46901, 16'd43264, 16'd39184, 16'd51359, 16'd41728, 16'd1258, 16'd24965, 16'd11183, 16'd22928});
	test_expansion(128'hdfc3641a8fc2564842de4ea74e4c9469, {16'd23532, 16'd62902, 16'd19511, 16'd54836, 16'd9525, 16'd52130, 16'd63904, 16'd37568, 16'd36358, 16'd50799, 16'd39813, 16'd44242, 16'd19030, 16'd14704, 16'd27124, 16'd20605, 16'd42083, 16'd7503, 16'd61731, 16'd61324, 16'd38164, 16'd35453, 16'd43778, 16'd50620, 16'd1408, 16'd37777});
	test_expansion(128'hd27200054265a51b48790d79a373ba37, {16'd12135, 16'd843, 16'd55242, 16'd64972, 16'd1169, 16'd56070, 16'd64789, 16'd50698, 16'd37003, 16'd63871, 16'd6070, 16'd51218, 16'd22645, 16'd55788, 16'd38192, 16'd9263, 16'd55380, 16'd63510, 16'd5524, 16'd62010, 16'd14372, 16'd48263, 16'd41565, 16'd14117, 16'd33443, 16'd47256});
	test_expansion(128'h6c08890524184c3b7924ea1c6448d4ab, {16'd52606, 16'd41571, 16'd9032, 16'd4901, 16'd29607, 16'd22233, 16'd7882, 16'd64433, 16'd1690, 16'd23800, 16'd47734, 16'd35984, 16'd5165, 16'd52809, 16'd29797, 16'd51467, 16'd22983, 16'd695, 16'd56102, 16'd47784, 16'd61810, 16'd31403, 16'd30952, 16'd11309, 16'd4117, 16'd7608});
	test_expansion(128'h15091a98bb2b6d1133a1e880f615c215, {16'd59264, 16'd5434, 16'd27964, 16'd38836, 16'd28648, 16'd9143, 16'd63413, 16'd51759, 16'd60376, 16'd36624, 16'd58667, 16'd48345, 16'd19706, 16'd59076, 16'd41513, 16'd47263, 16'd20550, 16'd27226, 16'd17073, 16'd47164, 16'd14743, 16'd54895, 16'd64686, 16'd59652, 16'd63362, 16'd56543});
	test_expansion(128'h0dabf4fa64af0e9cf7e32f5d3c0d6cfe, {16'd25492, 16'd38781, 16'd8569, 16'd8873, 16'd61642, 16'd25621, 16'd14746, 16'd23503, 16'd22292, 16'd46708, 16'd26014, 16'd37441, 16'd56797, 16'd37908, 16'd61288, 16'd31247, 16'd59157, 16'd43778, 16'd65144, 16'd59815, 16'd23204, 16'd303, 16'd49487, 16'd50677, 16'd60023, 16'd61512});
	test_expansion(128'h821961f8977220fc4fb1f8c0b91718a5, {16'd39135, 16'd59405, 16'd22033, 16'd10337, 16'd38714, 16'd9446, 16'd38353, 16'd51501, 16'd36972, 16'd47374, 16'd63928, 16'd49529, 16'd59630, 16'd9950, 16'd40601, 16'd86, 16'd65254, 16'd60778, 16'd61509, 16'd17504, 16'd48283, 16'd13287, 16'd14344, 16'd62241, 16'd36612, 16'd30514});
	test_expansion(128'h6fa5ec86123dde676eb7a071a4f08036, {16'd12589, 16'd65123, 16'd19038, 16'd1727, 16'd48672, 16'd23827, 16'd36566, 16'd52167, 16'd24018, 16'd38934, 16'd64731, 16'd63786, 16'd24951, 16'd57715, 16'd908, 16'd18123, 16'd57713, 16'd8231, 16'd5542, 16'd25750, 16'd41457, 16'd42432, 16'd25761, 16'd63954, 16'd34678, 16'd42793});
	test_expansion(128'h5d6a5b80d9653be0a4b7fade39385952, {16'd27084, 16'd41299, 16'd20582, 16'd31061, 16'd43667, 16'd2917, 16'd61330, 16'd3011, 16'd57217, 16'd15716, 16'd9255, 16'd5206, 16'd62975, 16'd58827, 16'd35417, 16'd23162, 16'd56543, 16'd35334, 16'd3617, 16'd57391, 16'd6074, 16'd56305, 16'd51117, 16'd23544, 16'd30316, 16'd27246});
	test_expansion(128'h036a3602b2b1fd5a746f5039b84971be, {16'd47151, 16'd10371, 16'd63223, 16'd39218, 16'd52346, 16'd37270, 16'd56581, 16'd5687, 16'd19029, 16'd5003, 16'd47018, 16'd18496, 16'd34331, 16'd2064, 16'd24348, 16'd19064, 16'd25468, 16'd49906, 16'd35737, 16'd25696, 16'd44994, 16'd3220, 16'd3919, 16'd48, 16'd21940, 16'd7580});
	test_expansion(128'hde036872a2e0bd6e22ac3a24e9bbdb7e, {16'd33760, 16'd16708, 16'd25204, 16'd11100, 16'd63205, 16'd31862, 16'd10574, 16'd29242, 16'd35963, 16'd31113, 16'd15159, 16'd27841, 16'd8437, 16'd26868, 16'd28687, 16'd131, 16'd26002, 16'd54488, 16'd29045, 16'd49255, 16'd63990, 16'd28517, 16'd59777, 16'd13776, 16'd14998, 16'd46115});
	test_expansion(128'hca9ed1937d07010393aedd937dab45c2, {16'd33006, 16'd21423, 16'd32089, 16'd34198, 16'd21649, 16'd40699, 16'd16269, 16'd36068, 16'd20732, 16'd5646, 16'd27106, 16'd44591, 16'd56500, 16'd28710, 16'd47038, 16'd27110, 16'd18232, 16'd56152, 16'd31909, 16'd7821, 16'd63797, 16'd63059, 16'd43600, 16'd58760, 16'd46982, 16'd24273});
	test_expansion(128'h2714efc628ae741d23389323eeeac233, {16'd48653, 16'd50109, 16'd2944, 16'd44264, 16'd60659, 16'd26917, 16'd6706, 16'd43146, 16'd58319, 16'd5349, 16'd35960, 16'd34146, 16'd55637, 16'd24009, 16'd30768, 16'd60512, 16'd60540, 16'd18197, 16'd16048, 16'd27066, 16'd59695, 16'd18339, 16'd26966, 16'd57443, 16'd10033, 16'd16279});
	test_expansion(128'h54ad4281929f3344041dfe104b4be44f, {16'd46303, 16'd34469, 16'd28144, 16'd36966, 16'd15602, 16'd42017, 16'd18811, 16'd61655, 16'd62778, 16'd39668, 16'd59748, 16'd34448, 16'd53039, 16'd22613, 16'd40168, 16'd54155, 16'd54408, 16'd56870, 16'd58027, 16'd53631, 16'd45228, 16'd17016, 16'd30331, 16'd9385, 16'd27699, 16'd45040});
	test_expansion(128'hc3dbef4bfac8ad85999401d2b231a738, {16'd59801, 16'd7629, 16'd14505, 16'd35568, 16'd51109, 16'd44060, 16'd9448, 16'd31013, 16'd10155, 16'd44068, 16'd42049, 16'd5497, 16'd46459, 16'd53748, 16'd7411, 16'd39222, 16'd4911, 16'd43686, 16'd48641, 16'd62502, 16'd20699, 16'd44739, 16'd30531, 16'd53638, 16'd19600, 16'd37794});
	test_expansion(128'h934a25ad3dd1617ce6f771d5f9c74616, {16'd23370, 16'd31508, 16'd34631, 16'd40595, 16'd61461, 16'd2563, 16'd17141, 16'd22034, 16'd47053, 16'd24722, 16'd51156, 16'd56506, 16'd48506, 16'd3061, 16'd11755, 16'd28656, 16'd42107, 16'd30451, 16'd51646, 16'd15061, 16'd42882, 16'd16251, 16'd20001, 16'd22389, 16'd41429, 16'd63185});
	test_expansion(128'h1e88572c043cb3ab0f88b4ba394ec6d3, {16'd50851, 16'd3934, 16'd59895, 16'd51722, 16'd60993, 16'd10419, 16'd58913, 16'd19368, 16'd27967, 16'd13953, 16'd44067, 16'd28854, 16'd38009, 16'd4130, 16'd64529, 16'd1262, 16'd22, 16'd43373, 16'd62403, 16'd30227, 16'd10113, 16'd41229, 16'd29077, 16'd8944, 16'd19389, 16'd57255});
	test_expansion(128'h44fb5f5153596834bea53167a8eded5f, {16'd54171, 16'd45192, 16'd54068, 16'd14580, 16'd29648, 16'd29255, 16'd40850, 16'd21621, 16'd12057, 16'd64069, 16'd3721, 16'd39270, 16'd4840, 16'd10662, 16'd23115, 16'd29027, 16'd58907, 16'd10824, 16'd55405, 16'd47750, 16'd16659, 16'd55750, 16'd61081, 16'd49664, 16'd54487, 16'd54957});
	test_expansion(128'h6b5e711fa550adf1ef7b9c74733b188d, {16'd38946, 16'd29878, 16'd1333, 16'd42373, 16'd19547, 16'd54480, 16'd42927, 16'd58024, 16'd10894, 16'd28424, 16'd43805, 16'd55043, 16'd12219, 16'd37722, 16'd16317, 16'd41285, 16'd39694, 16'd12553, 16'd59329, 16'd59323, 16'd60072, 16'd45520, 16'd10174, 16'd60558, 16'd55566, 16'd64702});
	test_expansion(128'h93b8db6f1cd6f5a050207bd74e9c64f5, {16'd40040, 16'd17708, 16'd3760, 16'd25758, 16'd41436, 16'd5303, 16'd36989, 16'd2733, 16'd4885, 16'd34617, 16'd54493, 16'd29814, 16'd10799, 16'd8746, 16'd9811, 16'd31581, 16'd8109, 16'd15539, 16'd5943, 16'd24674, 16'd20919, 16'd9825, 16'd13235, 16'd6316, 16'd53133, 16'd55705});
	test_expansion(128'h1b54de07a78cebd3e6a34e356a97e32d, {16'd55368, 16'd60592, 16'd37168, 16'd1315, 16'd65459, 16'd4981, 16'd22194, 16'd16553, 16'd10264, 16'd8150, 16'd41340, 16'd48122, 16'd30663, 16'd27869, 16'd52230, 16'd65397, 16'd25758, 16'd6799, 16'd4506, 16'd44585, 16'd9178, 16'd43823, 16'd61116, 16'd16370, 16'd15994, 16'd17658});
	test_expansion(128'hd1a7a99b05e89d70bdc5766b7d0ac2d8, {16'd25552, 16'd8088, 16'd17408, 16'd31473, 16'd15723, 16'd23742, 16'd15321, 16'd52994, 16'd38697, 16'd63307, 16'd13105, 16'd4409, 16'd38830, 16'd12788, 16'd32448, 16'd43097, 16'd22451, 16'd63188, 16'd62125, 16'd60859, 16'd34491, 16'd26506, 16'd53184, 16'd34290, 16'd32339, 16'd1880});
	test_expansion(128'ha089997a1be7ddea2a9758cb776a6d78, {16'd44437, 16'd19004, 16'd63374, 16'd10, 16'd28, 16'd62226, 16'd32810, 16'd17374, 16'd49289, 16'd34180, 16'd64272, 16'd36058, 16'd26055, 16'd1815, 16'd35043, 16'd21361, 16'd109, 16'd60915, 16'd23612, 16'd50168, 16'd15713, 16'd63718, 16'd27271, 16'd63265, 16'd31519, 16'd6128});
	test_expansion(128'h8e34eb653251fe0b51058f707bb2776f, {16'd20633, 16'd26294, 16'd38805, 16'd6775, 16'd62738, 16'd39756, 16'd14155, 16'd27861, 16'd61615, 16'd15717, 16'd64427, 16'd5850, 16'd44219, 16'd14700, 16'd12171, 16'd43565, 16'd57924, 16'd64974, 16'd3128, 16'd11222, 16'd29721, 16'd31524, 16'd61887, 16'd42370, 16'd2137, 16'd62702});
	test_expansion(128'hca250e1fb3b369927efdd2a27ca3e29d, {16'd3172, 16'd23207, 16'd5392, 16'd59772, 16'd25069, 16'd63411, 16'd7017, 16'd33446, 16'd16165, 16'd42449, 16'd63006, 16'd16765, 16'd25175, 16'd17512, 16'd44489, 16'd23390, 16'd47340, 16'd60268, 16'd45338, 16'd53853, 16'd53324, 16'd21065, 16'd41521, 16'd1276, 16'd8321, 16'd21023});
	test_expansion(128'h9e10ac757136582247bb1867fd3ccba9, {16'd55375, 16'd37817, 16'd13056, 16'd14342, 16'd24668, 16'd52095, 16'd10954, 16'd47259, 16'd350, 16'd6025, 16'd4248, 16'd42743, 16'd32320, 16'd51569, 16'd44734, 16'd23946, 16'd32369, 16'd48921, 16'd13377, 16'd23801, 16'd54526, 16'd15140, 16'd27986, 16'd51365, 16'd51956, 16'd22311});
	test_expansion(128'ha6522b810d4249e35e7139b61089ad03, {16'd23739, 16'd46641, 16'd11721, 16'd36332, 16'd15991, 16'd12426, 16'd47549, 16'd41729, 16'd11766, 16'd38528, 16'd28500, 16'd58835, 16'd2296, 16'd6212, 16'd64839, 16'd4453, 16'd50059, 16'd64351, 16'd60923, 16'd61465, 16'd25562, 16'd56397, 16'd53257, 16'd45090, 16'd8411, 16'd23697});
	test_expansion(128'h1fe5bec7f662e411de6eff5a4f467b26, {16'd41731, 16'd2553, 16'd48659, 16'd65353, 16'd57211, 16'd9997, 16'd57847, 16'd53865, 16'd16600, 16'd14958, 16'd34130, 16'd40889, 16'd7048, 16'd10839, 16'd19063, 16'd58984, 16'd16814, 16'd7399, 16'd55386, 16'd53933, 16'd61877, 16'd49284, 16'd38887, 16'd30107, 16'd37885, 16'd23421});
	test_expansion(128'h6ca44be537d0d2d107e26b4b16c98232, {16'd5605, 16'd53038, 16'd58999, 16'd3008, 16'd2148, 16'd29202, 16'd9406, 16'd37652, 16'd21456, 16'd64125, 16'd53900, 16'd61782, 16'd59046, 16'd28117, 16'd43153, 16'd60232, 16'd59762, 16'd26602, 16'd36743, 16'd5417, 16'd6867, 16'd55678, 16'd54150, 16'd898, 16'd11584, 16'd47963});
	test_expansion(128'h0c5d1612d357e3c45217e6c756f00334, {16'd12789, 16'd15295, 16'd10816, 16'd57536, 16'd50662, 16'd58029, 16'd6946, 16'd47737, 16'd7690, 16'd42165, 16'd25005, 16'd43340, 16'd59824, 16'd17893, 16'd10445, 16'd59493, 16'd38302, 16'd7503, 16'd64501, 16'd30703, 16'd31595, 16'd28540, 16'd13189, 16'd52752, 16'd920, 16'd10618});
	test_expansion(128'h728e7ec134f57c4d61f582c5a35ef6e6, {16'd43900, 16'd19858, 16'd43906, 16'd26280, 16'd12352, 16'd24753, 16'd29062, 16'd6954, 16'd17699, 16'd45802, 16'd35422, 16'd45074, 16'd30588, 16'd61397, 16'd3749, 16'd32350, 16'd11894, 16'd56348, 16'd50281, 16'd20260, 16'd5488, 16'd45084, 16'd32708, 16'd51625, 16'd62177, 16'd45149});
	test_expansion(128'h8f535b733f7c6521b3aa57abe14d70dc, {16'd17108, 16'd57647, 16'd10739, 16'd30283, 16'd49794, 16'd41618, 16'd30697, 16'd8778, 16'd21113, 16'd57932, 16'd62932, 16'd46122, 16'd48167, 16'd35315, 16'd34390, 16'd17399, 16'd62200, 16'd2781, 16'd22836, 16'd25295, 16'd58728, 16'd168, 16'd61653, 16'd56268, 16'd25242, 16'd54231});
	test_expansion(128'h0843740e9e3177291a061c2ac9cb8bc0, {16'd54636, 16'd50077, 16'd38414, 16'd56271, 16'd47179, 16'd32825, 16'd54046, 16'd15105, 16'd62222, 16'd45690, 16'd63610, 16'd56193, 16'd9885, 16'd50891, 16'd23923, 16'd22628, 16'd64890, 16'd45470, 16'd63662, 16'd45280, 16'd9816, 16'd29051, 16'd56364, 16'd42910, 16'd48162, 16'd25834});
	test_expansion(128'h485443d322556bdd39e14d46768b9617, {16'd41501, 16'd59876, 16'd44952, 16'd1555, 16'd34376, 16'd43395, 16'd50975, 16'd15719, 16'd22434, 16'd21408, 16'd130, 16'd57617, 16'd11464, 16'd50191, 16'd33600, 16'd15099, 16'd25327, 16'd48171, 16'd54601, 16'd34648, 16'd18606, 16'd52111, 16'd21917, 16'd25656, 16'd23642, 16'd16544});
	test_expansion(128'h2754eb14a6c49367afbf55b616dd0414, {16'd8704, 16'd39584, 16'd17634, 16'd8286, 16'd31442, 16'd6263, 16'd34046, 16'd5497, 16'd2975, 16'd48413, 16'd19933, 16'd48005, 16'd52398, 16'd32422, 16'd10310, 16'd41832, 16'd48373, 16'd22161, 16'd4758, 16'd52892, 16'd18598, 16'd55946, 16'd27925, 16'd4245, 16'd50889, 16'd34958});
	test_expansion(128'hfb59934a64387c47b927586d5fd4e785, {16'd50585, 16'd24951, 16'd41815, 16'd65101, 16'd42895, 16'd4677, 16'd37667, 16'd61787, 16'd28030, 16'd34384, 16'd40764, 16'd45074, 16'd32057, 16'd63798, 16'd45774, 16'd23855, 16'd26440, 16'd29650, 16'd24954, 16'd44612, 16'd49752, 16'd63577, 16'd19694, 16'd12953, 16'd32608, 16'd37333});
	test_expansion(128'h610cbe903193692aa5988bacef0e6794, {16'd47379, 16'd61550, 16'd38527, 16'd23465, 16'd8288, 16'd5449, 16'd26530, 16'd51266, 16'd12011, 16'd29644, 16'd8233, 16'd14172, 16'd36719, 16'd59832, 16'd53329, 16'd4890, 16'd60374, 16'd46319, 16'd23674, 16'd59682, 16'd55102, 16'd31064, 16'd15244, 16'd7122, 16'd6250, 16'd688});
	test_expansion(128'h6179eb2f16c99890aaab4169a2ad034d, {16'd360, 16'd11189, 16'd27165, 16'd981, 16'd53471, 16'd31497, 16'd6750, 16'd34126, 16'd62457, 16'd49280, 16'd61686, 16'd5403, 16'd64054, 16'd47070, 16'd21879, 16'd10686, 16'd23208, 16'd25294, 16'd5166, 16'd28501, 16'd44753, 16'd59524, 16'd32383, 16'd54906, 16'd35258, 16'd60704});
	test_expansion(128'hb1d9a7339989cbc7b0c3c87f082de999, {16'd34674, 16'd2564, 16'd12757, 16'd59150, 16'd50503, 16'd24846, 16'd9620, 16'd34134, 16'd18177, 16'd24846, 16'd45924, 16'd19248, 16'd237, 16'd24273, 16'd10826, 16'd18734, 16'd54830, 16'd30649, 16'd11980, 16'd65147, 16'd17367, 16'd11330, 16'd33355, 16'd9666, 16'd25977, 16'd55113});
	test_expansion(128'h0624e341658a4e719ecd77e43642f7a8, {16'd39252, 16'd13425, 16'd33338, 16'd32206, 16'd16313, 16'd64318, 16'd2037, 16'd218, 16'd38064, 16'd24910, 16'd61330, 16'd53388, 16'd55928, 16'd34559, 16'd58922, 16'd49249, 16'd21778, 16'd41504, 16'd53982, 16'd30385, 16'd36593, 16'd25707, 16'd56832, 16'd52330, 16'd34978, 16'd27627});
	test_expansion(128'he448108020ecc4e1b449f7e288d725a6, {16'd30634, 16'd36684, 16'd23242, 16'd40975, 16'd50600, 16'd59650, 16'd12995, 16'd60497, 16'd39792, 16'd62650, 16'd38897, 16'd50401, 16'd28304, 16'd568, 16'd21066, 16'd9021, 16'd53273, 16'd7281, 16'd35038, 16'd41373, 16'd62256, 16'd41696, 16'd27893, 16'd14397, 16'd28159, 16'd64407});
	test_expansion(128'hddd99239a0313f0428dea9066bee8d91, {16'd51221, 16'd36826, 16'd14717, 16'd57276, 16'd53117, 16'd30661, 16'd25021, 16'd15928, 16'd8594, 16'd47320, 16'd1776, 16'd10750, 16'd57592, 16'd51586, 16'd47122, 16'd60437, 16'd44483, 16'd45793, 16'd48308, 16'd13307, 16'd61243, 16'd1621, 16'd17079, 16'd5571, 16'd47892, 16'd34252});
	test_expansion(128'h90bcb505b27b399d0fd7248b4d144eb7, {16'd51860, 16'd38585, 16'd53367, 16'd51113, 16'd33816, 16'd51174, 16'd65396, 16'd51309, 16'd50428, 16'd25900, 16'd2735, 16'd47437, 16'd20727, 16'd59757, 16'd41958, 16'd54793, 16'd16685, 16'd9424, 16'd51918, 16'd54685, 16'd58579, 16'd15001, 16'd12114, 16'd5609, 16'd58643, 16'd55609});
	test_expansion(128'hd5b7583ff31ed71c34ef24c469cd3dab, {16'd28120, 16'd41242, 16'd30452, 16'd65126, 16'd44542, 16'd14174, 16'd40701, 16'd4116, 16'd49514, 16'd12263, 16'd64207, 16'd46433, 16'd15298, 16'd8623, 16'd48282, 16'd1794, 16'd2061, 16'd24426, 16'd43636, 16'd46267, 16'd46327, 16'd27902, 16'd53824, 16'd22597, 16'd53670, 16'd21371});
	test_expansion(128'hbedf9cee5f9f901a9c827e5aa64b93b9, {16'd58900, 16'd60635, 16'd35273, 16'd19398, 16'd50249, 16'd58147, 16'd24686, 16'd21093, 16'd17108, 16'd60367, 16'd33491, 16'd45899, 16'd28430, 16'd56406, 16'd29651, 16'd8279, 16'd61880, 16'd16339, 16'd57112, 16'd54613, 16'd16564, 16'd57728, 16'd63390, 16'd57711, 16'd54730, 16'd5275});
	test_expansion(128'h11babb6c3c09495e2f586643ce89e589, {16'd38792, 16'd4119, 16'd42521, 16'd23271, 16'd17384, 16'd48135, 16'd52186, 16'd39128, 16'd55414, 16'd53076, 16'd31354, 16'd28093, 16'd55844, 16'd32867, 16'd36095, 16'd2095, 16'd42576, 16'd55950, 16'd22601, 16'd5587, 16'd55357, 16'd35366, 16'd35928, 16'd48205, 16'd8396, 16'd12845});
	test_expansion(128'h394a854fe00910f8843e461e381af465, {16'd3353, 16'd44359, 16'd7088, 16'd39430, 16'd6946, 16'd3239, 16'd54780, 16'd63136, 16'd8761, 16'd24709, 16'd50296, 16'd39832, 16'd57764, 16'd58049, 16'd41603, 16'd23320, 16'd6958, 16'd41732, 16'd56484, 16'd32007, 16'd64741, 16'd5154, 16'd63401, 16'd50504, 16'd55486, 16'd39535});
	test_expansion(128'h6ad2b372ba9a301042f591f0241cb786, {16'd35827, 16'd32265, 16'd790, 16'd24391, 16'd33370, 16'd61044, 16'd43542, 16'd11628, 16'd43787, 16'd45610, 16'd26768, 16'd30849, 16'd29309, 16'd3572, 16'd23208, 16'd60705, 16'd27250, 16'd30198, 16'd40745, 16'd11067, 16'd16262, 16'd1818, 16'd63058, 16'd3422, 16'd47962, 16'd11208});
	test_expansion(128'h451e9aa8b6f2f8070f6907f891164100, {16'd33466, 16'd55246, 16'd11541, 16'd31732, 16'd392, 16'd56010, 16'd61182, 16'd28615, 16'd58389, 16'd32879, 16'd64099, 16'd39245, 16'd190, 16'd9877, 16'd13449, 16'd18134, 16'd58447, 16'd25056, 16'd19489, 16'd65224, 16'd39097, 16'd14397, 16'd29967, 16'd17987, 16'd47188, 16'd21518});
	test_expansion(128'hbffd8f93544feefa1990bfc41e587d0d, {16'd31661, 16'd55602, 16'd15394, 16'd9351, 16'd10448, 16'd5231, 16'd23216, 16'd63376, 16'd48896, 16'd54834, 16'd58947, 16'd44816, 16'd60745, 16'd54596, 16'd61641, 16'd57312, 16'd23112, 16'd11098, 16'd47542, 16'd52109, 16'd32926, 16'd22922, 16'd60129, 16'd7932, 16'd5886, 16'd59520});
	test_expansion(128'hda3cc78df3c69e345baf6bd8fd3fbb20, {16'd4249, 16'd42647, 16'd27068, 16'd7381, 16'd5434, 16'd64168, 16'd6201, 16'd41145, 16'd4976, 16'd18652, 16'd11411, 16'd33822, 16'd30372, 16'd33498, 16'd43826, 16'd11245, 16'd51561, 16'd16087, 16'd63361, 16'd46982, 16'd17023, 16'd42481, 16'd12369, 16'd59124, 16'd15588, 16'd64977});
	test_expansion(128'h5bf470c744833a53103c2394f5822856, {16'd49714, 16'd1798, 16'd32355, 16'd29392, 16'd24279, 16'd65024, 16'd13105, 16'd37247, 16'd48608, 16'd62185, 16'd23639, 16'd19749, 16'd22929, 16'd47808, 16'd19513, 16'd41486, 16'd15510, 16'd26073, 16'd46176, 16'd41859, 16'd50036, 16'd43817, 16'd34516, 16'd6655, 16'd24730, 16'd9313});
	test_expansion(128'hd8a65ba7d3c36999ff18bdfbad99ab33, {16'd18851, 16'd12923, 16'd35306, 16'd18789, 16'd55798, 16'd43048, 16'd35957, 16'd42808, 16'd27992, 16'd38827, 16'd59143, 16'd1200, 16'd40467, 16'd49277, 16'd1490, 16'd63137, 16'd39598, 16'd8712, 16'd24405, 16'd30001, 16'd15624, 16'd12061, 16'd16305, 16'd14167, 16'd31090, 16'd23881});
	test_expansion(128'h7f8bdfad5714e56a136ed339ae4ab9e9, {16'd17285, 16'd7046, 16'd61425, 16'd15556, 16'd26352, 16'd43221, 16'd11935, 16'd48930, 16'd16992, 16'd51255, 16'd57556, 16'd26211, 16'd4228, 16'd51239, 16'd7972, 16'd56364, 16'd5511, 16'd60330, 16'd9075, 16'd49185, 16'd19876, 16'd53530, 16'd1920, 16'd59799, 16'd32332, 16'd34547});
	test_expansion(128'h07289cfe9b0a55add74e70d9a2265f28, {16'd22044, 16'd11092, 16'd64081, 16'd10956, 16'd29277, 16'd59324, 16'd26717, 16'd36874, 16'd37275, 16'd35544, 16'd52275, 16'd63094, 16'd24294, 16'd32198, 16'd55139, 16'd48226, 16'd180, 16'd3488, 16'd58168, 16'd33128, 16'd12979, 16'd9782, 16'd44237, 16'd20677, 16'd3499, 16'd27915});
	test_expansion(128'h2a9e6ece6aaa6a93753d616b43856973, {16'd53426, 16'd62035, 16'd25094, 16'd38166, 16'd14798, 16'd1541, 16'd13077, 16'd37336, 16'd2549, 16'd33881, 16'd25730, 16'd5145, 16'd11291, 16'd64149, 16'd47699, 16'd37349, 16'd43470, 16'd27940, 16'd25924, 16'd39399, 16'd29931, 16'd62023, 16'd42882, 16'd42431, 16'd12371, 16'd37374});
	test_expansion(128'hbdd00c3155d1ee2dc9cf6ff0785ce8aa, {16'd35561, 16'd3192, 16'd58870, 16'd31068, 16'd6854, 16'd63722, 16'd19895, 16'd44317, 16'd26424, 16'd55658, 16'd35176, 16'd59865, 16'd63282, 16'd2589, 16'd55134, 16'd53516, 16'd43265, 16'd698, 16'd47654, 16'd49545, 16'd47674, 16'd4738, 16'd10764, 16'd63526, 16'd25334, 16'd8394});
	test_expansion(128'h63f12509148c10a94cd02ae918b305c8, {16'd59555, 16'd828, 16'd48413, 16'd19293, 16'd29652, 16'd62074, 16'd49916, 16'd54311, 16'd63688, 16'd40589, 16'd50286, 16'd49387, 16'd47121, 16'd13191, 16'd38457, 16'd46307, 16'd49783, 16'd35759, 16'd13827, 16'd6725, 16'd55909, 16'd58545, 16'd39547, 16'd18494, 16'd25731, 16'd41803});
	test_expansion(128'h1e64a8d30fb26a30e9f11d6da64a601a, {16'd57513, 16'd35721, 16'd15067, 16'd63331, 16'd12126, 16'd47265, 16'd10008, 16'd35687, 16'd47614, 16'd46014, 16'd29488, 16'd31374, 16'd28012, 16'd26972, 16'd51346, 16'd59154, 16'd36218, 16'd13292, 16'd6968, 16'd35472, 16'd9980, 16'd33917, 16'd25809, 16'd25075, 16'd934, 16'd54386});
	test_expansion(128'h9402fc24ebd9f31ef15c45588eed18db, {16'd5847, 16'd47761, 16'd23867, 16'd45170, 16'd40766, 16'd49113, 16'd6303, 16'd59630, 16'd3909, 16'd23509, 16'd5278, 16'd23381, 16'd5750, 16'd44565, 16'd7466, 16'd63703, 16'd61547, 16'd55870, 16'd6303, 16'd64424, 16'd33616, 16'd7250, 16'd56733, 16'd9556, 16'd24589, 16'd28823});
	test_expansion(128'h1f5dee942fd4582b640a7c41072877ae, {16'd65315, 16'd34787, 16'd29812, 16'd52595, 16'd21589, 16'd29247, 16'd46587, 16'd28914, 16'd47098, 16'd48857, 16'd52688, 16'd48988, 16'd58695, 16'd8628, 16'd44231, 16'd55745, 16'd28956, 16'd47994, 16'd35166, 16'd64282, 16'd13827, 16'd32828, 16'd50815, 16'd37360, 16'd1937, 16'd20008});
	test_expansion(128'h598c898e58cc3efea5fb6526033bdea4, {16'd33389, 16'd29812, 16'd25506, 16'd33483, 16'd36694, 16'd7293, 16'd36268, 16'd58943, 16'd59407, 16'd29764, 16'd30995, 16'd36317, 16'd5128, 16'd43774, 16'd39112, 16'd57309, 16'd52522, 16'd15732, 16'd60017, 16'd59890, 16'd25489, 16'd45067, 16'd30898, 16'd63251, 16'd4673, 16'd2700});
	test_expansion(128'h4987f264b0f0289527745f953b7a5905, {16'd9701, 16'd55338, 16'd28914, 16'd62710, 16'd64689, 16'd8341, 16'd62470, 16'd2465, 16'd24124, 16'd21781, 16'd34956, 16'd60926, 16'd4266, 16'd25708, 16'd37406, 16'd51401, 16'd4024, 16'd54968, 16'd36030, 16'd11781, 16'd45046, 16'd10479, 16'd39771, 16'd12564, 16'd30810, 16'd59055});
	test_expansion(128'hc1c82dcb4004941bdea04305ffa49f35, {16'd24271, 16'd58496, 16'd30984, 16'd35267, 16'd57880, 16'd40027, 16'd12390, 16'd32681, 16'd29962, 16'd40156, 16'd14346, 16'd43009, 16'd52340, 16'd38366, 16'd2577, 16'd27900, 16'd40140, 16'd62707, 16'd54572, 16'd46369, 16'd24608, 16'd47603, 16'd4272, 16'd35106, 16'd50588, 16'd1506});
	test_expansion(128'hce9f3bca2e4e547fbbe67637e8440fea, {16'd47907, 16'd52313, 16'd13895, 16'd61732, 16'd2730, 16'd50048, 16'd65205, 16'd38363, 16'd25657, 16'd44604, 16'd24048, 16'd65347, 16'd2028, 16'd28938, 16'd56701, 16'd64535, 16'd52197, 16'd31800, 16'd55472, 16'd35706, 16'd46376, 16'd26480, 16'd46967, 16'd14231, 16'd44398, 16'd29039});
	test_expansion(128'h012915e46a7a26f6c771f53c3585573c, {16'd56197, 16'd39817, 16'd63086, 16'd35775, 16'd56316, 16'd48991, 16'd29315, 16'd20858, 16'd10004, 16'd36182, 16'd51649, 16'd19249, 16'd56896, 16'd1624, 16'd6979, 16'd40733, 16'd28236, 16'd59407, 16'd14019, 16'd19649, 16'd56022, 16'd53765, 16'd40117, 16'd2935, 16'd19709, 16'd57685});
	test_expansion(128'h502f66aa86f983ca4fdd6ac3f480925a, {16'd46050, 16'd62857, 16'd9534, 16'd22487, 16'd23003, 16'd26498, 16'd7762, 16'd3660, 16'd21808, 16'd15954, 16'd30700, 16'd31158, 16'd18314, 16'd52124, 16'd40453, 16'd48760, 16'd51939, 16'd21972, 16'd28188, 16'd44802, 16'd13847, 16'd34824, 16'd6013, 16'd63533, 16'd41076, 16'd28623});
	test_expansion(128'h521f24d7c9ebc04fad369169dbf1ec63, {16'd64829, 16'd55395, 16'd55114, 16'd57178, 16'd53176, 16'd42607, 16'd38390, 16'd53607, 16'd1662, 16'd41178, 16'd31586, 16'd33782, 16'd29399, 16'd9197, 16'd35023, 16'd15002, 16'd25522, 16'd63179, 16'd28133, 16'd64612, 16'd61810, 16'd46111, 16'd63824, 16'd16802, 16'd33778, 16'd4758});
	test_expansion(128'h1501a39d7349885efd0fff9beed82ee7, {16'd47214, 16'd392, 16'd63036, 16'd21203, 16'd59098, 16'd16896, 16'd39021, 16'd59558, 16'd13529, 16'd15178, 16'd13140, 16'd35038, 16'd49681, 16'd60189, 16'd16128, 16'd56596, 16'd30263, 16'd56991, 16'd31861, 16'd40550, 16'd19302, 16'd51531, 16'd2014, 16'd59828, 16'd49196, 16'd1407});
	test_expansion(128'h2ac589a4dd79c9d767d50b9bb220df43, {16'd44910, 16'd19404, 16'd34930, 16'd55161, 16'd23353, 16'd32053, 16'd21963, 16'd43742, 16'd24583, 16'd11572, 16'd64793, 16'd60432, 16'd54342, 16'd40376, 16'd52586, 16'd45353, 16'd4888, 16'd47459, 16'd4818, 16'd50214, 16'd45478, 16'd40843, 16'd31910, 16'd35979, 16'd46962, 16'd8773});
	test_expansion(128'h71c5d1d7a05a5e8bb06f8e6368a8ab14, {16'd20822, 16'd427, 16'd40581, 16'd17904, 16'd26804, 16'd40661, 16'd54087, 16'd13994, 16'd10394, 16'd20311, 16'd35337, 16'd7232, 16'd23597, 16'd41111, 16'd14228, 16'd17384, 16'd46111, 16'd5748, 16'd41210, 16'd2707, 16'd24339, 16'd4855, 16'd47236, 16'd47573, 16'd42097, 16'd32737});
	test_expansion(128'h2a707aef782b9b72449e53e9f12c8017, {16'd17422, 16'd63921, 16'd44978, 16'd937, 16'd59121, 16'd45101, 16'd55444, 16'd25558, 16'd24207, 16'd5166, 16'd25270, 16'd36113, 16'd36814, 16'd13704, 16'd3590, 16'd51358, 16'd15813, 16'd3183, 16'd49543, 16'd3612, 16'd35365, 16'd43361, 16'd8800, 16'd59558, 16'd2160, 16'd12451});
	test_expansion(128'h3fded8e82f03ac9e696ff6d7a3f69b4b, {16'd23674, 16'd27645, 16'd34800, 16'd47853, 16'd45318, 16'd60526, 16'd45781, 16'd6502, 16'd57609, 16'd46396, 16'd40431, 16'd12045, 16'd53224, 16'd9263, 16'd58784, 16'd45590, 16'd57414, 16'd64452, 16'd36736, 16'd15022, 16'd58935, 16'd15915, 16'd24260, 16'd1906, 16'd44487, 16'd4461});
	test_expansion(128'h6dd022d9afa808e5aff64153fb2af272, {16'd19900, 16'd27410, 16'd60813, 16'd24317, 16'd3614, 16'd55628, 16'd48618, 16'd53176, 16'd943, 16'd38701, 16'd31115, 16'd35603, 16'd45463, 16'd11118, 16'd19656, 16'd41785, 16'd40546, 16'd24595, 16'd22417, 16'd42794, 16'd12011, 16'd35534, 16'd7169, 16'd64495, 16'd12187, 16'd34599});
	test_expansion(128'hc6708b554ace46aa36fb30fd76e3c10a, {16'd53199, 16'd58763, 16'd11912, 16'd44131, 16'd20810, 16'd26346, 16'd39108, 16'd55511, 16'd32509, 16'd28657, 16'd7808, 16'd57560, 16'd45808, 16'd58629, 16'd36398, 16'd31925, 16'd44796, 16'd27913, 16'd25106, 16'd63415, 16'd38407, 16'd49865, 16'd27278, 16'd5884, 16'd7828, 16'd56521});
	test_expansion(128'h6de7129bedcf680ca7495e45ffbe1a5d, {16'd22573, 16'd26561, 16'd39685, 16'd43692, 16'd56838, 16'd15296, 16'd11006, 16'd34669, 16'd29172, 16'd64978, 16'd8707, 16'd24996, 16'd9434, 16'd21117, 16'd61221, 16'd2698, 16'd63585, 16'd1097, 16'd4246, 16'd656, 16'd63254, 16'd16723, 16'd9554, 16'd28366, 16'd30931, 16'd41859});
	test_expansion(128'heade3112243872c48abb2834efe09498, {16'd40484, 16'd18401, 16'd28381, 16'd42190, 16'd25775, 16'd58249, 16'd64162, 16'd32976, 16'd1522, 16'd37151, 16'd13814, 16'd65345, 16'd43973, 16'd10270, 16'd41270, 16'd61014, 16'd11422, 16'd11356, 16'd6858, 16'd63775, 16'd54263, 16'd11599, 16'd26159, 16'd50710, 16'd42144, 16'd28704});
	test_expansion(128'h03e85554fcaed9e11e2f9f2991c452b9, {16'd20791, 16'd22023, 16'd25000, 16'd57655, 16'd33303, 16'd15511, 16'd50667, 16'd25338, 16'd17267, 16'd10754, 16'd31595, 16'd7419, 16'd15474, 16'd17833, 16'd22918, 16'd41587, 16'd24612, 16'd61228, 16'd16293, 16'd37812, 16'd31763, 16'd17326, 16'd12439, 16'd33909, 16'd44596, 16'd45265});
	test_expansion(128'h4300197f4a34aed344d14800f9bd4498, {16'd11849, 16'd4181, 16'd15255, 16'd21278, 16'd30760, 16'd16229, 16'd24378, 16'd7463, 16'd10471, 16'd55741, 16'd47786, 16'd15519, 16'd22564, 16'd64084, 16'd41768, 16'd10455, 16'd8006, 16'd58025, 16'd31226, 16'd50633, 16'd23590, 16'd33289, 16'd22549, 16'd43520, 16'd3834, 16'd3388});
	test_expansion(128'h627a90b5ab138860a13546f503d8b00a, {16'd13838, 16'd63896, 16'd39229, 16'd40240, 16'd32346, 16'd63432, 16'd41581, 16'd48748, 16'd62934, 16'd16365, 16'd22328, 16'd50008, 16'd37010, 16'd21923, 16'd40942, 16'd9332, 16'd27307, 16'd31644, 16'd5715, 16'd12192, 16'd38739, 16'd64085, 16'd26627, 16'd18789, 16'd52230, 16'd39367});
	test_expansion(128'hdcd813aa603506386363902b4aa41226, {16'd20808, 16'd20218, 16'd42311, 16'd49728, 16'd463, 16'd24858, 16'd4074, 16'd37374, 16'd62153, 16'd7298, 16'd19579, 16'd28437, 16'd29899, 16'd11566, 16'd38937, 16'd54329, 16'd59406, 16'd41230, 16'd14474, 16'd7616, 16'd64542, 16'd24665, 16'd21776, 16'd37455, 16'd61041, 16'd18530});
	test_expansion(128'h22a81a3573b9e56637f37ee7efdcee62, {16'd20982, 16'd45567, 16'd20570, 16'd46875, 16'd24660, 16'd31728, 16'd17330, 16'd20730, 16'd24286, 16'd45649, 16'd31733, 16'd29213, 16'd49565, 16'd49906, 16'd56864, 16'd12818, 16'd29462, 16'd19675, 16'd41126, 16'd52534, 16'd7436, 16'd730, 16'd9778, 16'd56572, 16'd55375, 16'd6973});
	test_expansion(128'h29f82a04193bf111ab9eb576c9f4e1a0, {16'd50141, 16'd50628, 16'd15460, 16'd34674, 16'd65021, 16'd63214, 16'd6573, 16'd8584, 16'd27941, 16'd56170, 16'd52781, 16'd44067, 16'd25668, 16'd56769, 16'd56388, 16'd21569, 16'd61127, 16'd7571, 16'd44790, 16'd26059, 16'd12566, 16'd59139, 16'd26242, 16'd9104, 16'd29154, 16'd35122});
	test_expansion(128'h18e6a94ae46b0999c013bef89dd083aa, {16'd43233, 16'd10892, 16'd59575, 16'd5256, 16'd5883, 16'd45795, 16'd9776, 16'd23881, 16'd47079, 16'd18860, 16'd6692, 16'd55703, 16'd56107, 16'd25201, 16'd3106, 16'd16906, 16'd42962, 16'd41333, 16'd16984, 16'd947, 16'd2899, 16'd40038, 16'd1969, 16'd17433, 16'd51792, 16'd18750});
	test_expansion(128'h20c6e9ddaa42d36b6c871e35a3908a23, {16'd49554, 16'd9838, 16'd8929, 16'd34847, 16'd11861, 16'd48657, 16'd20927, 16'd5848, 16'd864, 16'd45734, 16'd44369, 16'd45630, 16'd11244, 16'd46975, 16'd34065, 16'd416, 16'd26809, 16'd31466, 16'd51821, 16'd14354, 16'd5188, 16'd54397, 16'd62232, 16'd11391, 16'd26863, 16'd13085});
	test_expansion(128'h0b413974e634841b3039a299383a9dfe, {16'd59297, 16'd50388, 16'd45603, 16'd8078, 16'd27902, 16'd61811, 16'd45050, 16'd1134, 16'd47022, 16'd43115, 16'd12272, 16'd44252, 16'd10975, 16'd12192, 16'd37808, 16'd61925, 16'd23547, 16'd51211, 16'd19453, 16'd40334, 16'd53016, 16'd14662, 16'd22245, 16'd23878, 16'd54235, 16'd59272});
	test_expansion(128'h4610a98513fe2904c54122737069f75a, {16'd64218, 16'd32062, 16'd24430, 16'd51681, 16'd24573, 16'd6010, 16'd10823, 16'd25399, 16'd32612, 16'd18132, 16'd58731, 16'd24968, 16'd20280, 16'd6565, 16'd22759, 16'd7895, 16'd8695, 16'd38990, 16'd6022, 16'd54574, 16'd11992, 16'd25845, 16'd47222, 16'd3365, 16'd18342, 16'd56421});
	test_expansion(128'h306900281932d1b6bf385353958c026e, {16'd62733, 16'd52455, 16'd22345, 16'd38704, 16'd15981, 16'd3805, 16'd57426, 16'd8229, 16'd2678, 16'd57760, 16'd20388, 16'd4306, 16'd43801, 16'd22786, 16'd49460, 16'd60544, 16'd21785, 16'd43633, 16'd15112, 16'd15822, 16'd45368, 16'd63009, 16'd59367, 16'd7147, 16'd63770, 16'd61075});
	test_expansion(128'h796a104adf1b92123d7b37f1d224127d, {16'd17318, 16'd14763, 16'd23893, 16'd58422, 16'd5285, 16'd13996, 16'd60267, 16'd31161, 16'd16747, 16'd29405, 16'd61226, 16'd16669, 16'd36708, 16'd36199, 16'd53845, 16'd49851, 16'd57844, 16'd19152, 16'd51754, 16'd28623, 16'd11587, 16'd11311, 16'd6457, 16'd5880, 16'd20805, 16'd54818});
	test_expansion(128'h9c83ca8a905b1270926da3e6527e352a, {16'd14407, 16'd5518, 16'd57891, 16'd25232, 16'd40425, 16'd20709, 16'd58384, 16'd26185, 16'd55274, 16'd33605, 16'd43045, 16'd63538, 16'd24690, 16'd12475, 16'd59987, 16'd3421, 16'd8083, 16'd37506, 16'd27126, 16'd63328, 16'd29070, 16'd62653, 16'd34380, 16'd16150, 16'd3885, 16'd54604});
	test_expansion(128'h9164fd3c3bb88fda0df3c16e1c5f8959, {16'd55543, 16'd38537, 16'd3334, 16'd49511, 16'd32829, 16'd44471, 16'd2502, 16'd59530, 16'd27185, 16'd30663, 16'd43179, 16'd3306, 16'd17738, 16'd53622, 16'd40692, 16'd24566, 16'd65181, 16'd31560, 16'd29628, 16'd24214, 16'd58504, 16'd32071, 16'd61102, 16'd24986, 16'd9852, 16'd45780});
	test_expansion(128'h1b3a100c5c2706e5af3a7a1125bfce24, {16'd51180, 16'd64946, 16'd45162, 16'd53431, 16'd14916, 16'd57451, 16'd10770, 16'd20545, 16'd27709, 16'd37857, 16'd56340, 16'd8009, 16'd59345, 16'd5013, 16'd20037, 16'd55086, 16'd28136, 16'd61905, 16'd22266, 16'd50709, 16'd27146, 16'd61388, 16'd34310, 16'd16408, 16'd51783, 16'd63994});
	test_expansion(128'h64932764d515fa703eb2a0b0d5c91407, {16'd33567, 16'd25259, 16'd57723, 16'd38230, 16'd5803, 16'd63950, 16'd37454, 16'd13792, 16'd3639, 16'd4952, 16'd16207, 16'd31370, 16'd37553, 16'd47216, 16'd34382, 16'd59682, 16'd40505, 16'd49104, 16'd57684, 16'd1026, 16'd64591, 16'd64353, 16'd60316, 16'd8795, 16'd9947, 16'd17436});
	test_expansion(128'h33f0cd49dfea855109b8ba5507b95dee, {16'd57188, 16'd36249, 16'd10910, 16'd9663, 16'd59075, 16'd7852, 16'd6987, 16'd15376, 16'd15070, 16'd20915, 16'd38503, 16'd11603, 16'd48632, 16'd22385, 16'd39157, 16'd58669, 16'd5444, 16'd44250, 16'd10910, 16'd4912, 16'd10262, 16'd7571, 16'd47605, 16'd35538, 16'd33512, 16'd60362});
	test_expansion(128'hc55c3dbc147a82edbc4e5d17b1ddb172, {16'd60382, 16'd61863, 16'd52223, 16'd21736, 16'd23050, 16'd47928, 16'd40134, 16'd15371, 16'd56199, 16'd45810, 16'd55362, 16'd24945, 16'd10726, 16'd31561, 16'd6093, 16'd27702, 16'd4955, 16'd13796, 16'd26001, 16'd44763, 16'd3594, 16'd26436, 16'd16803, 16'd50957, 16'd30097, 16'd19525});
	test_expansion(128'h651deeb9a200b70ec069f3c164be284b, {16'd26336, 16'd21724, 16'd21633, 16'd20937, 16'd4113, 16'd1085, 16'd24587, 16'd45921, 16'd61579, 16'd64112, 16'd26157, 16'd23435, 16'd47920, 16'd21906, 16'd31430, 16'd48504, 16'd25914, 16'd6252, 16'd9410, 16'd63065, 16'd18386, 16'd20657, 16'd32004, 16'd47506, 16'd15604, 16'd44806});
	test_expansion(128'hf9bfeff026f903439e6d48ce0c42aded, {16'd7036, 16'd55789, 16'd38885, 16'd44273, 16'd45379, 16'd58169, 16'd56542, 16'd44136, 16'd50232, 16'd57968, 16'd46088, 16'd18997, 16'd3108, 16'd24859, 16'd11528, 16'd53765, 16'd45822, 16'd29849, 16'd55543, 16'd28322, 16'd60377, 16'd14561, 16'd36440, 16'd56413, 16'd22003, 16'd9373});
	test_expansion(128'h00cf7fccb3e73d6d572d161845bed431, {16'd22771, 16'd24011, 16'd3929, 16'd64797, 16'd17809, 16'd9708, 16'd44877, 16'd62627, 16'd52622, 16'd59760, 16'd15981, 16'd61990, 16'd58871, 16'd54507, 16'd41967, 16'd18658, 16'd57583, 16'd47402, 16'd38803, 16'd15739, 16'd8116, 16'd41886, 16'd8317, 16'd55690, 16'd46683, 16'd12821});
	test_expansion(128'hff4be854aca2ca42fba6099ab6d8d112, {16'd43696, 16'd34745, 16'd26949, 16'd23951, 16'd24893, 16'd18573, 16'd16324, 16'd52137, 16'd48099, 16'd56747, 16'd65394, 16'd56502, 16'd4232, 16'd832, 16'd24869, 16'd60428, 16'd4104, 16'd23911, 16'd47426, 16'd15349, 16'd58218, 16'd9528, 16'd59170, 16'd6614, 16'd15340, 16'd36260});
	test_expansion(128'h751b0c7335685a91275497527afa1db7, {16'd20706, 16'd55598, 16'd6727, 16'd60460, 16'd28085, 16'd14090, 16'd34495, 16'd2366, 16'd42065, 16'd57388, 16'd41919, 16'd42541, 16'd35060, 16'd17901, 16'd60424, 16'd51260, 16'd41990, 16'd26594, 16'd54202, 16'd23992, 16'd2308, 16'd30845, 16'd7, 16'd16465, 16'd12625, 16'd2044});
	test_expansion(128'h8edd3690cf5aa23936209268db4cfb44, {16'd4230, 16'd10904, 16'd43295, 16'd19353, 16'd49789, 16'd64831, 16'd44643, 16'd23256, 16'd18512, 16'd20496, 16'd39864, 16'd51373, 16'd53073, 16'd35105, 16'd41368, 16'd22971, 16'd29039, 16'd63072, 16'd9172, 16'd13038, 16'd21620, 16'd28049, 16'd38118, 16'd52232, 16'd18568, 16'd49107});
	test_expansion(128'ha3b27f39f93154995e3751f9f048356e, {16'd43515, 16'd2389, 16'd24797, 16'd59287, 16'd58136, 16'd7011, 16'd24911, 16'd23782, 16'd25288, 16'd64529, 16'd22115, 16'd60930, 16'd48830, 16'd60325, 16'd43186, 16'd23755, 16'd25217, 16'd50748, 16'd45844, 16'd25796, 16'd46139, 16'd5536, 16'd7396, 16'd46102, 16'd25230, 16'd11474});
	test_expansion(128'hcdfbca420fca1e62d3b327261a22cc5c, {16'd21796, 16'd29626, 16'd7591, 16'd58132, 16'd51498, 16'd1957, 16'd37378, 16'd55885, 16'd19093, 16'd50810, 16'd38668, 16'd20229, 16'd36392, 16'd17541, 16'd46936, 16'd63332, 16'd52741, 16'd461, 16'd44461, 16'd4317, 16'd44760, 16'd41339, 16'd2195, 16'd30257, 16'd14929, 16'd56012});
	test_expansion(128'h17034f555e3a21d8f2792cbfe932f67a, {16'd14181, 16'd63238, 16'd24248, 16'd54478, 16'd2250, 16'd37627, 16'd52794, 16'd58219, 16'd53366, 16'd27645, 16'd57702, 16'd60355, 16'd10079, 16'd52531, 16'd39617, 16'd31614, 16'd28318, 16'd12660, 16'd23015, 16'd45315, 16'd11767, 16'd26339, 16'd49448, 16'd4284, 16'd2814, 16'd23786});
	test_expansion(128'h8146b0144314e64934d18977c7bce9c0, {16'd30114, 16'd25850, 16'd4841, 16'd50804, 16'd21623, 16'd41755, 16'd2013, 16'd34910, 16'd6091, 16'd38730, 16'd46031, 16'd61219, 16'd57067, 16'd1021, 16'd21147, 16'd39969, 16'd11015, 16'd7989, 16'd14419, 16'd37382, 16'd30723, 16'd30315, 16'd18821, 16'd19296, 16'd20471, 16'd36343});
	test_expansion(128'hb8fc37199283d3967b0612ebbfb430af, {16'd35682, 16'd35317, 16'd50049, 16'd50975, 16'd47083, 16'd38403, 16'd14466, 16'd62343, 16'd1388, 16'd40459, 16'd27281, 16'd48167, 16'd62750, 16'd37301, 16'd39322, 16'd40756, 16'd44568, 16'd52187, 16'd18814, 16'd45362, 16'd63074, 16'd35913, 16'd9372, 16'd25264, 16'd16654, 16'd62309});
	test_expansion(128'h42c32c7855383c3879560c5bef605e0d, {16'd7858, 16'd36001, 16'd45727, 16'd23244, 16'd46555, 16'd21265, 16'd1864, 16'd41425, 16'd4273, 16'd4883, 16'd55387, 16'd60736, 16'd24993, 16'd52407, 16'd5429, 16'd9946, 16'd7749, 16'd61801, 16'd30504, 16'd23361, 16'd21948, 16'd2622, 16'd10729, 16'd6986, 16'd44025, 16'd59976});
	test_expansion(128'h48cb578fd3c97e908984131314f98180, {16'd25641, 16'd38792, 16'd63489, 16'd11625, 16'd64093, 16'd64831, 16'd24156, 16'd27332, 16'd10085, 16'd51329, 16'd57719, 16'd55573, 16'd64058, 16'd49257, 16'd60084, 16'd26985, 16'd37170, 16'd48845, 16'd58818, 16'd55767, 16'd47411, 16'd7897, 16'd15440, 16'd37407, 16'd50372, 16'd24152});
	test_expansion(128'h1e6ccb7db4e07a2b30066a27df2b8ed8, {16'd2614, 16'd58891, 16'd25365, 16'd55313, 16'd59697, 16'd12700, 16'd52528, 16'd20996, 16'd11915, 16'd10134, 16'd57560, 16'd60329, 16'd37966, 16'd35068, 16'd841, 16'd17197, 16'd7070, 16'd49842, 16'd19643, 16'd39091, 16'd3865, 16'd25823, 16'd27646, 16'd57204, 16'd12253, 16'd60751});
	test_expansion(128'he113e5bc220169288756ab0dc355fa4e, {16'd60693, 16'd46896, 16'd50054, 16'd35004, 16'd46110, 16'd41100, 16'd50647, 16'd39139, 16'd49872, 16'd23191, 16'd18737, 16'd6245, 16'd3703, 16'd37703, 16'd52986, 16'd48773, 16'd56736, 16'd50289, 16'd33586, 16'd39620, 16'd63175, 16'd31911, 16'd20996, 16'd18341, 16'd22787, 16'd43989});
	test_expansion(128'hebc47c36d66860bbca714bf031e5f64e, {16'd3486, 16'd63720, 16'd53628, 16'd64677, 16'd45465, 16'd59308, 16'd11822, 16'd16037, 16'd22429, 16'd51050, 16'd11066, 16'd30280, 16'd53321, 16'd65203, 16'd65009, 16'd48746, 16'd10289, 16'd12183, 16'd21119, 16'd56433, 16'd31111, 16'd61558, 16'd23605, 16'd5539, 16'd56175, 16'd56446});
	test_expansion(128'hbbc9c66096cfb611216418b5178567f9, {16'd61107, 16'd59829, 16'd6395, 16'd21701, 16'd608, 16'd19397, 16'd47473, 16'd61797, 16'd6723, 16'd47630, 16'd23118, 16'd33865, 16'd43760, 16'd51968, 16'd37800, 16'd41771, 16'd36718, 16'd5492, 16'd45233, 16'd31048, 16'd40393, 16'd18447, 16'd15022, 16'd8819, 16'd23890, 16'd34004});
	test_expansion(128'h9314d8161fb041072fa1ec51f8c7a8de, {16'd2810, 16'd45409, 16'd62014, 16'd48288, 16'd38610, 16'd13138, 16'd44633, 16'd28103, 16'd5562, 16'd42366, 16'd64478, 16'd32546, 16'd6134, 16'd14377, 16'd54679, 16'd13760, 16'd18681, 16'd47520, 16'd21430, 16'd14064, 16'd12214, 16'd61945, 16'd25642, 16'd51361, 16'd44151, 16'd41175});
	test_expansion(128'h62bcf9ffda7cf43f416d335bec7611f4, {16'd42581, 16'd53401, 16'd16914, 16'd55827, 16'd38095, 16'd48907, 16'd52320, 16'd40643, 16'd43345, 16'd40570, 16'd41666, 16'd15049, 16'd10746, 16'd13509, 16'd18883, 16'd15673, 16'd32624, 16'd33509, 16'd38340, 16'd62588, 16'd14632, 16'd45630, 16'd45481, 16'd35677, 16'd40514, 16'd52010});
	test_expansion(128'hc35fd1df4a7ce9779bae437c26fb8997, {16'd50470, 16'd31495, 16'd48323, 16'd4554, 16'd32427, 16'd60610, 16'd19293, 16'd33511, 16'd8473, 16'd13881, 16'd6570, 16'd28405, 16'd1752, 16'd4954, 16'd23685, 16'd45441, 16'd53103, 16'd29560, 16'd25420, 16'd45116, 16'd52742, 16'd40491, 16'd37915, 16'd58969, 16'd41148, 16'd29033});
	test_expansion(128'h2648f0ce1b03111de9e823ac2ee6aa07, {16'd28148, 16'd3923, 16'd32587, 16'd8209, 16'd24182, 16'd64185, 16'd45401, 16'd58538, 16'd54833, 16'd35289, 16'd65043, 16'd23897, 16'd630, 16'd4480, 16'd43505, 16'd64425, 16'd63924, 16'd19618, 16'd51801, 16'd64239, 16'd44529, 16'd9155, 16'd2141, 16'd40360, 16'd31797, 16'd12994});
	test_expansion(128'ha8c18af6752fb1ff8398f34e61696498, {16'd4679, 16'd47924, 16'd56010, 16'd56374, 16'd64943, 16'd40458, 16'd16667, 16'd65084, 16'd17512, 16'd11209, 16'd39417, 16'd25103, 16'd5434, 16'd29276, 16'd58107, 16'd2169, 16'd47614, 16'd24417, 16'd45578, 16'd4913, 16'd27145, 16'd43929, 16'd46197, 16'd19269, 16'd35093, 16'd14054});
	test_expansion(128'he8d5f1de0e1eda1e4281774d9362bdf0, {16'd14687, 16'd25396, 16'd12851, 16'd29136, 16'd33471, 16'd29828, 16'd33242, 16'd48244, 16'd13304, 16'd2828, 16'd44835, 16'd61663, 16'd23796, 16'd11875, 16'd33132, 16'd12893, 16'd9202, 16'd45894, 16'd64797, 16'd30212, 16'd11508, 16'd8379, 16'd40575, 16'd27482, 16'd48313, 16'd56039});
	test_expansion(128'h6bad4e4ba45dd7cac5a3aa9f53f8221d, {16'd15280, 16'd30687, 16'd4963, 16'd40279, 16'd19558, 16'd3582, 16'd9841, 16'd8376, 16'd6071, 16'd28308, 16'd52844, 16'd60386, 16'd53672, 16'd60681, 16'd42358, 16'd54813, 16'd4640, 16'd62974, 16'd63273, 16'd5060, 16'd63971, 16'd27147, 16'd35689, 16'd14539, 16'd49287, 16'd27460});
	test_expansion(128'h009853ffe3b180c46b0abc857fdbba4f, {16'd50638, 16'd4922, 16'd48404, 16'd58419, 16'd53554, 16'd20077, 16'd32537, 16'd41150, 16'd34743, 16'd37975, 16'd24829, 16'd54738, 16'd41568, 16'd20472, 16'd45265, 16'd60657, 16'd64837, 16'd53281, 16'd63579, 16'd16263, 16'd34566, 16'd57103, 16'd21000, 16'd36021, 16'd1243, 16'd25622});
	test_expansion(128'hb9c76b17031fe5347c8f04e3023fb4b1, {16'd13269, 16'd63039, 16'd4968, 16'd9301, 16'd40268, 16'd53020, 16'd32991, 16'd57762, 16'd43565, 16'd31090, 16'd33202, 16'd13611, 16'd38160, 16'd26414, 16'd51183, 16'd48364, 16'd32536, 16'd41654, 16'd62407, 16'd57971, 16'd38035, 16'd16809, 16'd6603, 16'd60674, 16'd7519, 16'd14355});
	test_expansion(128'hb6650564028025d2f6065f5c49960a36, {16'd5506, 16'd7896, 16'd47849, 16'd55533, 16'd32174, 16'd8387, 16'd1075, 16'd18172, 16'd36112, 16'd62441, 16'd51271, 16'd43509, 16'd11143, 16'd51048, 16'd62730, 16'd50913, 16'd36276, 16'd2121, 16'd51249, 16'd39723, 16'd29065, 16'd45627, 16'd10076, 16'd51774, 16'd18712, 16'd2902});
	test_expansion(128'ha30b713b2145815c54e00f15105522df, {16'd47784, 16'd44769, 16'd14453, 16'd55620, 16'd63774, 16'd34392, 16'd27667, 16'd747, 16'd28840, 16'd31014, 16'd51184, 16'd40082, 16'd4961, 16'd6380, 16'd8107, 16'd20846, 16'd33044, 16'd3266, 16'd27032, 16'd51585, 16'd63541, 16'd37173, 16'd43842, 16'd10720, 16'd1554, 16'd40530});
	test_expansion(128'h4d51da176c7a7e1d888fa6020b6537c7, {16'd49177, 16'd25723, 16'd16485, 16'd31559, 16'd12453, 16'd44438, 16'd37416, 16'd17880, 16'd16370, 16'd25947, 16'd11688, 16'd22560, 16'd43045, 16'd24504, 16'd55638, 16'd4785, 16'd16691, 16'd61489, 16'd63497, 16'd6044, 16'd55153, 16'd30532, 16'd3347, 16'd2808, 16'd8199, 16'd36734});
	test_expansion(128'h2b88ada416c2ab52289f68d324e13d67, {16'd44977, 16'd35391, 16'd52222, 16'd133, 16'd33547, 16'd55960, 16'd58370, 16'd41478, 16'd26403, 16'd24626, 16'd33831, 16'd25014, 16'd2950, 16'd42871, 16'd34005, 16'd4276, 16'd11676, 16'd50359, 16'd17644, 16'd28179, 16'd21808, 16'd52403, 16'd47973, 16'd33957, 16'd12300, 16'd62985});
	test_expansion(128'h1c4bbaf67e00c33e56a84e2c005e0fe7, {16'd39745, 16'd58043, 16'd41650, 16'd54092, 16'd1255, 16'd14249, 16'd13728, 16'd17354, 16'd45489, 16'd26301, 16'd62844, 16'd11982, 16'd42658, 16'd44521, 16'd46401, 16'd20997, 16'd8258, 16'd33516, 16'd9406, 16'd62809, 16'd29633, 16'd45354, 16'd63485, 16'd44329, 16'd59168, 16'd61906});
	test_expansion(128'hcdca3ce837e52e28009a4e42c5e34c2d, {16'd35359, 16'd33268, 16'd41103, 16'd33030, 16'd34221, 16'd10160, 16'd18042, 16'd21805, 16'd36922, 16'd62845, 16'd5070, 16'd60564, 16'd13327, 16'd29729, 16'd26238, 16'd42539, 16'd281, 16'd16861, 16'd11470, 16'd43512, 16'd2302, 16'd26055, 16'd45573, 16'd2028, 16'd38932, 16'd21409});
	test_expansion(128'ha37a351e91d84a2843dc69f2045f5752, {16'd53195, 16'd54821, 16'd52244, 16'd23484, 16'd28888, 16'd50281, 16'd34190, 16'd44880, 16'd25862, 16'd13651, 16'd15420, 16'd42992, 16'd45178, 16'd30540, 16'd6038, 16'd26616, 16'd33909, 16'd49597, 16'd15738, 16'd55767, 16'd6132, 16'd55913, 16'd57007, 16'd16877, 16'd29990, 16'd27857});
	test_expansion(128'h874d7f35e8a08d829fb74930b87ccec7, {16'd28986, 16'd34448, 16'd35335, 16'd12960, 16'd10833, 16'd57797, 16'd2099, 16'd14044, 16'd60530, 16'd51812, 16'd30809, 16'd47635, 16'd14064, 16'd23205, 16'd52970, 16'd38801, 16'd53434, 16'd54246, 16'd46008, 16'd56821, 16'd43438, 16'd25254, 16'd25579, 16'd13782, 16'd54153, 16'd10271});
	test_expansion(128'hae267a10ab133f91f47366716be4e148, {16'd279, 16'd55222, 16'd2773, 16'd4362, 16'd57405, 16'd63151, 16'd22388, 16'd31246, 16'd15833, 16'd3213, 16'd42174, 16'd22603, 16'd21596, 16'd6234, 16'd4561, 16'd22989, 16'd44518, 16'd33930, 16'd5394, 16'd39686, 16'd26706, 16'd49008, 16'd18765, 16'd18899, 16'd50174, 16'd58617});
	test_expansion(128'hf12af2064827ca74603d506910a315df, {16'd24380, 16'd4615, 16'd31987, 16'd23913, 16'd25055, 16'd33489, 16'd15909, 16'd54113, 16'd35629, 16'd12879, 16'd29805, 16'd18995, 16'd59574, 16'd27990, 16'd49610, 16'd47331, 16'd55814, 16'd46804, 16'd11481, 16'd36048, 16'd32177, 16'd25644, 16'd51651, 16'd323, 16'd44601, 16'd61590});
	test_expansion(128'h49ebe1f854d26d0001105254cf7f470b, {16'd41635, 16'd7742, 16'd21851, 16'd55984, 16'd15743, 16'd39191, 16'd50615, 16'd19832, 16'd30302, 16'd23244, 16'd53773, 16'd25078, 16'd34445, 16'd20055, 16'd48659, 16'd31799, 16'd4734, 16'd2777, 16'd19509, 16'd5367, 16'd62116, 16'd337, 16'd5025, 16'd9016, 16'd46770, 16'd51857});
	test_expansion(128'h15952d6883adebb57b5c5d8db289fcfe, {16'd12413, 16'd36546, 16'd62341, 16'd29000, 16'd19805, 16'd21693, 16'd9443, 16'd34930, 16'd54372, 16'd64879, 16'd16866, 16'd26044, 16'd47282, 16'd40028, 16'd33053, 16'd42468, 16'd12561, 16'd3377, 16'd3576, 16'd46103, 16'd50647, 16'd38077, 16'd25468, 16'd57248, 16'd20394, 16'd35146});
	test_expansion(128'h9786a608b29ffbeec66824f96c7a3bbf, {16'd24427, 16'd25630, 16'd34886, 16'd42659, 16'd17153, 16'd44472, 16'd42172, 16'd50110, 16'd39890, 16'd56452, 16'd29841, 16'd50945, 16'd647, 16'd64103, 16'd64286, 16'd13694, 16'd49032, 16'd57171, 16'd42274, 16'd43811, 16'd59284, 16'd11262, 16'd58056, 16'd40577, 16'd58761, 16'd11060});
	test_expansion(128'h4bdd52a76dc8f1151ffbc807a6347eab, {16'd53876, 16'd27599, 16'd62505, 16'd7201, 16'd39454, 16'd15486, 16'd40132, 16'd45592, 16'd22984, 16'd17561, 16'd27071, 16'd61721, 16'd7789, 16'd45533, 16'd31859, 16'd63300, 16'd63700, 16'd39528, 16'd28403, 16'd35574, 16'd56157, 16'd19259, 16'd61180, 16'd46415, 16'd57204, 16'd2682});
	test_expansion(128'hf65228f3466994672bf80d358a76878d, {16'd625, 16'd4093, 16'd25288, 16'd39842, 16'd25135, 16'd3278, 16'd59692, 16'd13799, 16'd28144, 16'd26942, 16'd47985, 16'd10537, 16'd64889, 16'd36438, 16'd47577, 16'd35869, 16'd20785, 16'd52426, 16'd23046, 16'd61958, 16'd16223, 16'd24045, 16'd1619, 16'd23804, 16'd44728, 16'd51492});
	test_expansion(128'h7dd892bb48d805652109850ab680dee0, {16'd23466, 16'd62024, 16'd18825, 16'd43861, 16'd64725, 16'd37681, 16'd25496, 16'd32847, 16'd11656, 16'd30036, 16'd49105, 16'd18545, 16'd14217, 16'd16210, 16'd23126, 16'd26543, 16'd63930, 16'd19942, 16'd14449, 16'd31914, 16'd29967, 16'd23566, 16'd31123, 16'd58146, 16'd44763, 16'd50600});
	test_expansion(128'h82cb31197562862e5ca12fadf7b3cd35, {16'd48224, 16'd8102, 16'd53093, 16'd13466, 16'd7053, 16'd29168, 16'd56683, 16'd7221, 16'd45147, 16'd11467, 16'd50167, 16'd18011, 16'd29341, 16'd51342, 16'd24081, 16'd4241, 16'd38883, 16'd5599, 16'd15435, 16'd1811, 16'd36557, 16'd26210, 16'd63920, 16'd22866, 16'd775, 16'd30599});
	test_expansion(128'h1c4d11eb3f2893731ac1e108fc95d640, {16'd52952, 16'd49600, 16'd9163, 16'd11346, 16'd57038, 16'd10410, 16'd24590, 16'd20509, 16'd40051, 16'd40716, 16'd36592, 16'd57233, 16'd55432, 16'd53768, 16'd17907, 16'd9037, 16'd45351, 16'd56169, 16'd63272, 16'd50746, 16'd25000, 16'd342, 16'd62032, 16'd7970, 16'd3067, 16'd60484});
	test_expansion(128'hb710bc617928c713586e7e356eb57d7a, {16'd2481, 16'd9964, 16'd62489, 16'd1581, 16'd19590, 16'd61189, 16'd19157, 16'd54506, 16'd6078, 16'd34983, 16'd43803, 16'd37338, 16'd30416, 16'd37933, 16'd28904, 16'd41491, 16'd10344, 16'd38991, 16'd34043, 16'd26171, 16'd186, 16'd59391, 16'd2964, 16'd52945, 16'd3694, 16'd46968});
	test_expansion(128'hf3dc37203365317bd8708c03ee472012, {16'd10375, 16'd27820, 16'd8822, 16'd56016, 16'd18539, 16'd60931, 16'd50811, 16'd29762, 16'd61461, 16'd46787, 16'd34964, 16'd48566, 16'd34307, 16'd52269, 16'd25512, 16'd54099, 16'd21593, 16'd51121, 16'd33969, 16'd24863, 16'd53022, 16'd29980, 16'd4316, 16'd9242, 16'd44661, 16'd5963});
	test_expansion(128'h760a36236c03c91dad064871943df315, {16'd17544, 16'd41336, 16'd35231, 16'd29781, 16'd19628, 16'd31903, 16'd2948, 16'd51620, 16'd63702, 16'd55110, 16'd6046, 16'd55301, 16'd31618, 16'd21268, 16'd1856, 16'd31960, 16'd3588, 16'd57841, 16'd59577, 16'd53072, 16'd50241, 16'd18851, 16'd63711, 16'd43771, 16'd14300, 16'd30456});
	test_expansion(128'h6fa5f60e10dba43c7e99aeb5d391bdb9, {16'd38841, 16'd13869, 16'd44194, 16'd49051, 16'd60, 16'd18036, 16'd47899, 16'd49800, 16'd2861, 16'd51870, 16'd3002, 16'd12009, 16'd7748, 16'd26354, 16'd49235, 16'd44944, 16'd7957, 16'd2411, 16'd14207, 16'd18013, 16'd9314, 16'd51350, 16'd38929, 16'd57953, 16'd43311, 16'd50349});
	test_expansion(128'h61963234be4f34b631cdbeff4e125b13, {16'd7825, 16'd45324, 16'd6684, 16'd59232, 16'd5304, 16'd60021, 16'd51381, 16'd47803, 16'd25573, 16'd1871, 16'd29704, 16'd37772, 16'd44806, 16'd12587, 16'd27665, 16'd22963, 16'd8795, 16'd38445, 16'd13758, 16'd63434, 16'd26594, 16'd35158, 16'd338, 16'd56631, 16'd23678, 16'd63984});
	test_expansion(128'hdeb192dc19c1327335d8c8c58c722ba1, {16'd42004, 16'd50129, 16'd15874, 16'd31346, 16'd51194, 16'd6674, 16'd58807, 16'd14448, 16'd45042, 16'd61954, 16'd22650, 16'd62800, 16'd5354, 16'd38023, 16'd33050, 16'd14164, 16'd40836, 16'd3219, 16'd31265, 16'd30148, 16'd44241, 16'd30765, 16'd19650, 16'd35791, 16'd49252, 16'd2318});
	test_expansion(128'h0fa7c7acd123cdad4092df97e0a3f6ad, {16'd35956, 16'd16792, 16'd4681, 16'd31095, 16'd39821, 16'd2506, 16'd10709, 16'd45856, 16'd48197, 16'd55868, 16'd40295, 16'd56720, 16'd46174, 16'd55323, 16'd45874, 16'd7850, 16'd42381, 16'd41218, 16'd61195, 16'd57298, 16'd5965, 16'd31566, 16'd19098, 16'd25998, 16'd17531, 16'd33521});
	test_expansion(128'h21dc04d4ffa44200c3494b0ac3d55d7d, {16'd2700, 16'd57520, 16'd7690, 16'd5212, 16'd34573, 16'd40341, 16'd6598, 16'd36212, 16'd26232, 16'd57306, 16'd31068, 16'd8384, 16'd15414, 16'd26472, 16'd62757, 16'd2148, 16'd15613, 16'd26372, 16'd58305, 16'd58933, 16'd26198, 16'd1615, 16'd32169, 16'd52178, 16'd49488, 16'd11581});
	test_expansion(128'h17ab21d69a13c11547bd7d1ee2e6226b, {16'd50202, 16'd51112, 16'd43878, 16'd1985, 16'd35348, 16'd34954, 16'd24492, 16'd4009, 16'd24700, 16'd15699, 16'd62767, 16'd16868, 16'd12752, 16'd1098, 16'd36921, 16'd894, 16'd8272, 16'd7446, 16'd53423, 16'd24467, 16'd43622, 16'd63411, 16'd16842, 16'd15325, 16'd12729, 16'd61282});
	test_expansion(128'h4b69cf160ad69d8aa33914288baa82e4, {16'd24137, 16'd42339, 16'd14759, 16'd8777, 16'd35988, 16'd27220, 16'd1247, 16'd46780, 16'd55643, 16'd9716, 16'd63340, 16'd5157, 16'd12211, 16'd8906, 16'd42135, 16'd61273, 16'd56106, 16'd20635, 16'd57005, 16'd49678, 16'd26244, 16'd17796, 16'd43476, 16'd30899, 16'd49141, 16'd34074});
	test_expansion(128'hd095b45626a067940532725007250961, {16'd62819, 16'd36025, 16'd8059, 16'd24332, 16'd49848, 16'd61508, 16'd40050, 16'd62681, 16'd46913, 16'd48954, 16'd41410, 16'd48334, 16'd34769, 16'd58128, 16'd35741, 16'd57391, 16'd7866, 16'd2613, 16'd47778, 16'd14293, 16'd11123, 16'd45520, 16'd24571, 16'd24784, 16'd38930, 16'd64708});
	test_expansion(128'hc152627c9813ab1a9fd204b0b2cb044c, {16'd55750, 16'd51628, 16'd57816, 16'd18272, 16'd54639, 16'd44165, 16'd12740, 16'd44000, 16'd62174, 16'd35, 16'd20385, 16'd55608, 16'd4181, 16'd37799, 16'd16405, 16'd8889, 16'd33954, 16'd49747, 16'd29148, 16'd4919, 16'd44054, 16'd31550, 16'd49194, 16'd64771, 16'd61661, 16'd11707});
	test_expansion(128'h4c4c0922bcab21e20d89ce9178b191c4, {16'd4914, 16'd29467, 16'd40179, 16'd3772, 16'd14050, 16'd25152, 16'd12607, 16'd11444, 16'd1524, 16'd20745, 16'd62591, 16'd58566, 16'd54479, 16'd30918, 16'd33385, 16'd47923, 16'd57374, 16'd20756, 16'd11622, 16'd37651, 16'd51193, 16'd14967, 16'd19209, 16'd4286, 16'd4880, 16'd34504});
	test_expansion(128'h20ea1cfa6e78b369214a8df6b996c8e6, {16'd13252, 16'd18015, 16'd50059, 16'd55525, 16'd25029, 16'd14955, 16'd60990, 16'd8215, 16'd47692, 16'd61459, 16'd51864, 16'd63106, 16'd18978, 16'd43109, 16'd10575, 16'd28829, 16'd44266, 16'd46313, 16'd12121, 16'd50128, 16'd48517, 16'd27061, 16'd15917, 16'd5820, 16'd31156, 16'd59300});
	test_expansion(128'h4be1892cac6ac42ae0b4c7a19130895b, {16'd20489, 16'd346, 16'd1256, 16'd44104, 16'd47126, 16'd43487, 16'd41686, 16'd46594, 16'd56461, 16'd63471, 16'd46705, 16'd13868, 16'd44131, 16'd39193, 16'd39740, 16'd32636, 16'd40697, 16'd59770, 16'd47440, 16'd42577, 16'd55411, 16'd46138, 16'd20945, 16'd4325, 16'd11639, 16'd10410});
	test_expansion(128'h07f40c43430676fc5cdb14ebdf8e3b6c, {16'd33701, 16'd28026, 16'd61597, 16'd36933, 16'd8882, 16'd7880, 16'd39695, 16'd29327, 16'd26954, 16'd2059, 16'd52464, 16'd5774, 16'd44966, 16'd20788, 16'd47330, 16'd24275, 16'd55764, 16'd61155, 16'd61563, 16'd18325, 16'd62934, 16'd7290, 16'd33078, 16'd26966, 16'd56229, 16'd56878});
	test_expansion(128'h99c429de402220c49fbdf1bbc64a5b88, {16'd38760, 16'd14029, 16'd24901, 16'd31675, 16'd27572, 16'd16797, 16'd32306, 16'd7561, 16'd60585, 16'd43463, 16'd39369, 16'd61601, 16'd44990, 16'd25866, 16'd47766, 16'd4316, 16'd10575, 16'd19882, 16'd46212, 16'd13732, 16'd31242, 16'd43736, 16'd20125, 16'd53920, 16'd59878, 16'd42202});
	test_expansion(128'h98713b33441e10d5888f461fa0deab59, {16'd44501, 16'd23027, 16'd58231, 16'd11893, 16'd20083, 16'd52934, 16'd59635, 16'd27452, 16'd39352, 16'd12240, 16'd5673, 16'd4961, 16'd14586, 16'd10864, 16'd3097, 16'd5661, 16'd47887, 16'd32641, 16'd5907, 16'd32434, 16'd8553, 16'd25493, 16'd51471, 16'd32327, 16'd31711, 16'd61582});
	test_expansion(128'h3489691a494e822c6007736cc1a6ed19, {16'd58409, 16'd61505, 16'd6765, 16'd36536, 16'd4039, 16'd47034, 16'd30146, 16'd10271, 16'd58309, 16'd9581, 16'd58931, 16'd34992, 16'd42561, 16'd1060, 16'd5792, 16'd38379, 16'd64517, 16'd34351, 16'd31529, 16'd47924, 16'd38497, 16'd47462, 16'd11416, 16'd35545, 16'd45838, 16'd57588});
	test_expansion(128'haabbe76a6eedee49a66e9e54607f0d55, {16'd52248, 16'd9605, 16'd21789, 16'd41194, 16'd54604, 16'd45509, 16'd33219, 16'd17242, 16'd37349, 16'd28695, 16'd36283, 16'd763, 16'd9421, 16'd56313, 16'd29979, 16'd42897, 16'd45730, 16'd61860, 16'd52585, 16'd47768, 16'd53527, 16'd8841, 16'd24426, 16'd37223, 16'd51530, 16'd57198});
	test_expansion(128'hfa30c3610cf55e0921976d7055557f17, {16'd19269, 16'd44572, 16'd48943, 16'd62542, 16'd39351, 16'd33183, 16'd15275, 16'd57168, 16'd45829, 16'd31790, 16'd41193, 16'd43918, 16'd28247, 16'd32992, 16'd25089, 16'd62553, 16'd19368, 16'd26789, 16'd34756, 16'd57584, 16'd65379, 16'd27005, 16'd42941, 16'd56408, 16'd33646, 16'd42160});
	test_expansion(128'h21768a54a684e9faca0c460a6b865755, {16'd24123, 16'd5384, 16'd46365, 16'd14195, 16'd3113, 16'd50253, 16'd24596, 16'd34186, 16'd43219, 16'd7149, 16'd61085, 16'd49330, 16'd14276, 16'd57171, 16'd29847, 16'd37862, 16'd47111, 16'd59471, 16'd21899, 16'd17703, 16'd63414, 16'd49030, 16'd53764, 16'd33560, 16'd5412, 16'd33463});
	test_expansion(128'h0996bec44b1aaadee270fddc9ca0ada4, {16'd46918, 16'd13636, 16'd16234, 16'd42560, 16'd61957, 16'd47660, 16'd62281, 16'd47735, 16'd23588, 16'd59501, 16'd26261, 16'd13572, 16'd17441, 16'd53786, 16'd33133, 16'd27736, 16'd61065, 16'd61258, 16'd683, 16'd20111, 16'd24923, 16'd12684, 16'd48706, 16'd14636, 16'd41081, 16'd29729});
	test_expansion(128'hb7894013119927522d7ffb5f7ac5d560, {16'd9017, 16'd55418, 16'd14470, 16'd12414, 16'd32271, 16'd26023, 16'd13950, 16'd57122, 16'd14950, 16'd35136, 16'd22259, 16'd50240, 16'd22939, 16'd731, 16'd43526, 16'd7281, 16'd27532, 16'd56843, 16'd45697, 16'd17555, 16'd41200, 16'd26957, 16'd41522, 16'd58304, 16'd32298, 16'd61743});
	test_expansion(128'h7c45f8f46a2430678715d601f4ef6bc6, {16'd48023, 16'd6314, 16'd47668, 16'd44279, 16'd55635, 16'd19880, 16'd51065, 16'd47869, 16'd48004, 16'd24917, 16'd11788, 16'd15085, 16'd19675, 16'd49774, 16'd42302, 16'd5053, 16'd36298, 16'd52926, 16'd3633, 16'd23314, 16'd28756, 16'd27531, 16'd30934, 16'd18075, 16'd47264, 16'd24449});
	test_expansion(128'h8389bbe22d3f388f7da0cbf9f7885e67, {16'd35772, 16'd12683, 16'd16881, 16'd12970, 16'd27760, 16'd24103, 16'd43322, 16'd37264, 16'd48888, 16'd18501, 16'd21610, 16'd62028, 16'd24148, 16'd50130, 16'd59634, 16'd25028, 16'd8852, 16'd58610, 16'd44624, 16'd47040, 16'd50128, 16'd58852, 16'd41826, 16'd45632, 16'd60356, 16'd9296});
	test_expansion(128'h0c0e0055ce0f33cf90890ce0e5b1a7f9, {16'd62157, 16'd29790, 16'd31632, 16'd60501, 16'd2712, 16'd55782, 16'd43406, 16'd44756, 16'd4282, 16'd23597, 16'd30246, 16'd37897, 16'd53767, 16'd50214, 16'd32869, 16'd58323, 16'd42264, 16'd41276, 16'd48315, 16'd36384, 16'd45416, 16'd7026, 16'd61705, 16'd36705, 16'd36003, 16'd22948});
	test_expansion(128'h61c2e9100fe3bb9cfc22304c2c4021f1, {16'd6542, 16'd29250, 16'd24859, 16'd29465, 16'd51374, 16'd48364, 16'd39289, 16'd35305, 16'd41946, 16'd56313, 16'd53387, 16'd18397, 16'd57183, 16'd2532, 16'd57817, 16'd27437, 16'd7918, 16'd56552, 16'd3645, 16'd916, 16'd54137, 16'd62784, 16'd159, 16'd17384, 16'd8628, 16'd27775});
	test_expansion(128'he183497b574026eda6192d5e682d057f, {16'd31029, 16'd30764, 16'd20343, 16'd17770, 16'd43863, 16'd64920, 16'd22410, 16'd2234, 16'd51342, 16'd49374, 16'd19195, 16'd42314, 16'd49550, 16'd13229, 16'd38938, 16'd13737, 16'd45406, 16'd12665, 16'd46573, 16'd65505, 16'd30464, 16'd34504, 16'd57413, 16'd62199, 16'd47020, 16'd45578});
	test_expansion(128'hd06c621f849be94e80dd51498c304416, {16'd7185, 16'd33921, 16'd25633, 16'd20329, 16'd51601, 16'd43385, 16'd59251, 16'd46642, 16'd5009, 16'd27582, 16'd59293, 16'd41565, 16'd6022, 16'd14811, 16'd57350, 16'd11334, 16'd21780, 16'd35282, 16'd28915, 16'd58695, 16'd26194, 16'd39041, 16'd56884, 16'd61467, 16'd1231, 16'd10333});
	test_expansion(128'h6f511c33539f9b527439d6fc237f804e, {16'd11986, 16'd14459, 16'd13769, 16'd48702, 16'd15245, 16'd7601, 16'd37594, 16'd61932, 16'd58360, 16'd23544, 16'd42079, 16'd37323, 16'd7603, 16'd62940, 16'd16525, 16'd34512, 16'd3990, 16'd8243, 16'd49511, 16'd16956, 16'd8286, 16'd19735, 16'd30680, 16'd12076, 16'd8730, 16'd42913});
	test_expansion(128'h4f8a186b057f30b6bacbb2af6066857b, {16'd47933, 16'd16505, 16'd47633, 16'd14461, 16'd44091, 16'd29040, 16'd13904, 16'd2019, 16'd17067, 16'd23425, 16'd52255, 16'd55106, 16'd41516, 16'd20232, 16'd35397, 16'd7075, 16'd60390, 16'd54909, 16'd2965, 16'd52092, 16'd62575, 16'd20238, 16'd18871, 16'd37044, 16'd42424, 16'd45426});
	test_expansion(128'h3f4349ac4b69fcfb6efecd8d2060664f, {16'd5727, 16'd30245, 16'd15238, 16'd62526, 16'd8841, 16'd46381, 16'd1450, 16'd54250, 16'd3346, 16'd13635, 16'd36813, 16'd64314, 16'd1015, 16'd19542, 16'd49152, 16'd52825, 16'd64809, 16'd32554, 16'd64475, 16'd61964, 16'd32903, 16'd25997, 16'd54765, 16'd57878, 16'd1372, 16'd60727});
	test_expansion(128'h7e8c9747b8663d2086165fb742b59642, {16'd1959, 16'd31001, 16'd61458, 16'd47976, 16'd21785, 16'd40678, 16'd42798, 16'd20287, 16'd7824, 16'd51482, 16'd59557, 16'd50257, 16'd47689, 16'd1411, 16'd3790, 16'd17761, 16'd60285, 16'd1311, 16'd59567, 16'd32479, 16'd25602, 16'd51059, 16'd59277, 16'd55844, 16'd54306, 16'd64883});
	test_expansion(128'ha6ba88214f9260667900151ad22338ed, {16'd23851, 16'd20414, 16'd39125, 16'd49222, 16'd33920, 16'd14632, 16'd15756, 16'd54661, 16'd61475, 16'd43959, 16'd32983, 16'd63951, 16'd51780, 16'd65521, 16'd30459, 16'd3476, 16'd6758, 16'd20133, 16'd64103, 16'd3841, 16'd1425, 16'd30234, 16'd4994, 16'd49712, 16'd31996, 16'd62370});
	test_expansion(128'h0433ee8a99a9dc6b2a93e7be34429b54, {16'd12100, 16'd2685, 16'd63219, 16'd17402, 16'd40305, 16'd9327, 16'd58320, 16'd30562, 16'd12956, 16'd19934, 16'd3417, 16'd54943, 16'd49346, 16'd3936, 16'd45129, 16'd54737, 16'd22374, 16'd6730, 16'd33547, 16'd8681, 16'd4614, 16'd17075, 16'd61539, 16'd52094, 16'd3757, 16'd21748});
	test_expansion(128'hd494ec151dcb85394e007126729b37b7, {16'd24700, 16'd18327, 16'd18543, 16'd27716, 16'd14271, 16'd18582, 16'd64810, 16'd14971, 16'd50517, 16'd33270, 16'd1048, 16'd50893, 16'd11660, 16'd45167, 16'd22136, 16'd5981, 16'd41719, 16'd61918, 16'd5530, 16'd65244, 16'd37407, 16'd47751, 16'd39273, 16'd40708, 16'd10436, 16'd46531});
	test_expansion(128'h9ae419a4dd0b55e8f5659c88455706a9, {16'd7026, 16'd20625, 16'd58603, 16'd65323, 16'd30964, 16'd26042, 16'd63918, 16'd47720, 16'd12041, 16'd41803, 16'd21433, 16'd53787, 16'd20587, 16'd26261, 16'd41244, 16'd23637, 16'd14914, 16'd17604, 16'd8263, 16'd23864, 16'd14130, 16'd47958, 16'd39616, 16'd9510, 16'd6872, 16'd24132});
	test_expansion(128'h5d032d6fd9df1796f4bb87d6323719c0, {16'd3047, 16'd4607, 16'd6392, 16'd42677, 16'd23469, 16'd42668, 16'd271, 16'd30140, 16'd57895, 16'd21792, 16'd971, 16'd8512, 16'd31084, 16'd30032, 16'd5290, 16'd16555, 16'd58636, 16'd44737, 16'd64801, 16'd33370, 16'd55676, 16'd22308, 16'd7483, 16'd63775, 16'd48694, 16'd20248});
	test_expansion(128'h953fccf91e5c998534896d57c0f76ff3, {16'd49491, 16'd52731, 16'd60021, 16'd64513, 16'd11131, 16'd12592, 16'd24899, 16'd3649, 16'd5555, 16'd5108, 16'd38630, 16'd16213, 16'd8540, 16'd26990, 16'd58223, 16'd1522, 16'd4464, 16'd46991, 16'd1814, 16'd29690, 16'd17272, 16'd42190, 16'd54155, 16'd21266, 16'd38594, 16'd25282});
	test_expansion(128'h6f891c134deb60ff46f22c6f3464f1bb, {16'd32345, 16'd55317, 16'd1835, 16'd16120, 16'd40870, 16'd55570, 16'd2917, 16'd64402, 16'd22693, 16'd34613, 16'd724, 16'd6005, 16'd51800, 16'd6339, 16'd60104, 16'd49739, 16'd22610, 16'd24531, 16'd5301, 16'd53337, 16'd25534, 16'd7125, 16'd46968, 16'd38250, 16'd45855, 16'd15810});
	test_expansion(128'h08f7bc6b4e666d5d484d7598d98a5aea, {16'd38264, 16'd48133, 16'd60879, 16'd15247, 16'd29265, 16'd22946, 16'd2072, 16'd14965, 16'd24886, 16'd53245, 16'd50814, 16'd29472, 16'd58809, 16'd28945, 16'd24314, 16'd59400, 16'd16583, 16'd43187, 16'd9386, 16'd34329, 16'd2165, 16'd65420, 16'd65073, 16'd30698, 16'd44027, 16'd9775});
	test_expansion(128'h1bbab5de31ea90ff729c0decf56da61a, {16'd5828, 16'd5060, 16'd23105, 16'd22440, 16'd45530, 16'd61859, 16'd25515, 16'd1317, 16'd19142, 16'd17681, 16'd4594, 16'd18346, 16'd65514, 16'd26105, 16'd46279, 16'd31407, 16'd16579, 16'd18276, 16'd40132, 16'd18747, 16'd59732, 16'd65259, 16'd54744, 16'd29350, 16'd2468, 16'd37062});
	test_expansion(128'he4f68ade4cd985fa2fae6adb512629ff, {16'd59435, 16'd48182, 16'd40180, 16'd19169, 16'd32408, 16'd27627, 16'd21716, 16'd34325, 16'd53713, 16'd56276, 16'd23026, 16'd45166, 16'd58173, 16'd57173, 16'd57659, 16'd62732, 16'd14371, 16'd1955, 16'd59521, 16'd51510, 16'd28662, 16'd58242, 16'd297, 16'd33801, 16'd43565, 16'd18633});
	test_expansion(128'h8cba566eb4d04616ff38c05a88fc0250, {16'd52397, 16'd389, 16'd18401, 16'd25678, 16'd25300, 16'd46448, 16'd24307, 16'd7011, 16'd17714, 16'd14683, 16'd12321, 16'd34913, 16'd54482, 16'd40675, 16'd6716, 16'd44287, 16'd60234, 16'd60767, 16'd23131, 16'd6209, 16'd26541, 16'd23749, 16'd44687, 16'd38544, 16'd17120, 16'd53881});
	test_expansion(128'hb2584e3c0b5d6aff194086beac35d61f, {16'd24939, 16'd11346, 16'd23724, 16'd17478, 16'd32494, 16'd34169, 16'd12036, 16'd45358, 16'd65323, 16'd63293, 16'd22778, 16'd29329, 16'd60543, 16'd2384, 16'd1337, 16'd25468, 16'd52152, 16'd28030, 16'd15984, 16'd31020, 16'd6843, 16'd30474, 16'd44108, 16'd5845, 16'd7119, 16'd20127});
	test_expansion(128'hadc232e0fc151b35414592d6450fae77, {16'd19293, 16'd32603, 16'd16863, 16'd29820, 16'd24522, 16'd51441, 16'd20187, 16'd10401, 16'd45735, 16'd1563, 16'd45457, 16'd16946, 16'd50125, 16'd6170, 16'd21094, 16'd39548, 16'd46281, 16'd9530, 16'd54927, 16'd28735, 16'd23635, 16'd25518, 16'd17332, 16'd32475, 16'd23935, 16'd12598});
	test_expansion(128'h2e3ad5371ab954e96122142235ffa527, {16'd21206, 16'd61358, 16'd56674, 16'd30171, 16'd63791, 16'd63055, 16'd11161, 16'd58731, 16'd25379, 16'd56864, 16'd53641, 16'd13946, 16'd42592, 16'd29229, 16'd34177, 16'd49619, 16'd18533, 16'd45246, 16'd18279, 16'd21015, 16'd19996, 16'd1499, 16'd47098, 16'd27570, 16'd58186, 16'd40533});
	test_expansion(128'h7e25e4b354aaeaf4c5ab026364d6bcb5, {16'd144, 16'd39368, 16'd31554, 16'd65029, 16'd15681, 16'd51106, 16'd56752, 16'd27991, 16'd54191, 16'd31560, 16'd12884, 16'd18960, 16'd63279, 16'd62435, 16'd17635, 16'd22486, 16'd21314, 16'd62692, 16'd56480, 16'd18669, 16'd10672, 16'd7611, 16'd2454, 16'd47008, 16'd15600, 16'd6610});
	test_expansion(128'hf3bfbda24143941bca6d025d61b44062, {16'd26022, 16'd37047, 16'd43109, 16'd5808, 16'd12463, 16'd18173, 16'd7620, 16'd43959, 16'd49172, 16'd562, 16'd6627, 16'd59912, 16'd11862, 16'd482, 16'd21448, 16'd5889, 16'd14331, 16'd63700, 16'd4464, 16'd58220, 16'd60219, 16'd16066, 16'd31416, 16'd46720, 16'd8205, 16'd22339});
	test_expansion(128'hb9d59d919af4521ae113587a7d5a794b, {16'd32428, 16'd49070, 16'd44158, 16'd13683, 16'd59033, 16'd35115, 16'd28581, 16'd28181, 16'd48234, 16'd13051, 16'd46323, 16'd17333, 16'd38035, 16'd45270, 16'd53010, 16'd10556, 16'd47468, 16'd51288, 16'd12107, 16'd24559, 16'd18701, 16'd41753, 16'd16014, 16'd12802, 16'd7301, 16'd6942});
	test_expansion(128'hf13a7a0a8d15ac1246f4c9ac46dd8062, {16'd14088, 16'd61237, 16'd65424, 16'd31421, 16'd4345, 16'd24633, 16'd12044, 16'd42305, 16'd12911, 16'd54382, 16'd53820, 16'd34435, 16'd5341, 16'd24988, 16'd51121, 16'd13323, 16'd64330, 16'd41532, 16'd19999, 16'd26226, 16'd38898, 16'd16057, 16'd7509, 16'd61317, 16'd39378, 16'd50645});
	test_expansion(128'h67b6d9c620249eaff7eaaac98ea7450b, {16'd6840, 16'd7798, 16'd39703, 16'd3351, 16'd53251, 16'd14334, 16'd4308, 16'd61366, 16'd63784, 16'd41919, 16'd34351, 16'd35466, 16'd47085, 16'd16860, 16'd18608, 16'd49159, 16'd43864, 16'd38619, 16'd46522, 16'd14248, 16'd41720, 16'd4249, 16'd17742, 16'd20682, 16'd34781, 16'd50879});
	test_expansion(128'ha64015dcfdefb6fb35665ce0bb2d2a3e, {16'd63009, 16'd10661, 16'd45036, 16'd10834, 16'd42561, 16'd61733, 16'd50153, 16'd52334, 16'd65058, 16'd13070, 16'd16252, 16'd14168, 16'd58430, 16'd60300, 16'd38446, 16'd35102, 16'd56479, 16'd314, 16'd46014, 16'd39496, 16'd32498, 16'd25470, 16'd17955, 16'd39257, 16'd25904, 16'd27813});
	test_expansion(128'h1196543eca19f2906217292500a7cf83, {16'd51643, 16'd20902, 16'd27291, 16'd54163, 16'd30394, 16'd12304, 16'd39125, 16'd18539, 16'd63902, 16'd27848, 16'd51448, 16'd39079, 16'd60190, 16'd56889, 16'd9285, 16'd52954, 16'd26714, 16'd40761, 16'd45270, 16'd22646, 16'd8231, 16'd27759, 16'd11616, 16'd10831, 16'd17738, 16'd61071});
	test_expansion(128'hb31e5a24a26c8d7caa6159410adb2cb6, {16'd22973, 16'd51101, 16'd49228, 16'd30837, 16'd26447, 16'd6592, 16'd56561, 16'd45649, 16'd34019, 16'd3124, 16'd24241, 16'd26526, 16'd59075, 16'd57498, 16'd19277, 16'd35838, 16'd33183, 16'd13798, 16'd326, 16'd40169, 16'd60887, 16'd23598, 16'd29029, 16'd18424, 16'd20375, 16'd12294});
	test_expansion(128'h36a4f61fc5a1f7d3271314a96da7afe3, {16'd15674, 16'd25884, 16'd61300, 16'd862, 16'd2038, 16'd13281, 16'd56780, 16'd29836, 16'd225, 16'd50466, 16'd56227, 16'd20307, 16'd62969, 16'd65114, 16'd36542, 16'd38316, 16'd22609, 16'd59323, 16'd28849, 16'd63143, 16'd15213, 16'd7991, 16'd21153, 16'd39317, 16'd40143, 16'd61426});
	test_expansion(128'h03eadcfc42af4a8f0ddddbc837c22683, {16'd12400, 16'd42824, 16'd59731, 16'd50073, 16'd64627, 16'd41296, 16'd62399, 16'd29799, 16'd45251, 16'd44581, 16'd52592, 16'd57380, 16'd63957, 16'd26750, 16'd31970, 16'd4649, 16'd28953, 16'd22141, 16'd21462, 16'd41984, 16'd23649, 16'd61776, 16'd2765, 16'd36898, 16'd50684, 16'd24344});
	test_expansion(128'h7108f04feb72b8d2e659c31ac27734b4, {16'd17882, 16'd23122, 16'd52276, 16'd1109, 16'd18154, 16'd53636, 16'd8729, 16'd46229, 16'd65005, 16'd43235, 16'd2115, 16'd5116, 16'd24772, 16'd65390, 16'd40429, 16'd45731, 16'd51319, 16'd20512, 16'd18886, 16'd14938, 16'd33384, 16'd23950, 16'd16985, 16'd44220, 16'd12389, 16'd19671});
	test_expansion(128'hbda0ed4e6889f92e4794c0cb47ffe1f3, {16'd12938, 16'd50600, 16'd8308, 16'd55717, 16'd42949, 16'd39919, 16'd27799, 16'd15252, 16'd34749, 16'd24775, 16'd27913, 16'd25751, 16'd28401, 16'd18665, 16'd4694, 16'd28802, 16'd29683, 16'd62808, 16'd20649, 16'd20309, 16'd15412, 16'd34039, 16'd34342, 16'd17088, 16'd41033, 16'd24964});
	test_expansion(128'h9aaff6644b6b835f9636a10e493478f8, {16'd43317, 16'd49328, 16'd24061, 16'd18012, 16'd59799, 16'd38327, 16'd30929, 16'd41956, 16'd49845, 16'd27449, 16'd9294, 16'd61619, 16'd60640, 16'd25619, 16'd38423, 16'd63577, 16'd47912, 16'd55277, 16'd34080, 16'd21810, 16'd46495, 16'd28491, 16'd51665, 16'd45382, 16'd6349, 16'd61669});
	test_expansion(128'h430fd2f57136de0ff88aa5f20bfb04f8, {16'd47684, 16'd32520, 16'd43079, 16'd52853, 16'd44377, 16'd1048, 16'd13104, 16'd59125, 16'd48117, 16'd25430, 16'd18060, 16'd11376, 16'd61812, 16'd12693, 16'd44205, 16'd33414, 16'd43726, 16'd14704, 16'd27354, 16'd25860, 16'd5472, 16'd3470, 16'd15875, 16'd55129, 16'd27875, 16'd46272});
	test_expansion(128'ha69012702fc2e455c5804e0455040978, {16'd19584, 16'd20625, 16'd59654, 16'd30181, 16'd14409, 16'd41949, 16'd51036, 16'd43514, 16'd25089, 16'd45771, 16'd10459, 16'd36716, 16'd36113, 16'd61766, 16'd7254, 16'd23510, 16'd6177, 16'd44178, 16'd43758, 16'd29949, 16'd59108, 16'd38180, 16'd16530, 16'd32233, 16'd15029, 16'd35357});
	test_expansion(128'h0371c50ad1aad9d7865f3e111e7d98ef, {16'd49882, 16'd41119, 16'd13568, 16'd20961, 16'd9612, 16'd24152, 16'd21124, 16'd57951, 16'd24462, 16'd17350, 16'd9325, 16'd26790, 16'd42835, 16'd10543, 16'd56951, 16'd50995, 16'd41055, 16'd21871, 16'd7153, 16'd50100, 16'd80, 16'd5358, 16'd50396, 16'd8523, 16'd55335, 16'd51710});
	test_expansion(128'h0610f88751ca0748550fafaa2d0050a9, {16'd6832, 16'd18471, 16'd37233, 16'd5734, 16'd12119, 16'd59195, 16'd17907, 16'd13735, 16'd16282, 16'd57363, 16'd3296, 16'd16782, 16'd804, 16'd27781, 16'd32222, 16'd31046, 16'd11675, 16'd10925, 16'd60165, 16'd33938, 16'd42111, 16'd53065, 16'd53932, 16'd17210, 16'd2690, 16'd20176});
	test_expansion(128'hb5cf1ce9352da0480ad87d47de016014, {16'd6072, 16'd40222, 16'd19616, 16'd59866, 16'd61749, 16'd58188, 16'd59884, 16'd13684, 16'd58647, 16'd36705, 16'd276, 16'd50450, 16'd8479, 16'd37140, 16'd6781, 16'd44348, 16'd8901, 16'd50290, 16'd44213, 16'd34571, 16'd64157, 16'd32798, 16'd25819, 16'd48271, 16'd10435, 16'd43641});
	test_expansion(128'h2a8c80e4be76d5ef6f3b99f2f11fcd7c, {16'd19957, 16'd41934, 16'd2241, 16'd25031, 16'd4649, 16'd15639, 16'd52143, 16'd42247, 16'd63397, 16'd5808, 16'd3329, 16'd35217, 16'd23662, 16'd15643, 16'd16120, 16'd63540, 16'd33297, 16'd46742, 16'd10757, 16'd62823, 16'd536, 16'd59409, 16'd51683, 16'd35448, 16'd34216, 16'd11254});
	test_expansion(128'h0eaba8ad6e6cfe321abcc46fe955c14f, {16'd7534, 16'd2645, 16'd61822, 16'd61855, 16'd23637, 16'd20906, 16'd21869, 16'd33656, 16'd25172, 16'd53388, 16'd3932, 16'd13512, 16'd25809, 16'd55790, 16'd14622, 16'd23103, 16'd7975, 16'd25196, 16'd33318, 16'd17343, 16'd65191, 16'd46901, 16'd38901, 16'd54981, 16'd35159, 16'd54005});
	test_expansion(128'hfd7a1ac37f43935a51f624276c6f1dc7, {16'd25452, 16'd4344, 16'd17727, 16'd50413, 16'd472, 16'd51161, 16'd211, 16'd36475, 16'd16709, 16'd5702, 16'd6332, 16'd62316, 16'd26278, 16'd14445, 16'd46924, 16'd30259, 16'd11186, 16'd12701, 16'd50495, 16'd51639, 16'd54849, 16'd61477, 16'd37212, 16'd56029, 16'd34627, 16'd22263});
	test_expansion(128'he1846d5bf624659bea9cc5aad904df83, {16'd41752, 16'd35461, 16'd17060, 16'd33558, 16'd43918, 16'd10520, 16'd28060, 16'd6479, 16'd46674, 16'd45362, 16'd22496, 16'd10276, 16'd10460, 16'd49900, 16'd58167, 16'd30227, 16'd65348, 16'd26858, 16'd1092, 16'd14713, 16'd13492, 16'd2451, 16'd35716, 16'd39664, 16'd47643, 16'd6629});
	test_expansion(128'h1901a75e780fb44d2b9593f7068d8314, {16'd15773, 16'd19751, 16'd58845, 16'd34543, 16'd19868, 16'd39385, 16'd15462, 16'd8967, 16'd1419, 16'd21148, 16'd39098, 16'd59775, 16'd16126, 16'd2547, 16'd40250, 16'd24053, 16'd47748, 16'd14142, 16'd47100, 16'd558, 16'd27406, 16'd4526, 16'd29362, 16'd14557, 16'd22729, 16'd21909});
	test_expansion(128'h1ffd10d1a5f31adf80530894b648bb39, {16'd30111, 16'd52962, 16'd50807, 16'd59745, 16'd11801, 16'd31531, 16'd2206, 16'd10875, 16'd37167, 16'd43231, 16'd21895, 16'd59800, 16'd28931, 16'd60338, 16'd31736, 16'd60408, 16'd18695, 16'd25801, 16'd38395, 16'd35494, 16'd24562, 16'd3994, 16'd59161, 16'd16946, 16'd57921, 16'd54088});
	test_expansion(128'h690eeb1204ee51da5316d7686a0cbe88, {16'd3177, 16'd54085, 16'd34387, 16'd63971, 16'd63130, 16'd30357, 16'd13295, 16'd6014, 16'd3879, 16'd13676, 16'd31539, 16'd35891, 16'd9878, 16'd7862, 16'd59555, 16'd4402, 16'd8804, 16'd38914, 16'd44351, 16'd3653, 16'd2657, 16'd20705, 16'd28029, 16'd31128, 16'd63780, 16'd52502});
	test_expansion(128'h9924bd84fde8884b238738d1d5ac85e0, {16'd52300, 16'd2560, 16'd30652, 16'd646, 16'd27460, 16'd24231, 16'd64606, 16'd51142, 16'd38461, 16'd1469, 16'd1475, 16'd9116, 16'd17848, 16'd40551, 16'd29521, 16'd2261, 16'd47150, 16'd829, 16'd49982, 16'd26685, 16'd57401, 16'd39672, 16'd50758, 16'd14064, 16'd59595, 16'd1153});
	test_expansion(128'he45fc1982ca249eff4de0fd2c7bf12b0, {16'd21225, 16'd9672, 16'd38324, 16'd19887, 16'd51713, 16'd64094, 16'd63651, 16'd4705, 16'd34382, 16'd51803, 16'd21620, 16'd50524, 16'd13272, 16'd30682, 16'd64632, 16'd44748, 16'd26280, 16'd56539, 16'd41180, 16'd19034, 16'd41344, 16'd8829, 16'd47324, 16'd19018, 16'd21082, 16'd31639});
	test_expansion(128'h961af09a8c5c1fdf18b059d94215e3ca, {16'd56919, 16'd23056, 16'd6085, 16'd4861, 16'd55272, 16'd10637, 16'd9394, 16'd36088, 16'd29033, 16'd4674, 16'd12519, 16'd30933, 16'd46434, 16'd63440, 16'd63017, 16'd1856, 16'd50441, 16'd33943, 16'd26107, 16'd27587, 16'd21115, 16'd43865, 16'd11599, 16'd14356, 16'd41537, 16'd23361});
	test_expansion(128'h297dd1df9e1f3bad94f6cf9a31c6e563, {16'd13240, 16'd11528, 16'd21586, 16'd20999, 16'd19189, 16'd29133, 16'd18426, 16'd26064, 16'd49823, 16'd6258, 16'd14611, 16'd24270, 16'd59475, 16'd27162, 16'd21480, 16'd60692, 16'd62135, 16'd17900, 16'd53726, 16'd30869, 16'd35168, 16'd36719, 16'd21214, 16'd18510, 16'd40122, 16'd57584});
	test_expansion(128'haa34010830dd4b8ae9cdee1e7faae039, {16'd23179, 16'd44518, 16'd63345, 16'd33926, 16'd52035, 16'd45576, 16'd13623, 16'd9709, 16'd15923, 16'd20196, 16'd8916, 16'd16460, 16'd47354, 16'd4351, 16'd60967, 16'd4223, 16'd28336, 16'd1257, 16'd62574, 16'd2581, 16'd19676, 16'd27123, 16'd4759, 16'd42192, 16'd6646, 16'd36019});
	test_expansion(128'h02d364f601a4adbdb6ce86a69b071578, {16'd10092, 16'd44698, 16'd9995, 16'd40574, 16'd36085, 16'd32176, 16'd12151, 16'd28388, 16'd41549, 16'd18481, 16'd37555, 16'd26913, 16'd4135, 16'd35965, 16'd24828, 16'd47854, 16'd23245, 16'd45919, 16'd54866, 16'd54643, 16'd6523, 16'd49843, 16'd38333, 16'd45701, 16'd14125, 16'd41356});
	test_expansion(128'h14eadaa351954aea28710447ae9f7ff8, {16'd16937, 16'd22199, 16'd65509, 16'd53828, 16'd2442, 16'd46435, 16'd5772, 16'd40925, 16'd34556, 16'd3764, 16'd24320, 16'd24955, 16'd36589, 16'd59143, 16'd36090, 16'd7236, 16'd22731, 16'd55283, 16'd38412, 16'd2649, 16'd39846, 16'd19516, 16'd54158, 16'd26638, 16'd26411, 16'd50714});
	test_expansion(128'h07dfb3af22184acde1cc73fdfdd59cfc, {16'd6099, 16'd14143, 16'd34069, 16'd51530, 16'd35084, 16'd58648, 16'd2759, 16'd5817, 16'd60803, 16'd32992, 16'd16633, 16'd41361, 16'd52157, 16'd30580, 16'd48771, 16'd16999, 16'd8605, 16'd59177, 16'd46605, 16'd40485, 16'd54153, 16'd62610, 16'd50077, 16'd46372, 16'd55331, 16'd43302});
	test_expansion(128'hdc8aa2ba6f7a7eb54956e315122cc529, {16'd32031, 16'd13461, 16'd47101, 16'd32591, 16'd31052, 16'd16674, 16'd61871, 16'd23083, 16'd7063, 16'd33171, 16'd10315, 16'd64302, 16'd41457, 16'd31143, 16'd13277, 16'd45220, 16'd22464, 16'd1944, 16'd1294, 16'd48946, 16'd20598, 16'd11556, 16'd51709, 16'd5249, 16'd22928, 16'd27857});
	test_expansion(128'hb87f2b791fef4c7bec64e69a3bbebef5, {16'd15003, 16'd23325, 16'd55508, 16'd40268, 16'd27194, 16'd47890, 16'd44811, 16'd26967, 16'd30526, 16'd19742, 16'd22268, 16'd63244, 16'd23822, 16'd5829, 16'd34905, 16'd1957, 16'd36083, 16'd14297, 16'd53386, 16'd37486, 16'd46915, 16'd14860, 16'd51918, 16'd23189, 16'd998, 16'd6040});
	test_expansion(128'h713361037afe035f1aeb5570e21391fc, {16'd274, 16'd29543, 16'd6303, 16'd13092, 16'd40102, 16'd22798, 16'd27651, 16'd7157, 16'd3939, 16'd11853, 16'd65095, 16'd58912, 16'd32685, 16'd55603, 16'd288, 16'd2688, 16'd36304, 16'd65003, 16'd53176, 16'd52492, 16'd6361, 16'd18106, 16'd171, 16'd21274, 16'd13361, 16'd17218});
	test_expansion(128'h32d046c855d0ad9c3968d7f4193ec6dc, {16'd29876, 16'd35955, 16'd2862, 16'd27589, 16'd30046, 16'd37565, 16'd11009, 16'd29347, 16'd56019, 16'd49147, 16'd37959, 16'd41701, 16'd9963, 16'd16508, 16'd63410, 16'd47237, 16'd37886, 16'd49590, 16'd58991, 16'd32819, 16'd26503, 16'd43928, 16'd24488, 16'd33440, 16'd61316, 16'd29565});
	test_expansion(128'h43893313a48a6193a8267d09afae7a88, {16'd61991, 16'd59678, 16'd45260, 16'd14648, 16'd37791, 16'd31769, 16'd51416, 16'd13342, 16'd50746, 16'd17383, 16'd39182, 16'd28423, 16'd10733, 16'd22821, 16'd44023, 16'd13779, 16'd41188, 16'd23873, 16'd34211, 16'd41771, 16'd8570, 16'd4988, 16'd42356, 16'd7231, 16'd5399, 16'd39084});
	test_expansion(128'hd9cf9325b4544663b1258c7a160d99dc, {16'd28533, 16'd21957, 16'd33276, 16'd22889, 16'd3535, 16'd42823, 16'd14595, 16'd63325, 16'd52340, 16'd12767, 16'd5444, 16'd6282, 16'd4891, 16'd51585, 16'd19795, 16'd26223, 16'd878, 16'd5829, 16'd52637, 16'd23330, 16'd62236, 16'd40128, 16'd28015, 16'd39980, 16'd44067, 16'd14579});
	test_expansion(128'heb2707c7d8f7cda5b1c517bf25adeae5, {16'd35863, 16'd37543, 16'd17092, 16'd14972, 16'd58957, 16'd60460, 16'd21569, 16'd10766, 16'd39596, 16'd36442, 16'd16540, 16'd56256, 16'd52799, 16'd40824, 16'd32730, 16'd3710, 16'd51629, 16'd4021, 16'd48186, 16'd8024, 16'd35918, 16'd25480, 16'd57174, 16'd19137, 16'd42616, 16'd9140});
	test_expansion(128'h55bb28af2dce2189a1debd1852f49619, {16'd48345, 16'd4604, 16'd2063, 16'd28135, 16'd30371, 16'd17608, 16'd51768, 16'd35972, 16'd14985, 16'd11284, 16'd42652, 16'd21283, 16'd50003, 16'd62041, 16'd3895, 16'd10926, 16'd38860, 16'd6267, 16'd5765, 16'd12806, 16'd40479, 16'd3350, 16'd43285, 16'd455, 16'd55074, 16'd6403});
	test_expansion(128'h1b2ac29b57eab31b5f0741baa86272af, {16'd28081, 16'd64080, 16'd46238, 16'd27000, 16'd33885, 16'd8809, 16'd11328, 16'd35087, 16'd50076, 16'd62547, 16'd49259, 16'd1740, 16'd36399, 16'd388, 16'd12801, 16'd45633, 16'd53505, 16'd14730, 16'd32614, 16'd51840, 16'd20345, 16'd55691, 16'd32731, 16'd32482, 16'd62680, 16'd6051});
	test_expansion(128'h017efce6075f498bab9988cc001d978b, {16'd33355, 16'd13590, 16'd40668, 16'd15835, 16'd22208, 16'd9142, 16'd2903, 16'd666, 16'd47227, 16'd11955, 16'd3956, 16'd4849, 16'd56587, 16'd45222, 16'd46936, 16'd47722, 16'd9732, 16'd53942, 16'd64628, 16'd27164, 16'd39830, 16'd62850, 16'd61141, 16'd45362, 16'd46742, 16'd24083});
	test_expansion(128'hd6cb39e19102f6f42c03e1248ebaf831, {16'd22411, 16'd52599, 16'd19303, 16'd47385, 16'd63286, 16'd35114, 16'd30898, 16'd53857, 16'd12643, 16'd34903, 16'd16071, 16'd5112, 16'd63153, 16'd12326, 16'd5351, 16'd54390, 16'd12397, 16'd37702, 16'd6091, 16'd9075, 16'd20955, 16'd9341, 16'd54070, 16'd7973, 16'd33877, 16'd3429});
	test_expansion(128'h590378d627e4409cec1ad455f9d7bd72, {16'd41502, 16'd13670, 16'd12858, 16'd53230, 16'd48067, 16'd51056, 16'd41794, 16'd10230, 16'd27072, 16'd27806, 16'd41215, 16'd2218, 16'd55787, 16'd5676, 16'd40664, 16'd38382, 16'd58469, 16'd43348, 16'd63631, 16'd46093, 16'd5577, 16'd47534, 16'd54991, 16'd47233, 16'd29114, 16'd19898});
	test_expansion(128'h8972522eee19f4567046ccc4a9102172, {16'd1244, 16'd58880, 16'd48559, 16'd41009, 16'd12062, 16'd42637, 16'd63071, 16'd65391, 16'd3838, 16'd50258, 16'd62763, 16'd7079, 16'd56082, 16'd23771, 16'd13558, 16'd16082, 16'd47259, 16'd4729, 16'd9665, 16'd30139, 16'd14452, 16'd43800, 16'd39552, 16'd65056, 16'd25016, 16'd43097});
	test_expansion(128'heaf4ab01edbc62443dee228d9e3ad011, {16'd39445, 16'd47562, 16'd46814, 16'd28903, 16'd39925, 16'd64753, 16'd33315, 16'd2740, 16'd8908, 16'd51201, 16'd18417, 16'd64820, 16'd3342, 16'd51051, 16'd11155, 16'd53116, 16'd18227, 16'd32166, 16'd35327, 16'd55501, 16'd5258, 16'd54319, 16'd16040, 16'd16244, 16'd58887, 16'd26849});
	test_expansion(128'h92aeb7be49d84e88ddf6d8bad28b76b4, {16'd34164, 16'd20912, 16'd46590, 16'd24497, 16'd10412, 16'd57486, 16'd40916, 16'd12494, 16'd54409, 16'd15363, 16'd17599, 16'd45443, 16'd36569, 16'd28746, 16'd55696, 16'd31832, 16'd41865, 16'd65315, 16'd47848, 16'd59308, 16'd58917, 16'd56818, 16'd53417, 16'd54645, 16'd58972, 16'd18211});
	test_expansion(128'hb9db77f0ab36d8d8e84aa417d150de73, {16'd9375, 16'd28730, 16'd18736, 16'd4805, 16'd49872, 16'd52149, 16'd63817, 16'd50297, 16'd12887, 16'd35521, 16'd16305, 16'd27107, 16'd12825, 16'd30963, 16'd63249, 16'd52717, 16'd47991, 16'd23680, 16'd11916, 16'd45761, 16'd5377, 16'd32241, 16'd48656, 16'd23258, 16'd63113, 16'd16612});
	test_expansion(128'h403674561c5a09fbf0a90e2a194a030a, {16'd29516, 16'd58215, 16'd47139, 16'd29783, 16'd45211, 16'd19939, 16'd54044, 16'd41885, 16'd5862, 16'd62284, 16'd11420, 16'd12012, 16'd63110, 16'd1948, 16'd15332, 16'd30350, 16'd14557, 16'd58112, 16'd54546, 16'd55778, 16'd20304, 16'd8406, 16'd31583, 16'd49092, 16'd8855, 16'd26711});
	test_expansion(128'hc30c94a242a59db37519ed628e775667, {16'd18149, 16'd24642, 16'd51940, 16'd27063, 16'd1125, 16'd50402, 16'd30974, 16'd47753, 16'd11797, 16'd45458, 16'd60066, 16'd55643, 16'd24425, 16'd40643, 16'd55274, 16'd22006, 16'd34203, 16'd29725, 16'd47632, 16'd18583, 16'd64719, 16'd57433, 16'd25932, 16'd55916, 16'd60704, 16'd7286});
	test_expansion(128'h22a0807494f321baf4d2c60460f37714, {16'd18109, 16'd3422, 16'd1657, 16'd18012, 16'd17023, 16'd64491, 16'd27922, 16'd48628, 16'd3535, 16'd4663, 16'd35181, 16'd19796, 16'd60262, 16'd5713, 16'd289, 16'd20746, 16'd65301, 16'd23387, 16'd45411, 16'd62326, 16'd52930, 16'd10060, 16'd11353, 16'd23237, 16'd43846, 16'd28222});
	test_expansion(128'h7dfe205fbb8642175b18cf4fa25e782f, {16'd50487, 16'd27014, 16'd53258, 16'd25844, 16'd9346, 16'd32010, 16'd38541, 16'd54474, 16'd54682, 16'd25229, 16'd29695, 16'd44752, 16'd14834, 16'd54976, 16'd12607, 16'd1730, 16'd14217, 16'd65341, 16'd16122, 16'd45491, 16'd16724, 16'd19912, 16'd43646, 16'd15074, 16'd65516, 16'd50420});
	test_expansion(128'h931f508ebfc58859a7669acbe503b952, {16'd3014, 16'd28563, 16'd16180, 16'd22918, 16'd51767, 16'd6112, 16'd12383, 16'd38005, 16'd36756, 16'd63074, 16'd22144, 16'd63868, 16'd5700, 16'd40928, 16'd3135, 16'd25019, 16'd29125, 16'd35503, 16'd52796, 16'd39231, 16'd28902, 16'd53717, 16'd44264, 16'd8803, 16'd18385, 16'd20541});
	test_expansion(128'h8a013ce6cf38b98ba4f553b5f0a9a082, {16'd16247, 16'd49388, 16'd53107, 16'd12755, 16'd27856, 16'd49970, 16'd32470, 16'd35969, 16'd4917, 16'd42935, 16'd24344, 16'd35298, 16'd16961, 16'd41525, 16'd25592, 16'd58017, 16'd54241, 16'd22915, 16'd39135, 16'd17151, 16'd26603, 16'd15143, 16'd12849, 16'd6631, 16'd38527, 16'd44586});
	test_expansion(128'h1f7a032248f30ad390f9bad4463f6a62, {16'd23859, 16'd6746, 16'd39809, 16'd8514, 16'd25952, 16'd48645, 16'd11612, 16'd44978, 16'd12887, 16'd4901, 16'd27443, 16'd27636, 16'd40723, 16'd47270, 16'd5290, 16'd9435, 16'd59853, 16'd26630, 16'd50158, 16'd13109, 16'd21999, 16'd49517, 16'd54440, 16'd53763, 16'd32791, 16'd38568});
	test_expansion(128'h8bf17248c64ead5e08df4078ac130f43, {16'd38792, 16'd25105, 16'd2773, 16'd2883, 16'd46357, 16'd62298, 16'd57594, 16'd50265, 16'd59700, 16'd46141, 16'd36472, 16'd2141, 16'd61987, 16'd40475, 16'd30732, 16'd3070, 16'd17089, 16'd14041, 16'd43227, 16'd16497, 16'd37868, 16'd17079, 16'd21932, 16'd32844, 16'd5664, 16'd19023});
	test_expansion(128'h39d1db4a92c4ee159109e3770425d84b, {16'd47012, 16'd28795, 16'd49442, 16'd41539, 16'd58802, 16'd10167, 16'd24135, 16'd41312, 16'd12382, 16'd64414, 16'd5001, 16'd58783, 16'd35634, 16'd2539, 16'd4231, 16'd29190, 16'd56166, 16'd49994, 16'd23366, 16'd29230, 16'd31850, 16'd22095, 16'd12826, 16'd3666, 16'd3748, 16'd40084});
	test_expansion(128'h61faaa67e2e8aea455be1b998607d394, {16'd2442, 16'd10566, 16'd55889, 16'd26442, 16'd13713, 16'd30348, 16'd18353, 16'd44106, 16'd8357, 16'd31239, 16'd21576, 16'd61644, 16'd63988, 16'd46913, 16'd40148, 16'd52536, 16'd27265, 16'd61447, 16'd37575, 16'd60312, 16'd27781, 16'd19550, 16'd41619, 16'd64552, 16'd6570, 16'd61607});
	test_expansion(128'he96e12f5e3ca40320710f4748d91cf6f, {16'd51023, 16'd5298, 16'd2271, 16'd52187, 16'd41205, 16'd58424, 16'd48917, 16'd29289, 16'd25773, 16'd64800, 16'd17353, 16'd3711, 16'd14467, 16'd23524, 16'd46642, 16'd45037, 16'd596, 16'd17532, 16'd49485, 16'd34740, 16'd53873, 16'd1799, 16'd59465, 16'd39035, 16'd40234, 16'd40308});
	test_expansion(128'h936c53eea167f91e610ac0277b2e8aa2, {16'd836, 16'd25648, 16'd10078, 16'd25218, 16'd40565, 16'd11923, 16'd43653, 16'd63340, 16'd30705, 16'd28729, 16'd60770, 16'd5531, 16'd64886, 16'd56297, 16'd50570, 16'd45803, 16'd55834, 16'd35019, 16'd36794, 16'd61832, 16'd14273, 16'd49146, 16'd51976, 16'd2420, 16'd28726, 16'd55827});
	test_expansion(128'hfb07b810bdabcc541ae570a753d8625e, {16'd40048, 16'd1428, 16'd31052, 16'd64639, 16'd47681, 16'd16140, 16'd53261, 16'd50104, 16'd1315, 16'd20119, 16'd44850, 16'd34910, 16'd8166, 16'd49870, 16'd24082, 16'd17807, 16'd55342, 16'd28681, 16'd34071, 16'd53995, 16'd58056, 16'd34845, 16'd8077, 16'd3520, 16'd39745, 16'd1883});
	test_expansion(128'hc738266aba59a55c8f09a147fadcde51, {16'd16566, 16'd1160, 16'd6638, 16'd20517, 16'd25928, 16'd52258, 16'd59163, 16'd62989, 16'd6345, 16'd30976, 16'd29206, 16'd35586, 16'd4861, 16'd52028, 16'd36589, 16'd31160, 16'd9784, 16'd44379, 16'd11234, 16'd42859, 16'd12422, 16'd5644, 16'd49991, 16'd65388, 16'd45556, 16'd58344});
	test_expansion(128'h05c4b91c98d7fa08b7416299efb24bb6, {16'd20807, 16'd31463, 16'd14024, 16'd47405, 16'd46414, 16'd15241, 16'd29223, 16'd27365, 16'd20106, 16'd32566, 16'd19922, 16'd5797, 16'd15165, 16'd31560, 16'd44239, 16'd26228, 16'd37905, 16'd38852, 16'd61264, 16'd22679, 16'd33434, 16'd24110, 16'd49392, 16'd65235, 16'd39761, 16'd61459});
	test_expansion(128'h6713a4ca43b95873f597e8300f69d8d4, {16'd47318, 16'd56371, 16'd22898, 16'd10422, 16'd4447, 16'd62640, 16'd49144, 16'd37594, 16'd17587, 16'd29696, 16'd48487, 16'd30933, 16'd52220, 16'd24528, 16'd6196, 16'd47546, 16'd27188, 16'd34967, 16'd11197, 16'd1570, 16'd18416, 16'd12329, 16'd10453, 16'd7844, 16'd8529, 16'd30489});
	test_expansion(128'hcfc8b27956e47db145a983738b2f634f, {16'd60962, 16'd14233, 16'd34764, 16'd51387, 16'd22689, 16'd65522, 16'd60996, 16'd47582, 16'd39767, 16'd56355, 16'd62779, 16'd4088, 16'd43907, 16'd8055, 16'd25511, 16'd58206, 16'd52665, 16'd57245, 16'd39412, 16'd61726, 16'd49779, 16'd64604, 16'd8005, 16'd41924, 16'd19591, 16'd48863});
	test_expansion(128'hea8b864ee4c62e88692294d31413319c, {16'd3837, 16'd3741, 16'd564, 16'd35881, 16'd55505, 16'd47410, 16'd59410, 16'd64036, 16'd32054, 16'd36602, 16'd63034, 16'd15420, 16'd31690, 16'd40275, 16'd16702, 16'd34578, 16'd45388, 16'd21625, 16'd33686, 16'd4246, 16'd1420, 16'd45592, 16'd19314, 16'd11061, 16'd23447, 16'd64968});
	test_expansion(128'h23fd0e1c47cec46d5ba6be6eb2b27f1c, {16'd63217, 16'd32975, 16'd2758, 16'd27397, 16'd47184, 16'd65144, 16'd16733, 16'd65396, 16'd50702, 16'd64316, 16'd40709, 16'd39450, 16'd24768, 16'd58687, 16'd51875, 16'd43982, 16'd43, 16'd9462, 16'd11092, 16'd43342, 16'd19964, 16'd16146, 16'd33430, 16'd8494, 16'd16252, 16'd49572});
	test_expansion(128'h91f92dadaaf952f0a352352feaef392e, {16'd34285, 16'd22278, 16'd40027, 16'd7163, 16'd31208, 16'd20825, 16'd22098, 16'd1504, 16'd14323, 16'd31671, 16'd58175, 16'd47298, 16'd45660, 16'd49537, 16'd58143, 16'd43392, 16'd40691, 16'd57308, 16'd21089, 16'd29394, 16'd60857, 16'd28410, 16'd34221, 16'd30504, 16'd31868, 16'd57283});
	test_expansion(128'h8930769e7e724a2cb25564fee6b87ec3, {16'd17161, 16'd11637, 16'd47273, 16'd13872, 16'd44671, 16'd62558, 16'd33435, 16'd43964, 16'd3319, 16'd47104, 16'd56889, 16'd53756, 16'd21041, 16'd62970, 16'd13538, 16'd44584, 16'd41376, 16'd51634, 16'd33607, 16'd40891, 16'd28780, 16'd59016, 16'd25913, 16'd61562, 16'd57683, 16'd32557});
	test_expansion(128'ha16255d3d54386ebc86caef68f038df7, {16'd31576, 16'd36031, 16'd61971, 16'd58584, 16'd47968, 16'd43781, 16'd23521, 16'd20871, 16'd39461, 16'd22319, 16'd37361, 16'd43369, 16'd35038, 16'd46402, 16'd48513, 16'd60892, 16'd59976, 16'd41652, 16'd52355, 16'd58154, 16'd64798, 16'd41117, 16'd35821, 16'd8746, 16'd16101, 16'd33818});
	test_expansion(128'h4d08088b438e3f7453ad16830ef6a838, {16'd2373, 16'd28184, 16'd38473, 16'd37430, 16'd15814, 16'd8633, 16'd8563, 16'd59722, 16'd6082, 16'd10345, 16'd22030, 16'd65120, 16'd11763, 16'd29485, 16'd21251, 16'd42460, 16'd16733, 16'd34704, 16'd18012, 16'd25771, 16'd14442, 16'd30386, 16'd60421, 16'd37315, 16'd46097, 16'd55214});
	test_expansion(128'hb41a51b3eb856eb6b23c08c4cf6b8b80, {16'd50477, 16'd60894, 16'd28847, 16'd42244, 16'd35766, 16'd60997, 16'd25294, 16'd9479, 16'd37386, 16'd7369, 16'd52510, 16'd10885, 16'd21966, 16'd34009, 16'd46666, 16'd26196, 16'd32764, 16'd2612, 16'd53739, 16'd37486, 16'd4808, 16'd12328, 16'd60437, 16'd64367, 16'd37941, 16'd37120});
	test_expansion(128'hb4f7bb9a5cee0ad0ea08add01b282ddc, {16'd59584, 16'd50718, 16'd35031, 16'd63460, 16'd56908, 16'd31862, 16'd37320, 16'd49596, 16'd6864, 16'd32727, 16'd57240, 16'd51479, 16'd61088, 16'd47793, 16'd8664, 16'd64277, 16'd6313, 16'd29512, 16'd13830, 16'd7158, 16'd58150, 16'd8652, 16'd509, 16'd29703, 16'd59481, 16'd54467});
	test_expansion(128'he6048f15a5c6cf4a0c556d7fc32a8b04, {16'd22472, 16'd22244, 16'd60853, 16'd12897, 16'd27287, 16'd63937, 16'd48664, 16'd33281, 16'd1072, 16'd43144, 16'd11937, 16'd10326, 16'd18553, 16'd22811, 16'd34722, 16'd778, 16'd43013, 16'd24429, 16'd43559, 16'd8793, 16'd7528, 16'd27473, 16'd16968, 16'd35910, 16'd7784, 16'd14433});
	test_expansion(128'hf6a89e9d82fc144b4ce4e801b8419447, {16'd63542, 16'd19563, 16'd25347, 16'd52364, 16'd10565, 16'd35682, 16'd7528, 16'd8387, 16'd47512, 16'd29129, 16'd31229, 16'd46853, 16'd9856, 16'd15649, 16'd13321, 16'd44398, 16'd1744, 16'd14798, 16'd29754, 16'd25989, 16'd31546, 16'd16237, 16'd49620, 16'd51880, 16'd22623, 16'd44555});
	test_expansion(128'h37e38947ba6a797e8c6909dafff5e3f0, {16'd47342, 16'd3670, 16'd47215, 16'd43563, 16'd11981, 16'd36758, 16'd37059, 16'd64674, 16'd16564, 16'd24965, 16'd45709, 16'd64585, 16'd1697, 16'd62586, 16'd9073, 16'd59147, 16'd33284, 16'd1671, 16'd11466, 16'd19649, 16'd36086, 16'd48236, 16'd46369, 16'd54022, 16'd27113, 16'd65030});
	test_expansion(128'ha0c2a0e152df0d290c5bc1c82907dddf, {16'd41600, 16'd63268, 16'd50192, 16'd504, 16'd4692, 16'd65056, 16'd36301, 16'd17420, 16'd40956, 16'd45446, 16'd53604, 16'd37433, 16'd7987, 16'd37054, 16'd21305, 16'd2021, 16'd51887, 16'd686, 16'd10558, 16'd30867, 16'd16160, 16'd52154, 16'd19285, 16'd33018, 16'd31435, 16'd30157});
	test_expansion(128'h7dd667a993104f79fa5c09dcd0b5004c, {16'd44541, 16'd21158, 16'd27246, 16'd18909, 16'd23422, 16'd25253, 16'd5923, 16'd22185, 16'd54763, 16'd27088, 16'd54997, 16'd18977, 16'd50087, 16'd14873, 16'd27570, 16'd61461, 16'd30283, 16'd8460, 16'd2389, 16'd15228, 16'd36845, 16'd29243, 16'd16019, 16'd58143, 16'd64288, 16'd8072});
	test_expansion(128'h912504d299c92ea6f406969fefee9dd4, {16'd61787, 16'd5792, 16'd26739, 16'd39911, 16'd2012, 16'd35666, 16'd18845, 16'd23768, 16'd35859, 16'd43672, 16'd28488, 16'd5643, 16'd31482, 16'd6995, 16'd40615, 16'd44637, 16'd57968, 16'd19571, 16'd43357, 16'd34804, 16'd51685, 16'd55767, 16'd39794, 16'd56863, 16'd13345, 16'd18676});
	test_expansion(128'hb8c0c3b8d350a797d31f8daa3b35c1b0, {16'd16350, 16'd1596, 16'd24428, 16'd23080, 16'd20799, 16'd13739, 16'd18596, 16'd27662, 16'd63826, 16'd22357, 16'd31543, 16'd36879, 16'd18425, 16'd20030, 16'd54324, 16'd21671, 16'd55359, 16'd5474, 16'd37913, 16'd33464, 16'd30090, 16'd33502, 16'd26436, 16'd9763, 16'd62125, 16'd53146});
	test_expansion(128'heb873d5d8f5edca141605a94d5b1c558, {16'd50030, 16'd13649, 16'd62829, 16'd54105, 16'd32918, 16'd56799, 16'd56160, 16'd44856, 16'd19181, 16'd24382, 16'd16845, 16'd22230, 16'd53471, 16'd1462, 16'd48763, 16'd21693, 16'd26815, 16'd20109, 16'd41029, 16'd61915, 16'd16629, 16'd50510, 16'd25191, 16'd19577, 16'd44232, 16'd23767});
	test_expansion(128'hea1053a65936512f253848ec29d6d4dd, {16'd37798, 16'd62098, 16'd23876, 16'd59008, 16'd15569, 16'd52077, 16'd29321, 16'd59070, 16'd51998, 16'd50739, 16'd24378, 16'd45685, 16'd44344, 16'd17216, 16'd20733, 16'd52834, 16'd22125, 16'd64037, 16'd28563, 16'd49923, 16'd35930, 16'd13573, 16'd17538, 16'd43803, 16'd62043, 16'd61830});
	test_expansion(128'h08da64a09bb57054b294f42249a1dcd6, {16'd52082, 16'd37657, 16'd25223, 16'd57814, 16'd18770, 16'd32783, 16'd11353, 16'd18929, 16'd7973, 16'd27480, 16'd52741, 16'd55268, 16'd16717, 16'd59897, 16'd50758, 16'd5417, 16'd27302, 16'd3815, 16'd62694, 16'd10415, 16'd13928, 16'd53224, 16'd34311, 16'd32337, 16'd57522, 16'd58519});
	test_expansion(128'hf385762ac09c9f213ea3b3d060c32f8a, {16'd26183, 16'd64510, 16'd59254, 16'd32189, 16'd56614, 16'd30399, 16'd39011, 16'd30013, 16'd17000, 16'd5764, 16'd28662, 16'd61895, 16'd25734, 16'd10453, 16'd63149, 16'd771, 16'd8967, 16'd43191, 16'd46552, 16'd60223, 16'd13049, 16'd32091, 16'd21266, 16'd35103, 16'd62618, 16'd18980});
	test_expansion(128'h7ecb705e356615830c1720f71b072adf, {16'd6909, 16'd52357, 16'd60156, 16'd5240, 16'd42145, 16'd18698, 16'd43319, 16'd59189, 16'd13472, 16'd6620, 16'd54130, 16'd62437, 16'd38679, 16'd37870, 16'd64049, 16'd39657, 16'd57578, 16'd63697, 16'd56899, 16'd11280, 16'd33142, 16'd50376, 16'd3966, 16'd32671, 16'd46149, 16'd30581});
	test_expansion(128'h9b25016b66c530eca07735b43a4ff260, {16'd40107, 16'd34085, 16'd50914, 16'd62601, 16'd63790, 16'd3494, 16'd36201, 16'd20453, 16'd46347, 16'd25642, 16'd59109, 16'd50159, 16'd37249, 16'd25490, 16'd3800, 16'd9741, 16'd56572, 16'd53474, 16'd21661, 16'd31144, 16'd30522, 16'd18606, 16'd59294, 16'd38017, 16'd10071, 16'd63851});
	test_expansion(128'h876c5067c89c131288a04c39a0d4029a, {16'd36121, 16'd48361, 16'd6090, 16'd6427, 16'd49674, 16'd43929, 16'd12109, 16'd57427, 16'd65410, 16'd1081, 16'd1011, 16'd28040, 16'd1502, 16'd55025, 16'd3261, 16'd319, 16'd51086, 16'd3562, 16'd49806, 16'd14302, 16'd62819, 16'd630, 16'd19570, 16'd40033, 16'd10432, 16'd16115});
	test_expansion(128'heefd00fa075018adec6a8e2f45e61e3c, {16'd50456, 16'd22470, 16'd57712, 16'd9903, 16'd14666, 16'd62842, 16'd7588, 16'd4948, 16'd18763, 16'd48296, 16'd50993, 16'd29872, 16'd5142, 16'd7548, 16'd62241, 16'd2012, 16'd36657, 16'd63065, 16'd38863, 16'd47220, 16'd9986, 16'd38076, 16'd18427, 16'd40007, 16'd44136, 16'd46719});
	test_expansion(128'h448e4a9c3cd16dde772b10c4a4177437, {16'd8304, 16'd18715, 16'd25346, 16'd1806, 16'd43932, 16'd39230, 16'd37569, 16'd14323, 16'd54051, 16'd12321, 16'd46767, 16'd6519, 16'd4794, 16'd3516, 16'd41797, 16'd63041, 16'd32503, 16'd17683, 16'd23131, 16'd18711, 16'd64581, 16'd13656, 16'd30026, 16'd20743, 16'd16932, 16'd56921});
	test_expansion(128'h7b72671122328a15b528a10caa75f01a, {16'd21357, 16'd52736, 16'd16486, 16'd33705, 16'd53701, 16'd30805, 16'd35637, 16'd13769, 16'd47818, 16'd25703, 16'd21646, 16'd11610, 16'd25974, 16'd23047, 16'd22387, 16'd36368, 16'd4814, 16'd3786, 16'd21752, 16'd4665, 16'd45344, 16'd49384, 16'd52820, 16'd30514, 16'd62910, 16'd9376});
	test_expansion(128'hb21c222ae2154aa18aa0102141bb1cce, {16'd4691, 16'd12895, 16'd40057, 16'd8799, 16'd47873, 16'd45715, 16'd16421, 16'd59600, 16'd22246, 16'd24443, 16'd11097, 16'd41278, 16'd11410, 16'd51941, 16'd35021, 16'd59090, 16'd24983, 16'd48281, 16'd3604, 16'd43440, 16'd60269, 16'd44082, 16'd47126, 16'd48620, 16'd35294, 16'd26877});
	test_expansion(128'h61da8c21600dfebc8e7cf8c2d600f852, {16'd43583, 16'd15990, 16'd17645, 16'd16123, 16'd61306, 16'd43540, 16'd12317, 16'd3965, 16'd33136, 16'd33491, 16'd39120, 16'd5491, 16'd38100, 16'd37203, 16'd31685, 16'd45074, 16'd29915, 16'd13854, 16'd6105, 16'd56642, 16'd39764, 16'd27015, 16'd14395, 16'd4742, 16'd9237, 16'd26880});
	test_expansion(128'hd14ea04902a717f428c0905016d6afe6, {16'd17778, 16'd60657, 16'd26336, 16'd36327, 16'd18956, 16'd28236, 16'd12502, 16'd58979, 16'd8023, 16'd42476, 16'd60602, 16'd50087, 16'd44178, 16'd46176, 16'd11999, 16'd25803, 16'd38321, 16'd12153, 16'd22149, 16'd47490, 16'd54936, 16'd30603, 16'd56655, 16'd3791, 16'd21843, 16'd37289});
	test_expansion(128'hc63ba5b0c36ffd4ac3da4dc8870b201b, {16'd24022, 16'd19300, 16'd35575, 16'd58706, 16'd18400, 16'd20022, 16'd65335, 16'd1464, 16'd19051, 16'd40016, 16'd30321, 16'd52972, 16'd41304, 16'd6033, 16'd13525, 16'd40744, 16'd32360, 16'd12788, 16'd37120, 16'd58946, 16'd1919, 16'd26015, 16'd12527, 16'd58732, 16'd8230, 16'd6124});
	test_expansion(128'h2368ef8c79eadf2cb88b4673a2828e22, {16'd39367, 16'd35647, 16'd48980, 16'd54241, 16'd65140, 16'd34977, 16'd12361, 16'd47870, 16'd51670, 16'd23755, 16'd47130, 16'd56176, 16'd52627, 16'd12928, 16'd27364, 16'd22967, 16'd31857, 16'd55338, 16'd29797, 16'd31828, 16'd7171, 16'd27176, 16'd64994, 16'd32117, 16'd39668, 16'd56623});
	test_expansion(128'hf3ee3dd2c72fc3a8a5e0c00b1fa86fbe, {16'd7483, 16'd11947, 16'd52986, 16'd35218, 16'd31934, 16'd56031, 16'd59745, 16'd22753, 16'd4837, 16'd36598, 16'd3107, 16'd3480, 16'd50949, 16'd23552, 16'd5453, 16'd23223, 16'd48929, 16'd37969, 16'd4609, 16'd12384, 16'd9903, 16'd49283, 16'd46439, 16'd46795, 16'd10726, 16'd56709});
	test_expansion(128'h6e96bcfea897b112b5f7d0bda19ea716, {16'd49356, 16'd34983, 16'd41291, 16'd49657, 16'd37997, 16'd51353, 16'd44123, 16'd44747, 16'd64398, 16'd62081, 16'd44351, 16'd52508, 16'd46156, 16'd41749, 16'd18342, 16'd18260, 16'd59864, 16'd33114, 16'd3992, 16'd52102, 16'd22969, 16'd48861, 16'd40764, 16'd44041, 16'd10302, 16'd18743});
	test_expansion(128'h04e4cce86c4901d7be18f00d82d0bde5, {16'd38656, 16'd47657, 16'd55341, 16'd21128, 16'd4894, 16'd55105, 16'd51500, 16'd63447, 16'd6604, 16'd19331, 16'd49012, 16'd39482, 16'd65505, 16'd34368, 16'd49201, 16'd12419, 16'd33052, 16'd41855, 16'd63332, 16'd14046, 16'd6169, 16'd7647, 16'd37562, 16'd38123, 16'd6660, 16'd31195});
	test_expansion(128'h3377ebcbcc3b9d3328a5986f723e718c, {16'd34753, 16'd48356, 16'd17053, 16'd59842, 16'd55908, 16'd55570, 16'd2719, 16'd4984, 16'd54368, 16'd40272, 16'd44208, 16'd58020, 16'd51220, 16'd4137, 16'd48360, 16'd44687, 16'd55254, 16'd30262, 16'd7207, 16'd60683, 16'd22148, 16'd34995, 16'd38381, 16'd51480, 16'd19905, 16'd4251});
	test_expansion(128'hf936bf6eaccab481c3d77d879a6a1c35, {16'd9206, 16'd48622, 16'd59995, 16'd46580, 16'd27710, 16'd17697, 16'd37627, 16'd37890, 16'd9267, 16'd37811, 16'd58214, 16'd45512, 16'd55343, 16'd14649, 16'd61814, 16'd55150, 16'd24370, 16'd21019, 16'd37567, 16'd14836, 16'd27407, 16'd52770, 16'd30677, 16'd55726, 16'd61200, 16'd61633});
	test_expansion(128'hccec0d7357bd4d90fef87b86f31a681d, {16'd63259, 16'd31991, 16'd12394, 16'd31953, 16'd42817, 16'd54636, 16'd62300, 16'd59598, 16'd60695, 16'd21579, 16'd59220, 16'd38374, 16'd28686, 16'd4479, 16'd11343, 16'd45821, 16'd46120, 16'd24515, 16'd35482, 16'd15916, 16'd3666, 16'd53404, 16'd26662, 16'd60312, 16'd38867, 16'd15631});
	test_expansion(128'h3e57ed46ccfd6eb949c1a38f60375c8e, {16'd34724, 16'd55828, 16'd26644, 16'd18235, 16'd44263, 16'd38740, 16'd32932, 16'd4988, 16'd26763, 16'd46396, 16'd45151, 16'd61177, 16'd2385, 16'd15639, 16'd4394, 16'd26212, 16'd60927, 16'd9276, 16'd48760, 16'd16156, 16'd42136, 16'd55731, 16'd34438, 16'd33363, 16'd44674, 16'd19975});
	test_expansion(128'h6de552e0e109ef017c11219a0267375e, {16'd15544, 16'd13980, 16'd64264, 16'd12641, 16'd47868, 16'd32964, 16'd8443, 16'd47178, 16'd4725, 16'd12448, 16'd3302, 16'd61352, 16'd58000, 16'd29813, 16'd29609, 16'd54515, 16'd24829, 16'd29222, 16'd25063, 16'd62572, 16'd58676, 16'd34450, 16'd20959, 16'd23623, 16'd4592, 16'd38507});
	test_expansion(128'h4710000402b49a5693746078e2bcc1f5, {16'd21269, 16'd42115, 16'd37382, 16'd4959, 16'd28560, 16'd50045, 16'd1356, 16'd18103, 16'd47768, 16'd27698, 16'd13789, 16'd20738, 16'd14423, 16'd61340, 16'd27637, 16'd30146, 16'd20787, 16'd55988, 16'd47931, 16'd50235, 16'd10314, 16'd50189, 16'd34538, 16'd5976, 16'd2053, 16'd7587});
	test_expansion(128'h47f0b7b50ea6e69c0e15383aade5df83, {16'd41626, 16'd17961, 16'd24117, 16'd64111, 16'd37872, 16'd54706, 16'd3054, 16'd5135, 16'd3486, 16'd53369, 16'd25882, 16'd37605, 16'd64479, 16'd24933, 16'd9021, 16'd11486, 16'd48790, 16'd34907, 16'd39739, 16'd41571, 16'd65114, 16'd61954, 16'd50436, 16'd13917, 16'd44938, 16'd23500});
	test_expansion(128'h81eb5eebc85ad725acf12bf4010da9ed, {16'd61767, 16'd46250, 16'd60849, 16'd61544, 16'd33527, 16'd56669, 16'd59522, 16'd36126, 16'd27108, 16'd47499, 16'd10595, 16'd36699, 16'd56688, 16'd4830, 16'd42624, 16'd26755, 16'd39817, 16'd32542, 16'd38504, 16'd35116, 16'd28904, 16'd22463, 16'd39907, 16'd2618, 16'd50384, 16'd44550});
	test_expansion(128'h69fa72f0d34a85c21cc83cd760d2fbec, {16'd56388, 16'd64505, 16'd21798, 16'd33765, 16'd55311, 16'd57619, 16'd33244, 16'd20036, 16'd31872, 16'd62769, 16'd56768, 16'd59181, 16'd63530, 16'd35997, 16'd30304, 16'd28196, 16'd51075, 16'd53176, 16'd15921, 16'd33436, 16'd29680, 16'd46602, 16'd8149, 16'd55308, 16'd13654, 16'd26033});
	test_expansion(128'h9b0b9f72383013dd8166c7d9b5c80fca, {16'd47272, 16'd50122, 16'd5002, 16'd23076, 16'd33762, 16'd62896, 16'd30002, 16'd320, 16'd29947, 16'd34860, 16'd39927, 16'd37161, 16'd11456, 16'd53951, 16'd61226, 16'd48266, 16'd45021, 16'd33264, 16'd51195, 16'd45417, 16'd47009, 16'd13535, 16'd29306, 16'd49386, 16'd34374, 16'd2902});
	test_expansion(128'h014a5154ccf50b73d52b5daf5a4ed831, {16'd24172, 16'd42139, 16'd3647, 16'd8809, 16'd52839, 16'd33133, 16'd52717, 16'd20997, 16'd56137, 16'd15007, 16'd28947, 16'd28818, 16'd46201, 16'd51758, 16'd5808, 16'd22167, 16'd6375, 16'd32315, 16'd58404, 16'd46725, 16'd2784, 16'd46320, 16'd42847, 16'd43812, 16'd12890, 16'd55442});
	test_expansion(128'h7e37bbab730d9352a31ac360efbb4044, {16'd29940, 16'd8210, 16'd3488, 16'd58849, 16'd2963, 16'd53703, 16'd39080, 16'd365, 16'd31273, 16'd17144, 16'd53051, 16'd59612, 16'd36510, 16'd30403, 16'd7052, 16'd46316, 16'd25903, 16'd32566, 16'd22009, 16'd58825, 16'd555, 16'd51073, 16'd36530, 16'd12143, 16'd10584, 16'd26583});
	test_expansion(128'hfe03e172c7cafb2eb04916715147c83a, {16'd47461, 16'd18612, 16'd21880, 16'd5740, 16'd57401, 16'd15418, 16'd50616, 16'd13173, 16'd46148, 16'd63310, 16'd15242, 16'd14776, 16'd41309, 16'd16723, 16'd20701, 16'd39393, 16'd64815, 16'd61277, 16'd51573, 16'd28031, 16'd30492, 16'd17395, 16'd22820, 16'd32931, 16'd42161, 16'd2592});
	test_expansion(128'h866efa8d4fd08feeaf4f1872ef38e7d0, {16'd61602, 16'd63722, 16'd14429, 16'd16421, 16'd64711, 16'd56230, 16'd44448, 16'd53934, 16'd16445, 16'd36439, 16'd54169, 16'd35143, 16'd55848, 16'd29324, 16'd54574, 16'd39786, 16'd33165, 16'd27255, 16'd45477, 16'd25190, 16'd38688, 16'd21018, 16'd16453, 16'd5262, 16'd57953, 16'd21242});
	test_expansion(128'h2f9a1b76eba0880d17284ab6a2d87fca, {16'd12937, 16'd12219, 16'd15905, 16'd23761, 16'd25090, 16'd39890, 16'd35640, 16'd49954, 16'd20181, 16'd18825, 16'd18040, 16'd55260, 16'd64709, 16'd30361, 16'd28348, 16'd16758, 16'd11527, 16'd17343, 16'd5207, 16'd48789, 16'd28477, 16'd11692, 16'd18676, 16'd5888, 16'd45226, 16'd19795});
	test_expansion(128'hc0b02c218533f5330a125dda4120c232, {16'd44322, 16'd65011, 16'd46948, 16'd16906, 16'd57359, 16'd46399, 16'd64180, 16'd5953, 16'd14782, 16'd30327, 16'd6046, 16'd838, 16'd45583, 16'd47755, 16'd16275, 16'd51100, 16'd13842, 16'd49274, 16'd36486, 16'd63155, 16'd55365, 16'd61620, 16'd15007, 16'd51073, 16'd17588, 16'd44865});
	test_expansion(128'h666130e4dfe068ed6891394006907a36, {16'd37164, 16'd29936, 16'd38965, 16'd2344, 16'd29577, 16'd20492, 16'd27133, 16'd55144, 16'd56920, 16'd327, 16'd31623, 16'd47872, 16'd27967, 16'd33481, 16'd43127, 16'd30249, 16'd2697, 16'd16588, 16'd32475, 16'd42786, 16'd65420, 16'd49281, 16'd38246, 16'd58867, 16'd61961, 16'd2007});
	test_expansion(128'h168b81b0e58881551056ceffa0cafe30, {16'd17835, 16'd14286, 16'd14741, 16'd29124, 16'd27678, 16'd15985, 16'd16530, 16'd18737, 16'd19835, 16'd18725, 16'd13423, 16'd44016, 16'd31489, 16'd50493, 16'd39344, 16'd57103, 16'd2377, 16'd9908, 16'd41262, 16'd48689, 16'd28834, 16'd25990, 16'd33608, 16'd6212, 16'd39427, 16'd879});
	test_expansion(128'h578f447a65fc5819d9e4941604a8e6e9, {16'd31734, 16'd23405, 16'd15186, 16'd49095, 16'd32432, 16'd31205, 16'd63560, 16'd17252, 16'd60005, 16'd64206, 16'd22858, 16'd4899, 16'd47976, 16'd62085, 16'd56546, 16'd52342, 16'd33281, 16'd19516, 16'd51696, 16'd16835, 16'd65337, 16'd27481, 16'd1074, 16'd33068, 16'd54005, 16'd11586});
	test_expansion(128'h0bf3c308ddb50edf35b63009cc0ae9dd, {16'd8400, 16'd56745, 16'd36903, 16'd35373, 16'd8341, 16'd33923, 16'd16473, 16'd33852, 16'd21883, 16'd48379, 16'd57581, 16'd27960, 16'd23352, 16'd37429, 16'd58570, 16'd43012, 16'd63800, 16'd52246, 16'd24346, 16'd38831, 16'd39881, 16'd30181, 16'd26672, 16'd41328, 16'd59768, 16'd50545});
	test_expansion(128'h69ac81b17b42ef9f6e5f7c78731eb3fb, {16'd58346, 16'd22366, 16'd13298, 16'd14119, 16'd50399, 16'd46077, 16'd53882, 16'd33967, 16'd1757, 16'd34600, 16'd14423, 16'd37475, 16'd20168, 16'd11259, 16'd57448, 16'd58487, 16'd42053, 16'd14732, 16'd7968, 16'd57643, 16'd51202, 16'd20414, 16'd30070, 16'd22626, 16'd2529, 16'd12312});
	test_expansion(128'h986b50c8e564e6a68ae61eb3f096ae0a, {16'd61004, 16'd22006, 16'd24613, 16'd49843, 16'd23096, 16'd39483, 16'd8364, 16'd23442, 16'd64952, 16'd18222, 16'd40512, 16'd61608, 16'd23558, 16'd46276, 16'd42804, 16'd17830, 16'd13521, 16'd27447, 16'd58030, 16'd7663, 16'd11518, 16'd53925, 16'd42730, 16'd19008, 16'd1564, 16'd55627});
	test_expansion(128'hd49a4a2491d282567d206c6e3568643f, {16'd29804, 16'd15165, 16'd10964, 16'd46179, 16'd12134, 16'd56054, 16'd33950, 16'd40834, 16'd53654, 16'd40760, 16'd31062, 16'd53083, 16'd47245, 16'd1281, 16'd58114, 16'd37514, 16'd61570, 16'd17152, 16'd48808, 16'd58035, 16'd28905, 16'd5409, 16'd2961, 16'd21781, 16'd54153, 16'd30342});
	test_expansion(128'hc9260ed066e8fe3562969b0ba0b159c2, {16'd47827, 16'd57917, 16'd55020, 16'd27452, 16'd2605, 16'd6318, 16'd3946, 16'd27880, 16'd6593, 16'd10285, 16'd50664, 16'd60838, 16'd4767, 16'd40899, 16'd45756, 16'd31820, 16'd49989, 16'd46075, 16'd55087, 16'd39284, 16'd17728, 16'd43622, 16'd23076, 16'd37397, 16'd32783, 16'd6294});
	test_expansion(128'h09b6d47d2ea769f4cfdb8e5cab913b32, {16'd24211, 16'd10977, 16'd18024, 16'd32688, 16'd6078, 16'd37358, 16'd18787, 16'd49629, 16'd11358, 16'd39697, 16'd23882, 16'd29484, 16'd62251, 16'd59769, 16'd56623, 16'd57593, 16'd28023, 16'd28124, 16'd34004, 16'd10211, 16'd37355, 16'd26519, 16'd36794, 16'd25751, 16'd16866, 16'd4265});
	test_expansion(128'hdcbf7fe2e18f5613bf2610649c5abaa2, {16'd32605, 16'd17812, 16'd27505, 16'd24380, 16'd2797, 16'd3764, 16'd26045, 16'd62187, 16'd47678, 16'd58852, 16'd14435, 16'd65374, 16'd12128, 16'd28415, 16'd63304, 16'd8207, 16'd19291, 16'd31724, 16'd45465, 16'd4652, 16'd21409, 16'd37563, 16'd49576, 16'd64631, 16'd56640, 16'd62966});
	test_expansion(128'hfa500fd76da3e6aa38bea90f0de536ff, {16'd10717, 16'd17281, 16'd63564, 16'd9078, 16'd45320, 16'd34720, 16'd54881, 16'd36001, 16'd18796, 16'd25350, 16'd15105, 16'd60451, 16'd23069, 16'd5437, 16'd62956, 16'd17331, 16'd48956, 16'd21432, 16'd2556, 16'd63217, 16'd29894, 16'd33041, 16'd33839, 16'd26734, 16'd59298, 16'd17015});
	test_expansion(128'h8a991609f42fc76d957e608d9fe3dc7a, {16'd1976, 16'd52008, 16'd11514, 16'd47597, 16'd27104, 16'd39598, 16'd26104, 16'd29001, 16'd10595, 16'd57916, 16'd65199, 16'd27219, 16'd42016, 16'd15824, 16'd36798, 16'd64512, 16'd18353, 16'd56478, 16'd39416, 16'd22026, 16'd54265, 16'd56990, 16'd61506, 16'd57857, 16'd9986, 16'd39834});
	test_expansion(128'h521650b92ca0acde7454ac7032c1d170, {16'd13789, 16'd63828, 16'd25398, 16'd3543, 16'd50411, 16'd18825, 16'd31683, 16'd19771, 16'd11750, 16'd52641, 16'd21928, 16'd15260, 16'd54233, 16'd29103, 16'd60308, 16'd7335, 16'd18563, 16'd57197, 16'd47844, 16'd31663, 16'd61211, 16'd26823, 16'd54257, 16'd52135, 16'd36218, 16'd36729});
	test_expansion(128'hf02e9f2c17caea123a2e11a96cd445bc, {16'd53906, 16'd65474, 16'd16572, 16'd3921, 16'd44148, 16'd20985, 16'd59544, 16'd6656, 16'd13257, 16'd24180, 16'd13424, 16'd14269, 16'd59604, 16'd48364, 16'd11674, 16'd22609, 16'd14493, 16'd62944, 16'd32608, 16'd30249, 16'd52890, 16'd7973, 16'd42896, 16'd65138, 16'd53449, 16'd35898});
	test_expansion(128'h3204046e80051e0fc26243e9d5a84d8a, {16'd58093, 16'd59181, 16'd63531, 16'd27626, 16'd26250, 16'd24585, 16'd33738, 16'd43941, 16'd25682, 16'd57184, 16'd49761, 16'd63905, 16'd9394, 16'd176, 16'd27612, 16'd65284, 16'd14949, 16'd26585, 16'd51689, 16'd43730, 16'd7443, 16'd53436, 16'd30742, 16'd20152, 16'd2221, 16'd26607});
	test_expansion(128'h3ac1734c2d5e7427ed0c6471a8b40256, {16'd45416, 16'd11935, 16'd62501, 16'd30420, 16'd42007, 16'd6562, 16'd4946, 16'd4104, 16'd55738, 16'd18038, 16'd41506, 16'd25909, 16'd27034, 16'd53051, 16'd28995, 16'd33480, 16'd20600, 16'd26328, 16'd59660, 16'd34740, 16'd52622, 16'd9946, 16'd52864, 16'd998, 16'd33971, 16'd37720});
	test_expansion(128'h19dc99b698b01f02dfb99064941b9bd3, {16'd10971, 16'd26482, 16'd25578, 16'd21243, 16'd54246, 16'd64874, 16'd36720, 16'd26949, 16'd17445, 16'd30404, 16'd22356, 16'd26234, 16'd54723, 16'd19842, 16'd14123, 16'd65203, 16'd62908, 16'd27025, 16'd10745, 16'd40849, 16'd10536, 16'd45169, 16'd9987, 16'd50351, 16'd14673, 16'd9775});
	test_expansion(128'heb8578ca0d4b52e259e70089111661ad, {16'd36101, 16'd51229, 16'd22782, 16'd39640, 16'd28712, 16'd41438, 16'd14259, 16'd36859, 16'd38360, 16'd37045, 16'd50491, 16'd44434, 16'd13375, 16'd62792, 16'd14692, 16'd15226, 16'd44032, 16'd12223, 16'd14090, 16'd28718, 16'd55989, 16'd4457, 16'd29562, 16'd44028, 16'd57582, 16'd21961});
	test_expansion(128'ha128a8945982838351828dc59c7b0e99, {16'd51317, 16'd7214, 16'd27051, 16'd26568, 16'd57097, 16'd51522, 16'd36455, 16'd59601, 16'd20239, 16'd36584, 16'd58050, 16'd26716, 16'd12533, 16'd33423, 16'd17900, 16'd38948, 16'd64002, 16'd34619, 16'd37388, 16'd31517, 16'd29896, 16'd37648, 16'd23224, 16'd5261, 16'd7866, 16'd58369});
	test_expansion(128'h0a696cc32403a4f6753e4639562b39f6, {16'd15972, 16'd30140, 16'd36105, 16'd46434, 16'd30807, 16'd17059, 16'd22267, 16'd39125, 16'd47714, 16'd16567, 16'd63644, 16'd27421, 16'd2060, 16'd14365, 16'd54714, 16'd27829, 16'd58672, 16'd2461, 16'd51334, 16'd46424, 16'd32032, 16'd34377, 16'd3336, 16'd40816, 16'd1064, 16'd33933});
	test_expansion(128'hcd2b80f8cbd9bd5851e47bf34ac3160c, {16'd54241, 16'd60144, 16'd63451, 16'd57218, 16'd1412, 16'd53573, 16'd47503, 16'd61019, 16'd7667, 16'd53176, 16'd16407, 16'd60509, 16'd26801, 16'd23642, 16'd24008, 16'd2028, 16'd65339, 16'd736, 16'd8338, 16'd480, 16'd34948, 16'd48042, 16'd38047, 16'd39065, 16'd58525, 16'd39981});
	test_expansion(128'ha4915c78c9ef9ecdbeb70db8bd28b055, {16'd5803, 16'd56427, 16'd9884, 16'd17530, 16'd9237, 16'd21033, 16'd28902, 16'd57542, 16'd54314, 16'd1474, 16'd38536, 16'd37245, 16'd9690, 16'd33003, 16'd56908, 16'd30675, 16'd52013, 16'd62429, 16'd40914, 16'd20986, 16'd51413, 16'd63024, 16'd56280, 16'd423, 16'd6366, 16'd51001});
	test_expansion(128'h55133eda59a3b8af282090911de6f6a3, {16'd58265, 16'd55560, 16'd29569, 16'd47889, 16'd63142, 16'd47016, 16'd27768, 16'd20200, 16'd34504, 16'd19477, 16'd40125, 16'd37680, 16'd43372, 16'd33705, 16'd30607, 16'd44219, 16'd11096, 16'd57757, 16'd5957, 16'd17740, 16'd32837, 16'd31667, 16'd49269, 16'd36103, 16'd6966, 16'd10275});
	test_expansion(128'h12b212ae21e77572a9441620023c6c1f, {16'd32314, 16'd61363, 16'd61485, 16'd25722, 16'd19625, 16'd61768, 16'd26263, 16'd47738, 16'd44286, 16'd36021, 16'd46885, 16'd36078, 16'd17488, 16'd28399, 16'd41359, 16'd62227, 16'd11704, 16'd48151, 16'd30490, 16'd65480, 16'd41419, 16'd63498, 16'd47769, 16'd49712, 16'd43327, 16'd16578});
	test_expansion(128'h052d41556ca10bc5c6a7cdee50f15602, {16'd33319, 16'd13555, 16'd20054, 16'd15487, 16'd1998, 16'd15178, 16'd26458, 16'd7982, 16'd44410, 16'd46853, 16'd55764, 16'd9034, 16'd38503, 16'd31892, 16'd20295, 16'd28013, 16'd51430, 16'd247, 16'd48257, 16'd29664, 16'd9654, 16'd64460, 16'd62676, 16'd38024, 16'd54110, 16'd59935});
	test_expansion(128'hdc5ffbf871a2f32c20344210add13227, {16'd62810, 16'd41314, 16'd38338, 16'd8424, 16'd22909, 16'd41903, 16'd56126, 16'd39640, 16'd61508, 16'd44196, 16'd29023, 16'd22299, 16'd2927, 16'd28919, 16'd60685, 16'd23702, 16'd1267, 16'd35727, 16'd11295, 16'd8892, 16'd2596, 16'd58576, 16'd30886, 16'd23228, 16'd12880, 16'd3568});
	test_expansion(128'hb5da4a8e4825af09934f7b8c716cea64, {16'd47604, 16'd61002, 16'd18357, 16'd36991, 16'd2823, 16'd34808, 16'd23203, 16'd25204, 16'd16283, 16'd30467, 16'd21504, 16'd64939, 16'd3842, 16'd25032, 16'd40030, 16'd47322, 16'd18572, 16'd31378, 16'd11912, 16'd34024, 16'd11566, 16'd17104, 16'd27154, 16'd56851, 16'd50783, 16'd2396});
	test_expansion(128'he5f497583ed7c594fd18c3b77b0f1493, {16'd18978, 16'd8870, 16'd21666, 16'd31057, 16'd52112, 16'd11703, 16'd61214, 16'd46371, 16'd59524, 16'd57106, 16'd54398, 16'd41036, 16'd40141, 16'd25177, 16'd40349, 16'd7083, 16'd29017, 16'd46816, 16'd55197, 16'd48804, 16'd9496, 16'd11021, 16'd41166, 16'd37932, 16'd44666, 16'd42870});
	test_expansion(128'he62756d27939a475b89e1ba668b3cba6, {16'd38387, 16'd2178, 16'd34525, 16'd20161, 16'd41979, 16'd25377, 16'd22064, 16'd138, 16'd36506, 16'd1012, 16'd42089, 16'd46031, 16'd55784, 16'd36052, 16'd27037, 16'd8403, 16'd11454, 16'd58174, 16'd37219, 16'd36056, 16'd34832, 16'd35050, 16'd30289, 16'd50932, 16'd4449, 16'd47417});
	test_expansion(128'hab58aeb5475f2815279ff28a9917a653, {16'd57920, 16'd32996, 16'd15817, 16'd59526, 16'd23543, 16'd14662, 16'd25575, 16'd14019, 16'd24427, 16'd45845, 16'd36779, 16'd43205, 16'd41700, 16'd23402, 16'd58255, 16'd35516, 16'd24092, 16'd11439, 16'd266, 16'd24137, 16'd43952, 16'd40850, 16'd7524, 16'd19597, 16'd31288, 16'd44355});
	test_expansion(128'h181739568a809998f85e31f2313241cf, {16'd48813, 16'd27114, 16'd11312, 16'd17763, 16'd16502, 16'd3490, 16'd55212, 16'd18269, 16'd41595, 16'd29992, 16'd60015, 16'd20024, 16'd32195, 16'd49408, 16'd43927, 16'd30765, 16'd11396, 16'd47428, 16'd17062, 16'd2399, 16'd57095, 16'd48989, 16'd37046, 16'd54760, 16'd48425, 16'd62522});
	test_expansion(128'hf28656cb57824c0e9825b2c41605198f, {16'd33787, 16'd52931, 16'd34273, 16'd10951, 16'd52349, 16'd25544, 16'd16133, 16'd50152, 16'd458, 16'd28743, 16'd7875, 16'd35350, 16'd50857, 16'd23123, 16'd24565, 16'd12236, 16'd46135, 16'd53419, 16'd58890, 16'd20172, 16'd61386, 16'd3303, 16'd20796, 16'd33022, 16'd36034, 16'd60406});
	test_expansion(128'h447cecc34af0c616c1008007dcea27bb, {16'd22666, 16'd45940, 16'd65237, 16'd54365, 16'd9020, 16'd43240, 16'd54215, 16'd58277, 16'd27076, 16'd37368, 16'd25360, 16'd64440, 16'd46215, 16'd46597, 16'd12233, 16'd32201, 16'd51757, 16'd13138, 16'd54199, 16'd17291, 16'd47215, 16'd21042, 16'd19779, 16'd35181, 16'd40079, 16'd59693});
	test_expansion(128'hf991bdf936beb9f9feb69cd7c6eae903, {16'd46456, 16'd39155, 16'd6619, 16'd166, 16'd46804, 16'd56816, 16'd35671, 16'd9519, 16'd47121, 16'd31373, 16'd63429, 16'd32322, 16'd30278, 16'd11671, 16'd3517, 16'd27308, 16'd1036, 16'd25229, 16'd41332, 16'd29359, 16'd55741, 16'd27657, 16'd26163, 16'd33125, 16'd34293, 16'd52711});
	test_expansion(128'h52588c3b6f7618dec59028e851fa7ec3, {16'd7189, 16'd17320, 16'd55526, 16'd7653, 16'd33281, 16'd26759, 16'd15185, 16'd46722, 16'd47750, 16'd38992, 16'd50897, 16'd51603, 16'd40578, 16'd52589, 16'd27927, 16'd41430, 16'd20006, 16'd50732, 16'd31724, 16'd15146, 16'd59887, 16'd11947, 16'd48630, 16'd56630, 16'd60505, 16'd10553});
	test_expansion(128'hb38f455259c4e6c4145d7791247c0d39, {16'd32508, 16'd65141, 16'd63581, 16'd13661, 16'd36587, 16'd29747, 16'd12403, 16'd39323, 16'd30495, 16'd41551, 16'd11771, 16'd5958, 16'd52493, 16'd56593, 16'd28179, 16'd46627, 16'd64035, 16'd58922, 16'd26854, 16'd55512, 16'd55921, 16'd5017, 16'd7028, 16'd49882, 16'd3237, 16'd51326});
	test_expansion(128'hda39bdc54e53a91deccf29abdf9e1a65, {16'd59859, 16'd62447, 16'd11069, 16'd8169, 16'd48349, 16'd26567, 16'd32848, 16'd3888, 16'd8224, 16'd60732, 16'd192, 16'd32045, 16'd27648, 16'd42205, 16'd13974, 16'd28534, 16'd57418, 16'd58780, 16'd6819, 16'd24397, 16'd33321, 16'd55688, 16'd32745, 16'd5254, 16'd38493, 16'd42695});
	test_expansion(128'h9f34b542393f456ad5cd1d2b0b9c75ee, {16'd15398, 16'd31191, 16'd32865, 16'd44719, 16'd5030, 16'd49179, 16'd29229, 16'd20218, 16'd53959, 16'd60629, 16'd2344, 16'd58854, 16'd38000, 16'd26558, 16'd61439, 16'd44052, 16'd52758, 16'd2402, 16'd39847, 16'd8904, 16'd25172, 16'd7891, 16'd42059, 16'd33072, 16'd15118, 16'd3117});
	test_expansion(128'ha31a3c3238142d4900808dc4f62aaf3c, {16'd26179, 16'd46189, 16'd56282, 16'd44749, 16'd36669, 16'd29390, 16'd33144, 16'd57309, 16'd18902, 16'd33650, 16'd64360, 16'd9261, 16'd64797, 16'd62691, 16'd31208, 16'd25982, 16'd1179, 16'd42310, 16'd31269, 16'd23970, 16'd7743, 16'd61745, 16'd29329, 16'd50179, 16'd2735, 16'd58085});
	test_expansion(128'hbb004dfa42caa515d9613c3196ead413, {16'd57240, 16'd52857, 16'd54773, 16'd7252, 16'd35557, 16'd33844, 16'd34753, 16'd1252, 16'd17256, 16'd22296, 16'd25034, 16'd9304, 16'd37464, 16'd21218, 16'd38748, 16'd18713, 16'd52821, 16'd21573, 16'd32474, 16'd3921, 16'd2879, 16'd58586, 16'd65178, 16'd943, 16'd24269, 16'd61922});
	test_expansion(128'hf61b68c7f2c72b96216ff4e3f1b613be, {16'd59689, 16'd54885, 16'd12984, 16'd4559, 16'd41360, 16'd65375, 16'd55359, 16'd37277, 16'd17338, 16'd43984, 16'd18682, 16'd17849, 16'd5038, 16'd17078, 16'd39515, 16'd12402, 16'd57569, 16'd24297, 16'd26860, 16'd47307, 16'd3753, 16'd64585, 16'd27543, 16'd37408, 16'd40509, 16'd39070});
	test_expansion(128'h6c0b0be1d855797e8b65ef5b22175524, {16'd52889, 16'd49682, 16'd193, 16'd56853, 16'd61318, 16'd64974, 16'd41372, 16'd3499, 16'd63601, 16'd35677, 16'd58913, 16'd48723, 16'd25073, 16'd19962, 16'd45104, 16'd43341, 16'd15286, 16'd25525, 16'd47480, 16'd33119, 16'd26357, 16'd33858, 16'd51332, 16'd13960, 16'd6850, 16'd21333});
	test_expansion(128'h12c8adb63e048a866822f01334f54cfe, {16'd44732, 16'd61919, 16'd15085, 16'd25192, 16'd61551, 16'd33021, 16'd6730, 16'd54149, 16'd11041, 16'd43249, 16'd26241, 16'd26250, 16'd51104, 16'd27397, 16'd25155, 16'd21163, 16'd16255, 16'd25628, 16'd41028, 16'd55216, 16'd51444, 16'd38014, 16'd24488, 16'd51128, 16'd434, 16'd18542});
	test_expansion(128'h78985561580e3d3a322cead7cf9225d0, {16'd45112, 16'd63187, 16'd55669, 16'd19521, 16'd18962, 16'd57940, 16'd13247, 16'd15361, 16'd59062, 16'd65029, 16'd18101, 16'd5917, 16'd54423, 16'd15725, 16'd47315, 16'd9607, 16'd29505, 16'd28369, 16'd27617, 16'd10418, 16'd37866, 16'd25646, 16'd31071, 16'd45420, 16'd15780, 16'd6649});
	test_expansion(128'h7f78d299413598b41b68b5c901a21ab2, {16'd53745, 16'd11441, 16'd20201, 16'd29652, 16'd12011, 16'd35307, 16'd20447, 16'd20980, 16'd10815, 16'd26201, 16'd64636, 16'd21444, 16'd28455, 16'd3210, 16'd1339, 16'd51214, 16'd52710, 16'd58182, 16'd32022, 16'd57987, 16'd24248, 16'd24189, 16'd42212, 16'd18127, 16'd37664, 16'd51047});
	test_expansion(128'hd863fdc4c8553b4341514d7fdbc84c25, {16'd48538, 16'd25850, 16'd30000, 16'd60863, 16'd35130, 16'd6154, 16'd15169, 16'd13391, 16'd24708, 16'd44474, 16'd40442, 16'd27874, 16'd63957, 16'd5041, 16'd57886, 16'd64529, 16'd23429, 16'd41202, 16'd28696, 16'd14802, 16'd28838, 16'd26794, 16'd10870, 16'd19851, 16'd39361, 16'd26216});
	test_expansion(128'h83209eefff0c26ed67a8b17678952388, {16'd48814, 16'd50718, 16'd19707, 16'd36258, 16'd2871, 16'd32200, 16'd25540, 16'd44454, 16'd48187, 16'd26047, 16'd63298, 16'd64536, 16'd25704, 16'd17276, 16'd14259, 16'd13967, 16'd28778, 16'd39436, 16'd26563, 16'd45559, 16'd12027, 16'd4953, 16'd9429, 16'd46033, 16'd26819, 16'd59});
	test_expansion(128'ha174104a02558de60fbaeb333c4ec7e7, {16'd34628, 16'd1829, 16'd30650, 16'd7373, 16'd18462, 16'd27511, 16'd9260, 16'd50099, 16'd10774, 16'd4090, 16'd2894, 16'd36626, 16'd61429, 16'd45291, 16'd18040, 16'd35646, 16'd55541, 16'd23016, 16'd14981, 16'd44023, 16'd42253, 16'd10291, 16'd34962, 16'd6097, 16'd15853, 16'd19765});
	test_expansion(128'h755d66816273fb3f9cb2da17c6fbe6a4, {16'd44092, 16'd61880, 16'd44456, 16'd1272, 16'd45291, 16'd29712, 16'd24401, 16'd44408, 16'd24109, 16'd44497, 16'd3107, 16'd16386, 16'd31887, 16'd55066, 16'd33218, 16'd4513, 16'd63427, 16'd40354, 16'd18498, 16'd43656, 16'd29634, 16'd39325, 16'd24950, 16'd41840, 16'd36274, 16'd14540});
	test_expansion(128'h8b166546665f7da1edd8bd831986dcdf, {16'd41014, 16'd30365, 16'd8851, 16'd33023, 16'd27134, 16'd18176, 16'd63801, 16'd59872, 16'd4109, 16'd7832, 16'd10655, 16'd58708, 16'd14854, 16'd39891, 16'd1944, 16'd41898, 16'd8917, 16'd50233, 16'd59220, 16'd20590, 16'd57467, 16'd56774, 16'd17417, 16'd22951, 16'd29130, 16'd23730});
	test_expansion(128'h31ce19c92e8f2ec72a70c2741842efc2, {16'd47102, 16'd34468, 16'd49318, 16'd52143, 16'd1813, 16'd34185, 16'd32996, 16'd14859, 16'd19735, 16'd54401, 16'd49344, 16'd18746, 16'd14533, 16'd27817, 16'd19697, 16'd48789, 16'd34429, 16'd16794, 16'd8970, 16'd61507, 16'd40382, 16'd58672, 16'd1190, 16'd10279, 16'd25810, 16'd54278});
	test_expansion(128'h9fccc03b59fc674c9d040531d0dbd14c, {16'd24446, 16'd37090, 16'd32241, 16'd19715, 16'd60275, 16'd32230, 16'd10750, 16'd6940, 16'd6201, 16'd3682, 16'd44010, 16'd59516, 16'd22443, 16'd53915, 16'd45576, 16'd20251, 16'd36164, 16'd38030, 16'd2193, 16'd42120, 16'd41699, 16'd15658, 16'd58995, 16'd9017, 16'd39241, 16'd1779});
	test_expansion(128'h69f14e314e1ccfda35ec9888c6525032, {16'd25187, 16'd26344, 16'd59987, 16'd12936, 16'd23940, 16'd34595, 16'd40558, 16'd40369, 16'd15648, 16'd21887, 16'd42134, 16'd38339, 16'd56636, 16'd25695, 16'd14101, 16'd20140, 16'd14597, 16'd19530, 16'd40643, 16'd34387, 16'd57386, 16'd47855, 16'd55124, 16'd16511, 16'd6965, 16'd15798});
	test_expansion(128'he142c7ebe5d076fe01c65c2a4678b8b3, {16'd17154, 16'd10240, 16'd51565, 16'd59588, 16'd64772, 16'd6668, 16'd45438, 16'd50369, 16'd24896, 16'd21509, 16'd14166, 16'd11121, 16'd42908, 16'd59185, 16'd30576, 16'd51167, 16'd38264, 16'd3142, 16'd28180, 16'd41375, 16'd42256, 16'd54547, 16'd62749, 16'd32828, 16'd24748, 16'd50399});
	test_expansion(128'heb8197011517fa712c9975202b628683, {16'd57892, 16'd48841, 16'd43480, 16'd44367, 16'd40345, 16'd29142, 16'd4371, 16'd63181, 16'd47226, 16'd14671, 16'd64185, 16'd47996, 16'd23751, 16'd22090, 16'd56511, 16'd28123, 16'd9133, 16'd28022, 16'd25665, 16'd38531, 16'd39982, 16'd28387, 16'd11081, 16'd46632, 16'd29730, 16'd37772});
	test_expansion(128'h1938eee45d3f42abd7eab1042feaf6ca, {16'd65528, 16'd33777, 16'd47677, 16'd17705, 16'd54888, 16'd56144, 16'd7740, 16'd4144, 16'd51053, 16'd30642, 16'd32836, 16'd46643, 16'd21553, 16'd15711, 16'd37707, 16'd9631, 16'd47648, 16'd43857, 16'd4289, 16'd29941, 16'd22045, 16'd42423, 16'd34557, 16'd55684, 16'd15889, 16'd37197});
	test_expansion(128'h39deed73047e1c417db3fb59bb583162, {16'd30045, 16'd30979, 16'd18445, 16'd24553, 16'd3126, 16'd6231, 16'd62241, 16'd28402, 16'd30503, 16'd26578, 16'd43239, 16'd27161, 16'd30463, 16'd22912, 16'd57456, 16'd40746, 16'd59661, 16'd32635, 16'd61549, 16'd5772, 16'd32049, 16'd9988, 16'd62403, 16'd2922, 16'd52687, 16'd13022});
	test_expansion(128'h9f6e09d067ac1cb1e450cfbd2dcb977f, {16'd25566, 16'd20179, 16'd14653, 16'd39290, 16'd57778, 16'd15509, 16'd53702, 16'd56231, 16'd30010, 16'd11929, 16'd16469, 16'd56720, 16'd54452, 16'd52998, 16'd37151, 16'd51464, 16'd7391, 16'd34860, 16'd37588, 16'd14402, 16'd23660, 16'd6400, 16'd27855, 16'd29123, 16'd32302, 16'd26812});
	test_expansion(128'h7f8f0f04fd33573cd5cc054063adc33a, {16'd52007, 16'd18036, 16'd4518, 16'd19389, 16'd20615, 16'd23958, 16'd17438, 16'd39248, 16'd30488, 16'd19246, 16'd42257, 16'd40864, 16'd36410, 16'd14947, 16'd7077, 16'd8370, 16'd49418, 16'd48519, 16'd9764, 16'd26612, 16'd27986, 16'd61350, 16'd54227, 16'd4256, 16'd32166, 16'd50165});
	test_expansion(128'h994cc0d780a7763f42b83001c5f5e4a8, {16'd52430, 16'd55721, 16'd25283, 16'd51695, 16'd30152, 16'd41712, 16'd18894, 16'd411, 16'd7131, 16'd34966, 16'd7949, 16'd60917, 16'd60037, 16'd55806, 16'd31542, 16'd9812, 16'd64981, 16'd17486, 16'd15775, 16'd47213, 16'd51830, 16'd22109, 16'd34506, 16'd53336, 16'd55332, 16'd11257});
	test_expansion(128'hd0dd63773b3f5a0e063dac3933136144, {16'd10386, 16'd44360, 16'd30124, 16'd50555, 16'd14556, 16'd34638, 16'd37832, 16'd4768, 16'd40623, 16'd55646, 16'd28953, 16'd11595, 16'd6918, 16'd8738, 16'd38733, 16'd51042, 16'd13417, 16'd39246, 16'd2882, 16'd43238, 16'd5490, 16'd5972, 16'd33014, 16'd63273, 16'd17990, 16'd20280});
	test_expansion(128'hcf04ef93d01ebbf896509d9220857866, {16'd18211, 16'd15034, 16'd18724, 16'd52361, 16'd30514, 16'd41457, 16'd47754, 16'd18693, 16'd25463, 16'd20321, 16'd37857, 16'd55874, 16'd32418, 16'd57579, 16'd21160, 16'd12917, 16'd25256, 16'd30172, 16'd48968, 16'd39451, 16'd47816, 16'd48915, 16'd298, 16'd26932, 16'd44846, 16'd30915});
	test_expansion(128'hf0245950e15511f0c681932790150dcd, {16'd22304, 16'd39517, 16'd5006, 16'd22701, 16'd57227, 16'd4936, 16'd20422, 16'd24760, 16'd16415, 16'd63070, 16'd34366, 16'd64012, 16'd18868, 16'd55615, 16'd1839, 16'd34728, 16'd5517, 16'd43641, 16'd25820, 16'd22264, 16'd7107, 16'd48104, 16'd29042, 16'd19925, 16'd46432, 16'd1874});
	test_expansion(128'h904702b857a592aacb0f7c08bf6fb011, {16'd56006, 16'd43958, 16'd36322, 16'd4813, 16'd28850, 16'd9017, 16'd62177, 16'd35039, 16'd60352, 16'd36279, 16'd57115, 16'd46781, 16'd13895, 16'd51395, 16'd40861, 16'd38764, 16'd28818, 16'd62285, 16'd16987, 16'd28337, 16'd15975, 16'd14562, 16'd57633, 16'd49889, 16'd61335, 16'd10585});
	test_expansion(128'h523daf68d7f32cdf1ed975c778a4ac1a, {16'd28216, 16'd4103, 16'd21561, 16'd2262, 16'd26770, 16'd11115, 16'd56008, 16'd37745, 16'd10426, 16'd58213, 16'd47105, 16'd36543, 16'd39447, 16'd5125, 16'd6945, 16'd12283, 16'd10983, 16'd9988, 16'd53895, 16'd39777, 16'd46909, 16'd28189, 16'd11749, 16'd50634, 16'd19585, 16'd8088});
	test_expansion(128'h55bb4b2633e1217c95aba312dd8f1c81, {16'd36334, 16'd46752, 16'd35334, 16'd4301, 16'd56074, 16'd40890, 16'd60577, 16'd31094, 16'd48423, 16'd38901, 16'd35373, 16'd47006, 16'd35778, 16'd13386, 16'd42958, 16'd22568, 16'd9820, 16'd35066, 16'd3590, 16'd36816, 16'd55443, 16'd24064, 16'd6619, 16'd20754, 16'd33355, 16'd64489});
	test_expansion(128'heb91b35e1c73df3db8bbc2d6acc01fe0, {16'd9320, 16'd31136, 16'd34472, 16'd16349, 16'd52775, 16'd1701, 16'd17286, 16'd58712, 16'd45092, 16'd12157, 16'd33019, 16'd54495, 16'd237, 16'd10885, 16'd55715, 16'd26452, 16'd14351, 16'd28570, 16'd30655, 16'd34049, 16'd10559, 16'd36560, 16'd14876, 16'd205, 16'd16547, 16'd59501});
	test_expansion(128'h11298c7fa474fa7a9f2676d8dff082de, {16'd41174, 16'd24556, 16'd30220, 16'd36987, 16'd62789, 16'd4775, 16'd8959, 16'd58337, 16'd34338, 16'd64981, 16'd57932, 16'd62179, 16'd6329, 16'd52901, 16'd16637, 16'd910, 16'd27710, 16'd12940, 16'd42170, 16'd25864, 16'd32770, 16'd45843, 16'd63799, 16'd27429, 16'd64990, 16'd13808});
	test_expansion(128'h62a6b2e64577745dc20e4490794541b3, {16'd12224, 16'd10380, 16'd35574, 16'd61101, 16'd8345, 16'd801, 16'd57976, 16'd22603, 16'd41025, 16'd16288, 16'd44940, 16'd46971, 16'd7702, 16'd32824, 16'd46466, 16'd24568, 16'd11986, 16'd63246, 16'd51386, 16'd33906, 16'd27231, 16'd5393, 16'd50458, 16'd31850, 16'd1935, 16'd33347});
	test_expansion(128'hebeb6129c64823a5f7e1083b14c831ae, {16'd60962, 16'd43583, 16'd38152, 16'd35802, 16'd58667, 16'd48507, 16'd14953, 16'd40936, 16'd64637, 16'd3169, 16'd14781, 16'd11047, 16'd17841, 16'd63821, 16'd28700, 16'd43021, 16'd38308, 16'd51923, 16'd17957, 16'd3150, 16'd6449, 16'd27580, 16'd47722, 16'd65329, 16'd56909, 16'd28377});
	test_expansion(128'h9a64e46b9d1a9fd6d8474ad524a854c6, {16'd11217, 16'd58600, 16'd46394, 16'd61955, 16'd63498, 16'd9846, 16'd20089, 16'd49292, 16'd38604, 16'd53222, 16'd16856, 16'd14985, 16'd43001, 16'd63730, 16'd3319, 16'd1609, 16'd50690, 16'd11693, 16'd33183, 16'd12257, 16'd10946, 16'd53418, 16'd22801, 16'd56937, 16'd51043, 16'd10864});
	test_expansion(128'h879d9046b7da75a689f930e466412bb2, {16'd338, 16'd6835, 16'd7679, 16'd58203, 16'd55234, 16'd52796, 16'd32707, 16'd10937, 16'd60508, 16'd51382, 16'd26803, 16'd48135, 16'd7815, 16'd54679, 16'd42067, 16'd58136, 16'd7363, 16'd22858, 16'd52263, 16'd41740, 16'd15781, 16'd19919, 16'd43652, 16'd19253, 16'd55340, 16'd60303});
	test_expansion(128'h445b2ca15887fb44d29a6f41344b4e17, {16'd16303, 16'd64124, 16'd40280, 16'd15164, 16'd39033, 16'd51279, 16'd23053, 16'd29840, 16'd37636, 16'd13990, 16'd64415, 16'd1100, 16'd44191, 16'd1946, 16'd37815, 16'd6546, 16'd50597, 16'd43648, 16'd57307, 16'd16725, 16'd11670, 16'd55718, 16'd49388, 16'd2688, 16'd9785, 16'd54382});
	test_expansion(128'h7e44f59184cce1e5eeb5e62f9f6a648d, {16'd59569, 16'd51816, 16'd43809, 16'd51934, 16'd40825, 16'd48331, 16'd51291, 16'd19526, 16'd12401, 16'd28012, 16'd39509, 16'd60424, 16'd14307, 16'd3803, 16'd35304, 16'd23884, 16'd1682, 16'd39378, 16'd14330, 16'd54690, 16'd42854, 16'd23274, 16'd17646, 16'd40166, 16'd44667, 16'd36529});
	test_expansion(128'h6447807de270ff5b10c8464d974b4f17, {16'd45123, 16'd39567, 16'd19852, 16'd33974, 16'd6990, 16'd40010, 16'd21461, 16'd43476, 16'd10153, 16'd19599, 16'd57117, 16'd57942, 16'd9392, 16'd58417, 16'd23382, 16'd7959, 16'd24103, 16'd12754, 16'd36416, 16'd55340, 16'd34490, 16'd13014, 16'd27298, 16'd35047, 16'd19898, 16'd11192});
	test_expansion(128'h1316a2d72b7eca58b00ac63b1ebf6465, {16'd45251, 16'd39363, 16'd49160, 16'd31336, 16'd45686, 16'd9224, 16'd59066, 16'd4382, 16'd3743, 16'd61721, 16'd46604, 16'd46571, 16'd47863, 16'd17385, 16'd40989, 16'd53919, 16'd16483, 16'd15843, 16'd14532, 16'd31280, 16'd3639, 16'd53257, 16'd10947, 16'd48667, 16'd24217, 16'd64823});
	test_expansion(128'h47ee273723c1d6aa64c66b4694f3c609, {16'd62230, 16'd52571, 16'd62341, 16'd51502, 16'd30219, 16'd25629, 16'd52910, 16'd3389, 16'd60305, 16'd44919, 16'd18237, 16'd41529, 16'd18963, 16'd52353, 16'd32334, 16'd26730, 16'd61955, 16'd21884, 16'd23398, 16'd36182, 16'd4880, 16'd38294, 16'd57443, 16'd50156, 16'd14889, 16'd34111});
	test_expansion(128'h591434fb9a21c97cecbbd9a84ab04608, {16'd61429, 16'd5114, 16'd20757, 16'd16800, 16'd48709, 16'd44922, 16'd19989, 16'd49940, 16'd32173, 16'd41732, 16'd48023, 16'd49863, 16'd46480, 16'd23376, 16'd53438, 16'd2546, 16'd4060, 16'd60241, 16'd54959, 16'd42962, 16'd4443, 16'd21093, 16'd32064, 16'd39267, 16'd58030, 16'd57140});
	test_expansion(128'h6ecd6c579f8c41f255655fdbd10aff98, {16'd10539, 16'd27438, 16'd48044, 16'd47229, 16'd63202, 16'd43163, 16'd33653, 16'd49622, 16'd57136, 16'd54762, 16'd55604, 16'd48092, 16'd35530, 16'd52830, 16'd26530, 16'd28219, 16'd55030, 16'd57710, 16'd6013, 16'd10042, 16'd31975, 16'd18658, 16'd36046, 16'd7726, 16'd50579, 16'd63087});
	test_expansion(128'h06c01f92960a2cb75a65ac6ad5e8b89a, {16'd21048, 16'd33999, 16'd14926, 16'd47287, 16'd17297, 16'd56318, 16'd8590, 16'd41602, 16'd28495, 16'd9703, 16'd29642, 16'd40411, 16'd55859, 16'd22995, 16'd4258, 16'd63495, 16'd17286, 16'd56207, 16'd7523, 16'd37787, 16'd28374, 16'd57278, 16'd34259, 16'd37978, 16'd45164, 16'd16078});
	test_expansion(128'hf90f0f7ed45495cad455b24684b011f1, {16'd52918, 16'd65034, 16'd56617, 16'd22294, 16'd12373, 16'd14599, 16'd23512, 16'd385, 16'd45900, 16'd53047, 16'd55208, 16'd348, 16'd24213, 16'd46971, 16'd48479, 16'd15467, 16'd60013, 16'd55072, 16'd2921, 16'd25919, 16'd35904, 16'd5438, 16'd45625, 16'd7148, 16'd32467, 16'd36686});
	test_expansion(128'h175167f1b30fd98891b3fe43b4c8c901, {16'd26361, 16'd65533, 16'd33756, 16'd41597, 16'd60195, 16'd53501, 16'd11878, 16'd20649, 16'd56380, 16'd8150, 16'd58482, 16'd7143, 16'd40140, 16'd59150, 16'd16024, 16'd4173, 16'd2947, 16'd34005, 16'd20443, 16'd57506, 16'd14038, 16'd28016, 16'd14848, 16'd62539, 16'd35953, 16'd8915});
	test_expansion(128'heebec3c402bd86560cd3361ef0c3099a, {16'd25073, 16'd63355, 16'd10198, 16'd59693, 16'd15345, 16'd28580, 16'd57291, 16'd45286, 16'd15424, 16'd43712, 16'd53344, 16'd43046, 16'd1329, 16'd32001, 16'd56099, 16'd8156, 16'd20248, 16'd7219, 16'd26270, 16'd62153, 16'd53344, 16'd45553, 16'd38874, 16'd27573, 16'd32829, 16'd44047});
	test_expansion(128'h24ae63bc83ae0dd8701b0814efa4d6fd, {16'd18950, 16'd42168, 16'd7463, 16'd55094, 16'd4292, 16'd2415, 16'd11987, 16'd47433, 16'd42450, 16'd11132, 16'd33403, 16'd1976, 16'd58839, 16'd35549, 16'd50810, 16'd24941, 16'd52113, 16'd54654, 16'd14680, 16'd43981, 16'd29882, 16'd46597, 16'd33942, 16'd49647, 16'd31775, 16'd58789});
	test_expansion(128'h24d88e18b384cc10a838963c0b9c1717, {16'd21497, 16'd2016, 16'd6020, 16'd23562, 16'd46776, 16'd55038, 16'd11191, 16'd13450, 16'd63195, 16'd41647, 16'd25459, 16'd16482, 16'd21926, 16'd37172, 16'd57335, 16'd29144, 16'd52969, 16'd48704, 16'd31791, 16'd51318, 16'd18914, 16'd29625, 16'd11053, 16'd38647, 16'd53178, 16'd52461});
	test_expansion(128'h38a32374980a93efe013ca826d81f0c4, {16'd7308, 16'd4584, 16'd7016, 16'd33238, 16'd63560, 16'd32797, 16'd52912, 16'd19356, 16'd7723, 16'd8892, 16'd60313, 16'd8326, 16'd21858, 16'd40448, 16'd18652, 16'd34590, 16'd42970, 16'd1511, 16'd43382, 16'd35796, 16'd21832, 16'd18476, 16'd5927, 16'd47471, 16'd38673, 16'd58406});
	test_expansion(128'hee4e2ad4bda182c68eee75d37444f309, {16'd55992, 16'd6436, 16'd64657, 16'd52054, 16'd20082, 16'd13653, 16'd5138, 16'd340, 16'd46456, 16'd6919, 16'd22773, 16'd55578, 16'd31199, 16'd4095, 16'd52089, 16'd16010, 16'd36149, 16'd21178, 16'd17358, 16'd25474, 16'd45209, 16'd7562, 16'd19417, 16'd8521, 16'd39072, 16'd16431});
	test_expansion(128'h5c6aa5b57e36ccc4e6c50e65c88b03a5, {16'd9430, 16'd36581, 16'd47717, 16'd19557, 16'd17697, 16'd16150, 16'd10595, 16'd6944, 16'd36567, 16'd19907, 16'd41286, 16'd32175, 16'd37176, 16'd40643, 16'd29887, 16'd22236, 16'd28657, 16'd12821, 16'd4525, 16'd53963, 16'd60000, 16'd4658, 16'd56865, 16'd57539, 16'd17914, 16'd60265});
	test_expansion(128'h337f2a83dc91c7e149882a87a9d26f79, {16'd61339, 16'd35993, 16'd61068, 16'd39635, 16'd36865, 16'd4987, 16'd41066, 16'd34680, 16'd4112, 16'd37415, 16'd60342, 16'd25509, 16'd56807, 16'd47975, 16'd37909, 16'd4352, 16'd10471, 16'd30629, 16'd64969, 16'd60930, 16'd25824, 16'd15792, 16'd42797, 16'd23355, 16'd63570, 16'd53858});
	test_expansion(128'he03fe945fd93b980e3617d4332945f83, {16'd18470, 16'd14151, 16'd57989, 16'd50873, 16'd2170, 16'd24200, 16'd51213, 16'd33953, 16'd5547, 16'd16198, 16'd49710, 16'd64087, 16'd46567, 16'd53534, 16'd7571, 16'd56236, 16'd17000, 16'd36413, 16'd62687, 16'd42527, 16'd13084, 16'd58214, 16'd49646, 16'd63953, 16'd57, 16'd30269});
	test_expansion(128'hd06e131da3aa00c79137d70cee4547b2, {16'd18105, 16'd11611, 16'd60856, 16'd47056, 16'd1865, 16'd46946, 16'd37046, 16'd48531, 16'd41949, 16'd2955, 16'd40671, 16'd21867, 16'd3930, 16'd744, 16'd33552, 16'd10070, 16'd60814, 16'd14721, 16'd9290, 16'd53764, 16'd27892, 16'd2118, 16'd57221, 16'd32672, 16'd59424, 16'd63967});
	test_expansion(128'h6e672ebc940e4fe54ba1fc679f55cbb6, {16'd19875, 16'd9824, 16'd43327, 16'd40074, 16'd49073, 16'd1291, 16'd20878, 16'd20862, 16'd17454, 16'd59177, 16'd749, 16'd8534, 16'd55065, 16'd57205, 16'd27884, 16'd48831, 16'd7474, 16'd43427, 16'd56832, 16'd1240, 16'd23273, 16'd12008, 16'd51804, 16'd20578, 16'd55917, 16'd7858});
	test_expansion(128'h9c2336d9b33c94e37164c0893eda00d0, {16'd38564, 16'd60020, 16'd943, 16'd28265, 16'd35552, 16'd35365, 16'd10747, 16'd40382, 16'd47344, 16'd26410, 16'd28211, 16'd35240, 16'd21127, 16'd64092, 16'd48004, 16'd1912, 16'd4912, 16'd36381, 16'd6200, 16'd41496, 16'd52783, 16'd26611, 16'd21696, 16'd1785, 16'd32842, 16'd53568});
	test_expansion(128'h29e1a4f044f34228c6e03ec35dfb90d6, {16'd28493, 16'd49813, 16'd31170, 16'd38521, 16'd53124, 16'd49027, 16'd3329, 16'd10650, 16'd62815, 16'd29550, 16'd62409, 16'd30203, 16'd5057, 16'd10637, 16'd59901, 16'd1566, 16'd29583, 16'd46630, 16'd61703, 16'd54007, 16'd34404, 16'd36891, 16'd38764, 16'd30458, 16'd31343, 16'd52745});
	test_expansion(128'hb561c640cdad621f9027c471b35f5e3b, {16'd60581, 16'd21630, 16'd43783, 16'd46673, 16'd29383, 16'd11141, 16'd58052, 16'd41833, 16'd64049, 16'd61100, 16'd53036, 16'd52530, 16'd1074, 16'd42367, 16'd50809, 16'd27469, 16'd55593, 16'd21538, 16'd25411, 16'd13455, 16'd37527, 16'd47376, 16'd48682, 16'd14997, 16'd62663, 16'd48665});
	test_expansion(128'h9c806ec434efab439b4afb7ae9836383, {16'd38309, 16'd54118, 16'd31851, 16'd36139, 16'd7927, 16'd31855, 16'd40902, 16'd58334, 16'd63753, 16'd64025, 16'd44738, 16'd47634, 16'd63962, 16'd50386, 16'd45441, 16'd35558, 16'd40274, 16'd56269, 16'd41655, 16'd54159, 16'd29045, 16'd37137, 16'd63485, 16'd63314, 16'd7841, 16'd47573});
	test_expansion(128'ha959efe3fcc2106087e02ac1cbf2ea5b, {16'd47230, 16'd39047, 16'd57456, 16'd10654, 16'd6893, 16'd17836, 16'd62996, 16'd23592, 16'd42550, 16'd17945, 16'd32102, 16'd4572, 16'd43507, 16'd58237, 16'd55013, 16'd5032, 16'd3327, 16'd42348, 16'd24122, 16'd27260, 16'd24936, 16'd56347, 16'd2660, 16'd61270, 16'd6828, 16'd51045});
	test_expansion(128'hbe3af408acba32d18a9f70e3efeb8bac, {16'd11539, 16'd6419, 16'd19268, 16'd64587, 16'd43764, 16'd15362, 16'd42750, 16'd17647, 16'd64932, 16'd43525, 16'd60828, 16'd6904, 16'd37330, 16'd50349, 16'd35898, 16'd14380, 16'd3012, 16'd12745, 16'd32891, 16'd5865, 16'd14246, 16'd39287, 16'd27334, 16'd5706, 16'd47997, 16'd20757});
	test_expansion(128'he0bd115b9dafc11365e547adc06e8bd6, {16'd9972, 16'd57758, 16'd15012, 16'd49772, 16'd898, 16'd19192, 16'd35471, 16'd4291, 16'd14324, 16'd45920, 16'd41249, 16'd58007, 16'd2714, 16'd15365, 16'd32749, 16'd26494, 16'd56465, 16'd23676, 16'd16141, 16'd47149, 16'd6818, 16'd15699, 16'd1981, 16'd53380, 16'd57289, 16'd3133});
	test_expansion(128'he3d00efaa232200081e35c4a84ea9eb7, {16'd28235, 16'd8052, 16'd38243, 16'd56198, 16'd773, 16'd49104, 16'd27678, 16'd54919, 16'd45830, 16'd63097, 16'd31267, 16'd9285, 16'd48435, 16'd24420, 16'd20694, 16'd34581, 16'd29407, 16'd4387, 16'd2861, 16'd14248, 16'd51337, 16'd54476, 16'd15469, 16'd43800, 16'd10385, 16'd61030});
	test_expansion(128'h422eb7bd9c9e4abdd388ba612a2b8e91, {16'd17249, 16'd25180, 16'd32916, 16'd23438, 16'd699, 16'd56367, 16'd39053, 16'd28027, 16'd61952, 16'd11891, 16'd17102, 16'd36261, 16'd22486, 16'd3616, 16'd23825, 16'd31500, 16'd33306, 16'd24024, 16'd58328, 16'd38843, 16'd28405, 16'd24006, 16'd19991, 16'd29075, 16'd6029, 16'd9072});
	test_expansion(128'had10fa8b119c68c9c552175fa6a473fd, {16'd38717, 16'd49764, 16'd51043, 16'd13714, 16'd4338, 16'd5060, 16'd18295, 16'd8281, 16'd60954, 16'd8266, 16'd15022, 16'd32243, 16'd2464, 16'd61325, 16'd38049, 16'd31081, 16'd44411, 16'd9335, 16'd24214, 16'd52836, 16'd10623, 16'd55522, 16'd44228, 16'd43961, 16'd17562, 16'd35568});
	test_expansion(128'h506d0b2710d40929f26b49bdbae0c8bd, {16'd18214, 16'd13729, 16'd18194, 16'd10415, 16'd13458, 16'd12320, 16'd60340, 16'd37769, 16'd3989, 16'd17205, 16'd1660, 16'd18748, 16'd30116, 16'd14016, 16'd304, 16'd32379, 16'd65305, 16'd27162, 16'd53412, 16'd39272, 16'd62132, 16'd26055, 16'd48217, 16'd14598, 16'd35000, 16'd45862});
	test_expansion(128'he4f434208e1ab5c6da868617098a7fb1, {16'd36831, 16'd6687, 16'd33889, 16'd186, 16'd28458, 16'd3938, 16'd30494, 16'd49417, 16'd4499, 16'd62087, 16'd49673, 16'd53345, 16'd63619, 16'd62032, 16'd3982, 16'd13382, 16'd11582, 16'd39113, 16'd50604, 16'd56079, 16'd28008, 16'd16116, 16'd22220, 16'd8203, 16'd44204, 16'd49168});
	test_expansion(128'h813c6e50fa0b8184e51edd8346e4f611, {16'd27533, 16'd17550, 16'd9364, 16'd15478, 16'd28586, 16'd59155, 16'd11334, 16'd23138, 16'd45819, 16'd43380, 16'd47049, 16'd10745, 16'd25067, 16'd59655, 16'd59663, 16'd50354, 16'd356, 16'd62191, 16'd28373, 16'd30580, 16'd53574, 16'd26321, 16'd14414, 16'd63796, 16'd632, 16'd37282});
	test_expansion(128'h8b45607968ad22adb587a99e27ffef0d, {16'd36078, 16'd16192, 16'd55686, 16'd24274, 16'd9605, 16'd34398, 16'd9631, 16'd25107, 16'd51770, 16'd1387, 16'd34979, 16'd5701, 16'd43220, 16'd21849, 16'd45654, 16'd38360, 16'd57248, 16'd51142, 16'd10307, 16'd11637, 16'd17690, 16'd22855, 16'd23392, 16'd47526, 16'd31751, 16'd42405});
	test_expansion(128'h30f80316268e388423cc2bbb3ab858c2, {16'd29628, 16'd41466, 16'd32556, 16'd16343, 16'd32867, 16'd36535, 16'd62264, 16'd37256, 16'd7166, 16'd40803, 16'd42068, 16'd36389, 16'd18758, 16'd47989, 16'd4464, 16'd44998, 16'd38465, 16'd61106, 16'd50061, 16'd12299, 16'd6774, 16'd56340, 16'd44905, 16'd59054, 16'd10087, 16'd25191});
	test_expansion(128'hba9bfca559157b1137eaabc59ca755a7, {16'd496, 16'd31856, 16'd25835, 16'd56834, 16'd3890, 16'd26186, 16'd15880, 16'd41523, 16'd32002, 16'd1723, 16'd50193, 16'd30506, 16'd42095, 16'd5418, 16'd15673, 16'd37105, 16'd24860, 16'd14253, 16'd4451, 16'd2647, 16'd45644, 16'd35740, 16'd9766, 16'd50625, 16'd14615, 16'd4650});
	test_expansion(128'ha7dcacd468203a4b08313978cc242dc6, {16'd14519, 16'd47419, 16'd15599, 16'd28237, 16'd49058, 16'd60222, 16'd20287, 16'd2198, 16'd15694, 16'd11332, 16'd46488, 16'd32968, 16'd30721, 16'd34409, 16'd13648, 16'd38760, 16'd22908, 16'd28004, 16'd12587, 16'd47275, 16'd43824, 16'd34785, 16'd46034, 16'd30259, 16'd52255, 16'd62799});
	test_expansion(128'h48778bee1b2548745c76ca25fede4421, {16'd53789, 16'd57974, 16'd36072, 16'd900, 16'd31588, 16'd13144, 16'd57750, 16'd36804, 16'd4034, 16'd22985, 16'd25361, 16'd30342, 16'd60029, 16'd1983, 16'd37873, 16'd26985, 16'd35530, 16'd27601, 16'd55337, 16'd31497, 16'd21810, 16'd36232, 16'd48688, 16'd55208, 16'd31411, 16'd48911});
	test_expansion(128'hcc360a81e9e156cf025315b6e1595e39, {16'd14368, 16'd38131, 16'd61786, 16'd38858, 16'd14801, 16'd44215, 16'd8745, 16'd53472, 16'd38444, 16'd50429, 16'd12412, 16'd5336, 16'd25473, 16'd53604, 16'd42531, 16'd50625, 16'd19503, 16'd1160, 16'd53660, 16'd42052, 16'd43514, 16'd30192, 16'd57620, 16'd24719, 16'd5804, 16'd8197});
	test_expansion(128'h14dbc17cc42e5253fec97aad72a173f5, {16'd22464, 16'd33127, 16'd15973, 16'd14047, 16'd43691, 16'd20568, 16'd42750, 16'd39670, 16'd18564, 16'd35625, 16'd49083, 16'd36218, 16'd23735, 16'd32092, 16'd58368, 16'd59758, 16'd27442, 16'd51845, 16'd14906, 16'd63797, 16'd56711, 16'd31711, 16'd2619, 16'd53564, 16'd52502, 16'd52653});
	test_expansion(128'h49c3e39937a659a069cf7cb1bb35f653, {16'd12922, 16'd9825, 16'd65047, 16'd11465, 16'd19538, 16'd7584, 16'd60599, 16'd40853, 16'd9928, 16'd56582, 16'd3346, 16'd11963, 16'd31411, 16'd39187, 16'd20170, 16'd57859, 16'd2030, 16'd36504, 16'd49957, 16'd4288, 16'd63877, 16'd4116, 16'd15242, 16'd5194, 16'd34339, 16'd20599});
	test_expansion(128'h7b7810b695893f6dc65d6a7ff678838b, {16'd6952, 16'd12501, 16'd17877, 16'd1224, 16'd52363, 16'd10886, 16'd53334, 16'd36714, 16'd17641, 16'd56562, 16'd47106, 16'd52396, 16'd39771, 16'd31684, 16'd29775, 16'd43999, 16'd17904, 16'd19153, 16'd4856, 16'd55084, 16'd24244, 16'd40874, 16'd14780, 16'd53457, 16'd47685, 16'd52498});
	test_expansion(128'h5ffc2438196a4d3434c06ea8e61aa2ed, {16'd4369, 16'd11062, 16'd36003, 16'd10873, 16'd64039, 16'd53666, 16'd60232, 16'd62488, 16'd51575, 16'd21300, 16'd27266, 16'd40676, 16'd47521, 16'd58406, 16'd19526, 16'd63023, 16'd38379, 16'd16525, 16'd46548, 16'd38405, 16'd16865, 16'd58335, 16'd26684, 16'd30765, 16'd33044, 16'd31667});
	test_expansion(128'he029283248288a3991cd8ed803a2d0ab, {16'd53693, 16'd23430, 16'd22966, 16'd63202, 16'd25291, 16'd46174, 16'd15923, 16'd23982, 16'd20469, 16'd10756, 16'd12930, 16'd33697, 16'd5502, 16'd9377, 16'd64017, 16'd41709, 16'd34313, 16'd30294, 16'd30208, 16'd19751, 16'd65299, 16'd23206, 16'd19043, 16'd3642, 16'd41522, 16'd62887});
	test_expansion(128'hb42e2a11b0fbed904af21b84d07d73ec, {16'd5947, 16'd64987, 16'd64727, 16'd12268, 16'd31846, 16'd16871, 16'd39110, 16'd65109, 16'd53344, 16'd42322, 16'd18944, 16'd48504, 16'd11647, 16'd32952, 16'd51753, 16'd19564, 16'd12622, 16'd6920, 16'd3744, 16'd51476, 16'd29342, 16'd21916, 16'd23161, 16'd23946, 16'd63688, 16'd44976});
	test_expansion(128'h6adf2295393e836cf78ef91c78fd55e9, {16'd6195, 16'd33643, 16'd18868, 16'd50538, 16'd33640, 16'd4992, 16'd32412, 16'd3373, 16'd20565, 16'd58165, 16'd51791, 16'd2435, 16'd53291, 16'd62268, 16'd12485, 16'd14050, 16'd35028, 16'd25038, 16'd27083, 16'd54132, 16'd33443, 16'd27329, 16'd52198, 16'd17076, 16'd14087, 16'd51331});
	test_expansion(128'h4b837410b438bc5068632fd4c0a62c5d, {16'd19368, 16'd50664, 16'd21320, 16'd52649, 16'd30049, 16'd1594, 16'd59688, 16'd58791, 16'd23526, 16'd16956, 16'd40285, 16'd63590, 16'd59341, 16'd34658, 16'd63494, 16'd45778, 16'd31983, 16'd44990, 16'd42277, 16'd51015, 16'd24236, 16'd17789, 16'd52464, 16'd50165, 16'd30544, 16'd6552});
	test_expansion(128'ha86b7adc2b78ee9e2b21898708eef3dd, {16'd15043, 16'd49744, 16'd2812, 16'd6927, 16'd45631, 16'd23279, 16'd28153, 16'd20502, 16'd9432, 16'd27159, 16'd10928, 16'd9650, 16'd34149, 16'd60497, 16'd42112, 16'd57920, 16'd51206, 16'd9841, 16'd18536, 16'd21249, 16'd40811, 16'd36517, 16'd23659, 16'd8191, 16'd50219, 16'd64788});
	test_expansion(128'h7810dc14d0cf1c1e563d26fc38f02770, {16'd58162, 16'd4808, 16'd10280, 16'd28985, 16'd48255, 16'd57863, 16'd37035, 16'd41554, 16'd15318, 16'd11149, 16'd12720, 16'd18332, 16'd24740, 16'd16670, 16'd38582, 16'd25317, 16'd5441, 16'd44453, 16'd21340, 16'd65082, 16'd37353, 16'd48318, 16'd450, 16'd64083, 16'd31090, 16'd8112});
	test_expansion(128'h2c2fb9472b234a72b794c7ee038780b8, {16'd62131, 16'd40233, 16'd32674, 16'd2217, 16'd32526, 16'd64432, 16'd37727, 16'd44544, 16'd17442, 16'd43342, 16'd51365, 16'd46582, 16'd44314, 16'd49139, 16'd27950, 16'd28219, 16'd29061, 16'd12962, 16'd5605, 16'd41188, 16'd7653, 16'd40076, 16'd51176, 16'd48945, 16'd25091, 16'd3466});
	test_expansion(128'h60d7cba694c30d0021436a2fbd771ea2, {16'd20256, 16'd25530, 16'd48751, 16'd30165, 16'd50425, 16'd6566, 16'd38858, 16'd1533, 16'd5868, 16'd8509, 16'd49570, 16'd49343, 16'd20638, 16'd49001, 16'd24635, 16'd21905, 16'd63966, 16'd23460, 16'd1230, 16'd6013, 16'd2074, 16'd58161, 16'd25057, 16'd15296, 16'd12110, 16'd13141});
	test_expansion(128'h0a88ff1814811d1925a54351e5418248, {16'd12247, 16'd63074, 16'd33795, 16'd17405, 16'd60133, 16'd42196, 16'd20040, 16'd28321, 16'd61297, 16'd64059, 16'd41802, 16'd16467, 16'd58978, 16'd61385, 16'd22222, 16'd7325, 16'd7498, 16'd14769, 16'd51549, 16'd54384, 16'd40219, 16'd1347, 16'd65294, 16'd22646, 16'd31278, 16'd62053});
	test_expansion(128'h5f58f05192c0a0cb115251ae3e509e3d, {16'd36104, 16'd20968, 16'd25308, 16'd40978, 16'd32089, 16'd53311, 16'd19831, 16'd44084, 16'd22630, 16'd17135, 16'd6243, 16'd27968, 16'd44118, 16'd58994, 16'd16953, 16'd37169, 16'd29067, 16'd43114, 16'd50813, 16'd8229, 16'd59097, 16'd14254, 16'd6495, 16'd40230, 16'd41720, 16'd29008});
	test_expansion(128'hcbd137f7f015accfc5b6b55e1349015b, {16'd64252, 16'd62890, 16'd34463, 16'd25600, 16'd36654, 16'd49792, 16'd15642, 16'd26194, 16'd23079, 16'd61466, 16'd11013, 16'd49647, 16'd26517, 16'd142, 16'd48495, 16'd12706, 16'd15971, 16'd51669, 16'd38362, 16'd40042, 16'd59651, 16'd55984, 16'd2493, 16'd20106, 16'd17067, 16'd19010});
	test_expansion(128'hd8d87d4fa8979f50af0d36f02743b9cc, {16'd59033, 16'd30393, 16'd28911, 16'd17761, 16'd34033, 16'd48689, 16'd19164, 16'd55781, 16'd24039, 16'd42401, 16'd63388, 16'd53895, 16'd42461, 16'd41991, 16'd3767, 16'd28643, 16'd34843, 16'd13112, 16'd26902, 16'd38056, 16'd61206, 16'd13141, 16'd14283, 16'd60028, 16'd18493, 16'd46520});
	test_expansion(128'h002c193d1ff5f480c75e7cfc44f8cee9, {16'd57164, 16'd32234, 16'd30696, 16'd53650, 16'd9621, 16'd62294, 16'd46020, 16'd27654, 16'd63454, 16'd34697, 16'd58942, 16'd9331, 16'd19752, 16'd58252, 16'd13203, 16'd16690, 16'd14751, 16'd22554, 16'd8913, 16'd60604, 16'd51120, 16'd38970, 16'd3398, 16'd3819, 16'd7511, 16'd63944});
	test_expansion(128'h079a7beacb1ac1cb674c639ca38e9b60, {16'd25667, 16'd40920, 16'd50320, 16'd17446, 16'd37805, 16'd56174, 16'd58999, 16'd26120, 16'd61534, 16'd29550, 16'd7489, 16'd11953, 16'd49014, 16'd34469, 16'd28152, 16'd37687, 16'd43817, 16'd48002, 16'd17893, 16'd38881, 16'd64050, 16'd47075, 16'd38992, 16'd58326, 16'd25341, 16'd2602});
	test_expansion(128'h6d791897f4069fcd1d3d19cdff3da2cf, {16'd60101, 16'd6950, 16'd58365, 16'd39606, 16'd48213, 16'd61191, 16'd56554, 16'd38594, 16'd33763, 16'd14025, 16'd63411, 16'd18261, 16'd55262, 16'd42349, 16'd41178, 16'd23560, 16'd18052, 16'd1236, 16'd62748, 16'd41226, 16'd36441, 16'd19554, 16'd42276, 16'd54569, 16'd26345, 16'd1267});
	test_expansion(128'heb18b87ff65f73d5e82dfda7187238a3, {16'd27595, 16'd9343, 16'd33656, 16'd4746, 16'd6755, 16'd28887, 16'd1298, 16'd64053, 16'd20777, 16'd57247, 16'd20405, 16'd45401, 16'd46570, 16'd11794, 16'd54578, 16'd4617, 16'd14648, 16'd54584, 16'd19545, 16'd22630, 16'd36656, 16'd39980, 16'd31606, 16'd990, 16'd33833, 16'd61323});
	test_expansion(128'h1b05650f8aea32a5e82f339a87adc1a4, {16'd25759, 16'd45896, 16'd41432, 16'd29226, 16'd64682, 16'd19237, 16'd9527, 16'd6735, 16'd55213, 16'd7606, 16'd62449, 16'd21431, 16'd27142, 16'd51880, 16'd4350, 16'd63625, 16'd38168, 16'd22853, 16'd8328, 16'd28876, 16'd36731, 16'd42663, 16'd50686, 16'd31713, 16'd43086, 16'd21679});
	test_expansion(128'hdaab707d0b66a6d8dd0233eb127d5a06, {16'd15490, 16'd18826, 16'd61371, 16'd6924, 16'd55242, 16'd41279, 16'd57544, 16'd17351, 16'd8234, 16'd4249, 16'd1149, 16'd20236, 16'd20905, 16'd29511, 16'd21852, 16'd47322, 16'd15896, 16'd54671, 16'd357, 16'd1583, 16'd54985, 16'd22037, 16'd36884, 16'd20896, 16'd6611, 16'd11612});
	test_expansion(128'h58907033374b76be66282c86e72941f3, {16'd42347, 16'd6810, 16'd7255, 16'd60561, 16'd24349, 16'd59693, 16'd45878, 16'd26251, 16'd11161, 16'd47892, 16'd25734, 16'd52218, 16'd42457, 16'd63051, 16'd2273, 16'd49679, 16'd22275, 16'd28838, 16'd31731, 16'd40857, 16'd32924, 16'd33173, 16'd16281, 16'd60800, 16'd11152, 16'd35686});
	test_expansion(128'h003a2814d9cc34badf1daee58d33fec5, {16'd20376, 16'd60577, 16'd22990, 16'd12080, 16'd25739, 16'd2399, 16'd40846, 16'd4713, 16'd10426, 16'd12442, 16'd32097, 16'd6503, 16'd52265, 16'd38807, 16'd53113, 16'd30546, 16'd61705, 16'd15539, 16'd61442, 16'd21844, 16'd35590, 16'd38064, 16'd10002, 16'd55166, 16'd38024, 16'd2893});
	test_expansion(128'hc2ab3abf6d851e97983e98352bcde28e, {16'd22017, 16'd33804, 16'd55364, 16'd24640, 16'd49823, 16'd47938, 16'd1739, 16'd10101, 16'd60026, 16'd7277, 16'd34176, 16'd13921, 16'd20000, 16'd23629, 16'd47723, 16'd39845, 16'd61364, 16'd28441, 16'd23221, 16'd62670, 16'd63098, 16'd39274, 16'd63134, 16'd13074, 16'd12627, 16'd2380});
	test_expansion(128'h13695574f4d158d9879674eff98df261, {16'd60354, 16'd38029, 16'd19149, 16'd61073, 16'd56342, 16'd50722, 16'd56193, 16'd29626, 16'd15952, 16'd3479, 16'd39895, 16'd15385, 16'd26670, 16'd5853, 16'd19259, 16'd15251, 16'd28263, 16'd47687, 16'd16273, 16'd59309, 16'd45112, 16'd56846, 16'd7091, 16'd56167, 16'd34349, 16'd4231});
	test_expansion(128'h946335dab93e4253edc8135f5827dcc4, {16'd30073, 16'd42119, 16'd42263, 16'd3291, 16'd25954, 16'd38510, 16'd9281, 16'd57259, 16'd30930, 16'd23783, 16'd39944, 16'd25155, 16'd33374, 16'd43353, 16'd54251, 16'd49549, 16'd35719, 16'd28918, 16'd61723, 16'd3361, 16'd34634, 16'd44192, 16'd7586, 16'd64832, 16'd19617, 16'd37602});
	test_expansion(128'hd64a233dfb5b282c711cc3951c11f1fb, {16'd7204, 16'd55093, 16'd64085, 16'd19656, 16'd2617, 16'd5315, 16'd5674, 16'd33174, 16'd50307, 16'd63047, 16'd17426, 16'd32519, 16'd14627, 16'd46307, 16'd22855, 16'd59376, 16'd16810, 16'd61599, 16'd54822, 16'd7762, 16'd16789, 16'd20785, 16'd21648, 16'd2891, 16'd31173, 16'd1067});
	test_expansion(128'h9924917ff5e72a455d31521047499e50, {16'd14892, 16'd38775, 16'd24730, 16'd49433, 16'd63632, 16'd24347, 16'd36118, 16'd37352, 16'd15470, 16'd52071, 16'd42961, 16'd59541, 16'd65149, 16'd63294, 16'd25146, 16'd62706, 16'd21472, 16'd62220, 16'd46665, 16'd6566, 16'd56841, 16'd4006, 16'd52240, 16'd61484, 16'd50059, 16'd3816});
	test_expansion(128'h9e8f0dd7789796742204a6840c149d82, {16'd32765, 16'd3139, 16'd62717, 16'd32874, 16'd21442, 16'd10144, 16'd22891, 16'd33306, 16'd53751, 16'd46717, 16'd26413, 16'd24010, 16'd50914, 16'd53471, 16'd35251, 16'd58249, 16'd52145, 16'd18493, 16'd17550, 16'd49346, 16'd25157, 16'd22883, 16'd32486, 16'd10597, 16'd46995, 16'd20546});
	test_expansion(128'hfdb6294a63f6d089c62bc73871120b2a, {16'd31593, 16'd11894, 16'd43457, 16'd24017, 16'd15926, 16'd10818, 16'd22957, 16'd33979, 16'd3320, 16'd40250, 16'd33526, 16'd45913, 16'd6075, 16'd39455, 16'd17413, 16'd46818, 16'd7454, 16'd13900, 16'd39787, 16'd50912, 16'd39156, 16'd65254, 16'd61788, 16'd19948, 16'd13168, 16'd62142});
	test_expansion(128'h6034dd529e2bf9a24792489e26311329, {16'd61775, 16'd63841, 16'd34113, 16'd38448, 16'd7758, 16'd28214, 16'd14371, 16'd20292, 16'd21024, 16'd58016, 16'd26887, 16'd10678, 16'd9696, 16'd5390, 16'd27449, 16'd38065, 16'd27201, 16'd27397, 16'd15751, 16'd9043, 16'd59397, 16'd49959, 16'd54715, 16'd9379, 16'd2506, 16'd1168});
	test_expansion(128'hec1d4e404da2dfdb3b4d5f2a7751944e, {16'd28877, 16'd31122, 16'd10386, 16'd46034, 16'd63701, 16'd19492, 16'd2783, 16'd12204, 16'd48873, 16'd13029, 16'd23486, 16'd17619, 16'd47617, 16'd34485, 16'd52236, 16'd7891, 16'd52510, 16'd57884, 16'd41097, 16'd14813, 16'd22373, 16'd48783, 16'd7390, 16'd28335, 16'd43459, 16'd55409});
	test_expansion(128'hb83744b63b484d2b965718ddea6e0924, {16'd43424, 16'd19411, 16'd44750, 16'd43253, 16'd52745, 16'd20227, 16'd31697, 16'd62459, 16'd29731, 16'd31087, 16'd37064, 16'd60616, 16'd11203, 16'd39609, 16'd50394, 16'd950, 16'd43435, 16'd14014, 16'd64600, 16'd25589, 16'd20244, 16'd49843, 16'd27829, 16'd3432, 16'd57845, 16'd18968});
	test_expansion(128'hd714b08e0a914d9164b3f2ff0546929e, {16'd59075, 16'd41703, 16'd44078, 16'd25244, 16'd32378, 16'd39703, 16'd55053, 16'd55847, 16'd62486, 16'd31965, 16'd2115, 16'd47383, 16'd61976, 16'd63259, 16'd63971, 16'd64271, 16'd58489, 16'd65313, 16'd59932, 16'd45078, 16'd44957, 16'd45866, 16'd15055, 16'd33600, 16'd65050, 16'd39416});
	test_expansion(128'h28ad63900f98a04e9b71af701894e859, {16'd51861, 16'd64855, 16'd32868, 16'd61154, 16'd48052, 16'd11919, 16'd1097, 16'd10647, 16'd35803, 16'd41186, 16'd51514, 16'd28889, 16'd3770, 16'd57260, 16'd40440, 16'd54397, 16'd26028, 16'd38031, 16'd698, 16'd32684, 16'd10737, 16'd33998, 16'd15358, 16'd43133, 16'd26032, 16'd12114});
	test_expansion(128'hab95543534d129a5a2c454dcb616f5cc, {16'd4372, 16'd28012, 16'd31179, 16'd28155, 16'd15261, 16'd25886, 16'd41288, 16'd16699, 16'd43682, 16'd60480, 16'd28507, 16'd9495, 16'd40594, 16'd55208, 16'd32862, 16'd54506, 16'd19551, 16'd60830, 16'd485, 16'd53668, 16'd37222, 16'd41283, 16'd65425, 16'd46674, 16'd49197, 16'd58402});
	test_expansion(128'h331beed885ac3899a76bdbd1e4432f03, {16'd33165, 16'd903, 16'd65179, 16'd49085, 16'd10571, 16'd1938, 16'd40965, 16'd51128, 16'd40847, 16'd58112, 16'd35175, 16'd24391, 16'd45215, 16'd53136, 16'd13759, 16'd238, 16'd44245, 16'd23660, 16'd23434, 16'd21932, 16'd32858, 16'd54293, 16'd64370, 16'd19463, 16'd43618, 16'd20741});
	test_expansion(128'h4797c060ffe5440d7fe9e414244e52ab, {16'd13058, 16'd23856, 16'd41919, 16'd38889, 16'd54609, 16'd58665, 16'd44148, 16'd3216, 16'd46086, 16'd2138, 16'd13354, 16'd15627, 16'd65327, 16'd16093, 16'd9523, 16'd8057, 16'd14377, 16'd44379, 16'd47255, 16'd52306, 16'd11985, 16'd486, 16'd56851, 16'd50099, 16'd2453, 16'd26879});
	test_expansion(128'h131b342f4150de618bae8212cf4fdf15, {16'd38467, 16'd54086, 16'd65194, 16'd26535, 16'd30604, 16'd2170, 16'd62090, 16'd29350, 16'd25849, 16'd25286, 16'd32554, 16'd55751, 16'd43881, 16'd10749, 16'd6676, 16'd5227, 16'd31958, 16'd43575, 16'd2299, 16'd64909, 16'd49441, 16'd29784, 16'd52127, 16'd56106, 16'd32009, 16'd44255});
	test_expansion(128'h21d8936f5fadd9f7fd1c8016012fad44, {16'd35240, 16'd15269, 16'd12245, 16'd15673, 16'd21853, 16'd28994, 16'd7718, 16'd58212, 16'd33869, 16'd14455, 16'd44659, 16'd28960, 16'd58315, 16'd39281, 16'd37779, 16'd36160, 16'd64680, 16'd49221, 16'd17114, 16'd43477, 16'd33395, 16'd21141, 16'd41920, 16'd30515, 16'd7526, 16'd19313});
	test_expansion(128'h786d370ec05d849f9f79da47589ec923, {16'd27860, 16'd59360, 16'd9344, 16'd9141, 16'd38248, 16'd49437, 16'd61108, 16'd22877, 16'd34853, 16'd20497, 16'd4603, 16'd8657, 16'd57721, 16'd50060, 16'd33663, 16'd24796, 16'd16613, 16'd4602, 16'd28425, 16'd25467, 16'd59644, 16'd38597, 16'd21368, 16'd29229, 16'd52885, 16'd44410});
	test_expansion(128'h894e281fc288da0ba24852c58ebd729a, {16'd21763, 16'd25714, 16'd18282, 16'd32217, 16'd41049, 16'd20473, 16'd24158, 16'd40929, 16'd62071, 16'd63683, 16'd38765, 16'd46828, 16'd31032, 16'd44737, 16'd7849, 16'd37690, 16'd10227, 16'd45191, 16'd50824, 16'd18033, 16'd14132, 16'd16311, 16'd37235, 16'd6008, 16'd9007, 16'd40102});
	test_expansion(128'h9199d42517c8a71acf05cb26faadc66a, {16'd34826, 16'd39942, 16'd54065, 16'd21576, 16'd65370, 16'd27547, 16'd29011, 16'd13614, 16'd61047, 16'd11624, 16'd25296, 16'd39479, 16'd47745, 16'd19388, 16'd56963, 16'd16676, 16'd64948, 16'd19100, 16'd51344, 16'd45254, 16'd31703, 16'd33824, 16'd46885, 16'd41083, 16'd61828, 16'd13640});
	test_expansion(128'hefcba538a147be786a2ebd255b6d39cb, {16'd30759, 16'd3604, 16'd60129, 16'd41634, 16'd48252, 16'd33689, 16'd27943, 16'd2235, 16'd35815, 16'd24694, 16'd14857, 16'd19244, 16'd918, 16'd24363, 16'd63460, 16'd53917, 16'd15742, 16'd639, 16'd5553, 16'd19850, 16'd5222, 16'd24343, 16'd38783, 16'd22414, 16'd52147, 16'd17052});
	test_expansion(128'h58bbd07ea32a5586c3a5ad636fa26942, {16'd41908, 16'd9584, 16'd39133, 16'd42981, 16'd49732, 16'd12644, 16'd32417, 16'd11277, 16'd39804, 16'd22047, 16'd24714, 16'd44866, 16'd20012, 16'd64357, 16'd37655, 16'd60576, 16'd51074, 16'd63718, 16'd58176, 16'd17039, 16'd7552, 16'd6018, 16'd17719, 16'd11655, 16'd9377, 16'd37223});
	test_expansion(128'hb297ab959e2764a84fef68c7553ea69e, {16'd10994, 16'd48722, 16'd33182, 16'd511, 16'd12762, 16'd10809, 16'd38456, 16'd56968, 16'd42982, 16'd15017, 16'd48961, 16'd44335, 16'd19017, 16'd46944, 16'd33716, 16'd49437, 16'd50210, 16'd7560, 16'd58993, 16'd29201, 16'd22528, 16'd29690, 16'd44229, 16'd54837, 16'd34349, 16'd60309});
	test_expansion(128'hbe083e0c419924752c88a57d3fad1000, {16'd16203, 16'd57420, 16'd21373, 16'd16788, 16'd51683, 16'd20645, 16'd44981, 16'd15758, 16'd25731, 16'd11758, 16'd2690, 16'd63628, 16'd20598, 16'd22188, 16'd36089, 16'd23455, 16'd2467, 16'd18077, 16'd1390, 16'd32215, 16'd54997, 16'd100, 16'd20213, 16'd5549, 16'd27561, 16'd42496});
	test_expansion(128'h2a15e3fe84af13618f024bf49b072890, {16'd11364, 16'd54498, 16'd18917, 16'd53461, 16'd14268, 16'd57384, 16'd8807, 16'd31982, 16'd3396, 16'd18747, 16'd36994, 16'd38378, 16'd26413, 16'd51699, 16'd14815, 16'd20523, 16'd1723, 16'd23815, 16'd8737, 16'd10640, 16'd36399, 16'd26633, 16'd48557, 16'd18694, 16'd29165, 16'd49370});
	test_expansion(128'h947b1db5f41e25ee7e592a7e8dd6e96f, {16'd2747, 16'd35855, 16'd11729, 16'd60255, 16'd62661, 16'd28644, 16'd33137, 16'd49365, 16'd28633, 16'd32725, 16'd10931, 16'd17015, 16'd36789, 16'd18721, 16'd51007, 16'd51657, 16'd47264, 16'd62862, 16'd26178, 16'd31290, 16'd42819, 16'd50077, 16'd13928, 16'd36296, 16'd6676, 16'd50357});
	test_expansion(128'h7a1a3056dc7d1158b08d8c7fb8864ef0, {16'd7053, 16'd30035, 16'd54753, 16'd6131, 16'd41996, 16'd54740, 16'd21259, 16'd7628, 16'd4231, 16'd49769, 16'd34788, 16'd1916, 16'd61241, 16'd53220, 16'd43885, 16'd44698, 16'd64738, 16'd60199, 16'd45492, 16'd45696, 16'd42769, 16'd38613, 16'd26668, 16'd42867, 16'd9206, 16'd3981});
	test_expansion(128'hd86f46c8e1153443f9b793fb19b966d3, {16'd49525, 16'd32612, 16'd18250, 16'd53608, 16'd36043, 16'd53528, 16'd59890, 16'd28691, 16'd16851, 16'd49449, 16'd33224, 16'd26002, 16'd34486, 16'd63766, 16'd1878, 16'd44416, 16'd10955, 16'd7363, 16'd51086, 16'd44628, 16'd26603, 16'd26879, 16'd13970, 16'd46963, 16'd62798, 16'd23585});
	test_expansion(128'h47752164c0f1c4df04452d93d4135285, {16'd47844, 16'd31883, 16'd33327, 16'd27841, 16'd47885, 16'd34074, 16'd38102, 16'd48600, 16'd32672, 16'd64347, 16'd56717, 16'd41237, 16'd53152, 16'd45373, 16'd6731, 16'd55083, 16'd41780, 16'd61964, 16'd34501, 16'd48347, 16'd59199, 16'd23254, 16'd8164, 16'd43305, 16'd9498, 16'd10121});
	test_expansion(128'hb58c9133c9a1cd6346389c0822765a7d, {16'd59288, 16'd6207, 16'd9549, 16'd23556, 16'd53358, 16'd18673, 16'd19450, 16'd62086, 16'd46684, 16'd4260, 16'd63075, 16'd53395, 16'd46559, 16'd51504, 16'd65126, 16'd51011, 16'd52291, 16'd58443, 16'd13881, 16'd3549, 16'd46597, 16'd31081, 16'd38794, 16'd57598, 16'd51258, 16'd63254});
	test_expansion(128'ha74deebd5e9eb2599c5ff06721e85f93, {16'd31195, 16'd55730, 16'd25921, 16'd52810, 16'd30859, 16'd50415, 16'd39609, 16'd44932, 16'd17739, 16'd58276, 16'd22669, 16'd17137, 16'd58387, 16'd38955, 16'd39102, 16'd6213, 16'd62725, 16'd11935, 16'd10428, 16'd36813, 16'd57102, 16'd45713, 16'd4577, 16'd48540, 16'd46109, 16'd21269});
	test_expansion(128'h184405f6ae4ae274e074aec313ba443b, {16'd57902, 16'd35189, 16'd2133, 16'd51363, 16'd44637, 16'd62679, 16'd42896, 16'd8036, 16'd53405, 16'd1853, 16'd33873, 16'd20902, 16'd47640, 16'd39001, 16'd17498, 16'd63405, 16'd39697, 16'd37797, 16'd27884, 16'd39970, 16'd42743, 16'd31587, 16'd29806, 16'd48695, 16'd25742, 16'd61840});
	test_expansion(128'h8a72bb8facfa9a0f773248167e1c87ad, {16'd21960, 16'd35330, 16'd36705, 16'd3095, 16'd18389, 16'd28565, 16'd27351, 16'd7972, 16'd61460, 16'd20340, 16'd31652, 16'd7927, 16'd6365, 16'd48907, 16'd30124, 16'd63932, 16'd59985, 16'd62959, 16'd27108, 16'd1656, 16'd46856, 16'd4055, 16'd38078, 16'd38576, 16'd38518, 16'd12464});
	test_expansion(128'h57d63db4a1cdacd5a571fe06feb9259f, {16'd13538, 16'd9506, 16'd5421, 16'd38264, 16'd46312, 16'd11614, 16'd55164, 16'd3072, 16'd13846, 16'd54446, 16'd3421, 16'd28505, 16'd17584, 16'd266, 16'd13727, 16'd39237, 16'd32111, 16'd34790, 16'd28770, 16'd22680, 16'd10253, 16'd7175, 16'd8620, 16'd51476, 16'd22106, 16'd24850});
	test_expansion(128'hd6085d5ce7e0f10d1edaaf6f7e5f2e0e, {16'd16423, 16'd36974, 16'd4509, 16'd60681, 16'd21762, 16'd38125, 16'd54472, 16'd44375, 16'd42354, 16'd27712, 16'd19627, 16'd11959, 16'd55864, 16'd2714, 16'd40862, 16'd26362, 16'd2321, 16'd31698, 16'd10387, 16'd35619, 16'd40471, 16'd31541, 16'd10230, 16'd25768, 16'd252, 16'd5906});
	test_expansion(128'h4df2e5fe5f198c85398c10bd65bc2d8a, {16'd56642, 16'd27379, 16'd38159, 16'd61476, 16'd42316, 16'd30283, 16'd11323, 16'd55131, 16'd16473, 16'd59074, 16'd18575, 16'd44911, 16'd58632, 16'd43760, 16'd35826, 16'd14202, 16'd25665, 16'd57081, 16'd54855, 16'd40100, 16'd38149, 16'd36264, 16'd24186, 16'd9905, 16'd3424, 16'd21386});
	test_expansion(128'h9617d5c167b166f88c86c8893a086eb8, {16'd31253, 16'd12123, 16'd33679, 16'd35344, 16'd41455, 16'd9597, 16'd40299, 16'd29623, 16'd47632, 16'd20691, 16'd62107, 16'd35934, 16'd58511, 16'd9882, 16'd52959, 16'd22970, 16'd38687, 16'd50836, 16'd15340, 16'd11361, 16'd18743, 16'd6573, 16'd25945, 16'd43360, 16'd62034, 16'd55324});
	test_expansion(128'h367cd23916fddc74e8b8270960becd87, {16'd42972, 16'd30399, 16'd56787, 16'd65024, 16'd32530, 16'd856, 16'd31262, 16'd49233, 16'd267, 16'd8626, 16'd49461, 16'd9531, 16'd41268, 16'd43475, 16'd29698, 16'd39311, 16'd13496, 16'd52606, 16'd9523, 16'd59506, 16'd20800, 16'd12982, 16'd14078, 16'd42766, 16'd28326, 16'd64183});
	test_expansion(128'h1609019bfc7bbdac302fae9b762b47a9, {16'd49356, 16'd31154, 16'd18035, 16'd39925, 16'd22945, 16'd22122, 16'd14183, 16'd28920, 16'd26643, 16'd22725, 16'd24354, 16'd52003, 16'd48558, 16'd36992, 16'd10984, 16'd9979, 16'd44503, 16'd32247, 16'd28381, 16'd46325, 16'd58639, 16'd36067, 16'd25296, 16'd2772, 16'd51450, 16'd49941});
	test_expansion(128'hf53ebaa1ddecbd1dc424333a6ef1917c, {16'd35576, 16'd34901, 16'd58338, 16'd4907, 16'd57936, 16'd28985, 16'd2616, 16'd10590, 16'd33308, 16'd58709, 16'd7730, 16'd22220, 16'd8051, 16'd60680, 16'd2553, 16'd41463, 16'd1004, 16'd60794, 16'd59074, 16'd16279, 16'd9770, 16'd41011, 16'd7282, 16'd46018, 16'd59865, 16'd53090});
	test_expansion(128'hb3878d15df53d47b7cccbf209ffaba1b, {16'd40052, 16'd46115, 16'd15453, 16'd30905, 16'd33955, 16'd17137, 16'd63303, 16'd51558, 16'd22707, 16'd4570, 16'd33363, 16'd20943, 16'd55447, 16'd3427, 16'd6069, 16'd45535, 16'd31171, 16'd21026, 16'd55718, 16'd1772, 16'd65357, 16'd58702, 16'd52210, 16'd45982, 16'd64111, 16'd64070});
	test_expansion(128'h3a8130d7065645447e7dcfbf5a8b89ef, {16'd10937, 16'd21159, 16'd38611, 16'd9528, 16'd48931, 16'd26457, 16'd55293, 16'd5307, 16'd40153, 16'd18090, 16'd54917, 16'd62692, 16'd9690, 16'd41008, 16'd4757, 16'd22253, 16'd10797, 16'd5960, 16'd57576, 16'd34515, 16'd33056, 16'd60417, 16'd45265, 16'd42880, 16'd21141, 16'd39443});
	test_expansion(128'h07adb49e385118e4d4965e19b69606f8, {16'd357, 16'd6737, 16'd26360, 16'd12360, 16'd61635, 16'd57391, 16'd48578, 16'd25414, 16'd47146, 16'd20708, 16'd40992, 16'd16425, 16'd37564, 16'd62540, 16'd35323, 16'd17153, 16'd34851, 16'd65022, 16'd34924, 16'd23337, 16'd14407, 16'd64057, 16'd44625, 16'd50826, 16'd38009, 16'd43505});
	test_expansion(128'h5c91ab7a619c4a309d06321199acfff4, {16'd26115, 16'd15155, 16'd59125, 16'd45404, 16'd30661, 16'd27486, 16'd59984, 16'd57211, 16'd33027, 16'd18215, 16'd45594, 16'd4113, 16'd56850, 16'd37995, 16'd63927, 16'd10097, 16'd17153, 16'd44613, 16'd15486, 16'd10557, 16'd32007, 16'd37230, 16'd20180, 16'd63483, 16'd31709, 16'd36784});
	test_expansion(128'hae61e05f530ad6d3e98c3711f908d01a, {16'd47215, 16'd42806, 16'd10396, 16'd22040, 16'd53987, 16'd9771, 16'd19667, 16'd51844, 16'd43865, 16'd39934, 16'd12752, 16'd62681, 16'd42412, 16'd54944, 16'd47352, 16'd7299, 16'd45210, 16'd53889, 16'd7523, 16'd49995, 16'd46745, 16'd16132, 16'd47005, 16'd13509, 16'd34256, 16'd34205});
	test_expansion(128'h148e59082152798e984c2b57a5f7439f, {16'd53118, 16'd16698, 16'd35242, 16'd13226, 16'd19745, 16'd23788, 16'd5017, 16'd26384, 16'd14992, 16'd45557, 16'd14364, 16'd2307, 16'd59789, 16'd12961, 16'd12068, 16'd56962, 16'd12523, 16'd27087, 16'd50266, 16'd18012, 16'd3530, 16'd37896, 16'd21936, 16'd41898, 16'd64754, 16'd38502});
	test_expansion(128'h97a00c8f9e53654d9645815cd4fc83b9, {16'd18779, 16'd46352, 16'd44499, 16'd13934, 16'd60494, 16'd25490, 16'd49060, 16'd37301, 16'd25445, 16'd6855, 16'd28283, 16'd6623, 16'd18608, 16'd47298, 16'd53888, 16'd61045, 16'd43157, 16'd52688, 16'd15543, 16'd12043, 16'd34387, 16'd62768, 16'd48403, 16'd19470, 16'd43905, 16'd22702});
	test_expansion(128'hd1d69875a402386ee589d61faaa83310, {16'd2304, 16'd22124, 16'd51425, 16'd11101, 16'd25233, 16'd4846, 16'd23065, 16'd9329, 16'd55544, 16'd9090, 16'd3598, 16'd27274, 16'd26719, 16'd63423, 16'd32603, 16'd48459, 16'd37452, 16'd59107, 16'd65290, 16'd24137, 16'd2058, 16'd32543, 16'd17422, 16'd6789, 16'd15770, 16'd7918});
	test_expansion(128'hd2399243bcc80a785786a5bb09169d07, {16'd55193, 16'd43285, 16'd8761, 16'd58533, 16'd27569, 16'd29569, 16'd35784, 16'd20444, 16'd40072, 16'd28169, 16'd57718, 16'd30596, 16'd16119, 16'd60349, 16'd49559, 16'd36602, 16'd15253, 16'd26514, 16'd5721, 16'd41468, 16'd28107, 16'd2774, 16'd18214, 16'd47301, 16'd45603, 16'd50986});
	test_expansion(128'h00cb116f47da077eb46b2dd8a8e1810d, {16'd28791, 16'd7269, 16'd56476, 16'd6365, 16'd20437, 16'd33144, 16'd31901, 16'd18700, 16'd61299, 16'd61758, 16'd52798, 16'd48804, 16'd61098, 16'd47023, 16'd3056, 16'd8117, 16'd50460, 16'd63590, 16'd43231, 16'd53538, 16'd3148, 16'd30054, 16'd8876, 16'd20212, 16'd8353, 16'd40271});
	test_expansion(128'h1afdc6833aa1d1afb921f9b508f61747, {16'd15513, 16'd51453, 16'd55261, 16'd57172, 16'd20346, 16'd17867, 16'd54036, 16'd48231, 16'd18444, 16'd52591, 16'd14561, 16'd35400, 16'd51609, 16'd42899, 16'd37796, 16'd5191, 16'd62805, 16'd27141, 16'd40294, 16'd12062, 16'd6030, 16'd22141, 16'd27016, 16'd4367, 16'd26088, 16'd32057});
	test_expansion(128'hcf405f67e37ee306a2538df8fb1d9686, {16'd39508, 16'd56208, 16'd34554, 16'd39723, 16'd27738, 16'd53614, 16'd60444, 16'd39747, 16'd16194, 16'd31367, 16'd24555, 16'd6035, 16'd46838, 16'd53211, 16'd64207, 16'd22678, 16'd41025, 16'd63035, 16'd6272, 16'd13702, 16'd63517, 16'd54900, 16'd30304, 16'd35761, 16'd26538, 16'd45262});
	test_expansion(128'h51d7c84a6de703451fa8153ee836b08f, {16'd4385, 16'd8316, 16'd9137, 16'd59537, 16'd48139, 16'd40760, 16'd42917, 16'd8865, 16'd16509, 16'd1754, 16'd39156, 16'd16641, 16'd40876, 16'd8383, 16'd32753, 16'd26396, 16'd23812, 16'd29377, 16'd45096, 16'd38435, 16'd30051, 16'd25563, 16'd42369, 16'd58146, 16'd15505, 16'd38550});
	test_expansion(128'h91027bee6d9e00cf832f5f32f1d40030, {16'd14747, 16'd20183, 16'd7862, 16'd60555, 16'd57481, 16'd34665, 16'd52956, 16'd32102, 16'd53198, 16'd44848, 16'd15997, 16'd10408, 16'd62015, 16'd13755, 16'd57006, 16'd52757, 16'd11746, 16'd3694, 16'd16256, 16'd37556, 16'd5365, 16'd61265, 16'd6153, 16'd61331, 16'd32184, 16'd59724});
	test_expansion(128'h205f51c0e15f98fe98aab76ac9defad2, {16'd54503, 16'd3315, 16'd52904, 16'd33117, 16'd9721, 16'd15184, 16'd11040, 16'd65408, 16'd62246, 16'd24620, 16'd16479, 16'd64485, 16'd46950, 16'd50619, 16'd26543, 16'd43962, 16'd32022, 16'd63518, 16'd46014, 16'd17496, 16'd42061, 16'd14756, 16'd52254, 16'd65138, 16'd60842, 16'd57035});
	test_expansion(128'h49f6557f655b1f0539a357efb81e80dd, {16'd42896, 16'd11871, 16'd54275, 16'd23646, 16'd45756, 16'd7197, 16'd45754, 16'd26692, 16'd1675, 16'd40776, 16'd35585, 16'd43372, 16'd25515, 16'd18345, 16'd53750, 16'd12022, 16'd49204, 16'd36752, 16'd58231, 16'd38006, 16'd2117, 16'd63197, 16'd15273, 16'd27729, 16'd34613, 16'd54061});
	test_expansion(128'h4be47e864940fd89ee0ef2fa1bceab35, {16'd51843, 16'd52333, 16'd342, 16'd7333, 16'd56293, 16'd14714, 16'd34548, 16'd35972, 16'd39162, 16'd5283, 16'd13862, 16'd39200, 16'd38046, 16'd42866, 16'd25992, 16'd45086, 16'd1681, 16'd7525, 16'd40871, 16'd25194, 16'd43374, 16'd36964, 16'd30768, 16'd52298, 16'd33619, 16'd54756});
	test_expansion(128'h52a5618da37974c73130e3602ca5dddf, {16'd7953, 16'd3522, 16'd39194, 16'd14227, 16'd60257, 16'd12925, 16'd57628, 16'd25903, 16'd31111, 16'd30168, 16'd60697, 16'd47851, 16'd31263, 16'd28211, 16'd35851, 16'd47375, 16'd9195, 16'd54146, 16'd437, 16'd58776, 16'd64886, 16'd55513, 16'd25480, 16'd14796, 16'd13904, 16'd51893});
	test_expansion(128'he90f75b8e58a3635a155d4581f4487aa, {16'd48675, 16'd59393, 16'd1406, 16'd50306, 16'd56355, 16'd23863, 16'd5276, 16'd26541, 16'd50051, 16'd62112, 16'd33002, 16'd63670, 16'd7130, 16'd12132, 16'd64087, 16'd9994, 16'd33557, 16'd28557, 16'd61407, 16'd42540, 16'd37095, 16'd16479, 16'd28538, 16'd39104, 16'd49304, 16'd41390});
	test_expansion(128'he364c5a65b529080c6962365052788c5, {16'd34593, 16'd43138, 16'd47764, 16'd2133, 16'd20950, 16'd28228, 16'd17693, 16'd59838, 16'd4707, 16'd35512, 16'd24889, 16'd32348, 16'd23872, 16'd63207, 16'd30599, 16'd5667, 16'd17130, 16'd18500, 16'd25041, 16'd12492, 16'd5731, 16'd31137, 16'd31895, 16'd17577, 16'd46437, 16'd61623});
	test_expansion(128'h07eb228608de771718b783098a3e6de9, {16'd199, 16'd16709, 16'd6984, 16'd40676, 16'd52593, 16'd51708, 16'd44573, 16'd13986, 16'd30346, 16'd43491, 16'd7380, 16'd47549, 16'd12800, 16'd56366, 16'd2599, 16'd58231, 16'd57363, 16'd14842, 16'd4625, 16'd38283, 16'd17159, 16'd16789, 16'd24640, 16'd29234, 16'd1605, 16'd11651});
	test_expansion(128'ha61ccb430f349b3a2ce9d2f41b5651fe, {16'd24696, 16'd37276, 16'd6988, 16'd31355, 16'd6979, 16'd817, 16'd12024, 16'd4220, 16'd47726, 16'd25487, 16'd21027, 16'd16955, 16'd59385, 16'd52122, 16'd27997, 16'd40119, 16'd21397, 16'd40024, 16'd12099, 16'd42321, 16'd41046, 16'd8902, 16'd22066, 16'd30509, 16'd37898, 16'd27298});
	test_expansion(128'h1d52abe5e8ca2acc1170e0a1b7e773b5, {16'd34383, 16'd338, 16'd8377, 16'd51590, 16'd27981, 16'd15602, 16'd19613, 16'd52706, 16'd39899, 16'd28340, 16'd10041, 16'd53307, 16'd55194, 16'd65483, 16'd61746, 16'd31311, 16'd17008, 16'd8906, 16'd30527, 16'd24948, 16'd17146, 16'd50099, 16'd41502, 16'd57394, 16'd33007, 16'd15629});
	test_expansion(128'hb6b8c791e71a05c5ff99006ab94cadd6, {16'd44081, 16'd61404, 16'd26097, 16'd48320, 16'd23145, 16'd63726, 16'd25701, 16'd45952, 16'd6774, 16'd32415, 16'd19601, 16'd52797, 16'd3691, 16'd35968, 16'd15032, 16'd64491, 16'd27244, 16'd39587, 16'd37423, 16'd20347, 16'd3553, 16'd42685, 16'd9424, 16'd33028, 16'd44602, 16'd33044});
	test_expansion(128'hca8ff508ce41f318938183574c307d68, {16'd48827, 16'd32592, 16'd64776, 16'd27433, 16'd58170, 16'd61519, 16'd65432, 16'd8378, 16'd26775, 16'd55044, 16'd12449, 16'd36728, 16'd43267, 16'd27262, 16'd21577, 16'd58475, 16'd45989, 16'd10519, 16'd11167, 16'd19572, 16'd65224, 16'd11955, 16'd1714, 16'd1798, 16'd1742, 16'd6527});
	test_expansion(128'hc72d1f1254460ea23ceb9dc72adc19d4, {16'd54748, 16'd19529, 16'd45324, 16'd52259, 16'd7514, 16'd21574, 16'd4416, 16'd33306, 16'd65379, 16'd12675, 16'd26841, 16'd57017, 16'd40747, 16'd23950, 16'd64957, 16'd56661, 16'd28105, 16'd53136, 16'd45312, 16'd50056, 16'd390, 16'd11672, 16'd48928, 16'd35816, 16'd46824, 16'd11443});
	test_expansion(128'hb1edfee3cf6a7f802b55237771ffef93, {16'd1138, 16'd56032, 16'd1344, 16'd17885, 16'd51581, 16'd48773, 16'd20428, 16'd44077, 16'd17963, 16'd21907, 16'd51052, 16'd23114, 16'd2204, 16'd49541, 16'd37866, 16'd39702, 16'd19222, 16'd13659, 16'd23953, 16'd9106, 16'd5597, 16'd46652, 16'd13939, 16'd59174, 16'd65090, 16'd50704});
	test_expansion(128'h435e7b024ab01a31fe6f65b5ae0caa68, {16'd15514, 16'd48542, 16'd63269, 16'd51666, 16'd21776, 16'd55546, 16'd65046, 16'd64028, 16'd34748, 16'd17680, 16'd58566, 16'd29017, 16'd50885, 16'd27733, 16'd23832, 16'd6941, 16'd64608, 16'd64660, 16'd56720, 16'd11824, 16'd19973, 16'd2642, 16'd59135, 16'd8011, 16'd35151, 16'd40632});
	test_expansion(128'h2e51cee918658fd5d2acf049c35830f0, {16'd40719, 16'd13787, 16'd37137, 16'd30637, 16'd47617, 16'd2813, 16'd57533, 16'd37786, 16'd55650, 16'd33810, 16'd31259, 16'd22463, 16'd2912, 16'd13325, 16'd25406, 16'd56358, 16'd42964, 16'd57582, 16'd39030, 16'd58351, 16'd6290, 16'd31395, 16'd55179, 16'd63503, 16'd9056, 16'd53935});
	test_expansion(128'he183ca4aafa9d7ecccbd83284490b42e, {16'd46114, 16'd16661, 16'd21241, 16'd8267, 16'd50275, 16'd49860, 16'd31792, 16'd38771, 16'd27194, 16'd26206, 16'd53349, 16'd23112, 16'd51965, 16'd27892, 16'd10199, 16'd63297, 16'd14047, 16'd39091, 16'd42670, 16'd3503, 16'd64332, 16'd58321, 16'd48281, 16'd22395, 16'd54913, 16'd16948});
	test_expansion(128'h9a50c0e95167cd9e1c8d7b9e315a9e01, {16'd62400, 16'd11481, 16'd1290, 16'd52327, 16'd6899, 16'd20254, 16'd3285, 16'd41599, 16'd59636, 16'd53887, 16'd50093, 16'd11360, 16'd58006, 16'd1016, 16'd47027, 16'd48530, 16'd58632, 16'd38416, 16'd26512, 16'd15881, 16'd57993, 16'd54731, 16'd53915, 16'd37021, 16'd12410, 16'd12928});
	test_expansion(128'h40f1aa089a604a4d9975bf5c25906f59, {16'd22363, 16'd48906, 16'd59805, 16'd8915, 16'd17791, 16'd5979, 16'd40736, 16'd7285, 16'd10539, 16'd43636, 16'd10866, 16'd24308, 16'd35876, 16'd2752, 16'd3525, 16'd14428, 16'd23919, 16'd58825, 16'd57122, 16'd41439, 16'd15643, 16'd60213, 16'd61401, 16'd3274, 16'd30136, 16'd47167});
	test_expansion(128'ha7e1fc2e5c0184c743478b4a790562e6, {16'd57066, 16'd32903, 16'd47130, 16'd11677, 16'd12362, 16'd16501, 16'd35160, 16'd13378, 16'd62668, 16'd46606, 16'd57789, 16'd30419, 16'd658, 16'd57648, 16'd56705, 16'd60656, 16'd53006, 16'd42559, 16'd12912, 16'd57508, 16'd64141, 16'd14365, 16'd54092, 16'd32344, 16'd15149, 16'd58731});
	test_expansion(128'hbc8672901f01e2040c63693cba526170, {16'd32688, 16'd65327, 16'd10601, 16'd25547, 16'd56055, 16'd16568, 16'd12129, 16'd41151, 16'd16641, 16'd38581, 16'd34266, 16'd9899, 16'd44086, 16'd22357, 16'd24789, 16'd61041, 16'd47946, 16'd38866, 16'd58805, 16'd15969, 16'd55610, 16'd29324, 16'd12755, 16'd49081, 16'd33676, 16'd5426});
	test_expansion(128'h8f0d4836e77189a8102fd97e2b085328, {16'd16408, 16'd59236, 16'd53524, 16'd40365, 16'd56464, 16'd5966, 16'd15982, 16'd61609, 16'd1988, 16'd15348, 16'd9188, 16'd50419, 16'd19850, 16'd45035, 16'd13726, 16'd59574, 16'd1529, 16'd2659, 16'd28749, 16'd17154, 16'd20052, 16'd52967, 16'd43321, 16'd47297, 16'd30578, 16'd38313});
	test_expansion(128'h7e1f51f0e73d9da4d24d5f8480d8bc39, {16'd2174, 16'd25461, 16'd30420, 16'd42810, 16'd54254, 16'd54972, 16'd60187, 16'd4298, 16'd43429, 16'd34143, 16'd55453, 16'd41624, 16'd36047, 16'd18232, 16'd5305, 16'd17793, 16'd33320, 16'd50393, 16'd1053, 16'd31451, 16'd42594, 16'd36430, 16'd26584, 16'd29876, 16'd26238, 16'd45133});
	test_expansion(128'he85b32af103ebd1aeee408e187a3feb8, {16'd21384, 16'd60647, 16'd50854, 16'd42252, 16'd59221, 16'd59171, 16'd25848, 16'd25227, 16'd54450, 16'd46051, 16'd827, 16'd5632, 16'd21489, 16'd18698, 16'd29251, 16'd1044, 16'd58443, 16'd42805, 16'd13183, 16'd43651, 16'd17757, 16'd27022, 16'd40652, 16'd50752, 16'd10522, 16'd17747});
	test_expansion(128'ha7125cbf2f92abd2f427431d9696842e, {16'd32378, 16'd24897, 16'd1204, 16'd55332, 16'd1123, 16'd42997, 16'd43968, 16'd41143, 16'd31123, 16'd51353, 16'd49651, 16'd6582, 16'd57737, 16'd12549, 16'd21093, 16'd6907, 16'd52543, 16'd52524, 16'd61846, 16'd29821, 16'd56027, 16'd456, 16'd38714, 16'd30626, 16'd45098, 16'd20674});
	test_expansion(128'hde54a1f8326d99784c60b68eb6d3148b, {16'd41702, 16'd5377, 16'd48258, 16'd64381, 16'd56819, 16'd50023, 16'd17247, 16'd47403, 16'd24859, 16'd45302, 16'd21801, 16'd13001, 16'd36949, 16'd64596, 16'd6241, 16'd3282, 16'd21235, 16'd44604, 16'd10942, 16'd617, 16'd61058, 16'd48131, 16'd49307, 16'd50118, 16'd37098, 16'd33277});
	test_expansion(128'hf4d0aa4846f9f4d66140a663ebf2deec, {16'd15790, 16'd2841, 16'd31718, 16'd21365, 16'd9636, 16'd39335, 16'd19362, 16'd57846, 16'd30277, 16'd64491, 16'd1582, 16'd6219, 16'd6606, 16'd14902, 16'd11628, 16'd63256, 16'd32903, 16'd26465, 16'd44467, 16'd32605, 16'd34541, 16'd18796, 16'd41102, 16'd2368, 16'd25113, 16'd40834});
	test_expansion(128'hbfa4056485d455b1c69f0a14a5c01ece, {16'd38583, 16'd63769, 16'd54002, 16'd17223, 16'd58240, 16'd26175, 16'd42582, 16'd13239, 16'd55329, 16'd55720, 16'd38652, 16'd53070, 16'd27756, 16'd16797, 16'd60067, 16'd7702, 16'd29571, 16'd32098, 16'd14757, 16'd2264, 16'd10901, 16'd7590, 16'd28970, 16'd10444, 16'd57965, 16'd62873});
	test_expansion(128'hf956ba8b1ea8b39a8b48f0081867fc90, {16'd63366, 16'd55751, 16'd3029, 16'd10090, 16'd34940, 16'd39851, 16'd63376, 16'd22251, 16'd26971, 16'd27322, 16'd51396, 16'd32329, 16'd45508, 16'd17400, 16'd54576, 16'd44146, 16'd2289, 16'd62170, 16'd61638, 16'd13050, 16'd13770, 16'd17063, 16'd38640, 16'd27487, 16'd12217, 16'd35970});
	test_expansion(128'h5e09dbcaa0568e0f7ba6d9048268fb57, {16'd49321, 16'd18821, 16'd55753, 16'd38558, 16'd11018, 16'd37757, 16'd60919, 16'd8416, 16'd16614, 16'd32549, 16'd825, 16'd25778, 16'd21938, 16'd34474, 16'd41756, 16'd39542, 16'd61175, 16'd12561, 16'd20520, 16'd46552, 16'd30, 16'd32443, 16'd50601, 16'd55702, 16'd20865, 16'd43986});
	test_expansion(128'h3e3ef636df916e89ec94c3e6c9330b0c, {16'd6873, 16'd41999, 16'd3009, 16'd60125, 16'd9938, 16'd45089, 16'd46321, 16'd2822, 16'd37698, 16'd50045, 16'd7339, 16'd41456, 16'd3224, 16'd38761, 16'd20255, 16'd62391, 16'd5010, 16'd52173, 16'd33188, 16'd38826, 16'd6896, 16'd40104, 16'd54667, 16'd58722, 16'd46017, 16'd27135});
	test_expansion(128'h2b038a0cbeb50c2a25be837723b0156c, {16'd62177, 16'd48097, 16'd31753, 16'd60932, 16'd18351, 16'd63595, 16'd7757, 16'd30404, 16'd16137, 16'd6897, 16'd64558, 16'd63862, 16'd57153, 16'd1204, 16'd49321, 16'd43550, 16'd56350, 16'd60945, 16'd55593, 16'd41496, 16'd47246, 16'd12229, 16'd64446, 16'd269, 16'd22019, 16'd29591});
	test_expansion(128'hddb6b74530b86f207f566b76d145a88b, {16'd50429, 16'd63160, 16'd30831, 16'd44599, 16'd24974, 16'd27603, 16'd60147, 16'd62077, 16'd48230, 16'd42745, 16'd30271, 16'd18256, 16'd18555, 16'd30956, 16'd40260, 16'd35944, 16'd33689, 16'd42676, 16'd21089, 16'd24297, 16'd31163, 16'd40801, 16'd4189, 16'd11521, 16'd28590, 16'd41217});
	test_expansion(128'h0fc8eb82b6dd5e5fefa3ccfe27858461, {16'd46599, 16'd26507, 16'd45106, 16'd12681, 16'd13819, 16'd51677, 16'd24197, 16'd15225, 16'd1680, 16'd9911, 16'd16372, 16'd35470, 16'd18586, 16'd62907, 16'd29938, 16'd8065, 16'd34401, 16'd59670, 16'd8465, 16'd40959, 16'd11247, 16'd13378, 16'd38461, 16'd21920, 16'd20219, 16'd5499});
	test_expansion(128'hb39b7a3b1d45c89b99a6b2465e8310f2, {16'd48835, 16'd29726, 16'd55389, 16'd6900, 16'd46935, 16'd24846, 16'd30693, 16'd46562, 16'd29518, 16'd53447, 16'd11870, 16'd41038, 16'd56944, 16'd29128, 16'd64385, 16'd38787, 16'd1668, 16'd41702, 16'd51551, 16'd30408, 16'd36159, 16'd26563, 16'd19392, 16'd17218, 16'd36284, 16'd55870});
	test_expansion(128'hefd119842d312f09252b13f6b118ef9b, {16'd55572, 16'd37140, 16'd62876, 16'd42582, 16'd50954, 16'd30454, 16'd25118, 16'd47707, 16'd56136, 16'd45525, 16'd32135, 16'd3259, 16'd46881, 16'd59268, 16'd30869, 16'd4195, 16'd31077, 16'd48117, 16'd41731, 16'd12908, 16'd53498, 16'd3608, 16'd53540, 16'd54026, 16'd56217, 16'd48828});
	test_expansion(128'h609cf8da206a6f0c5fa786fc2fc684d5, {16'd57045, 16'd13813, 16'd32889, 16'd24192, 16'd3121, 16'd62506, 16'd39015, 16'd50436, 16'd35955, 16'd8801, 16'd65021, 16'd46063, 16'd11408, 16'd10010, 16'd26331, 16'd63578, 16'd13626, 16'd3510, 16'd47539, 16'd7171, 16'd21643, 16'd33444, 16'd16241, 16'd58844, 16'd9762, 16'd24605});
	test_expansion(128'h26ff9129c7e30c12c4d0b4ae5146d388, {16'd50202, 16'd46319, 16'd19054, 16'd53269, 16'd8576, 16'd59649, 16'd21426, 16'd2693, 16'd18761, 16'd60190, 16'd21674, 16'd40356, 16'd6070, 16'd58092, 16'd60391, 16'd56243, 16'd31861, 16'd42015, 16'd58378, 16'd60736, 16'd21608, 16'd53613, 16'd26697, 16'd41536, 16'd43062, 16'd2599});
	test_expansion(128'hab20f455f7f89672e8cd09fe189c9f41, {16'd26522, 16'd37104, 16'd37145, 16'd3310, 16'd25608, 16'd3128, 16'd29017, 16'd29178, 16'd26620, 16'd46829, 16'd28091, 16'd19317, 16'd6119, 16'd57459, 16'd46080, 16'd34369, 16'd8063, 16'd57886, 16'd14351, 16'd15959, 16'd65246, 16'd31151, 16'd19072, 16'd14837, 16'd11828, 16'd25752});
	test_expansion(128'h60aa729b776d6f47467e342a5340a432, {16'd23726, 16'd12289, 16'd53515, 16'd36225, 16'd20182, 16'd33981, 16'd39754, 16'd14882, 16'd59796, 16'd61762, 16'd36059, 16'd6056, 16'd54436, 16'd1436, 16'd38433, 16'd56011, 16'd18677, 16'd56358, 16'd22789, 16'd4504, 16'd33381, 16'd30829, 16'd17373, 16'd33255, 16'd16009, 16'd19324});
	test_expansion(128'h56475f1d844c67989f27a01a4b2f93a0, {16'd18968, 16'd54712, 16'd17874, 16'd31731, 16'd33483, 16'd18824, 16'd9359, 16'd19545, 16'd56551, 16'd14454, 16'd14945, 16'd37672, 16'd13, 16'd61401, 16'd33712, 16'd49376, 16'd5419, 16'd54579, 16'd34344, 16'd14364, 16'd32993, 16'd42924, 16'd40362, 16'd42823, 16'd44409, 16'd29082});
	test_expansion(128'hcdc8a28911a27b66de0234ff1a4729a2, {16'd37388, 16'd47521, 16'd24698, 16'd48303, 16'd3048, 16'd32626, 16'd48006, 16'd6312, 16'd13266, 16'd541, 16'd45781, 16'd22010, 16'd46677, 16'd25671, 16'd14840, 16'd10123, 16'd3257, 16'd55330, 16'd43954, 16'd16968, 16'd53810, 16'd56513, 16'd48132, 16'd50955, 16'd14570, 16'd42629});
	test_expansion(128'h52746fc4d78798d5a221c3c6a37e4293, {16'd28499, 16'd26310, 16'd47654, 16'd18956, 16'd10050, 16'd47484, 16'd52133, 16'd6626, 16'd54855, 16'd9416, 16'd41806, 16'd54018, 16'd56341, 16'd24749, 16'd51302, 16'd8828, 16'd61524, 16'd24905, 16'd11801, 16'd4271, 16'd4993, 16'd28679, 16'd57038, 16'd17228, 16'd32941, 16'd14034});
	test_expansion(128'h01ae0be1411335989f3d8b3e75fc0909, {16'd33293, 16'd59563, 16'd23323, 16'd24693, 16'd55168, 16'd28040, 16'd1877, 16'd11090, 16'd36326, 16'd14886, 16'd29660, 16'd62615, 16'd29359, 16'd60384, 16'd18358, 16'd43398, 16'd26652, 16'd4120, 16'd55263, 16'd62116, 16'd39019, 16'd10258, 16'd39340, 16'd6718, 16'd37721, 16'd57130});
	test_expansion(128'he13e3cef38d22a8afdc2a7afc9993226, {16'd62004, 16'd6015, 16'd26648, 16'd31366, 16'd45868, 16'd44323, 16'd55472, 16'd50192, 16'd38977, 16'd49403, 16'd35716, 16'd12467, 16'd43114, 16'd13521, 16'd5273, 16'd43741, 16'd13238, 16'd61591, 16'd9801, 16'd61059, 16'd127, 16'd56750, 16'd61861, 16'd51766, 16'd35938, 16'd42437});
	test_expansion(128'hce516c5f6117106ee85ca8e8cd946454, {16'd30253, 16'd54557, 16'd19959, 16'd65170, 16'd52228, 16'd64781, 16'd56147, 16'd49224, 16'd37953, 16'd6843, 16'd53451, 16'd17851, 16'd63904, 16'd43179, 16'd37940, 16'd28301, 16'd60412, 16'd9904, 16'd9707, 16'd28643, 16'd3545, 16'd49165, 16'd5537, 16'd13850, 16'd26550, 16'd43053});
	test_expansion(128'ha77d1f8b89a7e08df350fc5c930ccb8e, {16'd18036, 16'd12704, 16'd12763, 16'd3117, 16'd17925, 16'd54304, 16'd36366, 16'd17571, 16'd11082, 16'd24776, 16'd8604, 16'd45832, 16'd32589, 16'd18932, 16'd38726, 16'd4224, 16'd44798, 16'd1675, 16'd35191, 16'd35958, 16'd40787, 16'd59786, 16'd34532, 16'd36884, 16'd16160, 16'd37633});
	test_expansion(128'hccc8f07fa808db76eee38e6d3780cac2, {16'd53121, 16'd24034, 16'd14485, 16'd53757, 16'd7054, 16'd11115, 16'd33332, 16'd27699, 16'd21535, 16'd23313, 16'd50542, 16'd10377, 16'd50474, 16'd36040, 16'd22559, 16'd21979, 16'd18095, 16'd27210, 16'd61979, 16'd14105, 16'd20318, 16'd59560, 16'd44777, 16'd51825, 16'd38091, 16'd65123});
	test_expansion(128'hdc1d90665139cf25cf4fc1c7928065ec, {16'd46170, 16'd26089, 16'd44166, 16'd36628, 16'd7567, 16'd40688, 16'd52553, 16'd3912, 16'd48670, 16'd13329, 16'd63272, 16'd9362, 16'd44901, 16'd42685, 16'd60971, 16'd5290, 16'd47780, 16'd58472, 16'd2825, 16'd56247, 16'd20048, 16'd32974, 16'd58684, 16'd44646, 16'd30593, 16'd7345});
	test_expansion(128'hb4756821dda151b38517f0616007997d, {16'd36209, 16'd13346, 16'd59934, 16'd54720, 16'd12544, 16'd464, 16'd36969, 16'd14966, 16'd18583, 16'd50833, 16'd1091, 16'd17892, 16'd54393, 16'd32763, 16'd37713, 16'd40878, 16'd61370, 16'd30750, 16'd36063, 16'd29125, 16'd56893, 16'd9798, 16'd15674, 16'd57594, 16'd47169, 16'd51499});
	test_expansion(128'hd1b5e6f50feeb99084d571f48666d95c, {16'd45808, 16'd47018, 16'd13623, 16'd51667, 16'd11897, 16'd19049, 16'd35299, 16'd41776, 16'd35778, 16'd40746, 16'd36731, 16'd27582, 16'd59830, 16'd23025, 16'd21332, 16'd20808, 16'd14507, 16'd40077, 16'd61644, 16'd62198, 16'd59584, 16'd2710, 16'd30455, 16'd30078, 16'd44624, 16'd51835});
	test_expansion(128'h1a02f3cbaa8981c6539f2bdccf64c045, {16'd35805, 16'd63411, 16'd3859, 16'd20195, 16'd44488, 16'd24105, 16'd40933, 16'd45991, 16'd18094, 16'd34531, 16'd18633, 16'd51313, 16'd16980, 16'd11381, 16'd46397, 16'd32772, 16'd31718, 16'd45159, 16'd29004, 16'd31280, 16'd17982, 16'd54465, 16'd6530, 16'd56646, 16'd36008, 16'd15129});
	test_expansion(128'hb2e1985b341d115c543c1003dc922deb, {16'd64708, 16'd27919, 16'd54917, 16'd25438, 16'd41939, 16'd19317, 16'd22703, 16'd49289, 16'd5431, 16'd53622, 16'd31754, 16'd47896, 16'd58015, 16'd144, 16'd35806, 16'd42373, 16'd47331, 16'd48423, 16'd11747, 16'd61831, 16'd48784, 16'd31684, 16'd41459, 16'd21833, 16'd16128, 16'd25672});
	test_expansion(128'hd52f509599ab063d4393e75bb8cb8c81, {16'd56981, 16'd55681, 16'd61186, 16'd54609, 16'd39933, 16'd28400, 16'd51752, 16'd42610, 16'd21076, 16'd11408, 16'd27086, 16'd50161, 16'd17667, 16'd18308, 16'd53566, 16'd3072, 16'd11371, 16'd63490, 16'd61162, 16'd62410, 16'd62286, 16'd32321, 16'd37751, 16'd60691, 16'd64955, 16'd7042});
	test_expansion(128'h04adc226dae563fadf422fda7674959c, {16'd33989, 16'd18662, 16'd52932, 16'd48835, 16'd46829, 16'd62363, 16'd58670, 16'd1964, 16'd46805, 16'd288, 16'd60442, 16'd44426, 16'd59519, 16'd23349, 16'd54588, 16'd53243, 16'd6485, 16'd45157, 16'd11907, 16'd49705, 16'd1460, 16'd53304, 16'd24552, 16'd52354, 16'd54778, 16'd33618});
	test_expansion(128'h8c2a8375a00bee90f36312dd1fcc9c4a, {16'd57204, 16'd29195, 16'd40051, 16'd10820, 16'd36580, 16'd1647, 16'd52095, 16'd59980, 16'd35991, 16'd32874, 16'd59910, 16'd59726, 16'd55361, 16'd14817, 16'd17921, 16'd20255, 16'd38234, 16'd48918, 16'd16492, 16'd34507, 16'd8472, 16'd60361, 16'd14438, 16'd35633, 16'd30253, 16'd63679});
	test_expansion(128'h2d71e5bd0bef99a89abb8fd766079279, {16'd3653, 16'd16338, 16'd51848, 16'd34813, 16'd49632, 16'd35417, 16'd372, 16'd47364, 16'd43041, 16'd38115, 16'd46301, 16'd59623, 16'd10738, 16'd53384, 16'd25914, 16'd34053, 16'd58625, 16'd6718, 16'd45923, 16'd59752, 16'd22832, 16'd18924, 16'd24143, 16'd14912, 16'd23335, 16'd61095});
	test_expansion(128'h5f8b04f694b8e5d5301e636a6cbbb704, {16'd10111, 16'd39513, 16'd32337, 16'd55429, 16'd25825, 16'd53782, 16'd16581, 16'd31175, 16'd34664, 16'd6109, 16'd39372, 16'd12711, 16'd34497, 16'd9742, 16'd44694, 16'd5021, 16'd7738, 16'd59486, 16'd14143, 16'd60073, 16'd929, 16'd62795, 16'd5893, 16'd9795, 16'd53948, 16'd41822});
	test_expansion(128'hfed35e879c29995b54611e85b4cec87c, {16'd48180, 16'd57455, 16'd39443, 16'd36738, 16'd26908, 16'd41453, 16'd17953, 16'd2792, 16'd39855, 16'd25772, 16'd8242, 16'd3848, 16'd26351, 16'd42224, 16'd331, 16'd14976, 16'd65494, 16'd12981, 16'd20900, 16'd26575, 16'd13175, 16'd1410, 16'd2417, 16'd2333, 16'd25018, 16'd40341});
	test_expansion(128'h5e9dab56e4760dab4393e0bdb3d72a8a, {16'd58980, 16'd47408, 16'd64930, 16'd9061, 16'd14130, 16'd36006, 16'd42429, 16'd3042, 16'd36465, 16'd32590, 16'd58599, 16'd41553, 16'd28611, 16'd21238, 16'd1114, 16'd51323, 16'd56873, 16'd15292, 16'd2501, 16'd27510, 16'd9515, 16'd23721, 16'd54127, 16'd52709, 16'd46322, 16'd36211});
	test_expansion(128'hc80e3873053f87d6114674b4812f279a, {16'd45285, 16'd64048, 16'd49531, 16'd40273, 16'd54390, 16'd53757, 16'd37328, 16'd60986, 16'd57663, 16'd56044, 16'd28549, 16'd10959, 16'd25488, 16'd6657, 16'd51844, 16'd59318, 16'd63688, 16'd149, 16'd15458, 16'd32785, 16'd36773, 16'd11441, 16'd7078, 16'd29308, 16'd704, 16'd503});
	test_expansion(128'haaa5819d7f6d713523e870ec111d7eaa, {16'd60021, 16'd44044, 16'd13461, 16'd45720, 16'd5461, 16'd33222, 16'd49136, 16'd24609, 16'd186, 16'd13083, 16'd12097, 16'd48872, 16'd27209, 16'd39358, 16'd63321, 16'd50588, 16'd26845, 16'd25309, 16'd49428, 16'd63420, 16'd47497, 16'd26720, 16'd2034, 16'd56119, 16'd15225, 16'd27836});
	test_expansion(128'h99322460ba77ef3bf1b73f36aadd4be0, {16'd33168, 16'd35070, 16'd47521, 16'd26929, 16'd3668, 16'd62461, 16'd49440, 16'd31030, 16'd98, 16'd22522, 16'd18104, 16'd47671, 16'd58582, 16'd45683, 16'd60738, 16'd48686, 16'd50020, 16'd59838, 16'd12518, 16'd40337, 16'd36462, 16'd8684, 16'd7374, 16'd14286, 16'd32532, 16'd19375});
	test_expansion(128'h64feb5645586db395e6d63a617ef4989, {16'd201, 16'd44534, 16'd35045, 16'd60263, 16'd49988, 16'd41323, 16'd25843, 16'd49891, 16'd10697, 16'd7478, 16'd37802, 16'd52154, 16'd48577, 16'd62433, 16'd40626, 16'd56009, 16'd30919, 16'd47736, 16'd38102, 16'd44368, 16'd660, 16'd6060, 16'd9287, 16'd61050, 16'd46222, 16'd48248});
	test_expansion(128'h47eca6483f088966f61a7da877473cfc, {16'd64680, 16'd62107, 16'd42690, 16'd43297, 16'd6998, 16'd63152, 16'd18323, 16'd25769, 16'd40692, 16'd23507, 16'd13414, 16'd33921, 16'd40915, 16'd3376, 16'd37840, 16'd58770, 16'd5123, 16'd6088, 16'd55602, 16'd49835, 16'd10651, 16'd31313, 16'd64916, 16'd15962, 16'd5830, 16'd2391});
	test_expansion(128'hd603b16cfe7168f0c0a738cd00e0c1bb, {16'd46366, 16'd32847, 16'd54762, 16'd9016, 16'd42396, 16'd52056, 16'd21362, 16'd50008, 16'd13722, 16'd9352, 16'd7459, 16'd51949, 16'd14030, 16'd55100, 16'd23656, 16'd1173, 16'd3181, 16'd31043, 16'd8459, 16'd59095, 16'd53137, 16'd59399, 16'd15463, 16'd55842, 16'd56175, 16'd58460});
	test_expansion(128'h97d224178e001df362e95dfc5fe158a5, {16'd40113, 16'd63194, 16'd52572, 16'd20398, 16'd9565, 16'd56670, 16'd42816, 16'd857, 16'd26956, 16'd2886, 16'd10572, 16'd60829, 16'd61913, 16'd58657, 16'd39383, 16'd39029, 16'd21145, 16'd15941, 16'd61849, 16'd21068, 16'd2462, 16'd30622, 16'd9012, 16'd15695, 16'd12545, 16'd1453});
	test_expansion(128'he320e0a5c7f0f67167fc074969a7ff0e, {16'd16000, 16'd1354, 16'd1524, 16'd34639, 16'd10985, 16'd26555, 16'd27356, 16'd34876, 16'd38272, 16'd21160, 16'd563, 16'd64852, 16'd44311, 16'd8690, 16'd11061, 16'd30363, 16'd39592, 16'd20655, 16'd63506, 16'd13001, 16'd2513, 16'd28804, 16'd49750, 16'd55089, 16'd5562, 16'd3879});
	test_expansion(128'he99384daf1e5be46d62751d9a09f5989, {16'd60716, 16'd61649, 16'd60636, 16'd3024, 16'd61472, 16'd21399, 16'd15792, 16'd8806, 16'd43125, 16'd39229, 16'd15304, 16'd18313, 16'd28501, 16'd54859, 16'd6409, 16'd5290, 16'd4315, 16'd43545, 16'd11301, 16'd23054, 16'd51668, 16'd52265, 16'd14081, 16'd1541, 16'd41484, 16'd50664});
	test_expansion(128'h85550b48e3f1fff9108cdbf1856e70e3, {16'd16772, 16'd54396, 16'd4994, 16'd58341, 16'd16123, 16'd490, 16'd56806, 16'd26977, 16'd18099, 16'd13950, 16'd38730, 16'd58921, 16'd17405, 16'd47191, 16'd14931, 16'd58067, 16'd52877, 16'd65297, 16'd65331, 16'd53593, 16'd56057, 16'd43294, 16'd51120, 16'd19170, 16'd65136, 16'd39089});
	test_expansion(128'hac34c38d1b646b25065c58ee58bcb0db, {16'd54842, 16'd47690, 16'd19851, 16'd59293, 16'd12653, 16'd33918, 16'd30904, 16'd60430, 16'd5158, 16'd64172, 16'd2270, 16'd33208, 16'd16774, 16'd55466, 16'd56017, 16'd46214, 16'd43920, 16'd47236, 16'd18308, 16'd59862, 16'd9120, 16'd2880, 16'd45957, 16'd15080, 16'd59541, 16'd34142});
	test_expansion(128'h077279cef15380e74ca6a259b620e313, {16'd52022, 16'd34621, 16'd62812, 16'd35264, 16'd5994, 16'd46563, 16'd23348, 16'd36346, 16'd21925, 16'd9722, 16'd39815, 16'd53673, 16'd33544, 16'd9313, 16'd15592, 16'd57443, 16'd19146, 16'd65099, 16'd35749, 16'd35453, 16'd41229, 16'd8193, 16'd10987, 16'd20360, 16'd49089, 16'd64943});
	test_expansion(128'h610516bd5106ee9c008821fa96f2bc88, {16'd18783, 16'd11670, 16'd54145, 16'd24967, 16'd6875, 16'd52038, 16'd60088, 16'd8215, 16'd62707, 16'd58398, 16'd14107, 16'd2226, 16'd42250, 16'd48721, 16'd37821, 16'd35782, 16'd38145, 16'd39355, 16'd32744, 16'd38432, 16'd28795, 16'd48702, 16'd21829, 16'd11622, 16'd32291, 16'd30180});
	test_expansion(128'hd8d733fb07ba04089b6c44361c0f5d92, {16'd24216, 16'd21719, 16'd13673, 16'd11363, 16'd26139, 16'd34512, 16'd40280, 16'd7655, 16'd3881, 16'd11046, 16'd32418, 16'd41915, 16'd19348, 16'd12317, 16'd57523, 16'd31007, 16'd16752, 16'd51000, 16'd43280, 16'd59524, 16'd30631, 16'd24714, 16'd35017, 16'd29746, 16'd22184, 16'd5934});
	test_expansion(128'h5df4f6880b2dfaa28f0172c7f76af796, {16'd3781, 16'd9915, 16'd30616, 16'd62889, 16'd23531, 16'd47900, 16'd3486, 16'd18749, 16'd54811, 16'd59359, 16'd61098, 16'd27708, 16'd49686, 16'd40383, 16'd59068, 16'd7578, 16'd35349, 16'd3378, 16'd9726, 16'd46183, 16'd3971, 16'd65004, 16'd13656, 16'd11373, 16'd5328, 16'd65513});
	test_expansion(128'h0e36c6c0e88897af360644a039ff9868, {16'd64377, 16'd44755, 16'd22444, 16'd2964, 16'd31213, 16'd980, 16'd65063, 16'd24204, 16'd4942, 16'd4116, 16'd30642, 16'd20084, 16'd14598, 16'd6547, 16'd52602, 16'd32529, 16'd32013, 16'd58339, 16'd47883, 16'd38456, 16'd46463, 16'd61949, 16'd30708, 16'd8983, 16'd24620, 16'd34785});
	test_expansion(128'hbdd5149f7d681eb95270353fb800f1cf, {16'd16120, 16'd58701, 16'd46260, 16'd35423, 16'd17947, 16'd2651, 16'd39768, 16'd41095, 16'd5850, 16'd58747, 16'd23664, 16'd25413, 16'd63823, 16'd31789, 16'd20608, 16'd51892, 16'd43891, 16'd53120, 16'd9834, 16'd61195, 16'd49782, 16'd44932, 16'd43865, 16'd1700, 16'd23913, 16'd52930});
	test_expansion(128'h9f87ab633e4a7ac743bf2b384a878ff2, {16'd58059, 16'd59340, 16'd36340, 16'd37875, 16'd51705, 16'd35734, 16'd2653, 16'd19067, 16'd59354, 16'd63349, 16'd43605, 16'd46876, 16'd61188, 16'd62791, 16'd42467, 16'd64785, 16'd38746, 16'd35934, 16'd1398, 16'd53083, 16'd9719, 16'd22295, 16'd31213, 16'd17310, 16'd44680, 16'd50803});
	test_expansion(128'hcc8853a3ad22916648d54d22128692e4, {16'd8496, 16'd35627, 16'd39343, 16'd3134, 16'd36961, 16'd53515, 16'd5183, 16'd41197, 16'd1076, 16'd49348, 16'd60283, 16'd61394, 16'd6196, 16'd60554, 16'd17090, 16'd17968, 16'd12903, 16'd24991, 16'd48737, 16'd60805, 16'd36851, 16'd63114, 16'd43157, 16'd22243, 16'd14022, 16'd13125});
	test_expansion(128'h5d26245359133b403c2d7421afe86e29, {16'd45335, 16'd7602, 16'd29585, 16'd13511, 16'd39084, 16'd3991, 16'd2359, 16'd27726, 16'd62230, 16'd48310, 16'd6882, 16'd5310, 16'd2615, 16'd43366, 16'd15581, 16'd39712, 16'd28675, 16'd50734, 16'd64433, 16'd16191, 16'd1875, 16'd27716, 16'd55980, 16'd32651, 16'd45791, 16'd57252});
	test_expansion(128'h23aad5364d8a450d3a62b47537528824, {16'd64956, 16'd18457, 16'd54865, 16'd49951, 16'd34020, 16'd36766, 16'd45808, 16'd9395, 16'd23018, 16'd20189, 16'd7782, 16'd46007, 16'd41502, 16'd26713, 16'd12773, 16'd53882, 16'd26438, 16'd58572, 16'd58291, 16'd47391, 16'd10800, 16'd29521, 16'd33790, 16'd2872, 16'd26615, 16'd17060});
	test_expansion(128'hdf6b77a1be5ca9e487223a01a9bda8ed, {16'd22031, 16'd48898, 16'd10440, 16'd38861, 16'd538, 16'd24529, 16'd51897, 16'd25644, 16'd22364, 16'd15901, 16'd15501, 16'd58082, 16'd46566, 16'd27019, 16'd21826, 16'd50080, 16'd19738, 16'd53934, 16'd36025, 16'd1120, 16'd33347, 16'd32813, 16'd42221, 16'd38706, 16'd4010, 16'd3183});
	test_expansion(128'heae5d1396f4949c88f5055d0f77e69c6, {16'd6456, 16'd41684, 16'd25826, 16'd53841, 16'd16160, 16'd7132, 16'd53576, 16'd22016, 16'd64228, 16'd39202, 16'd18107, 16'd4289, 16'd17876, 16'd11860, 16'd19228, 16'd19658, 16'd2575, 16'd45979, 16'd36261, 16'd21626, 16'd63328, 16'd42365, 16'd12468, 16'd11316, 16'd55101, 16'd51518});
	test_expansion(128'h115a1f7539a510ce6ce893144b3a6ed6, {16'd50619, 16'd8489, 16'd45065, 16'd44836, 16'd20488, 16'd58708, 16'd49970, 16'd41061, 16'd16474, 16'd2022, 16'd3924, 16'd56330, 16'd23560, 16'd61944, 16'd30515, 16'd8477, 16'd49625, 16'd43265, 16'd30639, 16'd55601, 16'd10729, 16'd24770, 16'd3274, 16'd32312, 16'd39821, 16'd28418});
	test_expansion(128'hea7e978bd660dba220ef79d7fa5d607d, {16'd6117, 16'd61645, 16'd32943, 16'd50772, 16'd61633, 16'd8319, 16'd7320, 16'd35322, 16'd25405, 16'd6393, 16'd62951, 16'd18844, 16'd60271, 16'd18112, 16'd9140, 16'd37518, 16'd55452, 16'd52921, 16'd44211, 16'd17632, 16'd42553, 16'd21897, 16'd56269, 16'd21286, 16'd54982, 16'd41794});
	test_expansion(128'h6a3e6efdbe4df5dce6f8d00ae0e28591, {16'd3124, 16'd12378, 16'd60496, 16'd21700, 16'd63427, 16'd24601, 16'd4670, 16'd19325, 16'd565, 16'd40617, 16'd60897, 16'd22458, 16'd57795, 16'd64211, 16'd24269, 16'd48957, 16'd17005, 16'd39506, 16'd30721, 16'd20494, 16'd3066, 16'd20485, 16'd64331, 16'd13839, 16'd35724, 16'd10399});
	test_expansion(128'hda8568f5b7d870e81e6c5233cbaf2581, {16'd44812, 16'd51927, 16'd40066, 16'd21848, 16'd15771, 16'd4623, 16'd47789, 16'd42170, 16'd7650, 16'd54090, 16'd30207, 16'd41894, 16'd23351, 16'd52401, 16'd28030, 16'd31501, 16'd56232, 16'd30575, 16'd40857, 16'd29152, 16'd19684, 16'd60868, 16'd4915, 16'd11533, 16'd55327, 16'd62678});
	test_expansion(128'h2ad806f174be3f317286ff06034c5973, {16'd46010, 16'd3439, 16'd38193, 16'd9411, 16'd13175, 16'd13953, 16'd47594, 16'd8704, 16'd39972, 16'd21550, 16'd12398, 16'd11074, 16'd3904, 16'd30267, 16'd32194, 16'd24681, 16'd12403, 16'd20853, 16'd65478, 16'd23973, 16'd12813, 16'd61148, 16'd14770, 16'd10393, 16'd24918, 16'd58389});
	test_expansion(128'h339ab2690b7017cb89e4fbb39fdc1f77, {16'd27667, 16'd37062, 16'd60547, 16'd24711, 16'd50653, 16'd778, 16'd44096, 16'd39264, 16'd50712, 16'd20270, 16'd20394, 16'd26999, 16'd65512, 16'd7399, 16'd52614, 16'd25509, 16'd26728, 16'd38367, 16'd50116, 16'd39344, 16'd37559, 16'd56015, 16'd49808, 16'd34843, 16'd24677, 16'd4863});
	test_expansion(128'h53d5d56e3b15f3eec3139cb8847380e9, {16'd33300, 16'd31350, 16'd6548, 16'd22983, 16'd1836, 16'd59815, 16'd27894, 16'd18704, 16'd16447, 16'd34688, 16'd6114, 16'd21527, 16'd25869, 16'd8463, 16'd627, 16'd31390, 16'd8299, 16'd54712, 16'd58509, 16'd34382, 16'd27456, 16'd25726, 16'd41671, 16'd55250, 16'd44289, 16'd37965});
	test_expansion(128'hd9fd66b5cd34c18f79508120b6474a13, {16'd46644, 16'd36857, 16'd24365, 16'd49469, 16'd24857, 16'd31744, 16'd60144, 16'd35166, 16'd2879, 16'd22993, 16'd44839, 16'd33545, 16'd25366, 16'd43176, 16'd23807, 16'd20489, 16'd56871, 16'd61624, 16'd54689, 16'd49901, 16'd6188, 16'd53209, 16'd19881, 16'd60281, 16'd43142, 16'd45621});
	test_expansion(128'h8db0d88c9b89acbe7ba979c5b103a068, {16'd62156, 16'd17037, 16'd52555, 16'd19486, 16'd51316, 16'd56268, 16'd57269, 16'd16194, 16'd43808, 16'd55157, 16'd2991, 16'd19482, 16'd60793, 16'd44851, 16'd3396, 16'd6032, 16'd59232, 16'd29300, 16'd2602, 16'd55880, 16'd19263, 16'd47713, 16'd39728, 16'd9726, 16'd57561, 16'd28081});
	test_expansion(128'h4c17429003f5955bab3d839826cd22fc, {16'd16510, 16'd57989, 16'd35675, 16'd57651, 16'd15407, 16'd39783, 16'd3101, 16'd20715, 16'd48989, 16'd13520, 16'd35357, 16'd65315, 16'd51152, 16'd32863, 16'd16426, 16'd1567, 16'd5887, 16'd48917, 16'd22970, 16'd35135, 16'd23155, 16'd7555, 16'd39560, 16'd40793, 16'd39866, 16'd2801});
	test_expansion(128'h4a4a835c8a320df71e52209baf6ee45f, {16'd41066, 16'd39452, 16'd56956, 16'd40699, 16'd63557, 16'd254, 16'd23302, 16'd7475, 16'd63688, 16'd52377, 16'd21861, 16'd14667, 16'd5367, 16'd19280, 16'd49391, 16'd65016, 16'd26168, 16'd12271, 16'd6781, 16'd14136, 16'd29856, 16'd18478, 16'd39781, 16'd46247, 16'd61533, 16'd7086});
	test_expansion(128'h9626e6bc9d3e2656f63b782b8206b8f2, {16'd21842, 16'd64988, 16'd45594, 16'd47718, 16'd34120, 16'd2250, 16'd60358, 16'd60847, 16'd31735, 16'd45880, 16'd5239, 16'd37380, 16'd62914, 16'd21336, 16'd45024, 16'd1996, 16'd16442, 16'd12827, 16'd30821, 16'd5284, 16'd57723, 16'd32661, 16'd39250, 16'd24798, 16'd15983, 16'd27429});
	test_expansion(128'h37f90e5b9ada84c8b55d596925c14627, {16'd37331, 16'd18312, 16'd24110, 16'd29614, 16'd34265, 16'd53634, 16'd57213, 16'd35475, 16'd45934, 16'd22636, 16'd17221, 16'd31122, 16'd61838, 16'd33777, 16'd24092, 16'd45764, 16'd35129, 16'd63758, 16'd36940, 16'd28322, 16'd41009, 16'd27121, 16'd8202, 16'd2810, 16'd13896, 16'd31614});
	test_expansion(128'hd73a5a4acc575107858f23b54a58d29e, {16'd54331, 16'd44096, 16'd3328, 16'd39728, 16'd8496, 16'd45595, 16'd51146, 16'd44868, 16'd49569, 16'd41849, 16'd20747, 16'd6787, 16'd55867, 16'd27652, 16'd53647, 16'd58981, 16'd34774, 16'd28358, 16'd62075, 16'd53414, 16'd1656, 16'd45935, 16'd33435, 16'd15037, 16'd62902, 16'd12524});
	test_expansion(128'he7064e509bb8e9faa66239821084b2a8, {16'd7258, 16'd18229, 16'd30225, 16'd39314, 16'd35987, 16'd48174, 16'd43556, 16'd54293, 16'd7879, 16'd59263, 16'd43182, 16'd39998, 16'd3546, 16'd53120, 16'd6082, 16'd62230, 16'd53097, 16'd42064, 16'd38610, 16'd61134, 16'd36275, 16'd45194, 16'd57224, 16'd4872, 16'd31754, 16'd54224});
	test_expansion(128'hcc8005243e98b8c6db5ad9324c838ce7, {16'd35782, 16'd4156, 16'd47183, 16'd24594, 16'd21170, 16'd4161, 16'd53511, 16'd42974, 16'd39106, 16'd10224, 16'd51220, 16'd9183, 16'd34894, 16'd55925, 16'd25956, 16'd20319, 16'd7607, 16'd46205, 16'd31587, 16'd42192, 16'd51426, 16'd30821, 16'd41352, 16'd20461, 16'd32871, 16'd4135});
	test_expansion(128'h14427d13637feaa70cd549e6d81862f1, {16'd43780, 16'd62714, 16'd42870, 16'd50607, 16'd21327, 16'd43101, 16'd48721, 16'd35144, 16'd35090, 16'd47909, 16'd63254, 16'd48621, 16'd17041, 16'd17036, 16'd34187, 16'd10977, 16'd45675, 16'd48088, 16'd59911, 16'd1351, 16'd4357, 16'd45951, 16'd18432, 16'd32558, 16'd18464, 16'd39509});
	test_expansion(128'ha4112535209f4ee6f32a18bdb46ce6b2, {16'd1009, 16'd62845, 16'd19653, 16'd35550, 16'd33246, 16'd43847, 16'd44269, 16'd38138, 16'd1581, 16'd29244, 16'd13159, 16'd33030, 16'd3429, 16'd1649, 16'd18230, 16'd18579, 16'd20947, 16'd10305, 16'd51440, 16'd9922, 16'd19033, 16'd44608, 16'd63076, 16'd12073, 16'd43351, 16'd61621});
	test_expansion(128'h0e92c243329b8168b2c73753a341ccce, {16'd6309, 16'd39173, 16'd40089, 16'd40163, 16'd21928, 16'd47601, 16'd63157, 16'd14722, 16'd53969, 16'd58784, 16'd32115, 16'd15411, 16'd27834, 16'd30809, 16'd45067, 16'd18993, 16'd48496, 16'd3384, 16'd12546, 16'd41591, 16'd54399, 16'd64854, 16'd40651, 16'd8467, 16'd50772, 16'd56542});
	test_expansion(128'h485d09b19b36044ec9c100394deb7c8d, {16'd64230, 16'd27445, 16'd49247, 16'd51780, 16'd2310, 16'd52903, 16'd36199, 16'd51599, 16'd45167, 16'd6532, 16'd46230, 16'd32043, 16'd29932, 16'd42481, 16'd1969, 16'd64334, 16'd36110, 16'd59740, 16'd6829, 16'd36858, 16'd55771, 16'd29638, 16'd1643, 16'd11814, 16'd56705, 16'd8190});
	test_expansion(128'h0aa1cf3a57fd7dec39a2b6b6e86fde23, {16'd40500, 16'd7561, 16'd30600, 16'd51191, 16'd33260, 16'd10487, 16'd23570, 16'd60160, 16'd31095, 16'd59610, 16'd40369, 16'd3142, 16'd35584, 16'd29625, 16'd15734, 16'd28196, 16'd8789, 16'd28793, 16'd27512, 16'd60594, 16'd34929, 16'd52571, 16'd9844, 16'd57327, 16'd17806, 16'd61339});
	test_expansion(128'h41ac3de6aff0e3116aebde408df73e4f, {16'd56101, 16'd48687, 16'd55083, 16'd25607, 16'd65254, 16'd150, 16'd6783, 16'd46878, 16'd18304, 16'd38436, 16'd39251, 16'd25268, 16'd23461, 16'd56086, 16'd55000, 16'd19344, 16'd27492, 16'd55062, 16'd36261, 16'd25600, 16'd44515, 16'd11931, 16'd24325, 16'd4530, 16'd31344, 16'd40261});
	test_expansion(128'hfce0a0f6df859a2fe9fe4f7a498d3401, {16'd62685, 16'd24180, 16'd15263, 16'd478, 16'd61064, 16'd49767, 16'd18228, 16'd15272, 16'd45573, 16'd59547, 16'd27452, 16'd10717, 16'd38001, 16'd30037, 16'd25876, 16'd8609, 16'd16387, 16'd22781, 16'd56214, 16'd39359, 16'd57411, 16'd48410, 16'd41050, 16'd63609, 16'd28563, 16'd5734});
	test_expansion(128'h9434d07bc4091218a4276486ec0ba7a5, {16'd23225, 16'd26705, 16'd59689, 16'd28441, 16'd31024, 16'd14116, 16'd4734, 16'd57988, 16'd36541, 16'd22895, 16'd57723, 16'd19868, 16'd35164, 16'd18354, 16'd11519, 16'd59538, 16'd62820, 16'd46790, 16'd47124, 16'd27966, 16'd52317, 16'd25216, 16'd11366, 16'd31558, 16'd50602, 16'd2764});
	test_expansion(128'hd16dcc5460f19fc4edd46d6a05f9c2ed, {16'd12820, 16'd13386, 16'd18829, 16'd28807, 16'd60012, 16'd14098, 16'd58064, 16'd55425, 16'd59304, 16'd58956, 16'd40860, 16'd22929, 16'd2804, 16'd21725, 16'd341, 16'd39541, 16'd44971, 16'd4086, 16'd51613, 16'd37284, 16'd11494, 16'd55558, 16'd50091, 16'd17642, 16'd28741, 16'd11636});
	test_expansion(128'h51b279ba97ea5b7139b932486b58fdc3, {16'd31506, 16'd39925, 16'd55046, 16'd30094, 16'd32722, 16'd56677, 16'd6198, 16'd16543, 16'd50739, 16'd29090, 16'd42636, 16'd35914, 16'd19512, 16'd30117, 16'd6988, 16'd22179, 16'd20070, 16'd46187, 16'd10433, 16'd50245, 16'd3828, 16'd62534, 16'd51803, 16'd41183, 16'd18726, 16'd58725});
	test_expansion(128'hcb47823a62b5f5b7545c483cc6f2ea2f, {16'd3288, 16'd2438, 16'd14402, 16'd64331, 16'd63973, 16'd59750, 16'd54212, 16'd18816, 16'd21848, 16'd63265, 16'd61414, 16'd61195, 16'd25097, 16'd22159, 16'd44258, 16'd53025, 16'd26404, 16'd35586, 16'd35687, 16'd17426, 16'd62129, 16'd17949, 16'd27246, 16'd45442, 16'd34246, 16'd4833});
	test_expansion(128'h63b4fca993cfeecabcd5f26cc8507b61, {16'd36209, 16'd6292, 16'd51993, 16'd50957, 16'd7960, 16'd5068, 16'd16283, 16'd65476, 16'd5539, 16'd38519, 16'd8578, 16'd26479, 16'd32196, 16'd31138, 16'd48872, 16'd29896, 16'd22459, 16'd46874, 16'd44788, 16'd62079, 16'd43086, 16'd53097, 16'd37676, 16'd13257, 16'd57420, 16'd30174});
	test_expansion(128'h0c0d2951a76ddce9326b9ad970e09bde, {16'd58032, 16'd11729, 16'd17526, 16'd55619, 16'd58775, 16'd10173, 16'd36460, 16'd15403, 16'd18357, 16'd8658, 16'd50018, 16'd22394, 16'd23987, 16'd1220, 16'd1576, 16'd16009, 16'd64190, 16'd63424, 16'd35732, 16'd30766, 16'd34611, 16'd27962, 16'd32112, 16'd6214, 16'd8718, 16'd56610});
	test_expansion(128'h2eaa3964e98c1ba3962f63767bc79b59, {16'd51608, 16'd28353, 16'd4483, 16'd50048, 16'd18496, 16'd65402, 16'd36680, 16'd28225, 16'd40816, 16'd23885, 16'd16897, 16'd30686, 16'd35258, 16'd61624, 16'd63365, 16'd45479, 16'd5710, 16'd1079, 16'd29896, 16'd49598, 16'd39528, 16'd17625, 16'd46119, 16'd14455, 16'd2774, 16'd51943});
	test_expansion(128'ha7e1ee20c84607c91cd712f294682970, {16'd20433, 16'd62541, 16'd43347, 16'd50512, 16'd43518, 16'd43604, 16'd26605, 16'd5037, 16'd42426, 16'd57162, 16'd51476, 16'd19638, 16'd7610, 16'd63443, 16'd43391, 16'd36168, 16'd20817, 16'd47643, 16'd55138, 16'd58049, 16'd55166, 16'd54631, 16'd38821, 16'd58973, 16'd56614, 16'd22250});
	test_expansion(128'hb4fe67fcafd92fe908c8528721ef05e0, {16'd33170, 16'd796, 16'd32530, 16'd18702, 16'd22091, 16'd52135, 16'd13757, 16'd14724, 16'd49746, 16'd17400, 16'd1618, 16'd45294, 16'd45006, 16'd63971, 16'd51277, 16'd25873, 16'd42553, 16'd27303, 16'd38141, 16'd26631, 16'd59230, 16'd53502, 16'd38290, 16'd6083, 16'd20372, 16'd13163});
	test_expansion(128'hc23b85d30b7c64f0d7ad83aa8662dd81, {16'd9576, 16'd52507, 16'd42813, 16'd37608, 16'd5261, 16'd33800, 16'd21992, 16'd35972, 16'd5556, 16'd37173, 16'd22120, 16'd50765, 16'd32470, 16'd21758, 16'd38066, 16'd1891, 16'd35768, 16'd39358, 16'd12044, 16'd37179, 16'd59422, 16'd15204, 16'd10549, 16'd22758, 16'd18173, 16'd38209});
	test_expansion(128'hb2ab0e8cf2782ff2053e2bb892f72c62, {16'd28603, 16'd24913, 16'd63059, 16'd54318, 16'd34105, 16'd15950, 16'd57686, 16'd26112, 16'd41737, 16'd46102, 16'd12134, 16'd47957, 16'd44512, 16'd52579, 16'd18222, 16'd56208, 16'd52676, 16'd60307, 16'd16313, 16'd55173, 16'd53444, 16'd20102, 16'd31290, 16'd22879, 16'd51695, 16'd8273});
	test_expansion(128'ha22878a6287d25bebf4392f0184bb9c5, {16'd43398, 16'd62867, 16'd9713, 16'd61778, 16'd65470, 16'd49807, 16'd55003, 16'd47179, 16'd13250, 16'd3557, 16'd15958, 16'd46576, 16'd1018, 16'd52415, 16'd49529, 16'd65069, 16'd64055, 16'd25276, 16'd3365, 16'd19532, 16'd60115, 16'd14654, 16'd12449, 16'd34635, 16'd49706, 16'd5952});
	test_expansion(128'h0d8e79401da3d74a51508c0bd00f43cb, {16'd23040, 16'd49525, 16'd45072, 16'd62095, 16'd39024, 16'd10007, 16'd27792, 16'd1205, 16'd4144, 16'd12310, 16'd39435, 16'd45843, 16'd38568, 16'd16633, 16'd58231, 16'd61489, 16'd11305, 16'd4357, 16'd37461, 16'd24711, 16'd12493, 16'd50142, 16'd14588, 16'd27641, 16'd18050, 16'd41067});
	test_expansion(128'h87460bc9c2f5b2962edc571130a062a6, {16'd48251, 16'd50699, 16'd37153, 16'd52520, 16'd24163, 16'd42344, 16'd16030, 16'd15133, 16'd52131, 16'd62862, 16'd53108, 16'd36491, 16'd5475, 16'd19953, 16'd37495, 16'd38628, 16'd63613, 16'd8190, 16'd16855, 16'd43845, 16'd63939, 16'd39787, 16'd56126, 16'd3045, 16'd32410, 16'd54779});
	test_expansion(128'hdcea2f16706cfac054ac65cc2fc4a7b4, {16'd17137, 16'd12131, 16'd8237, 16'd54339, 16'd28035, 16'd23268, 16'd2232, 16'd10773, 16'd16906, 16'd42796, 16'd32164, 16'd539, 16'd10336, 16'd12745, 16'd24535, 16'd40852, 16'd63563, 16'd42543, 16'd58511, 16'd12226, 16'd55475, 16'd34992, 16'd15974, 16'd996, 16'd18592, 16'd22805});
	test_expansion(128'haf985a256da94229936f9e3e8d5db094, {16'd10001, 16'd26044, 16'd13695, 16'd45128, 16'd17876, 16'd49687, 16'd6249, 16'd34512, 16'd37667, 16'd2350, 16'd20949, 16'd37024, 16'd6656, 16'd27222, 16'd6111, 16'd63837, 16'd1501, 16'd14907, 16'd6788, 16'd2516, 16'd10975, 16'd11150, 16'd14721, 16'd64568, 16'd15627, 16'd31505});
	test_expansion(128'h51f236bb716e1b9680e6bc467184987b, {16'd328, 16'd6420, 16'd48698, 16'd4671, 16'd60863, 16'd29846, 16'd27425, 16'd7166, 16'd25312, 16'd36966, 16'd3346, 16'd17825, 16'd36652, 16'd18811, 16'd8822, 16'd53044, 16'd62273, 16'd43958, 16'd56371, 16'd53492, 16'd59603, 16'd26033, 16'd46707, 16'd27292, 16'd9216, 16'd36411});
	test_expansion(128'h28cf215a95dd5fb74f5ddbfcc8c78b96, {16'd47260, 16'd42420, 16'd28852, 16'd23042, 16'd54281, 16'd60637, 16'd3966, 16'd52390, 16'd46953, 16'd8593, 16'd9022, 16'd55279, 16'd12023, 16'd62536, 16'd2210, 16'd46962, 16'd12978, 16'd24196, 16'd56418, 16'd62435, 16'd57119, 16'd1899, 16'd33128, 16'd24363, 16'd19421, 16'd61954});
	test_expansion(128'h6af84df9a0e5f61e37b694fef93bceef, {16'd12773, 16'd8306, 16'd28404, 16'd48476, 16'd14167, 16'd39312, 16'd29121, 16'd44972, 16'd15877, 16'd62675, 16'd5466, 16'd24189, 16'd20021, 16'd53255, 16'd62220, 16'd61491, 16'd54003, 16'd3052, 16'd63080, 16'd9629, 16'd43453, 16'd19229, 16'd35768, 16'd54809, 16'd48403, 16'd54169});
	test_expansion(128'h8b514a6f3b6c3188fd73b903e5bd1437, {16'd14082, 16'd27239, 16'd63881, 16'd20016, 16'd38990, 16'd9946, 16'd39792, 16'd22478, 16'd396, 16'd43706, 16'd15710, 16'd7519, 16'd42745, 16'd42204, 16'd38575, 16'd47725, 16'd18586, 16'd2146, 16'd18648, 16'd9593, 16'd10318, 16'd33950, 16'd28986, 16'd64441, 16'd378, 16'd20364});
	test_expansion(128'hba98d012d4175093c2da76e87315a7e9, {16'd36709, 16'd3924, 16'd16406, 16'd48619, 16'd51370, 16'd35591, 16'd29486, 16'd8444, 16'd7755, 16'd50613, 16'd36800, 16'd56065, 16'd62943, 16'd34883, 16'd1078, 16'd1201, 16'd43642, 16'd43550, 16'd48647, 16'd32713, 16'd39305, 16'd50942, 16'd36407, 16'd10483, 16'd35510, 16'd26866});
	test_expansion(128'h7a4c1516465165a2a9c1c5f9c192795a, {16'd50055, 16'd37915, 16'd42715, 16'd15958, 16'd44929, 16'd33985, 16'd57888, 16'd42404, 16'd27950, 16'd24589, 16'd15897, 16'd61304, 16'd14442, 16'd61862, 16'd53266, 16'd40547, 16'd23041, 16'd44677, 16'd57738, 16'd37950, 16'd58225, 16'd17490, 16'd28831, 16'd34682, 16'd17740, 16'd39066});
	test_expansion(128'h36fc13b39f7981ba354b7f7f0c73f232, {16'd31503, 16'd13506, 16'd5085, 16'd29001, 16'd24188, 16'd10130, 16'd31586, 16'd9083, 16'd3655, 16'd35697, 16'd19604, 16'd36695, 16'd62617, 16'd35631, 16'd46897, 16'd46798, 16'd11469, 16'd7222, 16'd9639, 16'd30437, 16'd16481, 16'd1164, 16'd34726, 16'd10131, 16'd37769, 16'd9665});
	test_expansion(128'h1d9825e4da091b357cbbefdab86958ea, {16'd21272, 16'd22665, 16'd9667, 16'd20455, 16'd18556, 16'd319, 16'd38051, 16'd12501, 16'd26203, 16'd45405, 16'd1455, 16'd15465, 16'd65102, 16'd62795, 16'd46425, 16'd36559, 16'd24888, 16'd135, 16'd53013, 16'd19325, 16'd15515, 16'd27997, 16'd57653, 16'd33555, 16'd38362, 16'd56487});
	test_expansion(128'h5dc9af82ef77562f4eb0dc9bff84edc0, {16'd64331, 16'd8258, 16'd34140, 16'd47583, 16'd6690, 16'd19237, 16'd25476, 16'd19433, 16'd43393, 16'd49814, 16'd24723, 16'd44899, 16'd20338, 16'd2399, 16'd16662, 16'd59623, 16'd45072, 16'd49349, 16'd44755, 16'd17723, 16'd21851, 16'd36124, 16'd40512, 16'd26753, 16'd28047, 16'd34378});
	test_expansion(128'h5b7c87b5daa16e6750b38c6aa5dde764, {16'd1929, 16'd40330, 16'd15654, 16'd15491, 16'd47339, 16'd60769, 16'd47172, 16'd3082, 16'd32896, 16'd18930, 16'd29357, 16'd37606, 16'd10277, 16'd36383, 16'd23126, 16'd22677, 16'd8663, 16'd27922, 16'd8722, 16'd32254, 16'd45482, 16'd5560, 16'd35554, 16'd57421, 16'd32355, 16'd13236});
	test_expansion(128'h85b3d057cbb0fab30d0d8b13a3b4cd4c, {16'd58650, 16'd49788, 16'd14607, 16'd54710, 16'd47197, 16'd23514, 16'd41674, 16'd20935, 16'd12775, 16'd4639, 16'd35254, 16'd49086, 16'd183, 16'd36849, 16'd56056, 16'd12518, 16'd20380, 16'd17920, 16'd10541, 16'd585, 16'd21290, 16'd24850, 16'd51632, 16'd47056, 16'd37811, 16'd18871});
	test_expansion(128'h0b47901e4907b03c38e8dafce80f273e, {16'd47002, 16'd51517, 16'd22971, 16'd39507, 16'd9797, 16'd60535, 16'd27237, 16'd58299, 16'd552, 16'd16854, 16'd54937, 16'd49950, 16'd39808, 16'd58976, 16'd53335, 16'd22941, 16'd47809, 16'd56585, 16'd13161, 16'd60318, 16'd25188, 16'd50451, 16'd42825, 16'd63984, 16'd13824, 16'd41420});
	test_expansion(128'h5de5f891da16d9f081510fd020f18809, {16'd10433, 16'd50268, 16'd39553, 16'd43025, 16'd20363, 16'd41951, 16'd10131, 16'd31841, 16'd17388, 16'd49127, 16'd2726, 16'd50271, 16'd15615, 16'd29137, 16'd22154, 16'd39106, 16'd44150, 16'd43688, 16'd13404, 16'd10278, 16'd44766, 16'd15280, 16'd8353, 16'd15168, 16'd42902, 16'd19002});
	test_expansion(128'h2c6325c72e9a1e1138aba65934457f60, {16'd36839, 16'd21465, 16'd48632, 16'd32589, 16'd47710, 16'd64986, 16'd61314, 16'd37446, 16'd36515, 16'd29, 16'd34374, 16'd43657, 16'd27018, 16'd3707, 16'd49116, 16'd20481, 16'd13921, 16'd30105, 16'd44409, 16'd16355, 16'd15513, 16'd25444, 16'd55088, 16'd50779, 16'd4339, 16'd56988});
	test_expansion(128'h5c929ac95ad3c6d2b13f583168ed739f, {16'd42715, 16'd15429, 16'd16580, 16'd34283, 16'd37858, 16'd20253, 16'd65341, 16'd8642, 16'd45037, 16'd56894, 16'd23682, 16'd58947, 16'd16907, 16'd36034, 16'd13001, 16'd35348, 16'd39277, 16'd26642, 16'd13894, 16'd44026, 16'd38398, 16'd35908, 16'd41856, 16'd26491, 16'd26833, 16'd870});
	test_expansion(128'h1c42f7b9a933bcf2e52e0a81a86986ad, {16'd34667, 16'd5950, 16'd44909, 16'd57141, 16'd57694, 16'd15567, 16'd540, 16'd32813, 16'd35635, 16'd61908, 16'd44602, 16'd33376, 16'd12083, 16'd24923, 16'd11796, 16'd57522, 16'd24943, 16'd46744, 16'd29977, 16'd24186, 16'd12061, 16'd57944, 16'd64687, 16'd11482, 16'd30045, 16'd7522});
	test_expansion(128'hf183d29fe49cb34b7b5fdd3d2ab1f708, {16'd15396, 16'd11841, 16'd37401, 16'd27699, 16'd39604, 16'd60347, 16'd56961, 16'd11545, 16'd61514, 16'd52197, 16'd27252, 16'd33262, 16'd45303, 16'd15567, 16'd19993, 16'd31303, 16'd1317, 16'd11957, 16'd6603, 16'd20145, 16'd12009, 16'd61264, 16'd27364, 16'd15122, 16'd28535, 16'd9359});
	test_expansion(128'h04b1e3ec2c0ff40e1897e4d199cbfa50, {16'd52263, 16'd14577, 16'd58910, 16'd26889, 16'd52990, 16'd52041, 16'd46798, 16'd5486, 16'd65050, 16'd53275, 16'd17354, 16'd17385, 16'd63613, 16'd45197, 16'd2251, 16'd51639, 16'd27901, 16'd36325, 16'd33720, 16'd19210, 16'd61540, 16'd46658, 16'd35506, 16'd38958, 16'd7894, 16'd26319});
	test_expansion(128'h4f7f9ac0d65ba1be84c0808788dcc59e, {16'd24013, 16'd64602, 16'd32984, 16'd23553, 16'd36074, 16'd41270, 16'd63273, 16'd38501, 16'd8037, 16'd30751, 16'd2511, 16'd4097, 16'd6809, 16'd9983, 16'd34173, 16'd3586, 16'd53777, 16'd14084, 16'd12509, 16'd39332, 16'd58252, 16'd44455, 16'd45384, 16'd7390, 16'd59595, 16'd32373});
	test_expansion(128'h02648498a5f44810cb6ccd0ddf94d37c, {16'd3188, 16'd10907, 16'd12532, 16'd41261, 16'd28547, 16'd6320, 16'd5468, 16'd29727, 16'd18617, 16'd1933, 16'd53101, 16'd43363, 16'd41667, 16'd46088, 16'd8870, 16'd55692, 16'd15916, 16'd63228, 16'd55904, 16'd51849, 16'd65215, 16'd48287, 16'd18272, 16'd2428, 16'd25069, 16'd14364});
	test_expansion(128'h09f6156493813d1d0bfe82c104156e3d, {16'd51914, 16'd56105, 16'd45072, 16'd35967, 16'd44971, 16'd53963, 16'd35242, 16'd54340, 16'd40376, 16'd60398, 16'd63685, 16'd46234, 16'd11496, 16'd1668, 16'd59233, 16'd55462, 16'd1830, 16'd23889, 16'd63526, 16'd55099, 16'd41824, 16'd10514, 16'd50842, 16'd2925, 16'd20591, 16'd45598});
	test_expansion(128'hac1d98110b140dedcf5743a0b8658107, {16'd29587, 16'd19315, 16'd4935, 16'd34549, 16'd9194, 16'd31736, 16'd41960, 16'd19705, 16'd51170, 16'd43379, 16'd28884, 16'd28818, 16'd32000, 16'd27573, 16'd33229, 16'd8188, 16'd63610, 16'd33266, 16'd9387, 16'd13924, 16'd52749, 16'd57073, 16'd27473, 16'd38773, 16'd48654, 16'd13235});
	test_expansion(128'h516d57f7cb5e4753eb65c5869baea10a, {16'd41432, 16'd26039, 16'd15206, 16'd23200, 16'd58096, 16'd17773, 16'd58654, 16'd24056, 16'd8514, 16'd25765, 16'd58502, 16'd45321, 16'd26866, 16'd55197, 16'd59917, 16'd52683, 16'd46114, 16'd58460, 16'd3499, 16'd28331, 16'd47888, 16'd25511, 16'd16955, 16'd4176, 16'd17556, 16'd60708});
	test_expansion(128'h237a10726c81c10f9f197bd697b79560, {16'd22381, 16'd7764, 16'd25350, 16'd14174, 16'd52721, 16'd42489, 16'd52418, 16'd47511, 16'd60552, 16'd37367, 16'd25133, 16'd39302, 16'd26355, 16'd36978, 16'd30646, 16'd39269, 16'd25898, 16'd13600, 16'd23558, 16'd41187, 16'd21336, 16'd4308, 16'd12620, 16'd9048, 16'd12130, 16'd39597});
	test_expansion(128'hef96aa12ed3addc882e313db226a0f71, {16'd56427, 16'd23555, 16'd6982, 16'd64073, 16'd59206, 16'd59645, 16'd11233, 16'd55894, 16'd8044, 16'd58799, 16'd35992, 16'd37345, 16'd17978, 16'd35363, 16'd57146, 16'd39649, 16'd39333, 16'd13937, 16'd20207, 16'd47261, 16'd33207, 16'd40267, 16'd26065, 16'd62214, 16'd53135, 16'd48261});
	test_expansion(128'he83f2496c224df20c589db9ed62d41f4, {16'd26343, 16'd29514, 16'd61377, 16'd58433, 16'd39909, 16'd62242, 16'd31866, 16'd3267, 16'd41663, 16'd60956, 16'd36709, 16'd10836, 16'd63148, 16'd51148, 16'd39178, 16'd24058, 16'd418, 16'd34966, 16'd20367, 16'd5109, 16'd57304, 16'd31834, 16'd16425, 16'd5509, 16'd52111, 16'd29474});
	test_expansion(128'h582d26ca5a68229a488e3dd08c09ac6f, {16'd5672, 16'd39585, 16'd9151, 16'd3715, 16'd14476, 16'd39845, 16'd42544, 16'd10658, 16'd51046, 16'd26411, 16'd30421, 16'd31453, 16'd19533, 16'd37920, 16'd49322, 16'd45594, 16'd41237, 16'd15166, 16'd9114, 16'd34988, 16'd11404, 16'd20105, 16'd35666, 16'd60433, 16'd14685, 16'd14181});
	test_expansion(128'h3323b2f59b869e081479018a3eae8572, {16'd56465, 16'd8881, 16'd23451, 16'd19615, 16'd64267, 16'd4139, 16'd13097, 16'd32681, 16'd40537, 16'd22060, 16'd24104, 16'd12492, 16'd14028, 16'd51082, 16'd8641, 16'd2928, 16'd6582, 16'd42604, 16'd51193, 16'd2740, 16'd34612, 16'd5475, 16'd49706, 16'd45186, 16'd21648, 16'd40144});
	test_expansion(128'h2dc3bebfae3291f13a8c788365c8d831, {16'd27424, 16'd18920, 16'd56731, 16'd4383, 16'd28621, 16'd30909, 16'd9295, 16'd31707, 16'd48920, 16'd15779, 16'd9296, 16'd54837, 16'd12463, 16'd29146, 16'd48150, 16'd18813, 16'd39057, 16'd49846, 16'd33848, 16'd19192, 16'd51397, 16'd61492, 16'd53778, 16'd28383, 16'd47511, 16'd17566});
	test_expansion(128'haf37772a23151e14af3be8b71fee56d0, {16'd42984, 16'd58273, 16'd61421, 16'd21681, 16'd4812, 16'd58100, 16'd61645, 16'd30468, 16'd44586, 16'd30430, 16'd34792, 16'd11134, 16'd16371, 16'd36120, 16'd43537, 16'd33380, 16'd37737, 16'd24120, 16'd60071, 16'd63393, 16'd41133, 16'd4445, 16'd43343, 16'd17870, 16'd20183, 16'd15702});
	test_expansion(128'hfef526ab181bf30e5d562e382a3a3805, {16'd44719, 16'd57701, 16'd52345, 16'd3098, 16'd59923, 16'd26803, 16'd34626, 16'd9184, 16'd52136, 16'd22135, 16'd14654, 16'd65120, 16'd10789, 16'd22497, 16'd6048, 16'd44860, 16'd61098, 16'd23911, 16'd41481, 16'd36240, 16'd20871, 16'd1769, 16'd26122, 16'd5889, 16'd60991, 16'd6201});
	test_expansion(128'h7563e554aab708d935925565669709f8, {16'd41890, 16'd65467, 16'd64088, 16'd5203, 16'd23978, 16'd26375, 16'd17290, 16'd25783, 16'd31837, 16'd38383, 16'd24111, 16'd10417, 16'd4935, 16'd50960, 16'd5812, 16'd4256, 16'd61889, 16'd13987, 16'd12070, 16'd46292, 16'd41916, 16'd5677, 16'd30426, 16'd49276, 16'd35795, 16'd6226});
	test_expansion(128'hb207b65ce9d018577da7b1415f4c0572, {16'd1183, 16'd20983, 16'd64719, 16'd38557, 16'd4477, 16'd57191, 16'd31034, 16'd41199, 16'd16005, 16'd50903, 16'd30185, 16'd10139, 16'd31738, 16'd56043, 16'd31314, 16'd27598, 16'd40372, 16'd12707, 16'd4094, 16'd1961, 16'd42410, 16'd25753, 16'd4968, 16'd23251, 16'd41719, 16'd35724});
	test_expansion(128'hf95d58aa48bebab03a91dfeb1bfd14dc, {16'd925, 16'd3582, 16'd31985, 16'd34128, 16'd12915, 16'd56939, 16'd40279, 16'd34420, 16'd10509, 16'd1665, 16'd44646, 16'd16011, 16'd13252, 16'd27845, 16'd20288, 16'd3791, 16'd1901, 16'd23815, 16'd28619, 16'd16945, 16'd59688, 16'd2986, 16'd56153, 16'd60223, 16'd21487, 16'd15982});
	test_expansion(128'h69bb385ccb2d55ebefc99e0a5bca8510, {16'd13139, 16'd65007, 16'd45374, 16'd5291, 16'd29441, 16'd45174, 16'd11003, 16'd51360, 16'd27657, 16'd14454, 16'd24292, 16'd3248, 16'd2434, 16'd14102, 16'd53268, 16'd516, 16'd34374, 16'd10432, 16'd11127, 16'd20633, 16'd36591, 16'd11832, 16'd60532, 16'd33066, 16'd27716, 16'd4880});
	test_expansion(128'h1569d543cbb779fb117534886ea45fe6, {16'd17316, 16'd64789, 16'd31780, 16'd56250, 16'd56575, 16'd33859, 16'd21835, 16'd44599, 16'd25280, 16'd869, 16'd9815, 16'd38578, 16'd39160, 16'd43089, 16'd13395, 16'd18539, 16'd54005, 16'd143, 16'd52725, 16'd47893, 16'd63807, 16'd56256, 16'd28303, 16'd34084, 16'd37772, 16'd1063});
	test_expansion(128'h50d181c0e011f5d1aad240005aea300d, {16'd9064, 16'd2716, 16'd55658, 16'd63843, 16'd56341, 16'd55855, 16'd3192, 16'd29529, 16'd38366, 16'd35099, 16'd487, 16'd63697, 16'd42169, 16'd6816, 16'd24287, 16'd47750, 16'd25885, 16'd56672, 16'd52884, 16'd24571, 16'd9574, 16'd17440, 16'd16604, 16'd1740, 16'd64525, 16'd1650});
	test_expansion(128'ha6d03a888a2728193c743e275e7b233b, {16'd29074, 16'd52559, 16'd3039, 16'd51439, 16'd34613, 16'd39260, 16'd58493, 16'd49050, 16'd23402, 16'd48984, 16'd19059, 16'd35939, 16'd23933, 16'd42575, 16'd11409, 16'd554, 16'd47143, 16'd6639, 16'd35528, 16'd44395, 16'd10168, 16'd8528, 16'd28575, 16'd10750, 16'd34439, 16'd45132});
	test_expansion(128'hb19329c1946108fbff0d60ba93629155, {16'd42676, 16'd32625, 16'd26321, 16'd39129, 16'd4397, 16'd59337, 16'd24068, 16'd34354, 16'd11504, 16'd17741, 16'd41240, 16'd12450, 16'd45984, 16'd21730, 16'd28173, 16'd57905, 16'd57952, 16'd50691, 16'd4250, 16'd64006, 16'd58834, 16'd14805, 16'd8686, 16'd54875, 16'd48721, 16'd51857});
	test_expansion(128'h521f5c6151a942dba7df688872b80ab9, {16'd12895, 16'd35372, 16'd51776, 16'd23401, 16'd13438, 16'd34938, 16'd13619, 16'd63059, 16'd36765, 16'd57647, 16'd5330, 16'd25300, 16'd43591, 16'd32900, 16'd41052, 16'd62092, 16'd60931, 16'd61572, 16'd5352, 16'd27256, 16'd46001, 16'd49272, 16'd43720, 16'd4137, 16'd28024, 16'd29111});
	test_expansion(128'h1585a8f8ae1bbbbd9dd29ce7126bd95f, {16'd60824, 16'd13219, 16'd12873, 16'd28657, 16'd25532, 16'd12052, 16'd7757, 16'd42232, 16'd17029, 16'd35762, 16'd18547, 16'd2042, 16'd2037, 16'd13300, 16'd49200, 16'd60781, 16'd14548, 16'd19358, 16'd20461, 16'd61837, 16'd35849, 16'd33730, 16'd40856, 16'd18043, 16'd41774, 16'd14475});
	test_expansion(128'haef0be344573d0bd3b196dfc9c1ac401, {16'd47917, 16'd19884, 16'd42422, 16'd14668, 16'd33207, 16'd47472, 16'd7101, 16'd137, 16'd39217, 16'd17384, 16'd26924, 16'd9884, 16'd59781, 16'd3823, 16'd7008, 16'd8829, 16'd40710, 16'd44191, 16'd11821, 16'd31378, 16'd53526, 16'd62244, 16'd53524, 16'd20010, 16'd26053, 16'd18747});
	test_expansion(128'hb1949f3cb8f6af0c8530afe340ed3083, {16'd61578, 16'd32710, 16'd23783, 16'd14906, 16'd33542, 16'd61967, 16'd1426, 16'd16677, 16'd55294, 16'd61604, 16'd41566, 16'd27475, 16'd29573, 16'd39872, 16'd20194, 16'd15293, 16'd51650, 16'd63633, 16'd44020, 16'd39253, 16'd29838, 16'd31182, 16'd5520, 16'd13345, 16'd33464, 16'd4142});
	test_expansion(128'h548e01676d50b67af1d55659488e835b, {16'd11551, 16'd11572, 16'd9557, 16'd21509, 16'd56312, 16'd13502, 16'd47332, 16'd17536, 16'd14206, 16'd15515, 16'd1654, 16'd36364, 16'd39023, 16'd27820, 16'd54710, 16'd11748, 16'd5401, 16'd52809, 16'd32541, 16'd3493, 16'd19422, 16'd13786, 16'd60855, 16'd15203, 16'd13316, 16'd34387});
	test_expansion(128'hec4f7ed12f33de72d7f74473d49b8afd, {16'd2444, 16'd59674, 16'd24537, 16'd1624, 16'd28650, 16'd63710, 16'd8922, 16'd31493, 16'd52581, 16'd48214, 16'd11221, 16'd29611, 16'd28472, 16'd19507, 16'd19916, 16'd30529, 16'd50998, 16'd30411, 16'd1855, 16'd7113, 16'd1722, 16'd41951, 16'd29427, 16'd34533, 16'd54890, 16'd24178});
	test_expansion(128'h4f586ae02050a03db3f9117f0509f1f7, {16'd56429, 16'd6465, 16'd40823, 16'd53519, 16'd19542, 16'd54095, 16'd44393, 16'd19259, 16'd57809, 16'd15759, 16'd53913, 16'd41638, 16'd38505, 16'd31991, 16'd41576, 16'd13979, 16'd31395, 16'd49244, 16'd50987, 16'd11470, 16'd51138, 16'd27401, 16'd5802, 16'd64789, 16'd2576, 16'd22530});
	test_expansion(128'h6d662efd945a0f9cbc721587b25e71cd, {16'd23925, 16'd55649, 16'd35632, 16'd39353, 16'd11429, 16'd4490, 16'd46744, 16'd51809, 16'd3060, 16'd50373, 16'd34360, 16'd57235, 16'd5388, 16'd7716, 16'd39326, 16'd39179, 16'd32266, 16'd29881, 16'd12538, 16'd28120, 16'd61926, 16'd16164, 16'd22894, 16'd16116, 16'd5959, 16'd25145});
	test_expansion(128'h89ac511af71de118311a86a6c10306fe, {16'd31113, 16'd14796, 16'd7066, 16'd52519, 16'd25440, 16'd29472, 16'd40045, 16'd6127, 16'd28147, 16'd11419, 16'd54956, 16'd2978, 16'd39233, 16'd27752, 16'd12999, 16'd44658, 16'd50926, 16'd44572, 16'd26537, 16'd5250, 16'd21362, 16'd52712, 16'd16853, 16'd17795, 16'd6443, 16'd51183});
	test_expansion(128'h2f1ebed4c6335ae6ace659ea76bb361d, {16'd57374, 16'd60026, 16'd54800, 16'd21990, 16'd62368, 16'd30646, 16'd16027, 16'd33662, 16'd63994, 16'd11526, 16'd44887, 16'd41799, 16'd28077, 16'd980, 16'd46220, 16'd20556, 16'd53743, 16'd10201, 16'd23468, 16'd40432, 16'd19133, 16'd6549, 16'd10968, 16'd14671, 16'd8025, 16'd38690});
	test_expansion(128'hb23c6e1660293cdf7df42016d8986022, {16'd1135, 16'd59802, 16'd64041, 16'd44314, 16'd44123, 16'd13339, 16'd54161, 16'd42446, 16'd4983, 16'd22264, 16'd62447, 16'd340, 16'd59706, 16'd8917, 16'd52062, 16'd28869, 16'd5351, 16'd18698, 16'd56690, 16'd49116, 16'd34688, 16'd1081, 16'd56723, 16'd22875, 16'd42433, 16'd35441});
	test_expansion(128'h1695879a27cf0203acadbb36e24648f1, {16'd38688, 16'd14354, 16'd62963, 16'd57496, 16'd52762, 16'd61457, 16'd58959, 16'd15000, 16'd5227, 16'd63353, 16'd29193, 16'd33427, 16'd51609, 16'd18999, 16'd36150, 16'd59054, 16'd34150, 16'd13324, 16'd12048, 16'd33668, 16'd56450, 16'd20084, 16'd50531, 16'd12376, 16'd59583, 16'd41360});
	test_expansion(128'h6680033d2e32a30ea25b841e4570be35, {16'd31839, 16'd48187, 16'd30805, 16'd28589, 16'd24493, 16'd65332, 16'd64831, 16'd35329, 16'd28854, 16'd57142, 16'd37273, 16'd35488, 16'd3932, 16'd12593, 16'd26009, 16'd54545, 16'd63217, 16'd63085, 16'd46818, 16'd50556, 16'd32366, 16'd33377, 16'd12712, 16'd32148, 16'd23986, 16'd50801});
	test_expansion(128'hdd842bea7b9b306409610d731d266258, {16'd43971, 16'd51966, 16'd64452, 16'd57199, 16'd30496, 16'd24093, 16'd57692, 16'd6217, 16'd61166, 16'd43756, 16'd54636, 16'd4056, 16'd3072, 16'd4475, 16'd41627, 16'd16679, 16'd40379, 16'd45136, 16'd29032, 16'd7630, 16'd19912, 16'd37595, 16'd17044, 16'd9878, 16'd45865, 16'd64148});
	test_expansion(128'hfde6ba160144e07beee2cd204fc6c091, {16'd3159, 16'd61964, 16'd34172, 16'd43908, 16'd50563, 16'd8277, 16'd6901, 16'd28475, 16'd22803, 16'd21328, 16'd31182, 16'd12506, 16'd59448, 16'd30992, 16'd34778, 16'd61424, 16'd24438, 16'd26147, 16'd1220, 16'd47540, 16'd33980, 16'd34707, 16'd53427, 16'd25453, 16'd44778, 16'd64036});
	test_expansion(128'h39456fdb7ccdb8ef2a448fa23fd0aa0d, {16'd32672, 16'd56725, 16'd19820, 16'd24958, 16'd64530, 16'd56746, 16'd8616, 16'd32516, 16'd6611, 16'd22041, 16'd54809, 16'd18644, 16'd6245, 16'd46415, 16'd18188, 16'd40505, 16'd59775, 16'd50069, 16'd39789, 16'd61782, 16'd64358, 16'd61198, 16'd18856, 16'd46965, 16'd21651, 16'd11546});
	test_expansion(128'h605b7e7925f6ad4c8388708e802d4193, {16'd27143, 16'd29215, 16'd3688, 16'd60736, 16'd36959, 16'd1237, 16'd37814, 16'd31378, 16'd37581, 16'd56710, 16'd58852, 16'd22859, 16'd57160, 16'd36402, 16'd9325, 16'd59726, 16'd51965, 16'd5811, 16'd694, 16'd35415, 16'd27084, 16'd42205, 16'd27380, 16'd47899, 16'd39934, 16'd27765});
	test_expansion(128'h30529fde3d73224b83b857d4284b9761, {16'd64179, 16'd16950, 16'd43741, 16'd1108, 16'd64109, 16'd20424, 16'd3812, 16'd40821, 16'd31266, 16'd59255, 16'd25382, 16'd49370, 16'd34960, 16'd20221, 16'd15153, 16'd65195, 16'd31998, 16'd8528, 16'd26370, 16'd52117, 16'd8995, 16'd51366, 16'd34838, 16'd15438, 16'd3183, 16'd5491});
	test_expansion(128'ha25b2568b700cf811238f66b1dc54332, {16'd50020, 16'd49992, 16'd58480, 16'd29327, 16'd50948, 16'd31402, 16'd39283, 16'd47558, 16'd1412, 16'd63178, 16'd31442, 16'd3105, 16'd40559, 16'd43309, 16'd19752, 16'd24873, 16'd61522, 16'd29189, 16'd560, 16'd30504, 16'd440, 16'd12662, 16'd52562, 16'd12925, 16'd57834, 16'd30922});
	test_expansion(128'hf504cc814574acb46c4d0fe91c4d5433, {16'd16146, 16'd4272, 16'd62514, 16'd13366, 16'd48077, 16'd3929, 16'd59577, 16'd25807, 16'd44189, 16'd59343, 16'd32895, 16'd33563, 16'd61928, 16'd45794, 16'd28589, 16'd7412, 16'd42223, 16'd27244, 16'd51137, 16'd47156, 16'd6337, 16'd31238, 16'd21329, 16'd21016, 16'd49938, 16'd56369});
	test_expansion(128'h90e4a1c1ddf81200f36817ed7b39eecd, {16'd8604, 16'd1156, 16'd26504, 16'd12798, 16'd11294, 16'd55523, 16'd27225, 16'd58291, 16'd14764, 16'd42218, 16'd7422, 16'd14018, 16'd12554, 16'd44122, 16'd20154, 16'd62258, 16'd64884, 16'd42307, 16'd38860, 16'd29677, 16'd17785, 16'd37977, 16'd38748, 16'd63285, 16'd6530, 16'd36});
	test_expansion(128'h0f8ee7da42497dceb48895302b0c3a26, {16'd54034, 16'd11387, 16'd28277, 16'd51611, 16'd55001, 16'd42288, 16'd5699, 16'd6281, 16'd61348, 16'd26292, 16'd50951, 16'd37635, 16'd42182, 16'd51217, 16'd16612, 16'd52911, 16'd24534, 16'd45425, 16'd46056, 16'd36130, 16'd58647, 16'd53947, 16'd27663, 16'd12530, 16'd45460, 16'd13865});
	test_expansion(128'h3eca1507b0c247c4a892801ca4291ecb, {16'd17679, 16'd49357, 16'd10728, 16'd1428, 16'd52807, 16'd46328, 16'd64752, 16'd26872, 16'd40933, 16'd5662, 16'd21231, 16'd24164, 16'd50950, 16'd7664, 16'd35794, 16'd37295, 16'd65034, 16'd55245, 16'd51560, 16'd15278, 16'd50012, 16'd47196, 16'd31847, 16'd32178, 16'd48349, 16'd61348});
	test_expansion(128'hda65b7aafbdb8625109490860c92e1bb, {16'd50507, 16'd57678, 16'd18837, 16'd8787, 16'd50955, 16'd7202, 16'd43667, 16'd29633, 16'd1290, 16'd47156, 16'd14667, 16'd27592, 16'd38538, 16'd59591, 16'd18079, 16'd14053, 16'd38051, 16'd30953, 16'd48310, 16'd7120, 16'd1274, 16'd40290, 16'd1183, 16'd4082, 16'd24155, 16'd12432});
	test_expansion(128'hd07fd6d845855cf764bf0aa1515c4da1, {16'd57570, 16'd44262, 16'd54168, 16'd29312, 16'd37026, 16'd35308, 16'd41817, 16'd16349, 16'd23978, 16'd15544, 16'd21170, 16'd57516, 16'd64747, 16'd34134, 16'd22822, 16'd41860, 16'd38981, 16'd31644, 16'd43698, 16'd32572, 16'd39358, 16'd39089, 16'd61562, 16'd60745, 16'd49676, 16'd32038});
	test_expansion(128'h4a7bb9ae4f91e1a8cb59b3408442a23c, {16'd65338, 16'd13943, 16'd12312, 16'd18709, 16'd61635, 16'd4166, 16'd248, 16'd36316, 16'd16033, 16'd6035, 16'd51407, 16'd46560, 16'd26263, 16'd23030, 16'd63815, 16'd2108, 16'd37802, 16'd22862, 16'd362, 16'd3370, 16'd57017, 16'd22349, 16'd31054, 16'd10983, 16'd54354, 16'd52829});
	test_expansion(128'h9671c1311a8f0b85e43d260d649a82ce, {16'd26200, 16'd47674, 16'd11805, 16'd30459, 16'd30415, 16'd42235, 16'd41037, 16'd27457, 16'd24039, 16'd54815, 16'd30384, 16'd36205, 16'd45707, 16'd60998, 16'd2276, 16'd57631, 16'd52444, 16'd4590, 16'd20695, 16'd40714, 16'd57494, 16'd32785, 16'd9401, 16'd32120, 16'd3343, 16'd33635});
	test_expansion(128'h0470d21cdd23d8e30114f0963a9cc64c, {16'd7923, 16'd13756, 16'd33098, 16'd52464, 16'd33912, 16'd63753, 16'd10892, 16'd55184, 16'd43173, 16'd63488, 16'd40625, 16'd18302, 16'd8564, 16'd41919, 16'd17956, 16'd50324, 16'd18265, 16'd25151, 16'd8385, 16'd27361, 16'd46320, 16'd3015, 16'd43899, 16'd64137, 16'd37191, 16'd59822});
	test_expansion(128'h97bbb361d7ecb32ced01ee8958e5b9d3, {16'd52577, 16'd60885, 16'd24961, 16'd37304, 16'd17200, 16'd22440, 16'd22895, 16'd61240, 16'd11552, 16'd34389, 16'd21639, 16'd49157, 16'd37972, 16'd11101, 16'd23244, 16'd7013, 16'd11559, 16'd49672, 16'd9168, 16'd29017, 16'd41927, 16'd6687, 16'd35883, 16'd45074, 16'd51142, 16'd62442});
	test_expansion(128'h93af31fa04ae43e74c40a666d60da96d, {16'd1405, 16'd46280, 16'd45573, 16'd18194, 16'd26983, 16'd64166, 16'd19406, 16'd22562, 16'd1922, 16'd6415, 16'd62000, 16'd46288, 16'd17949, 16'd30703, 16'd36006, 16'd44170, 16'd10454, 16'd2292, 16'd41935, 16'd22120, 16'd58912, 16'd46735, 16'd41264, 16'd41092, 16'd23025, 16'd12899});
	test_expansion(128'h0dd4e1adbfccb565cc219f8fe0531337, {16'd7793, 16'd20302, 16'd44614, 16'd46697, 16'd28066, 16'd5944, 16'd9292, 16'd38142, 16'd46191, 16'd44566, 16'd25540, 16'd32061, 16'd41014, 16'd58665, 16'd7268, 16'd4947, 16'd64116, 16'd64294, 16'd40617, 16'd20098, 16'd27544, 16'd38237, 16'd28902, 16'd36673, 16'd39243, 16'd17058});
	test_expansion(128'he57f6e8c41050955a6ed5e1ea4ac51eb, {16'd26690, 16'd57741, 16'd2690, 16'd31693, 16'd4514, 16'd24452, 16'd12747, 16'd50233, 16'd23101, 16'd18917, 16'd51901, 16'd64501, 16'd11598, 16'd8178, 16'd31736, 16'd17674, 16'd23291, 16'd48046, 16'd47029, 16'd2338, 16'd23665, 16'd42030, 16'd6266, 16'd27403, 16'd25611, 16'd14894});
	test_expansion(128'h057cdbcd2fdc5349e57b8dd1f34977dd, {16'd34738, 16'd22025, 16'd46445, 16'd38066, 16'd55665, 16'd2752, 16'd34975, 16'd64716, 16'd30017, 16'd44115, 16'd64734, 16'd22496, 16'd36300, 16'd61391, 16'd15991, 16'd36143, 16'd55082, 16'd19936, 16'd49579, 16'd34991, 16'd50112, 16'd6997, 16'd35368, 16'd62483, 16'd31037, 16'd29422});
	test_expansion(128'h1ce9d6e2dd8a6a241200dfa92a1e64e9, {16'd13240, 16'd48966, 16'd42001, 16'd12184, 16'd20281, 16'd36899, 16'd32935, 16'd30681, 16'd36746, 16'd5107, 16'd51620, 16'd10136, 16'd18977, 16'd62466, 16'd688, 16'd40843, 16'd25680, 16'd54746, 16'd37731, 16'd2973, 16'd6281, 16'd4038, 16'd48859, 16'd23276, 16'd59773, 16'd57710});
	test_expansion(128'h5344d3e299f1996c10a39f54f9de01a7, {16'd20837, 16'd13111, 16'd13243, 16'd43610, 16'd17453, 16'd17051, 16'd49068, 16'd7136, 16'd51885, 16'd16660, 16'd28369, 16'd53449, 16'd28282, 16'd64703, 16'd64599, 16'd2931, 16'd30000, 16'd60606, 16'd40125, 16'd48978, 16'd30956, 16'd53934, 16'd34698, 16'd63144, 16'd43029, 16'd16343});
	test_expansion(128'h93625706dc0b9ae14ad700a148ce8033, {16'd41590, 16'd25911, 16'd9948, 16'd23297, 16'd43946, 16'd1517, 16'd24041, 16'd52202, 16'd34678, 16'd31650, 16'd41551, 16'd17216, 16'd34297, 16'd43981, 16'd44692, 16'd1568, 16'd27013, 16'd3768, 16'd62880, 16'd62635, 16'd23870, 16'd49606, 16'd12382, 16'd11584, 16'd63776, 16'd36492});
	test_expansion(128'h9aafb2e499a46073f2decc3fc1c76d50, {16'd47530, 16'd56195, 16'd63108, 16'd53041, 16'd10408, 16'd10732, 16'd57266, 16'd18563, 16'd47699, 16'd46913, 16'd60518, 16'd34783, 16'd30212, 16'd51599, 16'd9014, 16'd8705, 16'd37810, 16'd27696, 16'd13924, 16'd21060, 16'd3118, 16'd55565, 16'd17586, 16'd24695, 16'd29859, 16'd20040});
	test_expansion(128'h88e104d06a33a4b48f5a59c5c356788d, {16'd22526, 16'd4125, 16'd7758, 16'd34711, 16'd15237, 16'd63378, 16'd58694, 16'd35258, 16'd64325, 16'd61084, 16'd41148, 16'd10174, 16'd43167, 16'd42714, 16'd43798, 16'd4569, 16'd59636, 16'd43702, 16'd31620, 16'd30650, 16'd54742, 16'd33981, 16'd27014, 16'd47465, 16'd43596, 16'd29814});
	test_expansion(128'h519e78cbeba00419cb33efe6c98cdd41, {16'd60972, 16'd38351, 16'd2408, 16'd11397, 16'd37771, 16'd27901, 16'd51194, 16'd5168, 16'd41060, 16'd21341, 16'd40026, 16'd27993, 16'd65527, 16'd62738, 16'd11339, 16'd64670, 16'd47255, 16'd60363, 16'd64864, 16'd28585, 16'd20145, 16'd44824, 16'd12408, 16'd62991, 16'd33570, 16'd26785});
	test_expansion(128'h5b377f3d10cfa1efb1539efcf9e3ce2b, {16'd28099, 16'd2151, 16'd6833, 16'd42767, 16'd34915, 16'd51995, 16'd50580, 16'd65498, 16'd61474, 16'd28984, 16'd42450, 16'd33282, 16'd44676, 16'd7257, 16'd11485, 16'd38973, 16'd40787, 16'd13555, 16'd51541, 16'd12185, 16'd21915, 16'd20472, 16'd39637, 16'd22613, 16'd7302, 16'd11065});
	test_expansion(128'h7f838a2fcebaaa4b59c16a434090adf0, {16'd16549, 16'd63032, 16'd8515, 16'd45921, 16'd38703, 16'd17309, 16'd41350, 16'd21784, 16'd9632, 16'd30224, 16'd3279, 16'd2922, 16'd32822, 16'd45130, 16'd50597, 16'd62633, 16'd18762, 16'd30285, 16'd20001, 16'd8413, 16'd48308, 16'd7642, 16'd32606, 16'd13466, 16'd25870, 16'd26463});
	test_expansion(128'h6c5ffe1b9b0b0095533b04671e80531b, {16'd60667, 16'd49202, 16'd8928, 16'd49534, 16'd43585, 16'd37774, 16'd21871, 16'd29173, 16'd18020, 16'd9008, 16'd15889, 16'd41948, 16'd55918, 16'd54284, 16'd59210, 16'd13820, 16'd58977, 16'd24418, 16'd33517, 16'd6033, 16'd5727, 16'd58626, 16'd59019, 16'd29407, 16'd12988, 16'd33661});
	test_expansion(128'h52c5ab64898174778354334917b1e24b, {16'd12900, 16'd21405, 16'd8548, 16'd31945, 16'd33978, 16'd10022, 16'd25694, 16'd8337, 16'd34025, 16'd41836, 16'd33193, 16'd7465, 16'd34182, 16'd21955, 16'd17752, 16'd21930, 16'd56849, 16'd13935, 16'd22004, 16'd34792, 16'd25341, 16'd28429, 16'd62314, 16'd3578, 16'd5078, 16'd28422});
	test_expansion(128'h1adaf7fe5b09487695173b45eab3cacf, {16'd13233, 16'd9470, 16'd18289, 16'd22597, 16'd28654, 16'd10535, 16'd50459, 16'd21589, 16'd24482, 16'd11951, 16'd52330, 16'd59049, 16'd37499, 16'd9709, 16'd11702, 16'd19726, 16'd64818, 16'd57848, 16'd28870, 16'd54404, 16'd24458, 16'd12290, 16'd8420, 16'd26025, 16'd9619, 16'd52372});
	test_expansion(128'hfe72e6ea4a623fecb47de5d79baf920a, {16'd2527, 16'd45589, 16'd15016, 16'd20923, 16'd60374, 16'd35179, 16'd44893, 16'd19389, 16'd39026, 16'd21514, 16'd8666, 16'd36854, 16'd21247, 16'd6401, 16'd26996, 16'd16451, 16'd9044, 16'd57633, 16'd23033, 16'd2911, 16'd17274, 16'd28558, 16'd34206, 16'd35045, 16'd3652, 16'd33465});
	test_expansion(128'h6d1956ae529494b241c65b21709e6182, {16'd10307, 16'd13975, 16'd15232, 16'd43744, 16'd28368, 16'd9147, 16'd28813, 16'd65432, 16'd13966, 16'd23015, 16'd56101, 16'd49339, 16'd18761, 16'd42490, 16'd63722, 16'd64767, 16'd3447, 16'd28510, 16'd4252, 16'd43605, 16'd39147, 16'd46421, 16'd53041, 16'd18191, 16'd20947, 16'd760});
	test_expansion(128'ha7a38997a1bf54b0fa390a3a4e34e1de, {16'd45102, 16'd29704, 16'd35440, 16'd43450, 16'd35671, 16'd22384, 16'd11112, 16'd49241, 16'd12675, 16'd27410, 16'd22715, 16'd9477, 16'd38233, 16'd11611, 16'd34343, 16'd30010, 16'd11422, 16'd40218, 16'd38474, 16'd49322, 16'd48802, 16'd18027, 16'd53510, 16'd24073, 16'd28675, 16'd53050});
	test_expansion(128'h980a0074c2ed454c8aa045949861c9fd, {16'd60943, 16'd52658, 16'd18277, 16'd53833, 16'd48428, 16'd59162, 16'd49600, 16'd23454, 16'd26820, 16'd39775, 16'd39968, 16'd41546, 16'd56892, 16'd22970, 16'd42876, 16'd46447, 16'd39184, 16'd53426, 16'd14223, 16'd52640, 16'd56974, 16'd39801, 16'd34684, 16'd15227, 16'd36999, 16'd39895});
	test_expansion(128'hed9045bee533640b3fe0d5e7951379c8, {16'd30611, 16'd12387, 16'd10277, 16'd11046, 16'd52511, 16'd27255, 16'd19227, 16'd12253, 16'd7038, 16'd4614, 16'd61361, 16'd24186, 16'd46456, 16'd16238, 16'd1785, 16'd6345, 16'd157, 16'd55382, 16'd39012, 16'd44798, 16'd46131, 16'd18829, 16'd4516, 16'd36263, 16'd51806, 16'd41612});
	test_expansion(128'hd5b432d540a24bd2e595f6ca81526371, {16'd14034, 16'd20334, 16'd52975, 16'd5773, 16'd33909, 16'd12336, 16'd7403, 16'd48783, 16'd48710, 16'd38373, 16'd12831, 16'd4045, 16'd14687, 16'd21416, 16'd27028, 16'd27778, 16'd38168, 16'd27828, 16'd59926, 16'd23829, 16'd6033, 16'd20081, 16'd64813, 16'd23100, 16'd4790, 16'd35756});
	test_expansion(128'hf081994c5d97b9c39e82a841cdc0b9f6, {16'd24081, 16'd56389, 16'd23192, 16'd25105, 16'd56834, 16'd1922, 16'd36088, 16'd28942, 16'd3104, 16'd7569, 16'd61023, 16'd34669, 16'd30362, 16'd42171, 16'd6516, 16'd53457, 16'd28765, 16'd33590, 16'd52966, 16'd10346, 16'd9367, 16'd16019, 16'd62017, 16'd23203, 16'd65490, 16'd53510});
	test_expansion(128'h09f7efb87c37c1a1a35be6eeb034402c, {16'd708, 16'd59178, 16'd53528, 16'd46055, 16'd7244, 16'd20200, 16'd46037, 16'd6512, 16'd19853, 16'd20166, 16'd34284, 16'd56102, 16'd17363, 16'd63072, 16'd62945, 16'd3915, 16'd38109, 16'd60363, 16'd48158, 16'd16064, 16'd36005, 16'd46716, 16'd48152, 16'd27936, 16'd31174, 16'd4918});
	test_expansion(128'h6d0e40ec71ef8bc54b475cb1aaef9f06, {16'd17879, 16'd38272, 16'd20498, 16'd16167, 16'd59298, 16'd4941, 16'd56671, 16'd63082, 16'd40073, 16'd26822, 16'd1721, 16'd54319, 16'd48998, 16'd1666, 16'd30605, 16'd2533, 16'd56467, 16'd56914, 16'd525, 16'd26545, 16'd36661, 16'd42939, 16'd946, 16'd21983, 16'd58716, 16'd45738});
	test_expansion(128'h5ec7947bdac9282391cdfaa5e97c1507, {16'd61251, 16'd6188, 16'd61963, 16'd60175, 16'd61824, 16'd30424, 16'd20630, 16'd29294, 16'd53249, 16'd35879, 16'd5201, 16'd49597, 16'd62300, 16'd32045, 16'd10890, 16'd54646, 16'd65460, 16'd45691, 16'd35451, 16'd37512, 16'd17574, 16'd13381, 16'd28925, 16'd41277, 16'd33223, 16'd32660});
	test_expansion(128'h8655df433044e76bd8d47d9048d6e7b3, {16'd47200, 16'd19227, 16'd15971, 16'd5196, 16'd44203, 16'd17088, 16'd47859, 16'd12855, 16'd16250, 16'd17431, 16'd53035, 16'd59434, 16'd4457, 16'd51559, 16'd65490, 16'd26459, 16'd12761, 16'd22055, 16'd32741, 16'd48861, 16'd7672, 16'd17309, 16'd56277, 16'd16433, 16'd23029, 16'd41281});
	test_expansion(128'hdf7b86595f599d8832a9c526ff490cdc, {16'd16363, 16'd63705, 16'd19322, 16'd31491, 16'd60810, 16'd36900, 16'd54108, 16'd60571, 16'd44472, 16'd31569, 16'd47874, 16'd49966, 16'd40865, 16'd11257, 16'd60632, 16'd27851, 16'd10404, 16'd24578, 16'd6491, 16'd8745, 16'd3580, 16'd39550, 16'd20779, 16'd31228, 16'd53209, 16'd6491});
	test_expansion(128'h7c345a1fb6c5d11a13221ebd19cf677e, {16'd7949, 16'd31482, 16'd11620, 16'd60752, 16'd16005, 16'd42173, 16'd62157, 16'd59368, 16'd48243, 16'd59145, 16'd42434, 16'd60120, 16'd14994, 16'd2514, 16'd38753, 16'd62329, 16'd60612, 16'd12294, 16'd15736, 16'd45257, 16'd10580, 16'd63488, 16'd45831, 16'd50943, 16'd4247, 16'd39006});
	test_expansion(128'h7198c8c18c975aba276bbf4f9033cf7b, {16'd44555, 16'd8354, 16'd47996, 16'd61309, 16'd30977, 16'd46130, 16'd39875, 16'd24834, 16'd34585, 16'd19915, 16'd40138, 16'd40652, 16'd44182, 16'd35800, 16'd63996, 16'd49504, 16'd3118, 16'd21919, 16'd45039, 16'd33166, 16'd27891, 16'd51260, 16'd27066, 16'd11612, 16'd15101, 16'd17652});
	test_expansion(128'h01eb9816e21f6c1d7d6d73d3db6f1e4d, {16'd1950, 16'd51547, 16'd40643, 16'd28399, 16'd39957, 16'd11464, 16'd51704, 16'd63894, 16'd65356, 16'd38238, 16'd34080, 16'd58542, 16'd378, 16'd11658, 16'd20452, 16'd34890, 16'd31267, 16'd44954, 16'd32031, 16'd52938, 16'd6084, 16'd19101, 16'd41090, 16'd50489, 16'd62584, 16'd36604});
	test_expansion(128'h23f394cc433bffc07c9f478309c6e9b6, {16'd25952, 16'd62902, 16'd37105, 16'd4047, 16'd60272, 16'd15187, 16'd52683, 16'd63, 16'd48821, 16'd65324, 16'd34086, 16'd16900, 16'd17367, 16'd63149, 16'd28331, 16'd31974, 16'd28662, 16'd37008, 16'd12555, 16'd4722, 16'd14728, 16'd6152, 16'd40572, 16'd40986, 16'd2295, 16'd20131});
	test_expansion(128'h718c7913048ff13c9533865190bfbf3a, {16'd57369, 16'd29974, 16'd63991, 16'd3761, 16'd5017, 16'd38685, 16'd53129, 16'd55277, 16'd59288, 16'd23711, 16'd12785, 16'd18667, 16'd30920, 16'd43705, 16'd32307, 16'd61125, 16'd50288, 16'd41886, 16'd57646, 16'd32814, 16'd53046, 16'd44941, 16'd13647, 16'd26728, 16'd9376, 16'd55351});
	test_expansion(128'hc82cdbabddc03d1c382319357f8dffa5, {16'd5560, 16'd12481, 16'd7748, 16'd11152, 16'd32211, 16'd58790, 16'd63967, 16'd44343, 16'd12928, 16'd1366, 16'd16055, 16'd55904, 16'd56657, 16'd27139, 16'd65296, 16'd2848, 16'd36783, 16'd61751, 16'd53792, 16'd60104, 16'd45435, 16'd53667, 16'd53858, 16'd9952, 16'd31562, 16'd10716});
	test_expansion(128'h72e713f0b8b2bd17e59614f99d73fc83, {16'd2962, 16'd10715, 16'd50943, 16'd22744, 16'd32761, 16'd55245, 16'd65327, 16'd24682, 16'd28835, 16'd17447, 16'd23145, 16'd12353, 16'd32874, 16'd51072, 16'd27853, 16'd58303, 16'd42715, 16'd11545, 16'd43481, 16'd44479, 16'd24247, 16'd19520, 16'd37702, 16'd59503, 16'd599, 16'd32909});
	test_expansion(128'hd4d047d8e9dc252551a8c5a1f641e845, {16'd37966, 16'd60345, 16'd4803, 16'd16689, 16'd50814, 16'd64785, 16'd24383, 16'd38457, 16'd48112, 16'd377, 16'd55467, 16'd9605, 16'd60360, 16'd40185, 16'd32480, 16'd36306, 16'd38522, 16'd10330, 16'd34714, 16'd57994, 16'd10147, 16'd36037, 16'd59845, 16'd19450, 16'd53503, 16'd26456});
	test_expansion(128'h27d8e6bee44e18a0de24bbc0b0fa4f55, {16'd46585, 16'd3972, 16'd39807, 16'd35101, 16'd18976, 16'd6279, 16'd43105, 16'd14581, 16'd704, 16'd59669, 16'd40892, 16'd64615, 16'd52694, 16'd34730, 16'd64491, 16'd46732, 16'd39046, 16'd3052, 16'd24899, 16'd30794, 16'd59583, 16'd64918, 16'd2903, 16'd39687, 16'd24752, 16'd21305});
	test_expansion(128'h0615568f315569eb7753d30de674bbd8, {16'd52296, 16'd16905, 16'd2087, 16'd21, 16'd8061, 16'd13010, 16'd34469, 16'd22683, 16'd133, 16'd42449, 16'd45219, 16'd45060, 16'd65022, 16'd30714, 16'd22364, 16'd20550, 16'd58501, 16'd22024, 16'd18902, 16'd29090, 16'd62063, 16'd15796, 16'd5557, 16'd35426, 16'd18695, 16'd56414});
	test_expansion(128'hef3e65074992283f54bba6675b6b4d7a, {16'd23061, 16'd47199, 16'd42007, 16'd8109, 16'd45377, 16'd39922, 16'd36307, 16'd27712, 16'd39219, 16'd61621, 16'd13211, 16'd17795, 16'd56724, 16'd51962, 16'd62170, 16'd62014, 16'd31690, 16'd54433, 16'd44169, 16'd50474, 16'd9410, 16'd54290, 16'd53501, 16'd17621, 16'd61945, 16'd52632});
	test_expansion(128'h107fbe7748bbb2d2f1c3ab59b84e935b, {16'd27514, 16'd62142, 16'd54327, 16'd35030, 16'd41005, 16'd64097, 16'd19130, 16'd22892, 16'd7574, 16'd42323, 16'd14804, 16'd12838, 16'd49377, 16'd57442, 16'd44404, 16'd55693, 16'd61126, 16'd56152, 16'd40090, 16'd44571, 16'd26106, 16'd60035, 16'd34320, 16'd31670, 16'd24625, 16'd38023});
	test_expansion(128'h466186f4df358278bb5357435de33267, {16'd52620, 16'd6614, 16'd61616, 16'd36368, 16'd14261, 16'd21909, 16'd25726, 16'd4005, 16'd30602, 16'd10134, 16'd32233, 16'd37307, 16'd36073, 16'd42215, 16'd64977, 16'd4904, 16'd45795, 16'd52088, 16'd2524, 16'd38111, 16'd14198, 16'd10596, 16'd36877, 16'd33799, 16'd1246, 16'd33269});
	test_expansion(128'h71486e373c9cda307b68d41fb4f091b2, {16'd49715, 16'd46819, 16'd5759, 16'd12733, 16'd55349, 16'd35798, 16'd7094, 16'd41473, 16'd35633, 16'd26784, 16'd46880, 16'd6940, 16'd21629, 16'd48079, 16'd39970, 16'd7942, 16'd21464, 16'd13659, 16'd22884, 16'd24374, 16'd17430, 16'd62087, 16'd50889, 16'd60993, 16'd3745, 16'd7860});
	test_expansion(128'hbdca3551560cddcbe4a23deaff2cc9f8, {16'd55889, 16'd39758, 16'd4130, 16'd36646, 16'd40766, 16'd58922, 16'd4696, 16'd33574, 16'd62604, 16'd27392, 16'd39830, 16'd18944, 16'd58679, 16'd63601, 16'd10774, 16'd38362, 16'd45242, 16'd34304, 16'd11733, 16'd8470, 16'd59484, 16'd40839, 16'd41195, 16'd53358, 16'd22638, 16'd50027});
	test_expansion(128'h9a6ffb26a7da1a02751b8b3e8950f915, {16'd32149, 16'd3444, 16'd59475, 16'd30832, 16'd62677, 16'd36608, 16'd44484, 16'd53273, 16'd20278, 16'd33879, 16'd11341, 16'd29875, 16'd56557, 16'd58093, 16'd34157, 16'd10431, 16'd1685, 16'd22131, 16'd6454, 16'd18209, 16'd40206, 16'd41600, 16'd56878, 16'd3571, 16'd12378, 16'd3312});
	test_expansion(128'hd89907b892b76821596a44685e9e7b9f, {16'd12299, 16'd4515, 16'd62525, 16'd43644, 16'd54703, 16'd17503, 16'd11513, 16'd27712, 16'd64048, 16'd55365, 16'd23000, 16'd22029, 16'd51469, 16'd209, 16'd38725, 16'd38545, 16'd47050, 16'd48525, 16'd21495, 16'd45328, 16'd42660, 16'd39512, 16'd62458, 16'd1987, 16'd36263, 16'd11326});
	test_expansion(128'h011ac850fa0f4c07fb55076c7ae382a2, {16'd61557, 16'd21401, 16'd1854, 16'd6959, 16'd57867, 16'd37946, 16'd56656, 16'd61720, 16'd732, 16'd21868, 16'd17971, 16'd15495, 16'd36718, 16'd17954, 16'd11684, 16'd25173, 16'd3426, 16'd59065, 16'd37881, 16'd60758, 16'd47392, 16'd10031, 16'd15631, 16'd31265, 16'd50374, 16'd64895});
	test_expansion(128'h08f308e4fdddfbd7369378a4b15f50aa, {16'd2278, 16'd38689, 16'd41871, 16'd62539, 16'd4686, 16'd44951, 16'd34335, 16'd6192, 16'd42015, 16'd45463, 16'd60252, 16'd40685, 16'd33674, 16'd5474, 16'd38452, 16'd56616, 16'd33299, 16'd28481, 16'd46435, 16'd43583, 16'd23527, 16'd24081, 16'd57803, 16'd36042, 16'd57137, 16'd32281});
	test_expansion(128'h270396363c86acdd088071c485124ad4, {16'd21809, 16'd65104, 16'd49198, 16'd23971, 16'd11130, 16'd31371, 16'd20020, 16'd20435, 16'd20351, 16'd50746, 16'd8018, 16'd5010, 16'd41744, 16'd40498, 16'd1033, 16'd24724, 16'd60461, 16'd42241, 16'd34423, 16'd49636, 16'd26962, 16'd39240, 16'd50708, 16'd10969, 16'd38739, 16'd37674});
	test_expansion(128'h73477e1ff6a9c49b97d2771af1d0464a, {16'd10521, 16'd22612, 16'd30244, 16'd8056, 16'd22260, 16'd43241, 16'd44896, 16'd10325, 16'd55999, 16'd27434, 16'd25002, 16'd28094, 16'd40164, 16'd64940, 16'd52412, 16'd63833, 16'd22955, 16'd43189, 16'd23383, 16'd63146, 16'd64468, 16'd63448, 16'd65143, 16'd545, 16'd44947, 16'd29623});
	test_expansion(128'hc0781b2f428c32644d5d96c8bb80ace9, {16'd9424, 16'd32776, 16'd22430, 16'd49641, 16'd64499, 16'd56241, 16'd31064, 16'd8840, 16'd50128, 16'd53577, 16'd49650, 16'd16054, 16'd20963, 16'd31571, 16'd48238, 16'd6373, 16'd54130, 16'd9128, 16'd33011, 16'd4219, 16'd30803, 16'd10091, 16'd19812, 16'd49245, 16'd32275, 16'd15220});
	test_expansion(128'hf77ec7f578597b6fc6410c2098b51ce9, {16'd10345, 16'd56055, 16'd61623, 16'd43053, 16'd59076, 16'd36778, 16'd822, 16'd61088, 16'd47694, 16'd28573, 16'd9487, 16'd32370, 16'd10742, 16'd27824, 16'd49583, 16'd38857, 16'd12766, 16'd29044, 16'd3852, 16'd39595, 16'd42107, 16'd10748, 16'd59408, 16'd50837, 16'd63813, 16'd36363});
	test_expansion(128'h8b3085c20fc9454d3a8e543c8b95bbf1, {16'd64080, 16'd7038, 16'd17027, 16'd35028, 16'd55075, 16'd23260, 16'd50225, 16'd31781, 16'd58308, 16'd54332, 16'd24314, 16'd37711, 16'd13162, 16'd31816, 16'd62282, 16'd45822, 16'd30559, 16'd63931, 16'd6280, 16'd57863, 16'd61605, 16'd891, 16'd44205, 16'd31411, 16'd63306, 16'd6462});
	test_expansion(128'h0b70f92df1a0487025432028a131998b, {16'd33787, 16'd60446, 16'd53716, 16'd2044, 16'd13078, 16'd62988, 16'd756, 16'd19078, 16'd49030, 16'd30407, 16'd41341, 16'd51455, 16'd34890, 16'd50604, 16'd54292, 16'd11871, 16'd47646, 16'd42129, 16'd43699, 16'd36914, 16'd51219, 16'd8357, 16'd19088, 16'd4571, 16'd31067, 16'd16707});
	test_expansion(128'h3506f87deebf67ce0a2f0167ed602698, {16'd51373, 16'd1917, 16'd44096, 16'd58243, 16'd17461, 16'd20363, 16'd55610, 16'd57590, 16'd65340, 16'd5165, 16'd58014, 16'd61658, 16'd23643, 16'd50269, 16'd58893, 16'd44459, 16'd61860, 16'd47577, 16'd56140, 16'd30339, 16'd26993, 16'd42874, 16'd27978, 16'd14289, 16'd62164, 16'd64785});
	test_expansion(128'hb0ca3204ff10caf57f2194c94634f35e, {16'd3953, 16'd56667, 16'd40520, 16'd18709, 16'd23599, 16'd22167, 16'd20963, 16'd45636, 16'd10240, 16'd53621, 16'd24882, 16'd44205, 16'd11496, 16'd15433, 16'd497, 16'd42458, 16'd31623, 16'd33057, 16'd6555, 16'd45475, 16'd63759, 16'd20368, 16'd17280, 16'd49369, 16'd5932, 16'd31985});
	test_expansion(128'h0514cf0b23294d48f07ed940c5559313, {16'd51237, 16'd7970, 16'd60492, 16'd3012, 16'd62086, 16'd39241, 16'd10863, 16'd3568, 16'd21789, 16'd7875, 16'd36588, 16'd64320, 16'd37181, 16'd15410, 16'd43836, 16'd28764, 16'd59745, 16'd44853, 16'd24132, 16'd60046, 16'd63913, 16'd30680, 16'd52068, 16'd15490, 16'd33088, 16'd12424});
	test_expansion(128'hff7181ed8eec5f601586a8cbb3b56081, {16'd52079, 16'd38229, 16'd35039, 16'd55061, 16'd22548, 16'd60889, 16'd46484, 16'd53182, 16'd29830, 16'd55189, 16'd28632, 16'd9198, 16'd65224, 16'd46232, 16'd52255, 16'd35817, 16'd23032, 16'd62130, 16'd52693, 16'd60576, 16'd6980, 16'd21891, 16'd61776, 16'd55721, 16'd37994, 16'd22600});
	test_expansion(128'h9fbb1fd133bc907b8f94115601da5cb6, {16'd32900, 16'd26690, 16'd26077, 16'd15521, 16'd25976, 16'd27187, 16'd44622, 16'd59837, 16'd19626, 16'd8967, 16'd47943, 16'd17229, 16'd41116, 16'd64106, 16'd39573, 16'd49284, 16'd23097, 16'd36934, 16'd7780, 16'd11743, 16'd28491, 16'd646, 16'd26929, 16'd55988, 16'd20162, 16'd44425});
	test_expansion(128'hcc980b1987b26611362ec89ca671a492, {16'd7638, 16'd1405, 16'd749, 16'd12882, 16'd49603, 16'd7045, 16'd41877, 16'd12980, 16'd32463, 16'd32492, 16'd47462, 16'd14852, 16'd32858, 16'd40694, 16'd44159, 16'd28032, 16'd64731, 16'd27152, 16'd57247, 16'd4255, 16'd32698, 16'd21453, 16'd59736, 16'd31037, 16'd2889, 16'd43911});
	test_expansion(128'h2458188b2448a1dfa251c6ebdb0aee3a, {16'd28228, 16'd51951, 16'd10732, 16'd31314, 16'd62968, 16'd47825, 16'd61423, 16'd39886, 16'd18712, 16'd39217, 16'd32239, 16'd47780, 16'd56729, 16'd33585, 16'd9222, 16'd47110, 16'd14217, 16'd56205, 16'd50596, 16'd25009, 16'd13005, 16'd16703, 16'd26936, 16'd5564, 16'd31578, 16'd33269});
	test_expansion(128'h9cb6b20e4522e872bf551c72a17d4d8d, {16'd25478, 16'd57128, 16'd31189, 16'd2402, 16'd550, 16'd34107, 16'd30933, 16'd38104, 16'd6204, 16'd54295, 16'd27693, 16'd25762, 16'd6849, 16'd63717, 16'd46146, 16'd22382, 16'd27076, 16'd23445, 16'd4084, 16'd62654, 16'd39345, 16'd21182, 16'd2139, 16'd58606, 16'd63360, 16'd36109});
	test_expansion(128'h8063cd202aafde9f87845783f3dacd6b, {16'd14083, 16'd54499, 16'd11708, 16'd53795, 16'd8773, 16'd38851, 16'd43688, 16'd44437, 16'd48878, 16'd30511, 16'd53779, 16'd26246, 16'd56040, 16'd58044, 16'd40868, 16'd36603, 16'd4751, 16'd55484, 16'd61261, 16'd48810, 16'd612, 16'd32222, 16'd60018, 16'd20570, 16'd33814, 16'd9644});
	test_expansion(128'h590c4d806bd9ed2506d510361340fdb2, {16'd58531, 16'd62746, 16'd61095, 16'd57273, 16'd22224, 16'd51420, 16'd28566, 16'd34052, 16'd44950, 16'd20139, 16'd51784, 16'd62676, 16'd49644, 16'd15657, 16'd17278, 16'd16547, 16'd39402, 16'd7377, 16'd6832, 16'd45147, 16'd35325, 16'd42496, 16'd17472, 16'd45638, 16'd18028, 16'd38820});
	test_expansion(128'had49a29e1cc8196cc7a351b90226628d, {16'd1100, 16'd37638, 16'd56266, 16'd55816, 16'd12682, 16'd22146, 16'd19782, 16'd23755, 16'd45153, 16'd22103, 16'd37113, 16'd37703, 16'd63032, 16'd17661, 16'd46310, 16'd32004, 16'd20330, 16'd36231, 16'd61354, 16'd19241, 16'd30635, 16'd59893, 16'd2155, 16'd35028, 16'd24563, 16'd46348});
	test_expansion(128'h6a327043d66eb42a79b313d80636cc81, {16'd2007, 16'd27044, 16'd57358, 16'd37067, 16'd29883, 16'd5620, 16'd3205, 16'd19935, 16'd14068, 16'd58558, 16'd45376, 16'd35194, 16'd17485, 16'd49967, 16'd28093, 16'd16784, 16'd53493, 16'd20238, 16'd58207, 16'd3012, 16'd35976, 16'd65131, 16'd56891, 16'd21349, 16'd47106, 16'd20061});
	test_expansion(128'h8b5d0b8dad1acac6a7e8dbcf8d17a317, {16'd30463, 16'd63455, 16'd13455, 16'd42305, 16'd36957, 16'd21832, 16'd47864, 16'd8453, 16'd30335, 16'd50617, 16'd57929, 16'd30029, 16'd6953, 16'd17549, 16'd44186, 16'd63449, 16'd25886, 16'd23634, 16'd8240, 16'd27339, 16'd19607, 16'd41227, 16'd45109, 16'd2528, 16'd19095, 16'd41742});
	test_expansion(128'h80bcf29e3a15e860e17bed8a7f9fb1a5, {16'd45765, 16'd13028, 16'd38137, 16'd29157, 16'd63157, 16'd25839, 16'd40474, 16'd10314, 16'd38560, 16'd20594, 16'd9111, 16'd19605, 16'd20700, 16'd53679, 16'd44148, 16'd58904, 16'd6156, 16'd17492, 16'd46187, 16'd13953, 16'd53089, 16'd10342, 16'd21216, 16'd27339, 16'd57697, 16'd9129});
	test_expansion(128'haa8d2ada9402efddfca9d71e74a9d1c2, {16'd44014, 16'd58480, 16'd53199, 16'd50899, 16'd14022, 16'd322, 16'd36232, 16'd63714, 16'd8510, 16'd61468, 16'd13163, 16'd56296, 16'd23886, 16'd50186, 16'd27583, 16'd54514, 16'd15205, 16'd35181, 16'd26160, 16'd8366, 16'd1980, 16'd47482, 16'd40074, 16'd54178, 16'd5143, 16'd46480});
	test_expansion(128'h70a752cbfc8b05027a8d2bce07a40416, {16'd30002, 16'd13764, 16'd21034, 16'd61988, 16'd39369, 16'd37702, 16'd57224, 16'd32707, 16'd12520, 16'd2435, 16'd57345, 16'd21337, 16'd32643, 16'd47995, 16'd30040, 16'd45440, 16'd4132, 16'd33280, 16'd59917, 16'd63280, 16'd26671, 16'd3612, 16'd65493, 16'd15931, 16'd12881, 16'd58819});
	test_expansion(128'h882db8dc7604f92419b4911d9309ecfe, {16'd14531, 16'd5119, 16'd51457, 16'd29193, 16'd12833, 16'd56408, 16'd62442, 16'd10054, 16'd33804, 16'd3132, 16'd9149, 16'd23407, 16'd8402, 16'd3076, 16'd61736, 16'd34033, 16'd54373, 16'd11055, 16'd63005, 16'd64739, 16'd43188, 16'd13993, 16'd54779, 16'd44921, 16'd8235, 16'd20200});
	test_expansion(128'h30229518db921e05d3ae2877b570486d, {16'd48304, 16'd12860, 16'd17389, 16'd24462, 16'd51062, 16'd35580, 16'd46778, 16'd8521, 16'd33013, 16'd53068, 16'd16139, 16'd8344, 16'd40319, 16'd18251, 16'd8323, 16'd59399, 16'd63518, 16'd49970, 16'd5184, 16'd38490, 16'd54232, 16'd17056, 16'd36870, 16'd25974, 16'd30660, 16'd27044});
	test_expansion(128'h6ba0f1022e98efd00d5d993e47b5506e, {16'd33856, 16'd25189, 16'd6631, 16'd50424, 16'd53299, 16'd3617, 16'd65337, 16'd16395, 16'd10276, 16'd15014, 16'd8304, 16'd27828, 16'd33145, 16'd17723, 16'd40388, 16'd37606, 16'd15457, 16'd8456, 16'd41575, 16'd63340, 16'd61092, 16'd39673, 16'd45734, 16'd30919, 16'd48437, 16'd29098});
	test_expansion(128'hfecdc2399d2a1a4a283a78fbf1fb651a, {16'd24529, 16'd3404, 16'd32176, 16'd38442, 16'd39589, 16'd33334, 16'd7503, 16'd37624, 16'd59077, 16'd51353, 16'd39478, 16'd14935, 16'd46310, 16'd38145, 16'd60842, 16'd5416, 16'd56329, 16'd27173, 16'd47385, 16'd43109, 16'd51445, 16'd62935, 16'd9160, 16'd2511, 16'd10280, 16'd29192});
	test_expansion(128'ha78c2aa56e33b8dd51a7f357078c510f, {16'd25423, 16'd30638, 16'd50628, 16'd19010, 16'd39066, 16'd41269, 16'd7515, 16'd51122, 16'd15992, 16'd59677, 16'd21900, 16'd33068, 16'd27156, 16'd49701, 16'd32421, 16'd35487, 16'd22360, 16'd16692, 16'd52303, 16'd63952, 16'd25353, 16'd55589, 16'd29306, 16'd26934, 16'd27705, 16'd21395});
	test_expansion(128'h2f2f3d3a21e27e6c3cb8c17f13981905, {16'd53490, 16'd54911, 16'd2476, 16'd9199, 16'd60681, 16'd36702, 16'd13236, 16'd40255, 16'd7063, 16'd15398, 16'd25874, 16'd3320, 16'd33330, 16'd40306, 16'd21124, 16'd53464, 16'd13819, 16'd63865, 16'd48470, 16'd59472, 16'd13269, 16'd14575, 16'd50565, 16'd36390, 16'd49928, 16'd10751});
	test_expansion(128'hbeb3383c6af95d1f2cac0ceff70c936d, {16'd13313, 16'd47940, 16'd38447, 16'd51680, 16'd33432, 16'd7375, 16'd64163, 16'd58886, 16'd57235, 16'd16555, 16'd17307, 16'd51778, 16'd39231, 16'd10418, 16'd9549, 16'd27973, 16'd16298, 16'd30576, 16'd7085, 16'd61386, 16'd63553, 16'd14227, 16'd9755, 16'd56492, 16'd27777, 16'd50167});
	test_expansion(128'h171b9f37c8ba33184ddd457d7acd591a, {16'd30220, 16'd5891, 16'd7885, 16'd22246, 16'd12876, 16'd28388, 16'd65033, 16'd11428, 16'd36103, 16'd57632, 16'd58627, 16'd5832, 16'd50302, 16'd27044, 16'd45543, 16'd9625, 16'd9398, 16'd57298, 16'd37678, 16'd17889, 16'd20857, 16'd11556, 16'd64526, 16'd58874, 16'd12108, 16'd40639});
	test_expansion(128'h666a7abb61f7856069a41f0dee39134d, {16'd31691, 16'd58721, 16'd21139, 16'd7477, 16'd25368, 16'd57056, 16'd44402, 16'd10537, 16'd52505, 16'd52182, 16'd4744, 16'd4053, 16'd53159, 16'd25557, 16'd8283, 16'd14258, 16'd56949, 16'd457, 16'd3094, 16'd63035, 16'd43549, 16'd43407, 16'd48797, 16'd26523, 16'd10922, 16'd5586});
	test_expansion(128'h2d01874b1bea5c49e415d9fb5ba9fcb7, {16'd9944, 16'd62303, 16'd2638, 16'd26586, 16'd34679, 16'd500, 16'd34974, 16'd39959, 16'd16541, 16'd17521, 16'd42591, 16'd47666, 16'd37746, 16'd29797, 16'd49009, 16'd10532, 16'd7082, 16'd20429, 16'd57634, 16'd9851, 16'd42145, 16'd46237, 16'd8546, 16'd36888, 16'd6329, 16'd3433});
	test_expansion(128'hb920e711a59706865187afd4981ae373, {16'd40846, 16'd18691, 16'd47530, 16'd10801, 16'd64111, 16'd37947, 16'd62709, 16'd18456, 16'd53781, 16'd30366, 16'd8060, 16'd8168, 16'd10619, 16'd3984, 16'd28747, 16'd46773, 16'd38799, 16'd11488, 16'd36809, 16'd1316, 16'd20201, 16'd54130, 16'd48503, 16'd9774, 16'd8813, 16'd52354});
	test_expansion(128'h0a500f120ecf2fde411a87b2ce8dda7b, {16'd43305, 16'd44568, 16'd42880, 16'd29672, 16'd16878, 16'd47411, 16'd10676, 16'd45582, 16'd35765, 16'd52310, 16'd24123, 16'd26952, 16'd11066, 16'd40577, 16'd26631, 16'd58133, 16'd12291, 16'd39239, 16'd55464, 16'd57953, 16'd1504, 16'd9052, 16'd17414, 16'd11325, 16'd11035, 16'd3275});
	test_expansion(128'hbb4a66ef4845efde04337d457344459d, {16'd26397, 16'd54031, 16'd32818, 16'd33842, 16'd18522, 16'd48174, 16'd23234, 16'd14250, 16'd62024, 16'd44819, 16'd5012, 16'd1601, 16'd47089, 16'd56061, 16'd62061, 16'd55419, 16'd23051, 16'd49378, 16'd63637, 16'd9746, 16'd47619, 16'd44650, 16'd46481, 16'd55249, 16'd47055, 16'd26553});
	test_expansion(128'h4889b33f4471fc49126567931b97cd8d, {16'd63083, 16'd28815, 16'd1009, 16'd39107, 16'd32029, 16'd40978, 16'd44706, 16'd19846, 16'd25379, 16'd32313, 16'd45196, 16'd41697, 16'd6445, 16'd41540, 16'd8149, 16'd28780, 16'd32638, 16'd56383, 16'd12667, 16'd51959, 16'd19718, 16'd11991, 16'd1761, 16'd9171, 16'd44169, 16'd47235});
	test_expansion(128'haf40ca7763f8e1a1d8426aed6e66d9a6, {16'd30166, 16'd57234, 16'd20873, 16'd25134, 16'd30824, 16'd56201, 16'd648, 16'd38559, 16'd55452, 16'd30690, 16'd54788, 16'd1389, 16'd33945, 16'd13244, 16'd22787, 16'd46074, 16'd3191, 16'd46568, 16'd12760, 16'd49761, 16'd63375, 16'd29596, 16'd48614, 16'd2352, 16'd62206, 16'd5515});
	test_expansion(128'h253bc0afe82d678ed4fce8e00bc28797, {16'd5346, 16'd38997, 16'd14486, 16'd58073, 16'd24940, 16'd58743, 16'd55867, 16'd5022, 16'd20021, 16'd55730, 16'd20158, 16'd3995, 16'd43584, 16'd56885, 16'd18101, 16'd30688, 16'd2153, 16'd24338, 16'd22648, 16'd7950, 16'd52757, 16'd48170, 16'd40543, 16'd52906, 16'd59200, 16'd48973});
	test_expansion(128'he53b3fad49c16d86093e27a50b92277e, {16'd61545, 16'd57543, 16'd37504, 16'd20348, 16'd34251, 16'd8559, 16'd55275, 16'd15957, 16'd52123, 16'd29519, 16'd15430, 16'd27349, 16'd62572, 16'd57586, 16'd6166, 16'd26252, 16'd11745, 16'd62956, 16'd5725, 16'd64562, 16'd34955, 16'd19812, 16'd2117, 16'd35014, 16'd34133, 16'd52730});
	test_expansion(128'ha3af46b291683339a27dfd8f6a74053e, {16'd1562, 16'd47636, 16'd53574, 16'd26105, 16'd35601, 16'd29472, 16'd55868, 16'd43016, 16'd21739, 16'd58470, 16'd32075, 16'd62840, 16'd52617, 16'd43694, 16'd17754, 16'd37247, 16'd16287, 16'd62090, 16'd33160, 16'd27486, 16'd2678, 16'd15070, 16'd5743, 16'd37136, 16'd50181, 16'd53603});
	test_expansion(128'h84f5f77874907de9c1404effd4b1b592, {16'd41864, 16'd34949, 16'd23319, 16'd56939, 16'd37494, 16'd64030, 16'd29698, 16'd39878, 16'd52792, 16'd4484, 16'd64643, 16'd1987, 16'd20424, 16'd37729, 16'd6120, 16'd51792, 16'd61267, 16'd29907, 16'd60774, 16'd59059, 16'd40022, 16'd17235, 16'd50881, 16'd62266, 16'd28654, 16'd6928});
	test_expansion(128'h484d65041097283ade5131daba0502f3, {16'd34967, 16'd349, 16'd24206, 16'd7026, 16'd48271, 16'd2460, 16'd17249, 16'd4016, 16'd44558, 16'd21052, 16'd40389, 16'd48742, 16'd40037, 16'd13095, 16'd64176, 16'd62669, 16'd63472, 16'd39338, 16'd55740, 16'd29952, 16'd39178, 16'd41842, 16'd44716, 16'd31033, 16'd43756, 16'd46069});
	test_expansion(128'hbd747bc6af51072a0a14741131a18ac5, {16'd12902, 16'd52831, 16'd54619, 16'd31374, 16'd22224, 16'd50741, 16'd35000, 16'd8099, 16'd22228, 16'd44317, 16'd43744, 16'd3526, 16'd62972, 16'd62465, 16'd33956, 16'd24681, 16'd13179, 16'd19314, 16'd33392, 16'd37465, 16'd38564, 16'd47832, 16'd49005, 16'd28036, 16'd55731, 16'd4070});
	test_expansion(128'h28a2b137a6286fe9c8e92cd4d29d4f42, {16'd31040, 16'd59089, 16'd24276, 16'd31768, 16'd33340, 16'd43301, 16'd23466, 16'd43874, 16'd46310, 16'd62837, 16'd40170, 16'd32063, 16'd36943, 16'd19353, 16'd28055, 16'd57112, 16'd58190, 16'd31359, 16'd59644, 16'd38848, 16'd50845, 16'd3678, 16'd63985, 16'd33930, 16'd2537, 16'd33455});
	test_expansion(128'ha08a7eaa7c30e90ea3811a92e4070bd9, {16'd12449, 16'd61854, 16'd16129, 16'd42969, 16'd42787, 16'd36181, 16'd39659, 16'd16821, 16'd27424, 16'd8014, 16'd24777, 16'd9421, 16'd405, 16'd142, 16'd46842, 16'd18624, 16'd23085, 16'd46069, 16'd43866, 16'd45698, 16'd32039, 16'd12594, 16'd60046, 16'd6215, 16'd44513, 16'd20908});
	test_expansion(128'h2e9a453f3f249bb8104efa0bc8a3289a, {16'd45702, 16'd12914, 16'd36921, 16'd63038, 16'd7205, 16'd5205, 16'd47355, 16'd51530, 16'd26466, 16'd39140, 16'd37654, 16'd54995, 16'd56430, 16'd14210, 16'd64384, 16'd31894, 16'd42789, 16'd52498, 16'd30539, 16'd18040, 16'd45019, 16'd50984, 16'd24525, 16'd42040, 16'd57607, 16'd51712});
	test_expansion(128'hecd8caeb408c1d64c388bb135de64c9e, {16'd64268, 16'd40469, 16'd31165, 16'd22727, 16'd64843, 16'd28481, 16'd11236, 16'd45330, 16'd53589, 16'd26641, 16'd38185, 16'd15869, 16'd13661, 16'd23321, 16'd6392, 16'd22661, 16'd60329, 16'd30864, 16'd55874, 16'd39959, 16'd41935, 16'd12895, 16'd52848, 16'd21124, 16'd2004, 16'd1420});
	test_expansion(128'he794e32773d60e94b96310a9670af413, {16'd28459, 16'd6358, 16'd49828, 16'd4838, 16'd37770, 16'd63186, 16'd49377, 16'd8883, 16'd58252, 16'd49431, 16'd12121, 16'd39511, 16'd20474, 16'd41271, 16'd29083, 16'd50603, 16'd38560, 16'd23359, 16'd42268, 16'd42970, 16'd4671, 16'd27234, 16'd35533, 16'd14421, 16'd35707, 16'd18772});
	test_expansion(128'ha74f3a8cbfecad6af11775e43c2893af, {16'd55009, 16'd11862, 16'd60276, 16'd12613, 16'd57573, 16'd17987, 16'd53669, 16'd15592, 16'd35945, 16'd60087, 16'd32735, 16'd7367, 16'd3351, 16'd16986, 16'd39972, 16'd49, 16'd34856, 16'd19990, 16'd55673, 16'd5296, 16'd38107, 16'd19946, 16'd11908, 16'd65377, 16'd25786, 16'd4127});
	test_expansion(128'h19929ba212a08920dfc98831c0ccecde, {16'd6002, 16'd58156, 16'd18430, 16'd56589, 16'd32225, 16'd46165, 16'd8437, 16'd42537, 16'd5671, 16'd40932, 16'd8819, 16'd57470, 16'd26685, 16'd30114, 16'd46837, 16'd45645, 16'd52306, 16'd38842, 16'd25236, 16'd3218, 16'd14156, 16'd15795, 16'd28527, 16'd37963, 16'd22960, 16'd33780});
	test_expansion(128'h86c2a9d628f5d923cc9b99c6c9082fb7, {16'd15565, 16'd29011, 16'd42178, 16'd17419, 16'd15139, 16'd41545, 16'd39282, 16'd19998, 16'd46968, 16'd10878, 16'd32434, 16'd43766, 16'd44565, 16'd1034, 16'd53986, 16'd20950, 16'd64851, 16'd30353, 16'd36562, 16'd14523, 16'd18, 16'd15742, 16'd16320, 16'd19395, 16'd44938, 16'd12034});
	test_expansion(128'h86288a7332eeb00e53891f084145287e, {16'd54918, 16'd12564, 16'd51937, 16'd63267, 16'd27070, 16'd62591, 16'd53562, 16'd32849, 16'd23066, 16'd21345, 16'd55291, 16'd64637, 16'd50436, 16'd62934, 16'd10280, 16'd8971, 16'd36728, 16'd20872, 16'd26455, 16'd39823, 16'd4799, 16'd52266, 16'd23768, 16'd7577, 16'd45175, 16'd31673});
	test_expansion(128'hdd93dacd74c46465de7a2e9ab7cee044, {16'd9031, 16'd18063, 16'd33772, 16'd55236, 16'd2449, 16'd13338, 16'd53970, 16'd22524, 16'd45765, 16'd41575, 16'd59143, 16'd54171, 16'd17591, 16'd64431, 16'd20549, 16'd17217, 16'd34324, 16'd5695, 16'd7778, 16'd15613, 16'd42254, 16'd48487, 16'd28253, 16'd51001, 16'd48386, 16'd20308});
	test_expansion(128'h0a194ca955a29c61abdd99a9b55151f3, {16'd18585, 16'd27408, 16'd30222, 16'd25928, 16'd61436, 16'd362, 16'd60277, 16'd7688, 16'd53682, 16'd36100, 16'd44180, 16'd8098, 16'd48372, 16'd4364, 16'd45645, 16'd22777, 16'd61947, 16'd55946, 16'd56049, 16'd47455, 16'd22504, 16'd47903, 16'd10746, 16'd36316, 16'd24122, 16'd5977});
	test_expansion(128'h018d5c9a6eff9846a39de4e3c4b5b403, {16'd54518, 16'd39225, 16'd41916, 16'd32131, 16'd24459, 16'd57439, 16'd22833, 16'd22926, 16'd40150, 16'd52557, 16'd31607, 16'd43760, 16'd7832, 16'd65384, 16'd25351, 16'd63368, 16'd58718, 16'd10967, 16'd9523, 16'd48176, 16'd39056, 16'd50857, 16'd47426, 16'd21469, 16'd7850, 16'd50522});
	test_expansion(128'hbe3c700fdf515146a060d7fbe8ba00ff, {16'd49852, 16'd47702, 16'd46822, 16'd43052, 16'd47157, 16'd3011, 16'd37686, 16'd36895, 16'd24615, 16'd30491, 16'd1873, 16'd24789, 16'd34715, 16'd53893, 16'd61849, 16'd27954, 16'd4689, 16'd18298, 16'd43177, 16'd19559, 16'd12459, 16'd28809, 16'd52517, 16'd26191, 16'd56869, 16'd309});
	test_expansion(128'h59a865920fbd21259187a91e5438cf8b, {16'd15568, 16'd46346, 16'd16673, 16'd7874, 16'd28543, 16'd63694, 16'd37527, 16'd15889, 16'd3024, 16'd42479, 16'd62069, 16'd931, 16'd7318, 16'd55582, 16'd25305, 16'd32719, 16'd13503, 16'd898, 16'd7587, 16'd36195, 16'd22994, 16'd10845, 16'd21493, 16'd11899, 16'd55840, 16'd34456});
	test_expansion(128'h06b1b95722ca4e953d0c519de93eecf1, {16'd13580, 16'd34804, 16'd15680, 16'd22483, 16'd19690, 16'd10062, 16'd53101, 16'd7814, 16'd5862, 16'd22910, 16'd36741, 16'd56010, 16'd47314, 16'd13005, 16'd41165, 16'd43644, 16'd6817, 16'd20349, 16'd63369, 16'd37943, 16'd10095, 16'd43487, 16'd45575, 16'd33663, 16'd32442, 16'd3195});
	test_expansion(128'h2432690a2ccbec0de65fdd5c855ee7a7, {16'd10107, 16'd50162, 16'd29394, 16'd12455, 16'd10363, 16'd3693, 16'd60900, 16'd55900, 16'd4544, 16'd26860, 16'd27403, 16'd10662, 16'd21002, 16'd48497, 16'd40094, 16'd50600, 16'd48992, 16'd12644, 16'd29099, 16'd7692, 16'd44143, 16'd30565, 16'd44577, 16'd51275, 16'd64212, 16'd11867});
	test_expansion(128'h0eaa4ca51b2557ddf56221b4cbf73984, {16'd25640, 16'd14957, 16'd23488, 16'd14327, 16'd47070, 16'd8781, 16'd62586, 16'd7559, 16'd60186, 16'd64088, 16'd16900, 16'd35939, 16'd26620, 16'd20618, 16'd40193, 16'd64819, 16'd60246, 16'd11589, 16'd35538, 16'd31076, 16'd32031, 16'd34482, 16'd26100, 16'd26517, 16'd17454, 16'd62321});
	test_expansion(128'hab4a3c366f1e1a23049bc0f69c8a1d69, {16'd49409, 16'd43243, 16'd31199, 16'd63207, 16'd57031, 16'd25603, 16'd21961, 16'd16871, 16'd15430, 16'd27000, 16'd43386, 16'd44797, 16'd26270, 16'd1910, 16'd25877, 16'd36798, 16'd25076, 16'd10243, 16'd29612, 16'd14413, 16'd50997, 16'd36737, 16'd58028, 16'd22883, 16'd52579, 16'd3523});
	test_expansion(128'h05bb699ea781086d041f2ecc85b59a10, {16'd19233, 16'd41913, 16'd44152, 16'd9806, 16'd18883, 16'd39122, 16'd18754, 16'd21732, 16'd25629, 16'd7306, 16'd6964, 16'd31373, 16'd56756, 16'd62456, 16'd60449, 16'd65120, 16'd65126, 16'd2231, 16'd48470, 16'd19159, 16'd387, 16'd11375, 16'd27695, 16'd6966, 16'd20572, 16'd39771});
	test_expansion(128'h8cd288c2de69c8538b34152ebb3c909b, {16'd60805, 16'd27299, 16'd39535, 16'd48238, 16'd25096, 16'd30085, 16'd46810, 16'd8352, 16'd64328, 16'd46305, 16'd42107, 16'd18462, 16'd61357, 16'd39339, 16'd57014, 16'd17479, 16'd1498, 16'd30735, 16'd44892, 16'd37723, 16'd40088, 16'd11204, 16'd12691, 16'd58238, 16'd65148, 16'd14264});
	test_expansion(128'h7a4f75144f91f3de08234e0240d53c56, {16'd16357, 16'd10545, 16'd52168, 16'd23306, 16'd3436, 16'd34002, 16'd50596, 16'd1312, 16'd38935, 16'd12475, 16'd9911, 16'd15659, 16'd9078, 16'd62296, 16'd49142, 16'd18108, 16'd63481, 16'd20792, 16'd4384, 16'd32199, 16'd42197, 16'd653, 16'd64420, 16'd52949, 16'd26845, 16'd27739});
	test_expansion(128'hc515d4025024a71dd9858106b7c3ebd9, {16'd31840, 16'd10073, 16'd24282, 16'd63930, 16'd25809, 16'd9284, 16'd8156, 16'd6720, 16'd57355, 16'd55238, 16'd39474, 16'd9721, 16'd52537, 16'd42428, 16'd42519, 16'd2750, 16'd56531, 16'd3362, 16'd6674, 16'd42098, 16'd19022, 16'd3844, 16'd14863, 16'd42513, 16'd24439, 16'd37376});
	test_expansion(128'he23c00d06efe72bced6508fde16e4899, {16'd38084, 16'd58324, 16'd19126, 16'd27840, 16'd49046, 16'd24424, 16'd42493, 16'd23626, 16'd36997, 16'd13413, 16'd45106, 16'd29868, 16'd20576, 16'd29501, 16'd60062, 16'd52257, 16'd63906, 16'd40904, 16'd37624, 16'd47196, 16'd58680, 16'd62322, 16'd38266, 16'd4624, 16'd62533, 16'd31764});
	test_expansion(128'h7ead2e330c237f5dbe080f2e52eac613, {16'd4831, 16'd5934, 16'd52699, 16'd59369, 16'd22316, 16'd22907, 16'd63547, 16'd30225, 16'd49834, 16'd41966, 16'd32367, 16'd62368, 16'd41334, 16'd19093, 16'd4686, 16'd5766, 16'd39253, 16'd60251, 16'd27808, 16'd17589, 16'd10355, 16'd27107, 16'd50995, 16'd37858, 16'd33392, 16'd33481});
	test_expansion(128'hf36aa7a3303d7e9ed5bd1bab940dcb2f, {16'd35668, 16'd10775, 16'd56450, 16'd19351, 16'd1565, 16'd58953, 16'd37650, 16'd43719, 16'd13213, 16'd14268, 16'd42325, 16'd51592, 16'd32287, 16'd18326, 16'd61828, 16'd63566, 16'd10019, 16'd37404, 16'd23183, 16'd39018, 16'd16969, 16'd50796, 16'd8197, 16'd35481, 16'd56320, 16'd44229});
	test_expansion(128'he8b0af64cc9adb0d5d129fa7a3d1aa15, {16'd49061, 16'd15314, 16'd57073, 16'd35875, 16'd57562, 16'd38639, 16'd37775, 16'd59739, 16'd3512, 16'd6036, 16'd33623, 16'd33795, 16'd62716, 16'd655, 16'd62747, 16'd37555, 16'd7214, 16'd11981, 16'd4267, 16'd58014, 16'd46640, 16'd29595, 16'd34266, 16'd25619, 16'd11535, 16'd3367});
	test_expansion(128'h457412225b82794f2abd6cb6ab11d53a, {16'd61459, 16'd39838, 16'd8844, 16'd26129, 16'd57476, 16'd11835, 16'd29186, 16'd23168, 16'd12217, 16'd61989, 16'd30153, 16'd53327, 16'd13133, 16'd18032, 16'd56296, 16'd36343, 16'd62439, 16'd39021, 16'd37439, 16'd30293, 16'd19128, 16'd264, 16'd59249, 16'd17650, 16'd28968, 16'd30357});
	test_expansion(128'h756b43be2ffa26f7debe49740f2c9b70, {16'd10687, 16'd23972, 16'd54586, 16'd22123, 16'd24310, 16'd35818, 16'd20016, 16'd20350, 16'd8881, 16'd46412, 16'd63481, 16'd29158, 16'd26890, 16'd46551, 16'd22235, 16'd37190, 16'd61867, 16'd12037, 16'd15510, 16'd53332, 16'd41209, 16'd41987, 16'd36130, 16'd34509, 16'd34946, 16'd16053});
	test_expansion(128'hf29e9a0050a19a108f7ea87a849648fb, {16'd7997, 16'd39432, 16'd6027, 16'd56045, 16'd19440, 16'd55834, 16'd34978, 16'd34150, 16'd59934, 16'd5538, 16'd2212, 16'd56806, 16'd24588, 16'd29189, 16'd54573, 16'd28052, 16'd44647, 16'd31035, 16'd40597, 16'd26689, 16'd35560, 16'd58928, 16'd4689, 16'd15489, 16'd29258, 16'd53978});
	test_expansion(128'hc514cf2d30052f92184125a5d98dbb70, {16'd42406, 16'd2154, 16'd28130, 16'd19986, 16'd32288, 16'd44849, 16'd42317, 16'd15395, 16'd32559, 16'd13997, 16'd6790, 16'd44694, 16'd17680, 16'd41723, 16'd18598, 16'd4894, 16'd56982, 16'd983, 16'd63977, 16'd197, 16'd22299, 16'd38927, 16'd29060, 16'd35390, 16'd47158, 16'd53819});
	test_expansion(128'ha4c5e3f7bf7785956c49813072178be3, {16'd38718, 16'd6824, 16'd14626, 16'd14531, 16'd25912, 16'd46105, 16'd37112, 16'd53931, 16'd29682, 16'd26921, 16'd20735, 16'd7732, 16'd35160, 16'd3721, 16'd18860, 16'd24354, 16'd18380, 16'd31591, 16'd57689, 16'd43072, 16'd47179, 16'd23769, 16'd12855, 16'd18475, 16'd13364, 16'd58606});
	test_expansion(128'h405f16e5bc491fab754ca4ec9342d4a4, {16'd21371, 16'd61537, 16'd6285, 16'd32141, 16'd22767, 16'd42427, 16'd18926, 16'd15727, 16'd11334, 16'd33187, 16'd34137, 16'd60780, 16'd12943, 16'd58290, 16'd33979, 16'd45237, 16'd56434, 16'd26712, 16'd52389, 16'd18463, 16'd31810, 16'd52258, 16'd46274, 16'd40982, 16'd25050, 16'd5252});
	test_expansion(128'hac8e40722dc418d63b6cfe985a0e0def, {16'd63558, 16'd29513, 16'd29422, 16'd7950, 16'd29463, 16'd12879, 16'd65489, 16'd64912, 16'd53571, 16'd29743, 16'd7094, 16'd61141, 16'd44127, 16'd47253, 16'd32374, 16'd5023, 16'd20148, 16'd11775, 16'd47242, 16'd45094, 16'd22131, 16'd30433, 16'd36650, 16'd7639, 16'd21316, 16'd24810});
	test_expansion(128'h939cb12942b2624e5f9635f9123c541b, {16'd53484, 16'd34881, 16'd23121, 16'd22945, 16'd38736, 16'd26884, 16'd31185, 16'd39408, 16'd59323, 16'd26143, 16'd39723, 16'd37808, 16'd165, 16'd11119, 16'd14821, 16'd53247, 16'd14320, 16'd62882, 16'd26907, 16'd56705, 16'd25450, 16'd10220, 16'd35820, 16'd47526, 16'd1184, 16'd57707});
	test_expansion(128'h33104e14f3932237624505fc04e97b3d, {16'd43398, 16'd34422, 16'd56868, 16'd22506, 16'd18448, 16'd22902, 16'd5876, 16'd49124, 16'd24945, 16'd41159, 16'd58359, 16'd38728, 16'd2654, 16'd20903, 16'd58624, 16'd52440, 16'd54755, 16'd65456, 16'd11334, 16'd32389, 16'd13404, 16'd8837, 16'd40287, 16'd36824, 16'd43658, 16'd65236});
	test_expansion(128'h5860f379fa5fa908d5869c8ad2b66740, {16'd57498, 16'd28008, 16'd9398, 16'd37391, 16'd21895, 16'd3234, 16'd30855, 16'd51511, 16'd63939, 16'd62387, 16'd22269, 16'd23051, 16'd42524, 16'd44431, 16'd48177, 16'd36607, 16'd1485, 16'd37566, 16'd30708, 16'd31254, 16'd30882, 16'd51387, 16'd24899, 16'd24862, 16'd13464, 16'd25144});
	test_expansion(128'h025b3de007d0a7ee6ae95d189e2fec0c, {16'd59661, 16'd56096, 16'd10563, 16'd63909, 16'd63296, 16'd16864, 16'd56242, 16'd35411, 16'd49352, 16'd28394, 16'd21187, 16'd64289, 16'd1835, 16'd52800, 16'd49439, 16'd63358, 16'd10099, 16'd57406, 16'd45060, 16'd46719, 16'd30380, 16'd21894, 16'd5158, 16'd20527, 16'd11217, 16'd16711});
	test_expansion(128'h99e84fcd15eceefedffbdca5e5cd5196, {16'd25397, 16'd5257, 16'd623, 16'd39757, 16'd21063, 16'd23127, 16'd54898, 16'd96, 16'd20372, 16'd1996, 16'd4154, 16'd14439, 16'd19626, 16'd7945, 16'd4012, 16'd47140, 16'd52343, 16'd23491, 16'd10597, 16'd44517, 16'd4326, 16'd24825, 16'd65023, 16'd58489, 16'd3094, 16'd5315});
	test_expansion(128'h5d6aef772651d8fd2948950d13408b14, {16'd3569, 16'd25745, 16'd60625, 16'd40046, 16'd46852, 16'd26850, 16'd46976, 16'd56290, 16'd38864, 16'd26045, 16'd42655, 16'd45017, 16'd43572, 16'd63895, 16'd7239, 16'd52241, 16'd61598, 16'd19725, 16'd20157, 16'd34650, 16'd25583, 16'd32840, 16'd50173, 16'd37023, 16'd12908, 16'd2372});
	test_expansion(128'h565072b3d20cdf4c037ca0957f71cea3, {16'd33101, 16'd259, 16'd1312, 16'd23635, 16'd42274, 16'd43144, 16'd15837, 16'd17579, 16'd677, 16'd52358, 16'd10826, 16'd3921, 16'd46952, 16'd13026, 16'd48053, 16'd28191, 16'd62259, 16'd7094, 16'd11427, 16'd12495, 16'd31753, 16'd3512, 16'd29321, 16'd52444, 16'd101, 16'd50641});
	test_expansion(128'hae20b3c655f666643f5cbecb5ed6ebc2, {16'd35475, 16'd40914, 16'd64548, 16'd46366, 16'd49723, 16'd31746, 16'd41783, 16'd59047, 16'd16419, 16'd58190, 16'd40032, 16'd6542, 16'd5820, 16'd15834, 16'd23679, 16'd42248, 16'd16675, 16'd39867, 16'd6602, 16'd51440, 16'd40275, 16'd2255, 16'd33352, 16'd56779, 16'd30532, 16'd32594});
	test_expansion(128'hcaa97b5818af87b5bb6be15f713d86a7, {16'd32638, 16'd15173, 16'd180, 16'd33146, 16'd47503, 16'd43405, 16'd9475, 16'd35008, 16'd25777, 16'd45044, 16'd52878, 16'd16917, 16'd50959, 16'd29713, 16'd28348, 16'd18399, 16'd27631, 16'd7224, 16'd16772, 16'd9294, 16'd59838, 16'd12696, 16'd42396, 16'd64289, 16'd35038, 16'd29334});
	test_expansion(128'h86542418a78e3050429b1238fddf0db5, {16'd52166, 16'd58431, 16'd20017, 16'd32077, 16'd23245, 16'd53367, 16'd34446, 16'd42063, 16'd33692, 16'd8593, 16'd3050, 16'd26393, 16'd6892, 16'd51824, 16'd57669, 16'd12265, 16'd21855, 16'd33955, 16'd10841, 16'd9255, 16'd20216, 16'd8227, 16'd10210, 16'd54532, 16'd29572, 16'd31549});
	test_expansion(128'he8ec7a77f9ecbf703d3b83d36513e8d1, {16'd27979, 16'd58015, 16'd14412, 16'd48208, 16'd23183, 16'd37027, 16'd57104, 16'd64753, 16'd55865, 16'd52542, 16'd4741, 16'd7117, 16'd41564, 16'd16702, 16'd55478, 16'd297, 16'd23850, 16'd31958, 16'd46134, 16'd610, 16'd51, 16'd9951, 16'd40833, 16'd64115, 16'd33412, 16'd62419});
	test_expansion(128'hfa622bbe470f5ffa6b9c915fbbf18b36, {16'd20664, 16'd20154, 16'd47093, 16'd30014, 16'd10445, 16'd13179, 16'd33812, 16'd62680, 16'd13207, 16'd64580, 16'd41260, 16'd23256, 16'd43564, 16'd6805, 16'd28124, 16'd34598, 16'd2570, 16'd13697, 16'd62479, 16'd5913, 16'd15804, 16'd64799, 16'd38209, 16'd29300, 16'd35923, 16'd48605});
	test_expansion(128'hf7c3c8f8371ad584160fe94f26e07c6b, {16'd6973, 16'd37353, 16'd18138, 16'd48068, 16'd47579, 16'd37010, 16'd23740, 16'd18911, 16'd9007, 16'd54862, 16'd59872, 16'd8507, 16'd25224, 16'd56297, 16'd41084, 16'd4427, 16'd42233, 16'd64521, 16'd2482, 16'd8445, 16'd32481, 16'd6465, 16'd23049, 16'd50866, 16'd64376, 16'd53843});
	test_expansion(128'hb7395ae2028e569b23504b109178ea9d, {16'd50793, 16'd50199, 16'd62670, 16'd15056, 16'd49260, 16'd21710, 16'd8874, 16'd34274, 16'd16846, 16'd20724, 16'd13481, 16'd52452, 16'd46438, 16'd39909, 16'd26697, 16'd56186, 16'd8129, 16'd65172, 16'd33096, 16'd28679, 16'd15094, 16'd19863, 16'd10268, 16'd32299, 16'd40711, 16'd5503});
	test_expansion(128'h7afe837843baa87ff5637f8e76c5b7db, {16'd59462, 16'd23815, 16'd20934, 16'd35703, 16'd3915, 16'd17034, 16'd43599, 16'd39338, 16'd37383, 16'd2877, 16'd16918, 16'd35236, 16'd22300, 16'd42487, 16'd16577, 16'd18884, 16'd7977, 16'd53780, 16'd25450, 16'd64957, 16'd982, 16'd37230, 16'd32309, 16'd39610, 16'd13798, 16'd41864});
	test_expansion(128'h50bb3eebeab11c3145d6447a2572db4e, {16'd34437, 16'd35865, 16'd11072, 16'd13462, 16'd64800, 16'd45159, 16'd9325, 16'd25987, 16'd37662, 16'd22350, 16'd61828, 16'd4309, 16'd34006, 16'd25039, 16'd3816, 16'd57981, 16'd21852, 16'd14012, 16'd61616, 16'd44051, 16'd53058, 16'd55043, 16'd9655, 16'd28157, 16'd26992, 16'd47148});
	test_expansion(128'hf7b6af87abc454c4445b205e854baf91, {16'd39925, 16'd26676, 16'd31011, 16'd59704, 16'd27903, 16'd41324, 16'd36314, 16'd52876, 16'd43452, 16'd30187, 16'd19520, 16'd52681, 16'd5172, 16'd23874, 16'd28349, 16'd24597, 16'd45020, 16'd54046, 16'd25815, 16'd9432, 16'd17533, 16'd37932, 16'd58217, 16'd18613, 16'd18385, 16'd31383});
	test_expansion(128'h255610a5cd67850f535499afa93ef090, {16'd12596, 16'd5849, 16'd21607, 16'd42840, 16'd12797, 16'd48210, 16'd51930, 16'd16020, 16'd3896, 16'd56653, 16'd49827, 16'd14180, 16'd34110, 16'd65256, 16'd62501, 16'd6648, 16'd13607, 16'd23145, 16'd38243, 16'd3939, 16'd7063, 16'd30433, 16'd48901, 16'd33609, 16'd62564, 16'd20130});
	test_expansion(128'haf9b69d64602bbcc138cfca65911414d, {16'd63203, 16'd53611, 16'd1646, 16'd62358, 16'd45608, 16'd2369, 16'd13417, 16'd1939, 16'd28653, 16'd42161, 16'd38551, 16'd12349, 16'd41299, 16'd13119, 16'd39609, 16'd17810, 16'd62392, 16'd3160, 16'd45902, 16'd28446, 16'd9920, 16'd50258, 16'd49386, 16'd63025, 16'd34286, 16'd6363});
	test_expansion(128'h7cbe2ef0553244fb6e3d9476d8640948, {16'd64951, 16'd32502, 16'd3411, 16'd57713, 16'd31266, 16'd26020, 16'd30703, 16'd42376, 16'd24454, 16'd60333, 16'd50575, 16'd16357, 16'd33190, 16'd40808, 16'd50154, 16'd50558, 16'd49591, 16'd16928, 16'd55082, 16'd57718, 16'd1117, 16'd27382, 16'd20102, 16'd29449, 16'd64758, 16'd63127});
	test_expansion(128'hd2d3bea7c350f351397006aa695a6351, {16'd45656, 16'd39001, 16'd52237, 16'd60540, 16'd59792, 16'd39551, 16'd23298, 16'd44093, 16'd21158, 16'd1910, 16'd59397, 16'd11285, 16'd24102, 16'd42401, 16'd64837, 16'd51232, 16'd33019, 16'd28680, 16'd61624, 16'd25232, 16'd60510, 16'd45974, 16'd16351, 16'd28733, 16'd19773, 16'd24586});
	test_expansion(128'h74bafd840c61402beb33eac7c29a16f5, {16'd751, 16'd9724, 16'd9773, 16'd13166, 16'd17341, 16'd3092, 16'd4111, 16'd30445, 16'd63202, 16'd48889, 16'd50606, 16'd41363, 16'd30668, 16'd62613, 16'd40504, 16'd9906, 16'd65314, 16'd55931, 16'd27400, 16'd27622, 16'd64258, 16'd26735, 16'd7093, 16'd57154, 16'd9895, 16'd16412});
	test_expansion(128'h80d9fe382a7da297a12076ad62aa9cfc, {16'd39128, 16'd19434, 16'd58290, 16'd9941, 16'd49462, 16'd22891, 16'd13377, 16'd62204, 16'd42729, 16'd18357, 16'd19604, 16'd45302, 16'd23109, 16'd24272, 16'd54858, 16'd61690, 16'd23921, 16'd32523, 16'd43742, 16'd17394, 16'd2758, 16'd24240, 16'd40244, 16'd6460, 16'd24094, 16'd42735});
	test_expansion(128'h114f8bbfc9fa05dfbb201129e8ed27b8, {16'd32003, 16'd63411, 16'd9103, 16'd19633, 16'd15882, 16'd62604, 16'd5911, 16'd13063, 16'd27553, 16'd97, 16'd51885, 16'd40212, 16'd16309, 16'd65155, 16'd43860, 16'd52230, 16'd56528, 16'd54619, 16'd53313, 16'd54365, 16'd7562, 16'd63709, 16'd28670, 16'd28760, 16'd39011, 16'd58121});
	test_expansion(128'hb2d98d315bb97e6fb5f97ae08792150b, {16'd28855, 16'd43751, 16'd49458, 16'd34022, 16'd25950, 16'd56164, 16'd24072, 16'd9687, 16'd4143, 16'd1008, 16'd8709, 16'd57637, 16'd15336, 16'd44098, 16'd58551, 16'd6588, 16'd48702, 16'd54083, 16'd57553, 16'd29930, 16'd23915, 16'd64878, 16'd4810, 16'd62719, 16'd35492, 16'd4240});
	test_expansion(128'h2f85f1b31a69aa2c1030bcb170421df3, {16'd62115, 16'd24808, 16'd61188, 16'd8684, 16'd27877, 16'd50203, 16'd18291, 16'd47825, 16'd8456, 16'd52932, 16'd43976, 16'd29776, 16'd52519, 16'd44607, 16'd20727, 16'd65505, 16'd57449, 16'd39776, 16'd51526, 16'd55889, 16'd9322, 16'd33635, 16'd20718, 16'd44245, 16'd4896, 16'd32736});
	test_expansion(128'hbeeaa96a37938aa723b31f00aa32ad88, {16'd32515, 16'd48450, 16'd9371, 16'd26952, 16'd24212, 16'd28910, 16'd64487, 16'd43254, 16'd49956, 16'd44516, 16'd44851, 16'd33353, 16'd26692, 16'd42090, 16'd19464, 16'd25145, 16'd35838, 16'd33028, 16'd41621, 16'd29460, 16'd54248, 16'd52504, 16'd54257, 16'd35517, 16'd52969, 16'd50202});
	test_expansion(128'h9f2455df9d4033e35382ad376fe7e9b0, {16'd5256, 16'd35654, 16'd14793, 16'd61868, 16'd24544, 16'd60168, 16'd4493, 16'd30647, 16'd54268, 16'd1092, 16'd7055, 16'd53405, 16'd2332, 16'd64617, 16'd33009, 16'd5288, 16'd12301, 16'd58628, 16'd55323, 16'd50094, 16'd61954, 16'd54578, 16'd50682, 16'd215, 16'd56801, 16'd21627});
	test_expansion(128'h3baad58ba9b3487f88ce13cf182af78f, {16'd38586, 16'd12269, 16'd6549, 16'd50316, 16'd6831, 16'd40251, 16'd41714, 16'd56471, 16'd55894, 16'd45490, 16'd34979, 16'd2420, 16'd26652, 16'd44371, 16'd33698, 16'd49125, 16'd49509, 16'd48158, 16'd47023, 16'd42016, 16'd46522, 16'd48019, 16'd42243, 16'd9340, 16'd217, 16'd19022});
	test_expansion(128'h98407fbe0bb605a9bf38d76fd0c25783, {16'd64330, 16'd51721, 16'd21353, 16'd12360, 16'd45532, 16'd10918, 16'd41620, 16'd28310, 16'd794, 16'd29291, 16'd61502, 16'd53220, 16'd2090, 16'd60477, 16'd22074, 16'd32189, 16'd39057, 16'd42855, 16'd40830, 16'd24690, 16'd20029, 16'd55447, 16'd12626, 16'd52225, 16'd47289, 16'd62336});
	test_expansion(128'he322b81be7959fd4972d75128e164f01, {16'd49517, 16'd25767, 16'd4621, 16'd44531, 16'd25393, 16'd27088, 16'd61336, 16'd31008, 16'd65070, 16'd13318, 16'd20369, 16'd18722, 16'd43304, 16'd42127, 16'd31257, 16'd38209, 16'd5650, 16'd8698, 16'd38031, 16'd980, 16'd1012, 16'd55628, 16'd53352, 16'd26791, 16'd45124, 16'd60899});
	test_expansion(128'hf00bc46e979b697a3dbfecc70edc6d22, {16'd51600, 16'd8042, 16'd63636, 16'd36290, 16'd51372, 16'd26912, 16'd8979, 16'd29919, 16'd44865, 16'd60267, 16'd49281, 16'd25294, 16'd52702, 16'd6839, 16'd63452, 16'd39861, 16'd18944, 16'd23630, 16'd25854, 16'd12359, 16'd49782, 16'd6362, 16'd324, 16'd21691, 16'd41104, 16'd37759});
	test_expansion(128'hd8415af4f1cd663ba4715d44a06ad309, {16'd54093, 16'd22608, 16'd12626, 16'd64044, 16'd46676, 16'd24780, 16'd63447, 16'd30025, 16'd41351, 16'd26119, 16'd30210, 16'd26006, 16'd30485, 16'd20776, 16'd60645, 16'd18345, 16'd65475, 16'd30252, 16'd39193, 16'd39266, 16'd51734, 16'd10062, 16'd43616, 16'd61961, 16'd8916, 16'd41775});
	test_expansion(128'hd40a202c7cc2a4dcc75ed68f62ad52e9, {16'd13961, 16'd54365, 16'd18195, 16'd16769, 16'd39798, 16'd2300, 16'd63440, 16'd46632, 16'd44743, 16'd5885, 16'd41641, 16'd41614, 16'd13706, 16'd37747, 16'd6658, 16'd43488, 16'd19990, 16'd53133, 16'd60313, 16'd47733, 16'd49287, 16'd28511, 16'd45031, 16'd22356, 16'd38434, 16'd41777});
	test_expansion(128'hc9b3a77619d20bcd87a17882a38926b0, {16'd9472, 16'd17524, 16'd49778, 16'd17059, 16'd19358, 16'd52015, 16'd51429, 16'd31594, 16'd59118, 16'd36194, 16'd34880, 16'd64268, 16'd56768, 16'd25376, 16'd18816, 16'd963, 16'd2596, 16'd61296, 16'd14282, 16'd53695, 16'd51113, 16'd8226, 16'd14762, 16'd20823, 16'd65339, 16'd47227});
	test_expansion(128'h03de9f5abb7020b7ab8fac0663105799, {16'd39671, 16'd7884, 16'd15446, 16'd34340, 16'd20124, 16'd62990, 16'd6701, 16'd6076, 16'd18911, 16'd48519, 16'd18782, 16'd24548, 16'd34582, 16'd6104, 16'd11055, 16'd62220, 16'd25413, 16'd60187, 16'd61957, 16'd45624, 16'd45720, 16'd43500, 16'd28314, 16'd1499, 16'd17701, 16'd32277});
	test_expansion(128'haf91b1123d0c8ed0a447bdb5a777a0c9, {16'd58235, 16'd43898, 16'd58943, 16'd45138, 16'd37293, 16'd28659, 16'd47377, 16'd34126, 16'd2872, 16'd19291, 16'd11389, 16'd19613, 16'd34428, 16'd12244, 16'd60188, 16'd30217, 16'd38904, 16'd26852, 16'd30287, 16'd30239, 16'd53957, 16'd34010, 16'd9556, 16'd13108, 16'd39324, 16'd39940});
	test_expansion(128'hca4507ecc85770b13e46b3af194f4353, {16'd58538, 16'd30566, 16'd12775, 16'd36145, 16'd16358, 16'd25645, 16'd60055, 16'd27445, 16'd16799, 16'd17920, 16'd4301, 16'd35718, 16'd48677, 16'd65461, 16'd59140, 16'd679, 16'd19211, 16'd57911, 16'd21588, 16'd38147, 16'd39134, 16'd43447, 16'd41798, 16'd7737, 16'd63896, 16'd33541});
	test_expansion(128'h1c29c390368b1ab8dc8869b7175aed1d, {16'd33586, 16'd37003, 16'd17612, 16'd31617, 16'd31262, 16'd4796, 16'd46124, 16'd15629, 16'd30891, 16'd1412, 16'd13950, 16'd57804, 16'd13460, 16'd35198, 16'd37584, 16'd32689, 16'd50808, 16'd20622, 16'd13522, 16'd7475, 16'd17778, 16'd60846, 16'd37280, 16'd5614, 16'd12356, 16'd46479});
	test_expansion(128'he3edb3bcdcf8714efb15de41b5ca7fad, {16'd57045, 16'd28848, 16'd3382, 16'd58669, 16'd4233, 16'd44470, 16'd35895, 16'd10150, 16'd16148, 16'd60419, 16'd58998, 16'd18892, 16'd5392, 16'd37089, 16'd45448, 16'd35798, 16'd2743, 16'd12341, 16'd4276, 16'd42553, 16'd65055, 16'd65348, 16'd2728, 16'd48130, 16'd32770, 16'd8547});
	test_expansion(128'h5e370972d435080416bbbe8fe52616e3, {16'd42560, 16'd57185, 16'd43266, 16'd62815, 16'd36594, 16'd38272, 16'd32992, 16'd64897, 16'd56040, 16'd60784, 16'd11987, 16'd6965, 16'd45316, 16'd39597, 16'd13186, 16'd18232, 16'd28037, 16'd17328, 16'd2516, 16'd23424, 16'd6318, 16'd38354, 16'd32880, 16'd18535, 16'd995, 16'd49282});
	test_expansion(128'hfffbb429c2c6a39bae6188201183d137, {16'd27412, 16'd58815, 16'd26831, 16'd20450, 16'd30901, 16'd43281, 16'd12014, 16'd48244, 16'd57854, 16'd24623, 16'd31784, 16'd54603, 16'd23505, 16'd19246, 16'd7538, 16'd49974, 16'd51, 16'd52651, 16'd7973, 16'd36552, 16'd61405, 16'd23139, 16'd20256, 16'd26201, 16'd4932, 16'd59899});
	test_expansion(128'h62c0a714d55f5e25fa8fcaeca82f6138, {16'd11522, 16'd29327, 16'd6756, 16'd12925, 16'd24246, 16'd64568, 16'd50236, 16'd50975, 16'd7493, 16'd59844, 16'd24039, 16'd49146, 16'd16198, 16'd17424, 16'd7189, 16'd38079, 16'd32981, 16'd43085, 16'd19197, 16'd40089, 16'd28150, 16'd22078, 16'd46119, 16'd65389, 16'd64619, 16'd52084});
	test_expansion(128'hc1ae7299200d693c1abd48d8bdb828af, {16'd53885, 16'd48174, 16'd55868, 16'd591, 16'd20938, 16'd25910, 16'd43839, 16'd29041, 16'd30205, 16'd58546, 16'd1339, 16'd15285, 16'd39958, 16'd47532, 16'd47126, 16'd15231, 16'd35435, 16'd38643, 16'd62375, 16'd9018, 16'd48194, 16'd29009, 16'd9932, 16'd55851, 16'd18208, 16'd25294});
	test_expansion(128'h2c551af55971bd7a76fbd04ecd6663e7, {16'd32050, 16'd33306, 16'd1322, 16'd55741, 16'd42624, 16'd34050, 16'd40567, 16'd8728, 16'd4445, 16'd32077, 16'd28881, 16'd34396, 16'd36666, 16'd57456, 16'd26632, 16'd10477, 16'd8177, 16'd33188, 16'd12754, 16'd48963, 16'd21476, 16'd63396, 16'd9550, 16'd24797, 16'd3513, 16'd32780});
	test_expansion(128'h31891ba7e68eb96e14378b84b4ff9943, {16'd63002, 16'd37554, 16'd58922, 16'd42605, 16'd8507, 16'd34430, 16'd37892, 16'd43455, 16'd39909, 16'd45751, 16'd32710, 16'd24112, 16'd49502, 16'd14599, 16'd2668, 16'd3871, 16'd58547, 16'd50648, 16'd36356, 16'd32993, 16'd4936, 16'd862, 16'd55134, 16'd27947, 16'd46386, 16'd14219});
	test_expansion(128'he82eb752e1fa6cf2a4d4f7ec7f4254c1, {16'd27862, 16'd9719, 16'd22006, 16'd1117, 16'd56402, 16'd45435, 16'd7338, 16'd55877, 16'd58367, 16'd54432, 16'd58938, 16'd2195, 16'd35375, 16'd59743, 16'd11418, 16'd51766, 16'd30514, 16'd57331, 16'd22501, 16'd23864, 16'd33185, 16'd41717, 16'd54528, 16'd8160, 16'd49016, 16'd12217});
	test_expansion(128'h59083ec7a916e22739342ce568732748, {16'd4896, 16'd10443, 16'd34720, 16'd60082, 16'd49723, 16'd23660, 16'd13124, 16'd6860, 16'd1403, 16'd6583, 16'd60507, 16'd9249, 16'd5695, 16'd42302, 16'd35817, 16'd19943, 16'd32416, 16'd36091, 16'd55534, 16'd41212, 16'd3919, 16'd5466, 16'd29844, 16'd26217, 16'd2364, 16'd32835});
	test_expansion(128'heead9244b5f6744036aaddc9ebc96853, {16'd23832, 16'd24691, 16'd42550, 16'd65166, 16'd15222, 16'd16033, 16'd41978, 16'd27052, 16'd29111, 16'd64830, 16'd45716, 16'd27406, 16'd59885, 16'd7813, 16'd29518, 16'd54519, 16'd8611, 16'd43849, 16'd42306, 16'd31760, 16'd2945, 16'd57444, 16'd49981, 16'd56044, 16'd27768, 16'd37657});
	test_expansion(128'h634fd80b673d8d658fb0dbb81a237113, {16'd63575, 16'd14644, 16'd17475, 16'd42859, 16'd57805, 16'd28894, 16'd34273, 16'd58068, 16'd17277, 16'd33042, 16'd3780, 16'd64708, 16'd56827, 16'd57501, 16'd6646, 16'd33440, 16'd18265, 16'd3365, 16'd42846, 16'd26124, 16'd58787, 16'd61862, 16'd62039, 16'd17101, 16'd46570, 16'd20303});
	test_expansion(128'h9a06c72986ac63c9b3993dead660b049, {16'd17922, 16'd13799, 16'd37556, 16'd2350, 16'd49936, 16'd50087, 16'd32614, 16'd40127, 16'd11817, 16'd25003, 16'd6606, 16'd51007, 16'd11744, 16'd41056, 16'd33217, 16'd737, 16'd30333, 16'd19103, 16'd41468, 16'd53801, 16'd50003, 16'd27545, 16'd44839, 16'd20266, 16'd57235, 16'd30733});
	test_expansion(128'h7a39582feeb9ce786ba73e7c6a172899, {16'd35464, 16'd7009, 16'd54963, 16'd45818, 16'd41788, 16'd28504, 16'd2839, 16'd14111, 16'd40883, 16'd29017, 16'd53474, 16'd45632, 16'd52247, 16'd18285, 16'd62488, 16'd4657, 16'd63334, 16'd29045, 16'd11172, 16'd33297, 16'd16298, 16'd28527, 16'd7394, 16'd3388, 16'd8925, 16'd5000});
	test_expansion(128'haf801592d7315c17ebd50505385117c1, {16'd24785, 16'd17878, 16'd32133, 16'd24105, 16'd45556, 16'd64120, 16'd18470, 16'd54036, 16'd60363, 16'd35899, 16'd40830, 16'd54728, 16'd51787, 16'd44250, 16'd55166, 16'd56395, 16'd26206, 16'd63561, 16'd19605, 16'd11735, 16'd49157, 16'd63514, 16'd61376, 16'd49512, 16'd37142, 16'd21229});
	test_expansion(128'h06dd493471336ddb694cac87cad3e691, {16'd49762, 16'd31826, 16'd23100, 16'd63167, 16'd13709, 16'd30242, 16'd40455, 16'd14099, 16'd47500, 16'd48867, 16'd64425, 16'd27108, 16'd33289, 16'd63527, 16'd22640, 16'd52684, 16'd25451, 16'd15831, 16'd17772, 16'd49065, 16'd21221, 16'd20234, 16'd63413, 16'd63753, 16'd41356, 16'd19132});
	test_expansion(128'he6d78b367282ed636f6991a4f3d9b8a3, {16'd63985, 16'd47616, 16'd32992, 16'd17926, 16'd7932, 16'd49083, 16'd40713, 16'd30025, 16'd10908, 16'd51461, 16'd24175, 16'd13259, 16'd2327, 16'd5278, 16'd7547, 16'd20474, 16'd14868, 16'd42766, 16'd27685, 16'd45809, 16'd24029, 16'd15777, 16'd58891, 16'd55031, 16'd56395, 16'd59070});
	test_expansion(128'h9543059472d341a159dfc15d1b3e0778, {16'd49422, 16'd59634, 16'd6228, 16'd56713, 16'd44840, 16'd19235, 16'd57081, 16'd38972, 16'd23038, 16'd30266, 16'd26117, 16'd46977, 16'd48051, 16'd47398, 16'd54584, 16'd54321, 16'd12918, 16'd52259, 16'd20332, 16'd10071, 16'd65059, 16'd48638, 16'd21801, 16'd6368, 16'd62851, 16'd30698});
	test_expansion(128'h85ef49ee009f39b67ac67fc76beb3aa3, {16'd20595, 16'd43695, 16'd64230, 16'd16286, 16'd48597, 16'd58987, 16'd34980, 16'd46285, 16'd15102, 16'd52357, 16'd45187, 16'd6550, 16'd34376, 16'd47774, 16'd43231, 16'd63022, 16'd32356, 16'd27755, 16'd55159, 16'd7387, 16'd46338, 16'd58770, 16'd48356, 16'd15444, 16'd20267, 16'd64835});
	test_expansion(128'hae865550dd522fb75a75260d520a00e4, {16'd46840, 16'd30773, 16'd63256, 16'd61981, 16'd40323, 16'd26868, 16'd10704, 16'd22037, 16'd49210, 16'd9301, 16'd26203, 16'd62667, 16'd20656, 16'd31320, 16'd48959, 16'd1666, 16'd54708, 16'd19537, 16'd61898, 16'd52641, 16'd16491, 16'd11975, 16'd27408, 16'd16068, 16'd2275, 16'd6946});
	test_expansion(128'h12b6f9ab112238223ed56e0f334d42af, {16'd11157, 16'd45966, 16'd45944, 16'd7097, 16'd38288, 16'd30333, 16'd44999, 16'd1910, 16'd52004, 16'd54467, 16'd31259, 16'd57376, 16'd39344, 16'd7721, 16'd52682, 16'd38988, 16'd9449, 16'd88, 16'd36366, 16'd14616, 16'd56309, 16'd7678, 16'd14524, 16'd61861, 16'd49318, 16'd40892});
	test_expansion(128'h6503a4facf61e1ff53f08992aaea369b, {16'd15685, 16'd6407, 16'd32012, 16'd59025, 16'd20149, 16'd40929, 16'd46778, 16'd25262, 16'd26318, 16'd63527, 16'd4444, 16'd45161, 16'd15445, 16'd27142, 16'd27923, 16'd16034, 16'd36451, 16'd40131, 16'd29852, 16'd56619, 16'd62286, 16'd10743, 16'd25700, 16'd46954, 16'd64020, 16'd22212});
	test_expansion(128'h23dab1a300b26c64e88696487e4b0ead, {16'd14382, 16'd48080, 16'd46442, 16'd4473, 16'd35761, 16'd42350, 16'd27528, 16'd11559, 16'd24911, 16'd54413, 16'd28994, 16'd33993, 16'd26706, 16'd11611, 16'd42660, 16'd43099, 16'd31732, 16'd15698, 16'd16766, 16'd41044, 16'd27280, 16'd27140, 16'd8998, 16'd32453, 16'd874, 16'd26342});
	test_expansion(128'h8cae69cb85e9712ab7bcd5508f02361c, {16'd48609, 16'd285, 16'd42684, 16'd3923, 16'd40949, 16'd62803, 16'd37334, 16'd22765, 16'd57080, 16'd63626, 16'd8674, 16'd28401, 16'd20302, 16'd1374, 16'd23940, 16'd23165, 16'd56678, 16'd56569, 16'd58720, 16'd6260, 16'd32704, 16'd6845, 16'd46140, 16'd5583, 16'd18847, 16'd38547});
	test_expansion(128'h388078904aa8a9afef5117db3a587b18, {16'd15700, 16'd14052, 16'd30669, 16'd40286, 16'd14776, 16'd49196, 16'd34570, 16'd24537, 16'd1254, 16'd13733, 16'd132, 16'd8389, 16'd22942, 16'd10772, 16'd11809, 16'd44697, 16'd26561, 16'd34237, 16'd23645, 16'd20814, 16'd15569, 16'd65441, 16'd56646, 16'd17810, 16'd48634, 16'd39759});
	test_expansion(128'hfb748cd59e32393fccd4d023146313c9, {16'd63058, 16'd10528, 16'd7988, 16'd2593, 16'd60382, 16'd61467, 16'd3985, 16'd21378, 16'd39710, 16'd28313, 16'd10887, 16'd30010, 16'd58494, 16'd31553, 16'd19813, 16'd23808, 16'd58106, 16'd24481, 16'd56247, 16'd30584, 16'd40963, 16'd11370, 16'd50574, 16'd27079, 16'd3156, 16'd44794});
	test_expansion(128'ha71a9e2cf73b86866b53eb36f410435b, {16'd9485, 16'd3037, 16'd40737, 16'd48203, 16'd6223, 16'd38313, 16'd11037, 16'd35528, 16'd9266, 16'd26718, 16'd34575, 16'd3799, 16'd52286, 16'd38897, 16'd19832, 16'd1046, 16'd29333, 16'd15674, 16'd64493, 16'd34166, 16'd23904, 16'd62385, 16'd48638, 16'd19475, 16'd42112, 16'd1342});
	test_expansion(128'h7fbfd359aa1132b07fe3a774d41ddf97, {16'd32311, 16'd11657, 16'd10460, 16'd4334, 16'd53940, 16'd24902, 16'd46320, 16'd32337, 16'd49910, 16'd56218, 16'd12101, 16'd50267, 16'd11314, 16'd25195, 16'd33548, 16'd29908, 16'd60219, 16'd2892, 16'd35650, 16'd16574, 16'd40557, 16'd24386, 16'd38307, 16'd11322, 16'd27107, 16'd57649});
	test_expansion(128'hbcbf815217157ad46b45ea5e5437f783, {16'd6979, 16'd29748, 16'd11338, 16'd55002, 16'd64322, 16'd53442, 16'd34328, 16'd2338, 16'd36184, 16'd61604, 16'd53924, 16'd33398, 16'd51356, 16'd25846, 16'd45098, 16'd62243, 16'd36897, 16'd35403, 16'd12312, 16'd4385, 16'd24409, 16'd16345, 16'd46188, 16'd43858, 16'd47743, 16'd7444});
	test_expansion(128'h833cbfadc05ff9acf73c50611feb864a, {16'd36925, 16'd59656, 16'd58978, 16'd4186, 16'd63386, 16'd55335, 16'd22265, 16'd57792, 16'd16980, 16'd12446, 16'd23040, 16'd26910, 16'd1495, 16'd2527, 16'd16655, 16'd8618, 16'd32160, 16'd36108, 16'd57492, 16'd55457, 16'd44126, 16'd28803, 16'd39723, 16'd7000, 16'd16919, 16'd28973});
	test_expansion(128'h161653289cecf921c2ce80f61f0f8b2d, {16'd45226, 16'd14796, 16'd29795, 16'd25343, 16'd52788, 16'd28016, 16'd50095, 16'd14754, 16'd63542, 16'd8054, 16'd61137, 16'd52362, 16'd21146, 16'd39983, 16'd40939, 16'd51917, 16'd64427, 16'd26263, 16'd55378, 16'd10770, 16'd42863, 16'd59627, 16'd63192, 16'd39123, 16'd13009, 16'd54178});
	test_expansion(128'h114d48af5be6afed7e729aee372a4d16, {16'd8577, 16'd16646, 16'd42609, 16'd10472, 16'd417, 16'd805, 16'd26153, 16'd32712, 16'd53745, 16'd6860, 16'd44244, 16'd15464, 16'd28163, 16'd9958, 16'd22566, 16'd35610, 16'd25158, 16'd9263, 16'd2024, 16'd63027, 16'd19547, 16'd64486, 16'd61247, 16'd11052, 16'd39737, 16'd8199});
	test_expansion(128'h35e3528de92eafec3e59de4c56f722bc, {16'd55097, 16'd3965, 16'd59339, 16'd23183, 16'd16473, 16'd25193, 16'd59190, 16'd19331, 16'd13495, 16'd63272, 16'd9735, 16'd56407, 16'd41750, 16'd2493, 16'd55360, 16'd4370, 16'd51125, 16'd39800, 16'd20005, 16'd115, 16'd16324, 16'd46123, 16'd33674, 16'd19496, 16'd24900, 16'd22499});
	test_expansion(128'hacd4ddc190e9d1c2c15423366985fd2d, {16'd23920, 16'd27505, 16'd61112, 16'd57646, 16'd49288, 16'd31256, 16'd63263, 16'd21101, 16'd26250, 16'd5843, 16'd57063, 16'd33923, 16'd34509, 16'd32551, 16'd14939, 16'd17710, 16'd53531, 16'd48817, 16'd17271, 16'd55529, 16'd10258, 16'd36972, 16'd30080, 16'd31944, 16'd46104, 16'd37766});
	test_expansion(128'h343f73a11d7c411f5e674fc4e0feaed9, {16'd14807, 16'd37578, 16'd15450, 16'd21042, 16'd23331, 16'd1644, 16'd18938, 16'd3660, 16'd26895, 16'd54018, 16'd11503, 16'd30790, 16'd61602, 16'd4699, 16'd12235, 16'd45703, 16'd27149, 16'd7276, 16'd41493, 16'd45424, 16'd39445, 16'd59776, 16'd7152, 16'd6767, 16'd34151, 16'd29604});
	test_expansion(128'h26be3d523b2c091154a370a58470098f, {16'd1986, 16'd48120, 16'd9577, 16'd47922, 16'd38099, 16'd44793, 16'd26433, 16'd61490, 16'd2515, 16'd37174, 16'd62354, 16'd60561, 16'd49475, 16'd16780, 16'd7563, 16'd26020, 16'd3135, 16'd36380, 16'd59619, 16'd7524, 16'd15017, 16'd35, 16'd31366, 16'd64129, 16'd17925, 16'd46478});
	test_expansion(128'h14219c76c1f607d4ee4619dc37ebf2eb, {16'd4754, 16'd33046, 16'd60195, 16'd37848, 16'd35202, 16'd21329, 16'd56467, 16'd40377, 16'd30648, 16'd65058, 16'd27551, 16'd59912, 16'd26679, 16'd23957, 16'd13810, 16'd54734, 16'd51534, 16'd58200, 16'd36557, 16'd58916, 16'd30305, 16'd45899, 16'd54506, 16'd17674, 16'd15050, 16'd7893});
	test_expansion(128'hce2b2a2fd1ca5645b72274fabf6ed0a6, {16'd48360, 16'd49131, 16'd40866, 16'd64296, 16'd38654, 16'd8152, 16'd9627, 16'd7165, 16'd42526, 16'd58122, 16'd43238, 16'd28344, 16'd35272, 16'd23674, 16'd29438, 16'd63611, 16'd36489, 16'd33273, 16'd5146, 16'd20549, 16'd26272, 16'd64081, 16'd6488, 16'd57911, 16'd20832, 16'd32808});
	test_expansion(128'hc09bc014fd121b5ec098c14704c0829a, {16'd40903, 16'd55809, 16'd58975, 16'd8777, 16'd58912, 16'd45688, 16'd3798, 16'd24174, 16'd45284, 16'd65470, 16'd58332, 16'd15687, 16'd30949, 16'd27013, 16'd28134, 16'd56314, 16'd9484, 16'd32082, 16'd59469, 16'd15671, 16'd17964, 16'd30789, 16'd24615, 16'd40463, 16'd58690, 16'd55368});
	test_expansion(128'heeef3409163720756311c28fa13f2dab, {16'd19210, 16'd21801, 16'd11950, 16'd62875, 16'd30280, 16'd22698, 16'd7565, 16'd50445, 16'd62327, 16'd23444, 16'd10101, 16'd30748, 16'd5855, 16'd32462, 16'd43384, 16'd14377, 16'd17525, 16'd55323, 16'd65505, 16'd43827, 16'd52277, 16'd55030, 16'd12306, 16'd35150, 16'd28912, 16'd34253});
	test_expansion(128'he06b3875d0d861e63807887ff97ec5b0, {16'd22819, 16'd31935, 16'd1247, 16'd47323, 16'd38509, 16'd10492, 16'd32309, 16'd4013, 16'd53134, 16'd17541, 16'd16200, 16'd44034, 16'd5578, 16'd39042, 16'd48154, 16'd20889, 16'd12179, 16'd7712, 16'd2826, 16'd51000, 16'd38764, 16'd20164, 16'd23164, 16'd58946, 16'd9292, 16'd49609});
	test_expansion(128'hcafd203b0cbd925edd7c2be2e4ed8daf, {16'd63443, 16'd18483, 16'd59345, 16'd22399, 16'd59186, 16'd43318, 16'd30258, 16'd48290, 16'd56568, 16'd64380, 16'd54296, 16'd43504, 16'd31045, 16'd56271, 16'd16861, 16'd28278, 16'd6121, 16'd33294, 16'd3928, 16'd318, 16'd31794, 16'd62744, 16'd24532, 16'd52021, 16'd31894, 16'd32124});
	test_expansion(128'h3dfe08810b36af4684d63d4d52ee2a4a, {16'd19832, 16'd36291, 16'd45801, 16'd15526, 16'd24046, 16'd36434, 16'd16939, 16'd9461, 16'd33624, 16'd40077, 16'd5668, 16'd55844, 16'd34158, 16'd48298, 16'd2939, 16'd64213, 16'd5631, 16'd37436, 16'd47005, 16'd56910, 16'd38829, 16'd42253, 16'd31476, 16'd60630, 16'd35235, 16'd24234});
	test_expansion(128'h1d812ba80f27fd6fabf7cb293578d3f7, {16'd50137, 16'd46320, 16'd49164, 16'd15113, 16'd47237, 16'd7627, 16'd58864, 16'd35310, 16'd63794, 16'd17454, 16'd714, 16'd11625, 16'd37028, 16'd18376, 16'd63965, 16'd52167, 16'd28773, 16'd36342, 16'd6674, 16'd14376, 16'd62642, 16'd4943, 16'd26240, 16'd62686, 16'd2326, 16'd32747});
	test_expansion(128'h0d8aa5281797a81d4ee5a39b374db752, {16'd23808, 16'd45469, 16'd13593, 16'd9445, 16'd56706, 16'd575, 16'd43269, 16'd2101, 16'd11186, 16'd15054, 16'd23174, 16'd11039, 16'd50464, 16'd64463, 16'd60945, 16'd10329, 16'd32889, 16'd25163, 16'd33854, 16'd47289, 16'd38375, 16'd57044, 16'd58740, 16'd116, 16'd6472, 16'd56966});
	test_expansion(128'h50d4a20e8e2d20181dba044c97dd71fa, {16'd48382, 16'd56617, 16'd13052, 16'd10562, 16'd56071, 16'd49755, 16'd33193, 16'd32403, 16'd31218, 16'd25176, 16'd38951, 16'd33492, 16'd8620, 16'd7955, 16'd44535, 16'd50444, 16'd136, 16'd17378, 16'd25589, 16'd16502, 16'd27968, 16'd1305, 16'd1215, 16'd1830, 16'd15194, 16'd6369});
	test_expansion(128'hfcfeba905d3bb4ac6f09ff77a52bd031, {16'd59885, 16'd26528, 16'd21058, 16'd13308, 16'd10665, 16'd51804, 16'd39926, 16'd21457, 16'd41229, 16'd64808, 16'd20563, 16'd39106, 16'd52930, 16'd62532, 16'd8030, 16'd15919, 16'd365, 16'd41902, 16'd40978, 16'd54476, 16'd23367, 16'd38313, 16'd1726, 16'd35613, 16'd347, 16'd23352});
	test_expansion(128'h0da17e5358541dc54d33f1a7614e4c41, {16'd47408, 16'd25470, 16'd51970, 16'd19271, 16'd6053, 16'd34990, 16'd43365, 16'd58385, 16'd55423, 16'd35174, 16'd45669, 16'd29447, 16'd32061, 16'd30696, 16'd51066, 16'd24213, 16'd12522, 16'd62734, 16'd54652, 16'd38222, 16'd30701, 16'd60251, 16'd2041, 16'd36805, 16'd12210, 16'd1323});
	test_expansion(128'h71535402c7227e82dfc5ca7d96edda17, {16'd39071, 16'd2296, 16'd52737, 16'd42073, 16'd24057, 16'd29914, 16'd924, 16'd34311, 16'd332, 16'd59796, 16'd28814, 16'd19164, 16'd35390, 16'd38278, 16'd36360, 16'd32921, 16'd62842, 16'd17070, 16'd31032, 16'd13760, 16'd9108, 16'd28043, 16'd31074, 16'd23848, 16'd30084, 16'd29791});
	test_expansion(128'h6f2289807112ecbc6e9139a026409a7b, {16'd42681, 16'd44209, 16'd1664, 16'd35445, 16'd19748, 16'd8625, 16'd61067, 16'd18261, 16'd58994, 16'd33839, 16'd39850, 16'd55792, 16'd407, 16'd62203, 16'd756, 16'd46719, 16'd25638, 16'd37580, 16'd61736, 16'd30997, 16'd57632, 16'd33514, 16'd3156, 16'd2523, 16'd22577, 16'd14994});
	test_expansion(128'hb1e1e813760c50f7fbd34129f3d693b3, {16'd25204, 16'd32571, 16'd56951, 16'd44838, 16'd29824, 16'd22623, 16'd18553, 16'd59406, 16'd27582, 16'd48931, 16'd15239, 16'd62558, 16'd29422, 16'd32937, 16'd33613, 16'd45191, 16'd4399, 16'd6004, 16'd10237, 16'd48236, 16'd879, 16'd4480, 16'd55648, 16'd27299, 16'd39474, 16'd47768});
	test_expansion(128'hf50fc10034ec91fdb8ea7589f4a9797f, {16'd36979, 16'd43819, 16'd17314, 16'd47161, 16'd1496, 16'd37733, 16'd38066, 16'd27512, 16'd12354, 16'd56088, 16'd60145, 16'd28257, 16'd9316, 16'd64292, 16'd15609, 16'd20993, 16'd3244, 16'd16718, 16'd28891, 16'd22468, 16'd54793, 16'd45904, 16'd36480, 16'd35786, 16'd29946, 16'd32070});
	test_expansion(128'h819b5fb6158da2ae445ec09b0961e8cb, {16'd10358, 16'd63720, 16'd45527, 16'd54362, 16'd64193, 16'd9920, 16'd32619, 16'd51664, 16'd13635, 16'd50447, 16'd13535, 16'd11552, 16'd31401, 16'd50208, 16'd36704, 16'd30759, 16'd50020, 16'd40284, 16'd33219, 16'd10010, 16'd57370, 16'd48420, 16'd28979, 16'd52320, 16'd52872, 16'd60570});
	test_expansion(128'h350ddbf14090701dca8ec4a6a811ef65, {16'd18690, 16'd53950, 16'd29318, 16'd51151, 16'd26564, 16'd57041, 16'd65426, 16'd50014, 16'd42279, 16'd46382, 16'd58533, 16'd27341, 16'd47094, 16'd10860, 16'd28509, 16'd50437, 16'd46964, 16'd31896, 16'd24221, 16'd16886, 16'd55121, 16'd15827, 16'd33292, 16'd43539, 16'd55484, 16'd24268});
	test_expansion(128'h174c17bd0fbab6b6904fa7851b62ea29, {16'd37546, 16'd33508, 16'd4840, 16'd33044, 16'd8303, 16'd53932, 16'd29066, 16'd502, 16'd6983, 16'd45936, 16'd10247, 16'd4653, 16'd39467, 16'd54175, 16'd6989, 16'd52382, 16'd54851, 16'd8321, 16'd20579, 16'd31750, 16'd32454, 16'd19643, 16'd23507, 16'd56704, 16'd11885, 16'd3748});
	test_expansion(128'h51d6054430ec34cb262837904177a119, {16'd9087, 16'd20851, 16'd34457, 16'd38491, 16'd53991, 16'd22900, 16'd50187, 16'd28359, 16'd45951, 16'd63799, 16'd53594, 16'd11425, 16'd13742, 16'd59073, 16'd36339, 16'd57837, 16'd38109, 16'd107, 16'd48785, 16'd9381, 16'd16578, 16'd2362, 16'd26429, 16'd49183, 16'd8898, 16'd52767});
	test_expansion(128'hc37fe108f409ac13985d093f89ae8eeb, {16'd12504, 16'd7681, 16'd28923, 16'd36591, 16'd33333, 16'd45955, 16'd59521, 16'd4016, 16'd55056, 16'd36449, 16'd52066, 16'd51106, 16'd11377, 16'd18819, 16'd918, 16'd8680, 16'd23558, 16'd31845, 16'd34310, 16'd28338, 16'd62104, 16'd56848, 16'd17084, 16'd4251, 16'd47003, 16'd29801});
	test_expansion(128'h157ca7ff2c45c6211a7cd8943f499a31, {16'd45390, 16'd9824, 16'd49945, 16'd35673, 16'd58394, 16'd55467, 16'd23439, 16'd37983, 16'd44537, 16'd44300, 16'd24237, 16'd19770, 16'd31329, 16'd51580, 16'd50169, 16'd1037, 16'd31678, 16'd24664, 16'd35816, 16'd31298, 16'd63410, 16'd18259, 16'd23458, 16'd22932, 16'd45900, 16'd60119});
	test_expansion(128'h49cda6ea81ef5ae0216298e04a2f3f4f, {16'd58156, 16'd41958, 16'd43352, 16'd2412, 16'd44954, 16'd29273, 16'd27308, 16'd4426, 16'd43407, 16'd30488, 16'd29590, 16'd14934, 16'd49758, 16'd48475, 16'd44203, 16'd10629, 16'd35597, 16'd61604, 16'd44421, 16'd47946, 16'd57858, 16'd11083, 16'd17160, 16'd25738, 16'd33002, 16'd4399});
	test_expansion(128'h2e8fd0d017d980d7eec0f131feeefdda, {16'd21048, 16'd13395, 16'd16855, 16'd11031, 16'd18228, 16'd9733, 16'd50503, 16'd53534, 16'd24579, 16'd46377, 16'd44774, 16'd52953, 16'd62143, 16'd56596, 16'd14861, 16'd38487, 16'd47094, 16'd33077, 16'd2605, 16'd45269, 16'd43219, 16'd18203, 16'd24934, 16'd16496, 16'd57590, 16'd37691});
	test_expansion(128'hdeff64b741137f050c7ed766b1589087, {16'd43354, 16'd57762, 16'd961, 16'd3054, 16'd44884, 16'd24515, 16'd42163, 16'd1115, 16'd13543, 16'd29140, 16'd62431, 16'd45117, 16'd61499, 16'd18339, 16'd908, 16'd28840, 16'd4961, 16'd54411, 16'd19430, 16'd23483, 16'd7272, 16'd12880, 16'd2637, 16'd25224, 16'd14108, 16'd46238});
	test_expansion(128'hf29a590cdc80424e2e9a3dc3e42c5187, {16'd57706, 16'd10446, 16'd60342, 16'd48161, 16'd7548, 16'd13209, 16'd45582, 16'd30702, 16'd17624, 16'd12205, 16'd64896, 16'd13204, 16'd48477, 16'd34861, 16'd61271, 16'd40989, 16'd7426, 16'd64197, 16'd48529, 16'd16830, 16'd31306, 16'd64755, 16'd23360, 16'd61836, 16'd26217, 16'd61629});
	test_expansion(128'hfb26e89d091d73e3579bd52a058973f2, {16'd1559, 16'd38193, 16'd20140, 16'd60380, 16'd57789, 16'd20044, 16'd18171, 16'd27773, 16'd4143, 16'd44518, 16'd28144, 16'd3817, 16'd54844, 16'd34559, 16'd34153, 16'd41983, 16'd8524, 16'd53507, 16'd47380, 16'd26632, 16'd1693, 16'd6629, 16'd62651, 16'd2556, 16'd26960, 16'd53495});
	test_expansion(128'hc6ec4d49b13699c886f682266a08f7df, {16'd29028, 16'd2550, 16'd1211, 16'd4907, 16'd33516, 16'd59257, 16'd32530, 16'd12461, 16'd3755, 16'd47504, 16'd41470, 16'd59142, 16'd19111, 16'd53684, 16'd33564, 16'd6724, 16'd32918, 16'd31413, 16'd60178, 16'd16972, 16'd18606, 16'd48165, 16'd39436, 16'd47209, 16'd9061, 16'd19686});
	test_expansion(128'h1f7537e0d22dc11a5af7a05279dd67ff, {16'd238, 16'd17284, 16'd11838, 16'd408, 16'd61842, 16'd63049, 16'd23965, 16'd37066, 16'd58421, 16'd8682, 16'd6847, 16'd21972, 16'd45956, 16'd31188, 16'd1268, 16'd24547, 16'd7465, 16'd20243, 16'd12465, 16'd61541, 16'd5341, 16'd38877, 16'd65389, 16'd7270, 16'd22368, 16'd35129});
	test_expansion(128'h4ac02b9c824b2f6e179cbe7307e3a30b, {16'd26056, 16'd35573, 16'd43096, 16'd55275, 16'd18540, 16'd47131, 16'd1406, 16'd64157, 16'd56665, 16'd7503, 16'd65, 16'd48653, 16'd60619, 16'd36504, 16'd52121, 16'd4168, 16'd22581, 16'd45197, 16'd52721, 16'd50183, 16'd39764, 16'd60209, 16'd64520, 16'd44141, 16'd61205, 16'd55147});
	test_expansion(128'h05d815d1855cdf5bd48c5dfd2a683db4, {16'd38884, 16'd28155, 16'd57628, 16'd30682, 16'd7230, 16'd18813, 16'd57918, 16'd51835, 16'd42346, 16'd58383, 16'd2810, 16'd11380, 16'd3793, 16'd2991, 16'd56961, 16'd12229, 16'd50591, 16'd52290, 16'd34821, 16'd18750, 16'd63100, 16'd22224, 16'd16143, 16'd12681, 16'd49559, 16'd62120});
	test_expansion(128'h28bcca56446b2500b26a048ed6645d01, {16'd41247, 16'd37953, 16'd29599, 16'd49544, 16'd55796, 16'd61240, 16'd48549, 16'd56959, 16'd48897, 16'd3076, 16'd1386, 16'd9385, 16'd27403, 16'd45999, 16'd17741, 16'd13760, 16'd27510, 16'd19643, 16'd63329, 16'd40585, 16'd53319, 16'd9581, 16'd13400, 16'd6297, 16'd62668, 16'd1309});
	test_expansion(128'h249998fbec875c4921bdc06b7926f0e5, {16'd10910, 16'd55145, 16'd23036, 16'd55889, 16'd3261, 16'd65174, 16'd39487, 16'd64804, 16'd13505, 16'd31442, 16'd60910, 16'd33610, 16'd48361, 16'd29041, 16'd33347, 16'd10345, 16'd10689, 16'd42939, 16'd19928, 16'd58715, 16'd13228, 16'd54230, 16'd24240, 16'd49818, 16'd14855, 16'd60037});
	test_expansion(128'h8e69fa2319249fbead2d76bff64ec4d1, {16'd33742, 16'd26242, 16'd31025, 16'd39926, 16'd16277, 16'd52751, 16'd13822, 16'd6319, 16'd49739, 16'd26887, 16'd46838, 16'd49046, 16'd18248, 16'd56128, 16'd39670, 16'd19828, 16'd47687, 16'd59492, 16'd2721, 16'd12999, 16'd4465, 16'd43368, 16'd46111, 16'd32263, 16'd35543, 16'd54304});
	test_expansion(128'haa7051aba4315287ac1a357830f52d10, {16'd16789, 16'd27446, 16'd49422, 16'd52188, 16'd5352, 16'd61287, 16'd61478, 16'd56083, 16'd61308, 16'd30911, 16'd5542, 16'd41316, 16'd7683, 16'd28872, 16'd30784, 16'd26549, 16'd14477, 16'd33728, 16'd55961, 16'd61638, 16'd2546, 16'd26385, 16'd35698, 16'd48677, 16'd20528, 16'd10727});
	test_expansion(128'hec1268a7078647e68ff205aceb33bf94, {16'd55023, 16'd22613, 16'd26594, 16'd32489, 16'd25380, 16'd34049, 16'd60406, 16'd37682, 16'd59420, 16'd16012, 16'd33289, 16'd45054, 16'd31999, 16'd54498, 16'd11346, 16'd50934, 16'd21759, 16'd5359, 16'd58877, 16'd37414, 16'd22375, 16'd3725, 16'd33502, 16'd983, 16'd19522, 16'd7868});
	test_expansion(128'h4fc39486ba498ab65baeff3eb8ee0727, {16'd18560, 16'd19849, 16'd58339, 16'd65412, 16'd20312, 16'd42536, 16'd35582, 16'd51194, 16'd60626, 16'd6961, 16'd53822, 16'd10063, 16'd6918, 16'd42254, 16'd11635, 16'd27768, 16'd52002, 16'd44559, 16'd48487, 16'd63551, 16'd28577, 16'd38250, 16'd33746, 16'd60570, 16'd24142, 16'd33530});
	test_expansion(128'h21367112601999e7a03d370a4c6a970d, {16'd52007, 16'd6429, 16'd1019, 16'd41336, 16'd63231, 16'd43476, 16'd9429, 16'd47978, 16'd46226, 16'd13935, 16'd58207, 16'd58058, 16'd59953, 16'd13917, 16'd42394, 16'd59632, 16'd56842, 16'd32928, 16'd16532, 16'd1199, 16'd40940, 16'd3148, 16'd47343, 16'd13675, 16'd46881, 16'd21206});
	test_expansion(128'hf578c2c37e073d5ca0e4ed9c258550fd, {16'd39852, 16'd27764, 16'd45732, 16'd34026, 16'd11522, 16'd36288, 16'd19619, 16'd2826, 16'd43386, 16'd20731, 16'd58938, 16'd1150, 16'd39898, 16'd56782, 16'd40080, 16'd48409, 16'd3643, 16'd17569, 16'd27505, 16'd33827, 16'd52263, 16'd57657, 16'd58554, 16'd24299, 16'd52551, 16'd46245});
	test_expansion(128'h7983362c4df60e7059eb4b834b71da30, {16'd4870, 16'd49721, 16'd36215, 16'd44173, 16'd13900, 16'd8831, 16'd38463, 16'd51050, 16'd62517, 16'd58931, 16'd3410, 16'd13759, 16'd34313, 16'd51033, 16'd37695, 16'd1763, 16'd30433, 16'd37267, 16'd19271, 16'd7116, 16'd4048, 16'd27287, 16'd43205, 16'd4613, 16'd23925, 16'd42987});
	test_expansion(128'h88fcdf83ed215a0cd3b44ed98e8f5d77, {16'd12078, 16'd21372, 16'd53789, 16'd52251, 16'd42610, 16'd28393, 16'd18155, 16'd55580, 16'd59183, 16'd50721, 16'd12742, 16'd59773, 16'd13122, 16'd27293, 16'd59730, 16'd17285, 16'd9220, 16'd8333, 16'd37385, 16'd29188, 16'd34280, 16'd60491, 16'd19413, 16'd29372, 16'd6470, 16'd50669});
	test_expansion(128'h0346f15e0df5e72a7f62637c1fd4da62, {16'd2665, 16'd20090, 16'd59403, 16'd63638, 16'd41959, 16'd29010, 16'd27245, 16'd6307, 16'd34397, 16'd28806, 16'd10668, 16'd62794, 16'd7258, 16'd21681, 16'd18635, 16'd63840, 16'd57074, 16'd46487, 16'd47458, 16'd60936, 16'd5137, 16'd25529, 16'd23373, 16'd52927, 16'd29865, 16'd25350});
	test_expansion(128'h48bb68a63d05c01d721aa3b320f199d5, {16'd52548, 16'd5084, 16'd5115, 16'd32246, 16'd4012, 16'd7077, 16'd31335, 16'd5948, 16'd21182, 16'd51880, 16'd21648, 16'd58621, 16'd8245, 16'd9501, 16'd12690, 16'd32960, 16'd60426, 16'd30607, 16'd40648, 16'd9883, 16'd58958, 16'd29640, 16'd12391, 16'd40526, 16'd27076, 16'd5554});
	test_expansion(128'h76e0bc09c1df8ef72a014717f57f2bd8, {16'd59141, 16'd43455, 16'd34430, 16'd41766, 16'd47480, 16'd13811, 16'd62515, 16'd33922, 16'd12699, 16'd55508, 16'd55222, 16'd51651, 16'd57689, 16'd59974, 16'd25461, 16'd8918, 16'd8008, 16'd58931, 16'd64708, 16'd55727, 16'd32654, 16'd8130, 16'd45306, 16'd45243, 16'd48787, 16'd33238});
	test_expansion(128'hd7620f55bd25ac432394678d27cef5df, {16'd15716, 16'd1590, 16'd32141, 16'd39596, 16'd65073, 16'd13822, 16'd2661, 16'd27003, 16'd23810, 16'd54931, 16'd26940, 16'd47102, 16'd21221, 16'd23155, 16'd17938, 16'd12149, 16'd33571, 16'd2215, 16'd49243, 16'd42371, 16'd25680, 16'd17671, 16'd8029, 16'd19850, 16'd26465, 16'd62694});
	test_expansion(128'hb63dd4e9d860078666e9f130d0644e12, {16'd63224, 16'd15234, 16'd43665, 16'd22944, 16'd47532, 16'd28315, 16'd32617, 16'd32349, 16'd10996, 16'd1974, 16'd24160, 16'd2428, 16'd15321, 16'd2597, 16'd2024, 16'd17780, 16'd16041, 16'd36554, 16'd39990, 16'd25843, 16'd26229, 16'd60022, 16'd44308, 16'd31588, 16'd22798, 16'd44822});
	test_expansion(128'h986f5d7656bc1c6960375fea94a2fed9, {16'd52349, 16'd47054, 16'd22033, 16'd26079, 16'd8837, 16'd35379, 16'd1522, 16'd19907, 16'd63507, 16'd59795, 16'd9903, 16'd56840, 16'd13663, 16'd5090, 16'd62356, 16'd34764, 16'd58514, 16'd35597, 16'd35512, 16'd30787, 16'd64486, 16'd8165, 16'd22407, 16'd29078, 16'd58402, 16'd41622});
	test_expansion(128'h4ca66e891653a56aabc0997065500093, {16'd55082, 16'd30259, 16'd8459, 16'd61621, 16'd1208, 16'd60827, 16'd42114, 16'd21578, 16'd18395, 16'd27445, 16'd28493, 16'd59127, 16'd20353, 16'd60668, 16'd47358, 16'd40472, 16'd4739, 16'd21771, 16'd22447, 16'd36490, 16'd35099, 16'd18675, 16'd20243, 16'd18442, 16'd60187, 16'd45941});
	test_expansion(128'hf5cbf2c160cfe388f1c4a0b8e4bd9fa1, {16'd62491, 16'd60295, 16'd44574, 16'd41128, 16'd50242, 16'd31037, 16'd23187, 16'd40459, 16'd7744, 16'd62582, 16'd60385, 16'd64501, 16'd25638, 16'd63530, 16'd11310, 16'd18544, 16'd40594, 16'd48632, 16'd48146, 16'd2206, 16'd24796, 16'd50294, 16'd35664, 16'd7603, 16'd17604, 16'd17749});
	test_expansion(128'hd846f8e02e3d0c75bc2fde63d4f8175a, {16'd36517, 16'd12501, 16'd31363, 16'd53809, 16'd45950, 16'd2598, 16'd3748, 16'd61955, 16'd31300, 16'd18785, 16'd50964, 16'd14543, 16'd63775, 16'd21437, 16'd5110, 16'd13789, 16'd10839, 16'd40951, 16'd7685, 16'd25931, 16'd14499, 16'd27175, 16'd27095, 16'd47874, 16'd16728, 16'd28194});
	test_expansion(128'hd5ac8f972e243ed2db57a5ed8d745cee, {16'd46986, 16'd16188, 16'd4523, 16'd11453, 16'd42148, 16'd14254, 16'd13939, 16'd59654, 16'd60376, 16'd18620, 16'd48396, 16'd4567, 16'd147, 16'd50787, 16'd43080, 16'd40671, 16'd110, 16'd9335, 16'd26313, 16'd28474, 16'd35728, 16'd51014, 16'd40577, 16'd26745, 16'd40454, 16'd17337});
	test_expansion(128'h6717c3396eeac41399d3daad0b2f1f7d, {16'd38049, 16'd22329, 16'd43964, 16'd27135, 16'd60507, 16'd23357, 16'd18262, 16'd3149, 16'd25137, 16'd27769, 16'd61713, 16'd49481, 16'd26289, 16'd4532, 16'd1138, 16'd54638, 16'd3250, 16'd1759, 16'd64292, 16'd32937, 16'd42118, 16'd11119, 16'd42922, 16'd59391, 16'd13381, 16'd27762});
	test_expansion(128'h16ce4fd1b1570f1e39b4d357588feca9, {16'd21108, 16'd16754, 16'd14917, 16'd58361, 16'd16290, 16'd30035, 16'd3255, 16'd40108, 16'd26592, 16'd36782, 16'd17410, 16'd59798, 16'd24452, 16'd39781, 16'd36698, 16'd30456, 16'd31152, 16'd56402, 16'd51972, 16'd64365, 16'd58591, 16'd31898, 16'd5376, 16'd46522, 16'd16683, 16'd11058});
	test_expansion(128'h393c33350ece6d603fc90869291e0d8d, {16'd8373, 16'd56602, 16'd16965, 16'd26197, 16'd2810, 16'd14776, 16'd52644, 16'd52919, 16'd3064, 16'd18850, 16'd40463, 16'd29926, 16'd63973, 16'd50470, 16'd6732, 16'd46476, 16'd50888, 16'd54668, 16'd34761, 16'd61463, 16'd60342, 16'd44110, 16'd7005, 16'd40471, 16'd42037, 16'd60507});
	test_expansion(128'h23938d2542129e0acffc791ecc906606, {16'd24026, 16'd52987, 16'd46239, 16'd11343, 16'd40239, 16'd59948, 16'd41453, 16'd27693, 16'd48523, 16'd15089, 16'd34946, 16'd44129, 16'd38115, 16'd12160, 16'd42516, 16'd15393, 16'd15120, 16'd36285, 16'd15677, 16'd14412, 16'd61823, 16'd44840, 16'd1340, 16'd16628, 16'd600, 16'd58745});
	test_expansion(128'h56095b37b091456e7bab421aaeb57ae0, {16'd3465, 16'd2038, 16'd30851, 16'd6686, 16'd266, 16'd30883, 16'd38486, 16'd63766, 16'd21013, 16'd45172, 16'd60225, 16'd64901, 16'd2631, 16'd48016, 16'd30174, 16'd2412, 16'd11441, 16'd19003, 16'd63393, 16'd10296, 16'd32957, 16'd27806, 16'd38189, 16'd26032, 16'd37507, 16'd36309});
	test_expansion(128'h616fd83ea9310baf689fa62b2e1c57ae, {16'd30783, 16'd268, 16'd12967, 16'd15481, 16'd20638, 16'd55249, 16'd51121, 16'd26083, 16'd9453, 16'd41718, 16'd38566, 16'd48920, 16'd19933, 16'd39413, 16'd33125, 16'd32578, 16'd59176, 16'd2181, 16'd53043, 16'd58423, 16'd42270, 16'd19099, 16'd5484, 16'd3448, 16'd37301, 16'd62564});
	test_expansion(128'hd4667b6a38abfe32787ca07dd36906d4, {16'd19330, 16'd25778, 16'd44275, 16'd42729, 16'd31964, 16'd61389, 16'd9981, 16'd39810, 16'd51184, 16'd27753, 16'd1399, 16'd12042, 16'd37323, 16'd20436, 16'd10269, 16'd19427, 16'd57543, 16'd63000, 16'd65283, 16'd11945, 16'd4598, 16'd52589, 16'd19376, 16'd42551, 16'd30942, 16'd20299});
	test_expansion(128'h226ca49f32667e37cf65f0a1d1f360f2, {16'd50496, 16'd24446, 16'd34911, 16'd35544, 16'd51611, 16'd51701, 16'd16460, 16'd45046, 16'd23354, 16'd28974, 16'd61273, 16'd51498, 16'd50584, 16'd1309, 16'd2694, 16'd8064, 16'd64357, 16'd66, 16'd55752, 16'd2494, 16'd54175, 16'd19764, 16'd23430, 16'd32555, 16'd36741, 16'd36716});
	test_expansion(128'h120837e3eacfea2dfe7a291846a51cde, {16'd20309, 16'd33080, 16'd60443, 16'd49555, 16'd26390, 16'd51395, 16'd45494, 16'd57185, 16'd23943, 16'd56566, 16'd54709, 16'd1553, 16'd25257, 16'd12441, 16'd40026, 16'd33478, 16'd28792, 16'd37099, 16'd23163, 16'd45801, 16'd519, 16'd27013, 16'd1126, 16'd31474, 16'd21383, 16'd21995});
	test_expansion(128'h1b833bce57c38458195d9e47b4cba172, {16'd8034, 16'd3585, 16'd27464, 16'd46213, 16'd6722, 16'd40570, 16'd62011, 16'd58536, 16'd2145, 16'd26393, 16'd31006, 16'd37220, 16'd21019, 16'd46353, 16'd36652, 16'd40041, 16'd54082, 16'd18407, 16'd41798, 16'd24869, 16'd47625, 16'd7365, 16'd6783, 16'd36268, 16'd42440, 16'd43718});
	test_expansion(128'h9f7f616fd7b5c44fdbb830fe357df8a9, {16'd46902, 16'd22499, 16'd43985, 16'd23889, 16'd21457, 16'd13414, 16'd55842, 16'd38226, 16'd41284, 16'd56057, 16'd37797, 16'd11812, 16'd10583, 16'd13175, 16'd7435, 16'd11703, 16'd57498, 16'd57801, 16'd4918, 16'd47270, 16'd50466, 16'd9960, 16'd584, 16'd19589, 16'd46572, 16'd17104});
	test_expansion(128'h27428e44e77e334c61b32435e0f6133a, {16'd21965, 16'd44266, 16'd25643, 16'd51634, 16'd9912, 16'd6027, 16'd7705, 16'd5683, 16'd38698, 16'd60647, 16'd62000, 16'd46652, 16'd40995, 16'd4223, 16'd26920, 16'd2770, 16'd10762, 16'd36624, 16'd24450, 16'd41365, 16'd60548, 16'd48167, 16'd50230, 16'd11877, 16'd47611, 16'd56725});
	test_expansion(128'hae02d189c47255f4530b76a8a0c11938, {16'd3944, 16'd18434, 16'd47095, 16'd47139, 16'd38991, 16'd1714, 16'd36284, 16'd47148, 16'd6547, 16'd41217, 16'd44527, 16'd24113, 16'd9465, 16'd20253, 16'd44106, 16'd52335, 16'd41096, 16'd37914, 16'd44079, 16'd50100, 16'd56852, 16'd6578, 16'd45921, 16'd19907, 16'd14008, 16'd56410});
	test_expansion(128'h921bc1aee3ab5fdc0062a788276c1c21, {16'd54441, 16'd43819, 16'd40836, 16'd30790, 16'd22707, 16'd58602, 16'd28111, 16'd6913, 16'd34404, 16'd26932, 16'd7573, 16'd12855, 16'd23103, 16'd57502, 16'd64024, 16'd7783, 16'd50225, 16'd31681, 16'd12765, 16'd48333, 16'd52404, 16'd14425, 16'd63001, 16'd61683, 16'd55653, 16'd48787});
	test_expansion(128'h540c7c51516217ff2b0e88821fee0191, {16'd50646, 16'd62937, 16'd9288, 16'd4148, 16'd20069, 16'd41511, 16'd55270, 16'd2103, 16'd43812, 16'd6339, 16'd54251, 16'd227, 16'd1068, 16'd5252, 16'd40432, 16'd16808, 16'd52203, 16'd41061, 16'd40742, 16'd19470, 16'd964, 16'd2973, 16'd29047, 16'd44647, 16'd21333, 16'd4550});
	test_expansion(128'h9a23f45e4bd0fb2072f0d1ac393610b5, {16'd58785, 16'd28953, 16'd35946, 16'd13798, 16'd56844, 16'd6315, 16'd1065, 16'd56087, 16'd13622, 16'd5120, 16'd18725, 16'd4878, 16'd48909, 16'd47085, 16'd32875, 16'd25220, 16'd8874, 16'd47413, 16'd9250, 16'd23415, 16'd7772, 16'd16374, 16'd46355, 16'd43615, 16'd60481, 16'd59234});
	test_expansion(128'hff4fdfe01eb27f691b7785219cf80527, {16'd1461, 16'd24933, 16'd12689, 16'd29612, 16'd31722, 16'd62206, 16'd36802, 16'd7619, 16'd52468, 16'd21136, 16'd64921, 16'd40141, 16'd62710, 16'd41660, 16'd51066, 16'd2817, 16'd555, 16'd49533, 16'd49451, 16'd48913, 16'd54974, 16'd52044, 16'd33740, 16'd35688, 16'd32029, 16'd50646});
	test_expansion(128'h27e0e6066a5c21166a5cba670a865bcd, {16'd25642, 16'd38489, 16'd63074, 16'd35124, 16'd58452, 16'd26402, 16'd56459, 16'd14297, 16'd29461, 16'd45942, 16'd64048, 16'd30931, 16'd62850, 16'd52718, 16'd7161, 16'd25968, 16'd55693, 16'd55774, 16'd54843, 16'd12430, 16'd19507, 16'd48056, 16'd5259, 16'd61956, 16'd43714, 16'd3349});
	test_expansion(128'he8a3a99a1e11cc71c3ecfd3aa0b6f12f, {16'd28724, 16'd45278, 16'd31690, 16'd10997, 16'd2229, 16'd30169, 16'd5531, 16'd61998, 16'd20856, 16'd49506, 16'd65221, 16'd29677, 16'd46540, 16'd4168, 16'd11769, 16'd40824, 16'd57309, 16'd64877, 16'd8881, 16'd33242, 16'd52814, 16'd43536, 16'd50348, 16'd33033, 16'd5106, 16'd17153});
	test_expansion(128'h768d7dafa4e1fbc808f7a57d8a9a6cb2, {16'd291, 16'd31836, 16'd59137, 16'd40825, 16'd43105, 16'd45300, 16'd17396, 16'd49159, 16'd36723, 16'd63360, 16'd25266, 16'd36452, 16'd39775, 16'd53200, 16'd645, 16'd1469, 16'd24697, 16'd5832, 16'd42409, 16'd61977, 16'd48199, 16'd31148, 16'd12738, 16'd10603, 16'd46502, 16'd44559});
	test_expansion(128'hb143dc8f34f14582df509f31f02a7231, {16'd23354, 16'd35693, 16'd50919, 16'd54466, 16'd23940, 16'd9092, 16'd35574, 16'd63777, 16'd48466, 16'd8122, 16'd57036, 16'd30799, 16'd56624, 16'd53810, 16'd11524, 16'd11417, 16'd62559, 16'd50536, 16'd2793, 16'd34704, 16'd43018, 16'd17577, 16'd62222, 16'd6567, 16'd44428, 16'd54303});
	test_expansion(128'h0c6c32d6cfb077d86673e8c3dc19f911, {16'd13447, 16'd1499, 16'd45541, 16'd10039, 16'd62795, 16'd52254, 16'd11682, 16'd13246, 16'd6679, 16'd55563, 16'd29998, 16'd54429, 16'd36484, 16'd41927, 16'd284, 16'd39205, 16'd11376, 16'd13015, 16'd8895, 16'd41857, 16'd41453, 16'd17058, 16'd46933, 16'd59421, 16'd62717, 16'd46438});
	test_expansion(128'h47589e97f5155480cca11b8b737f2806, {16'd48750, 16'd33943, 16'd62972, 16'd57929, 16'd57268, 16'd59397, 16'd25750, 16'd23632, 16'd30579, 16'd56692, 16'd53940, 16'd65108, 16'd48326, 16'd63835, 16'd35440, 16'd53967, 16'd51717, 16'd26174, 16'd51641, 16'd47208, 16'd19582, 16'd23513, 16'd2148, 16'd33602, 16'd17847, 16'd17002});
	test_expansion(128'he71dff640b4245a07dae309e8d93e6a3, {16'd50934, 16'd16653, 16'd30982, 16'd17268, 16'd33584, 16'd24990, 16'd684, 16'd56190, 16'd41870, 16'd36180, 16'd55801, 16'd42817, 16'd24111, 16'd32559, 16'd22680, 16'd38254, 16'd2368, 16'd26036, 16'd25900, 16'd20947, 16'd57797, 16'd15063, 16'd9978, 16'd25579, 16'd17604, 16'd47525});
	test_expansion(128'h133bd6f94afe92de7addb03e6f57f8c9, {16'd31827, 16'd22486, 16'd5930, 16'd53872, 16'd64737, 16'd56133, 16'd30626, 16'd22314, 16'd7405, 16'd37301, 16'd5639, 16'd29218, 16'd14772, 16'd759, 16'd52844, 16'd16224, 16'd27177, 16'd64731, 16'd13110, 16'd1543, 16'd63158, 16'd50027, 16'd41488, 16'd741, 16'd64046, 16'd42065});
	test_expansion(128'hda0ac9c47085099985e686f1b24a7ceb, {16'd53720, 16'd2295, 16'd22055, 16'd27296, 16'd9756, 16'd55674, 16'd22580, 16'd50422, 16'd14919, 16'd37587, 16'd7635, 16'd3072, 16'd46704, 16'd58001, 16'd38758, 16'd48449, 16'd8372, 16'd30892, 16'd28510, 16'd47796, 16'd27306, 16'd17348, 16'd64519, 16'd20433, 16'd41565, 16'd27737});
	test_expansion(128'h6b3de17d71c89a174aa2953cd0d48c15, {16'd47347, 16'd25176, 16'd55355, 16'd5796, 16'd3999, 16'd39059, 16'd58464, 16'd23417, 16'd60730, 16'd20793, 16'd63075, 16'd55726, 16'd41960, 16'd10440, 16'd40907, 16'd55903, 16'd17116, 16'd15529, 16'd5429, 16'd57587, 16'd53275, 16'd4069, 16'd11692, 16'd13584, 16'd2709, 16'd60512});
	test_expansion(128'hc310037631fe137d3cf292e431079df2, {16'd43121, 16'd59756, 16'd1198, 16'd24088, 16'd24886, 16'd64574, 16'd38884, 16'd8542, 16'd52860, 16'd10790, 16'd60761, 16'd16084, 16'd13299, 16'd29367, 16'd40426, 16'd57078, 16'd20257, 16'd20243, 16'd41881, 16'd16637, 16'd42528, 16'd38727, 16'd64841, 16'd37547, 16'd58054, 16'd59416});
	test_expansion(128'h5f23a9084bc6d4c0023f7fddf01658f0, {16'd59979, 16'd50769, 16'd60317, 16'd63718, 16'd35324, 16'd22127, 16'd8442, 16'd7180, 16'd64843, 16'd47870, 16'd3086, 16'd12668, 16'd1676, 16'd52380, 16'd61669, 16'd8483, 16'd61303, 16'd2362, 16'd21751, 16'd18723, 16'd12126, 16'd46575, 16'd2403, 16'd35689, 16'd22723, 16'd42797});
	test_expansion(128'hbb44f0269d7968dced2d9d0dd8e62861, {16'd45889, 16'd55692, 16'd19191, 16'd30626, 16'd3526, 16'd53651, 16'd10859, 16'd9678, 16'd32323, 16'd45169, 16'd34156, 16'd45955, 16'd30130, 16'd30014, 16'd15783, 16'd16171, 16'd48379, 16'd57277, 16'd23842, 16'd36734, 16'd7181, 16'd29217, 16'd25387, 16'd35754, 16'd2825, 16'd34820});
	test_expansion(128'hca142251bf2edf84c5e504926d7e4580, {16'd12579, 16'd43305, 16'd33559, 16'd54932, 16'd49936, 16'd3137, 16'd41906, 16'd47044, 16'd14913, 16'd40624, 16'd51099, 16'd18132, 16'd34116, 16'd6422, 16'd51784, 16'd65431, 16'd25183, 16'd4705, 16'd21484, 16'd53138, 16'd1897, 16'd55789, 16'd49235, 16'd5550, 16'd2163, 16'd4803});
	test_expansion(128'hf19c1813d22e62b2eea72468713b9c8a, {16'd7911, 16'd26298, 16'd51155, 16'd36883, 16'd4091, 16'd35197, 16'd20022, 16'd57954, 16'd42781, 16'd40886, 16'd17881, 16'd53613, 16'd49524, 16'd49112, 16'd6665, 16'd615, 16'd22600, 16'd63441, 16'd23042, 16'd59683, 16'd62090, 16'd11273, 16'd17484, 16'd53101, 16'd25806, 16'd41013});
	test_expansion(128'hf800d20600fb708b14fd75b1e330776c, {16'd47487, 16'd23695, 16'd63104, 16'd15864, 16'd21911, 16'd2270, 16'd29046, 16'd26899, 16'd27312, 16'd29945, 16'd20277, 16'd21739, 16'd42012, 16'd9514, 16'd59759, 16'd63684, 16'd58034, 16'd20851, 16'd32285, 16'd19368, 16'd22070, 16'd6839, 16'd61289, 16'd26735, 16'd38047, 16'd63361});
	test_expansion(128'h825388eb993a9ac74c7c9161ebe31fa6, {16'd35413, 16'd39863, 16'd15381, 16'd22331, 16'd35641, 16'd49602, 16'd11247, 16'd64477, 16'd21406, 16'd43923, 16'd19349, 16'd20630, 16'd45346, 16'd18459, 16'd60835, 16'd36049, 16'd63334, 16'd26607, 16'd19895, 16'd36963, 16'd37182, 16'd37855, 16'd29837, 16'd10423, 16'd4474, 16'd44767});
	test_expansion(128'h7d0f78659e04a03c1345803ca41de1dc, {16'd13920, 16'd33241, 16'd51440, 16'd50656, 16'd45038, 16'd10345, 16'd54916, 16'd50052, 16'd2831, 16'd15010, 16'd13052, 16'd62998, 16'd37913, 16'd31178, 16'd41609, 16'd30083, 16'd38838, 16'd60396, 16'd59283, 16'd51989, 16'd15718, 16'd21470, 16'd52499, 16'd51466, 16'd37337, 16'd17480});
	test_expansion(128'h077ff498d996b9a44c832e5b2bd2b323, {16'd64005, 16'd58978, 16'd63217, 16'd46625, 16'd53846, 16'd18445, 16'd57349, 16'd65162, 16'd23556, 16'd17479, 16'd58536, 16'd643, 16'd41810, 16'd44286, 16'd64125, 16'd20394, 16'd42636, 16'd65040, 16'd19807, 16'd11892, 16'd35464, 16'd5675, 16'd8496, 16'd10397, 16'd63582, 16'd56509});
	test_expansion(128'hcebdd2c20c68da89bdea03db253b715e, {16'd27122, 16'd6000, 16'd40787, 16'd10300, 16'd55118, 16'd46188, 16'd13420, 16'd30522, 16'd25306, 16'd2442, 16'd40042, 16'd48892, 16'd31385, 16'd21421, 16'd20819, 16'd2824, 16'd18053, 16'd7634, 16'd38525, 16'd34762, 16'd54320, 16'd11200, 16'd63792, 16'd50965, 16'd3940, 16'd55422});
	test_expansion(128'h7e8d43373399a06694eb25ca45c19a2b, {16'd27250, 16'd4338, 16'd2235, 16'd54490, 16'd48585, 16'd47723, 16'd7870, 16'd60318, 16'd10961, 16'd58073, 16'd34971, 16'd31439, 16'd44812, 16'd232, 16'd24206, 16'd4919, 16'd51001, 16'd35587, 16'd26243, 16'd18466, 16'd8649, 16'd6740, 16'd14718, 16'd9274, 16'd52044, 16'd27668});
	test_expansion(128'h78e5dad3121e840c80128aedc49bc86e, {16'd7018, 16'd13033, 16'd47737, 16'd5879, 16'd482, 16'd16631, 16'd50948, 16'd48565, 16'd50514, 16'd56277, 16'd7479, 16'd61584, 16'd60720, 16'd37755, 16'd14418, 16'd61973, 16'd23055, 16'd14132, 16'd42384, 16'd22695, 16'd61338, 16'd54669, 16'd14973, 16'd50629, 16'd519, 16'd42627});
	test_expansion(128'h9bd848e4c9f07da2c765f72a6379d814, {16'd1218, 16'd58781, 16'd27105, 16'd49401, 16'd50378, 16'd30259, 16'd5215, 16'd62904, 16'd54321, 16'd58821, 16'd39398, 16'd22339, 16'd11822, 16'd44231, 16'd8949, 16'd20817, 16'd24079, 16'd26927, 16'd48373, 16'd57205, 16'd21875, 16'd14322, 16'd28941, 16'd23205, 16'd22364, 16'd59231});
	test_expansion(128'hfb87cd24057d87fedba454b2f351d029, {16'd7707, 16'd7073, 16'd6123, 16'd38339, 16'd63283, 16'd55576, 16'd61873, 16'd53056, 16'd47914, 16'd50398, 16'd17057, 16'd37537, 16'd11156, 16'd11842, 16'd44948, 16'd28181, 16'd45923, 16'd7607, 16'd19, 16'd34049, 16'd24685, 16'd4465, 16'd25862, 16'd24385, 16'd1684, 16'd20274});
	test_expansion(128'h497c0cfd27da35517eeb515caa505f43, {16'd6817, 16'd47998, 16'd49536, 16'd27374, 16'd25012, 16'd33778, 16'd54296, 16'd34278, 16'd3372, 16'd43011, 16'd29876, 16'd30581, 16'd48035, 16'd60070, 16'd18524, 16'd64147, 16'd63265, 16'd43283, 16'd15659, 16'd32359, 16'd19223, 16'd3528, 16'd31634, 16'd16162, 16'd19365, 16'd54768});
	test_expansion(128'h8d329ea2b98b469fcd4e24120b56e0f3, {16'd22292, 16'd27528, 16'd53372, 16'd24993, 16'd26293, 16'd65180, 16'd55231, 16'd27180, 16'd54729, 16'd34217, 16'd37271, 16'd47167, 16'd1797, 16'd31099, 16'd15604, 16'd30265, 16'd56594, 16'd29064, 16'd39682, 16'd15337, 16'd37622, 16'd53451, 16'd19580, 16'd12836, 16'd17158, 16'd26712});
	test_expansion(128'h9c1d60e80599bd056fcd9b332224c832, {16'd12036, 16'd47452, 16'd36952, 16'd39769, 16'd21712, 16'd4573, 16'd43790, 16'd37985, 16'd61841, 16'd25846, 16'd34310, 16'd4162, 16'd42200, 16'd23180, 16'd60936, 16'd50607, 16'd41101, 16'd25562, 16'd49446, 16'd50495, 16'd65052, 16'd40093, 16'd8785, 16'd55679, 16'd62162, 16'd7486});
	test_expansion(128'h815a7557b39a961c6ea1258cd7f0c406, {16'd6939, 16'd38145, 16'd57853, 16'd2329, 16'd21466, 16'd62708, 16'd20559, 16'd42041, 16'd58362, 16'd27023, 16'd41910, 16'd46536, 16'd30854, 16'd38662, 16'd31458, 16'd21150, 16'd40679, 16'd1124, 16'd15425, 16'd63378, 16'd6395, 16'd30733, 16'd3796, 16'd61969, 16'd28529, 16'd3334});
	test_expansion(128'h0b5d25117e5aa8ee76b83312f40263e9, {16'd11152, 16'd34881, 16'd39334, 16'd19941, 16'd16147, 16'd32634, 16'd39175, 16'd35479, 16'd10400, 16'd2794, 16'd14035, 16'd24834, 16'd5596, 16'd36234, 16'd63034, 16'd54583, 16'd18324, 16'd23408, 16'd9066, 16'd1950, 16'd1692, 16'd60704, 16'd4571, 16'd48743, 16'd56002, 16'd44242});
	test_expansion(128'hcb1d457a8f214e6b0785696635a713e9, {16'd704, 16'd34909, 16'd57415, 16'd15227, 16'd46731, 16'd13665, 16'd36269, 16'd52482, 16'd12402, 16'd51501, 16'd38752, 16'd25539, 16'd25162, 16'd61700, 16'd40201, 16'd20621, 16'd12346, 16'd8738, 16'd22748, 16'd21955, 16'd16505, 16'd63751, 16'd8577, 16'd44100, 16'd41812, 16'd5237});
	test_expansion(128'haf6fef40b60d9d9f097588cd86accc56, {16'd41930, 16'd10105, 16'd2420, 16'd31773, 16'd38328, 16'd52172, 16'd64797, 16'd36960, 16'd14938, 16'd24356, 16'd26859, 16'd13814, 16'd48500, 16'd24659, 16'd59654, 16'd46216, 16'd10897, 16'd40897, 16'd11976, 16'd42727, 16'd18709, 16'd5420, 16'd11293, 16'd46791, 16'd38965, 16'd58089});
	test_expansion(128'h167084cb9da9aa8d6cb1d0e1241413e7, {16'd48915, 16'd11490, 16'd8979, 16'd60295, 16'd57344, 16'd39781, 16'd47703, 16'd62317, 16'd33958, 16'd46511, 16'd63171, 16'd21241, 16'd45587, 16'd14413, 16'd1703, 16'd55081, 16'd41975, 16'd16936, 16'd45283, 16'd59336, 16'd30997, 16'd45, 16'd34677, 16'd57340, 16'd62156, 16'd25931});
	test_expansion(128'h05d1b0610d747b0d2d0d220e00362700, {16'd16161, 16'd35333, 16'd9452, 16'd351, 16'd6807, 16'd48085, 16'd55002, 16'd31376, 16'd34706, 16'd53564, 16'd6618, 16'd7411, 16'd53765, 16'd27783, 16'd31214, 16'd32993, 16'd32213, 16'd29596, 16'd47992, 16'd11233, 16'd8223, 16'd27036, 16'd13583, 16'd35364, 16'd55971, 16'd40918});
	test_expansion(128'hbc34efbc111f26981d8556c61ad91315, {16'd64201, 16'd28710, 16'd26385, 16'd39022, 16'd38843, 16'd1191, 16'd18735, 16'd2677, 16'd45018, 16'd63707, 16'd3233, 16'd65055, 16'd64025, 16'd43478, 16'd14071, 16'd41912, 16'd55818, 16'd13591, 16'd3743, 16'd10576, 16'd24957, 16'd45777, 16'd38536, 16'd31123, 16'd33114, 16'd22064});
	test_expansion(128'h08b72b9ca483a8488c97b4049d26b03e, {16'd58283, 16'd22451, 16'd33321, 16'd53919, 16'd38755, 16'd42781, 16'd28528, 16'd52283, 16'd20888, 16'd59188, 16'd2909, 16'd21353, 16'd6683, 16'd64295, 16'd14361, 16'd1909, 16'd4391, 16'd47952, 16'd5827, 16'd19362, 16'd62483, 16'd43249, 16'd32760, 16'd34612, 16'd25178, 16'd62008});
	test_expansion(128'hc83a6bbb72b58c14beed1cdb144bd0c2, {16'd55145, 16'd31691, 16'd45968, 16'd52292, 16'd29949, 16'd44464, 16'd6247, 16'd45914, 16'd7372, 16'd45788, 16'd53974, 16'd43202, 16'd49442, 16'd26387, 16'd45657, 16'd48942, 16'd44076, 16'd62898, 16'd32532, 16'd64459, 16'd50400, 16'd3511, 16'd53783, 16'd922, 16'd19588, 16'd62259});
	test_expansion(128'h94fff2a3df4d0e69db29011a717b9385, {16'd48479, 16'd33377, 16'd10388, 16'd58528, 16'd51495, 16'd24094, 16'd39310, 16'd27521, 16'd28357, 16'd62325, 16'd46474, 16'd59260, 16'd22397, 16'd51089, 16'd12900, 16'd37630, 16'd36541, 16'd37929, 16'd19841, 16'd38899, 16'd52522, 16'd55664, 16'd17063, 16'd3506, 16'd21458, 16'd50265});
	test_expansion(128'he62b63527b58ee88c94f1596e4612c9e, {16'd51271, 16'd56888, 16'd26028, 16'd52313, 16'd59702, 16'd60433, 16'd849, 16'd65144, 16'd63334, 16'd31289, 16'd35512, 16'd61696, 16'd48793, 16'd11099, 16'd63101, 16'd16649, 16'd5488, 16'd8749, 16'd13140, 16'd62879, 16'd25754, 16'd36693, 16'd56942, 16'd3708, 16'd52836, 16'd55657});
	test_expansion(128'h516ed37d2f115635a3441ac80db51062, {16'd6793, 16'd53769, 16'd16575, 16'd52902, 16'd59473, 16'd37524, 16'd21876, 16'd37158, 16'd59689, 16'd23580, 16'd34334, 16'd41512, 16'd7466, 16'd19351, 16'd15530, 16'd23735, 16'd55465, 16'd11086, 16'd65311, 16'd63277, 16'd23994, 16'd18581, 16'd17668, 16'd38593, 16'd16985, 16'd50709});
	test_expansion(128'hc046b340bdf67315dc4761a7599a9611, {16'd42748, 16'd37152, 16'd26246, 16'd24613, 16'd37759, 16'd1190, 16'd30102, 16'd39149, 16'd7464, 16'd48244, 16'd5337, 16'd18687, 16'd19861, 16'd29986, 16'd44632, 16'd38254, 16'd47710, 16'd40911, 16'd35252, 16'd61571, 16'd27692, 16'd36060, 16'd65056, 16'd41716, 16'd855, 16'd63236});
	test_expansion(128'hc095d5343ecf25ecd8e6f712e2bfcc58, {16'd59119, 16'd26620, 16'd56521, 16'd49642, 16'd22832, 16'd18613, 16'd37470, 16'd47228, 16'd14673, 16'd22994, 16'd12969, 16'd52114, 16'd63953, 16'd15394, 16'd162, 16'd51740, 16'd18826, 16'd10081, 16'd37479, 16'd28866, 16'd36153, 16'd59551, 16'd11971, 16'd25337, 16'd49348, 16'd12548});
	test_expansion(128'h9c7537bed518ba965b96972ec77347b7, {16'd7348, 16'd6533, 16'd43913, 16'd22729, 16'd32532, 16'd14384, 16'd3129, 16'd64130, 16'd48815, 16'd4567, 16'd41779, 16'd1454, 16'd35815, 16'd34343, 16'd35585, 16'd42949, 16'd34823, 16'd39215, 16'd7006, 16'd48158, 16'd38959, 16'd16123, 16'd4930, 16'd36449, 16'd19425, 16'd27642});
	test_expansion(128'h9be14ba0289d299e010ee10f0dacd549, {16'd58964, 16'd16293, 16'd60963, 16'd33988, 16'd42922, 16'd55003, 16'd62169, 16'd23222, 16'd18794, 16'd47722, 16'd53602, 16'd51113, 16'd29222, 16'd59638, 16'd46521, 16'd16829, 16'd31086, 16'd29219, 16'd5965, 16'd25470, 16'd51622, 16'd64320, 16'd28839, 16'd50717, 16'd42294, 16'd56669});
	test_expansion(128'h2c262a52f62dfde706428cc621a4aa58, {16'd25307, 16'd38819, 16'd4085, 16'd64759, 16'd18886, 16'd51023, 16'd2104, 16'd25815, 16'd52008, 16'd44509, 16'd13238, 16'd32507, 16'd19869, 16'd56255, 16'd60859, 16'd1062, 16'd19814, 16'd51885, 16'd18255, 16'd22688, 16'd60612, 16'd52314, 16'd22839, 16'd11467, 16'd35400, 16'd34350});
	test_expansion(128'h20561c275844c35896e7a6fa6448dd6b, {16'd4289, 16'd59079, 16'd42823, 16'd1992, 16'd48277, 16'd27324, 16'd41081, 16'd12828, 16'd9109, 16'd61559, 16'd761, 16'd44377, 16'd54074, 16'd719, 16'd53245, 16'd38986, 16'd39600, 16'd30137, 16'd46871, 16'd53681, 16'd47823, 16'd33102, 16'd46471, 16'd20416, 16'd31088, 16'd29951});
	test_expansion(128'h8a53fd5aaa2af99d09a9eec38555624b, {16'd43794, 16'd62029, 16'd33675, 16'd8868, 16'd7761, 16'd58885, 16'd52564, 16'd63265, 16'd12075, 16'd3819, 16'd3117, 16'd8586, 16'd59689, 16'd15423, 16'd33437, 16'd47237, 16'd31878, 16'd49806, 16'd55929, 16'd28032, 16'd29425, 16'd25517, 16'd28161, 16'd4506, 16'd48127, 16'd47240});
	test_expansion(128'h7882425a17cf4f65610274d5a9f0bcbd, {16'd18995, 16'd12811, 16'd17607, 16'd35178, 16'd23711, 16'd44691, 16'd57241, 16'd18281, 16'd27879, 16'd51373, 16'd18874, 16'd45881, 16'd55715, 16'd36459, 16'd31231, 16'd1002, 16'd51526, 16'd49110, 16'd24372, 16'd16358, 16'd23985, 16'd8678, 16'd60294, 16'd28539, 16'd59785, 16'd65462});
	test_expansion(128'hfd7385c95cf14910fe036aaa74932f91, {16'd687, 16'd18251, 16'd29302, 16'd45875, 16'd28900, 16'd20143, 16'd27084, 16'd3924, 16'd13982, 16'd198, 16'd19282, 16'd14652, 16'd8081, 16'd46527, 16'd46556, 16'd36785, 16'd48820, 16'd62087, 16'd49251, 16'd20424, 16'd24658, 16'd44097, 16'd11459, 16'd1763, 16'd22740, 16'd48092});
	test_expansion(128'hdae4bd52da74d4a3eaff9db2b4006e6f, {16'd561, 16'd37094, 16'd11760, 16'd54536, 16'd36414, 16'd52087, 16'd37422, 16'd42729, 16'd21678, 16'd51804, 16'd48365, 16'd50469, 16'd64654, 16'd22681, 16'd8867, 16'd64184, 16'd24918, 16'd34382, 16'd45967, 16'd32983, 16'd47924, 16'd60269, 16'd29495, 16'd21756, 16'd20553, 16'd65484});
	test_expansion(128'h58cd63c873cac8b8d93e313bc94e76e3, {16'd35321, 16'd15656, 16'd16457, 16'd64746, 16'd42619, 16'd7320, 16'd48076, 16'd50567, 16'd25672, 16'd44132, 16'd61011, 16'd62780, 16'd2393, 16'd29833, 16'd31796, 16'd13999, 16'd18788, 16'd47416, 16'd56045, 16'd60190, 16'd5006, 16'd43891, 16'd6244, 16'd58289, 16'd57520, 16'd30573});
	test_expansion(128'h6b78b4ca2d14d41eaddc460378e76ed2, {16'd30315, 16'd19212, 16'd50890, 16'd59825, 16'd61180, 16'd46967, 16'd30046, 16'd56916, 16'd24890, 16'd16290, 16'd25690, 16'd20969, 16'd27703, 16'd59475, 16'd17857, 16'd36894, 16'd11664, 16'd46462, 16'd15810, 16'd57991, 16'd47279, 16'd59728, 16'd30494, 16'd29020, 16'd62380, 16'd20780});
	test_expansion(128'h97037b451c3ca2caecd87f7920bfa582, {16'd57795, 16'd17500, 16'd13231, 16'd13075, 16'd58658, 16'd62649, 16'd26031, 16'd62492, 16'd205, 16'd7194, 16'd48777, 16'd54790, 16'd56728, 16'd9775, 16'd18489, 16'd61679, 16'd50777, 16'd15970, 16'd62664, 16'd45091, 16'd35147, 16'd45808, 16'd6218, 16'd61696, 16'd18883, 16'd58888});
	test_expansion(128'h3b654899f102aab3b26d7d211748bdef, {16'd4973, 16'd2372, 16'd41494, 16'd58568, 16'd50537, 16'd50438, 16'd3054, 16'd23998, 16'd47076, 16'd30062, 16'd65017, 16'd64786, 16'd53492, 16'd59687, 16'd64573, 16'd41698, 16'd14045, 16'd13425, 16'd38675, 16'd32732, 16'd3292, 16'd3962, 16'd59434, 16'd11842, 16'd48931, 16'd47197});
	test_expansion(128'hfb2db411fe3671b73131db2dc932427d, {16'd37570, 16'd7520, 16'd4036, 16'd48885, 16'd39769, 16'd44737, 16'd62041, 16'd26207, 16'd11025, 16'd13162, 16'd5260, 16'd62894, 16'd46292, 16'd54639, 16'd63862, 16'd61829, 16'd45650, 16'd41839, 16'd9823, 16'd38547, 16'd17774, 16'd18263, 16'd8214, 16'd24742, 16'd25829, 16'd1382});
	test_expansion(128'hb3a5fda482941f64fb0046f5c3f74534, {16'd43047, 16'd13169, 16'd46954, 16'd55630, 16'd34366, 16'd15604, 16'd5706, 16'd1211, 16'd36460, 16'd36861, 16'd55773, 16'd24318, 16'd63536, 16'd60958, 16'd64384, 16'd25348, 16'd38466, 16'd61188, 16'd57233, 16'd40832, 16'd8507, 16'd52677, 16'd50802, 16'd49511, 16'd29091, 16'd60521});
	test_expansion(128'h325345cc006aceffa0966555c51efc09, {16'd40121, 16'd25120, 16'd7548, 16'd50705, 16'd50206, 16'd6192, 16'd11037, 16'd20693, 16'd21751, 16'd55883, 16'd13164, 16'd3996, 16'd46541, 16'd39453, 16'd32946, 16'd42589, 16'd39485, 16'd37830, 16'd61704, 16'd13586, 16'd28183, 16'd38246, 16'd60830, 16'd65075, 16'd14958, 16'd35790});
	test_expansion(128'hb27bb0e332a773c309d309fc2b2a4eff, {16'd4363, 16'd36449, 16'd4828, 16'd27937, 16'd12252, 16'd21658, 16'd42213, 16'd32986, 16'd17714, 16'd63610, 16'd1467, 16'd37998, 16'd38028, 16'd6322, 16'd53711, 16'd25916, 16'd500, 16'd21843, 16'd2745, 16'd23829, 16'd23642, 16'd22398, 16'd57777, 16'd37484, 16'd35017, 16'd54082});
	test_expansion(128'h564c8d03fed53313e4d492cf8044b01b, {16'd39739, 16'd29211, 16'd4149, 16'd27215, 16'd42091, 16'd25131, 16'd11961, 16'd20920, 16'd38165, 16'd33545, 16'd27998, 16'd23668, 16'd27174, 16'd41900, 16'd44008, 16'd19892, 16'd51227, 16'd10779, 16'd21243, 16'd18573, 16'd15124, 16'd2117, 16'd65132, 16'd51981, 16'd50482, 16'd6886});
	test_expansion(128'h7956d180c91b22b8bfc3d12dbb505077, {16'd15689, 16'd25194, 16'd14246, 16'd27241, 16'd9054, 16'd38461, 16'd65416, 16'd32743, 16'd51414, 16'd5625, 16'd24972, 16'd33767, 16'd35648, 16'd16331, 16'd44629, 16'd49194, 16'd11132, 16'd56200, 16'd20070, 16'd6870, 16'd8861, 16'd31004, 16'd49150, 16'd25172, 16'd26265, 16'd31558});
	test_expansion(128'h6c4a37ee11b22943f8b0f524e43f84ed, {16'd42599, 16'd14780, 16'd60376, 16'd24208, 16'd33236, 16'd42230, 16'd23330, 16'd64148, 16'd56300, 16'd50334, 16'd12935, 16'd18743, 16'd31780, 16'd63440, 16'd34730, 16'd27786, 16'd62686, 16'd36976, 16'd24729, 16'd50598, 16'd61274, 16'd17180, 16'd48530, 16'd25825, 16'd23270, 16'd30891});
	test_expansion(128'hec74da69cd01fabc003f19ad4d18bafa, {16'd21432, 16'd60786, 16'd45063, 16'd26373, 16'd41065, 16'd36511, 16'd64566, 16'd19031, 16'd23904, 16'd24970, 16'd12969, 16'd34858, 16'd60969, 16'd25062, 16'd53502, 16'd44375, 16'd63843, 16'd60632, 16'd33126, 16'd48881, 16'd14438, 16'd42361, 16'd57891, 16'd3640, 16'd30563, 16'd4169});
	test_expansion(128'h2379aca7d4b08aac26009b58157fef65, {16'd28641, 16'd17445, 16'd23686, 16'd15364, 16'd28111, 16'd54688, 16'd11876, 16'd49290, 16'd33503, 16'd58238, 16'd488, 16'd29391, 16'd42568, 16'd21817, 16'd6777, 16'd36467, 16'd62211, 16'd32133, 16'd2555, 16'd38954, 16'd27664, 16'd6789, 16'd21639, 16'd39884, 16'd7717, 16'd10283});
	test_expansion(128'h6664db6ede8128e7c3060013badde080, {16'd402, 16'd34527, 16'd36075, 16'd59258, 16'd21551, 16'd46496, 16'd7726, 16'd35776, 16'd14205, 16'd37256, 16'd29513, 16'd25521, 16'd27989, 16'd40182, 16'd31537, 16'd55162, 16'd11551, 16'd6885, 16'd37453, 16'd1668, 16'd62709, 16'd43590, 16'd35060, 16'd42998, 16'd55416, 16'd32159});
	test_expansion(128'h052f6522d679aacea90db55984e96ce5, {16'd14966, 16'd51153, 16'd51501, 16'd24804, 16'd4147, 16'd64160, 16'd4479, 16'd12263, 16'd46100, 16'd32278, 16'd44843, 16'd62596, 16'd33902, 16'd2937, 16'd216, 16'd40041, 16'd65024, 16'd15535, 16'd53775, 16'd7262, 16'd20143, 16'd8882, 16'd25148, 16'd29833, 16'd24279, 16'd47594});
	test_expansion(128'ha570fd960d717332274b6ced26020a35, {16'd38029, 16'd61133, 16'd4629, 16'd12470, 16'd16243, 16'd62591, 16'd49931, 16'd63606, 16'd13645, 16'd7832, 16'd10697, 16'd8775, 16'd43552, 16'd6734, 16'd48706, 16'd43592, 16'd4898, 16'd34224, 16'd4776, 16'd30268, 16'd24582, 16'd48792, 16'd65257, 16'd50051, 16'd34068, 16'd5435});
	test_expansion(128'h7e1d9a53818ce226ae6ed7d71cf43536, {16'd57453, 16'd9777, 16'd28155, 16'd40407, 16'd41182, 16'd65497, 16'd16647, 16'd60609, 16'd18741, 16'd37904, 16'd46668, 16'd5393, 16'd5799, 16'd60426, 16'd51808, 16'd62649, 16'd11362, 16'd2670, 16'd28926, 16'd24924, 16'd18701, 16'd64392, 16'd55999, 16'd9635, 16'd45356, 16'd30053});
	test_expansion(128'he1ac28cfbdd3af4a7da23ff23609d0a7, {16'd36315, 16'd60670, 16'd28844, 16'd45388, 16'd23575, 16'd28866, 16'd51174, 16'd48990, 16'd63256, 16'd39980, 16'd55438, 16'd29003, 16'd39330, 16'd1787, 16'd34902, 16'd46167, 16'd32220, 16'd24452, 16'd9737, 16'd662, 16'd27661, 16'd43523, 16'd56767, 16'd55556, 16'd33439, 16'd622});
	test_expansion(128'h68b6abd6a5696898a3d9c7e795ecba02, {16'd55372, 16'd36108, 16'd44279, 16'd58342, 16'd42497, 16'd57259, 16'd13449, 16'd28110, 16'd46518, 16'd46799, 16'd3434, 16'd64052, 16'd12394, 16'd49546, 16'd34949, 16'd6409, 16'd56953, 16'd8748, 16'd33955, 16'd38404, 16'd42174, 16'd5546, 16'd7637, 16'd45431, 16'd28264, 16'd36905});
	test_expansion(128'h21bf698eecdf5368321cb2f0dd90efba, {16'd19347, 16'd52475, 16'd32530, 16'd56573, 16'd28256, 16'd43488, 16'd41533, 16'd3846, 16'd35037, 16'd44887, 16'd9265, 16'd39860, 16'd39511, 16'd12180, 16'd13554, 16'd59252, 16'd2082, 16'd56664, 16'd43942, 16'd33592, 16'd57622, 16'd46386, 16'd19124, 16'd42380, 16'd59430, 16'd60266});
	test_expansion(128'h1d549d17464200991ce6462529e55a9b, {16'd49810, 16'd29251, 16'd52332, 16'd46631, 16'd19651, 16'd25079, 16'd42963, 16'd62609, 16'd14961, 16'd27013, 16'd44997, 16'd16923, 16'd49678, 16'd12959, 16'd2837, 16'd31024, 16'd36750, 16'd38663, 16'd26676, 16'd1039, 16'd17943, 16'd32014, 16'd27944, 16'd18557, 16'd49342, 16'd5931});
	test_expansion(128'hcdda6ef32a25dc3ce41e0c6576b2cebe, {16'd10446, 16'd24704, 16'd59705, 16'd13982, 16'd14839, 16'd60488, 16'd23537, 16'd65154, 16'd36501, 16'd61785, 16'd46893, 16'd1360, 16'd52039, 16'd7539, 16'd18948, 16'd15024, 16'd24014, 16'd49314, 16'd16247, 16'd29200, 16'd9861, 16'd17841, 16'd17614, 16'd51481, 16'd61662, 16'd37251});
	test_expansion(128'hec78870269175f8bf0531d7bd2878c4c, {16'd52088, 16'd61417, 16'd27258, 16'd12322, 16'd53190, 16'd16044, 16'd40368, 16'd54945, 16'd29924, 16'd59615, 16'd23718, 16'd54157, 16'd50518, 16'd24386, 16'd50181, 16'd58020, 16'd53954, 16'd60758, 16'd10996, 16'd64108, 16'd21174, 16'd64894, 16'd20165, 16'd14560, 16'd16150, 16'd46382});
	test_expansion(128'h35696dcc889a893c765eb82ee60ca16e, {16'd55304, 16'd11131, 16'd28548, 16'd16011, 16'd29279, 16'd53896, 16'd57998, 16'd40363, 16'd7146, 16'd26706, 16'd42607, 16'd56735, 16'd40375, 16'd48469, 16'd47452, 16'd27542, 16'd27827, 16'd3487, 16'd29728, 16'd56683, 16'd8478, 16'd61777, 16'd48568, 16'd29135, 16'd35879, 16'd10258});
	test_expansion(128'h84a3de5fe0eb903f9a283649ac499463, {16'd42744, 16'd20128, 16'd22374, 16'd38153, 16'd47701, 16'd55358, 16'd49485, 16'd45921, 16'd50021, 16'd30534, 16'd8178, 16'd8292, 16'd45641, 16'd29057, 16'd36519, 16'd62098, 16'd47548, 16'd4733, 16'd59033, 16'd5339, 16'd4999, 16'd27394, 16'd8533, 16'd8984, 16'd3112, 16'd14814});
	test_expansion(128'h29daf74ebf8e18219e5c7fb535da1f56, {16'd16426, 16'd60238, 16'd21546, 16'd48633, 16'd5093, 16'd34237, 16'd49922, 16'd63246, 16'd54550, 16'd41047, 16'd21504, 16'd63051, 16'd2474, 16'd49852, 16'd41161, 16'd25378, 16'd9910, 16'd33981, 16'd25346, 16'd25548, 16'd40617, 16'd17066, 16'd43342, 16'd39886, 16'd16370, 16'd5847});
	test_expansion(128'h7dd7d1467c4744305c35e0eb411db6c1, {16'd35562, 16'd26575, 16'd29800, 16'd57666, 16'd10163, 16'd40147, 16'd62240, 16'd39414, 16'd46725, 16'd56960, 16'd50018, 16'd18564, 16'd18387, 16'd42158, 16'd48551, 16'd29241, 16'd23770, 16'd28689, 16'd17822, 16'd37632, 16'd36160, 16'd41571, 16'd26349, 16'd33104, 16'd48182, 16'd2833});
	test_expansion(128'h1ac22a6a36fb958ce4ff3f5c60f928b0, {16'd55589, 16'd36480, 16'd17796, 16'd33675, 16'd63206, 16'd24023, 16'd40959, 16'd22905, 16'd16032, 16'd54191, 16'd16163, 16'd54836, 16'd14003, 16'd34467, 16'd8179, 16'd48945, 16'd20423, 16'd45544, 16'd40190, 16'd56278, 16'd42607, 16'd22235, 16'd8894, 16'd371, 16'd17072, 16'd37708});
	test_expansion(128'h318cb780ef16cab4f1c3ff6a7172ad67, {16'd32868, 16'd41139, 16'd37321, 16'd43369, 16'd38854, 16'd51689, 16'd21886, 16'd40992, 16'd48173, 16'd53483, 16'd19543, 16'd9430, 16'd11967, 16'd28279, 16'd8055, 16'd5915, 16'd16095, 16'd34020, 16'd50321, 16'd12461, 16'd46128, 16'd63675, 16'd7285, 16'd4521, 16'd63096, 16'd57192});
	test_expansion(128'h113114d742e508b912f9bf418260a026, {16'd27178, 16'd19772, 16'd45634, 16'd61707, 16'd64338, 16'd2797, 16'd37558, 16'd32192, 16'd4754, 16'd1355, 16'd24375, 16'd28147, 16'd48689, 16'd5307, 16'd188, 16'd48559, 16'd49959, 16'd37059, 16'd25910, 16'd8708, 16'd34392, 16'd27136, 16'd460, 16'd35677, 16'd7548, 16'd60177});
	test_expansion(128'hd2fbabe6d6b63ba5694a4c172d0f4cff, {16'd30, 16'd32188, 16'd61766, 16'd37730, 16'd48898, 16'd45865, 16'd30317, 16'd38765, 16'd63759, 16'd9719, 16'd5294, 16'd61207, 16'd50126, 16'd22000, 16'd17954, 16'd55984, 16'd39605, 16'd52530, 16'd15313, 16'd27175, 16'd35458, 16'd37733, 16'd44207, 16'd55152, 16'd15205, 16'd42344});
	test_expansion(128'h309236837d29228bc2888aee51d2d4a7, {16'd43263, 16'd35942, 16'd33686, 16'd23992, 16'd13283, 16'd32951, 16'd41342, 16'd9748, 16'd9487, 16'd52648, 16'd27160, 16'd10767, 16'd12241, 16'd43764, 16'd40100, 16'd28724, 16'd57968, 16'd44449, 16'd22845, 16'd39888, 16'd48898, 16'd10713, 16'd54178, 16'd4628, 16'd30646, 16'd49188});
	test_expansion(128'h4f7a29ee8a9fbd6653fae9261b18ed43, {16'd52766, 16'd11228, 16'd64052, 16'd11631, 16'd49929, 16'd18359, 16'd6452, 16'd50314, 16'd12625, 16'd48137, 16'd42384, 16'd27666, 16'd13974, 16'd60424, 16'd5554, 16'd43804, 16'd24010, 16'd32979, 16'd57558, 16'd18532, 16'd4372, 16'd46015, 16'd37047, 16'd12720, 16'd65270, 16'd60252});
	test_expansion(128'hfda7099f7b81e67a70293ad7a8ec5329, {16'd20489, 16'd9620, 16'd6466, 16'd28051, 16'd12749, 16'd38082, 16'd6872, 16'd17322, 16'd24523, 16'd51806, 16'd4792, 16'd24423, 16'd59734, 16'd32282, 16'd16334, 16'd40997, 16'd19493, 16'd44286, 16'd15344, 16'd49291, 16'd14916, 16'd4462, 16'd1955, 16'd30002, 16'd37777, 16'd19243});
	test_expansion(128'h6f3e439a828f974ce5152eac88398184, {16'd17871, 16'd64791, 16'd42500, 16'd47316, 16'd6588, 16'd33865, 16'd21711, 16'd7736, 16'd30733, 16'd13899, 16'd17954, 16'd45036, 16'd51624, 16'd25776, 16'd25665, 16'd4596, 16'd41240, 16'd9515, 16'd8032, 16'd19181, 16'd62054, 16'd30494, 16'd2161, 16'd35530, 16'd28833, 16'd30145});
	test_expansion(128'h09dc98caa80a9b9a0f36a7c4768b4d5d, {16'd15354, 16'd31086, 16'd54424, 16'd22678, 16'd33029, 16'd43036, 16'd6492, 16'd27060, 16'd31361, 16'd1253, 16'd8496, 16'd44082, 16'd22801, 16'd26824, 16'd56718, 16'd12788, 16'd57663, 16'd62258, 16'd46323, 16'd27711, 16'd59047, 16'd63457, 16'd57002, 16'd62543, 16'd52260, 16'd9711});
	test_expansion(128'h4dad73918a6b072f595a8a56a2c621f3, {16'd44045, 16'd30158, 16'd32832, 16'd20778, 16'd58877, 16'd12492, 16'd49499, 16'd56703, 16'd19516, 16'd17199, 16'd4606, 16'd17313, 16'd20171, 16'd18151, 16'd56198, 16'd42587, 16'd8820, 16'd21335, 16'd52224, 16'd18900, 16'd5053, 16'd23671, 16'd64089, 16'd8985, 16'd31208, 16'd10645});
	test_expansion(128'h06a77b1773334d7f536db1e960b208bb, {16'd61156, 16'd3610, 16'd45893, 16'd45113, 16'd22167, 16'd42648, 16'd57961, 16'd40986, 16'd52839, 16'd4705, 16'd60431, 16'd9848, 16'd12660, 16'd7095, 16'd32635, 16'd45545, 16'd35274, 16'd51404, 16'd63842, 16'd43938, 16'd17411, 16'd9664, 16'd51464, 16'd6842, 16'd48010, 16'd9829});
	test_expansion(128'h3a274b0cb49d67f2ca165c15ed42630a, {16'd59794, 16'd9486, 16'd4468, 16'd22991, 16'd46590, 16'd28692, 16'd9241, 16'd37471, 16'd50327, 16'd51786, 16'd5034, 16'd46666, 16'd37635, 16'd9592, 16'd43566, 16'd36751, 16'd35484, 16'd18808, 16'd46715, 16'd60339, 16'd30220, 16'd6788, 16'd9715, 16'd51160, 16'd65271, 16'd4023});
	test_expansion(128'h4a06fffdbb3c72c30db2319464023e32, {16'd39250, 16'd6926, 16'd35621, 16'd56292, 16'd7870, 16'd15255, 16'd11294, 16'd31684, 16'd2314, 16'd59318, 16'd61084, 16'd35184, 16'd53777, 16'd17867, 16'd18827, 16'd58115, 16'd11577, 16'd43832, 16'd35817, 16'd8552, 16'd15092, 16'd57777, 16'd50343, 16'd27434, 16'd12955, 16'd33670});
	test_expansion(128'hdab78940a8a3a3353a51c5ccf95336ae, {16'd3131, 16'd39162, 16'd64118, 16'd12936, 16'd56671, 16'd58359, 16'd49229, 16'd4846, 16'd41081, 16'd14144, 16'd23821, 16'd13425, 16'd23439, 16'd50717, 16'd56745, 16'd61040, 16'd23862, 16'd45316, 16'd26493, 16'd54989, 16'd11683, 16'd22746, 16'd52925, 16'd5447, 16'd34082, 16'd56964});
	test_expansion(128'h6babccb58230dab6644d891b6be591aa, {16'd63279, 16'd21763, 16'd27493, 16'd64850, 16'd8794, 16'd42073, 16'd47936, 16'd60695, 16'd9750, 16'd56168, 16'd14729, 16'd25858, 16'd49402, 16'd34759, 16'd20401, 16'd65296, 16'd17154, 16'd8120, 16'd32219, 16'd17644, 16'd23623, 16'd47667, 16'd51567, 16'd9043, 16'd6332, 16'd2425});
	test_expansion(128'hdb5c45d2480342fbb69e0c50deb3514d, {16'd20438, 16'd60662, 16'd45857, 16'd214, 16'd36734, 16'd45197, 16'd57943, 16'd52519, 16'd26680, 16'd12613, 16'd36817, 16'd41864, 16'd42521, 16'd31248, 16'd53837, 16'd16591, 16'd15404, 16'd15264, 16'd29378, 16'd15824, 16'd30225, 16'd34290, 16'd15713, 16'd12397, 16'd1676, 16'd19759});
	test_expansion(128'h764755f5a303b894e27aec26c3e226fe, {16'd62783, 16'd65252, 16'd46879, 16'd23880, 16'd41311, 16'd16203, 16'd48262, 16'd22323, 16'd21583, 16'd45983, 16'd27041, 16'd33730, 16'd35533, 16'd16924, 16'd23597, 16'd48045, 16'd46439, 16'd63970, 16'd52100, 16'd18396, 16'd5718, 16'd33690, 16'd7498, 16'd41199, 16'd23102, 16'd23999});
	test_expansion(128'h51f2f6114ae18029b0b38d3b5a34a5b5, {16'd60397, 16'd43109, 16'd52399, 16'd55854, 16'd1458, 16'd51183, 16'd43618, 16'd43795, 16'd27102, 16'd60327, 16'd61688, 16'd13811, 16'd62606, 16'd17455, 16'd17435, 16'd50120, 16'd28156, 16'd10950, 16'd25562, 16'd9076, 16'd15599, 16'd2391, 16'd63235, 16'd19962, 16'd56514, 16'd40803});
	test_expansion(128'h739b91088b3fc53ab6d8206a771bb792, {16'd55190, 16'd40341, 16'd25155, 16'd26626, 16'd48336, 16'd53562, 16'd12320, 16'd19880, 16'd19307, 16'd35940, 16'd33016, 16'd8743, 16'd37501, 16'd40017, 16'd41730, 16'd2309, 16'd64592, 16'd2137, 16'd17579, 16'd61619, 16'd47978, 16'd36016, 16'd8935, 16'd51307, 16'd34964, 16'd3065});
	test_expansion(128'h2894a42ecbf35f908620b164fe7178fd, {16'd19338, 16'd52898, 16'd26129, 16'd17947, 16'd49975, 16'd41449, 16'd33113, 16'd2369, 16'd56801, 16'd48863, 16'd3252, 16'd6490, 16'd15106, 16'd54184, 16'd56389, 16'd31887, 16'd53110, 16'd29747, 16'd25429, 16'd20616, 16'd18456, 16'd40507, 16'd11681, 16'd522, 16'd25690, 16'd8914});
	test_expansion(128'h058b778357ece0b23a041e97d7a30915, {16'd23531, 16'd7135, 16'd26657, 16'd51270, 16'd63092, 16'd45724, 16'd15314, 16'd24251, 16'd51671, 16'd11213, 16'd34202, 16'd15921, 16'd19691, 16'd61743, 16'd6912, 16'd29212, 16'd34630, 16'd6793, 16'd10423, 16'd44649, 16'd52916, 16'd24872, 16'd27039, 16'd34977, 16'd64335, 16'd5763});
	test_expansion(128'h5c752fcacbcf799e5c8696550be8f4da, {16'd47819, 16'd25104, 16'd32064, 16'd48808, 16'd27361, 16'd57631, 16'd33630, 16'd20643, 16'd50996, 16'd7986, 16'd5955, 16'd47309, 16'd19324, 16'd11931, 16'd57640, 16'd7185, 16'd8294, 16'd33084, 16'd12682, 16'd45928, 16'd1324, 16'd3367, 16'd32824, 16'd49584, 16'd22395, 16'd62887});
	test_expansion(128'hcfb4a178dc770aa65dc0a09caeeef216, {16'd50183, 16'd20942, 16'd16062, 16'd39846, 16'd11732, 16'd35333, 16'd32218, 16'd50606, 16'd23408, 16'd7257, 16'd1424, 16'd16182, 16'd49344, 16'd64167, 16'd37199, 16'd5219, 16'd27624, 16'd64380, 16'd59239, 16'd52231, 16'd54261, 16'd22344, 16'd427, 16'd22473, 16'd21261, 16'd52040});
	test_expansion(128'hce2b0496e958092c351411a6d204be35, {16'd63128, 16'd20589, 16'd33758, 16'd51585, 16'd55264, 16'd59596, 16'd21966, 16'd7241, 16'd64206, 16'd32021, 16'd48492, 16'd64879, 16'd41200, 16'd17174, 16'd40537, 16'd4733, 16'd52450, 16'd52615, 16'd48567, 16'd50634, 16'd50845, 16'd63558, 16'd16021, 16'd15099, 16'd59491, 16'd19050});
	test_expansion(128'h59f0086f109250a9ea1ed6b29d717ac6, {16'd58975, 16'd27579, 16'd6289, 16'd23943, 16'd39102, 16'd41191, 16'd19955, 16'd26169, 16'd63108, 16'd47643, 16'd29498, 16'd6469, 16'd57245, 16'd47414, 16'd3494, 16'd63798, 16'd58763, 16'd41666, 16'd64291, 16'd5059, 16'd57606, 16'd42989, 16'd19990, 16'd12122, 16'd3787, 16'd14222});
	test_expansion(128'hb926dab0a983e7e190c7a26718f40629, {16'd32194, 16'd18963, 16'd41697, 16'd43277, 16'd7829, 16'd48550, 16'd63645, 16'd20345, 16'd707, 16'd49945, 16'd37505, 16'd52540, 16'd23946, 16'd29501, 16'd14767, 16'd10086, 16'd498, 16'd54182, 16'd50037, 16'd32812, 16'd5085, 16'd38654, 16'd32624, 16'd18492, 16'd10641, 16'd29283});
	test_expansion(128'h496aef89cecc14f28d457cc2e8305626, {16'd99, 16'd17683, 16'd34174, 16'd34762, 16'd36617, 16'd26257, 16'd23473, 16'd30556, 16'd6536, 16'd36336, 16'd49185, 16'd17058, 16'd65388, 16'd22222, 16'd46967, 16'd1087, 16'd28943, 16'd48218, 16'd12815, 16'd13803, 16'd22176, 16'd60032, 16'd59346, 16'd43060, 16'd17372, 16'd17338});
	test_expansion(128'h5cb6db5f41b93ea64c8aa8cb95680974, {16'd7106, 16'd36784, 16'd60111, 16'd7798, 16'd20077, 16'd62028, 16'd38309, 16'd43589, 16'd5379, 16'd9573, 16'd18276, 16'd2217, 16'd44533, 16'd33165, 16'd22350, 16'd45700, 16'd14382, 16'd44884, 16'd37814, 16'd40105, 16'd3201, 16'd26066, 16'd27983, 16'd45015, 16'd33751, 16'd3222});
	test_expansion(128'he4ce05d03eb7640b389bc1b42b1bb813, {16'd30289, 16'd61034, 16'd37757, 16'd7972, 16'd45896, 16'd35609, 16'd61442, 16'd20287, 16'd22921, 16'd40939, 16'd40621, 16'd38562, 16'd22508, 16'd54827, 16'd64874, 16'd30627, 16'd39342, 16'd54357, 16'd48071, 16'd5124, 16'd32001, 16'd12392, 16'd32896, 16'd22000, 16'd54414, 16'd52075});
	test_expansion(128'hc341857a5aff5fe3f9ebd605095aefba, {16'd36028, 16'd53857, 16'd8917, 16'd59489, 16'd32987, 16'd8710, 16'd25931, 16'd8011, 16'd54296, 16'd50997, 16'd54036, 16'd11476, 16'd678, 16'd23990, 16'd60993, 16'd27968, 16'd56933, 16'd11027, 16'd60719, 16'd64156, 16'd6586, 16'd16596, 16'd42965, 16'd4985, 16'd54366, 16'd3383});
	test_expansion(128'h2f273396ed3efc3a373ad44eab21794a, {16'd4217, 16'd47592, 16'd5199, 16'd32094, 16'd41002, 16'd3532, 16'd38292, 16'd27283, 16'd22944, 16'd27629, 16'd28907, 16'd61924, 16'd27493, 16'd13568, 16'd29537, 16'd59362, 16'd8410, 16'd50823, 16'd45236, 16'd17587, 16'd12339, 16'd64205, 16'd62105, 16'd30826, 16'd33799, 16'd33398});
	test_expansion(128'h424ab97214f77450e656324698b3c29c, {16'd47723, 16'd26532, 16'd14487, 16'd20921, 16'd10789, 16'd37956, 16'd45888, 16'd19670, 16'd15831, 16'd48971, 16'd41729, 16'd15052, 16'd48452, 16'd38729, 16'd12997, 16'd2290, 16'd32308, 16'd53921, 16'd11982, 16'd50407, 16'd34580, 16'd56839, 16'd47990, 16'd1108, 16'd22102, 16'd49048});
	test_expansion(128'hee180c6917f29775dfd95c45f6f69a19, {16'd57638, 16'd57294, 16'd30968, 16'd20518, 16'd13047, 16'd2256, 16'd6882, 16'd60079, 16'd40620, 16'd40717, 16'd63503, 16'd50032, 16'd2549, 16'd50230, 16'd22425, 16'd37523, 16'd34421, 16'd39214, 16'd42581, 16'd41061, 16'd29479, 16'd6289, 16'd9152, 16'd23580, 16'd37427, 16'd52258});
	test_expansion(128'h81022308e8c1546310d4896f1983f6bb, {16'd56161, 16'd16281, 16'd3143, 16'd29591, 16'd12657, 16'd35722, 16'd23553, 16'd49371, 16'd13891, 16'd52269, 16'd39943, 16'd17277, 16'd54949, 16'd25575, 16'd21684, 16'd48498, 16'd65099, 16'd39003, 16'd10955, 16'd36456, 16'd54559, 16'd54082, 16'd54526, 16'd5160, 16'd15248, 16'd17684});
	test_expansion(128'hde5d8fa05f1a653d0195fc59c312bb0f, {16'd65222, 16'd21584, 16'd42587, 16'd32581, 16'd9058, 16'd4202, 16'd36626, 16'd3356, 16'd60271, 16'd31352, 16'd2117, 16'd23486, 16'd55950, 16'd30870, 16'd36735, 16'd17371, 16'd45749, 16'd55650, 16'd21706, 16'd15531, 16'd4830, 16'd60392, 16'd5052, 16'd36555, 16'd11963, 16'd1636});
	test_expansion(128'h05cba974ed307f7a78cb117abac8d403, {16'd34865, 16'd43016, 16'd51450, 16'd39687, 16'd32832, 16'd56407, 16'd23792, 16'd18185, 16'd34275, 16'd25332, 16'd37203, 16'd17319, 16'd9903, 16'd16798, 16'd21935, 16'd4021, 16'd64509, 16'd12148, 16'd47192, 16'd31120, 16'd11839, 16'd39179, 16'd56474, 16'd17657, 16'd11417, 16'd12628});
	test_expansion(128'heec3479bfb3cf55fdb187e233b0f7326, {16'd36717, 16'd20304, 16'd28616, 16'd49269, 16'd9201, 16'd33221, 16'd16442, 16'd19769, 16'd46275, 16'd1544, 16'd42733, 16'd736, 16'd46387, 16'd29752, 16'd52222, 16'd25094, 16'd1171, 16'd48721, 16'd34926, 16'd15392, 16'd22092, 16'd34525, 16'd46463, 16'd53929, 16'd45487, 16'd28248});
	test_expansion(128'h284b138b181fa77a2236b86e3925833e, {16'd45698, 16'd12282, 16'd60557, 16'd59496, 16'd49380, 16'd61058, 16'd55464, 16'd3621, 16'd54225, 16'd39484, 16'd36161, 16'd55087, 16'd19281, 16'd58076, 16'd52597, 16'd3377, 16'd58677, 16'd14218, 16'd63365, 16'd661, 16'd14804, 16'd28341, 16'd61973, 16'd15372, 16'd1738, 16'd56642});
	test_expansion(128'hb0ebcf318916a74ac319dd18e0372510, {16'd20051, 16'd20355, 16'd27823, 16'd61295, 16'd62219, 16'd62543, 16'd3815, 16'd24897, 16'd36959, 16'd16009, 16'd23672, 16'd33310, 16'd62535, 16'd29141, 16'd36730, 16'd62041, 16'd38287, 16'd14904, 16'd47217, 16'd31373, 16'd28709, 16'd62018, 16'd30841, 16'd64662, 16'd24387, 16'd39324});
	test_expansion(128'h487e80221e30602b5404dae20d9d846d, {16'd48724, 16'd37946, 16'd42169, 16'd57168, 16'd38934, 16'd50243, 16'd62854, 16'd39971, 16'd39224, 16'd46499, 16'd17462, 16'd5163, 16'd45487, 16'd53256, 16'd25643, 16'd11670, 16'd21806, 16'd42951, 16'd22746, 16'd42821, 16'd7965, 16'd9103, 16'd30321, 16'd17829, 16'd14589, 16'd36920});
	test_expansion(128'he72300d07e6d27909c43a9a3921acfb0, {16'd48680, 16'd9065, 16'd45425, 16'd56421, 16'd32934, 16'd7247, 16'd36502, 16'd59112, 16'd41813, 16'd63782, 16'd2239, 16'd8117, 16'd3838, 16'd38797, 16'd15245, 16'd45635, 16'd13908, 16'd32434, 16'd5519, 16'd48773, 16'd51375, 16'd14284, 16'd53192, 16'd17101, 16'd38930, 16'd30002});
	test_expansion(128'h957352a10e0a8d432b59095a5c0c48d8, {16'd37763, 16'd57383, 16'd3495, 16'd44298, 16'd613, 16'd16137, 16'd64629, 16'd60212, 16'd58285, 16'd17329, 16'd11801, 16'd43919, 16'd30064, 16'd45817, 16'd31128, 16'd37557, 16'd29417, 16'd65149, 16'd5705, 16'd64807, 16'd62237, 16'd3393, 16'd21862, 16'd21089, 16'd59961, 16'd31499});
	test_expansion(128'h68b3967a2203714c12c2049331842c3a, {16'd9809, 16'd60477, 16'd274, 16'd34912, 16'd8717, 16'd31022, 16'd55459, 16'd35654, 16'd34992, 16'd37383, 16'd63774, 16'd43020, 16'd14450, 16'd20905, 16'd36683, 16'd20866, 16'd62428, 16'd22289, 16'd46054, 16'd35892, 16'd22152, 16'd4047, 16'd4994, 16'd62876, 16'd17550, 16'd56827});
	test_expansion(128'hfcf8e61a931d4d5bff99a4b2afbeb82f, {16'd10906, 16'd37113, 16'd25745, 16'd44703, 16'd6665, 16'd4293, 16'd2513, 16'd3412, 16'd53185, 16'd9011, 16'd8151, 16'd45439, 16'd6186, 16'd42016, 16'd24327, 16'd47737, 16'd58875, 16'd21131, 16'd61805, 16'd23193, 16'd57069, 16'd58769, 16'd42625, 16'd35473, 16'd54460, 16'd39411});
	test_expansion(128'hc57f3e642010a91cb1792b5a846cd8b5, {16'd20534, 16'd36832, 16'd24399, 16'd13265, 16'd9879, 16'd45470, 16'd3257, 16'd12439, 16'd37323, 16'd51078, 16'd42699, 16'd44843, 16'd13012, 16'd29972, 16'd44981, 16'd60140, 16'd41379, 16'd42354, 16'd25504, 16'd23158, 16'd265, 16'd25389, 16'd47928, 16'd12943, 16'd57532, 16'd31390});
	test_expansion(128'hc2d00a4326707e1e1ff6177431ee4252, {16'd3727, 16'd16514, 16'd59103, 16'd59682, 16'd41949, 16'd4942, 16'd30233, 16'd17247, 16'd4279, 16'd25689, 16'd9405, 16'd44021, 16'd28147, 16'd48466, 16'd33268, 16'd63060, 16'd52642, 16'd10375, 16'd63864, 16'd48842, 16'd14778, 16'd19307, 16'd20757, 16'd3992, 16'd17553, 16'd34011});
	test_expansion(128'h63a3b6cb02e81df886f43c61a483813c, {16'd50750, 16'd22963, 16'd3036, 16'd49525, 16'd20518, 16'd14425, 16'd29655, 16'd35657, 16'd41325, 16'd54855, 16'd18669, 16'd57399, 16'd47438, 16'd59143, 16'd36324, 16'd65224, 16'd23348, 16'd56194, 16'd23004, 16'd53502, 16'd10797, 16'd39539, 16'd5576, 16'd18010, 16'd8780, 16'd32206});
	test_expansion(128'hff3a4d866d5c9ce5edad74ef5a464365, {16'd25634, 16'd12540, 16'd39471, 16'd46128, 16'd55091, 16'd58990, 16'd32044, 16'd16648, 16'd9795, 16'd10678, 16'd18407, 16'd34300, 16'd5004, 16'd20599, 16'd1696, 16'd31589, 16'd7684, 16'd64000, 16'd5614, 16'd49216, 16'd9521, 16'd41959, 16'd63604, 16'd31590, 16'd48874, 16'd13227});
	test_expansion(128'h15f1149961b91b0ef7cb7ecaddb7a133, {16'd61327, 16'd20161, 16'd20495, 16'd37726, 16'd27399, 16'd63611, 16'd58814, 16'd65424, 16'd60059, 16'd60019, 16'd61184, 16'd29784, 16'd42772, 16'd27024, 16'd44849, 16'd9185, 16'd582, 16'd40415, 16'd5739, 16'd31291, 16'd23849, 16'd1016, 16'd50131, 16'd28693, 16'd34362, 16'd58554});
	test_expansion(128'hd928cd9a19c62aa7eeca004befc16fee, {16'd42206, 16'd64478, 16'd11560, 16'd25716, 16'd25016, 16'd32217, 16'd35769, 16'd12447, 16'd60265, 16'd16591, 16'd13669, 16'd38343, 16'd49157, 16'd18793, 16'd49854, 16'd2143, 16'd46947, 16'd49023, 16'd49805, 16'd59200, 16'd29961, 16'd50561, 16'd58234, 16'd10018, 16'd24046, 16'd60836});
	test_expansion(128'hcd12c3a2c805405004bb28a6e2afa43a, {16'd39774, 16'd25186, 16'd51200, 16'd59811, 16'd47055, 16'd62498, 16'd29591, 16'd22957, 16'd55663, 16'd46742, 16'd15235, 16'd3504, 16'd24255, 16'd5071, 16'd61717, 16'd25125, 16'd37205, 16'd7860, 16'd48372, 16'd2317, 16'd26865, 16'd27591, 16'd29412, 16'd55333, 16'd50519, 16'd50934});
	test_expansion(128'hfcadcbbe9645203f6b3996cd665a482b, {16'd30317, 16'd41272, 16'd8077, 16'd5161, 16'd47616, 16'd57705, 16'd1024, 16'd56069, 16'd58595, 16'd38983, 16'd63037, 16'd2566, 16'd43894, 16'd30812, 16'd6231, 16'd41693, 16'd17703, 16'd34937, 16'd2552, 16'd55254, 16'd22425, 16'd45774, 16'd63342, 16'd37279, 16'd59232, 16'd2264});
	test_expansion(128'hefd60211975795df24f26faf8c0b116c, {16'd30799, 16'd35174, 16'd64489, 16'd29934, 16'd28280, 16'd22632, 16'd13508, 16'd18421, 16'd42608, 16'd37733, 16'd22997, 16'd6781, 16'd49959, 16'd42769, 16'd8169, 16'd32428, 16'd3371, 16'd17513, 16'd31691, 16'd8971, 16'd6950, 16'd24487, 16'd15273, 16'd41269, 16'd11221, 16'd20121});
	test_expansion(128'h8f30a719a9e65e7e913eeb151e1b3d0a, {16'd11059, 16'd28884, 16'd31710, 16'd13829, 16'd60121, 16'd34319, 16'd7302, 16'd25916, 16'd43840, 16'd38857, 16'd4693, 16'd17544, 16'd40362, 16'd5165, 16'd25639, 16'd29516, 16'd56435, 16'd60322, 16'd10655, 16'd37589, 16'd48548, 16'd5662, 16'd1945, 16'd48126, 16'd51578, 16'd63403});
	test_expansion(128'hd4e7776970a77c9f55a59e0f8a40e521, {16'd20284, 16'd57489, 16'd44040, 16'd64412, 16'd44775, 16'd56517, 16'd36129, 16'd52093, 16'd31092, 16'd12106, 16'd7326, 16'd37749, 16'd20942, 16'd50145, 16'd8366, 16'd7663, 16'd13714, 16'd61977, 16'd14277, 16'd54243, 16'd6197, 16'd43148, 16'd25907, 16'd61795, 16'd11186, 16'd57030});
	test_expansion(128'h32e8cac4d648df26f5e173b19c6e90ac, {16'd33827, 16'd11814, 16'd30634, 16'd19446, 16'd17373, 16'd1375, 16'd58576, 16'd61442, 16'd16560, 16'd15965, 16'd34240, 16'd19496, 16'd46228, 16'd55381, 16'd14898, 16'd40608, 16'd21113, 16'd11294, 16'd55988, 16'd2910, 16'd24827, 16'd49638, 16'd16669, 16'd53087, 16'd2457, 16'd43674});
	test_expansion(128'hdf46dd92a884e052b50c9836dc4f5408, {16'd54816, 16'd17448, 16'd42900, 16'd24479, 16'd17375, 16'd23457, 16'd13534, 16'd55708, 16'd57642, 16'd50273, 16'd35787, 16'd10188, 16'd61438, 16'd18872, 16'd32619, 16'd17177, 16'd9770, 16'd8268, 16'd24844, 16'd18444, 16'd58282, 16'd53225, 16'd15777, 16'd60695, 16'd19155, 16'd20262});
	test_expansion(128'hfaea8a29470aa8267103a59c3e754acd, {16'd23954, 16'd14835, 16'd35891, 16'd24557, 16'd49296, 16'd8216, 16'd38325, 16'd45784, 16'd36689, 16'd53264, 16'd27352, 16'd60636, 16'd17573, 16'd58640, 16'd46130, 16'd37258, 16'd33497, 16'd17933, 16'd26432, 16'd54984, 16'd38132, 16'd61504, 16'd53872, 16'd40941, 16'd3106, 16'd2093});
	test_expansion(128'hc43f156fa5a3ad2bf3d4b555b933fcb4, {16'd1097, 16'd54199, 16'd3387, 16'd18340, 16'd30006, 16'd52653, 16'd18258, 16'd56582, 16'd63895, 16'd64268, 16'd28377, 16'd22214, 16'd29839, 16'd31416, 16'd44252, 16'd400, 16'd45, 16'd1783, 16'd10348, 16'd50465, 16'd41007, 16'd149, 16'd22866, 16'd33789, 16'd62938, 16'd14918});
	test_expansion(128'h9317c18ae2afdda5513884b3f99e6145, {16'd17962, 16'd30110, 16'd5233, 16'd46100, 16'd32175, 16'd19150, 16'd1784, 16'd10045, 16'd11369, 16'd63938, 16'd1051, 16'd36001, 16'd46542, 16'd32601, 16'd7235, 16'd10929, 16'd33891, 16'd13098, 16'd15372, 16'd43917, 16'd14853, 16'd25324, 16'd34069, 16'd32058, 16'd31030, 16'd8499});
	test_expansion(128'h9d57e0de32d78e89277de0852980d3a7, {16'd37969, 16'd5348, 16'd46728, 16'd43994, 16'd58517, 16'd530, 16'd62031, 16'd12933, 16'd31735, 16'd5539, 16'd28403, 16'd52155, 16'd64762, 16'd8466, 16'd15784, 16'd14808, 16'd3304, 16'd12960, 16'd60451, 16'd7251, 16'd10278, 16'd56840, 16'd61610, 16'd7076, 16'd19550, 16'd763});
	test_expansion(128'h5abb45fbb8d720e30c4994f0c56fb6fd, {16'd7739, 16'd22587, 16'd57716, 16'd17586, 16'd34106, 16'd13982, 16'd3250, 16'd37349, 16'd38181, 16'd37816, 16'd46578, 16'd29512, 16'd43339, 16'd22219, 16'd1881, 16'd28811, 16'd63592, 16'd18230, 16'd20864, 16'd5157, 16'd48729, 16'd4541, 16'd647, 16'd58186, 16'd64168, 16'd14947});
	test_expansion(128'ha37bfc1f2bdb5a99b9dbbd4a627253ad, {16'd8124, 16'd29701, 16'd13318, 16'd8022, 16'd63384, 16'd29514, 16'd51071, 16'd24180, 16'd13748, 16'd38003, 16'd21946, 16'd5253, 16'd46392, 16'd55140, 16'd33400, 16'd46765, 16'd13508, 16'd30754, 16'd2867, 16'd5546, 16'd26967, 16'd63234, 16'd65150, 16'd58267, 16'd5817, 16'd30354});
	test_expansion(128'h9c227fdfde864ad72dcb313894001ef5, {16'd27427, 16'd38201, 16'd31494, 16'd40437, 16'd15848, 16'd41980, 16'd29520, 16'd11018, 16'd64376, 16'd57669, 16'd52354, 16'd23376, 16'd34182, 16'd31243, 16'd15552, 16'd12744, 16'd61961, 16'd13287, 16'd162, 16'd61174, 16'd11955, 16'd7620, 16'd41969, 16'd267, 16'd3006, 16'd46313});
	test_expansion(128'h7c8b47c0d78dc5e8fa8ec262a3a11596, {16'd63317, 16'd13550, 16'd17072, 16'd26247, 16'd44917, 16'd19718, 16'd35281, 16'd26335, 16'd15453, 16'd9133, 16'd15424, 16'd44813, 16'd22934, 16'd6139, 16'd52176, 16'd52202, 16'd51487, 16'd21083, 16'd26007, 16'd5090, 16'd36759, 16'd59059, 16'd29757, 16'd55505, 16'd34629, 16'd27076});
	test_expansion(128'h7b84e792eff6fd36f4b7c9ffd1a16618, {16'd35929, 16'd8825, 16'd5538, 16'd19265, 16'd4209, 16'd35383, 16'd25449, 16'd52358, 16'd48779, 16'd52026, 16'd54512, 16'd5086, 16'd37009, 16'd23407, 16'd21336, 16'd41619, 16'd64030, 16'd48837, 16'd8937, 16'd8228, 16'd11527, 16'd927, 16'd57828, 16'd59844, 16'd46667, 16'd46065});
	test_expansion(128'h9d326442bf091b12ab69d804fb899ad3, {16'd28878, 16'd32402, 16'd20921, 16'd19787, 16'd32092, 16'd34346, 16'd52015, 16'd21550, 16'd29608, 16'd1391, 16'd41341, 16'd55260, 16'd42987, 16'd35240, 16'd33489, 16'd16728, 16'd45288, 16'd30295, 16'd49954, 16'd4320, 16'd56482, 16'd58467, 16'd27694, 16'd7690, 16'd28760, 16'd2976});
	test_expansion(128'h6e64808ea48183993ceda166490a1201, {16'd61464, 16'd63824, 16'd57895, 16'd60678, 16'd31442, 16'd32533, 16'd8206, 16'd20186, 16'd3322, 16'd10550, 16'd56632, 16'd24641, 16'd27007, 16'd26305, 16'd64178, 16'd21924, 16'd13118, 16'd64256, 16'd7656, 16'd3242, 16'd14338, 16'd41811, 16'd44278, 16'd51427, 16'd44026, 16'd54620});
	test_expansion(128'h8e1f788b6d543ce3e6a3218474158526, {16'd50944, 16'd64641, 16'd15197, 16'd26022, 16'd14252, 16'd7762, 16'd20525, 16'd10790, 16'd43822, 16'd16491, 16'd17540, 16'd50848, 16'd40419, 16'd57976, 16'd35137, 16'd11926, 16'd54375, 16'd812, 16'd41948, 16'd31562, 16'd6322, 16'd44213, 16'd40836, 16'd34748, 16'd7557, 16'd37198});
	test_expansion(128'hdf0a25e42909fbeae0cd360cbae97c8f, {16'd28581, 16'd28634, 16'd59700, 16'd34018, 16'd56974, 16'd4859, 16'd5719, 16'd35827, 16'd8638, 16'd44237, 16'd57542, 16'd37263, 16'd30219, 16'd24206, 16'd19486, 16'd19847, 16'd18877, 16'd25848, 16'd45625, 16'd18642, 16'd41259, 16'd57096, 16'd45769, 16'd22782, 16'd11946, 16'd51012});
	test_expansion(128'h5263c1cd57884b7873725af274a4d904, {16'd7884, 16'd46913, 16'd38446, 16'd55846, 16'd47560, 16'd36173, 16'd25355, 16'd15487, 16'd30736, 16'd65326, 16'd848, 16'd2306, 16'd29255, 16'd48638, 16'd17727, 16'd58547, 16'd62157, 16'd28705, 16'd41490, 16'd30815, 16'd46403, 16'd1754, 16'd4094, 16'd34169, 16'd46261, 16'd38341});
	test_expansion(128'h8dcc89fb637906cade4cf41d842a7676, {16'd18819, 16'd15172, 16'd23309, 16'd38261, 16'd33457, 16'd62322, 16'd22571, 16'd14087, 16'd646, 16'd57084, 16'd12903, 16'd63053, 16'd27297, 16'd44834, 16'd9666, 16'd21528, 16'd63492, 16'd36626, 16'd13939, 16'd46226, 16'd18441, 16'd40571, 16'd42833, 16'd49559, 16'd38290, 16'd51176});
	test_expansion(128'hc5c2447ded3d24bee2f56f0eef55f336, {16'd26935, 16'd20245, 16'd10177, 16'd45083, 16'd15505, 16'd5248, 16'd7916, 16'd34219, 16'd46312, 16'd37450, 16'd42898, 16'd50461, 16'd2141, 16'd34081, 16'd53317, 16'd50733, 16'd43889, 16'd20886, 16'd39932, 16'd57980, 16'd24127, 16'd28112, 16'd34580, 16'd24819, 16'd1879, 16'd59534});
	test_expansion(128'h2a6ac50a2f7dc3bae838c08d5379496f, {16'd37431, 16'd13343, 16'd2352, 16'd28425, 16'd34253, 16'd39712, 16'd49487, 16'd34555, 16'd7430, 16'd23998, 16'd26365, 16'd33360, 16'd25432, 16'd31748, 16'd6966, 16'd22140, 16'd12889, 16'd28379, 16'd12105, 16'd30061, 16'd55370, 16'd11122, 16'd36918, 16'd23518, 16'd60526, 16'd14173});
	test_expansion(128'hb8091ca20301daa503c3fc0350aa5e89, {16'd50067, 16'd8599, 16'd47942, 16'd24214, 16'd55766, 16'd19906, 16'd58610, 16'd28875, 16'd25593, 16'd25363, 16'd63712, 16'd43093, 16'd11997, 16'd11343, 16'd61126, 16'd159, 16'd8815, 16'd25051, 16'd48649, 16'd29956, 16'd44289, 16'd46735, 16'd37323, 16'd38543, 16'd61045, 16'd11650});
	test_expansion(128'h529a49d9e24ecb89ed1d8c40325ae339, {16'd38615, 16'd64832, 16'd13084, 16'd47638, 16'd60139, 16'd36457, 16'd1746, 16'd32351, 16'd47404, 16'd50738, 16'd17920, 16'd35553, 16'd65187, 16'd38886, 16'd52226, 16'd21155, 16'd48775, 16'd47059, 16'd22515, 16'd53240, 16'd48490, 16'd31116, 16'd23954, 16'd49790, 16'd17032, 16'd9333});
	test_expansion(128'h19cacafb6337e150c2877117c772af5c, {16'd43674, 16'd38397, 16'd54344, 16'd27221, 16'd61855, 16'd64686, 16'd31626, 16'd13259, 16'd3954, 16'd27071, 16'd18371, 16'd28492, 16'd60196, 16'd54665, 16'd57635, 16'd10960, 16'd61192, 16'd55868, 16'd1842, 16'd15417, 16'd50034, 16'd53461, 16'd52219, 16'd28555, 16'd13125, 16'd34682});
	test_expansion(128'h48a92b234b807ea3c27e6dd09a22ec2f, {16'd32883, 16'd21178, 16'd6993, 16'd63736, 16'd13997, 16'd17586, 16'd10282, 16'd8437, 16'd1103, 16'd2509, 16'd32541, 16'd63406, 16'd17622, 16'd17984, 16'd2827, 16'd38388, 16'd10850, 16'd63079, 16'd43032, 16'd38631, 16'd60012, 16'd33114, 16'd54002, 16'd36800, 16'd45280, 16'd59560});
	test_expansion(128'h89ad9200fd9e8ef02f800f1c504f4faf, {16'd40886, 16'd11868, 16'd14646, 16'd26084, 16'd11623, 16'd10007, 16'd5654, 16'd62074, 16'd36411, 16'd24588, 16'd13815, 16'd16632, 16'd8031, 16'd39887, 16'd25884, 16'd12133, 16'd61765, 16'd13599, 16'd18891, 16'd12219, 16'd59520, 16'd62539, 16'd5273, 16'd61443, 16'd29554, 16'd30561});
	test_expansion(128'had00e28dfda43804e62f30cd777a2e91, {16'd10713, 16'd41872, 16'd63471, 16'd42728, 16'd31457, 16'd9479, 16'd35672, 16'd54286, 16'd63589, 16'd47121, 16'd32722, 16'd25746, 16'd7305, 16'd40538, 16'd43176, 16'd43610, 16'd15057, 16'd62507, 16'd14833, 16'd923, 16'd60099, 16'd63493, 16'd7179, 16'd25189, 16'd35754, 16'd16124});
	test_expansion(128'hfb3ca87b73094aea980b8f1580261e1f, {16'd7819, 16'd46390, 16'd43377, 16'd60614, 16'd20404, 16'd11779, 16'd49116, 16'd18582, 16'd64921, 16'd37804, 16'd19796, 16'd60414, 16'd57104, 16'd52148, 16'd55479, 16'd34130, 16'd28183, 16'd13173, 16'd11304, 16'd1493, 16'd36074, 16'd8592, 16'd36580, 16'd27733, 16'd11680, 16'd55947});
	test_expansion(128'h6c17b14eb21cafc5b9e92edc70fee38b, {16'd15465, 16'd15790, 16'd47291, 16'd33142, 16'd52801, 16'd14470, 16'd55047, 16'd62213, 16'd56569, 16'd25140, 16'd32509, 16'd30911, 16'd32568, 16'd40456, 16'd9101, 16'd52243, 16'd25710, 16'd36196, 16'd16683, 16'd18829, 16'd11937, 16'd51634, 16'd28203, 16'd4109, 16'd22582, 16'd60954});
	test_expansion(128'h3dc4da0fd8bf687077e8c9b8882888e8, {16'd4273, 16'd18136, 16'd38160, 16'd32006, 16'd24091, 16'd13694, 16'd32930, 16'd31304, 16'd16653, 16'd18798, 16'd17465, 16'd12037, 16'd54193, 16'd12272, 16'd40744, 16'd25267, 16'd22087, 16'd10419, 16'd47466, 16'd62810, 16'd33344, 16'd29875, 16'd44997, 16'd7654, 16'd15694, 16'd45440});
	test_expansion(128'h8766029878bb7a55353967cfd9a313fd, {16'd21402, 16'd1312, 16'd62824, 16'd52286, 16'd10903, 16'd60091, 16'd48052, 16'd59823, 16'd39713, 16'd23661, 16'd40300, 16'd62117, 16'd23985, 16'd50007, 16'd35973, 16'd16175, 16'd62326, 16'd34051, 16'd37385, 16'd16105, 16'd59309, 16'd47734, 16'd23234, 16'd53189, 16'd21730, 16'd8799});
	test_expansion(128'h7e3d8726f6f2360d7984b3766552515c, {16'd42939, 16'd44684, 16'd50217, 16'd35433, 16'd28767, 16'd1453, 16'd12104, 16'd32471, 16'd48021, 16'd65159, 16'd394, 16'd23407, 16'd39681, 16'd53783, 16'd2358, 16'd35521, 16'd46125, 16'd41821, 16'd19397, 16'd6049, 16'd47982, 16'd43527, 16'd37300, 16'd36872, 16'd41664, 16'd29033});
	test_expansion(128'h0d13cca76e9b07b55495fbca8d071891, {16'd52679, 16'd62934, 16'd9687, 16'd49859, 16'd30262, 16'd32495, 16'd705, 16'd20350, 16'd61897, 16'd34986, 16'd2689, 16'd12880, 16'd9729, 16'd1178, 16'd42614, 16'd12522, 16'd21859, 16'd11520, 16'd30665, 16'd43808, 16'd7286, 16'd9925, 16'd2395, 16'd30818, 16'd37790, 16'd35173});
	test_expansion(128'h0e19324a4a149edc577c5f82cabf11d6, {16'd10242, 16'd35413, 16'd30272, 16'd9818, 16'd33473, 16'd27006, 16'd25864, 16'd45460, 16'd51298, 16'd22357, 16'd52941, 16'd13744, 16'd6178, 16'd24642, 16'd28353, 16'd38, 16'd61071, 16'd48948, 16'd37741, 16'd61143, 16'd61791, 16'd53794, 16'd53374, 16'd57600, 16'd61356, 16'd37506});
	test_expansion(128'h19253ed8cc26b883c1abb2ee436dfd8e, {16'd23559, 16'd18513, 16'd65347, 16'd39505, 16'd44336, 16'd52815, 16'd19425, 16'd21356, 16'd61973, 16'd24685, 16'd35953, 16'd21840, 16'd13469, 16'd23456, 16'd1623, 16'd9121, 16'd59972, 16'd24511, 16'd1683, 16'd11525, 16'd39743, 16'd28349, 16'd40666, 16'd19312, 16'd59629, 16'd62605});
	test_expansion(128'h070ff4d65b58294a8ac573719219d47b, {16'd55121, 16'd27493, 16'd63724, 16'd54193, 16'd64942, 16'd64823, 16'd48149, 16'd17871, 16'd48931, 16'd26, 16'd6821, 16'd20951, 16'd9435, 16'd47324, 16'd13043, 16'd33749, 16'd1193, 16'd15833, 16'd35658, 16'd29597, 16'd12294, 16'd53884, 16'd30247, 16'd27555, 16'd59689, 16'd11635});
	test_expansion(128'hdbbf18b843a265c4125997a0bc8d3498, {16'd38359, 16'd14868, 16'd6144, 16'd9202, 16'd11536, 16'd24564, 16'd49883, 16'd19205, 16'd23013, 16'd48613, 16'd48491, 16'd52755, 16'd50322, 16'd64645, 16'd58558, 16'd12694, 16'd11961, 16'd4785, 16'd52701, 16'd42853, 16'd1948, 16'd63240, 16'd16175, 16'd41491, 16'd15812, 16'd4711});
	test_expansion(128'h0201271f5c2813247b779e49084251e8, {16'd26182, 16'd29409, 16'd21558, 16'd64334, 16'd56910, 16'd46632, 16'd7313, 16'd10164, 16'd60428, 16'd58169, 16'd31211, 16'd52571, 16'd45900, 16'd32381, 16'd27393, 16'd58738, 16'd27312, 16'd31731, 16'd21307, 16'd9496, 16'd15353, 16'd39602, 16'd633, 16'd6204, 16'd23042, 16'd19811});
	test_expansion(128'h55ad055cb9902c311f56b3e8ed03c138, {16'd37655, 16'd43516, 16'd17236, 16'd11349, 16'd49054, 16'd60708, 16'd30261, 16'd53623, 16'd8307, 16'd59361, 16'd62464, 16'd54268, 16'd6970, 16'd63763, 16'd52033, 16'd63979, 16'd23329, 16'd30667, 16'd2460, 16'd11815, 16'd35938, 16'd32096, 16'd63403, 16'd35172, 16'd23605, 16'd33037});
	test_expansion(128'h386fab21e2a05ce212600fcda105cc1d, {16'd14847, 16'd15652, 16'd56388, 16'd59072, 16'd34690, 16'd36406, 16'd32185, 16'd11357, 16'd24171, 16'd44455, 16'd5482, 16'd54585, 16'd35027, 16'd62965, 16'd16823, 16'd11719, 16'd28324, 16'd36713, 16'd21385, 16'd53441, 16'd40743, 16'd20195, 16'd4952, 16'd10417, 16'd48950, 16'd2315});
	test_expansion(128'hf2248461982c894b2815789340d0af58, {16'd41899, 16'd4871, 16'd41023, 16'd6849, 16'd3455, 16'd19563, 16'd26335, 16'd41294, 16'd3641, 16'd30507, 16'd54883, 16'd45743, 16'd65349, 16'd60350, 16'd45144, 16'd63479, 16'd30943, 16'd6028, 16'd24792, 16'd19220, 16'd44005, 16'd38791, 16'd62210, 16'd53469, 16'd2449, 16'd9283});
	test_expansion(128'h3201e95b396cb76cdd7f04742443437d, {16'd41512, 16'd53755, 16'd2318, 16'd39616, 16'd58869, 16'd52033, 16'd61828, 16'd38811, 16'd13459, 16'd15262, 16'd3172, 16'd23532, 16'd4425, 16'd43853, 16'd50446, 16'd20797, 16'd17842, 16'd58876, 16'd18054, 16'd38403, 16'd59601, 16'd53392, 16'd10491, 16'd7991, 16'd4816, 16'd45794});
	test_expansion(128'h7c2237a4f092988aeba99d4e2b2d1ed1, {16'd36516, 16'd647, 16'd7691, 16'd1714, 16'd336, 16'd52642, 16'd41642, 16'd17777, 16'd26009, 16'd65107, 16'd28580, 16'd2319, 16'd19403, 16'd4869, 16'd20675, 16'd59589, 16'd48603, 16'd33330, 16'd8814, 16'd22036, 16'd50217, 16'd32116, 16'd47704, 16'd49157, 16'd9811, 16'd20966});
	test_expansion(128'h01160b5d8cd8cc38b9bc53ba693fb9ee, {16'd43815, 16'd8466, 16'd7361, 16'd48252, 16'd17797, 16'd37183, 16'd60506, 16'd40689, 16'd55597, 16'd15488, 16'd18032, 16'd49979, 16'd21369, 16'd19144, 16'd49404, 16'd9407, 16'd56894, 16'd61920, 16'd7713, 16'd3316, 16'd7830, 16'd58938, 16'd50482, 16'd19803, 16'd48424, 16'd1552});
	test_expansion(128'hf042129916d434898c63671d8bfd1d43, {16'd28633, 16'd36656, 16'd50976, 16'd19171, 16'd25897, 16'd12834, 16'd30959, 16'd52158, 16'd46398, 16'd43930, 16'd17633, 16'd51392, 16'd64254, 16'd31625, 16'd35076, 16'd8953, 16'd59390, 16'd22010, 16'd5815, 16'd59113, 16'd32203, 16'd32656, 16'd7901, 16'd54946, 16'd13141, 16'd12160});
	test_expansion(128'h22947e54e3bf08e63e05c49dd999515a, {16'd55553, 16'd23113, 16'd62646, 16'd51959, 16'd23168, 16'd11887, 16'd14308, 16'd36378, 16'd36454, 16'd19119, 16'd65115, 16'd46932, 16'd58546, 16'd2025, 16'd22952, 16'd41427, 16'd51498, 16'd33047, 16'd29509, 16'd34366, 16'd34554, 16'd39475, 16'd34948, 16'd44801, 16'd58661, 16'd45277});
	test_expansion(128'h65dbe6fc0b387600e289fcf45b2ce8cb, {16'd59387, 16'd40093, 16'd54270, 16'd3100, 16'd30671, 16'd41428, 16'd35249, 16'd15517, 16'd50739, 16'd62149, 16'd37942, 16'd59174, 16'd36147, 16'd7222, 16'd50864, 16'd19133, 16'd33001, 16'd5220, 16'd29366, 16'd41929, 16'd47835, 16'd25443, 16'd4154, 16'd47024, 16'd40976, 16'd14118});
	test_expansion(128'ha2e8608faf7311e99ff2709b20665e6e, {16'd64865, 16'd24424, 16'd17035, 16'd35528, 16'd58291, 16'd47853, 16'd3814, 16'd58648, 16'd2286, 16'd8851, 16'd26850, 16'd18080, 16'd19557, 16'd6741, 16'd32463, 16'd30384, 16'd51116, 16'd16709, 16'd9429, 16'd43680, 16'd47563, 16'd65266, 16'd57071, 16'd5323, 16'd3749, 16'd50824});
	test_expansion(128'hdb43a8217b7b798f0bb4df68d5fe2f76, {16'd48141, 16'd58376, 16'd14399, 16'd10530, 16'd20386, 16'd11219, 16'd31116, 16'd37891, 16'd3238, 16'd17750, 16'd5413, 16'd24165, 16'd33211, 16'd37313, 16'd36166, 16'd24494, 16'd36271, 16'd59737, 16'd61953, 16'd30879, 16'd4614, 16'd30052, 16'd44852, 16'd9830, 16'd40554, 16'd12819});
	test_expansion(128'hc089846f76ef45716068753d9ec2b1b5, {16'd1514, 16'd63253, 16'd27937, 16'd4884, 16'd52741, 16'd55385, 16'd48867, 16'd57628, 16'd23575, 16'd23171, 16'd30500, 16'd307, 16'd18984, 16'd42316, 16'd4206, 16'd59624, 16'd10159, 16'd33214, 16'd54585, 16'd12537, 16'd48644, 16'd48066, 16'd34240, 16'd59258, 16'd17850, 16'd65283});
	test_expansion(128'h49aead0fc5711251f4302a0fd56cefd4, {16'd8900, 16'd28197, 16'd6550, 16'd52332, 16'd21664, 16'd444, 16'd45237, 16'd1831, 16'd9583, 16'd21284, 16'd13191, 16'd52623, 16'd60416, 16'd26626, 16'd50891, 16'd38334, 16'd2796, 16'd30334, 16'd1242, 16'd38528, 16'd62108, 16'd15068, 16'd63370, 16'd11848, 16'd46306, 16'd23533});
	test_expansion(128'h445458c55a344c0fc87a7d59e77b6d9a, {16'd18280, 16'd56687, 16'd7295, 16'd34316, 16'd14308, 16'd32783, 16'd586, 16'd16534, 16'd13236, 16'd63944, 16'd54973, 16'd45466, 16'd13753, 16'd46928, 16'd41125, 16'd63980, 16'd31971, 16'd18451, 16'd18854, 16'd30921, 16'd16320, 16'd29792, 16'd42365, 16'd45441, 16'd54375, 16'd55546});
	test_expansion(128'h4e1ccd49d64081975d0079e9fded2e0c, {16'd3723, 16'd63822, 16'd19115, 16'd36846, 16'd60126, 16'd63602, 16'd39859, 16'd24404, 16'd36612, 16'd51719, 16'd26627, 16'd22472, 16'd26630, 16'd56627, 16'd2151, 16'd50954, 16'd30590, 16'd2768, 16'd62403, 16'd55375, 16'd21507, 16'd22642, 16'd59048, 16'd64165, 16'd18467, 16'd47759});
	test_expansion(128'h95e6730abe6760036481a855a9e4477b, {16'd42, 16'd20508, 16'd36976, 16'd11846, 16'd44883, 16'd39028, 16'd63031, 16'd41610, 16'd13806, 16'd20269, 16'd60899, 16'd7118, 16'd51420, 16'd50813, 16'd15747, 16'd61315, 16'd21516, 16'd32359, 16'd14211, 16'd62461, 16'd33573, 16'd65067, 16'd54966, 16'd8442, 16'd18840, 16'd18626});
	test_expansion(128'h8706380a0134be77dabc82e951ab08c2, {16'd51827, 16'd15389, 16'd52393, 16'd7349, 16'd13691, 16'd62369, 16'd29188, 16'd59336, 16'd5098, 16'd17608, 16'd55666, 16'd35092, 16'd28596, 16'd22127, 16'd20607, 16'd38705, 16'd4765, 16'd45339, 16'd22079, 16'd3451, 16'd6921, 16'd57839, 16'd24638, 16'd62797, 16'd31923, 16'd51898});
	test_expansion(128'h2a6f86c3fd28ebcd054836ded35bb0cb, {16'd29542, 16'd4555, 16'd50778, 16'd9053, 16'd58300, 16'd17758, 16'd8832, 16'd41457, 16'd20482, 16'd19193, 16'd48501, 16'd9978, 16'd19090, 16'd54093, 16'd56335, 16'd56605, 16'd43153, 16'd6040, 16'd64113, 16'd49927, 16'd39821, 16'd14075, 16'd31426, 16'd44260, 16'd42483, 16'd7387});
	test_expansion(128'h4e6f69d77f63aaa3847376de2352d84e, {16'd48915, 16'd34870, 16'd18644, 16'd16913, 16'd11719, 16'd50624, 16'd18642, 16'd37741, 16'd62138, 16'd11274, 16'd48820, 16'd1350, 16'd11790, 16'd11066, 16'd3017, 16'd26430, 16'd38737, 16'd4899, 16'd65495, 16'd19417, 16'd13559, 16'd47105, 16'd20216, 16'd8930, 16'd46551, 16'd22637});
	test_expansion(128'h5b71d44437b5919a515e89d9d02420af, {16'd45730, 16'd64391, 16'd62161, 16'd62979, 16'd31443, 16'd4365, 16'd3711, 16'd16861, 16'd10298, 16'd51856, 16'd50593, 16'd8154, 16'd43917, 16'd2985, 16'd22493, 16'd32768, 16'd29470, 16'd54121, 16'd2653, 16'd53925, 16'd19921, 16'd59781, 16'd10271, 16'd25519, 16'd13064, 16'd46482});
	test_expansion(128'h238ea7f9322584a26abe8d4557124e5b, {16'd40281, 16'd50867, 16'd34942, 16'd57269, 16'd33422, 16'd33376, 16'd60809, 16'd35040, 16'd24366, 16'd12486, 16'd59757, 16'd46291, 16'd6646, 16'd14043, 16'd22172, 16'd25869, 16'd26914, 16'd17211, 16'd54304, 16'd14019, 16'd1474, 16'd1583, 16'd58289, 16'd24303, 16'd32683, 16'd1516});
	test_expansion(128'he0fa77e7aa8e05e9ac57ff7578df93d0, {16'd35262, 16'd22184, 16'd53220, 16'd30631, 16'd10695, 16'd39207, 16'd10702, 16'd8071, 16'd44844, 16'd44987, 16'd33466, 16'd7031, 16'd54333, 16'd54794, 16'd26132, 16'd13436, 16'd52395, 16'd65177, 16'd6606, 16'd54371, 16'd13142, 16'd5780, 16'd13143, 16'd32771, 16'd50515, 16'd280});
	test_expansion(128'h17a354cdbeb343cc1c8def3c2a529b82, {16'd34054, 16'd55233, 16'd65410, 16'd31725, 16'd35899, 16'd59693, 16'd49847, 16'd29547, 16'd64890, 16'd15222, 16'd34017, 16'd17619, 16'd18140, 16'd29416, 16'd35651, 16'd9686, 16'd36710, 16'd3081, 16'd17406, 16'd28634, 16'd5922, 16'd53964, 16'd4490, 16'd25617, 16'd57185, 16'd34809});
	test_expansion(128'h97f723f26b266ae68b137e981e7a30b8, {16'd61283, 16'd11312, 16'd33037, 16'd34202, 16'd43305, 16'd38493, 16'd47591, 16'd22225, 16'd29365, 16'd14400, 16'd17470, 16'd4594, 16'd52173, 16'd1018, 16'd56352, 16'd37307, 16'd62218, 16'd54967, 16'd29550, 16'd36758, 16'd44498, 16'd56909, 16'd44922, 16'd42622, 16'd37998, 16'd56410});
	test_expansion(128'hfefbc85cf0959449d3e9632c91bcb35a, {16'd60116, 16'd41650, 16'd5490, 16'd22649, 16'd45564, 16'd11956, 16'd64386, 16'd14919, 16'd55265, 16'd64973, 16'd8096, 16'd47804, 16'd41696, 16'd43297, 16'd22358, 16'd5624, 16'd18878, 16'd26445, 16'd6171, 16'd36269, 16'd54820, 16'd6515, 16'd48169, 16'd47704, 16'd17396, 16'd57046});
	test_expansion(128'hffdbb731ce984daee487cd6c25104496, {16'd21945, 16'd8448, 16'd6405, 16'd46343, 16'd44746, 16'd60062, 16'd7318, 16'd57514, 16'd22817, 16'd17043, 16'd39077, 16'd14095, 16'd42709, 16'd38521, 16'd46514, 16'd60900, 16'd58812, 16'd53684, 16'd24110, 16'd34599, 16'd55122, 16'd18033, 16'd47371, 16'd43162, 16'd62277, 16'd34899});
	test_expansion(128'hd2ad0e2cceb88a8ba2d8517578fa032e, {16'd54433, 16'd52444, 16'd17372, 16'd53865, 16'd51114, 16'd20807, 16'd33932, 16'd46906, 16'd59885, 16'd55952, 16'd44377, 16'd56561, 16'd3308, 16'd33853, 16'd47646, 16'd40746, 16'd51405, 16'd63269, 16'd60604, 16'd25251, 16'd16290, 16'd56782, 16'd50973, 16'd8170, 16'd63327, 16'd5983});
	test_expansion(128'h3cb6ea027b12e774f5269dc29c6b77cf, {16'd48979, 16'd61550, 16'd63166, 16'd24128, 16'd5796, 16'd36853, 16'd25883, 16'd29893, 16'd22605, 16'd63774, 16'd43387, 16'd48078, 16'd10321, 16'd34089, 16'd58618, 16'd34193, 16'd46546, 16'd17444, 16'd38193, 16'd11089, 16'd25405, 16'd12255, 16'd30833, 16'd62703, 16'd27869, 16'd6699});
	test_expansion(128'hf8de9399d069aef7641adbb2aadd3630, {16'd25881, 16'd49953, 16'd16550, 16'd13592, 16'd10057, 16'd2791, 16'd20073, 16'd55534, 16'd40766, 16'd51808, 16'd62079, 16'd10745, 16'd43243, 16'd19497, 16'd30939, 16'd37010, 16'd62459, 16'd26049, 16'd39103, 16'd9634, 16'd58208, 16'd21600, 16'd3019, 16'd19714, 16'd39849, 16'd56966});
	test_expansion(128'hb9d9242d7cf5a0a9ab417847bd279151, {16'd47373, 16'd35736, 16'd21899, 16'd48298, 16'd9763, 16'd29248, 16'd42952, 16'd12206, 16'd32948, 16'd29701, 16'd15402, 16'd3056, 16'd26610, 16'd39726, 16'd25382, 16'd63500, 16'd15439, 16'd35966, 16'd50644, 16'd54559, 16'd63799, 16'd46570, 16'd48920, 16'd32644, 16'd44042, 16'd3106});
	test_expansion(128'hfbf6193a6aaa99afe97b103c743985ad, {16'd22522, 16'd23907, 16'd459, 16'd45404, 16'd56029, 16'd60712, 16'd44421, 16'd58955, 16'd61204, 16'd18103, 16'd58160, 16'd14070, 16'd65463, 16'd45552, 16'd28030, 16'd3176, 16'd61073, 16'd9391, 16'd43807, 16'd59105, 16'd9784, 16'd54874, 16'd11996, 16'd64655, 16'd56396, 16'd41675});
	test_expansion(128'hfb10c556e615e443ae2940efde4fca47, {16'd38781, 16'd29708, 16'd50917, 16'd46432, 16'd38404, 16'd17234, 16'd64155, 16'd24781, 16'd27187, 16'd12983, 16'd13722, 16'd29649, 16'd16138, 16'd47991, 16'd29125, 16'd22889, 16'd32257, 16'd36425, 16'd4352, 16'd55456, 16'd50700, 16'd25575, 16'd53317, 16'd20678, 16'd42897, 16'd22600});
	test_expansion(128'h6eb77211504e05816d41d6481a1d9090, {16'd6845, 16'd2229, 16'd9043, 16'd50543, 16'd24261, 16'd9590, 16'd41205, 16'd19916, 16'd45725, 16'd44573, 16'd39476, 16'd3869, 16'd11275, 16'd11037, 16'd3691, 16'd25126, 16'd35098, 16'd8914, 16'd31658, 16'd39280, 16'd15555, 16'd60303, 16'd29804, 16'd1140, 16'd55194, 16'd5414});
	test_expansion(128'h608f7a1e4899c3a4a7955d0c4ec92008, {16'd48583, 16'd4816, 16'd9905, 16'd59390, 16'd1514, 16'd14814, 16'd15353, 16'd50349, 16'd15209, 16'd53199, 16'd14065, 16'd34287, 16'd60702, 16'd64990, 16'd41112, 16'd44026, 16'd19452, 16'd13832, 16'd16267, 16'd16326, 16'd42215, 16'd19005, 16'd5852, 16'd15083, 16'd32888, 16'd43796});
	test_expansion(128'h12e9b77af86ba81b6c35c86e341e7265, {16'd53488, 16'd11319, 16'd20011, 16'd56614, 16'd52031, 16'd791, 16'd65372, 16'd57591, 16'd20474, 16'd41840, 16'd50194, 16'd28589, 16'd65015, 16'd34414, 16'd8803, 16'd65217, 16'd34963, 16'd65090, 16'd43008, 16'd48969, 16'd60207, 16'd33853, 16'd1311, 16'd29186, 16'd44929, 16'd16878});
	test_expansion(128'h7590215c41958d26c84179126e6b9e36, {16'd44941, 16'd44136, 16'd4906, 16'd10798, 16'd34144, 16'd37318, 16'd59050, 16'd22947, 16'd54947, 16'd46156, 16'd9770, 16'd41116, 16'd5090, 16'd57002, 16'd50392, 16'd61281, 16'd16958, 16'd44896, 16'd24170, 16'd55555, 16'd49336, 16'd36830, 16'd60188, 16'd40443, 16'd14051, 16'd16405});
	test_expansion(128'hdce0e077e64169ccb7cb65f0c4785204, {16'd17620, 16'd48948, 16'd41483, 16'd53071, 16'd21033, 16'd29815, 16'd1297, 16'd62052, 16'd62806, 16'd27861, 16'd6062, 16'd45201, 16'd12330, 16'd14017, 16'd23474, 16'd29978, 16'd34577, 16'd59213, 16'd42199, 16'd4595, 16'd49890, 16'd7152, 16'd47635, 16'd44804, 16'd53491, 16'd18837});
	test_expansion(128'h10cb96678ee055a675baa944c9b24914, {16'd5775, 16'd15988, 16'd5856, 16'd25497, 16'd21844, 16'd55674, 16'd24536, 16'd64102, 16'd38722, 16'd33167, 16'd61327, 16'd34374, 16'd16534, 16'd58387, 16'd15360, 16'd40919, 16'd34181, 16'd62799, 16'd7764, 16'd25323, 16'd14687, 16'd13611, 16'd37635, 16'd29950, 16'd30062, 16'd20191});
	test_expansion(128'h7a14a70667ba8dc04bc600e56c7e7b74, {16'd53359, 16'd28794, 16'd54536, 16'd51984, 16'd35779, 16'd18878, 16'd35286, 16'd62018, 16'd61281, 16'd16950, 16'd29546, 16'd50746, 16'd9084, 16'd9304, 16'd22377, 16'd27154, 16'd58738, 16'd8273, 16'd27845, 16'd52896, 16'd7381, 16'd11608, 16'd54686, 16'd8754, 16'd22919, 16'd38528});
	test_expansion(128'h6b787bdcc9209ce6c70fdc912ab5de83, {16'd32735, 16'd15647, 16'd47966, 16'd19678, 16'd42935, 16'd56336, 16'd19976, 16'd61827, 16'd19294, 16'd4206, 16'd9763, 16'd2809, 16'd39455, 16'd46076, 16'd54212, 16'd16598, 16'd35092, 16'd36559, 16'd56650, 16'd13536, 16'd4898, 16'd31859, 16'd63749, 16'd23783, 16'd50287, 16'd14618});
	test_expansion(128'hca86dbe6e13c98afaffeaa6f1c65cb3b, {16'd14541, 16'd35329, 16'd24734, 16'd13186, 16'd54843, 16'd4357, 16'd53385, 16'd10466, 16'd42750, 16'd56778, 16'd24186, 16'd48721, 16'd57663, 16'd50790, 16'd61524, 16'd52375, 16'd28235, 16'd17822, 16'd59426, 16'd44205, 16'd4578, 16'd56237, 16'd41959, 16'd12996, 16'd23379, 16'd35334});
	test_expansion(128'h1fada7ff2e4b2099a7e0f9f7cc2fd387, {16'd22984, 16'd14167, 16'd53121, 16'd7928, 16'd5961, 16'd16501, 16'd38653, 16'd1609, 16'd44798, 16'd48238, 16'd44013, 16'd44646, 16'd28994, 16'd34238, 16'd16946, 16'd11401, 16'd14341, 16'd53775, 16'd18939, 16'd48111, 16'd3926, 16'd18322, 16'd8578, 16'd45274, 16'd2383, 16'd65452});
	test_expansion(128'h45c6d4106546780d9589f8c43d7be202, {16'd33853, 16'd200, 16'd36709, 16'd3593, 16'd60556, 16'd61104, 16'd16818, 16'd1413, 16'd25511, 16'd23426, 16'd11398, 16'd15823, 16'd3533, 16'd40865, 16'd16593, 16'd34141, 16'd63418, 16'd58984, 16'd30712, 16'd11588, 16'd17380, 16'd21910, 16'd19556, 16'd19027, 16'd54421, 16'd976});
	test_expansion(128'h69b7cdf0b46cd3ace948563189cd70df, {16'd12534, 16'd44582, 16'd19416, 16'd16984, 16'd28862, 16'd17838, 16'd31520, 16'd60562, 16'd9375, 16'd24287, 16'd48001, 16'd50867, 16'd33153, 16'd54040, 16'd56279, 16'd11428, 16'd52306, 16'd47209, 16'd52649, 16'd59653, 16'd41853, 16'd18116, 16'd58417, 16'd52826, 16'd13818, 16'd24742});
	test_expansion(128'hf71a8c9cf3a3fe02db42925ffe82aaab, {16'd30694, 16'd8599, 16'd7774, 16'd18054, 16'd37500, 16'd48797, 16'd17741, 16'd33964, 16'd22623, 16'd24763, 16'd50429, 16'd61943, 16'd52728, 16'd29359, 16'd42706, 16'd14216, 16'd14372, 16'd28384, 16'd39535, 16'd11846, 16'd8572, 16'd8891, 16'd21437, 16'd29329, 16'd41094, 16'd61299});
	test_expansion(128'h2ef261c7182799b1e7e1d8050326743d, {16'd9547, 16'd6170, 16'd42787, 16'd60285, 16'd12198, 16'd35620, 16'd39712, 16'd22406, 16'd34187, 16'd21293, 16'd941, 16'd53956, 16'd61348, 16'd13336, 16'd12564, 16'd29690, 16'd36504, 16'd23434, 16'd52553, 16'd20738, 16'd8106, 16'd31466, 16'd55295, 16'd18254, 16'd48925, 16'd58357});
	test_expansion(128'h9f3ea3df0b1a56afe8d976eabe6d028a, {16'd54991, 16'd40094, 16'd55031, 16'd1912, 16'd19490, 16'd39821, 16'd4660, 16'd22819, 16'd41031, 16'd6937, 16'd58023, 16'd45649, 16'd21565, 16'd47839, 16'd44034, 16'd50284, 16'd31611, 16'd59438, 16'd27481, 16'd32538, 16'd48699, 16'd25886, 16'd50923, 16'd37778, 16'd29478, 16'd48260});
	test_expansion(128'he966a9cb36a868b50cccbcc84ea86740, {16'd12068, 16'd12326, 16'd32813, 16'd23001, 16'd22585, 16'd24044, 16'd49391, 16'd17825, 16'd35622, 16'd25305, 16'd37662, 16'd10547, 16'd55858, 16'd22124, 16'd33212, 16'd32520, 16'd2802, 16'd43334, 16'd1101, 16'd29855, 16'd11588, 16'd59766, 16'd60264, 16'd28457, 16'd50056, 16'd54604});
	test_expansion(128'hb590bc256240f883ec82197cfaead33d, {16'd35044, 16'd2404, 16'd17168, 16'd10734, 16'd26158, 16'd27300, 16'd54946, 16'd39651, 16'd25496, 16'd22677, 16'd60483, 16'd48314, 16'd9044, 16'd53762, 16'd12999, 16'd7743, 16'd36222, 16'd57942, 16'd49982, 16'd25237, 16'd39394, 16'd37887, 16'd13638, 16'd46182, 16'd21880, 16'd53519});
	test_expansion(128'h28998f1f62e2f0b40679c65189f8b2de, {16'd53478, 16'd56224, 16'd29123, 16'd3579, 16'd63952, 16'd1158, 16'd59541, 16'd5799, 16'd36950, 16'd49019, 16'd63848, 16'd26767, 16'd34447, 16'd48825, 16'd47484, 16'd25566, 16'd33657, 16'd7724, 16'd34906, 16'd64264, 16'd18205, 16'd3661, 16'd34978, 16'd55094, 16'd708, 16'd58082});
	test_expansion(128'h1b59721e2f2b20f532a6745c0285fe2c, {16'd47054, 16'd3538, 16'd14357, 16'd22021, 16'd34451, 16'd1728, 16'd53833, 16'd25500, 16'd13741, 16'd12298, 16'd13776, 16'd20214, 16'd34311, 16'd40032, 16'd4430, 16'd511, 16'd27772, 16'd10353, 16'd23218, 16'd27654, 16'd1856, 16'd49503, 16'd62770, 16'd15479, 16'd21862, 16'd10322});
	test_expansion(128'h02b79ead9d2b34b82c035c6bf199ce52, {16'd27636, 16'd29960, 16'd31221, 16'd16950, 16'd42824, 16'd18614, 16'd9802, 16'd21481, 16'd49207, 16'd62109, 16'd63266, 16'd51150, 16'd18385, 16'd5676, 16'd51118, 16'd8205, 16'd12465, 16'd2472, 16'd29392, 16'd34107, 16'd47672, 16'd12703, 16'd22956, 16'd16064, 16'd13610, 16'd64537});
	test_expansion(128'h229dc73646181c30798a6248bc803d1d, {16'd32291, 16'd32875, 16'd58941, 16'd55528, 16'd17983, 16'd9559, 16'd59924, 16'd32626, 16'd14745, 16'd62944, 16'd46904, 16'd53182, 16'd30986, 16'd8197, 16'd50009, 16'd13496, 16'd9453, 16'd8165, 16'd21772, 16'd4398, 16'd7262, 16'd34888, 16'd40636, 16'd54627, 16'd40011, 16'd39920});
	test_expansion(128'h54d0109e201a61f34e6865807f4bcd8b, {16'd19390, 16'd58066, 16'd16523, 16'd57720, 16'd54103, 16'd18523, 16'd46212, 16'd25353, 16'd55206, 16'd47244, 16'd23862, 16'd54730, 16'd59468, 16'd58603, 16'd65251, 16'd31243, 16'd58172, 16'd31410, 16'd47399, 16'd32385, 16'd41861, 16'd17990, 16'd21363, 16'd6656, 16'd4966, 16'd59611});
	test_expansion(128'h18634d2ac1f3aa729d2dfd381288bdeb, {16'd3838, 16'd12846, 16'd5005, 16'd27505, 16'd36665, 16'd1226, 16'd23988, 16'd65011, 16'd35947, 16'd65330, 16'd54761, 16'd34686, 16'd14347, 16'd16844, 16'd18448, 16'd9737, 16'd11266, 16'd40483, 16'd22784, 16'd1034, 16'd4617, 16'd46153, 16'd42265, 16'd64489, 16'd57811, 16'd32027});
	test_expansion(128'hccbfd0441ebe033b156a5306dc5354a5, {16'd19411, 16'd15430, 16'd29758, 16'd49254, 16'd45235, 16'd31619, 16'd10763, 16'd60397, 16'd15913, 16'd33783, 16'd38533, 16'd10965, 16'd25229, 16'd43317, 16'd27946, 16'd43082, 16'd62951, 16'd10725, 16'd43876, 16'd60352, 16'd56465, 16'd31238, 16'd20096, 16'd45547, 16'd41792, 16'd2628});
	test_expansion(128'hed6f6dd45f8fc4abfc86d62b4a4c14d9, {16'd63444, 16'd55760, 16'd21179, 16'd6445, 16'd14061, 16'd10292, 16'd57004, 16'd5465, 16'd64134, 16'd55030, 16'd56607, 16'd11009, 16'd13436, 16'd6995, 16'd35892, 16'd57928, 16'd59439, 16'd43654, 16'd62749, 16'd15992, 16'd34579, 16'd9412, 16'd7591, 16'd54432, 16'd35408, 16'd22366});
	test_expansion(128'h3e1c74b19eb11b2ed58bd2b100546571, {16'd21236, 16'd63562, 16'd35251, 16'd17697, 16'd33324, 16'd41604, 16'd16963, 16'd29174, 16'd31073, 16'd18862, 16'd61986, 16'd53928, 16'd11464, 16'd28296, 16'd43667, 16'd26778, 16'd23577, 16'd30049, 16'd40199, 16'd15466, 16'd55063, 16'd5397, 16'd2180, 16'd60152, 16'd4000, 16'd27812});
	test_expansion(128'hc72d4ed3b76c3d36445510c5a841b613, {16'd13998, 16'd28965, 16'd56688, 16'd5223, 16'd26936, 16'd4284, 16'd5411, 16'd31792, 16'd2343, 16'd59091, 16'd10501, 16'd5302, 16'd51036, 16'd24069, 16'd34600, 16'd32211, 16'd37587, 16'd3314, 16'd51616, 16'd53600, 16'd29873, 16'd58183, 16'd64227, 16'd32731, 16'd38775, 16'd58750});
	test_expansion(128'hc3e682035476ae4355f473ee6020462a, {16'd51228, 16'd59820, 16'd58721, 16'd51811, 16'd41025, 16'd56233, 16'd21815, 16'd35666, 16'd17101, 16'd46194, 16'd34121, 16'd43879, 16'd44872, 16'd20079, 16'd26752, 16'd35993, 16'd24831, 16'd31101, 16'd11904, 16'd60857, 16'd16014, 16'd42291, 16'd65130, 16'd29123, 16'd54178, 16'd51208});
	test_expansion(128'h05800f90dec8d93298e4cb4c0d6fdaac, {16'd54820, 16'd23779, 16'd44252, 16'd26650, 16'd63220, 16'd47082, 16'd35846, 16'd29034, 16'd19396, 16'd30173, 16'd137, 16'd28386, 16'd47097, 16'd58706, 16'd36393, 16'd3495, 16'd18265, 16'd55948, 16'd47977, 16'd40039, 16'd44111, 16'd57661, 16'd39404, 16'd30977, 16'd30832, 16'd48519});
	test_expansion(128'hbc8e7f61a3eb40b75306bb09987a71ba, {16'd4994, 16'd2997, 16'd64889, 16'd37293, 16'd4398, 16'd16980, 16'd62428, 16'd58036, 16'd42193, 16'd18137, 16'd56137, 16'd45280, 16'd56030, 16'd34307, 16'd17922, 16'd52942, 16'd35523, 16'd30812, 16'd42298, 16'd2714, 16'd8729, 16'd27282, 16'd18481, 16'd58796, 16'd61807, 16'd32054});
	test_expansion(128'hf2b5482e23d60dace568ccbde5a198ea, {16'd11059, 16'd40195, 16'd21107, 16'd14349, 16'd4357, 16'd2345, 16'd32169, 16'd7443, 16'd59860, 16'd4003, 16'd1120, 16'd31790, 16'd6856, 16'd19667, 16'd64985, 16'd31195, 16'd2211, 16'd21066, 16'd4343, 16'd56262, 16'd53764, 16'd7025, 16'd7233, 16'd50049, 16'd51711, 16'd39315});
	test_expansion(128'h26ac951a98bbec059e1db1f18819f462, {16'd64448, 16'd23151, 16'd50293, 16'd54295, 16'd9210, 16'd11459, 16'd62875, 16'd48867, 16'd64967, 16'd29622, 16'd40730, 16'd6711, 16'd24885, 16'd1288, 16'd4290, 16'd24339, 16'd52721, 16'd46428, 16'd47839, 16'd6001, 16'd33256, 16'd38192, 16'd31690, 16'd42389, 16'd10536, 16'd42984});
	test_expansion(128'h6aedcdb00b1c9f48fea1931698bc8e5c, {16'd38876, 16'd38582, 16'd47735, 16'd11220, 16'd42453, 16'd12465, 16'd35226, 16'd50557, 16'd245, 16'd32157, 16'd65156, 16'd53639, 16'd22791, 16'd57679, 16'd13069, 16'd29222, 16'd45499, 16'd35139, 16'd1634, 16'd61776, 16'd7861, 16'd14727, 16'd21424, 16'd44904, 16'd42189, 16'd61201});
	test_expansion(128'hccfc837d2fafac31532b0fb62569a12a, {16'd41027, 16'd40834, 16'd51212, 16'd30063, 16'd62005, 16'd7111, 16'd29639, 16'd14387, 16'd60695, 16'd5386, 16'd44132, 16'd54870, 16'd29313, 16'd9251, 16'd34572, 16'd37471, 16'd51542, 16'd33984, 16'd45920, 16'd27532, 16'd2231, 16'd63876, 16'd39658, 16'd3182, 16'd20597, 16'd7826});
	test_expansion(128'h3a231d1a7cd30cde4dbe51a4f072e460, {16'd15050, 16'd5290, 16'd41217, 16'd1017, 16'd7039, 16'd4803, 16'd55131, 16'd53537, 16'd46882, 16'd54108, 16'd15206, 16'd25948, 16'd55434, 16'd58387, 16'd37950, 16'd15839, 16'd59281, 16'd47743, 16'd13200, 16'd25548, 16'd52804, 16'd53798, 16'd14883, 16'd30099, 16'd32318, 16'd15289});
	test_expansion(128'h562236deb9b0c3123ebcea87e394eba5, {16'd22241, 16'd11925, 16'd64134, 16'd40275, 16'd35030, 16'd41828, 16'd47772, 16'd26554, 16'd51713, 16'd59555, 16'd62570, 16'd8687, 16'd64946, 16'd56890, 16'd31616, 16'd59863, 16'd46224, 16'd25298, 16'd19457, 16'd45798, 16'd65255, 16'd30623, 16'd5331, 16'd30659, 16'd54695, 16'd59613});
	test_expansion(128'hc6e26e1cd534a36a2a5a2366a6ec664e, {16'd39951, 16'd22416, 16'd38678, 16'd41857, 16'd59115, 16'd58055, 16'd213, 16'd43932, 16'd55184, 16'd49236, 16'd22258, 16'd43573, 16'd27367, 16'd2541, 16'd29545, 16'd47178, 16'd26179, 16'd15361, 16'd25343, 16'd6488, 16'd50289, 16'd39823, 16'd24265, 16'd8895, 16'd52136, 16'd13999});
	test_expansion(128'h52be4c8a7dff3f6031b319e97c3716d7, {16'd44029, 16'd10325, 16'd42171, 16'd18098, 16'd43781, 16'd28289, 16'd41289, 16'd51807, 16'd7335, 16'd22209, 16'd25359, 16'd5164, 16'd31221, 16'd5531, 16'd32275, 16'd35469, 16'd50810, 16'd8760, 16'd25226, 16'd30232, 16'd52815, 16'd2429, 16'd46226, 16'd29943, 16'd44695, 16'd42062});
	test_expansion(128'h6abc7f1cc01c1ab24ed66222fc1a7eec, {16'd9350, 16'd49080, 16'd27622, 16'd48898, 16'd52911, 16'd35545, 16'd27373, 16'd54376, 16'd3137, 16'd18126, 16'd9956, 16'd60931, 16'd61765, 16'd229, 16'd1155, 16'd2255, 16'd12016, 16'd1207, 16'd13117, 16'd4450, 16'd52930, 16'd33135, 16'd34063, 16'd1713, 16'd355, 16'd37257});
	test_expansion(128'h686efcc9d7dd33a3401750624de34703, {16'd48762, 16'd33608, 16'd55847, 16'd7495, 16'd16580, 16'd64883, 16'd43175, 16'd29008, 16'd23641, 16'd28310, 16'd10777, 16'd44887, 16'd1396, 16'd8913, 16'd36428, 16'd46198, 16'd25309, 16'd47089, 16'd63086, 16'd31596, 16'd10472, 16'd25335, 16'd43066, 16'd49712, 16'd10509, 16'd48572});
	test_expansion(128'haa8ebcb8cd03a1fd6c264f5bf52c708e, {16'd59808, 16'd27166, 16'd4252, 16'd10798, 16'd45392, 16'd60000, 16'd20323, 16'd27267, 16'd32849, 16'd24186, 16'd24042, 16'd42940, 16'd11197, 16'd54988, 16'd58016, 16'd64203, 16'd54096, 16'd15429, 16'd35715, 16'd40009, 16'd2880, 16'd2573, 16'd30112, 16'd2462, 16'd46763, 16'd33811});
	test_expansion(128'h9aed034bc1daa85abfe1393bc94d83a9, {16'd58187, 16'd44615, 16'd46239, 16'd21188, 16'd41551, 16'd34763, 16'd41019, 16'd51729, 16'd23146, 16'd32103, 16'd57823, 16'd48728, 16'd29315, 16'd17578, 16'd9158, 16'd30182, 16'd29834, 16'd62231, 16'd20809, 16'd3442, 16'd58343, 16'd4239, 16'd57767, 16'd16424, 16'd34038, 16'd25196});
	test_expansion(128'h23214486957d9c6516191d197292f941, {16'd36804, 16'd60153, 16'd4020, 16'd8673, 16'd55310, 16'd33037, 16'd18358, 16'd6355, 16'd62557, 16'd15120, 16'd62160, 16'd7787, 16'd6840, 16'd24593, 16'd45149, 16'd59191, 16'd24551, 16'd56423, 16'd4086, 16'd14282, 16'd51648, 16'd53658, 16'd16165, 16'd23111, 16'd31245, 16'd65137});
	test_expansion(128'h2514cbc80c2e715028e780ed6e285491, {16'd9918, 16'd2004, 16'd12748, 16'd32210, 16'd45285, 16'd4397, 16'd12408, 16'd20528, 16'd44494, 16'd26876, 16'd37400, 16'd44548, 16'd112, 16'd61836, 16'd27406, 16'd41477, 16'd30635, 16'd1929, 16'd21102, 16'd21406, 16'd51581, 16'd32955, 16'd22110, 16'd30436, 16'd16292, 16'd52767});
	test_expansion(128'hae148a16b97fd611a41b97a7a99e47a8, {16'd15785, 16'd19881, 16'd37840, 16'd9827, 16'd28452, 16'd33097, 16'd61309, 16'd22375, 16'd58395, 16'd37451, 16'd50240, 16'd56186, 16'd56535, 16'd57533, 16'd47197, 16'd45774, 16'd52994, 16'd53003, 16'd56828, 16'd34815, 16'd47702, 16'd18150, 16'd20357, 16'd42154, 16'd17729, 16'd64001});
	test_expansion(128'h3e25f5a4738e00f02b2bffbe5344a0d7, {16'd30549, 16'd19866, 16'd33450, 16'd14409, 16'd41431, 16'd35588, 16'd26787, 16'd17556, 16'd57488, 16'd38966, 16'd57733, 16'd12873, 16'd54578, 16'd32836, 16'd21010, 16'd59115, 16'd46446, 16'd35554, 16'd49912, 16'd18587, 16'd1017, 16'd49496, 16'd604, 16'd50894, 16'd44743, 16'd35422});
	test_expansion(128'hbf28baa4729ceff2df91fa54d55587f6, {16'd53751, 16'd23658, 16'd48194, 16'd42939, 16'd6544, 16'd10703, 16'd60446, 16'd34819, 16'd64047, 16'd62964, 16'd51715, 16'd14125, 16'd52274, 16'd1003, 16'd23710, 16'd11510, 16'd64565, 16'd7206, 16'd2237, 16'd20645, 16'd14697, 16'd54466, 16'd49725, 16'd20226, 16'd5101, 16'd60409});
	test_expansion(128'hb49876b2930728f2554b3cb151be2444, {16'd42207, 16'd13043, 16'd56175, 16'd41406, 16'd54511, 16'd50299, 16'd40126, 16'd39141, 16'd10830, 16'd44912, 16'd46482, 16'd38358, 16'd58490, 16'd50526, 16'd29112, 16'd55242, 16'd55140, 16'd25673, 16'd44325, 16'd50896, 16'd8535, 16'd17242, 16'd49982, 16'd36942, 16'd36152, 16'd42601});
	test_expansion(128'hff12fbb3f46c4a4fd41fdf0a6455803e, {16'd6398, 16'd101, 16'd52514, 16'd64105, 16'd37534, 16'd45914, 16'd48718, 16'd16784, 16'd13627, 16'd657, 16'd51745, 16'd40746, 16'd29390, 16'd62970, 16'd620, 16'd42137, 16'd19486, 16'd6959, 16'd63302, 16'd37038, 16'd49033, 16'd34493, 16'd45605, 16'd48175, 16'd5383, 16'd8631});
	test_expansion(128'h54c20d84458c6c2ff3d7b46dc2a0ae9e, {16'd63456, 16'd50567, 16'd8755, 16'd9417, 16'd42348, 16'd511, 16'd29076, 16'd6864, 16'd6154, 16'd32280, 16'd53386, 16'd31003, 16'd62111, 16'd62645, 16'd12451, 16'd10926, 16'd46221, 16'd9829, 16'd31169, 16'd22353, 16'd14756, 16'd31955, 16'd7647, 16'd8432, 16'd58479, 16'd26086});
	test_expansion(128'hb1d883df2511791a860aee517a666f68, {16'd2930, 16'd28269, 16'd61249, 16'd57403, 16'd32947, 16'd29341, 16'd53027, 16'd10299, 16'd19429, 16'd23842, 16'd57647, 16'd21190, 16'd47742, 16'd2446, 16'd58076, 16'd59079, 16'd62895, 16'd26702, 16'd36647, 16'd53138, 16'd18754, 16'd34112, 16'd12701, 16'd43506, 16'd16720, 16'd25377});
	test_expansion(128'hdebde833f557f72da92c90e956c61e1b, {16'd49117, 16'd62720, 16'd19438, 16'd17643, 16'd49015, 16'd63484, 16'd21289, 16'd22408, 16'd6990, 16'd17127, 16'd76, 16'd28328, 16'd22913, 16'd14190, 16'd39507, 16'd36309, 16'd53062, 16'd58725, 16'd10253, 16'd39865, 16'd35386, 16'd45712, 16'd27677, 16'd39086, 16'd9814, 16'd9059});
	test_expansion(128'hcbed4ae110c6b4eb92e3900a68c0652c, {16'd9909, 16'd53570, 16'd15034, 16'd1638, 16'd40957, 16'd2916, 16'd41173, 16'd44994, 16'd39268, 16'd48482, 16'd22301, 16'd26819, 16'd57137, 16'd25756, 16'd40613, 16'd61428, 16'd60936, 16'd47157, 16'd57635, 16'd6667, 16'd6646, 16'd28009, 16'd14291, 16'd33056, 16'd23025, 16'd10262});
	test_expansion(128'hfca8199f8cb5067a89d36ee8c33181ac, {16'd29038, 16'd7248, 16'd15064, 16'd39317, 16'd19824, 16'd21659, 16'd4054, 16'd54741, 16'd19354, 16'd35134, 16'd47162, 16'd31141, 16'd39136, 16'd16929, 16'd13784, 16'd3209, 16'd7440, 16'd63623, 16'd10917, 16'd25247, 16'd53599, 16'd23148, 16'd3127, 16'd44013, 16'd5804, 16'd49901});
	test_expansion(128'h9bd69bf682dc2f1c362e7991805da926, {16'd49733, 16'd28591, 16'd50779, 16'd63571, 16'd4156, 16'd58251, 16'd34819, 16'd64340, 16'd12061, 16'd5121, 16'd7552, 16'd35597, 16'd33718, 16'd49144, 16'd32335, 16'd13590, 16'd48570, 16'd14495, 16'd8083, 16'd32932, 16'd35436, 16'd55730, 16'd29339, 16'd43641, 16'd26854, 16'd36638});
	test_expansion(128'h3d50841e1008405f317396472f2254cb, {16'd10164, 16'd25745, 16'd38812, 16'd46009, 16'd17205, 16'd46367, 16'd40176, 16'd10842, 16'd57547, 16'd25296, 16'd48507, 16'd28887, 16'd63390, 16'd38466, 16'd30837, 16'd59406, 16'd27158, 16'd40761, 16'd26453, 16'd29582, 16'd1688, 16'd42305, 16'd62229, 16'd14211, 16'd14497, 16'd21570});
	test_expansion(128'h7cc6b37e183a0d4ea10741822d07ce26, {16'd20370, 16'd12898, 16'd56031, 16'd52939, 16'd63856, 16'd11300, 16'd38566, 16'd19003, 16'd11702, 16'd22717, 16'd41077, 16'd58525, 16'd5917, 16'd56858, 16'd39027, 16'd17333, 16'd41396, 16'd32113, 16'd63488, 16'd49905, 16'd30997, 16'd26290, 16'd38453, 16'd64473, 16'd28873, 16'd4972});
	test_expansion(128'h32624cd08de3c2b2322bc6f46f5b74be, {16'd14163, 16'd45585, 16'd54579, 16'd55117, 16'd51909, 16'd56234, 16'd9139, 16'd36160, 16'd15766, 16'd8341, 16'd37983, 16'd7162, 16'd16973, 16'd17131, 16'd48627, 16'd24857, 16'd11582, 16'd40678, 16'd47588, 16'd2806, 16'd19954, 16'd24482, 16'd34872, 16'd44885, 16'd43034, 16'd17404});
	test_expansion(128'h219a978f785402bf65888ab24c966944, {16'd19390, 16'd6775, 16'd26562, 16'd30540, 16'd47672, 16'd25456, 16'd61142, 16'd63526, 16'd32928, 16'd18472, 16'd50025, 16'd40523, 16'd322, 16'd28438, 16'd14376, 16'd36207, 16'd19856, 16'd58694, 16'd29060, 16'd53217, 16'd39391, 16'd28653, 16'd33863, 16'd58908, 16'd21245, 16'd10291});
	test_expansion(128'h82ad7ad1bffea62afc76f03b3f0c9de6, {16'd65321, 16'd53957, 16'd3693, 16'd8824, 16'd50910, 16'd31955, 16'd57528, 16'd27216, 16'd15879, 16'd50505, 16'd34837, 16'd18851, 16'd4621, 16'd11023, 16'd9944, 16'd33422, 16'd43181, 16'd43345, 16'd20503, 16'd63164, 16'd36058, 16'd28345, 16'd9619, 16'd57957, 16'd50873, 16'd41006});
	test_expansion(128'h2f8705bb5ff7e7cb7be2f679bfa10e39, {16'd26252, 16'd54509, 16'd44231, 16'd26065, 16'd53794, 16'd27530, 16'd45427, 16'd39221, 16'd27311, 16'd4905, 16'd53261, 16'd30318, 16'd63658, 16'd43946, 16'd52667, 16'd42405, 16'd25628, 16'd13756, 16'd10477, 16'd36471, 16'd45901, 16'd49971, 16'd17929, 16'd38882, 16'd50599, 16'd49901});
	test_expansion(128'hc00f0d4f2b33ecab61559e08717ff7a7, {16'd64365, 16'd4204, 16'd35829, 16'd54408, 16'd4080, 16'd47545, 16'd30011, 16'd4044, 16'd62764, 16'd24629, 16'd65493, 16'd18375, 16'd10322, 16'd60023, 16'd50974, 16'd48188, 16'd25129, 16'd1601, 16'd54212, 16'd46701, 16'd15377, 16'd14478, 16'd19886, 16'd61699, 16'd21190, 16'd46858});
	test_expansion(128'h7482bdaa25b0abb2b2ac902f5afef9df, {16'd39410, 16'd24290, 16'd38108, 16'd41869, 16'd9948, 16'd39719, 16'd15809, 16'd27228, 16'd62496, 16'd50894, 16'd27552, 16'd20537, 16'd11549, 16'd18610, 16'd56522, 16'd64303, 16'd49987, 16'd1306, 16'd32458, 16'd48612, 16'd29502, 16'd23554, 16'd53384, 16'd35965, 16'd13214, 16'd50424});
	test_expansion(128'he39cb24989659a064cb2de555c9e9d49, {16'd48527, 16'd15280, 16'd13627, 16'd27880, 16'd6293, 16'd30449, 16'd1997, 16'd32447, 16'd33518, 16'd45286, 16'd52828, 16'd1791, 16'd55187, 16'd62989, 16'd59140, 16'd745, 16'd57481, 16'd19027, 16'd46324, 16'd22104, 16'd32115, 16'd689, 16'd12566, 16'd50567, 16'd27984, 16'd31267});
	test_expansion(128'h26ffc588ad836b29fa0f613d0938c457, {16'd9641, 16'd38342, 16'd28634, 16'd3552, 16'd11974, 16'd5441, 16'd3439, 16'd36648, 16'd37511, 16'd18950, 16'd65144, 16'd24909, 16'd18591, 16'd60863, 16'd62888, 16'd10353, 16'd17642, 16'd28237, 16'd10163, 16'd61316, 16'd50319, 16'd10945, 16'd18037, 16'd53348, 16'd23125, 16'd63401});
	test_expansion(128'h63a28aa652fe3790b6b65db7e93fc6ae, {16'd14091, 16'd5840, 16'd60706, 16'd7570, 16'd25973, 16'd26177, 16'd5662, 16'd30621, 16'd3914, 16'd41305, 16'd32211, 16'd62387, 16'd44044, 16'd35887, 16'd17780, 16'd62143, 16'd18135, 16'd217, 16'd37657, 16'd12991, 16'd24025, 16'd1345, 16'd61052, 16'd55096, 16'd60087, 16'd29909});
	test_expansion(128'hed250515a5f2e52a3ff4c1bce3257f53, {16'd7553, 16'd17415, 16'd59664, 16'd38781, 16'd61218, 16'd19212, 16'd42071, 16'd1728, 16'd10806, 16'd64419, 16'd56291, 16'd54442, 16'd31455, 16'd40226, 16'd22000, 16'd24662, 16'd2770, 16'd47333, 16'd6994, 16'd22502, 16'd46236, 16'd50885, 16'd35796, 16'd40771, 16'd38421, 16'd44599});
	test_expansion(128'hb60289447cf2c3c26a118fc22fa37ed7, {16'd52587, 16'd26618, 16'd24963, 16'd22042, 16'd3424, 16'd15329, 16'd10591, 16'd46348, 16'd29683, 16'd33543, 16'd41848, 16'd29656, 16'd39085, 16'd62809, 16'd43089, 16'd22685, 16'd57455, 16'd41137, 16'd28407, 16'd24977, 16'd60026, 16'd16454, 16'd48777, 16'd56982, 16'd62779, 16'd31129});
	test_expansion(128'h07516c23059519e0e25106cc565050b0, {16'd12539, 16'd45800, 16'd55498, 16'd20928, 16'd21060, 16'd47909, 16'd61377, 16'd21630, 16'd56031, 16'd44075, 16'd46050, 16'd4582, 16'd4504, 16'd19496, 16'd41526, 16'd22483, 16'd19452, 16'd50829, 16'd14642, 16'd251, 16'd33338, 16'd64730, 16'd57555, 16'd8718, 16'd2811, 16'd60865});
	test_expansion(128'h5bcad377b420f980e6d1f151aa7df889, {16'd23182, 16'd2345, 16'd604, 16'd49624, 16'd52497, 16'd19717, 16'd58677, 16'd61548, 16'd43810, 16'd44448, 16'd37395, 16'd46782, 16'd34655, 16'd4507, 16'd27075, 16'd2405, 16'd65294, 16'd19871, 16'd36385, 16'd13155, 16'd28740, 16'd34363, 16'd35518, 16'd11491, 16'd111, 16'd60519});
	test_expansion(128'h985cfcfaf90caa3b701fabbe2534141e, {16'd48218, 16'd65454, 16'd17570, 16'd25299, 16'd21312, 16'd23857, 16'd62928, 16'd25093, 16'd41401, 16'd47214, 16'd33921, 16'd41586, 16'd56804, 16'd18770, 16'd30912, 16'd43455, 16'd15181, 16'd63586, 16'd24772, 16'd1015, 16'd50224, 16'd57171, 16'd60522, 16'd50302, 16'd52276, 16'd61134});
	test_expansion(128'h07d11e3661f81e01386a75914e24dd36, {16'd53876, 16'd6811, 16'd61565, 16'd49396, 16'd22586, 16'd12408, 16'd3908, 16'd45692, 16'd37820, 16'd45622, 16'd39813, 16'd3958, 16'd37969, 16'd18684, 16'd5820, 16'd7069, 16'd61004, 16'd23239, 16'd10842, 16'd51812, 16'd9131, 16'd47209, 16'd30417, 16'd31556, 16'd33173, 16'd18634});
	test_expansion(128'ha3cb99c735e7a45e692f4c5fa5d4b1f3, {16'd59974, 16'd4135, 16'd4492, 16'd5302, 16'd12956, 16'd20419, 16'd11993, 16'd58192, 16'd20707, 16'd17210, 16'd54122, 16'd26927, 16'd59585, 16'd63049, 16'd39730, 16'd61396, 16'd3095, 16'd47896, 16'd12733, 16'd21484, 16'd7916, 16'd55731, 16'd55260, 16'd56977, 16'd27701, 16'd14182});
	test_expansion(128'hec2c2acdb99ab0460b36736d746d72ad, {16'd42475, 16'd10212, 16'd57566, 16'd65298, 16'd21898, 16'd19179, 16'd803, 16'd34584, 16'd44656, 16'd62609, 16'd43062, 16'd11768, 16'd51349, 16'd31614, 16'd4203, 16'd3587, 16'd60284, 16'd51118, 16'd16197, 16'd21604, 16'd64597, 16'd10957, 16'd1890, 16'd30222, 16'd8416, 16'd45485});
	test_expansion(128'h40518da41b15494f6aa4e71f0cd11288, {16'd27586, 16'd64437, 16'd50156, 16'd52406, 16'd9442, 16'd34084, 16'd27286, 16'd29152, 16'd15802, 16'd23094, 16'd32131, 16'd27491, 16'd17907, 16'd18496, 16'd48666, 16'd22922, 16'd9078, 16'd40695, 16'd11020, 16'd20039, 16'd37547, 16'd25801, 16'd18221, 16'd7616, 16'd28585, 16'd24116});
	test_expansion(128'h7df1158e65499117a8f48394513eee91, {16'd34571, 16'd43894, 16'd50879, 16'd9592, 16'd39318, 16'd48057, 16'd47863, 16'd42056, 16'd47609, 16'd42960, 16'd19380, 16'd12183, 16'd20955, 16'd59165, 16'd29064, 16'd39235, 16'd27430, 16'd59421, 16'd34914, 16'd9911, 16'd36975, 16'd31302, 16'd22164, 16'd59712, 16'd30136, 16'd15680});
	test_expansion(128'h7f0becc0da9c5ac82d98367d30b09d7d, {16'd8538, 16'd1210, 16'd12681, 16'd42749, 16'd56048, 16'd22926, 16'd52459, 16'd33024, 16'd45125, 16'd52614, 16'd29162, 16'd55968, 16'd44288, 16'd24901, 16'd57526, 16'd61363, 16'd15057, 16'd37563, 16'd64832, 16'd3428, 16'd21215, 16'd18566, 16'd47536, 16'd45739, 16'd42147, 16'd5152});
	test_expansion(128'h3f69cc3ac925811690a464c153778ed5, {16'd8024, 16'd26971, 16'd41179, 16'd3989, 16'd19424, 16'd58623, 16'd28687, 16'd53162, 16'd19870, 16'd63763, 16'd32002, 16'd29027, 16'd28100, 16'd14625, 16'd58824, 16'd9376, 16'd56586, 16'd14185, 16'd36370, 16'd34339, 16'd52408, 16'd60460, 16'd38638, 16'd42188, 16'd34277, 16'd10709});
	test_expansion(128'hbb2708d9c23c0c2ac76db2663d82998d, {16'd23255, 16'd31052, 16'd47162, 16'd6374, 16'd31416, 16'd60690, 16'd21154, 16'd41714, 16'd60416, 16'd38789, 16'd63715, 16'd60779, 16'd50801, 16'd39803, 16'd48233, 16'd14147, 16'd55231, 16'd9036, 16'd45509, 16'd59677, 16'd2266, 16'd63177, 16'd25924, 16'd40188, 16'd37369, 16'd12186});
	test_expansion(128'h6b30c326b0ec7d01e5d20625233612d9, {16'd36388, 16'd17554, 16'd6914, 16'd16225, 16'd44123, 16'd35912, 16'd9227, 16'd15948, 16'd27970, 16'd36408, 16'd29254, 16'd22363, 16'd56174, 16'd6036, 16'd63992, 16'd50450, 16'd22569, 16'd21906, 16'd23183, 16'd47019, 16'd18093, 16'd17875, 16'd59996, 16'd21919, 16'd14640, 16'd49707});
	test_expansion(128'h5e02ac15711438eed9fc1917a50782ac, {16'd25927, 16'd5366, 16'd2752, 16'd58613, 16'd27380, 16'd65396, 16'd64296, 16'd3131, 16'd49803, 16'd28963, 16'd54908, 16'd53873, 16'd16862, 16'd58094, 16'd19107, 16'd5274, 16'd45043, 16'd63961, 16'd50528, 16'd51635, 16'd60913, 16'd6274, 16'd5231, 16'd26783, 16'd37736, 16'd9018});
	test_expansion(128'h0480e023dbff1af9e63a84818eb7258b, {16'd2408, 16'd35205, 16'd10966, 16'd8237, 16'd6971, 16'd64019, 16'd12861, 16'd33252, 16'd26334, 16'd40551, 16'd49264, 16'd10070, 16'd31533, 16'd13658, 16'd44655, 16'd19032, 16'd6798, 16'd43503, 16'd45977, 16'd16433, 16'd62660, 16'd27254, 16'd23981, 16'd51911, 16'd17782, 16'd6068});
	test_expansion(128'h2e62747beece621f8616f2aebcec8dde, {16'd12640, 16'd51199, 16'd28910, 16'd16320, 16'd13659, 16'd27796, 16'd43958, 16'd58098, 16'd16849, 16'd61544, 16'd43423, 16'd52480, 16'd49988, 16'd12179, 16'd17438, 16'd58719, 16'd30715, 16'd12602, 16'd17876, 16'd29484, 16'd11715, 16'd16246, 16'd64389, 16'd6537, 16'd24609, 16'd11545});
	test_expansion(128'hb1f71f0fc97d31252ef3f5fd7b8583d6, {16'd51597, 16'd57108, 16'd50427, 16'd33101, 16'd16119, 16'd30979, 16'd10608, 16'd21580, 16'd40552, 16'd3623, 16'd38774, 16'd48129, 16'd5968, 16'd26654, 16'd41097, 16'd48282, 16'd11900, 16'd61067, 16'd42860, 16'd25616, 16'd21377, 16'd25642, 16'd9121, 16'd17508, 16'd2745, 16'd31024});
	test_expansion(128'h6a767996f6ca22b191e5fa094c6bfe6d, {16'd21440, 16'd19373, 16'd52147, 16'd2114, 16'd18910, 16'd60969, 16'd9301, 16'd47539, 16'd35836, 16'd64093, 16'd15460, 16'd59939, 16'd34088, 16'd36664, 16'd54835, 16'd27944, 16'd20604, 16'd40933, 16'd63075, 16'd1672, 16'd34412, 16'd14945, 16'd5502, 16'd57370, 16'd35267, 16'd16973});
	test_expansion(128'ha608394f38bf8b0d7e70ad685c80d5a4, {16'd11004, 16'd18178, 16'd10608, 16'd25504, 16'd22456, 16'd48264, 16'd5830, 16'd51872, 16'd8728, 16'd20142, 16'd12400, 16'd41962, 16'd9500, 16'd22438, 16'd17894, 16'd54723, 16'd20900, 16'd28672, 16'd41759, 16'd42246, 16'd62900, 16'd8116, 16'd28578, 16'd5346, 16'd35024, 16'd49472});
	test_expansion(128'he0109df4c60adc6b64bf2c00d07e5b9d, {16'd54484, 16'd64284, 16'd31826, 16'd18891, 16'd54853, 16'd28433, 16'd50512, 16'd36997, 16'd35507, 16'd31121, 16'd23104, 16'd40459, 16'd62460, 16'd12115, 16'd46929, 16'd196, 16'd28473, 16'd33659, 16'd24870, 16'd46247, 16'd22187, 16'd54130, 16'd53873, 16'd7318, 16'd60342, 16'd12181});
	test_expansion(128'h43547cfefb49a080fd4e5c442714fa4f, {16'd3060, 16'd39805, 16'd25883, 16'd31563, 16'd21619, 16'd454, 16'd45232, 16'd37275, 16'd54601, 16'd47711, 16'd14905, 16'd27396, 16'd49529, 16'd22171, 16'd29932, 16'd20898, 16'd51034, 16'd7685, 16'd48905, 16'd49363, 16'd19032, 16'd63694, 16'd36518, 16'd21114, 16'd122, 16'd20210});
	test_expansion(128'hf18f6450477a6db1ea671f0140abde6e, {16'd10451, 16'd56981, 16'd64291, 16'd11885, 16'd46931, 16'd23935, 16'd22522, 16'd34200, 16'd433, 16'd19487, 16'd35604, 16'd18811, 16'd29824, 16'd20330, 16'd27036, 16'd35143, 16'd54999, 16'd26523, 16'd51198, 16'd33212, 16'd30007, 16'd35734, 16'd53154, 16'd19496, 16'd1774, 16'd61028});
	test_expansion(128'h74a2edfdeb092574fb720db9abf13129, {16'd29961, 16'd54638, 16'd44352, 16'd43397, 16'd22597, 16'd36030, 16'd36811, 16'd50101, 16'd62731, 16'd44774, 16'd23447, 16'd38575, 16'd38495, 16'd22122, 16'd8924, 16'd10912, 16'd23491, 16'd23294, 16'd9080, 16'd28755, 16'd25396, 16'd51482, 16'd3446, 16'd48141, 16'd44549, 16'd48588});
	test_expansion(128'hcbbf7ff69ed9e37f6525095ce9ec8712, {16'd39946, 16'd27849, 16'd38851, 16'd41827, 16'd4698, 16'd53580, 16'd23301, 16'd36750, 16'd59428, 16'd40707, 16'd54152, 16'd5224, 16'd4994, 16'd14868, 16'd62440, 16'd24179, 16'd55894, 16'd54870, 16'd32320, 16'd40668, 16'd15640, 16'd4897, 16'd23822, 16'd39751, 16'd34774, 16'd24842});
	test_expansion(128'h7cebbc3124767e3c82e7594792e835c5, {16'd46477, 16'd62459, 16'd2997, 16'd4416, 16'd6406, 16'd64278, 16'd20908, 16'd19584, 16'd27693, 16'd30669, 16'd61102, 16'd41232, 16'd23377, 16'd28798, 16'd23833, 16'd24664, 16'd60291, 16'd54879, 16'd44753, 16'd44624, 16'd46728, 16'd49052, 16'd12306, 16'd27894, 16'd65355, 16'd278});
	test_expansion(128'hc54eb8d7e4cb0b130173839f537e418a, {16'd47045, 16'd17119, 16'd30391, 16'd20934, 16'd20377, 16'd13334, 16'd51738, 16'd28025, 16'd6364, 16'd59234, 16'd22428, 16'd15059, 16'd43236, 16'd14723, 16'd8918, 16'd21497, 16'd24710, 16'd25113, 16'd14843, 16'd18289, 16'd55863, 16'd53107, 16'd18366, 16'd21409, 16'd38118, 16'd49748});
	test_expansion(128'h606c3d0d59f32b27ac115ca0a745ea34, {16'd34231, 16'd60619, 16'd65442, 16'd47421, 16'd40055, 16'd59650, 16'd12433, 16'd65246, 16'd48421, 16'd25624, 16'd31225, 16'd1925, 16'd27872, 16'd26298, 16'd45971, 16'd55189, 16'd26940, 16'd62541, 16'd13545, 16'd34190, 16'd29199, 16'd22318, 16'd8196, 16'd11876, 16'd54355, 16'd48329});
	test_expansion(128'h2eed6009b17fbcf6b72498c668a2eaa2, {16'd19226, 16'd64504, 16'd33903, 16'd52153, 16'd64970, 16'd27474, 16'd42939, 16'd15163, 16'd9612, 16'd26264, 16'd65064, 16'd40895, 16'd33201, 16'd48085, 16'd40451, 16'd17519, 16'd54521, 16'd1388, 16'd52751, 16'd39586, 16'd41809, 16'd40978, 16'd54238, 16'd11716, 16'd59081, 16'd30446});
	test_expansion(128'h606e0297396614740a2113719d6bba64, {16'd58660, 16'd54650, 16'd55654, 16'd25506, 16'd9754, 16'd20915, 16'd64404, 16'd1169, 16'd9606, 16'd24948, 16'd47352, 16'd29328, 16'd1068, 16'd48785, 16'd19131, 16'd4648, 16'd48110, 16'd30404, 16'd5862, 16'd21792, 16'd21691, 16'd19512, 16'd65497, 16'd46135, 16'd64348, 16'd34902});
	test_expansion(128'ha19c609c41b8fbddd00ad1702dbeee1d, {16'd46061, 16'd63178, 16'd58733, 16'd42653, 16'd3784, 16'd41084, 16'd3454, 16'd9541, 16'd49378, 16'd5043, 16'd8747, 16'd47501, 16'd12274, 16'd12057, 16'd503, 16'd3356, 16'd37036, 16'd26875, 16'd18954, 16'd12050, 16'd50957, 16'd57182, 16'd35649, 16'd31042, 16'd27072, 16'd60197});
	test_expansion(128'h8b6be94e1a57c879ea1f09293b5ad395, {16'd12674, 16'd21379, 16'd18302, 16'd9323, 16'd11070, 16'd10373, 16'd57684, 16'd55384, 16'd62443, 16'd37277, 16'd12652, 16'd26046, 16'd7966, 16'd44874, 16'd3063, 16'd32178, 16'd10000, 16'd45244, 16'd32904, 16'd59807, 16'd52911, 16'd8769, 16'd19691, 16'd54237, 16'd5192, 16'd22515});
	test_expansion(128'h9801a159c011679ec01af170970ba5c7, {16'd21945, 16'd16308, 16'd51424, 16'd6657, 16'd11254, 16'd50552, 16'd32022, 16'd57045, 16'd49379, 16'd17013, 16'd3171, 16'd42873, 16'd10526, 16'd65191, 16'd61120, 16'd24834, 16'd31582, 16'd33942, 16'd57629, 16'd61119, 16'd47321, 16'd4214, 16'd47691, 16'd13727, 16'd35697, 16'd56003});
	test_expansion(128'h4ce7a554b0158f61d27d072dcc5fc907, {16'd10181, 16'd31765, 16'd20559, 16'd50488, 16'd20230, 16'd55119, 16'd62904, 16'd12480, 16'd62155, 16'd56648, 16'd19690, 16'd28442, 16'd3419, 16'd42799, 16'd37912, 16'd62138, 16'd47536, 16'd36159, 16'd53776, 16'd57848, 16'd42521, 16'd56560, 16'd8704, 16'd22984, 16'd56292, 16'd22924});
	test_expansion(128'hd45268d6f43f4e3570297e00f5373477, {16'd34288, 16'd50773, 16'd15893, 16'd18711, 16'd9888, 16'd45186, 16'd57662, 16'd11755, 16'd64984, 16'd62917, 16'd24831, 16'd34058, 16'd536, 16'd20963, 16'd1864, 16'd10349, 16'd47600, 16'd17813, 16'd859, 16'd9268, 16'd53486, 16'd30191, 16'd62082, 16'd1950, 16'd40492, 16'd35127});
	test_expansion(128'h79acfaa1a0773d54e6226979a318531a, {16'd18752, 16'd55084, 16'd57315, 16'd18435, 16'd31257, 16'd53008, 16'd29185, 16'd19405, 16'd46495, 16'd13032, 16'd15162, 16'd19844, 16'd5888, 16'd15205, 16'd25250, 16'd14950, 16'd59337, 16'd36901, 16'd27919, 16'd58615, 16'd51021, 16'd18899, 16'd32922, 16'd23233, 16'd28236, 16'd31860});
	test_expansion(128'h11a347f92cfb3fc4ceab9785d9f49895, {16'd65022, 16'd37420, 16'd52711, 16'd42703, 16'd9783, 16'd25547, 16'd11220, 16'd16987, 16'd5947, 16'd56042, 16'd64122, 16'd49222, 16'd53989, 16'd23859, 16'd61312, 16'd27386, 16'd2421, 16'd37961, 16'd61030, 16'd47149, 16'd61073, 16'd50729, 16'd51642, 16'd57893, 16'd57943, 16'd35746});
	test_expansion(128'h3469415082bdb89f4835942162f452d9, {16'd1626, 16'd46513, 16'd5770, 16'd11037, 16'd57822, 16'd18888, 16'd37497, 16'd52380, 16'd62163, 16'd58861, 16'd9394, 16'd19903, 16'd23667, 16'd25197, 16'd11850, 16'd49379, 16'd14838, 16'd36868, 16'd10298, 16'd54658, 16'd55200, 16'd56805, 16'd38725, 16'd22391, 16'd25212, 16'd61598});
	test_expansion(128'hcfe286058540dcffa68a75c8569b1d1b, {16'd18819, 16'd34986, 16'd45931, 16'd31468, 16'd40320, 16'd27070, 16'd46559, 16'd41270, 16'd53255, 16'd18481, 16'd34289, 16'd56346, 16'd59969, 16'd5731, 16'd16244, 16'd19190, 16'd27069, 16'd15395, 16'd26095, 16'd24117, 16'd37397, 16'd39581, 16'd47823, 16'd22229, 16'd54759, 16'd23830});
	test_expansion(128'hb5da2f3c7ba715c560b30ef1fd2a71f6, {16'd53909, 16'd57499, 16'd58109, 16'd64815, 16'd26849, 16'd36965, 16'd30663, 16'd32445, 16'd51541, 16'd34851, 16'd19935, 16'd30445, 16'd54440, 16'd8503, 16'd51264, 16'd14091, 16'd4528, 16'd35758, 16'd64512, 16'd62739, 16'd14398, 16'd12840, 16'd25272, 16'd22304, 16'd5286, 16'd27203});
	test_expansion(128'h25d63d700d21677c0db2f81a57013676, {16'd43779, 16'd64764, 16'd10158, 16'd65416, 16'd32069, 16'd4095, 16'd14380, 16'd37103, 16'd121, 16'd13293, 16'd19795, 16'd49786, 16'd59035, 16'd15404, 16'd44586, 16'd28390, 16'd29462, 16'd30717, 16'd21683, 16'd20146, 16'd40259, 16'd19765, 16'd52054, 16'd53303, 16'd47816, 16'd29486});
	test_expansion(128'h94a8912e038690468a722ef02643fc54, {16'd62587, 16'd44861, 16'd47491, 16'd10240, 16'd15888, 16'd60254, 16'd21226, 16'd7000, 16'd21950, 16'd11471, 16'd12772, 16'd3321, 16'd27888, 16'd43141, 16'd38021, 16'd14017, 16'd65120, 16'd25455, 16'd37283, 16'd45550, 16'd22253, 16'd8393, 16'd18121, 16'd52765, 16'd25022, 16'd52797});
	test_expansion(128'hf1ba7aab02c6c8ecc2118730b65894aa, {16'd39789, 16'd24408, 16'd16868, 16'd27614, 16'd37721, 16'd45082, 16'd19524, 16'd52224, 16'd58055, 16'd48886, 16'd51851, 16'd60013, 16'd48089, 16'd24373, 16'd37370, 16'd3542, 16'd62900, 16'd37169, 16'd39020, 16'd13203, 16'd63066, 16'd28795, 16'd16097, 16'd48851, 16'd34551, 16'd14037});
	test_expansion(128'h0194e636c1e2e9f34db28d2b7ff6df99, {16'd35428, 16'd45206, 16'd25197, 16'd47085, 16'd1401, 16'd23526, 16'd13664, 16'd27853, 16'd49578, 16'd59390, 16'd56734, 16'd64528, 16'd20892, 16'd56552, 16'd48819, 16'd60869, 16'd10255, 16'd17587, 16'd36490, 16'd11057, 16'd54584, 16'd27281, 16'd63241, 16'd11376, 16'd50704, 16'd30585});
	test_expansion(128'hc7cd07452d05d0d8458cecd72549c1f2, {16'd32998, 16'd39268, 16'd1460, 16'd2985, 16'd27745, 16'd53319, 16'd46132, 16'd25403, 16'd11361, 16'd19179, 16'd37370, 16'd53726, 16'd18608, 16'd24800, 16'd56369, 16'd12413, 16'd34977, 16'd58882, 16'd30047, 16'd44925, 16'd24641, 16'd41776, 16'd40439, 16'd17487, 16'd58305, 16'd57561});
	test_expansion(128'h0367aadb62769f8df263a365ffaa7d43, {16'd36952, 16'd27815, 16'd65427, 16'd59250, 16'd24180, 16'd8324, 16'd15791, 16'd25270, 16'd60706, 16'd7612, 16'd45650, 16'd48935, 16'd61967, 16'd32190, 16'd19209, 16'd61750, 16'd14988, 16'd1856, 16'd6168, 16'd21027, 16'd39426, 16'd15389, 16'd61617, 16'd48851, 16'd10291, 16'd3130});
	test_expansion(128'h837c09b64a90e07436d679ad70b60564, {16'd55019, 16'd7251, 16'd59613, 16'd33739, 16'd64391, 16'd46806, 16'd39567, 16'd40687, 16'd43325, 16'd28254, 16'd1877, 16'd24796, 16'd50900, 16'd4867, 16'd8802, 16'd49029, 16'd2318, 16'd14805, 16'd46323, 16'd9705, 16'd1496, 16'd49924, 16'd14275, 16'd48456, 16'd16251, 16'd7253});
	test_expansion(128'h2296399c34ab4def006a96bc06ed8c69, {16'd33063, 16'd51717, 16'd3985, 16'd26455, 16'd37262, 16'd54010, 16'd43088, 16'd55667, 16'd42758, 16'd11320, 16'd43733, 16'd33625, 16'd28154, 16'd11672, 16'd43396, 16'd60454, 16'd23462, 16'd30398, 16'd33509, 16'd39863, 16'd2620, 16'd40737, 16'd60522, 16'd55291, 16'd50563, 16'd40534});
	test_expansion(128'h9fa4732cf873281ed0044af4a9791bd9, {16'd12606, 16'd52341, 16'd27021, 16'd38447, 16'd1162, 16'd30450, 16'd23714, 16'd61602, 16'd17796, 16'd22441, 16'd16599, 16'd14304, 16'd53942, 16'd27053, 16'd17479, 16'd15302, 16'd46816, 16'd31373, 16'd45305, 16'd9067, 16'd7721, 16'd42276, 16'd12381, 16'd28514, 16'd28495, 16'd9692});
	test_expansion(128'h8a0a8239fa9b5378ddb9f42237e113f1, {16'd43187, 16'd3770, 16'd41154, 16'd63867, 16'd58361, 16'd56568, 16'd42294, 16'd54514, 16'd22483, 16'd55466, 16'd22679, 16'd8483, 16'd29645, 16'd27233, 16'd5558, 16'd59904, 16'd34969, 16'd17845, 16'd24758, 16'd55681, 16'd25465, 16'd50536, 16'd52164, 16'd20465, 16'd13563, 16'd62885});
	test_expansion(128'h7078d7ccd8572a74757bb50d11eae576, {16'd4142, 16'd2078, 16'd44070, 16'd8138, 16'd28234, 16'd38230, 16'd2771, 16'd23617, 16'd18555, 16'd37908, 16'd52911, 16'd27505, 16'd22501, 16'd55299, 16'd10360, 16'd5512, 16'd30508, 16'd51568, 16'd63717, 16'd11247, 16'd60012, 16'd55648, 16'd61899, 16'd30434, 16'd54418, 16'd38243});
	test_expansion(128'h1c05fca39b1ac8ab640be8fecb9c7f85, {16'd40401, 16'd27461, 16'd38870, 16'd34173, 16'd53031, 16'd52332, 16'd22752, 16'd26845, 16'd3033, 16'd2283, 16'd24179, 16'd53951, 16'd44755, 16'd12315, 16'd14612, 16'd34547, 16'd4756, 16'd19741, 16'd22254, 16'd55962, 16'd14534, 16'd22170, 16'd63189, 16'd34667, 16'd60584, 16'd9751});
	test_expansion(128'he903e8078cbea8a589e17f65c7ef5321, {16'd65068, 16'd33158, 16'd13765, 16'd51554, 16'd58069, 16'd50563, 16'd42787, 16'd47815, 16'd55269, 16'd61869, 16'd62255, 16'd37711, 16'd37807, 16'd32596, 16'd16409, 16'd10173, 16'd64235, 16'd58481, 16'd64434, 16'd46812, 16'd38755, 16'd13638, 16'd41488, 16'd21984, 16'd64369, 16'd36632});
	test_expansion(128'he754e6b2ee5e7b67e79bd61aa18f6f23, {16'd3327, 16'd7636, 16'd63781, 16'd55383, 16'd15828, 16'd45877, 16'd36677, 16'd47661, 16'd13384, 16'd63200, 16'd31190, 16'd61319, 16'd15066, 16'd19122, 16'd27468, 16'd55109, 16'd21298, 16'd33330, 16'd921, 16'd33917, 16'd23485, 16'd9058, 16'd34144, 16'd8607, 16'd15573, 16'd27413});
	test_expansion(128'hf427499c5c950371bd7b1297571f40ab, {16'd62190, 16'd41461, 16'd48126, 16'd40116, 16'd49835, 16'd45488, 16'd22079, 16'd6744, 16'd14673, 16'd23377, 16'd49650, 16'd28677, 16'd35497, 16'd46918, 16'd25967, 16'd33537, 16'd36697, 16'd15666, 16'd56778, 16'd27573, 16'd40304, 16'd52566, 16'd19731, 16'd42014, 16'd10441, 16'd64855});
	test_expansion(128'h4c5f2a4e483a2fd3e364b5fd037cca76, {16'd9887, 16'd61105, 16'd54745, 16'd10977, 16'd5221, 16'd52641, 16'd14127, 16'd54387, 16'd50997, 16'd51443, 16'd37332, 16'd51456, 16'd46052, 16'd32759, 16'd34220, 16'd1554, 16'd20972, 16'd51700, 16'd4080, 16'd21732, 16'd34850, 16'd38118, 16'd29027, 16'd29411, 16'd18014, 16'd62417});
	test_expansion(128'hdbec50f6cb9918574c16a72d65bdea28, {16'd17872, 16'd63222, 16'd35374, 16'd25706, 16'd16921, 16'd45833, 16'd18232, 16'd63971, 16'd63738, 16'd35477, 16'd17990, 16'd7389, 16'd63083, 16'd37272, 16'd38930, 16'd3847, 16'd62532, 16'd25652, 16'd14105, 16'd52565, 16'd58780, 16'd47430, 16'd27056, 16'd21635, 16'd52882, 16'd38622});
	test_expansion(128'h797bf91b0b992d1e53d637024b7df855, {16'd48441, 16'd718, 16'd52755, 16'd23539, 16'd46996, 16'd57553, 16'd19760, 16'd32149, 16'd25028, 16'd4390, 16'd40860, 16'd14708, 16'd26297, 16'd5750, 16'd31364, 16'd13363, 16'd39195, 16'd53077, 16'd11611, 16'd54750, 16'd32068, 16'd11213, 16'd46427, 16'd21359, 16'd59785, 16'd22562});
	test_expansion(128'h673304e435dd6e409c1f62c1e75e380e, {16'd60704, 16'd18742, 16'd57469, 16'd34360, 16'd55873, 16'd37263, 16'd51181, 16'd5313, 16'd41108, 16'd745, 16'd39257, 16'd14, 16'd17833, 16'd9727, 16'd57236, 16'd43832, 16'd32228, 16'd32596, 16'd28771, 16'd61144, 16'd64725, 16'd30627, 16'd38782, 16'd49052, 16'd13133, 16'd53720});
	test_expansion(128'hb5296eebdb4fefe2292252a04a23bd5a, {16'd31726, 16'd23416, 16'd48995, 16'd42922, 16'd26616, 16'd45689, 16'd30433, 16'd36914, 16'd13972, 16'd59343, 16'd27988, 16'd27781, 16'd44754, 16'd43690, 16'd37060, 16'd46664, 16'd30616, 16'd60966, 16'd49820, 16'd48101, 16'd8933, 16'd9655, 16'd62981, 16'd5583, 16'd21554, 16'd4087});
	test_expansion(128'he41f383cbdccbcd2d34efb776ed26f91, {16'd18131, 16'd22411, 16'd28158, 16'd58258, 16'd19772, 16'd49018, 16'd59447, 16'd30768, 16'd25877, 16'd2486, 16'd53582, 16'd38727, 16'd35955, 16'd28197, 16'd14024, 16'd36500, 16'd40629, 16'd46182, 16'd30751, 16'd18332, 16'd2258, 16'd27354, 16'd29873, 16'd50062, 16'd19200, 16'd40074});
	test_expansion(128'hc0a659874f4e5a6acb20776f991ea792, {16'd31646, 16'd53699, 16'd23278, 16'd24187, 16'd19144, 16'd16127, 16'd56734, 16'd47593, 16'd49492, 16'd17222, 16'd23120, 16'd22341, 16'd10643, 16'd39336, 16'd64031, 16'd30339, 16'd32991, 16'd8997, 16'd20322, 16'd25874, 16'd30612, 16'd53039, 16'd30380, 16'd25694, 16'd35885, 16'd62568});
	test_expansion(128'hcf1df7cc362b2f78df6c8e5c7521b67c, {16'd6405, 16'd25002, 16'd13224, 16'd39356, 16'd29486, 16'd24756, 16'd41229, 16'd13871, 16'd10757, 16'd50098, 16'd58959, 16'd8184, 16'd19904, 16'd35879, 16'd45270, 16'd26860, 16'd45933, 16'd9918, 16'd41407, 16'd20861, 16'd63929, 16'd18339, 16'd41528, 16'd36635, 16'd4447, 16'd46110});
	test_expansion(128'h69e1c5e3886697a720f88ead02882d88, {16'd27195, 16'd56648, 16'd1523, 16'd53194, 16'd10724, 16'd5219, 16'd34682, 16'd51277, 16'd637, 16'd20105, 16'd41891, 16'd42387, 16'd64336, 16'd3901, 16'd7523, 16'd50906, 16'd17100, 16'd56530, 16'd54767, 16'd16129, 16'd28637, 16'd35070, 16'd38287, 16'd54659, 16'd54776, 16'd23139});
	test_expansion(128'hb1ce42d4be9d528cd0be16c9c799cc78, {16'd63727, 16'd14246, 16'd58026, 16'd49395, 16'd36981, 16'd39728, 16'd42106, 16'd24926, 16'd44792, 16'd35921, 16'd47156, 16'd37387, 16'd40017, 16'd35648, 16'd38845, 16'd14444, 16'd13706, 16'd62627, 16'd55758, 16'd23646, 16'd11756, 16'd62902, 16'd33491, 16'd29348, 16'd51189, 16'd22573});
	test_expansion(128'hc130609af48e8abfbc00e51e5a4fc411, {16'd36000, 16'd22721, 16'd55756, 16'd40896, 16'd19205, 16'd61746, 16'd62848, 16'd33949, 16'd57604, 16'd63092, 16'd4961, 16'd28335, 16'd23476, 16'd7486, 16'd15547, 16'd53524, 16'd19093, 16'd27055, 16'd60519, 16'd65114, 16'd34040, 16'd4539, 16'd14117, 16'd42967, 16'd55323, 16'd38565});
	test_expansion(128'hf3d1239751f55864c1d86a5f1b73eb26, {16'd12314, 16'd27774, 16'd5868, 16'd19783, 16'd63690, 16'd17570, 16'd13596, 16'd49994, 16'd46337, 16'd4307, 16'd41603, 16'd35, 16'd34450, 16'd64048, 16'd50166, 16'd6284, 16'd23805, 16'd39330, 16'd236, 16'd60127, 16'd59991, 16'd12085, 16'd2390, 16'd16461, 16'd2696, 16'd23518});
	test_expansion(128'h706d8b5531891cd3c74a54325baf5038, {16'd26439, 16'd65155, 16'd26305, 16'd21998, 16'd33832, 16'd43406, 16'd55400, 16'd22178, 16'd33, 16'd15139, 16'd40170, 16'd49130, 16'd20621, 16'd61007, 16'd58002, 16'd59674, 16'd36812, 16'd63611, 16'd12347, 16'd23815, 16'd34284, 16'd64116, 16'd53898, 16'd24531, 16'd50192, 16'd1137});
	test_expansion(128'hb9068a04c7a3eb77b88ede833b681e46, {16'd62337, 16'd12397, 16'd33829, 16'd51547, 16'd20477, 16'd31437, 16'd13271, 16'd21819, 16'd53259, 16'd28770, 16'd55217, 16'd34121, 16'd16150, 16'd13869, 16'd27247, 16'd42865, 16'd9173, 16'd4629, 16'd54467, 16'd64520, 16'd34607, 16'd39874, 16'd58353, 16'd59927, 16'd31850, 16'd53416});
	test_expansion(128'hfa2a6081fa22274d0f8a1ae28bd3d4a4, {16'd29303, 16'd35344, 16'd60178, 16'd14762, 16'd29739, 16'd42553, 16'd46917, 16'd26744, 16'd39968, 16'd47527, 16'd13739, 16'd9258, 16'd18261, 16'd34150, 16'd4735, 16'd62233, 16'd17234, 16'd51200, 16'd20599, 16'd25165, 16'd64530, 16'd23948, 16'd29275, 16'd30401, 16'd6288, 16'd40048});
	test_expansion(128'he5c8b4ea692e6a5c2cffcdc28be4296d, {16'd48587, 16'd54934, 16'd63668, 16'd58807, 16'd51980, 16'd19757, 16'd43017, 16'd60739, 16'd63657, 16'd18886, 16'd37754, 16'd24834, 16'd45741, 16'd45814, 16'd63646, 16'd37628, 16'd45394, 16'd53505, 16'd7989, 16'd56927, 16'd55896, 16'd33066, 16'd63375, 16'd59953, 16'd48346, 16'd48606});
	test_expansion(128'h4b57de2e1567fb72bdc396259faa347d, {16'd18419, 16'd36828, 16'd51868, 16'd5927, 16'd49827, 16'd6949, 16'd46539, 16'd20223, 16'd57123, 16'd51162, 16'd50394, 16'd34924, 16'd2164, 16'd63572, 16'd27000, 16'd37550, 16'd56906, 16'd44634, 16'd45193, 16'd51014, 16'd53459, 16'd43959, 16'd13755, 16'd63192, 16'd15548, 16'd14427});
	test_expansion(128'h9141c471717f36cf0bc1593d82a09814, {16'd63419, 16'd5669, 16'd48787, 16'd54858, 16'd13266, 16'd4180, 16'd4443, 16'd38579, 16'd12068, 16'd2561, 16'd27822, 16'd12659, 16'd45542, 16'd26469, 16'd42562, 16'd33621, 16'd54187, 16'd8653, 16'd5198, 16'd23205, 16'd56513, 16'd13124, 16'd48293, 16'd31296, 16'd10852, 16'd57018});
	test_expansion(128'h6beaf69b96fbfb337e420ee23f7937c1, {16'd38724, 16'd61697, 16'd39895, 16'd44029, 16'd40683, 16'd20710, 16'd61192, 16'd31789, 16'd59291, 16'd24794, 16'd13929, 16'd29054, 16'd50491, 16'd7150, 16'd27634, 16'd56561, 16'd16442, 16'd9331, 16'd29848, 16'd31050, 16'd52119, 16'd45051, 16'd43332, 16'd52512, 16'd42947, 16'd2264});
	test_expansion(128'h5867503a21f2370083db58f906caac20, {16'd1104, 16'd33826, 16'd41005, 16'd32845, 16'd30840, 16'd15895, 16'd23010, 16'd62472, 16'd5710, 16'd32948, 16'd16010, 16'd38340, 16'd32567, 16'd64572, 16'd7684, 16'd13423, 16'd64904, 16'd56681, 16'd26958, 16'd44992, 16'd20014, 16'd45245, 16'd27112, 16'd54341, 16'd44352, 16'd31107});
	test_expansion(128'h4dc01ea7c39e8492dfae3b053a71d303, {16'd1245, 16'd51327, 16'd7480, 16'd36719, 16'd51315, 16'd41251, 16'd50669, 16'd47984, 16'd56552, 16'd24588, 16'd57726, 16'd18816, 16'd21474, 16'd9003, 16'd61957, 16'd5760, 16'd46224, 16'd1781, 16'd18711, 16'd30952, 16'd63141, 16'd30813, 16'd62742, 16'd15611, 16'd61717, 16'd20807});
	test_expansion(128'h26c03f7a099040d060854c12e9dcb85f, {16'd1205, 16'd40651, 16'd32185, 16'd54861, 16'd11987, 16'd24797, 16'd33008, 16'd35750, 16'd56386, 16'd37996, 16'd27853, 16'd49651, 16'd22778, 16'd26857, 16'd17572, 16'd47758, 16'd20907, 16'd27866, 16'd46713, 16'd62312, 16'd35456, 16'd54841, 16'd10015, 16'd19440, 16'd47805, 16'd63844});
	test_expansion(128'h9ac9ffac9455a0892572ad1af372b5bb, {16'd5302, 16'd34052, 16'd59890, 16'd52307, 16'd45904, 16'd28093, 16'd14541, 16'd59498, 16'd60643, 16'd52977, 16'd39299, 16'd51897, 16'd26207, 16'd59954, 16'd60928, 16'd33222, 16'd10202, 16'd26852, 16'd60955, 16'd1065, 16'd50190, 16'd33191, 16'd16860, 16'd24673, 16'd35042, 16'd35328});
	test_expansion(128'hf804e329b0a54410ac594fcb613630ca, {16'd14704, 16'd28859, 16'd19236, 16'd19448, 16'd38168, 16'd51591, 16'd19971, 16'd10334, 16'd16286, 16'd1627, 16'd26150, 16'd28795, 16'd65337, 16'd64908, 16'd47583, 16'd50775, 16'd6747, 16'd23712, 16'd6142, 16'd44307, 16'd63440, 16'd452, 16'd5440, 16'd11822, 16'd49214, 16'd29005});
	test_expansion(128'haf536c43b278bc6428a9ac53566afcc1, {16'd44627, 16'd14669, 16'd4597, 16'd55432, 16'd61826, 16'd65251, 16'd38882, 16'd2414, 16'd44001, 16'd18513, 16'd48293, 16'd30612, 16'd51416, 16'd17713, 16'd19348, 16'd53818, 16'd624, 16'd24331, 16'd22420, 16'd62700, 16'd36683, 16'd33198, 16'd1547, 16'd56754, 16'd40428, 16'd8924});
	test_expansion(128'h721c7a8c0310cd749230ebb01e883a3b, {16'd53557, 16'd23754, 16'd46897, 16'd59301, 16'd56143, 16'd60951, 16'd8, 16'd60656, 16'd24670, 16'd47188, 16'd32839, 16'd1575, 16'd29295, 16'd24951, 16'd11318, 16'd53292, 16'd19600, 16'd26974, 16'd13448, 16'd55218, 16'd16482, 16'd54341, 16'd17160, 16'd51443, 16'd38814, 16'd22656});
	test_expansion(128'h1e6e4ea8dc0e9396ea47ebdebc7796b9, {16'd42023, 16'd9977, 16'd57923, 16'd6939, 16'd64988, 16'd32599, 16'd32435, 16'd42554, 16'd11496, 16'd56330, 16'd18191, 16'd57591, 16'd48184, 16'd8947, 16'd45006, 16'd39259, 16'd23664, 16'd58448, 16'd18868, 16'd14380, 16'd53768, 16'd18763, 16'd40278, 16'd27234, 16'd15689, 16'd26961});
	test_expansion(128'hd13a22d777c692ce26f3dc1ee4c17689, {16'd24739, 16'd19610, 16'd1208, 16'd33914, 16'd19474, 16'd1955, 16'd25001, 16'd45473, 16'd23402, 16'd40337, 16'd27248, 16'd13347, 16'd34620, 16'd27631, 16'd958, 16'd61397, 16'd46898, 16'd35313, 16'd57988, 16'd30311, 16'd3538, 16'd62889, 16'd6130, 16'd27747, 16'd61737, 16'd51317});
	test_expansion(128'hea7863a69dddefb13af864a3dfb150c7, {16'd9606, 16'd61165, 16'd23303, 16'd51004, 16'd2806, 16'd63532, 16'd29922, 16'd65007, 16'd11899, 16'd28546, 16'd22209, 16'd52123, 16'd9492, 16'd21723, 16'd15215, 16'd58319, 16'd13584, 16'd38605, 16'd17361, 16'd18679, 16'd1481, 16'd60369, 16'd26352, 16'd17217, 16'd35975, 16'd32644});
	test_expansion(128'h1925dc0d7f450594cbd528ce186c7135, {16'd17852, 16'd32765, 16'd18457, 16'd4876, 16'd10218, 16'd33744, 16'd15826, 16'd29063, 16'd65112, 16'd15308, 16'd49419, 16'd7355, 16'd26315, 16'd21921, 16'd17590, 16'd1282, 16'd56693, 16'd9293, 16'd13207, 16'd5441, 16'd2414, 16'd22882, 16'd40257, 16'd14206, 16'd38685, 16'd62044});
	test_expansion(128'h3b8953366de2774aa1945c318a5a99e5, {16'd27837, 16'd40333, 16'd54323, 16'd22058, 16'd60500, 16'd45021, 16'd64751, 16'd16270, 16'd24075, 16'd27733, 16'd29075, 16'd41356, 16'd22530, 16'd40168, 16'd42532, 16'd12888, 16'd50635, 16'd44622, 16'd52171, 16'd27096, 16'd5187, 16'd61573, 16'd13293, 16'd63126, 16'd61724, 16'd38233});
	test_expansion(128'hddc924a2eaa70a8e5a46a65a4aed5e7a, {16'd58693, 16'd2890, 16'd43108, 16'd43450, 16'd10354, 16'd7406, 16'd58703, 16'd5606, 16'd62225, 16'd51271, 16'd46240, 16'd14443, 16'd55509, 16'd21639, 16'd14204, 16'd54971, 16'd14448, 16'd63370, 16'd29020, 16'd16240, 16'd5870, 16'd46185, 16'd42660, 16'd20702, 16'd12111, 16'd31014});
	test_expansion(128'he6d96dba3efc0fdf52e343b0fc51bdfd, {16'd31480, 16'd32651, 16'd41819, 16'd57791, 16'd33991, 16'd64651, 16'd24083, 16'd3979, 16'd34566, 16'd29111, 16'd49074, 16'd38487, 16'd45146, 16'd28937, 16'd6373, 16'd31198, 16'd19020, 16'd33675, 16'd8487, 16'd8877, 16'd63590, 16'd22232, 16'd21440, 16'd16341, 16'd21805, 16'd59835});
	test_expansion(128'h5d4ed43625a9db18c001d6e3606ab4db, {16'd36406, 16'd15030, 16'd50367, 16'd35331, 16'd19700, 16'd31454, 16'd15118, 16'd47647, 16'd16605, 16'd27086, 16'd51755, 16'd10925, 16'd13131, 16'd57511, 16'd46135, 16'd52233, 16'd45284, 16'd62793, 16'd17838, 16'd4469, 16'd53062, 16'd6290, 16'd14910, 16'd49856, 16'd10151, 16'd8812});
	test_expansion(128'h2c590d6bcc203fab7d2f36b2aa9ce486, {16'd38099, 16'd65331, 16'd58560, 16'd60779, 16'd15322, 16'd13979, 16'd29612, 16'd64838, 16'd35401, 16'd63924, 16'd52833, 16'd29056, 16'd60375, 16'd12526, 16'd7490, 16'd2523, 16'd7354, 16'd64357, 16'd11453, 16'd20802, 16'd33972, 16'd6249, 16'd48032, 16'd64676, 16'd53563, 16'd42225});
	test_expansion(128'ha0d4ba9d15d1ab8d7d1ed4e58dc34be5, {16'd59875, 16'd12222, 16'd11381, 16'd11712, 16'd23047, 16'd42274, 16'd27998, 16'd27405, 16'd31339, 16'd59165, 16'd52337, 16'd52386, 16'd52833, 16'd26305, 16'd56182, 16'd5986, 16'd43376, 16'd43220, 16'd13694, 16'd60948, 16'd36160, 16'd14325, 16'd42081, 16'd48207, 16'd34645, 16'd1859});
	test_expansion(128'hd708df76efe35a2fec2759e9648adde3, {16'd59965, 16'd23321, 16'd55316, 16'd22849, 16'd7261, 16'd45630, 16'd57374, 16'd4225, 16'd38973, 16'd39929, 16'd49854, 16'd27435, 16'd34897, 16'd61770, 16'd42795, 16'd701, 16'd27089, 16'd33465, 16'd59665, 16'd23980, 16'd63820, 16'd15734, 16'd58308, 16'd170, 16'd49506, 16'd2233});
	test_expansion(128'h7326c18c6542b262388365ff41abe221, {16'd34016, 16'd2856, 16'd14398, 16'd14229, 16'd33734, 16'd21956, 16'd61625, 16'd34378, 16'd26446, 16'd54841, 16'd31975, 16'd17616, 16'd59896, 16'd9644, 16'd26528, 16'd40567, 16'd63306, 16'd61616, 16'd61560, 16'd59660, 16'd37793, 16'd3154, 16'd62557, 16'd27195, 16'd2615, 16'd19224});
	test_expansion(128'h42e64040bd9777663aa595606b6c4fae, {16'd23242, 16'd41930, 16'd41728, 16'd27307, 16'd47583, 16'd48941, 16'd63744, 16'd41731, 16'd30704, 16'd8651, 16'd54232, 16'd56896, 16'd19982, 16'd3660, 16'd8951, 16'd50951, 16'd14380, 16'd24055, 16'd47743, 16'd46326, 16'd64625, 16'd26449, 16'd26007, 16'd27695, 16'd48281, 16'd9356});
	test_expansion(128'h49d560e0b5bcb3e8fc665c752d4709d0, {16'd14918, 16'd12864, 16'd16298, 16'd58925, 16'd8404, 16'd53283, 16'd10686, 16'd9223, 16'd6017, 16'd52155, 16'd8097, 16'd58388, 16'd35018, 16'd10713, 16'd50143, 16'd40219, 16'd2436, 16'd43487, 16'd413, 16'd56480, 16'd52061, 16'd5423, 16'd59517, 16'd43552, 16'd25979, 16'd9346});
	test_expansion(128'h94209f95af8c78ae800abdb0bffbac66, {16'd8557, 16'd57869, 16'd9977, 16'd53106, 16'd8916, 16'd22079, 16'd56996, 16'd13437, 16'd63382, 16'd26408, 16'd23701, 16'd57368, 16'd24823, 16'd39181, 16'd45095, 16'd11000, 16'd45468, 16'd53521, 16'd50935, 16'd44989, 16'd52561, 16'd30438, 16'd54985, 16'd21432, 16'd49834, 16'd61201});
	test_expansion(128'hb5d23670d8129cdaca247e38581582dd, {16'd4254, 16'd40834, 16'd48594, 16'd43841, 16'd63991, 16'd6456, 16'd4497, 16'd33469, 16'd14210, 16'd55444, 16'd61328, 16'd46666, 16'd55822, 16'd19381, 16'd54909, 16'd12658, 16'd4123, 16'd3487, 16'd43719, 16'd53667, 16'd46230, 16'd21235, 16'd19853, 16'd36807, 16'd45635, 16'd24403});
	test_expansion(128'hffcfb3bb746dc9a40aaa36d897bb5572, {16'd6891, 16'd1878, 16'd60229, 16'd47241, 16'd16463, 16'd42406, 16'd31504, 16'd52567, 16'd45033, 16'd51229, 16'd5076, 16'd32022, 16'd13779, 16'd34034, 16'd11072, 16'd3960, 16'd58351, 16'd57075, 16'd1067, 16'd42090, 16'd36653, 16'd34778, 16'd61905, 16'd28540, 16'd44076, 16'd59277});
	test_expansion(128'h9398ade2ce63630a094a4c210294aa02, {16'd9221, 16'd16133, 16'd8976, 16'd2875, 16'd37526, 16'd50352, 16'd60097, 16'd47984, 16'd19532, 16'd30651, 16'd47228, 16'd26434, 16'd16294, 16'd60073, 16'd54173, 16'd12109, 16'd4849, 16'd19352, 16'd31040, 16'd42339, 16'd22084, 16'd60294, 16'd928, 16'd30973, 16'd27041, 16'd59920});
	test_expansion(128'h04d48e34060e6dfc8ad91ab57d9a5805, {16'd42064, 16'd41011, 16'd4784, 16'd36032, 16'd58218, 16'd6052, 16'd22550, 16'd33991, 16'd16782, 16'd22842, 16'd40019, 16'd60217, 16'd57112, 16'd6384, 16'd49318, 16'd42802, 16'd33690, 16'd60230, 16'd49447, 16'd58006, 16'd12934, 16'd53421, 16'd13054, 16'd7568, 16'd51058, 16'd41155});
	test_expansion(128'h504f23e10496ec64a83dc7e917231417, {16'd7237, 16'd62338, 16'd35510, 16'd45115, 16'd28009, 16'd39725, 16'd6480, 16'd18165, 16'd55123, 16'd23485, 16'd13623, 16'd30370, 16'd7685, 16'd65073, 16'd46904, 16'd59040, 16'd31557, 16'd24600, 16'd44118, 16'd25004, 16'd57696, 16'd8065, 16'd5204, 16'd52859, 16'd59211, 16'd52492});
	test_expansion(128'h2b965b96702faea42ef86f20179612ed, {16'd46123, 16'd2668, 16'd9918, 16'd14723, 16'd19608, 16'd30150, 16'd34704, 16'd40459, 16'd60559, 16'd48644, 16'd17712, 16'd60826, 16'd31309, 16'd13322, 16'd56336, 16'd16184, 16'd56856, 16'd32973, 16'd8886, 16'd37532, 16'd53320, 16'd20074, 16'd57672, 16'd33900, 16'd65142, 16'd7128});
	test_expansion(128'hfd39904956fb12e353eb866c40f9ef7d, {16'd32845, 16'd45358, 16'd40365, 16'd41839, 16'd34368, 16'd42371, 16'd38458, 16'd39267, 16'd38452, 16'd13410, 16'd28337, 16'd18267, 16'd49354, 16'd38315, 16'd27128, 16'd14660, 16'd7062, 16'd33893, 16'd55572, 16'd64475, 16'd38903, 16'd9580, 16'd12163, 16'd64118, 16'd18170, 16'd49743});
	test_expansion(128'hc1aec729eebd0e1baf5900ce3daad665, {16'd62690, 16'd63698, 16'd19681, 16'd40386, 16'd6206, 16'd21591, 16'd30769, 16'd11820, 16'd64385, 16'd63944, 16'd35095, 16'd49840, 16'd17415, 16'd59761, 16'd4597, 16'd30070, 16'd38642, 16'd12193, 16'd35461, 16'd14203, 16'd142, 16'd20371, 16'd15333, 16'd37413, 16'd55908, 16'd55672});
	test_expansion(128'hcafd38cde12165b6767b3435c038d36d, {16'd18259, 16'd24863, 16'd54302, 16'd62678, 16'd55352, 16'd36479, 16'd44317, 16'd45108, 16'd41887, 16'd12253, 16'd52310, 16'd35820, 16'd63921, 16'd10805, 16'd16133, 16'd32643, 16'd20559, 16'd26475, 16'd52506, 16'd12375, 16'd36188, 16'd49492, 16'd5990, 16'd40690, 16'd12599, 16'd14573});
	test_expansion(128'hfcfa6a9d8375af567394ed6933eafc25, {16'd40535, 16'd48909, 16'd59727, 16'd16940, 16'd2960, 16'd58966, 16'd52440, 16'd62607, 16'd26562, 16'd37882, 16'd60914, 16'd58571, 16'd62991, 16'd23231, 16'd59003, 16'd5859, 16'd27127, 16'd12508, 16'd14407, 16'd3849, 16'd6485, 16'd25127, 16'd1212, 16'd10923, 16'd27727, 16'd25868});
	test_expansion(128'heba7bbaaadfa8d3b6da3df60a4457ae2, {16'd25836, 16'd18045, 16'd8764, 16'd8956, 16'd61262, 16'd3822, 16'd22467, 16'd35287, 16'd10252, 16'd29326, 16'd6767, 16'd25781, 16'd41609, 16'd41892, 16'd54733, 16'd2274, 16'd54276, 16'd14719, 16'd27014, 16'd35799, 16'd34406, 16'd40169, 16'd28627, 16'd3522, 16'd62111, 16'd35658});
	test_expansion(128'h28831fae7b669b2e861128af774cb7f5, {16'd50591, 16'd32034, 16'd42246, 16'd65263, 16'd46015, 16'd27937, 16'd7146, 16'd59540, 16'd9695, 16'd14283, 16'd3336, 16'd65411, 16'd36942, 16'd23319, 16'd48526, 16'd15822, 16'd40575, 16'd53620, 16'd11319, 16'd59436, 16'd41186, 16'd45102, 16'd31230, 16'd38740, 16'd11942, 16'd5268});
	test_expansion(128'h5d038188564a520e4404ae7b3b7262c9, {16'd65157, 16'd16526, 16'd6864, 16'd49517, 16'd63142, 16'd31672, 16'd364, 16'd43726, 16'd32225, 16'd35664, 16'd55611, 16'd5183, 16'd42439, 16'd28141, 16'd16406, 16'd11405, 16'd21908, 16'd8929, 16'd54269, 16'd51164, 16'd8217, 16'd53675, 16'd23047, 16'd41089, 16'd55642, 16'd55005});
	test_expansion(128'h49b31968e4f1b987320bf5a4e86de762, {16'd42798, 16'd37822, 16'd62894, 16'd63211, 16'd30207, 16'd37, 16'd30681, 16'd6120, 16'd40492, 16'd10906, 16'd1616, 16'd6606, 16'd38733, 16'd16811, 16'd50630, 16'd15209, 16'd44826, 16'd21222, 16'd62949, 16'd51340, 16'd58054, 16'd32368, 16'd27412, 16'd47360, 16'd44087, 16'd49400});
	test_expansion(128'h578acc56d427044b26e97470a586d27e, {16'd45374, 16'd33520, 16'd47031, 16'd51110, 16'd38196, 16'd49586, 16'd37085, 16'd21133, 16'd6447, 16'd18812, 16'd40858, 16'd9297, 16'd50207, 16'd62134, 16'd548, 16'd7607, 16'd36615, 16'd19755, 16'd10358, 16'd56935, 16'd26615, 16'd51479, 16'd28697, 16'd36195, 16'd58987, 16'd40523});
	test_expansion(128'hfcc75c699648b553d6a7e35fec885b41, {16'd25899, 16'd12064, 16'd20967, 16'd58712, 16'd61640, 16'd43174, 16'd23192, 16'd16264, 16'd26677, 16'd2749, 16'd40097, 16'd25360, 16'd8108, 16'd21871, 16'd16218, 16'd56545, 16'd48064, 16'd43281, 16'd21507, 16'd63407, 16'd41994, 16'd51254, 16'd22257, 16'd55427, 16'd19921, 16'd2238});
	test_expansion(128'h40bb74684bdc3c14f2df1aa1a3324e50, {16'd27831, 16'd31086, 16'd26995, 16'd22715, 16'd8936, 16'd26581, 16'd7845, 16'd3633, 16'd43098, 16'd46242, 16'd41358, 16'd10040, 16'd28223, 16'd56722, 16'd36556, 16'd44994, 16'd13104, 16'd46410, 16'd62045, 16'd39455, 16'd25729, 16'd16456, 16'd39917, 16'd29956, 16'd38317, 16'd2958});
	test_expansion(128'h565f4e30c29372bf1d102abd1325c7f5, {16'd17356, 16'd38305, 16'd33496, 16'd23192, 16'd63896, 16'd47760, 16'd55589, 16'd50151, 16'd41600, 16'd20787, 16'd27796, 16'd58184, 16'd50966, 16'd57012, 16'd38816, 16'd10434, 16'd20387, 16'd37314, 16'd26804, 16'd6898, 16'd63137, 16'd3358, 16'd24318, 16'd7741, 16'd166, 16'd42413});
	test_expansion(128'h27443e5b58ed8fe1f8697ae9fe38aedd, {16'd35775, 16'd30510, 16'd20452, 16'd15382, 16'd44559, 16'd39769, 16'd37254, 16'd54761, 16'd10666, 16'd18278, 16'd35893, 16'd28915, 16'd17379, 16'd448, 16'd21460, 16'd8848, 16'd20755, 16'd28923, 16'd43608, 16'd50327, 16'd64382, 16'd35927, 16'd21715, 16'd19850, 16'd26818, 16'd17593});
	test_expansion(128'h703da1952f5c1c7aa1f6f40c936ec2f2, {16'd20258, 16'd40651, 16'd51248, 16'd29424, 16'd11462, 16'd38899, 16'd59918, 16'd36154, 16'd23950, 16'd34167, 16'd43358, 16'd30711, 16'd29913, 16'd60650, 16'd31417, 16'd38921, 16'd34727, 16'd56763, 16'd45265, 16'd19995, 16'd56406, 16'd33327, 16'd16716, 16'd46700, 16'd23826, 16'd24385});
	test_expansion(128'h79c1cc80a0fd4a6ffc9e5440b4d90b24, {16'd51596, 16'd29746, 16'd4926, 16'd63064, 16'd29800, 16'd30901, 16'd41202, 16'd29049, 16'd35541, 16'd27792, 16'd12271, 16'd39939, 16'd58287, 16'd50826, 16'd15391, 16'd55882, 16'd29475, 16'd48581, 16'd43167, 16'd7886, 16'd32637, 16'd21143, 16'd50638, 16'd55748, 16'd20641, 16'd17082});
	test_expansion(128'h680ffb2b06605bac8d1e5f6a8591413b, {16'd29698, 16'd57025, 16'd65120, 16'd46882, 16'd14648, 16'd61430, 16'd31223, 16'd20114, 16'd43798, 16'd20707, 16'd51441, 16'd31000, 16'd30779, 16'd13847, 16'd48274, 16'd6288, 16'd23603, 16'd64202, 16'd34456, 16'd5548, 16'd10963, 16'd35970, 16'd48193, 16'd31006, 16'd33760, 16'd17780});
	test_expansion(128'h068c9a3d71dd7db900e6a35c2261b79e, {16'd17086, 16'd42534, 16'd58963, 16'd52782, 16'd63209, 16'd36224, 16'd18797, 16'd35920, 16'd39111, 16'd42759, 16'd4650, 16'd64585, 16'd17584, 16'd15744, 16'd13436, 16'd24957, 16'd13484, 16'd29196, 16'd44105, 16'd39217, 16'd65499, 16'd4932, 16'd9000, 16'd25140, 16'd44373, 16'd13389});
	test_expansion(128'h698d205d7251f974368eba065bd71386, {16'd16331, 16'd25546, 16'd61728, 16'd51506, 16'd43365, 16'd14627, 16'd51615, 16'd49585, 16'd19034, 16'd16617, 16'd44156, 16'd21510, 16'd13083, 16'd56113, 16'd14492, 16'd51216, 16'd43015, 16'd3473, 16'd22335, 16'd31515, 16'd41093, 16'd21080, 16'd46567, 16'd17551, 16'd49341, 16'd18146});
	test_expansion(128'ha9bdbc713b8d6620dec2210889c856e5, {16'd28869, 16'd50006, 16'd46784, 16'd32542, 16'd260, 16'd33396, 16'd41575, 16'd35032, 16'd34192, 16'd24502, 16'd6630, 16'd15980, 16'd1033, 16'd4843, 16'd21325, 16'd63756, 16'd53356, 16'd10721, 16'd44496, 16'd64961, 16'd404, 16'd64302, 16'd39342, 16'd55516, 16'd28031, 16'd62506});
	test_expansion(128'h9d99e13cb33244ccbc61d777091b37b9, {16'd21724, 16'd51353, 16'd47761, 16'd54597, 16'd57267, 16'd62119, 16'd32562, 16'd9127, 16'd51514, 16'd25707, 16'd63909, 16'd40930, 16'd49578, 16'd4451, 16'd48653, 16'd9569, 16'd5632, 16'd36089, 16'd30984, 16'd34733, 16'd5752, 16'd4755, 16'd36436, 16'd9689, 16'd54592, 16'd32294});
	test_expansion(128'hcd763bdaccbd52ee5ec2554321fbca00, {16'd51696, 16'd35909, 16'd3395, 16'd21162, 16'd30479, 16'd784, 16'd19460, 16'd48254, 16'd9124, 16'd7880, 16'd14889, 16'd22701, 16'd28960, 16'd43271, 16'd24589, 16'd9455, 16'd22585, 16'd19058, 16'd29403, 16'd60746, 16'd31155, 16'd52410, 16'd38283, 16'd61864, 16'd5608, 16'd65300});
	test_expansion(128'h11c7f50b1fa3a82fbf69fb21735ca85b, {16'd56561, 16'd510, 16'd2577, 16'd15179, 16'd35357, 16'd43668, 16'd18778, 16'd33289, 16'd22769, 16'd46408, 16'd23218, 16'd8884, 16'd1870, 16'd6107, 16'd12630, 16'd29399, 16'd59881, 16'd5848, 16'd38291, 16'd50314, 16'd34689, 16'd56075, 16'd33293, 16'd54569, 16'd44542, 16'd45729});
	test_expansion(128'hdb53965391903257c4e51e36f5a78c13, {16'd21657, 16'd25531, 16'd56192, 16'd14828, 16'd37847, 16'd61735, 16'd55175, 16'd326, 16'd28785, 16'd31707, 16'd7438, 16'd56294, 16'd5656, 16'd9665, 16'd15092, 16'd2976, 16'd13963, 16'd35544, 16'd56763, 16'd10688, 16'd42733, 16'd60314, 16'd11407, 16'd28499, 16'd40312, 16'd17750});
	test_expansion(128'h85b761f74c8b5dd1163fb3b504351f08, {16'd11896, 16'd354, 16'd52685, 16'd16821, 16'd2325, 16'd49881, 16'd54449, 16'd43057, 16'd55953, 16'd31842, 16'd44203, 16'd59155, 16'd9849, 16'd20831, 16'd26538, 16'd31687, 16'd4121, 16'd24005, 16'd58748, 16'd4893, 16'd7441, 16'd44949, 16'd63914, 16'd2860, 16'd54288, 16'd28188});
	test_expansion(128'he09c7b18f43a56757a9d3f9dfe6a03a6, {16'd31618, 16'd384, 16'd34401, 16'd63273, 16'd35873, 16'd41170, 16'd38502, 16'd41342, 16'd51970, 16'd36695, 16'd4208, 16'd10663, 16'd7256, 16'd15823, 16'd20180, 16'd56000, 16'd56199, 16'd50541, 16'd40704, 16'd20693, 16'd15670, 16'd56215, 16'd42494, 16'd16778, 16'd44317, 16'd48678});
	test_expansion(128'hd24702bc9b64e808f8acce00865588a5, {16'd4715, 16'd48732, 16'd57201, 16'd11772, 16'd31, 16'd32156, 16'd12560, 16'd58101, 16'd17500, 16'd4412, 16'd37254, 16'd56393, 16'd9456, 16'd2471, 16'd28544, 16'd22313, 16'd42926, 16'd49137, 16'd406, 16'd55250, 16'd57637, 16'd59941, 16'd60998, 16'd15227, 16'd50922, 16'd3792});
	test_expansion(128'h0ea40874c6db4fe745e1bc08e3f3c7a0, {16'd45710, 16'd15442, 16'd14332, 16'd64030, 16'd52618, 16'd44764, 16'd6437, 16'd4950, 16'd53245, 16'd1234, 16'd11108, 16'd51480, 16'd10039, 16'd49900, 16'd57647, 16'd43773, 16'd54576, 16'd33105, 16'd2707, 16'd24217, 16'd24019, 16'd43667, 16'd48023, 16'd54264, 16'd7869, 16'd5911});
	test_expansion(128'hfe15b32bd1207d887c7d9558e67841aa, {16'd59643, 16'd9316, 16'd4207, 16'd59514, 16'd35785, 16'd46601, 16'd58497, 16'd33813, 16'd22989, 16'd55356, 16'd6935, 16'd31266, 16'd31010, 16'd28135, 16'd55386, 16'd38587, 16'd5909, 16'd34671, 16'd14411, 16'd32637, 16'd2131, 16'd43393, 16'd62699, 16'd28694, 16'd34214, 16'd50051});
	test_expansion(128'hf1520f488658c9e596dbff58eda9d8c6, {16'd57395, 16'd1538, 16'd20426, 16'd43329, 16'd4220, 16'd1464, 16'd11989, 16'd40621, 16'd24723, 16'd37195, 16'd24111, 16'd6440, 16'd59925, 16'd59922, 16'd50412, 16'd41001, 16'd24181, 16'd12038, 16'd29835, 16'd46495, 16'd51904, 16'd41665, 16'd36928, 16'd34787, 16'd57654, 16'd51747});
	test_expansion(128'h9904084060374760ddf8c0d92a0140b9, {16'd21103, 16'd56104, 16'd51645, 16'd25023, 16'd51749, 16'd27232, 16'd19340, 16'd29408, 16'd3949, 16'd23396, 16'd2852, 16'd22116, 16'd15407, 16'd20197, 16'd17253, 16'd37312, 16'd53062, 16'd52378, 16'd32955, 16'd50503, 16'd35224, 16'd52612, 16'd59262, 16'd37619, 16'd45864, 16'd15207});
	test_expansion(128'hbd4f8adc6835fd2ddc81717a7cfdc481, {16'd17966, 16'd50679, 16'd59419, 16'd26570, 16'd47225, 16'd40846, 16'd38202, 16'd17833, 16'd38034, 16'd55480, 16'd52615, 16'd3794, 16'd633, 16'd25728, 16'd11065, 16'd55370, 16'd62372, 16'd57641, 16'd4974, 16'd47019, 16'd933, 16'd14330, 16'd38551, 16'd26345, 16'd36042, 16'd41040});
	test_expansion(128'he3eaabb2202d3eac54515a51f1aed732, {16'd58235, 16'd46735, 16'd1269, 16'd64559, 16'd25009, 16'd4430, 16'd21534, 16'd63090, 16'd24831, 16'd20095, 16'd11602, 16'd56872, 16'd41308, 16'd11107, 16'd55487, 16'd40982, 16'd23596, 16'd30308, 16'd50420, 16'd57140, 16'd21163, 16'd17395, 16'd21676, 16'd38603, 16'd18330, 16'd50499});
	test_expansion(128'h6d3fad6ddd3b88b4bb5c633c8f6ef548, {16'd13311, 16'd43558, 16'd27029, 16'd25865, 16'd55045, 16'd26439, 16'd59023, 16'd24262, 16'd33873, 16'd23636, 16'd59411, 16'd40086, 16'd8879, 16'd21448, 16'd32822, 16'd54199, 16'd56162, 16'd48366, 16'd45378, 16'd20816, 16'd53038, 16'd14883, 16'd1321, 16'd36495, 16'd30899, 16'd16965});
	test_expansion(128'h2e0c3dc269dcaf8832b72ab9199bcc31, {16'd4424, 16'd18156, 16'd5074, 16'd22571, 16'd5852, 16'd38683, 16'd47654, 16'd30847, 16'd60631, 16'd54877, 16'd61158, 16'd12192, 16'd32506, 16'd63590, 16'd64648, 16'd23347, 16'd26991, 16'd1403, 16'd48249, 16'd61020, 16'd42465, 16'd64051, 16'd39892, 16'd23404, 16'd41324, 16'd55530});
	test_expansion(128'h4a9f2d0387e92c693b76230a5e50318b, {16'd3684, 16'd50936, 16'd10198, 16'd43747, 16'd19444, 16'd40724, 16'd33450, 16'd45244, 16'd14598, 16'd36835, 16'd62589, 16'd37950, 16'd18682, 16'd10876, 16'd19537, 16'd31716, 16'd60985, 16'd12642, 16'd15262, 16'd28812, 16'd6934, 16'd56260, 16'd32271, 16'd44284, 16'd44436, 16'd21760});
	test_expansion(128'h413cb996112295d0e3255568f1b2965b, {16'd7163, 16'd43647, 16'd50836, 16'd10238, 16'd8121, 16'd8984, 16'd58124, 16'd49351, 16'd41967, 16'd33814, 16'd48025, 16'd55481, 16'd61249, 16'd47694, 16'd56122, 16'd11376, 16'd20262, 16'd54102, 16'd34609, 16'd45302, 16'd21538, 16'd26841, 16'd9321, 16'd52805, 16'd48837, 16'd23308});
	test_expansion(128'h0218544e329930119baf178306764937, {16'd18315, 16'd29253, 16'd128, 16'd5160, 16'd59938, 16'd60187, 16'd29736, 16'd1094, 16'd28377, 16'd5237, 16'd6213, 16'd54593, 16'd39143, 16'd49397, 16'd52687, 16'd10204, 16'd26536, 16'd11763, 16'd34080, 16'd18837, 16'd48290, 16'd42564, 16'd54299, 16'd55882, 16'd47601, 16'd28537});
	test_expansion(128'h8d725fdda2970d8e55b788d29de5724e, {16'd22902, 16'd43348, 16'd10762, 16'd63290, 16'd25814, 16'd64510, 16'd61408, 16'd22090, 16'd8487, 16'd21655, 16'd14923, 16'd22436, 16'd18832, 16'd7256, 16'd57901, 16'd62654, 16'd3502, 16'd18435, 16'd28073, 16'd16077, 16'd23585, 16'd14048, 16'd46644, 16'd6294, 16'd3693, 16'd27735});
	test_expansion(128'ha39a0ba6d15028cd386f9314f8000b59, {16'd52052, 16'd48024, 16'd31591, 16'd37618, 16'd35063, 16'd52499, 16'd33747, 16'd36649, 16'd49726, 16'd51050, 16'd63520, 16'd38952, 16'd55729, 16'd37767, 16'd38339, 16'd57457, 16'd24404, 16'd2958, 16'd58932, 16'd24232, 16'd16637, 16'd63351, 16'd3333, 16'd1406, 16'd42021, 16'd5325});
	test_expansion(128'h80b1344fcb0500eabe717b3dacc543e8, {16'd47582, 16'd36356, 16'd7365, 16'd35640, 16'd31884, 16'd15929, 16'd40810, 16'd59811, 16'd57253, 16'd36463, 16'd30646, 16'd13222, 16'd65093, 16'd32914, 16'd4531, 16'd15667, 16'd64852, 16'd24936, 16'd43988, 16'd40044, 16'd11338, 16'd49028, 16'd59415, 16'd39632, 16'd11637, 16'd9687});
	test_expansion(128'h3b1b378ad9fbdde54fcdf28b8a147383, {16'd7121, 16'd17470, 16'd60616, 16'd64103, 16'd4734, 16'd14589, 16'd50107, 16'd9276, 16'd54530, 16'd11162, 16'd7986, 16'd22508, 16'd10728, 16'd44011, 16'd61801, 16'd58869, 16'd32115, 16'd30024, 16'd39481, 16'd35348, 16'd21298, 16'd41253, 16'd52182, 16'd18690, 16'd3608, 16'd57777});
	test_expansion(128'hc1565cad0a6b83316f96390ccf8c0f91, {16'd62116, 16'd52887, 16'd5060, 16'd13951, 16'd6328, 16'd25657, 16'd13510, 16'd10125, 16'd12060, 16'd43099, 16'd42960, 16'd12643, 16'd702, 16'd24214, 16'd3927, 16'd18724, 16'd29490, 16'd27866, 16'd34507, 16'd33557, 16'd23476, 16'd13333, 16'd36249, 16'd4718, 16'd39926, 16'd32610});
	test_expansion(128'h70a7fad947fc9346b87e08fcd8ab103a, {16'd60120, 16'd27774, 16'd64914, 16'd36120, 16'd35911, 16'd10895, 16'd3487, 16'd55807, 16'd10566, 16'd9564, 16'd45676, 16'd31272, 16'd26232, 16'd46357, 16'd59395, 16'd52332, 16'd17983, 16'd51911, 16'd14460, 16'd64155, 16'd29585, 16'd26913, 16'd11700, 16'd44291, 16'd61131, 16'd25285});
	test_expansion(128'h8eaaad0ac82116cf44e1fc2b51e51e82, {16'd21755, 16'd36713, 16'd34741, 16'd64114, 16'd2934, 16'd45714, 16'd17354, 16'd52245, 16'd20888, 16'd33863, 16'd41431, 16'd41445, 16'd3406, 16'd61971, 16'd60593, 16'd44941, 16'd10750, 16'd63027, 16'd51718, 16'd51998, 16'd13322, 16'd27621, 16'd56063, 16'd41021, 16'd834, 16'd54575});
	test_expansion(128'h25d247b5ab575384e2f08bc0bf2df75a, {16'd3470, 16'd8359, 16'd56259, 16'd44704, 16'd58996, 16'd63201, 16'd8209, 16'd48264, 16'd10186, 16'd39245, 16'd60135, 16'd55408, 16'd58728, 16'd17493, 16'd27523, 16'd4725, 16'd5908, 16'd63249, 16'd22567, 16'd41913, 16'd32628, 16'd46955, 16'd8261, 16'd30671, 16'd31746, 16'd57807});
	test_expansion(128'hd7d7c57aca093d49b38c7723cdf1b896, {16'd39636, 16'd32990, 16'd46238, 16'd58741, 16'd47281, 16'd52457, 16'd64203, 16'd44970, 16'd53050, 16'd49956, 16'd64181, 16'd31516, 16'd22857, 16'd29815, 16'd11229, 16'd11894, 16'd63989, 16'd22804, 16'd64450, 16'd3353, 16'd16548, 16'd41149, 16'd48118, 16'd26975, 16'd48070, 16'd1671});
	test_expansion(128'h1d4faed896302442395e65bfbfa85b40, {16'd56234, 16'd19486, 16'd41421, 16'd32228, 16'd41823, 16'd31098, 16'd42801, 16'd3887, 16'd51599, 16'd8429, 16'd45570, 16'd26599, 16'd34871, 16'd31101, 16'd61785, 16'd1700, 16'd41038, 16'd37552, 16'd40504, 16'd44301, 16'd59509, 16'd8396, 16'd13715, 16'd46837, 16'd39372, 16'd11855});
	test_expansion(128'h18e18637f09ab7d36da5973cc6c699a7, {16'd49591, 16'd44797, 16'd58188, 16'd58343, 16'd52673, 16'd45109, 16'd8891, 16'd62197, 16'd17404, 16'd22895, 16'd49540, 16'd33358, 16'd14343, 16'd59519, 16'd14598, 16'd16679, 16'd48127, 16'd17690, 16'd6096, 16'd22532, 16'd24664, 16'd9785, 16'd9066, 16'd47217, 16'd44938, 16'd63284});
	test_expansion(128'hb81deac8f0a9cebb0c40a23cc03e4e56, {16'd13643, 16'd10147, 16'd18779, 16'd38213, 16'd48107, 16'd45436, 16'd29031, 16'd29807, 16'd22512, 16'd23807, 16'd50326, 16'd35791, 16'd11815, 16'd30550, 16'd33357, 16'd14890, 16'd41980, 16'd15898, 16'd37470, 16'd30528, 16'd17974, 16'd61534, 16'd8471, 16'd57203, 16'd24104, 16'd33758});
	test_expansion(128'he4c8cee5a00956499b9149dfbcd5ee07, {16'd51094, 16'd23252, 16'd42156, 16'd23880, 16'd61859, 16'd31723, 16'd29693, 16'd3102, 16'd3589, 16'd34867, 16'd33818, 16'd27100, 16'd39468, 16'd16931, 16'd2591, 16'd37010, 16'd18887, 16'd29881, 16'd10376, 16'd10033, 16'd16545, 16'd5485, 16'd63999, 16'd44921, 16'd55683, 16'd51102});
	test_expansion(128'hf6b99dd0a59952eae6c14bd5b57c1741, {16'd57700, 16'd57033, 16'd28792, 16'd54379, 16'd38125, 16'd58977, 16'd56510, 16'd6390, 16'd16760, 16'd4380, 16'd59324, 16'd43432, 16'd1591, 16'd12894, 16'd27592, 16'd26210, 16'd39653, 16'd8854, 16'd58538, 16'd21870, 16'd30271, 16'd45861, 16'd34079, 16'd18966, 16'd38038, 16'd52436});
	test_expansion(128'ha1f604becca6beb7a2ada682c68f5bbc, {16'd27868, 16'd11606, 16'd6633, 16'd37903, 16'd10489, 16'd14954, 16'd15554, 16'd28060, 16'd35630, 16'd33230, 16'd26631, 16'd9422, 16'd24099, 16'd11797, 16'd29481, 16'd37884, 16'd13287, 16'd12184, 16'd21911, 16'd40609, 16'd42026, 16'd35791, 16'd37593, 16'd37443, 16'd24810, 16'd53006});
	test_expansion(128'h0ba5fde6b296fb5adf9829f9905346fb, {16'd39771, 16'd3963, 16'd36313, 16'd35107, 16'd13641, 16'd38612, 16'd52521, 16'd17503, 16'd46547, 16'd46573, 16'd33751, 16'd27339, 16'd44836, 16'd52611, 16'd15182, 16'd18434, 16'd45427, 16'd22491, 16'd62360, 16'd48615, 16'd10729, 16'd11690, 16'd62721, 16'd666, 16'd25056, 16'd11063});
	test_expansion(128'h8c5cfbab8295d0356d6c6f636500ff98, {16'd21896, 16'd11835, 16'd4583, 16'd28478, 16'd55874, 16'd52656, 16'd65195, 16'd59557, 16'd12793, 16'd64924, 16'd31204, 16'd44654, 16'd25491, 16'd35847, 16'd45274, 16'd35845, 16'd62059, 16'd13451, 16'd38776, 16'd10325, 16'd42783, 16'd58725, 16'd46033, 16'd567, 16'd320, 16'd31126});
	test_expansion(128'had7e52913889bba91ade17ea16af757a, {16'd20151, 16'd62311, 16'd13716, 16'd21012, 16'd49928, 16'd60468, 16'd27392, 16'd15432, 16'd31348, 16'd38332, 16'd47265, 16'd52088, 16'd35610, 16'd45653, 16'd9372, 16'd1107, 16'd12035, 16'd3155, 16'd6408, 16'd52287, 16'd30458, 16'd21307, 16'd20780, 16'd5235, 16'd63952, 16'd63499});
	test_expansion(128'hfdd7b1342a4d1203bd359af3016e2f4c, {16'd9377, 16'd37596, 16'd50154, 16'd37380, 16'd59989, 16'd21391, 16'd61142, 16'd56313, 16'd64349, 16'd33594, 16'd19905, 16'd49846, 16'd39570, 16'd56103, 16'd39303, 16'd49421, 16'd40013, 16'd46710, 16'd20161, 16'd7143, 16'd16505, 16'd15206, 16'd65299, 16'd9323, 16'd25737, 16'd7108});
	test_expansion(128'h325f97aeee5e3ff4c04c50b85d021a8f, {16'd62941, 16'd22867, 16'd28366, 16'd16800, 16'd58653, 16'd14523, 16'd1522, 16'd26967, 16'd56884, 16'd53427, 16'd7801, 16'd60565, 16'd40439, 16'd22129, 16'd47856, 16'd19694, 16'd25538, 16'd19319, 16'd58611, 16'd51101, 16'd12353, 16'd50843, 16'd42765, 16'd28015, 16'd30461, 16'd56402});
	test_expansion(128'ha00b2c9888ecd418339c4bca6ad4769a, {16'd39872, 16'd35304, 16'd60895, 16'd37176, 16'd55868, 16'd7256, 16'd47959, 16'd40003, 16'd18614, 16'd27304, 16'd20949, 16'd17236, 16'd54404, 16'd15530, 16'd21365, 16'd48006, 16'd52538, 16'd42336, 16'd22205, 16'd36401, 16'd21978, 16'd58087, 16'd55912, 16'd31076, 16'd42347, 16'd27524});
	test_expansion(128'h9c2c95d32f28707156be0529743d01be, {16'd61575, 16'd36402, 16'd11727, 16'd43758, 16'd47866, 16'd4109, 16'd30177, 16'd57492, 16'd59172, 16'd29773, 16'd57741, 16'd5335, 16'd37347, 16'd377, 16'd60675, 16'd22489, 16'd51647, 16'd58786, 16'd11236, 16'd3576, 16'd5272, 16'd62317, 16'd61680, 16'd28841, 16'd17568, 16'd57848});
	test_expansion(128'hde422c0eb6905a0abb92d432421fb2b9, {16'd41276, 16'd23558, 16'd4493, 16'd6576, 16'd2668, 16'd12269, 16'd49253, 16'd20047, 16'd64435, 16'd54787, 16'd23996, 16'd33829, 16'd8617, 16'd53819, 16'd42744, 16'd22827, 16'd57145, 16'd20353, 16'd35133, 16'd9483, 16'd20274, 16'd6005, 16'd14175, 16'd37669, 16'd2631, 16'd52265});
	test_expansion(128'h93ff708a8b13bd9af19f4cd145ac75d6, {16'd7298, 16'd63440, 16'd40542, 16'd23609, 16'd30222, 16'd54460, 16'd28978, 16'd13992, 16'd40067, 16'd22243, 16'd34592, 16'd5966, 16'd17911, 16'd44473, 16'd7816, 16'd25852, 16'd50764, 16'd32001, 16'd22720, 16'd40467, 16'd30339, 16'd40745, 16'd63369, 16'd38745, 16'd36247, 16'd361});
	test_expansion(128'hdd467f8e29fe343ae3dc84a63ab99c2b, {16'd59260, 16'd16360, 16'd12115, 16'd23362, 16'd36134, 16'd23604, 16'd58253, 16'd37865, 16'd20619, 16'd36346, 16'd2707, 16'd36541, 16'd6691, 16'd11966, 16'd58667, 16'd40528, 16'd58648, 16'd38393, 16'd7647, 16'd27166, 16'd10936, 16'd26236, 16'd25577, 16'd42619, 16'd54810, 16'd11116});
	test_expansion(128'h4a8ec42a6454b12705734f5cd2b0378d, {16'd17715, 16'd15258, 16'd29245, 16'd42032, 16'd59000, 16'd20881, 16'd24027, 16'd64998, 16'd19503, 16'd27707, 16'd18772, 16'd21523, 16'd6038, 16'd60249, 16'd1224, 16'd44331, 16'd37159, 16'd61451, 16'd13197, 16'd42490, 16'd35603, 16'd1306, 16'd32463, 16'd16268, 16'd37341, 16'd60972});
	test_expansion(128'h9cbd9bc7b20cf9d80ee2cdeb842d596a, {16'd21483, 16'd61119, 16'd36145, 16'd64734, 16'd6125, 16'd49177, 16'd50588, 16'd3732, 16'd47813, 16'd30980, 16'd33662, 16'd44705, 16'd47834, 16'd20849, 16'd1150, 16'd64210, 16'd47688, 16'd11133, 16'd30675, 16'd57967, 16'd59338, 16'd18575, 16'd18786, 16'd32280, 16'd26717, 16'd43547});
	test_expansion(128'h803bc6ce9902d3413e4ec441afa9d685, {16'd15307, 16'd39247, 16'd44268, 16'd38167, 16'd64035, 16'd45629, 16'd8234, 16'd27487, 16'd28500, 16'd4174, 16'd21623, 16'd6428, 16'd19993, 16'd61037, 16'd18778, 16'd15982, 16'd48382, 16'd38930, 16'd59651, 16'd63043, 16'd42362, 16'd39844, 16'd53369, 16'd32018, 16'd9509, 16'd428});
	test_expansion(128'h54ef1b2c7946869545275d863744b972, {16'd8938, 16'd41958, 16'd65195, 16'd62614, 16'd34200, 16'd45653, 16'd37890, 16'd14371, 16'd45125, 16'd8578, 16'd12503, 16'd45376, 16'd12311, 16'd49904, 16'd29894, 16'd60095, 16'd34418, 16'd45289, 16'd35863, 16'd8498, 16'd806, 16'd5210, 16'd50003, 16'd33381, 16'd3315, 16'd50521});
	test_expansion(128'h370d6458f231c3c07c026b7e488b8718, {16'd9270, 16'd47082, 16'd3953, 16'd8078, 16'd46869, 16'd1683, 16'd56992, 16'd46958, 16'd1105, 16'd29072, 16'd20690, 16'd29131, 16'd12469, 16'd44079, 16'd37497, 16'd14190, 16'd5503, 16'd56683, 16'd52339, 16'd34739, 16'd24087, 16'd29470, 16'd30880, 16'd28555, 16'd39926, 16'd35663});
	test_expansion(128'h72116f5d1c3ce9d6adcb1ee5de31d84d, {16'd49111, 16'd60109, 16'd18501, 16'd16392, 16'd13489, 16'd31430, 16'd50444, 16'd63948, 16'd61465, 16'd16321, 16'd52333, 16'd9292, 16'd33082, 16'd11942, 16'd12768, 16'd39319, 16'd36735, 16'd9481, 16'd21951, 16'd53347, 16'd5766, 16'd8111, 16'd63254, 16'd46583, 16'd13063, 16'd62382});
	test_expansion(128'h559c61ed696eb361947e80c649fa39e5, {16'd5883, 16'd1262, 16'd26146, 16'd4811, 16'd2727, 16'd40434, 16'd42048, 16'd61017, 16'd17693, 16'd10989, 16'd38041, 16'd40628, 16'd36291, 16'd938, 16'd15187, 16'd64642, 16'd29455, 16'd16495, 16'd10328, 16'd11332, 16'd15596, 16'd10972, 16'd63832, 16'd22321, 16'd57715, 16'd1897});
	test_expansion(128'hada92c65a0e06589807c934f2ffefd5f, {16'd12548, 16'd65510, 16'd39246, 16'd40343, 16'd10792, 16'd6763, 16'd42319, 16'd59474, 16'd48466, 16'd64412, 16'd28185, 16'd60710, 16'd65054, 16'd18364, 16'd59979, 16'd25547, 16'd51126, 16'd56437, 16'd32754, 16'd17690, 16'd50110, 16'd63733, 16'd64607, 16'd29814, 16'd14018, 16'd21757});
	test_expansion(128'hfdf788307a5b347661e52d57866590a4, {16'd35737, 16'd29474, 16'd14655, 16'd65248, 16'd56556, 16'd14645, 16'd39476, 16'd22213, 16'd23929, 16'd32966, 16'd30813, 16'd2305, 16'd8536, 16'd45097, 16'd21648, 16'd53329, 16'd13971, 16'd64279, 16'd44158, 16'd30770, 16'd25009, 16'd42286, 16'd28493, 16'd25545, 16'd6192, 16'd26590});
	test_expansion(128'hcbb5640ae79345c4f8ee06483d2f342e, {16'd50803, 16'd31045, 16'd35678, 16'd33614, 16'd31955, 16'd4155, 16'd56582, 16'd5593, 16'd61251, 16'd15344, 16'd53218, 16'd64032, 16'd59488, 16'd49573, 16'd13852, 16'd55184, 16'd40874, 16'd58217, 16'd31089, 16'd41408, 16'd12153, 16'd35795, 16'd28818, 16'd42350, 16'd43112, 16'd16104});
	test_expansion(128'h2e79c12e7a0051c4b640974f6c12b7e7, {16'd8272, 16'd31574, 16'd28329, 16'd3191, 16'd58859, 16'd28912, 16'd59116, 16'd41744, 16'd24888, 16'd28605, 16'd29073, 16'd49888, 16'd10927, 16'd31646, 16'd9501, 16'd2262, 16'd52572, 16'd56636, 16'd62784, 16'd63806, 16'd55089, 16'd17587, 16'd47854, 16'd23471, 16'd43185, 16'd43042});
	test_expansion(128'h279760e44496aa20afede2c87fe80adc, {16'd3507, 16'd45080, 16'd795, 16'd18401, 16'd55502, 16'd10186, 16'd24999, 16'd463, 16'd35298, 16'd44331, 16'd28703, 16'd23337, 16'd63221, 16'd63890, 16'd55558, 16'd37526, 16'd12506, 16'd57499, 16'd1624, 16'd48364, 16'd65206, 16'd31550, 16'd13926, 16'd1405, 16'd59317, 16'd35604});
	test_expansion(128'h972d06eb79a88b54f4424be065a85f56, {16'd57083, 16'd30279, 16'd61800, 16'd39240, 16'd40810, 16'd31462, 16'd51932, 16'd62172, 16'd43754, 16'd61947, 16'd41647, 16'd4303, 16'd18311, 16'd62410, 16'd45516, 16'd6120, 16'd58586, 16'd33574, 16'd41349, 16'd60992, 16'd20648, 16'd1319, 16'd64044, 16'd23991, 16'd25589, 16'd48903});
	test_expansion(128'h2bc0c8ba9dc80926abcb59c333743e89, {16'd64622, 16'd43274, 16'd18534, 16'd15348, 16'd34315, 16'd47140, 16'd22623, 16'd14108, 16'd1911, 16'd2770, 16'd32509, 16'd13759, 16'd9939, 16'd48385, 16'd24017, 16'd45983, 16'd38867, 16'd18797, 16'd50333, 16'd12463, 16'd7615, 16'd56548, 16'd27948, 16'd13918, 16'd65080, 16'd43150});
	test_expansion(128'h862fbed2374644aa1a1e914075c03569, {16'd52468, 16'd48687, 16'd55028, 16'd50687, 16'd16008, 16'd62792, 16'd10108, 16'd12694, 16'd3557, 16'd8772, 16'd22236, 16'd34823, 16'd43172, 16'd61396, 16'd48274, 16'd52820, 16'd48149, 16'd20505, 16'd16728, 16'd14981, 16'd61831, 16'd13254, 16'd15528, 16'd22574, 16'd41529, 16'd5384});
	test_expansion(128'hf5681888628f35277b8ed6dfb87b724a, {16'd45331, 16'd60592, 16'd37277, 16'd54611, 16'd42910, 16'd27789, 16'd26268, 16'd50439, 16'd59046, 16'd8196, 16'd5255, 16'd3112, 16'd42506, 16'd46916, 16'd21793, 16'd46926, 16'd44235, 16'd57540, 16'd33347, 16'd26711, 16'd12829, 16'd44, 16'd42557, 16'd62698, 16'd45720, 16'd15756});
	test_expansion(128'hc666f08f09a6dd77735c6d99f8a199d0, {16'd4372, 16'd3597, 16'd48241, 16'd45578, 16'd21647, 16'd53662, 16'd57954, 16'd15601, 16'd15637, 16'd3617, 16'd49022, 16'd62425, 16'd4716, 16'd26630, 16'd18409, 16'd44564, 16'd17197, 16'd18425, 16'd12794, 16'd28980, 16'd1842, 16'd50929, 16'd32875, 16'd35766, 16'd404, 16'd24116});
	test_expansion(128'h96872e98a7baae5faabf5b1c3357ac2d, {16'd16036, 16'd49601, 16'd33522, 16'd32035, 16'd60089, 16'd317, 16'd26081, 16'd7732, 16'd33164, 16'd24423, 16'd23578, 16'd57431, 16'd5423, 16'd55984, 16'd19487, 16'd25309, 16'd40619, 16'd38049, 16'd17082, 16'd50657, 16'd23080, 16'd11820, 16'd2776, 16'd54931, 16'd31266, 16'd53747});
	test_expansion(128'ha2c35f2b526d123d29bdbeeceb018629, {16'd32372, 16'd24535, 16'd27193, 16'd37991, 16'd52658, 16'd20222, 16'd31715, 16'd30624, 16'd24114, 16'd29817, 16'd32077, 16'd48460, 16'd12296, 16'd24867, 16'd21117, 16'd17952, 16'd39042, 16'd32746, 16'd15393, 16'd33597, 16'd58766, 16'd63722, 16'd65531, 16'd16237, 16'd7077, 16'd2109});
	test_expansion(128'hfdab1c8b9be06bc2bdbb0f5baed38241, {16'd52335, 16'd31003, 16'd6664, 16'd60492, 16'd13403, 16'd15779, 16'd22333, 16'd22774, 16'd60000, 16'd15255, 16'd56959, 16'd54973, 16'd1644, 16'd35114, 16'd13358, 16'd62654, 16'd8280, 16'd29951, 16'd32051, 16'd37996, 16'd30848, 16'd61865, 16'd28280, 16'd31563, 16'd31024, 16'd61665});
	test_expansion(128'h7e25ce7421ab7326a73d4d276f1ae32a, {16'd61188, 16'd49818, 16'd54843, 16'd40715, 16'd61321, 16'd60328, 16'd17129, 16'd34470, 16'd39111, 16'd13469, 16'd21203, 16'd19254, 16'd31558, 16'd22160, 16'd60234, 16'd12205, 16'd56100, 16'd54349, 16'd49521, 16'd37900, 16'd54836, 16'd38021, 16'd59901, 16'd49937, 16'd10565, 16'd50956});
	test_expansion(128'h56b116f72ca52eec0c58e729c4404d34, {16'd20183, 16'd26746, 16'd19733, 16'd906, 16'd55268, 16'd46397, 16'd18322, 16'd14390, 16'd36099, 16'd15689, 16'd10338, 16'd40760, 16'd54006, 16'd32585, 16'd39658, 16'd10415, 16'd8863, 16'd1585, 16'd60116, 16'd29186, 16'd21096, 16'd48141, 16'd7545, 16'd44871, 16'd28880, 16'd21702});
	test_expansion(128'h830243d6c0a8ff85220dec2d01d061e0, {16'd26556, 16'd53592, 16'd65403, 16'd10162, 16'd23972, 16'd3019, 16'd8944, 16'd44499, 16'd89, 16'd15530, 16'd10203, 16'd20864, 16'd47533, 16'd32255, 16'd39364, 16'd62070, 16'd4881, 16'd56207, 16'd63955, 16'd12242, 16'd144, 16'd37215, 16'd51166, 16'd57293, 16'd278, 16'd24053});
	test_expansion(128'hd5b31ec01ff4d697510287931f06146e, {16'd13952, 16'd33164, 16'd11839, 16'd40525, 16'd3295, 16'd57228, 16'd55986, 16'd11511, 16'd35427, 16'd32974, 16'd15486, 16'd7756, 16'd59169, 16'd30488, 16'd49871, 16'd2207, 16'd10630, 16'd62343, 16'd12373, 16'd51782, 16'd39293, 16'd10345, 16'd46855, 16'd18724, 16'd52312, 16'd51426});
	test_expansion(128'h56a79f1fa4eb7e2897a932ad2db94731, {16'd61006, 16'd55398, 16'd8265, 16'd26062, 16'd7904, 16'd64306, 16'd48298, 16'd16805, 16'd5254, 16'd16176, 16'd55139, 16'd57196, 16'd13478, 16'd6845, 16'd33450, 16'd11315, 16'd35376, 16'd43241, 16'd19919, 16'd21761, 16'd42244, 16'd17241, 16'd28283, 16'd13254, 16'd65131, 16'd33730});
	test_expansion(128'ha59a4425bacd0742938bf90e8687a6a4, {16'd13314, 16'd19884, 16'd50441, 16'd55389, 16'd60880, 16'd46221, 16'd7019, 16'd42841, 16'd4656, 16'd2982, 16'd44359, 16'd4769, 16'd15066, 16'd59105, 16'd45284, 16'd21263, 16'd30748, 16'd21462, 16'd28165, 16'd22170, 16'd1526, 16'd36874, 16'd27559, 16'd11043, 16'd53469, 16'd5037});
	test_expansion(128'h7be3ea68dc2e57c6eec0aa140de5e226, {16'd9837, 16'd55099, 16'd32324, 16'd40852, 16'd31896, 16'd34799, 16'd59988, 16'd12446, 16'd57561, 16'd55770, 16'd44434, 16'd1208, 16'd53407, 16'd13192, 16'd58497, 16'd18915, 16'd34544, 16'd9372, 16'd23080, 16'd36382, 16'd8489, 16'd36615, 16'd9418, 16'd3817, 16'd9207, 16'd2482});
	test_expansion(128'h1a601aeb621038a30dbbdc897344b1b8, {16'd18672, 16'd45390, 16'd60110, 16'd42680, 16'd35879, 16'd38236, 16'd47950, 16'd9610, 16'd32420, 16'd42800, 16'd53259, 16'd20698, 16'd28354, 16'd41766, 16'd13336, 16'd25691, 16'd65535, 16'd5706, 16'd45823, 16'd4550, 16'd38460, 16'd841, 16'd7230, 16'd45250, 16'd58623, 16'd12819});
	test_expansion(128'h262503bb625a84616ef31595f1b038cc, {16'd15603, 16'd3458, 16'd60759, 16'd41725, 16'd24135, 16'd37629, 16'd37367, 16'd25192, 16'd24837, 16'd32392, 16'd15413, 16'd41443, 16'd58574, 16'd19240, 16'd56779, 16'd63495, 16'd6464, 16'd2931, 16'd37639, 16'd39887, 16'd18822, 16'd41639, 16'd23551, 16'd57764, 16'd26088, 16'd13340});
	test_expansion(128'h5c4d19b6c5d326946e28590d090ccd24, {16'd40945, 16'd26325, 16'd16267, 16'd55129, 16'd52269, 16'd47954, 16'd19777, 16'd48518, 16'd16340, 16'd44664, 16'd35869, 16'd17951, 16'd36395, 16'd64164, 16'd11009, 16'd6858, 16'd5013, 16'd54991, 16'd41978, 16'd33629, 16'd26090, 16'd48141, 16'd52577, 16'd173, 16'd44460, 16'd21608});
	test_expansion(128'hf464b487f9369a11450f21faf5cdeca4, {16'd44704, 16'd13295, 16'd53836, 16'd46059, 16'd44434, 16'd49357, 16'd47965, 16'd11298, 16'd39540, 16'd25727, 16'd33415, 16'd45542, 16'd23484, 16'd24467, 16'd12923, 16'd23657, 16'd819, 16'd54979, 16'd13022, 16'd21798, 16'd4504, 16'd33553, 16'd6415, 16'd54082, 16'd15038, 16'd55328});
	test_expansion(128'h6b2fa4dbce12136b217e6d294ae4ae0b, {16'd61398, 16'd51400, 16'd23789, 16'd53310, 16'd19472, 16'd47576, 16'd44341, 16'd28255, 16'd18597, 16'd14165, 16'd30869, 16'd20726, 16'd21834, 16'd59948, 16'd20378, 16'd8645, 16'd56894, 16'd20731, 16'd36916, 16'd21464, 16'd19, 16'd27541, 16'd6278, 16'd4410, 16'd62413, 16'd55642});
	test_expansion(128'hfb3d2a6c49ae8ce435a0e8a9110f677f, {16'd22383, 16'd55999, 16'd63978, 16'd14208, 16'd46135, 16'd4999, 16'd9130, 16'd7588, 16'd15478, 16'd45430, 16'd15564, 16'd38838, 16'd32038, 16'd37751, 16'd10748, 16'd53023, 16'd14977, 16'd51515, 16'd15627, 16'd16248, 16'd11805, 16'd30031, 16'd15278, 16'd34027, 16'd20425, 16'd43050});
	test_expansion(128'h6256c1bb8688bef0c6ffd06e7820e988, {16'd48044, 16'd62076, 16'd15311, 16'd38678, 16'd37843, 16'd35821, 16'd41921, 16'd15379, 16'd15274, 16'd1056, 16'd31842, 16'd59185, 16'd37061, 16'd34008, 16'd45215, 16'd10837, 16'd13135, 16'd12738, 16'd26577, 16'd41727, 16'd37344, 16'd61029, 16'd20095, 16'd9342, 16'd18674, 16'd48937});
	test_expansion(128'he75eaa2ffaba29b87d0e7cb41cabd5fd, {16'd8500, 16'd1014, 16'd17640, 16'd44123, 16'd23333, 16'd25339, 16'd62905, 16'd54639, 16'd61620, 16'd13284, 16'd56459, 16'd19073, 16'd2154, 16'd8154, 16'd60218, 16'd64004, 16'd406, 16'd60432, 16'd18292, 16'd29398, 16'd60575, 16'd15909, 16'd55725, 16'd24581, 16'd41413, 16'd51223});
	test_expansion(128'h110346e6f2545d877bc3d3c6525a40f3, {16'd25325, 16'd33649, 16'd43682, 16'd1283, 16'd12401, 16'd25843, 16'd9237, 16'd64344, 16'd63347, 16'd12396, 16'd54974, 16'd36684, 16'd50942, 16'd32314, 16'd27471, 16'd41778, 16'd50306, 16'd42261, 16'd39052, 16'd57570, 16'd38340, 16'd26637, 16'd62595, 16'd57263, 16'd51644, 16'd15587});
	test_expansion(128'h2f635970acff070354c90af01f9cf6db, {16'd34796, 16'd28897, 16'd33560, 16'd62739, 16'd52358, 16'd24347, 16'd17301, 16'd11343, 16'd32991, 16'd20956, 16'd47618, 16'd7780, 16'd48538, 16'd23190, 16'd11079, 16'd20535, 16'd4921, 16'd31018, 16'd1954, 16'd58674, 16'd5078, 16'd34206, 16'd7574, 16'd41487, 16'd28480, 16'd17945});
	test_expansion(128'h19f2bde61b8739e99388b8d7442367ba, {16'd3880, 16'd19326, 16'd25239, 16'd30158, 16'd11879, 16'd41879, 16'd37632, 16'd55797, 16'd65512, 16'd47242, 16'd18279, 16'd15549, 16'd6272, 16'd11022, 16'd61274, 16'd7348, 16'd24567, 16'd54261, 16'd13119, 16'd19299, 16'd56757, 16'd8049, 16'd34954, 16'd32565, 16'd42289, 16'd26606});
	test_expansion(128'he5f60b8bd137cc6730b8c56ce7449738, {16'd49403, 16'd36683, 16'd31116, 16'd44698, 16'd31199, 16'd41228, 16'd4138, 16'd56964, 16'd47880, 16'd58090, 16'd27456, 16'd14754, 16'd50696, 16'd13015, 16'd37735, 16'd58047, 16'd314, 16'd52207, 16'd40503, 16'd49016, 16'd8834, 16'd17347, 16'd2535, 16'd14610, 16'd17920, 16'd41690});
	test_expansion(128'h16432fe728d10f3010674e8cfa242163, {16'd14766, 16'd64231, 16'd61405, 16'd28423, 16'd30397, 16'd18464, 16'd28769, 16'd54739, 16'd55754, 16'd30738, 16'd16145, 16'd59393, 16'd35000, 16'd3160, 16'd43324, 16'd28841, 16'd9824, 16'd35135, 16'd60678, 16'd40533, 16'd48718, 16'd53522, 16'd23083, 16'd28171, 16'd14884, 16'd60529});
	test_expansion(128'h7aa3555a3ae5326efac1b47d62497962, {16'd58454, 16'd22674, 16'd41262, 16'd459, 16'd6308, 16'd39888, 16'd48820, 16'd64333, 16'd50043, 16'd63101, 16'd45437, 16'd34996, 16'd43848, 16'd44799, 16'd21145, 16'd11047, 16'd64091, 16'd13956, 16'd37435, 16'd28474, 16'd3699, 16'd58072, 16'd28675, 16'd4145, 16'd46670, 16'd18681});
	test_expansion(128'h8073ceb5a5ed5156598e01c2c6e13983, {16'd8767, 16'd29730, 16'd65463, 16'd1534, 16'd58874, 16'd26674, 16'd7202, 16'd32823, 16'd61614, 16'd27023, 16'd22747, 16'd17827, 16'd26428, 16'd56059, 16'd53229, 16'd10865, 16'd59682, 16'd19404, 16'd32748, 16'd5460, 16'd37087, 16'd12478, 16'd58432, 16'd9119, 16'd49143, 16'd4295});
	test_expansion(128'h5902b92bee125db30abb4b31cae30ead, {16'd26883, 16'd32713, 16'd39666, 16'd56960, 16'd64813, 16'd13036, 16'd37554, 16'd34784, 16'd29586, 16'd15787, 16'd65022, 16'd25565, 16'd52927, 16'd33186, 16'd40287, 16'd36231, 16'd19360, 16'd14588, 16'd36393, 16'd63906, 16'd19926, 16'd23388, 16'd10064, 16'd50869, 16'd12263, 16'd10272});
	test_expansion(128'hb6892dab64f6727e46da7c4dca02426a, {16'd12943, 16'd51378, 16'd55820, 16'd20770, 16'd58660, 16'd34724, 16'd35487, 16'd30034, 16'd45064, 16'd3187, 16'd7555, 16'd7547, 16'd14723, 16'd53315, 16'd60762, 16'd13422, 16'd10622, 16'd14380, 16'd7946, 16'd57619, 16'd1113, 16'd3878, 16'd39558, 16'd36269, 16'd31193, 16'd65450});
	test_expansion(128'h7d305e4c74b1583ee106526efb4b37e6, {16'd16824, 16'd52757, 16'd18039, 16'd3996, 16'd40571, 16'd52870, 16'd18842, 16'd35046, 16'd23861, 16'd1749, 16'd10141, 16'd31625, 16'd64180, 16'd50699, 16'd24952, 16'd47573, 16'd64599, 16'd18831, 16'd10459, 16'd29147, 16'd3735, 16'd63904, 16'd22241, 16'd62385, 16'd5341, 16'd57369});
	test_expansion(128'hf71cc293de2807dc597fe230f4204478, {16'd60672, 16'd52893, 16'd15297, 16'd14289, 16'd56925, 16'd58511, 16'd28983, 16'd32102, 16'd57909, 16'd38611, 16'd47176, 16'd43147, 16'd10570, 16'd45258, 16'd60812, 16'd36844, 16'd50966, 16'd26923, 16'd43156, 16'd15911, 16'd33150, 16'd46199, 16'd24401, 16'd670, 16'd9135, 16'd35674});
	test_expansion(128'hbdaac6684b69e130c9f0aeb9fdd11266, {16'd6358, 16'd11773, 16'd47093, 16'd29345, 16'd27577, 16'd23270, 16'd9386, 16'd42790, 16'd15137, 16'd22282, 16'd27157, 16'd59555, 16'd58595, 16'd55245, 16'd54995, 16'd16143, 16'd30226, 16'd9923, 16'd3136, 16'd24045, 16'd16826, 16'd59787, 16'd25316, 16'd14241, 16'd11921, 16'd49759});
	test_expansion(128'h05b89445c79751807b0f9f69cc4fc1bd, {16'd6180, 16'd5160, 16'd20937, 16'd53295, 16'd61801, 16'd50934, 16'd18464, 16'd56616, 16'd2753, 16'd44181, 16'd22389, 16'd4934, 16'd9639, 16'd12225, 16'd26296, 16'd12552, 16'd59672, 16'd31364, 16'd45311, 16'd29420, 16'd1063, 16'd56002, 16'd21394, 16'd61705, 16'd28999, 16'd14481});
	test_expansion(128'hb8caa34f22e2205488e4c7e0c1ccb518, {16'd30662, 16'd25417, 16'd48781, 16'd48548, 16'd47424, 16'd35182, 16'd35960, 16'd27808, 16'd64460, 16'd10670, 16'd40428, 16'd39761, 16'd43001, 16'd19495, 16'd19296, 16'd48959, 16'd50445, 16'd64681, 16'd65438, 16'd64391, 16'd10630, 16'd34250, 16'd5151, 16'd32025, 16'd59870, 16'd7737});
	test_expansion(128'hdff8143fbe3b27840e1d18406a07b692, {16'd46311, 16'd24437, 16'd21401, 16'd25216, 16'd19096, 16'd2460, 16'd25272, 16'd63331, 16'd11118, 16'd6477, 16'd22427, 16'd25458, 16'd209, 16'd32894, 16'd2279, 16'd18874, 16'd25057, 16'd12464, 16'd39938, 16'd12051, 16'd51271, 16'd2201, 16'd63186, 16'd36192, 16'd26958, 16'd41747});
	test_expansion(128'h22bb466d105f45754c6f70c1da57a62d, {16'd59363, 16'd38790, 16'd25190, 16'd9253, 16'd37477, 16'd3129, 16'd55689, 16'd44223, 16'd3155, 16'd19025, 16'd5836, 16'd8438, 16'd12469, 16'd1904, 16'd54223, 16'd58639, 16'd46454, 16'd15502, 16'd4451, 16'd10887, 16'd57606, 16'd31957, 16'd37147, 16'd38298, 16'd38389, 16'd44408});
	test_expansion(128'h4e9f0d6dfc6435b9de982ccb08ef51fb, {16'd35372, 16'd18647, 16'd21294, 16'd52030, 16'd38325, 16'd41635, 16'd31339, 16'd3349, 16'd8932, 16'd26704, 16'd17161, 16'd42154, 16'd48115, 16'd57348, 16'd8937, 16'd480, 16'd22483, 16'd63675, 16'd55557, 16'd45444, 16'd12064, 16'd49814, 16'd14474, 16'd52966, 16'd2471, 16'd49318});
	test_expansion(128'hde80e59b033c9454f0e87d40e959519c, {16'd62455, 16'd34927, 16'd43854, 16'd5085, 16'd36838, 16'd13638, 16'd9629, 16'd37074, 16'd16178, 16'd33737, 16'd23582, 16'd48115, 16'd26950, 16'd33288, 16'd23402, 16'd44110, 16'd36805, 16'd18740, 16'd59170, 16'd34742, 16'd44141, 16'd6431, 16'd21160, 16'd13125, 16'd3909, 16'd26399});
	test_expansion(128'ha39cf75c7a0b1209459e825a6a0d535b, {16'd15337, 16'd25878, 16'd49296, 16'd33224, 16'd28419, 16'd47364, 16'd38980, 16'd12074, 16'd38280, 16'd6413, 16'd56299, 16'd65051, 16'd13178, 16'd4670, 16'd63193, 16'd5420, 16'd62202, 16'd28975, 16'd26607, 16'd31253, 16'd5727, 16'd5695, 16'd12660, 16'd46791, 16'd20699, 16'd35803});
	test_expansion(128'h85a5276b6163f017877fa82d16dc640c, {16'd15124, 16'd58739, 16'd1371, 16'd50208, 16'd53649, 16'd44217, 16'd49530, 16'd11998, 16'd53068, 16'd22761, 16'd9105, 16'd64629, 16'd56742, 16'd51475, 16'd55277, 16'd29379, 16'd40238, 16'd61988, 16'd10981, 16'd45562, 16'd11369, 16'd51185, 16'd2232, 16'd45094, 16'd3516, 16'd62354});
	test_expansion(128'h41ebbcc847460a302c36d657a599cf75, {16'd15169, 16'd63621, 16'd11606, 16'd12723, 16'd50260, 16'd46127, 16'd65111, 16'd23936, 16'd42265, 16'd37676, 16'd19180, 16'd65139, 16'd53092, 16'd36308, 16'd22824, 16'd6277, 16'd17662, 16'd42789, 16'd44879, 16'd46933, 16'd44649, 16'd65011, 16'd599, 16'd54362, 16'd53270, 16'd1249});
	test_expansion(128'h58a68db446a7e82ad39c0c4136fc43a5, {16'd14544, 16'd29548, 16'd33706, 16'd50441, 16'd20532, 16'd3836, 16'd58090, 16'd63060, 16'd50829, 16'd42781, 16'd53955, 16'd7905, 16'd55409, 16'd52060, 16'd30713, 16'd36696, 16'd34740, 16'd52965, 16'd1335, 16'd31324, 16'd5723, 16'd60228, 16'd49170, 16'd63005, 16'd52728, 16'd22738});
	test_expansion(128'hbf2d7b134121fe1df3efc6ec62a4874b, {16'd30362, 16'd47937, 16'd32697, 16'd56899, 16'd57744, 16'd37875, 16'd36175, 16'd10096, 16'd13286, 16'd28966, 16'd17040, 16'd45604, 16'd50606, 16'd37359, 16'd49239, 16'd9708, 16'd38089, 16'd57608, 16'd38096, 16'd55690, 16'd54732, 16'd23576, 16'd24506, 16'd15795, 16'd5506, 16'd45866});
	test_expansion(128'h082c2b1c83e1c3cf2bb5bc71a178e8a4, {16'd31611, 16'd44520, 16'd27642, 16'd18804, 16'd41713, 16'd63102, 16'd33287, 16'd22271, 16'd25743, 16'd16554, 16'd2497, 16'd20273, 16'd34754, 16'd18234, 16'd28052, 16'd50793, 16'd45633, 16'd12465, 16'd39412, 16'd11619, 16'd56604, 16'd23732, 16'd39117, 16'd2828, 16'd5220, 16'd62217});
	test_expansion(128'hf4eebe90fa8b3485bebfb45b75b84360, {16'd23143, 16'd2449, 16'd29264, 16'd6601, 16'd4349, 16'd33136, 16'd45202, 16'd55239, 16'd11707, 16'd56318, 16'd15636, 16'd51690, 16'd9563, 16'd39809, 16'd20995, 16'd62092, 16'd21254, 16'd36252, 16'd13359, 16'd600, 16'd44371, 16'd45272, 16'd4134, 16'd32934, 16'd48750, 16'd49449});
	test_expansion(128'h216dee5c41626ed87518e17377210ead, {16'd45533, 16'd50448, 16'd42543, 16'd23433, 16'd50764, 16'd19639, 16'd30476, 16'd61557, 16'd33498, 16'd45301, 16'd59866, 16'd24916, 16'd32675, 16'd45330, 16'd1517, 16'd2206, 16'd37634, 16'd12915, 16'd65136, 16'd37599, 16'd5098, 16'd45713, 16'd54716, 16'd40464, 16'd4581, 16'd22676});
	test_expansion(128'h10b1683085f05c963118a30a585a6676, {16'd45425, 16'd15344, 16'd602, 16'd55261, 16'd53112, 16'd43607, 16'd18092, 16'd20271, 16'd15349, 16'd6790, 16'd35145, 16'd10577, 16'd17396, 16'd36835, 16'd45718, 16'd51486, 16'd14721, 16'd10496, 16'd57812, 16'd3627, 16'd42773, 16'd52763, 16'd48151, 16'd23025, 16'd47162, 16'd3550});
	test_expansion(128'hf71d13f2a429be912da884149326d7a2, {16'd64397, 16'd32124, 16'd11776, 16'd341, 16'd15696, 16'd54420, 16'd57867, 16'd47303, 16'd52235, 16'd19805, 16'd19615, 16'd31461, 16'd56702, 16'd12840, 16'd19169, 16'd31464, 16'd20076, 16'd28828, 16'd11285, 16'd3242, 16'd55463, 16'd5745, 16'd29661, 16'd9296, 16'd56849, 16'd18720});
	test_expansion(128'h239fe3789d4991518592fc389f24a0fe, {16'd38510, 16'd52013, 16'd30946, 16'd34254, 16'd5522, 16'd8531, 16'd62073, 16'd19558, 16'd63952, 16'd62938, 16'd5671, 16'd56947, 16'd62449, 16'd63909, 16'd4396, 16'd2017, 16'd49257, 16'd58659, 16'd17374, 16'd9675, 16'd44519, 16'd48287, 16'd5335, 16'd33103, 16'd63541, 16'd50142});
	test_expansion(128'h152bd94bb23c11d72ea3b4c56a0fb790, {16'd5222, 16'd56841, 16'd6977, 16'd49556, 16'd47872, 16'd21779, 16'd38878, 16'd12047, 16'd50490, 16'd31315, 16'd64313, 16'd16168, 16'd25891, 16'd7328, 16'd18063, 16'd49292, 16'd25628, 16'd40267, 16'd41885, 16'd45823, 16'd63222, 16'd53465, 16'd41580, 16'd42103, 16'd52958, 16'd59581});
	test_expansion(128'h8ee40d4cd10f09f0f457ef5ab599bb83, {16'd62861, 16'd16830, 16'd6703, 16'd16373, 16'd1192, 16'd18537, 16'd28235, 16'd36288, 16'd45465, 16'd20437, 16'd39376, 16'd32406, 16'd761, 16'd2517, 16'd56362, 16'd43934, 16'd60266, 16'd18207, 16'd36990, 16'd18070, 16'd60734, 16'd51228, 16'd38708, 16'd35858, 16'd17879, 16'd60696});
	test_expansion(128'h98d3591ad758b3b6ace980266296c984, {16'd54848, 16'd46378, 16'd49525, 16'd58718, 16'd10966, 16'd8191, 16'd45024, 16'd50826, 16'd724, 16'd18358, 16'd223, 16'd31302, 16'd10544, 16'd13843, 16'd44043, 16'd47975, 16'd13701, 16'd62826, 16'd61830, 16'd20317, 16'd10157, 16'd49057, 16'd42245, 16'd10304, 16'd21820, 16'd58346});
	test_expansion(128'ha5ce3c4601b7807fd08f453611c0a77e, {16'd50710, 16'd51809, 16'd9116, 16'd56373, 16'd17844, 16'd44318, 16'd12124, 16'd50246, 16'd50898, 16'd49999, 16'd57889, 16'd37633, 16'd43482, 16'd46901, 16'd16756, 16'd44522, 16'd48643, 16'd50987, 16'd11915, 16'd52174, 16'd28200, 16'd59825, 16'd44659, 16'd10437, 16'd38711, 16'd18680});
	test_expansion(128'hbe1db1b7f60eb4fcb3c772ab33b30917, {16'd48625, 16'd57113, 16'd63619, 16'd57867, 16'd22294, 16'd27774, 16'd35315, 16'd6464, 16'd45694, 16'd46246, 16'd13899, 16'd29282, 16'd42121, 16'd48482, 16'd41999, 16'd29563, 16'd12425, 16'd38155, 16'd13778, 16'd9000, 16'd32596, 16'd3079, 16'd32081, 16'd26915, 16'd13971, 16'd6046});
	test_expansion(128'h18e1041dbc10a311d90776cdad7f2682, {16'd23584, 16'd22953, 16'd64757, 16'd15469, 16'd880, 16'd28835, 16'd49440, 16'd19804, 16'd15218, 16'd37386, 16'd13909, 16'd47971, 16'd51521, 16'd59052, 16'd32214, 16'd53404, 16'd40017, 16'd1539, 16'd31510, 16'd10130, 16'd50661, 16'd1309, 16'd63582, 16'd22656, 16'd10029, 16'd56105});
	test_expansion(128'h34f120d8a82b48b1a97e6b4591bc8c7c, {16'd16352, 16'd46207, 16'd61849, 16'd61065, 16'd28211, 16'd45487, 16'd9203, 16'd25499, 16'd61077, 16'd38088, 16'd18646, 16'd30891, 16'd1867, 16'd19553, 16'd34578, 16'd29901, 16'd47862, 16'd56772, 16'd18484, 16'd24861, 16'd28953, 16'd40815, 16'd34098, 16'd44803, 16'd47148, 16'd43436});
	test_expansion(128'hf94364ff3da46658dc4a442085b74098, {16'd9444, 16'd44611, 16'd47634, 16'd12716, 16'd52805, 16'd62974, 16'd26587, 16'd19446, 16'd57354, 16'd27983, 16'd38583, 16'd18287, 16'd32724, 16'd52612, 16'd53843, 16'd45553, 16'd49291, 16'd15597, 16'd54016, 16'd48010, 16'd18860, 16'd21649, 16'd7078, 16'd3992, 16'd21944, 16'd62553});
	test_expansion(128'hb084b3e3776de71a2c32293828648cd5, {16'd62190, 16'd17083, 16'd31366, 16'd38335, 16'd11363, 16'd42979, 16'd28900, 16'd9815, 16'd55773, 16'd974, 16'd35304, 16'd15795, 16'd64297, 16'd32424, 16'd33037, 16'd21520, 16'd53806, 16'd54457, 16'd15484, 16'd39997, 16'd63535, 16'd56840, 16'd5529, 16'd25304, 16'd59731, 16'd32443});
	test_expansion(128'h801cf79e35cc27889aad9f557a35758d, {16'd8118, 16'd30111, 16'd62127, 16'd52131, 16'd5054, 16'd31581, 16'd37994, 16'd22488, 16'd51310, 16'd64779, 16'd48815, 16'd35573, 16'd16257, 16'd29272, 16'd70, 16'd59831, 16'd47439, 16'd49498, 16'd43092, 16'd14859, 16'd5274, 16'd23029, 16'd29631, 16'd26680, 16'd52174, 16'd6813});
	test_expansion(128'h04eb8bcb4635f0b4a92bc098ffd69042, {16'd54987, 16'd18893, 16'd3736, 16'd46618, 16'd28069, 16'd4099, 16'd49781, 16'd22507, 16'd17253, 16'd1028, 16'd64639, 16'd63815, 16'd29568, 16'd65059, 16'd34162, 16'd48722, 16'd30115, 16'd26709, 16'd1282, 16'd52084, 16'd37280, 16'd7178, 16'd10963, 16'd42246, 16'd50234, 16'd9946});
	test_expansion(128'hac747b2b39e8b233648b3451f4e6311a, {16'd23826, 16'd3446, 16'd60306, 16'd17956, 16'd42646, 16'd50264, 16'd39185, 16'd63677, 16'd5386, 16'd45174, 16'd15140, 16'd49195, 16'd54862, 16'd48500, 16'd58153, 16'd5680, 16'd23415, 16'd60017, 16'd59783, 16'd55116, 16'd38957, 16'd63013, 16'd7709, 16'd17155, 16'd65323, 16'd23252});
	test_expansion(128'h3989166297b3a2175ef4c33dec6d48fd, {16'd54513, 16'd17022, 16'd19568, 16'd1071, 16'd22010, 16'd62797, 16'd12490, 16'd34112, 16'd38328, 16'd55934, 16'd35733, 16'd57485, 16'd24503, 16'd16994, 16'd3260, 16'd16708, 16'd15669, 16'd6005, 16'd46017, 16'd31398, 16'd62775, 16'd6013, 16'd45001, 16'd30324, 16'd7193, 16'd55242});
	test_expansion(128'he93632e5427375428b951f05b095b45a, {16'd23859, 16'd65399, 16'd42470, 16'd13562, 16'd58756, 16'd46602, 16'd44095, 16'd23260, 16'd34718, 16'd36817, 16'd39057, 16'd24644, 16'd60097, 16'd20818, 16'd18865, 16'd5489, 16'd43841, 16'd2378, 16'd16553, 16'd36661, 16'd6628, 16'd28893, 16'd23424, 16'd21597, 16'd62798, 16'd34444});
	test_expansion(128'hb7a2bc59dc9656b2b441875ecd9f3ff7, {16'd56025, 16'd63123, 16'd16799, 16'd59566, 16'd11278, 16'd11434, 16'd39372, 16'd6679, 16'd44288, 16'd10320, 16'd49990, 16'd50356, 16'd2461, 16'd61470, 16'd45489, 16'd4837, 16'd33208, 16'd49887, 16'd39300, 16'd58072, 16'd58696, 16'd19575, 16'd54372, 16'd988, 16'd17896, 16'd41580});
	test_expansion(128'h1e3fade2a5b1fbed8c7c1b2989395e2d, {16'd62152, 16'd13598, 16'd18474, 16'd29540, 16'd25684, 16'd1701, 16'd40286, 16'd42950, 16'd2357, 16'd28936, 16'd5262, 16'd25860, 16'd39038, 16'd36298, 16'd38972, 16'd50067, 16'd48812, 16'd8493, 16'd25084, 16'd11950, 16'd12577, 16'd5435, 16'd30414, 16'd45284, 16'd8269, 16'd64794});
	test_expansion(128'h062a3cbd9a5f4d0b36221c77e1b5daab, {16'd33572, 16'd50474, 16'd6880, 16'd6364, 16'd28656, 16'd1639, 16'd37378, 16'd51523, 16'd37804, 16'd62500, 16'd53140, 16'd28490, 16'd62352, 16'd55632, 16'd14720, 16'd43682, 16'd38368, 16'd36559, 16'd25665, 16'd50152, 16'd41198, 16'd54730, 16'd47058, 16'd28610, 16'd40237, 16'd14530});
	test_expansion(128'h12f4fdfb8c1506992352c6f566cf6695, {16'd28414, 16'd52424, 16'd19449, 16'd23591, 16'd27708, 16'd27857, 16'd15354, 16'd40963, 16'd54782, 16'd19449, 16'd51362, 16'd55166, 16'd15619, 16'd44462, 16'd40467, 16'd60678, 16'd4324, 16'd64757, 16'd3976, 16'd38731, 16'd1470, 16'd23138, 16'd60964, 16'd46345, 16'd46655, 16'd62943});
	test_expansion(128'hf70e124fbe28921ec119e4440a96beb2, {16'd60343, 16'd44210, 16'd27902, 16'd60092, 16'd42665, 16'd16173, 16'd4471, 16'd34264, 16'd9177, 16'd4275, 16'd19831, 16'd57013, 16'd38622, 16'd35063, 16'd28424, 16'd19963, 16'd47278, 16'd38245, 16'd27045, 16'd32186, 16'd57743, 16'd29204, 16'd35723, 16'd62488, 16'd50632, 16'd4305});
	test_expansion(128'hce47a205ebfa998a0103398461191c8e, {16'd12672, 16'd13180, 16'd48842, 16'd27471, 16'd10458, 16'd2098, 16'd62186, 16'd32280, 16'd3349, 16'd19660, 16'd56748, 16'd9821, 16'd18749, 16'd2164, 16'd45912, 16'd572, 16'd37674, 16'd47301, 16'd59589, 16'd1390, 16'd25873, 16'd59709, 16'd33363, 16'd20736, 16'd25440, 16'd21265});
	test_expansion(128'h9baa3e38154bc36e54556ea08cbf6b8d, {16'd14313, 16'd35026, 16'd38658, 16'd25020, 16'd11684, 16'd41738, 16'd11983, 16'd42902, 16'd8510, 16'd25474, 16'd31332, 16'd39509, 16'd62753, 16'd9203, 16'd59635, 16'd64595, 16'd41154, 16'd22593, 16'd53051, 16'd40513, 16'd15908, 16'd62247, 16'd29758, 16'd2063, 16'd7020, 16'd12753});
	test_expansion(128'h3f1da088b70d3f0982f2c13ad36a1367, {16'd46900, 16'd38148, 16'd49204, 16'd48806, 16'd3751, 16'd306, 16'd12470, 16'd53643, 16'd9487, 16'd64893, 16'd55812, 16'd21401, 16'd61053, 16'd57811, 16'd22768, 16'd41598, 16'd3111, 16'd54811, 16'd35221, 16'd56925, 16'd53383, 16'd63852, 16'd5036, 16'd12290, 16'd2966, 16'd41184});
	test_expansion(128'h9091018e915a46a434541f84521c8d5a, {16'd24521, 16'd51812, 16'd47091, 16'd1401, 16'd48040, 16'd12180, 16'd54864, 16'd5680, 16'd42041, 16'd14490, 16'd17173, 16'd54872, 16'd31000, 16'd2678, 16'd11386, 16'd46256, 16'd27326, 16'd43442, 16'd11497, 16'd27040, 16'd11984, 16'd6139, 16'd19495, 16'd53702, 16'd8959, 16'd54008});
	test_expansion(128'h2c3fe683c0d2a1d99858ac3e932b1014, {16'd38077, 16'd7315, 16'd42356, 16'd35035, 16'd55704, 16'd11586, 16'd58213, 16'd64161, 16'd42102, 16'd6232, 16'd19288, 16'd42227, 16'd6462, 16'd27213, 16'd48590, 16'd59767, 16'd485, 16'd53415, 16'd53871, 16'd41480, 16'd46288, 16'd25488, 16'd46381, 16'd51491, 16'd62099, 16'd49208});
	test_expansion(128'h6e63aaf77b01a65e41e4ee7272ec4672, {16'd17182, 16'd2546, 16'd23245, 16'd48385, 16'd4182, 16'd52155, 16'd60107, 16'd44183, 16'd5127, 16'd3038, 16'd15151, 16'd30219, 16'd24439, 16'd7494, 16'd64456, 16'd46103, 16'd4023, 16'd32311, 16'd22311, 16'd62955, 16'd41081, 16'd4649, 16'd33847, 16'd31626, 16'd14879, 16'd9906});
	test_expansion(128'hd81ef208b48e290f1ab17c839302be6c, {16'd24350, 16'd59459, 16'd37683, 16'd55164, 16'd50990, 16'd49615, 16'd65117, 16'd61012, 16'd55492, 16'd12825, 16'd17181, 16'd45879, 16'd43391, 16'd49739, 16'd18297, 16'd13676, 16'd55817, 16'd24371, 16'd39277, 16'd58910, 16'd16591, 16'd33003, 16'd6927, 16'd55690, 16'd23918, 16'd21003});
	test_expansion(128'h576d3000f93100ced44086f4d3f4b350, {16'd46742, 16'd36016, 16'd51214, 16'd31656, 16'd15725, 16'd36203, 16'd50292, 16'd42986, 16'd3656, 16'd44737, 16'd40649, 16'd56643, 16'd12809, 16'd54942, 16'd14057, 16'd60545, 16'd48663, 16'd9292, 16'd43371, 16'd25763, 16'd37010, 16'd18342, 16'd34144, 16'd18380, 16'd24330, 16'd16666});
	test_expansion(128'hd1f2a7a57fc864d7d8c0d88f8b9c851d, {16'd49390, 16'd59752, 16'd54287, 16'd57796, 16'd10028, 16'd61171, 16'd17806, 16'd38782, 16'd42677, 16'd56878, 16'd15817, 16'd64381, 16'd6069, 16'd27208, 16'd27772, 16'd29297, 16'd25342, 16'd15325, 16'd54674, 16'd53703, 16'd49688, 16'd12177, 16'd53204, 16'd45621, 16'd45833, 16'd30351});
	test_expansion(128'h3c255da537770cdf69a1c77fe57c0565, {16'd27014, 16'd22598, 16'd23248, 16'd51022, 16'd41976, 16'd55101, 16'd48071, 16'd33025, 16'd805, 16'd8308, 16'd43905, 16'd49874, 16'd35331, 16'd51815, 16'd5171, 16'd26294, 16'd7736, 16'd40856, 16'd46389, 16'd11187, 16'd47356, 16'd57691, 16'd10887, 16'd21314, 16'd30764, 16'd6964});
	test_expansion(128'hfc9c8e6793af52814d2eee5148e67073, {16'd9892, 16'd13888, 16'd11140, 16'd33826, 16'd27836, 16'd56517, 16'd43135, 16'd44051, 16'd19008, 16'd28074, 16'd29997, 16'd1834, 16'd46842, 16'd60291, 16'd37851, 16'd16478, 16'd20749, 16'd5833, 16'd50504, 16'd56806, 16'd59155, 16'd53187, 16'd31901, 16'd39272, 16'd55373, 16'd53197});
	test_expansion(128'h44b0cfda116e0d03f720650fa6d25aee, {16'd62641, 16'd7880, 16'd51952, 16'd53914, 16'd5217, 16'd13440, 16'd7455, 16'd41293, 16'd30575, 16'd48168, 16'd37926, 16'd45183, 16'd18219, 16'd39006, 16'd15433, 16'd18035, 16'd44311, 16'd60063, 16'd42665, 16'd7890, 16'd8053, 16'd28990, 16'd4102, 16'd17061, 16'd4166, 16'd978});
	test_expansion(128'h64d772998e2d12df4dd3b147fedd1be2, {16'd30577, 16'd4616, 16'd30571, 16'd19397, 16'd391, 16'd45532, 16'd35035, 16'd46074, 16'd31684, 16'd25137, 16'd40838, 16'd7512, 16'd26431, 16'd54224, 16'd33095, 16'd63370, 16'd55960, 16'd30348, 16'd30498, 16'd23593, 16'd40787, 16'd44378, 16'd3984, 16'd48338, 16'd52808, 16'd50643});
	test_expansion(128'h9628986e038ca775a6fc77ceb1ee6728, {16'd24120, 16'd12467, 16'd19701, 16'd32614, 16'd48339, 16'd34466, 16'd52067, 16'd12119, 16'd19595, 16'd27136, 16'd26287, 16'd44408, 16'd14795, 16'd32034, 16'd24330, 16'd46109, 16'd14260, 16'd35127, 16'd5088, 16'd35579, 16'd42849, 16'd2376, 16'd51237, 16'd12489, 16'd65333, 16'd19249});
	test_expansion(128'h5190d4edb1d7d15fcbddaac6018ec54f, {16'd51059, 16'd14274, 16'd41649, 16'd2813, 16'd55642, 16'd53179, 16'd57542, 16'd27321, 16'd52240, 16'd24633, 16'd60965, 16'd47126, 16'd24413, 16'd7335, 16'd50468, 16'd23648, 16'd9354, 16'd40534, 16'd9009, 16'd24378, 16'd23375, 16'd39858, 16'd6457, 16'd27371, 16'd19770, 16'd23111});
	test_expansion(128'h832e0c70fbb132f3b5ba2a4b2e08853e, {16'd41244, 16'd31101, 16'd50266, 16'd37303, 16'd31139, 16'd10532, 16'd54104, 16'd43494, 16'd34753, 16'd25107, 16'd51873, 16'd55023, 16'd50245, 16'd34464, 16'd53566, 16'd22757, 16'd35683, 16'd45300, 16'd50237, 16'd39626, 16'd771, 16'd16423, 16'd26216, 16'd46183, 16'd5739, 16'd26249});
	test_expansion(128'h6dba63fd350b2a4e188c8cfec626ba6e, {16'd24987, 16'd16040, 16'd31982, 16'd26634, 16'd16880, 16'd15044, 16'd40644, 16'd48732, 16'd39670, 16'd64468, 16'd40960, 16'd239, 16'd3741, 16'd31389, 16'd49813, 16'd33301, 16'd51971, 16'd14239, 16'd52325, 16'd40344, 16'd43143, 16'd40642, 16'd62043, 16'd39445, 16'd24577, 16'd61156});
	test_expansion(128'hbb418e383cb99e391743ffbb05ab8d54, {16'd28772, 16'd42217, 16'd20617, 16'd15629, 16'd24776, 16'd25466, 16'd42292, 16'd53233, 16'd58483, 16'd54931, 16'd8128, 16'd31946, 16'd37728, 16'd37009, 16'd21779, 16'd48177, 16'd59728, 16'd4700, 16'd53865, 16'd1485, 16'd33931, 16'd1076, 16'd30179, 16'd33643, 16'd57773, 16'd23261});
	test_expansion(128'h16a0d4a9259f562815b98a015a9baf39, {16'd10299, 16'd16365, 16'd13292, 16'd1890, 16'd60673, 16'd22602, 16'd34547, 16'd55534, 16'd53555, 16'd29099, 16'd46528, 16'd27555, 16'd27563, 16'd62814, 16'd39470, 16'd16247, 16'd59023, 16'd32321, 16'd47500, 16'd64995, 16'd5629, 16'd44172, 16'd28310, 16'd63377, 16'd43126, 16'd38883});
	test_expansion(128'hb093735bc82c4cfce523ef56c432fbce, {16'd40900, 16'd10719, 16'd50754, 16'd26897, 16'd26965, 16'd56374, 16'd61765, 16'd32841, 16'd42164, 16'd17527, 16'd5235, 16'd25590, 16'd55583, 16'd22128, 16'd14612, 16'd33590, 16'd35593, 16'd57005, 16'd27640, 16'd50999, 16'd55504, 16'd606, 16'd41711, 16'd15491, 16'd54493, 16'd1321});
	test_expansion(128'h5373bcf481beb529a3e06b0358a798f7, {16'd41515, 16'd19665, 16'd38732, 16'd37886, 16'd54628, 16'd57997, 16'd5720, 16'd34041, 16'd42580, 16'd4260, 16'd5049, 16'd55157, 16'd38349, 16'd15604, 16'd56004, 16'd40859, 16'd61461, 16'd20756, 16'd7115, 16'd27132, 16'd53156, 16'd3033, 16'd37202, 16'd59492, 16'd25037, 16'd34133});
	test_expansion(128'h4066cf70c95fb6e6182b24eacb19624b, {16'd36196, 16'd38635, 16'd29853, 16'd23224, 16'd56012, 16'd949, 16'd61221, 16'd20062, 16'd14781, 16'd2918, 16'd32253, 16'd14281, 16'd17991, 16'd7113, 16'd25220, 16'd63802, 16'd27313, 16'd13842, 16'd1024, 16'd13889, 16'd60279, 16'd55556, 16'd25125, 16'd38866, 16'd50288, 16'd17419});
	test_expansion(128'hab5c20d9fe790a5c89bd249d99313d83, {16'd15054, 16'd13661, 16'd30298, 16'd9194, 16'd15987, 16'd37644, 16'd52034, 16'd25048, 16'd29094, 16'd10095, 16'd56186, 16'd4462, 16'd18860, 16'd20329, 16'd57126, 16'd7677, 16'd46241, 16'd40831, 16'd30314, 16'd38820, 16'd33565, 16'd4631, 16'd60235, 16'd8270, 16'd11320, 16'd12558});
	test_expansion(128'h2c121716aca44457b842bb46324a0bce, {16'd59628, 16'd32333, 16'd47940, 16'd57903, 16'd13320, 16'd63249, 16'd14281, 16'd62065, 16'd14998, 16'd24894, 16'd4809, 16'd3227, 16'd40164, 16'd20271, 16'd39681, 16'd16909, 16'd1436, 16'd34303, 16'd6135, 16'd50650, 16'd61441, 16'd16427, 16'd16366, 16'd10589, 16'd37580, 16'd27421});
	test_expansion(128'h79fa53bfa0d8e66a1c16c824f0898313, {16'd46666, 16'd58217, 16'd43352, 16'd9307, 16'd25820, 16'd11972, 16'd21953, 16'd20160, 16'd16586, 16'd51813, 16'd24785, 16'd9266, 16'd61735, 16'd25047, 16'd20183, 16'd15869, 16'd56814, 16'd25099, 16'd27714, 16'd26051, 16'd15854, 16'd9507, 16'd12326, 16'd31900, 16'd15961, 16'd54501});
	test_expansion(128'h6e67a16664ca4f0d2470756f6f8ffebc, {16'd58305, 16'd45418, 16'd8114, 16'd35518, 16'd12759, 16'd5118, 16'd14648, 16'd38728, 16'd22187, 16'd60611, 16'd6470, 16'd60893, 16'd10680, 16'd37648, 16'd43533, 16'd6257, 16'd26356, 16'd2117, 16'd33303, 16'd36670, 16'd23549, 16'd25677, 16'd12949, 16'd53555, 16'd45459, 16'd996});
	test_expansion(128'h91bdbcb648a1bfd0912898c1dc9a8a64, {16'd55712, 16'd54144, 16'd53999, 16'd46927, 16'd65445, 16'd38929, 16'd27852, 16'd54402, 16'd44312, 16'd36664, 16'd973, 16'd11781, 16'd10158, 16'd54022, 16'd22814, 16'd51973, 16'd5634, 16'd35363, 16'd48352, 16'd826, 16'd52658, 16'd25439, 16'd64938, 16'd36401, 16'd43569, 16'd10480});
	test_expansion(128'hb5f33d11702634263817816c65b3b63d, {16'd12954, 16'd64159, 16'd65380, 16'd25639, 16'd2483, 16'd11627, 16'd26078, 16'd17689, 16'd21635, 16'd30992, 16'd55319, 16'd62510, 16'd16655, 16'd37270, 16'd28345, 16'd32977, 16'd11278, 16'd16204, 16'd25642, 16'd38858, 16'd20578, 16'd4261, 16'd21206, 16'd3979, 16'd32364, 16'd31595});
	test_expansion(128'h19ecb982d5447245f0f8e4fe4d078908, {16'd54832, 16'd33688, 16'd52946, 16'd24926, 16'd32333, 16'd22626, 16'd11056, 16'd49952, 16'd10783, 16'd60145, 16'd28936, 16'd65002, 16'd17706, 16'd2492, 16'd8807, 16'd20769, 16'd51739, 16'd34803, 16'd19221, 16'd59678, 16'd61286, 16'd26601, 16'd22131, 16'd25905, 16'd22572, 16'd16724});
	test_expansion(128'h09ccb0348c47b048a88e04823e0328e6, {16'd40373, 16'd46830, 16'd42881, 16'd64706, 16'd57706, 16'd41090, 16'd15022, 16'd62172, 16'd4448, 16'd54778, 16'd39297, 16'd41720, 16'd36258, 16'd40438, 16'd21757, 16'd55319, 16'd13260, 16'd16101, 16'd30229, 16'd25795, 16'd39707, 16'd41386, 16'd51958, 16'd37778, 16'd44502, 16'd8574});
	test_expansion(128'h109959e72f73abf76a72228081f028c7, {16'd7056, 16'd5169, 16'd47367, 16'd36088, 16'd61518, 16'd27404, 16'd15099, 16'd58252, 16'd56347, 16'd58265, 16'd25392, 16'd14941, 16'd27957, 16'd45384, 16'd1168, 16'd12146, 16'd13444, 16'd25473, 16'd32982, 16'd5895, 16'd62361, 16'd54202, 16'd23501, 16'd34378, 16'd44473, 16'd8010});
	test_expansion(128'h99b5645499ecf9b96f4bcc95b055d1f0, {16'd14817, 16'd32228, 16'd8318, 16'd59254, 16'd1253, 16'd32892, 16'd14173, 16'd26334, 16'd59967, 16'd44701, 16'd34212, 16'd38978, 16'd50199, 16'd3282, 16'd21234, 16'd54738, 16'd61296, 16'd25267, 16'd25931, 16'd27186, 16'd64422, 16'd5307, 16'd62287, 16'd30679, 16'd44063, 16'd32346});
	test_expansion(128'hef013af61c966e337378fca1db1073a9, {16'd14030, 16'd18407, 16'd56749, 16'd38844, 16'd42958, 16'd4413, 16'd51315, 16'd20914, 16'd33190, 16'd52800, 16'd13032, 16'd49790, 16'd18375, 16'd32306, 16'd29821, 16'd16351, 16'd36780, 16'd32925, 16'd50794, 16'd40322, 16'd30657, 16'd43369, 16'd54358, 16'd54480, 16'd35058, 16'd54031});
	test_expansion(128'hfba73357a4df80f23a2c20f86708560d, {16'd14224, 16'd64469, 16'd63656, 16'd4652, 16'd33495, 16'd28503, 16'd13399, 16'd37496, 16'd63595, 16'd56094, 16'd56712, 16'd38378, 16'd60781, 16'd49217, 16'd7617, 16'd17423, 16'd12927, 16'd10262, 16'd49556, 16'd18431, 16'd43447, 16'd28724, 16'd14271, 16'd56829, 16'd31802, 16'd3074});
	test_expansion(128'h36342e4a73f460f2348d3e9702029852, {16'd22664, 16'd2967, 16'd49347, 16'd32406, 16'd34853, 16'd58589, 16'd15878, 16'd16881, 16'd22938, 16'd24036, 16'd24005, 16'd53638, 16'd46402, 16'd38880, 16'd6394, 16'd52776, 16'd45801, 16'd12209, 16'd40010, 16'd15075, 16'd65122, 16'd25231, 16'd37914, 16'd14139, 16'd34419, 16'd61907});
	test_expansion(128'hb8a72372ea9ea8c766bc361d63e48a10, {16'd13055, 16'd64733, 16'd56793, 16'd11136, 16'd9351, 16'd26453, 16'd64782, 16'd18341, 16'd64120, 16'd26508, 16'd2939, 16'd65415, 16'd39954, 16'd9310, 16'd13156, 16'd2877, 16'd41962, 16'd25372, 16'd33173, 16'd52500, 16'd43707, 16'd48406, 16'd14296, 16'd14645, 16'd61252, 16'd45825});
	test_expansion(128'h492aff675b64a9fc8c62764712d16721, {16'd39213, 16'd50742, 16'd3366, 16'd61719, 16'd25400, 16'd15545, 16'd50537, 16'd64346, 16'd43649, 16'd56959, 16'd52480, 16'd57733, 16'd22866, 16'd11678, 16'd18430, 16'd35207, 16'd23060, 16'd20057, 16'd21089, 16'd12191, 16'd46157, 16'd8783, 16'd40364, 16'd22986, 16'd38053, 16'd60885});
	test_expansion(128'haca0e1ce9a0db96d7892aecae3753445, {16'd3476, 16'd42634, 16'd27535, 16'd28541, 16'd54673, 16'd54882, 16'd15620, 16'd4574, 16'd33109, 16'd1421, 16'd55075, 16'd22222, 16'd48597, 16'd9917, 16'd25688, 16'd38276, 16'd29439, 16'd12636, 16'd60718, 16'd43020, 16'd31135, 16'd13983, 16'd17522, 16'd61511, 16'd49673, 16'd10661});
	test_expansion(128'h284ed811bece39eed9b5afdbed2a0d3e, {16'd8965, 16'd39497, 16'd11299, 16'd28357, 16'd49550, 16'd46139, 16'd19362, 16'd34330, 16'd27990, 16'd7107, 16'd62031, 16'd163, 16'd54502, 16'd35930, 16'd17884, 16'd58350, 16'd51869, 16'd60931, 16'd19992, 16'd62371, 16'd58928, 16'd19056, 16'd46098, 16'd45079, 16'd20547, 16'd7412});
	test_expansion(128'h8a9253b5e1023f9cf720deaa02a4976d, {16'd55501, 16'd1466, 16'd21618, 16'd19016, 16'd46652, 16'd20517, 16'd7439, 16'd11115, 16'd26677, 16'd32375, 16'd2038, 16'd31453, 16'd46870, 16'd12687, 16'd40514, 16'd55047, 16'd54136, 16'd35438, 16'd29942, 16'd40528, 16'd59992, 16'd36558, 16'd2853, 16'd56726, 16'd6822, 16'd21250});
	test_expansion(128'h272e156161b388c2d836c84dcc99cf84, {16'd38296, 16'd20755, 16'd7101, 16'd54301, 16'd35537, 16'd43035, 16'd57967, 16'd4010, 16'd37523, 16'd2772, 16'd850, 16'd36177, 16'd33125, 16'd33459, 16'd39232, 16'd60227, 16'd37243, 16'd41976, 16'd50525, 16'd20851, 16'd55843, 16'd15217, 16'd37070, 16'd15525, 16'd9044, 16'd2835});
	test_expansion(128'hd934ebe854320dca07e9119d9043f780, {16'd22654, 16'd3250, 16'd64852, 16'd22617, 16'd56529, 16'd40832, 16'd52080, 16'd62206, 16'd33459, 16'd39675, 16'd11181, 16'd27585, 16'd45171, 16'd14972, 16'd2684, 16'd13814, 16'd16380, 16'd3607, 16'd32817, 16'd33766, 16'd32635, 16'd5538, 16'd27177, 16'd37565, 16'd44983, 16'd16141});
	test_expansion(128'hacee07dd2eb92aec25ed6678bc45e186, {16'd45679, 16'd59165, 16'd54534, 16'd20175, 16'd22641, 16'd59895, 16'd18250, 16'd43303, 16'd20081, 16'd3299, 16'd6711, 16'd29202, 16'd21926, 16'd2836, 16'd37848, 16'd1352, 16'd23671, 16'd22179, 16'd46194, 16'd63419, 16'd61757, 16'd37449, 16'd64129, 16'd19822, 16'd30574, 16'd7131});
	test_expansion(128'hd370fb22eabe0e277d2adbbb030c5bc6, {16'd7470, 16'd54744, 16'd5166, 16'd40283, 16'd52644, 16'd37557, 16'd13503, 16'd60538, 16'd36078, 16'd13749, 16'd3201, 16'd49058, 16'd40104, 16'd15748, 16'd56957, 16'd55539, 16'd49870, 16'd31932, 16'd55772, 16'd47203, 16'd8589, 16'd49806, 16'd11080, 16'd8275, 16'd11393, 16'd61548});
	test_expansion(128'hed147d93420cf6bc8fafa82269e5cf3c, {16'd46687, 16'd26463, 16'd20030, 16'd17373, 16'd46594, 16'd52231, 16'd32659, 16'd50289, 16'd47938, 16'd3396, 16'd63864, 16'd51694, 16'd58841, 16'd9162, 16'd37356, 16'd43835, 16'd49140, 16'd14594, 16'd61263, 16'd58403, 16'd25243, 16'd59266, 16'd47331, 16'd28864, 16'd63112, 16'd53570});
	test_expansion(128'hf1e48cf02277791bdfbd46b4ab007d74, {16'd48994, 16'd49464, 16'd15084, 16'd48150, 16'd35131, 16'd35818, 16'd63328, 16'd25215, 16'd53638, 16'd36506, 16'd19904, 16'd27891, 16'd16624, 16'd45645, 16'd7706, 16'd54511, 16'd55121, 16'd41839, 16'd11222, 16'd54202, 16'd46748, 16'd35773, 16'd6503, 16'd21673, 16'd60769, 16'd35440});
	test_expansion(128'h76fb593a59a6ba6ad3c9d27fa99cef5f, {16'd50230, 16'd50397, 16'd4813, 16'd37302, 16'd3676, 16'd5522, 16'd15338, 16'd14871, 16'd11266, 16'd31230, 16'd40818, 16'd45468, 16'd14643, 16'd34957, 16'd57232, 16'd38853, 16'd18296, 16'd53924, 16'd12967, 16'd7584, 16'd28592, 16'd63707, 16'd6655, 16'd30959, 16'd14766, 16'd5159});
	test_expansion(128'h594a708496cbcbb19f2b65109ea1cc17, {16'd24661, 16'd34241, 16'd502, 16'd50946, 16'd59319, 16'd32819, 16'd13132, 16'd59331, 16'd17654, 16'd38294, 16'd59689, 16'd24958, 16'd61941, 16'd49194, 16'd19645, 16'd8533, 16'd29253, 16'd39090, 16'd14994, 16'd43864, 16'd14869, 16'd28711, 16'd48919, 16'd11475, 16'd12988, 16'd54875});
	test_expansion(128'hdd9884f4b53c5532604427af2dd5de7d, {16'd43769, 16'd25911, 16'd16503, 16'd46559, 16'd15143, 16'd52519, 16'd22727, 16'd56396, 16'd5884, 16'd1157, 16'd36581, 16'd31030, 16'd41014, 16'd41474, 16'd16403, 16'd18439, 16'd24933, 16'd21458, 16'd65023, 16'd30460, 16'd34338, 16'd14313, 16'd43888, 16'd60684, 16'd25259, 16'd16815});
	test_expansion(128'hbf5cb34b6ebf89eb5adf1d1f60ed3afb, {16'd44700, 16'd51482, 16'd62935, 16'd38260, 16'd53984, 16'd20404, 16'd2239, 16'd44994, 16'd7294, 16'd3146, 16'd14541, 16'd19094, 16'd7468, 16'd17224, 16'd10373, 16'd57778, 16'd31228, 16'd54227, 16'd8742, 16'd59290, 16'd27697, 16'd39268, 16'd26306, 16'd26072, 16'd2469, 16'd53835});
	test_expansion(128'hc41b1b1c28cfbc22c600c04979ce96cc, {16'd55136, 16'd47980, 16'd7478, 16'd65045, 16'd25939, 16'd35343, 16'd24911, 16'd36320, 16'd28311, 16'd7681, 16'd43117, 16'd28575, 16'd53293, 16'd25132, 16'd32898, 16'd60462, 16'd19413, 16'd26204, 16'd41953, 16'd23317, 16'd55151, 16'd29094, 16'd26913, 16'd63339, 16'd26579, 16'd26502});
	test_expansion(128'hf3e5a180653ffcea90ebe2c50e3ac231, {16'd14133, 16'd5277, 16'd62376, 16'd24711, 16'd23218, 16'd64834, 16'd23320, 16'd63641, 16'd48106, 16'd51712, 16'd17750, 16'd30905, 16'd22, 16'd57421, 16'd8726, 16'd40139, 16'd5205, 16'd25268, 16'd57393, 16'd29407, 16'd27784, 16'd25458, 16'd10362, 16'd12528, 16'd3373, 16'd18925});
	test_expansion(128'h7ef5fddad4ce7233c466c509566a18f3, {16'd30569, 16'd20294, 16'd25097, 16'd18458, 16'd12524, 16'd57729, 16'd57932, 16'd9203, 16'd13319, 16'd42838, 16'd52626, 16'd61557, 16'd3664, 16'd29962, 16'd2656, 16'd49909, 16'd16957, 16'd43561, 16'd65151, 16'd62134, 16'd63078, 16'd18330, 16'd7397, 16'd34222, 16'd26134, 16'd19340});
	test_expansion(128'h4b4b0a01dc4b1ea45359c85e11cb1064, {16'd28439, 16'd18633, 16'd443, 16'd30096, 16'd24469, 16'd30237, 16'd59082, 16'd18857, 16'd33116, 16'd37920, 16'd41816, 16'd32161, 16'd50906, 16'd119, 16'd44408, 16'd51937, 16'd18947, 16'd64469, 16'd35921, 16'd38173, 16'd58007, 16'd65325, 16'd64769, 16'd43254, 16'd18899, 16'd45289});
	test_expansion(128'hc728b065eee8e678bd33c59e6159c1d2, {16'd24536, 16'd22142, 16'd2469, 16'd31648, 16'd12461, 16'd18323, 16'd31126, 16'd44722, 16'd32091, 16'd53682, 16'd45124, 16'd28051, 16'd28059, 16'd11281, 16'd7888, 16'd18639, 16'd38379, 16'd25137, 16'd64887, 16'd15074, 16'd56666, 16'd35685, 16'd42716, 16'd60665, 16'd22991, 16'd33729});
	test_expansion(128'h1043b9690b71a187a8cc55165f6109d5, {16'd46068, 16'd33207, 16'd29044, 16'd36343, 16'd15399, 16'd55041, 16'd46642, 16'd39461, 16'd10360, 16'd35511, 16'd6147, 16'd2776, 16'd52005, 16'd59161, 16'd56587, 16'd53976, 16'd61271, 16'd12647, 16'd65405, 16'd48466, 16'd49219, 16'd9593, 16'd22364, 16'd28242, 16'd56443, 16'd40530});
	test_expansion(128'he48766b3a245ba688f006d5ee5464200, {16'd38393, 16'd5770, 16'd19673, 16'd28978, 16'd11755, 16'd217, 16'd41361, 16'd833, 16'd9291, 16'd36645, 16'd14967, 16'd22457, 16'd53053, 16'd47975, 16'd50965, 16'd2411, 16'd23539, 16'd27894, 16'd46541, 16'd33175, 16'd32576, 16'd36119, 16'd51102, 16'd9258, 16'd10976, 16'd37353});
	test_expansion(128'hf5a9d273d733e1a40b7e85635a7f2180, {16'd11232, 16'd60972, 16'd3431, 16'd4301, 16'd35991, 16'd42452, 16'd11890, 16'd49150, 16'd15864, 16'd36553, 16'd22292, 16'd41209, 16'd25067, 16'd4245, 16'd11315, 16'd39530, 16'd49495, 16'd35558, 16'd28504, 16'd29753, 16'd37239, 16'd52966, 16'd2799, 16'd31677, 16'd47440, 16'd50500});
	test_expansion(128'h7f321e5523857d918846e8a6bc1968e6, {16'd36304, 16'd52452, 16'd27659, 16'd63897, 16'd65430, 16'd26946, 16'd40859, 16'd37325, 16'd1785, 16'd33444, 16'd64954, 16'd4855, 16'd63510, 16'd36098, 16'd24784, 16'd12191, 16'd31882, 16'd22205, 16'd64752, 16'd30449, 16'd18247, 16'd17335, 16'd1462, 16'd53082, 16'd46535, 16'd1089});
	test_expansion(128'hfcb250c83300e9ece336b803db632428, {16'd55871, 16'd18585, 16'd102, 16'd57660, 16'd24822, 16'd1539, 16'd45220, 16'd15337, 16'd39829, 16'd4766, 16'd20675, 16'd16701, 16'd8703, 16'd50650, 16'd64959, 16'd39827, 16'd11393, 16'd46652, 16'd8174, 16'd19284, 16'd61309, 16'd36872, 16'd33206, 16'd16000, 16'd42606, 16'd7532});
	test_expansion(128'h23cd97f85eb91d525a0bcf60e4f6b5d1, {16'd56863, 16'd45067, 16'd55431, 16'd39642, 16'd10158, 16'd24702, 16'd5247, 16'd64809, 16'd63640, 16'd13110, 16'd7901, 16'd12679, 16'd48768, 16'd59825, 16'd16411, 16'd6485, 16'd64572, 16'd354, 16'd58891, 16'd50319, 16'd42918, 16'd3156, 16'd50897, 16'd64741, 16'd32385, 16'd5427});
	test_expansion(128'h0a1d8cf6c97533546bc9a25e58a9001f, {16'd62786, 16'd58939, 16'd44972, 16'd65293, 16'd6092, 16'd55228, 16'd9470, 16'd10057, 16'd12215, 16'd51734, 16'd55442, 16'd9533, 16'd64330, 16'd12626, 16'd49968, 16'd22646, 16'd42335, 16'd30207, 16'd3272, 16'd45762, 16'd23972, 16'd54649, 16'd42014, 16'd30863, 16'd20178, 16'd51207});
	test_expansion(128'h4e4259ce925814e9e08dabb08f50074c, {16'd40333, 16'd59491, 16'd4674, 16'd30696, 16'd10069, 16'd61250, 16'd56460, 16'd38451, 16'd25308, 16'd5627, 16'd31140, 16'd26941, 16'd14988, 16'd21020, 16'd38735, 16'd21927, 16'd40106, 16'd18643, 16'd138, 16'd26978, 16'd23519, 16'd54416, 16'd21531, 16'd25279, 16'd63748, 16'd53927});
	test_expansion(128'h73d052e94aef7256fdeb52de02c43193, {16'd3171, 16'd64575, 16'd33177, 16'd16452, 16'd43094, 16'd4738, 16'd29894, 16'd62287, 16'd4127, 16'd23275, 16'd3768, 16'd40202, 16'd13172, 16'd40384, 16'd51685, 16'd48670, 16'd18986, 16'd58171, 16'd49845, 16'd15119, 16'd49071, 16'd978, 16'd61622, 16'd47121, 16'd8863, 16'd3165});
	test_expansion(128'h112d9b5e2236e87a5d334fd95a1b5248, {16'd3232, 16'd6372, 16'd12662, 16'd58534, 16'd28035, 16'd4220, 16'd40369, 16'd9834, 16'd38958, 16'd34427, 16'd43701, 16'd21559, 16'd46787, 16'd64197, 16'd55166, 16'd33209, 16'd12350, 16'd41717, 16'd53511, 16'd43546, 16'd235, 16'd21300, 16'd24766, 16'd13727, 16'd1671, 16'd61794});
	test_expansion(128'h5a72efb937c92bffd84852b034435886, {16'd14638, 16'd4153, 16'd23621, 16'd32917, 16'd11627, 16'd53158, 16'd30583, 16'd64997, 16'd13351, 16'd21818, 16'd40608, 16'd36967, 16'd2512, 16'd15460, 16'd32288, 16'd54360, 16'd4734, 16'd64313, 16'd64864, 16'd21638, 16'd47014, 16'd61234, 16'd6706, 16'd42090, 16'd20020, 16'd19939});
	test_expansion(128'hdbc97302f610b34a20411ef85f6c606b, {16'd29863, 16'd45241, 16'd22258, 16'd39381, 16'd55696, 16'd61118, 16'd47017, 16'd60906, 16'd33069, 16'd1363, 16'd27427, 16'd58689, 16'd14420, 16'd3486, 16'd57023, 16'd53969, 16'd4433, 16'd40738, 16'd2663, 16'd24388, 16'd1499, 16'd34198, 16'd65505, 16'd34138, 16'd47572, 16'd61006});
	test_expansion(128'he9002865bf8897c03e7a988e5efd4819, {16'd58328, 16'd56105, 16'd52730, 16'd53030, 16'd2760, 16'd42429, 16'd15704, 16'd33844, 16'd13928, 16'd12570, 16'd23535, 16'd10818, 16'd23255, 16'd48519, 16'd56362, 16'd13794, 16'd23761, 16'd639, 16'd57714, 16'd36518, 16'd47879, 16'd50192, 16'd30547, 16'd13206, 16'd52075, 16'd43313});
	test_expansion(128'h26595ea076427140abff1e35c74c17ec, {16'd5942, 16'd30090, 16'd52761, 16'd31628, 16'd36638, 16'd18886, 16'd25040, 16'd50419, 16'd10560, 16'd55963, 16'd32045, 16'd27820, 16'd28745, 16'd39526, 16'd43730, 16'd59095, 16'd62747, 16'd25589, 16'd48296, 16'd36551, 16'd40504, 16'd56162, 16'd29558, 16'd45360, 16'd55004, 16'd985});
	test_expansion(128'h0c4ffbc10ebac433281e19a608863dff, {16'd53147, 16'd51074, 16'd22633, 16'd783, 16'd29352, 16'd49450, 16'd46118, 16'd28321, 16'd25848, 16'd29084, 16'd40603, 16'd58137, 16'd53710, 16'd43845, 16'd12049, 16'd42059, 16'd2072, 16'd36571, 16'd64126, 16'd23571, 16'd38945, 16'd56802, 16'd60748, 16'd38779, 16'd26298, 16'd10913});
	test_expansion(128'hfc2c726f8586b91b392f522607ea936f, {16'd41698, 16'd16770, 16'd18608, 16'd45779, 16'd45750, 16'd20543, 16'd36661, 16'd21951, 16'd2903, 16'd12510, 16'd22031, 16'd7040, 16'd43234, 16'd38219, 16'd46431, 16'd19432, 16'd43420, 16'd29309, 16'd11047, 16'd64323, 16'd5305, 16'd30520, 16'd35917, 16'd50821, 16'd32577, 16'd54586});
	test_expansion(128'h6010bc36486b71835a2cdcacff993b00, {16'd19228, 16'd28832, 16'd46602, 16'd55528, 16'd44037, 16'd20717, 16'd4012, 16'd51092, 16'd48558, 16'd43672, 16'd53321, 16'd44450, 16'd26840, 16'd8996, 16'd12090, 16'd41534, 16'd65270, 16'd48522, 16'd26016, 16'd22981, 16'd49982, 16'd20004, 16'd10543, 16'd23444, 16'd46832, 16'd63245});
	test_expansion(128'h8dc0a7c305758f756e0949186a05f275, {16'd2993, 16'd44706, 16'd53062, 16'd47430, 16'd62110, 16'd8959, 16'd34110, 16'd703, 16'd34106, 16'd35792, 16'd3955, 16'd45275, 16'd14903, 16'd37810, 16'd18062, 16'd44087, 16'd1997, 16'd35703, 16'd64508, 16'd2944, 16'd11815, 16'd17911, 16'd38942, 16'd39122, 16'd46001, 16'd54475});
	test_expansion(128'he93554e9407fadb55d857b8291de881d, {16'd8291, 16'd23800, 16'd41550, 16'd50304, 16'd29732, 16'd17789, 16'd4985, 16'd12869, 16'd52248, 16'd36718, 16'd31616, 16'd32124, 16'd9688, 16'd21876, 16'd2546, 16'd23013, 16'd60824, 16'd29441, 16'd45143, 16'd25912, 16'd52943, 16'd5814, 16'd25249, 16'd59548, 16'd15274, 16'd16372});
	test_expansion(128'h4c3f150b683e10fb23791aa5cac09c0e, {16'd51253, 16'd27255, 16'd42704, 16'd18739, 16'd45338, 16'd31920, 16'd64615, 16'd47083, 16'd22699, 16'd50533, 16'd14623, 16'd33583, 16'd45085, 16'd60854, 16'd37565, 16'd61079, 16'd57600, 16'd24133, 16'd7983, 16'd36365, 16'd39280, 16'd4074, 16'd27795, 16'd16836, 16'd26999, 16'd62447});
	test_expansion(128'hf77f8093362624244c945b8a12915ae5, {16'd19273, 16'd65378, 16'd52333, 16'd59043, 16'd33919, 16'd22247, 16'd10965, 16'd62280, 16'd24882, 16'd15237, 16'd16738, 16'd413, 16'd25868, 16'd11081, 16'd63078, 16'd13205, 16'd26899, 16'd37230, 16'd24899, 16'd12428, 16'd63073, 16'd42896, 16'd50351, 16'd2611, 16'd49925, 16'd25468});
	test_expansion(128'h6f431c20503797c0b4bcd93eb8cd8868, {16'd22120, 16'd16516, 16'd57151, 16'd26150, 16'd51419, 16'd36578, 16'd25839, 16'd9617, 16'd39287, 16'd53868, 16'd37781, 16'd33805, 16'd51422, 16'd25068, 16'd691, 16'd27709, 16'd53632, 16'd34422, 16'd57418, 16'd54656, 16'd33917, 16'd61224, 16'd64828, 16'd10389, 16'd35778, 16'd50792});
	test_expansion(128'h32aa9866e3ccd60e3b08286190e056f8, {16'd30812, 16'd21393, 16'd62918, 16'd47287, 16'd7934, 16'd9373, 16'd20844, 16'd32642, 16'd51698, 16'd4024, 16'd21016, 16'd5717, 16'd58968, 16'd27203, 16'd41719, 16'd55967, 16'd13392, 16'd12148, 16'd17577, 16'd31874, 16'd27232, 16'd24539, 16'd21241, 16'd57359, 16'd18446, 16'd26049});
	test_expansion(128'hc464a666491f2d755ed82cd90e883146, {16'd11530, 16'd23308, 16'd14384, 16'd62577, 16'd32697, 16'd3601, 16'd44295, 16'd17998, 16'd36376, 16'd1618, 16'd39486, 16'd52975, 16'd44180, 16'd56542, 16'd47181, 16'd8598, 16'd60832, 16'd45966, 16'd53844, 16'd24299, 16'd19591, 16'd12445, 16'd22273, 16'd36920, 16'd61831, 16'd7575});
	test_expansion(128'h87b389e863c5b413779d1ee900fb376a, {16'd51308, 16'd26649, 16'd50997, 16'd21819, 16'd25074, 16'd3568, 16'd3894, 16'd55117, 16'd62082, 16'd64628, 16'd15391, 16'd21081, 16'd38303, 16'd54296, 16'd23880, 16'd55829, 16'd444, 16'd38343, 16'd13217, 16'd6299, 16'd58178, 16'd10262, 16'd61639, 16'd35803, 16'd48579, 16'd15639});
	test_expansion(128'h5000c36edcdad0edaf464c15607fea93, {16'd29351, 16'd21477, 16'd38772, 16'd22647, 16'd28661, 16'd50640, 16'd4783, 16'd45157, 16'd61471, 16'd20433, 16'd1707, 16'd34172, 16'd42140, 16'd40658, 16'd45457, 16'd3516, 16'd56500, 16'd64445, 16'd2435, 16'd41510, 16'd49789, 16'd43005, 16'd9002, 16'd21488, 16'd52031, 16'd7570});
	test_expansion(128'h2a02d92eaec16a5658959e7db2884fc7, {16'd31046, 16'd42950, 16'd61508, 16'd53770, 16'd63, 16'd30025, 16'd14695, 16'd47387, 16'd40208, 16'd9326, 16'd53836, 16'd58920, 16'd20046, 16'd60643, 16'd6492, 16'd52550, 16'd54862, 16'd27537, 16'd36286, 16'd28559, 16'd20157, 16'd26009, 16'd25015, 16'd45885, 16'd660, 16'd39414});
	test_expansion(128'h9cd92a8044b38e8544efb519a53e6312, {16'd16362, 16'd62738, 16'd2055, 16'd24905, 16'd32123, 16'd40890, 16'd63456, 16'd56078, 16'd42050, 16'd32608, 16'd3092, 16'd49491, 16'd8164, 16'd5160, 16'd50577, 16'd51022, 16'd62826, 16'd35372, 16'd55489, 16'd54090, 16'd3612, 16'd40404, 16'd60482, 16'd58689, 16'd39107, 16'd4396});
	test_expansion(128'h74d3216c506b99935acaaa3b7c609d69, {16'd27182, 16'd10591, 16'd22322, 16'd39960, 16'd49768, 16'd54713, 16'd27113, 16'd40087, 16'd5942, 16'd27410, 16'd39919, 16'd39696, 16'd19888, 16'd49138, 16'd33123, 16'd27794, 16'd43926, 16'd59823, 16'd14048, 16'd5678, 16'd64524, 16'd62230, 16'd44404, 16'd11967, 16'd907, 16'd16368});
	test_expansion(128'h3226968c82480e4347e0801b7b417762, {16'd13581, 16'd4179, 16'd43054, 16'd16144, 16'd55333, 16'd11853, 16'd17973, 16'd7652, 16'd18871, 16'd34012, 16'd10909, 16'd10668, 16'd41908, 16'd15604, 16'd11247, 16'd56480, 16'd61929, 16'd761, 16'd58417, 16'd59303, 16'd59766, 16'd62656, 16'd11744, 16'd28433, 16'd7342, 16'd41156});
	test_expansion(128'ha466e5c2bf950d3183ad8a44e4f7a4d7, {16'd57731, 16'd21903, 16'd40588, 16'd60941, 16'd30860, 16'd6063, 16'd28734, 16'd58266, 16'd3000, 16'd42476, 16'd20138, 16'd44474, 16'd40729, 16'd23701, 16'd23288, 16'd3954, 16'd18762, 16'd20760, 16'd50999, 16'd49141, 16'd44677, 16'd28985, 16'd39889, 16'd59864, 16'd25363, 16'd26869});
	test_expansion(128'h4ee8c8cf07739282e3a38d4e209226ee, {16'd54376, 16'd56050, 16'd55017, 16'd19328, 16'd39677, 16'd27990, 16'd22272, 16'd21720, 16'd39640, 16'd29463, 16'd15526, 16'd54919, 16'd53302, 16'd58959, 16'd50051, 16'd54059, 16'd1390, 16'd49764, 16'd3198, 16'd34056, 16'd43160, 16'd43787, 16'd39106, 16'd27160, 16'd5057, 16'd26152});
	test_expansion(128'h8d20de2deeb7b8dcaaca47ddcdd4779f, {16'd10699, 16'd32602, 16'd13842, 16'd22900, 16'd21166, 16'd12236, 16'd54806, 16'd37238, 16'd1673, 16'd7731, 16'd50237, 16'd13735, 16'd35033, 16'd15299, 16'd12178, 16'd27094, 16'd23007, 16'd58580, 16'd52557, 16'd39643, 16'd51095, 16'd46363, 16'd34956, 16'd28877, 16'd12177, 16'd42924});
	test_expansion(128'h568b3b9ee66ee29fe6da4551c53490b2, {16'd26341, 16'd34702, 16'd34657, 16'd39774, 16'd65109, 16'd21412, 16'd35406, 16'd24906, 16'd3950, 16'd49718, 16'd33868, 16'd34128, 16'd13931, 16'd34533, 16'd9214, 16'd47235, 16'd58980, 16'd44217, 16'd33898, 16'd33889, 16'd3294, 16'd48559, 16'd29947, 16'd1798, 16'd60796, 16'd45907});
	test_expansion(128'h36dd55e9da2f2c551e28dbb377ced1dd, {16'd44153, 16'd24675, 16'd17723, 16'd5543, 16'd49151, 16'd2839, 16'd53691, 16'd13916, 16'd33519, 16'd25303, 16'd8777, 16'd29709, 16'd11895, 16'd53547, 16'd64419, 16'd51122, 16'd13486, 16'd17794, 16'd5915, 16'd61606, 16'd313, 16'd28326, 16'd56564, 16'd60384, 16'd33510, 16'd28440});
	test_expansion(128'h82b525cda83f65b2697020998fa43e77, {16'd62494, 16'd59506, 16'd26522, 16'd40673, 16'd25096, 16'd13829, 16'd36356, 16'd64607, 16'd55346, 16'd17270, 16'd43665, 16'd63102, 16'd64663, 16'd6678, 16'd49671, 16'd14105, 16'd36891, 16'd58837, 16'd19922, 16'd35378, 16'd50296, 16'd50296, 16'd33698, 16'd64705, 16'd45840, 16'd14948});
	test_expansion(128'he459d7ef75e6e3d091f275f380ea8243, {16'd33061, 16'd55614, 16'd10520, 16'd2681, 16'd35308, 16'd46930, 16'd28332, 16'd59468, 16'd59158, 16'd39111, 16'd58605, 16'd28112, 16'd8039, 16'd60859, 16'd34150, 16'd37416, 16'd45648, 16'd256, 16'd10194, 16'd53735, 16'd60560, 16'd22025, 16'd806, 16'd47088, 16'd44587, 16'd22242});
	test_expansion(128'hf0edb1b52b200221262d02595afea8f2, {16'd45681, 16'd59960, 16'd23500, 16'd55722, 16'd41221, 16'd3830, 16'd11313, 16'd10009, 16'd54065, 16'd28189, 16'd22816, 16'd15653, 16'd62290, 16'd50444, 16'd53999, 16'd14612, 16'd42079, 16'd62342, 16'd34036, 16'd23660, 16'd39781, 16'd684, 16'd52315, 16'd22645, 16'd34529, 16'd34835});
	test_expansion(128'h4ac92551f8f8e2745c967c30082e3a5e, {16'd4969, 16'd11722, 16'd14034, 16'd28708, 16'd153, 16'd4199, 16'd36354, 16'd51078, 16'd27625, 16'd37913, 16'd15748, 16'd19176, 16'd57160, 16'd61158, 16'd58725, 16'd21324, 16'd2595, 16'd191, 16'd40951, 16'd42571, 16'd32698, 16'd34149, 16'd54302, 16'd46188, 16'd13281, 16'd17741});
	test_expansion(128'hbdf45d2a02724ede00f7049880b8e734, {16'd29072, 16'd47374, 16'd55425, 16'd1219, 16'd33912, 16'd29228, 16'd47679, 16'd63233, 16'd33163, 16'd14885, 16'd31370, 16'd40024, 16'd54547, 16'd23417, 16'd18826, 16'd20564, 16'd52430, 16'd36457, 16'd9061, 16'd60115, 16'd55173, 16'd64419, 16'd52661, 16'd3062, 16'd38862, 16'd25118});
	test_expansion(128'h4c7b897ad3d4a91d4ad68212ff48e93c, {16'd787, 16'd6555, 16'd62210, 16'd3921, 16'd4065, 16'd43552, 16'd51221, 16'd6845, 16'd44581, 16'd38636, 16'd42567, 16'd28235, 16'd23232, 16'd22785, 16'd4785, 16'd44631, 16'd37686, 16'd38693, 16'd25063, 16'd34345, 16'd46329, 16'd58294, 16'd38622, 16'd6219, 16'd16202, 16'd20638});
	test_expansion(128'h26646192d25d389de9b2d9a2da664997, {16'd19518, 16'd8417, 16'd18203, 16'd33723, 16'd42809, 16'd48057, 16'd17402, 16'd29568, 16'd38037, 16'd31021, 16'd54528, 16'd41631, 16'd853, 16'd27272, 16'd62, 16'd3260, 16'd1848, 16'd55124, 16'd49741, 16'd16368, 16'd35266, 16'd47718, 16'd50568, 16'd46290, 16'd29322, 16'd17663});
	test_expansion(128'h850913af0dd8bd52aa174756ff34e015, {16'd55311, 16'd10855, 16'd41570, 16'd2318, 16'd2430, 16'd17233, 16'd267, 16'd37418, 16'd35191, 16'd33587, 16'd37366, 16'd38056, 16'd53675, 16'd17870, 16'd61784, 16'd7512, 16'd20857, 16'd16572, 16'd27675, 16'd35713, 16'd16144, 16'd51289, 16'd49601, 16'd3667, 16'd1703, 16'd53907});
	test_expansion(128'h11573767e0c586204e9d191fd1ac87d6, {16'd6455, 16'd26032, 16'd54381, 16'd43225, 16'd22398, 16'd23263, 16'd20217, 16'd30060, 16'd40438, 16'd54499, 16'd50, 16'd64775, 16'd13394, 16'd55876, 16'd58078, 16'd20545, 16'd19268, 16'd50628, 16'd25163, 16'd12593, 16'd1730, 16'd50343, 16'd12527, 16'd29644, 16'd24144, 16'd29445});
	test_expansion(128'h8ee4f6b8c2dfee648d38c97bb7d76b01, {16'd32003, 16'd3231, 16'd34175, 16'd21784, 16'd46018, 16'd21936, 16'd54015, 16'd53325, 16'd37963, 16'd405, 16'd5420, 16'd29625, 16'd1943, 16'd43393, 16'd3721, 16'd58888, 16'd7524, 16'd15892, 16'd16874, 16'd63431, 16'd17805, 16'd2359, 16'd8864, 16'd51668, 16'd42059, 16'd52863});
	test_expansion(128'h1e1ee749a53750546ea09d32b5a39edd, {16'd23925, 16'd60361, 16'd4647, 16'd34846, 16'd12961, 16'd55401, 16'd44095, 16'd38627, 16'd708, 16'd57137, 16'd16160, 16'd45960, 16'd760, 16'd31526, 16'd49697, 16'd39722, 16'd33298, 16'd51219, 16'd20615, 16'd62455, 16'd15264, 16'd43044, 16'd37190, 16'd16594, 16'd32743, 16'd14152});
	test_expansion(128'h231fd44ef0aa2fd1d7d8a805089b63a7, {16'd18916, 16'd32698, 16'd29782, 16'd38474, 16'd44394, 16'd23155, 16'd549, 16'd59956, 16'd31477, 16'd27880, 16'd45592, 16'd22201, 16'd1230, 16'd23487, 16'd40205, 16'd50581, 16'd13060, 16'd6995, 16'd43483, 16'd17446, 16'd50512, 16'd26144, 16'd212, 16'd1068, 16'd33754, 16'd29751});
	test_expansion(128'h170825154cf547e55970821f8bbe69f9, {16'd31377, 16'd48467, 16'd20312, 16'd19340, 16'd47643, 16'd5117, 16'd47870, 16'd33466, 16'd56134, 16'd50115, 16'd27308, 16'd9052, 16'd46804, 16'd52129, 16'd9187, 16'd54583, 16'd33511, 16'd61684, 16'd41278, 16'd36227, 16'd27162, 16'd39963, 16'd46977, 16'd52152, 16'd30404, 16'd18556});
	test_expansion(128'h8581a0e2043e63ce4cd68c7fdd1fc590, {16'd21123, 16'd5467, 16'd27287, 16'd7928, 16'd16362, 16'd21388, 16'd38445, 16'd58521, 16'd60691, 16'd57388, 16'd34747, 16'd4817, 16'd4306, 16'd36912, 16'd22262, 16'd19389, 16'd52806, 16'd40871, 16'd33984, 16'd63208, 16'd50194, 16'd9523, 16'd26769, 16'd17159, 16'd9663, 16'd45282});
	test_expansion(128'h65a836772127e7652652b082d76d73d5, {16'd13244, 16'd6371, 16'd4532, 16'd4892, 16'd9682, 16'd29205, 16'd61567, 16'd46253, 16'd26140, 16'd24012, 16'd23774, 16'd27443, 16'd20471, 16'd20129, 16'd47439, 16'd6704, 16'd698, 16'd8085, 16'd46602, 16'd64282, 16'd33071, 16'd3919, 16'd3413, 16'd29447, 16'd372, 16'd9272});
	test_expansion(128'h6bb30dfb5e3251a8afa9b63dcad3148c, {16'd32304, 16'd7057, 16'd20793, 16'd34764, 16'd2696, 16'd51311, 16'd5601, 16'd16898, 16'd17729, 16'd32995, 16'd19374, 16'd57430, 16'd27053, 16'd57481, 16'd54429, 16'd8522, 16'd42856, 16'd49070, 16'd29279, 16'd29245, 16'd62301, 16'd44131, 16'd49386, 16'd53578, 16'd10570, 16'd24764});
	test_expansion(128'h8090a38977b5d73028938415b1eb8773, {16'd46240, 16'd47794, 16'd20122, 16'd35462, 16'd15441, 16'd3431, 16'd27917, 16'd787, 16'd34549, 16'd14033, 16'd13924, 16'd22123, 16'd4026, 16'd61098, 16'd40649, 16'd46850, 16'd15096, 16'd54649, 16'd23738, 16'd20558, 16'd40727, 16'd5702, 16'd31950, 16'd23303, 16'd55015, 16'd15187});
	test_expansion(128'h531a8dc1c3b0b1e85c7cbc144d783955, {16'd1021, 16'd46955, 16'd6784, 16'd11351, 16'd18235, 16'd18348, 16'd51938, 16'd8542, 16'd13094, 16'd27818, 16'd57060, 16'd8991, 16'd18341, 16'd6824, 16'd22545, 16'd54490, 16'd33365, 16'd39385, 16'd1601, 16'd64438, 16'd11544, 16'd2549, 16'd19319, 16'd52368, 16'd17525, 16'd57825});
	test_expansion(128'h9c1752ec707191101230a46b7a9bd302, {16'd18765, 16'd46583, 16'd60238, 16'd64550, 16'd44928, 16'd27282, 16'd25841, 16'd10008, 16'd1412, 16'd61303, 16'd37979, 16'd56040, 16'd50251, 16'd22952, 16'd47137, 16'd42918, 16'd46878, 16'd62402, 16'd38260, 16'd22544, 16'd24719, 16'd18842, 16'd41856, 16'd16261, 16'd31944, 16'd18625});
	test_expansion(128'h7a4c4e039344861b19e2a3915a4948d6, {16'd46339, 16'd25427, 16'd8333, 16'd36247, 16'd34198, 16'd39355, 16'd60279, 16'd28240, 16'd40682, 16'd33219, 16'd60869, 16'd52001, 16'd12515, 16'd8796, 16'd19483, 16'd46798, 16'd10972, 16'd42139, 16'd58960, 16'd56149, 16'd62708, 16'd53952, 16'd58513, 16'd54474, 16'd55304, 16'd42417});
	test_expansion(128'hc3e3351d4f9ace3af9c3fb4975d98a04, {16'd7059, 16'd38103, 16'd19739, 16'd14606, 16'd22747, 16'd59771, 16'd62586, 16'd65171, 16'd4655, 16'd34980, 16'd33639, 16'd10873, 16'd17495, 16'd48693, 16'd8338, 16'd10430, 16'd39265, 16'd9726, 16'd48458, 16'd31376, 16'd42316, 16'd19442, 16'd12136, 16'd28956, 16'd48798, 16'd56286});
	test_expansion(128'h453b6e194d8c517efad2b59ad4ad36f2, {16'd49488, 16'd40392, 16'd22635, 16'd3593, 16'd42821, 16'd23623, 16'd30716, 16'd633, 16'd54258, 16'd27100, 16'd24274, 16'd4383, 16'd48912, 16'd41276, 16'd39634, 16'd31497, 16'd56420, 16'd29376, 16'd37580, 16'd28471, 16'd32168, 16'd22888, 16'd29587, 16'd39179, 16'd27221, 16'd22551});
	test_expansion(128'h87a1339e44ecf90dbd920745cbc9e43d, {16'd23857, 16'd45405, 16'd18255, 16'd47780, 16'd61733, 16'd41693, 16'd30245, 16'd34780, 16'd47326, 16'd43876, 16'd54986, 16'd5050, 16'd35705, 16'd3377, 16'd7498, 16'd7971, 16'd54232, 16'd54350, 16'd36650, 16'd19528, 16'd135, 16'd6670, 16'd19530, 16'd52528, 16'd29311, 16'd33044});
	test_expansion(128'h8a62bfc3807d7efb228eba73f5a9ada5, {16'd61235, 16'd30809, 16'd4432, 16'd45412, 16'd53473, 16'd21238, 16'd44442, 16'd30354, 16'd55409, 16'd45705, 16'd55352, 16'd2387, 16'd23083, 16'd30714, 16'd19810, 16'd48360, 16'd24666, 16'd48830, 16'd40615, 16'd64145, 16'd38674, 16'd35524, 16'd48810, 16'd58864, 16'd47061, 16'd43001});
	test_expansion(128'ha61f54a03c9c3e588be92bfc14dcb024, {16'd27227, 16'd31372, 16'd13888, 16'd51425, 16'd55795, 16'd61394, 16'd8429, 16'd51503, 16'd61600, 16'd37263, 16'd15542, 16'd28851, 16'd30250, 16'd59202, 16'd48169, 16'd48320, 16'd5189, 16'd57096, 16'd38731, 16'd8681, 16'd63702, 16'd30162, 16'd6885, 16'd2900, 16'd55533, 16'd62959});
	test_expansion(128'hceab9e0fa2cca24bdfb90b5073f01df7, {16'd25850, 16'd39473, 16'd6047, 16'd4652, 16'd13566, 16'd3404, 16'd13246, 16'd28325, 16'd25325, 16'd61468, 16'd22829, 16'd22753, 16'd64890, 16'd48366, 16'd8456, 16'd43448, 16'd51979, 16'd37682, 16'd12544, 16'd44281, 16'd35613, 16'd60400, 16'd31549, 16'd35878, 16'd37714, 16'd14855});
	test_expansion(128'ha5251f4f29ddead26220a1fad9ae5444, {16'd14631, 16'd34080, 16'd49186, 16'd16968, 16'd25020, 16'd25108, 16'd39025, 16'd31328, 16'd43354, 16'd60245, 16'd16073, 16'd3987, 16'd48745, 16'd45785, 16'd34325, 16'd6721, 16'd16195, 16'd47164, 16'd57678, 16'd1331, 16'd65200, 16'd36121, 16'd2380, 16'd8052, 16'd20728, 16'd24175});
	test_expansion(128'hc6548012c6ee3627495da36f4df7e6ee, {16'd43921, 16'd23613, 16'd64619, 16'd30475, 16'd6931, 16'd61284, 16'd58840, 16'd51619, 16'd60316, 16'd64539, 16'd43739, 16'd27607, 16'd20592, 16'd1531, 16'd55059, 16'd24739, 16'd7267, 16'd28604, 16'd16525, 16'd54677, 16'd23584, 16'd21541, 16'd9263, 16'd57316, 16'd54231, 16'd58977});
	test_expansion(128'h54be4bdd68605be4fa2dc2856c501973, {16'd55944, 16'd21794, 16'd16872, 16'd26236, 16'd39995, 16'd32285, 16'd48778, 16'd34550, 16'd20791, 16'd51600, 16'd2823, 16'd7100, 16'd31907, 16'd28523, 16'd40076, 16'd46394, 16'd5078, 16'd25345, 16'd32670, 16'd23842, 16'd17854, 16'd48630, 16'd53038, 16'd46158, 16'd43085, 16'd2758});
	test_expansion(128'h5368cdb2620dee37c6ddce35ba6aaeff, {16'd42460, 16'd8679, 16'd13485, 16'd19384, 16'd54231, 16'd9150, 16'd19856, 16'd1660, 16'd25756, 16'd30005, 16'd24732, 16'd52532, 16'd16863, 16'd56576, 16'd14676, 16'd1675, 16'd46618, 16'd55050, 16'd25588, 16'd38868, 16'd63205, 16'd56654, 16'd13902, 16'd59435, 16'd10358, 16'd32610});
	test_expansion(128'h45bb9059d66e62546b6e25d2f4f0a28a, {16'd44209, 16'd3794, 16'd15309, 16'd52803, 16'd31431, 16'd50807, 16'd52302, 16'd59031, 16'd34287, 16'd15340, 16'd42554, 16'd49760, 16'd48346, 16'd27291, 16'd21273, 16'd45068, 16'd58245, 16'd21706, 16'd64450, 16'd46183, 16'd8189, 16'd33375, 16'd18893, 16'd41915, 16'd56135, 16'd33523});
	test_expansion(128'h56fa304a3e52ab0e927bba08fb7fa9e1, {16'd52246, 16'd39270, 16'd14750, 16'd42122, 16'd45129, 16'd6028, 16'd44864, 16'd53869, 16'd16611, 16'd21485, 16'd32238, 16'd55196, 16'd25751, 16'd45252, 16'd46165, 16'd56593, 16'd352, 16'd39596, 16'd56112, 16'd48214, 16'd26495, 16'd9808, 16'd52904, 16'd63082, 16'd60152, 16'd33702});
	test_expansion(128'h93664a051ea1bc2a0c3d8c5829f41738, {16'd20760, 16'd37954, 16'd46492, 16'd56599, 16'd3442, 16'd42189, 16'd32494, 16'd50104, 16'd11754, 16'd49126, 16'd59572, 16'd30832, 16'd28268, 16'd24210, 16'd7999, 16'd38537, 16'd44345, 16'd12983, 16'd7683, 16'd22837, 16'd6941, 16'd23869, 16'd3200, 16'd34610, 16'd6611, 16'd15079});
	test_expansion(128'hdf7bac3d76961df56735e73e7e934f05, {16'd36875, 16'd8245, 16'd61158, 16'd28746, 16'd44203, 16'd18407, 16'd7327, 16'd50172, 16'd45814, 16'd11304, 16'd50894, 16'd51766, 16'd42370, 16'd43185, 16'd18944, 16'd38352, 16'd53807, 16'd25979, 16'd17893, 16'd29000, 16'd52685, 16'd14754, 16'd27375, 16'd21623, 16'd54230, 16'd27238});
	test_expansion(128'h07147e2778c9191726a5a46fa016e291, {16'd32860, 16'd22053, 16'd24427, 16'd1468, 16'd28138, 16'd48719, 16'd3401, 16'd42502, 16'd43779, 16'd7997, 16'd48575, 16'd40439, 16'd48872, 16'd48519, 16'd47290, 16'd47241, 16'd44592, 16'd40772, 16'd13756, 16'd15167, 16'd17471, 16'd48976, 16'd58194, 16'd7264, 16'd7375, 16'd1537});
	test_expansion(128'hcf34f3db9e8bffa3ff17373ddc66f588, {16'd35432, 16'd45485, 16'd35115, 16'd42695, 16'd8594, 16'd58225, 16'd41823, 16'd4286, 16'd53327, 16'd58116, 16'd49600, 16'd7391, 16'd2328, 16'd9953, 16'd53319, 16'd27170, 16'd61993, 16'd44833, 16'd50644, 16'd57281, 16'd23753, 16'd1614, 16'd47559, 16'd40000, 16'd35374, 16'd18212});
	test_expansion(128'h12b618ece8c601341eded7f0d813c58d, {16'd51526, 16'd56093, 16'd45782, 16'd44239, 16'd15602, 16'd170, 16'd6353, 16'd56658, 16'd43579, 16'd55966, 16'd64047, 16'd35651, 16'd42640, 16'd756, 16'd28420, 16'd57189, 16'd39675, 16'd49034, 16'd43850, 16'd32381, 16'd34645, 16'd50898, 16'd47589, 16'd21143, 16'd24345, 16'd37514});
	test_expansion(128'hdb4712de008b7035e278b62bb72d700b, {16'd1863, 16'd50347, 16'd18228, 16'd53595, 16'd7365, 16'd51033, 16'd18474, 16'd6111, 16'd58187, 16'd21893, 16'd5874, 16'd32118, 16'd14037, 16'd26680, 16'd55033, 16'd57391, 16'd17255, 16'd26256, 16'd23283, 16'd40728, 16'd35566, 16'd5211, 16'd14244, 16'd2562, 16'd63829, 16'd53398});
	test_expansion(128'h2a24358c26099d40d4774cc9ecfe4d0a, {16'd14374, 16'd45552, 16'd25452, 16'd36504, 16'd35487, 16'd37667, 16'd52819, 16'd58252, 16'd7003, 16'd9197, 16'd13833, 16'd30362, 16'd44479, 16'd4943, 16'd3852, 16'd61954, 16'd26040, 16'd63272, 16'd40500, 16'd7307, 16'd16475, 16'd36554, 16'd50415, 16'd50157, 16'd5006, 16'd50095});
	test_expansion(128'h50080e5e7c6fffbcb0fc82e9f5036c4d, {16'd26457, 16'd51147, 16'd2487, 16'd28372, 16'd1598, 16'd21899, 16'd25023, 16'd54317, 16'd13448, 16'd59499, 16'd22771, 16'd22591, 16'd64675, 16'd43141, 16'd52117, 16'd30123, 16'd39738, 16'd26641, 16'd3200, 16'd51434, 16'd53437, 16'd61484, 16'd14119, 16'd61769, 16'd47324, 16'd312});
	test_expansion(128'hae1dfc4dc4c093b1153ac483ee96faf1, {16'd42576, 16'd41573, 16'd58866, 16'd16679, 16'd11585, 16'd15006, 16'd46736, 16'd44869, 16'd50243, 16'd62655, 16'd41558, 16'd778, 16'd47592, 16'd49077, 16'd36753, 16'd31339, 16'd30703, 16'd60863, 16'd44656, 16'd15363, 16'd54292, 16'd63335, 16'd27753, 16'd28009, 16'd35523, 16'd28995});
	test_expansion(128'ha5a708f6e7d04185c67344cec62db694, {16'd45241, 16'd30947, 16'd25689, 16'd3591, 16'd18293, 16'd579, 16'd11466, 16'd52166, 16'd13407, 16'd16398, 16'd43563, 16'd18536, 16'd41241, 16'd55012, 16'd34812, 16'd22284, 16'd21588, 16'd11980, 16'd46779, 16'd33361, 16'd42321, 16'd59280, 16'd53789, 16'd29514, 16'd23330, 16'd24687});
	test_expansion(128'h7b4376f06fd7fe3e5aa776b84b9ca3b6, {16'd10558, 16'd62829, 16'd941, 16'd65282, 16'd43271, 16'd35777, 16'd21018, 16'd11125, 16'd50803, 16'd19524, 16'd35763, 16'd32120, 16'd40661, 16'd37607, 16'd33927, 16'd40289, 16'd20783, 16'd9213, 16'd51437, 16'd22424, 16'd34415, 16'd39320, 16'd5578, 16'd18599, 16'd24527, 16'd9216});
	test_expansion(128'h625062d375e0d41ceb50c9b4c28c49ce, {16'd43060, 16'd41468, 16'd26957, 16'd16854, 16'd11197, 16'd54119, 16'd20109, 16'd41018, 16'd62657, 16'd8914, 16'd53514, 16'd27273, 16'd43753, 16'd56971, 16'd59515, 16'd39815, 16'd52587, 16'd53349, 16'd29259, 16'd33769, 16'd11882, 16'd53239, 16'd14228, 16'd6527, 16'd43596, 16'd35107});
	test_expansion(128'hd48f8236df85088956a213b4f3b6400b, {16'd3270, 16'd62580, 16'd5247, 16'd56673, 16'd30190, 16'd37071, 16'd45028, 16'd9253, 16'd48037, 16'd39884, 16'd35199, 16'd36170, 16'd22754, 16'd54685, 16'd40405, 16'd10555, 16'd27935, 16'd58823, 16'd61564, 16'd13365, 16'd36294, 16'd5969, 16'd26198, 16'd45389, 16'd2248, 16'd64686});
	test_expansion(128'hc030ec9329ac656b3180bdbc4de73f15, {16'd51165, 16'd7775, 16'd11847, 16'd25676, 16'd51747, 16'd62689, 16'd4070, 16'd5425, 16'd2861, 16'd2593, 16'd27044, 16'd62819, 16'd60686, 16'd48402, 16'd12655, 16'd1429, 16'd26407, 16'd9684, 16'd22317, 16'd9289, 16'd61238, 16'd61115, 16'd1622, 16'd44202, 16'd2411, 16'd14967});
	test_expansion(128'hc2748b85a1376a753560eb0365f05b85, {16'd60968, 16'd33116, 16'd34632, 16'd39812, 16'd26702, 16'd52829, 16'd31889, 16'd56585, 16'd30825, 16'd5891, 16'd11, 16'd52694, 16'd5362, 16'd35664, 16'd50514, 16'd32107, 16'd63212, 16'd49037, 16'd12098, 16'd50095, 16'd268, 16'd3463, 16'd44064, 16'd62021, 16'd31560, 16'd61639});
	test_expansion(128'h88f9879832e63a27cc2b7d06753e042b, {16'd18698, 16'd41972, 16'd35425, 16'd33162, 16'd17515, 16'd27187, 16'd47769, 16'd58943, 16'd65211, 16'd26820, 16'd4929, 16'd62948, 16'd34549, 16'd40046, 16'd23990, 16'd26337, 16'd22333, 16'd16824, 16'd63526, 16'd52918, 16'd16818, 16'd2197, 16'd58305, 16'd48292, 16'd50926, 16'd47452});
	test_expansion(128'ha984de47bbdac3bf4c0de3a19b031bf7, {16'd21098, 16'd53151, 16'd12636, 16'd25986, 16'd60235, 16'd5521, 16'd13948, 16'd26785, 16'd64210, 16'd56961, 16'd45925, 16'd34936, 16'd3942, 16'd58056, 16'd10279, 16'd65422, 16'd12952, 16'd23495, 16'd20522, 16'd26847, 16'd52808, 16'd58559, 16'd41724, 16'd2725, 16'd58068, 16'd5372});
	test_expansion(128'h13758b9e88dfe05cf8dd458da5cf7a4a, {16'd39409, 16'd6151, 16'd19861, 16'd49370, 16'd61166, 16'd58657, 16'd56035, 16'd25618, 16'd33769, 16'd33418, 16'd10744, 16'd4758, 16'd12905, 16'd8987, 16'd1055, 16'd9084, 16'd13828, 16'd15758, 16'd44104, 16'd48338, 16'd20424, 16'd56954, 16'd51664, 16'd43301, 16'd63230, 16'd60181});
	test_expansion(128'hc8beadf33c6c850425f887229fb5346f, {16'd38920, 16'd1948, 16'd24432, 16'd62733, 16'd34028, 16'd15681, 16'd52023, 16'd32510, 16'd52844, 16'd6637, 16'd14479, 16'd15138, 16'd8948, 16'd35904, 16'd48043, 16'd23554, 16'd7813, 16'd16182, 16'd61810, 16'd13094, 16'd32084, 16'd45698, 16'd44288, 16'd56647, 16'd37198, 16'd55031});
	test_expansion(128'h6a9c2a0c80174e28b070230121548f51, {16'd2435, 16'd64101, 16'd14723, 16'd30527, 16'd56492, 16'd43718, 16'd23136, 16'd46635, 16'd30110, 16'd55246, 16'd36745, 16'd3540, 16'd32518, 16'd521, 16'd17418, 16'd64329, 16'd21904, 16'd5460, 16'd47398, 16'd30627, 16'd63613, 16'd751, 16'd8830, 16'd41160, 16'd27194, 16'd37571});
	test_expansion(128'h541d3e62c55793fa0762b6c4c7816d93, {16'd26473, 16'd27521, 16'd17345, 16'd6774, 16'd196, 16'd17724, 16'd35402, 16'd61714, 16'd34449, 16'd12817, 16'd23737, 16'd13822, 16'd45857, 16'd14471, 16'd41008, 16'd34906, 16'd29859, 16'd24369, 16'd52657, 16'd25268, 16'd16318, 16'd40621, 16'd49390, 16'd61049, 16'd2541, 16'd52053});
	test_expansion(128'h7d9affc981baed54d8f7e3823f0bcd27, {16'd14597, 16'd23707, 16'd38376, 16'd63507, 16'd54145, 16'd15924, 16'd20017, 16'd63241, 16'd53412, 16'd53543, 16'd22672, 16'd3189, 16'd13083, 16'd63363, 16'd42683, 16'd64734, 16'd41755, 16'd26390, 16'd44775, 16'd6869, 16'd65292, 16'd58328, 16'd49339, 16'd17560, 16'd23180, 16'd51957});
	test_expansion(128'h428203cf6e7982a8a3be279e28d315b1, {16'd43590, 16'd56745, 16'd35349, 16'd32645, 16'd44920, 16'd28812, 16'd4760, 16'd12900, 16'd21764, 16'd12718, 16'd32436, 16'd3735, 16'd40681, 16'd49726, 16'd57256, 16'd52171, 16'd36353, 16'd24782, 16'd17190, 16'd35448, 16'd27693, 16'd63481, 16'd48485, 16'd51946, 16'd91, 16'd42552});
	test_expansion(128'hbe6373009b8f30aa551fe15e102ce178, {16'd10716, 16'd49769, 16'd21839, 16'd34881, 16'd7116, 16'd18408, 16'd24140, 16'd54630, 16'd32851, 16'd43223, 16'd34266, 16'd19927, 16'd59732, 16'd3669, 16'd46602, 16'd26390, 16'd11996, 16'd45324, 16'd40020, 16'd43372, 16'd43838, 16'd9174, 16'd17940, 16'd55495, 16'd16674, 16'd6878});
	test_expansion(128'h95ea92835589a13e85a2b3cf5a7b511b, {16'd54631, 16'd26810, 16'd42192, 16'd48567, 16'd65083, 16'd1784, 16'd63159, 16'd45128, 16'd15538, 16'd19771, 16'd46433, 16'd55590, 16'd3673, 16'd62937, 16'd16517, 16'd8674, 16'd1949, 16'd7010, 16'd29840, 16'd14955, 16'd51022, 16'd52149, 16'd45418, 16'd55335, 16'd23874, 16'd10438});
	test_expansion(128'h3616b1b4d440480b8f6998a173beab05, {16'd63860, 16'd40273, 16'd45114, 16'd12067, 16'd9758, 16'd17634, 16'd22274, 16'd19621, 16'd62943, 16'd24603, 16'd53821, 16'd26006, 16'd48, 16'd32245, 16'd51319, 16'd50961, 16'd48462, 16'd36030, 16'd11148, 16'd47529, 16'd51437, 16'd4826, 16'd53373, 16'd12891, 16'd32635, 16'd3917});
	test_expansion(128'h236e99c6d05452b898c3a619e384d166, {16'd1802, 16'd33451, 16'd63498, 16'd32565, 16'd12759, 16'd24328, 16'd23602, 16'd12466, 16'd5837, 16'd24507, 16'd46168, 16'd27659, 16'd23173, 16'd33220, 16'd3434, 16'd35479, 16'd44222, 16'd39851, 16'd18362, 16'd61649, 16'd16579, 16'd64020, 16'd43969, 16'd10590, 16'd53132, 16'd2284});
	test_expansion(128'h85505cc4713ff20835872b67d8fc048b, {16'd31630, 16'd23254, 16'd62880, 16'd21025, 16'd56159, 16'd32741, 16'd19545, 16'd22956, 16'd13263, 16'd5534, 16'd9142, 16'd37352, 16'd37967, 16'd30278, 16'd5582, 16'd44209, 16'd7521, 16'd39834, 16'd51231, 16'd59771, 16'd55045, 16'd64297, 16'd25149, 16'd5276, 16'd53715, 16'd9424});
	test_expansion(128'h648febac6ff7cb12be8f2ccd8be76d28, {16'd21887, 16'd12691, 16'd21320, 16'd65468, 16'd52942, 16'd58651, 16'd23595, 16'd41597, 16'd52739, 16'd10410, 16'd62765, 16'd63865, 16'd43579, 16'd15795, 16'd44600, 16'd8351, 16'd1446, 16'd21438, 16'd37822, 16'd30782, 16'd41480, 16'd43326, 16'd3463, 16'd56908, 16'd24929, 16'd22709});
	test_expansion(128'hd1e7859a5776fe54a3bde1337bae6005, {16'd63888, 16'd7250, 16'd24684, 16'd22566, 16'd57442, 16'd31757, 16'd38836, 16'd50648, 16'd30897, 16'd29232, 16'd51926, 16'd42930, 16'd25889, 16'd4818, 16'd35016, 16'd31020, 16'd50965, 16'd37060, 16'd60221, 16'd25767, 16'd25582, 16'd57288, 16'd58636, 16'd47843, 16'd37961, 16'd31429});
	test_expansion(128'hedf261adc25276f36e59ac159ea84906, {16'd19755, 16'd267, 16'd52062, 16'd23190, 16'd23850, 16'd40509, 16'd55380, 16'd37440, 16'd61453, 16'd409, 16'd49446, 16'd37593, 16'd20341, 16'd48920, 16'd45302, 16'd51457, 16'd64065, 16'd7297, 16'd21676, 16'd1067, 16'd21527, 16'd57595, 16'd43689, 16'd34942, 16'd43575, 16'd49516});
	test_expansion(128'h77445c45eb4013a8cd9a78eb8aa5af86, {16'd3568, 16'd32838, 16'd64226, 16'd47489, 16'd64190, 16'd57446, 16'd63618, 16'd58148, 16'd10131, 16'd339, 16'd12839, 16'd29197, 16'd7684, 16'd14343, 16'd62778, 16'd50671, 16'd31399, 16'd30073, 16'd11020, 16'd2768, 16'd56182, 16'd57322, 16'd44081, 16'd61382, 16'd41155, 16'd18184});
	test_expansion(128'hfe64fc92fb07bd2ecd29eedeb816ab8d, {16'd4165, 16'd61039, 16'd54726, 16'd17856, 16'd13473, 16'd6865, 16'd64541, 16'd59227, 16'd59457, 16'd29316, 16'd53520, 16'd39114, 16'd10587, 16'd48628, 16'd4062, 16'd4550, 16'd33742, 16'd7590, 16'd49064, 16'd41114, 16'd44077, 16'd51451, 16'd4967, 16'd45559, 16'd49367, 16'd55653});
	test_expansion(128'hf9c1275de56a1140c7b7603f624cd619, {16'd46352, 16'd13874, 16'd32921, 16'd58888, 16'd60856, 16'd2501, 16'd17904, 16'd16525, 16'd52334, 16'd58979, 16'd29856, 16'd62255, 16'd18272, 16'd23025, 16'd32206, 16'd40295, 16'd63899, 16'd44311, 16'd64118, 16'd43705, 16'd6922, 16'd8404, 16'd6341, 16'd10440, 16'd38049, 16'd901});
	test_expansion(128'hed9c2f35f30929c01a82446b6b70299b, {16'd35864, 16'd13558, 16'd1876, 16'd10311, 16'd11228, 16'd18214, 16'd16092, 16'd43541, 16'd57156, 16'd9913, 16'd22555, 16'd2101, 16'd61474, 16'd34371, 16'd62161, 16'd57445, 16'd59492, 16'd21646, 16'd57152, 16'd18717, 16'd52436, 16'd7766, 16'd56876, 16'd64963, 16'd38366, 16'd26670});
	test_expansion(128'h9f2dbc7e8bc6e64209b345fc20efe978, {16'd18099, 16'd23645, 16'd49237, 16'd27022, 16'd50218, 16'd7517, 16'd52114, 16'd23651, 16'd53861, 16'd7214, 16'd19987, 16'd17530, 16'd32774, 16'd33, 16'd29535, 16'd44228, 16'd17986, 16'd39020, 16'd58389, 16'd30648, 16'd20475, 16'd58472, 16'd53687, 16'd2388, 16'd60458, 16'd22491});
	test_expansion(128'h3facec2d032f33cbc19c27180ecb4cac, {16'd34845, 16'd18905, 16'd57175, 16'd4241, 16'd37248, 16'd63548, 16'd20088, 16'd33445, 16'd44507, 16'd14459, 16'd10090, 16'd26979, 16'd57892, 16'd31609, 16'd42154, 16'd8131, 16'd58167, 16'd21507, 16'd23855, 16'd11141, 16'd40548, 16'd29280, 16'd52566, 16'd53923, 16'd55703, 16'd21596});
	test_expansion(128'h2c3777dc99512d9bf0a825afc569c748, {16'd6074, 16'd37118, 16'd28864, 16'd31882, 16'd53915, 16'd35863, 16'd55353, 16'd24909, 16'd48502, 16'd61933, 16'd29371, 16'd9776, 16'd11572, 16'd48989, 16'd20738, 16'd46291, 16'd23995, 16'd42754, 16'd24245, 16'd48511, 16'd15883, 16'd45674, 16'd60238, 16'd40987, 16'd9669, 16'd157});
	test_expansion(128'h132f946fd7da1eff74f36b07eb5cf3d1, {16'd6095, 16'd27441, 16'd31402, 16'd31483, 16'd30034, 16'd42262, 16'd19015, 16'd53987, 16'd58982, 16'd939, 16'd27987, 16'd61882, 16'd49854, 16'd50334, 16'd63236, 16'd20176, 16'd47290, 16'd19347, 16'd8484, 16'd20324, 16'd63986, 16'd12667, 16'd58446, 16'd25080, 16'd48894, 16'd10108});
	test_expansion(128'h98aab7a3983226f55e0a260524386706, {16'd9781, 16'd62785, 16'd23072, 16'd13675, 16'd9890, 16'd13202, 16'd21650, 16'd46553, 16'd6196, 16'd36616, 16'd2500, 16'd14606, 16'd16450, 16'd21170, 16'd7577, 16'd24736, 16'd58947, 16'd65288, 16'd19196, 16'd11170, 16'd14037, 16'd64296, 16'd44455, 16'd43495, 16'd9208, 16'd2921});
	test_expansion(128'h5f77b74d26627abf5ccada1d00f8ee26, {16'd52793, 16'd64196, 16'd36164, 16'd43054, 16'd24499, 16'd51389, 16'd41707, 16'd11425, 16'd50847, 16'd35898, 16'd23545, 16'd64952, 16'd32149, 16'd21545, 16'd17923, 16'd36736, 16'd53784, 16'd15699, 16'd33106, 16'd21270, 16'd54082, 16'd13159, 16'd13209, 16'd15665, 16'd51559, 16'd52770});
	test_expansion(128'hbb2b88b151c1f9383e8b9bb7bb021d88, {16'd65041, 16'd50376, 16'd11065, 16'd55378, 16'd3446, 16'd43555, 16'd10149, 16'd31142, 16'd60702, 16'd4453, 16'd43375, 16'd10400, 16'd57645, 16'd4243, 16'd10612, 16'd16431, 16'd27131, 16'd51504, 16'd24617, 16'd19477, 16'd5023, 16'd54455, 16'd58142, 16'd58585, 16'd64307, 16'd37074});
	test_expansion(128'hba63d1d1ac4e892790b163745ece73be, {16'd34505, 16'd62417, 16'd60212, 16'd28303, 16'd55392, 16'd37362, 16'd33152, 16'd40624, 16'd21733, 16'd38050, 16'd29101, 16'd11330, 16'd40914, 16'd61440, 16'd50831, 16'd4251, 16'd37516, 16'd60879, 16'd47648, 16'd45996, 16'd18955, 16'd29713, 16'd42949, 16'd56350, 16'd61529, 16'd23218});
	test_expansion(128'h2c45c6f5e43ec88a7f3cedf29255b10e, {16'd56560, 16'd55374, 16'd39189, 16'd49802, 16'd55242, 16'd27000, 16'd22529, 16'd30478, 16'd62206, 16'd55454, 16'd47589, 16'd29812, 16'd35393, 16'd49465, 16'd44309, 16'd62581, 16'd27101, 16'd35039, 16'd33977, 16'd64735, 16'd38079, 16'd61433, 16'd49898, 16'd56816, 16'd16099, 16'd62511});
	test_expansion(128'hacb02dd9dd1b661c1d9a663d67b9df82, {16'd12170, 16'd29514, 16'd23762, 16'd12314, 16'd41072, 16'd59443, 16'd11689, 16'd7940, 16'd29897, 16'd27337, 16'd12856, 16'd29015, 16'd23192, 16'd40966, 16'd31742, 16'd42187, 16'd42448, 16'd23165, 16'd63225, 16'd4657, 16'd35474, 16'd27140, 16'd42645, 16'd52797, 16'd28456, 16'd24609});
	test_expansion(128'hb2c31dc23f97a017decb7c2b9cdab58c, {16'd13134, 16'd36509, 16'd40927, 16'd10916, 16'd58075, 16'd25971, 16'd6547, 16'd14062, 16'd48596, 16'd32173, 16'd49087, 16'd25780, 16'd44010, 16'd52930, 16'd35115, 16'd37858, 16'd5123, 16'd56214, 16'd18980, 16'd15505, 16'd24409, 16'd30755, 16'd1150, 16'd641, 16'd47702, 16'd55745});
	test_expansion(128'h6779823a0649b8e79c1d9a696a440b4a, {16'd36824, 16'd47782, 16'd14922, 16'd32977, 16'd2871, 16'd7038, 16'd19675, 16'd44100, 16'd56791, 16'd31394, 16'd11911, 16'd36747, 16'd43552, 16'd42669, 16'd51382, 16'd43828, 16'd21089, 16'd11587, 16'd10335, 16'd35767, 16'd21239, 16'd64171, 16'd39822, 16'd15451, 16'd1146, 16'd4563});
	test_expansion(128'he6adca4e54609f295943f3f82782ef09, {16'd39068, 16'd31817, 16'd49052, 16'd15138, 16'd26810, 16'd895, 16'd36731, 16'd29473, 16'd57756, 16'd38624, 16'd16694, 16'd42918, 16'd47279, 16'd64256, 16'd38297, 16'd61277, 16'd65505, 16'd11451, 16'd50682, 16'd16167, 16'd44634, 16'd38869, 16'd24651, 16'd62971, 16'd136, 16'd58931});
	test_expansion(128'ha0952a832aaff681a28417a0ababd1ab, {16'd13245, 16'd62513, 16'd34554, 16'd63481, 16'd2276, 16'd48232, 16'd11826, 16'd15070, 16'd64132, 16'd46225, 16'd51320, 16'd58242, 16'd23623, 16'd43297, 16'd33875, 16'd55847, 16'd15764, 16'd25273, 16'd22534, 16'd37103, 16'd28740, 16'd29225, 16'd53209, 16'd23424, 16'd63198, 16'd612});
	test_expansion(128'h19735c0d8de43c59f0ebee0d536d8617, {16'd41150, 16'd32305, 16'd3705, 16'd37192, 16'd34036, 16'd22853, 16'd18109, 16'd19582, 16'd47795, 16'd46521, 16'd14544, 16'd6098, 16'd18318, 16'd6170, 16'd26595, 16'd32496, 16'd17068, 16'd2324, 16'd32336, 16'd55329, 16'd26056, 16'd2101, 16'd45570, 16'd31693, 16'd63925, 16'd5842});
	test_expansion(128'h8918c56836dc5c0f980200c4921f1e0e, {16'd7972, 16'd15866, 16'd16638, 16'd4010, 16'd46476, 16'd1642, 16'd24101, 16'd49209, 16'd63648, 16'd45477, 16'd2646, 16'd17000, 16'd27337, 16'd10085, 16'd60032, 16'd47452, 16'd23125, 16'd62944, 16'd60395, 16'd52350, 16'd33946, 16'd52243, 16'd29585, 16'd61924, 16'd4537, 16'd9485});
	test_expansion(128'h53e43cdea6c96a3fb46cb65402df7b20, {16'd23041, 16'd28367, 16'd6205, 16'd4315, 16'd36891, 16'd19617, 16'd2655, 16'd36506, 16'd17110, 16'd5197, 16'd10654, 16'd23660, 16'd33292, 16'd6989, 16'd8954, 16'd40037, 16'd42353, 16'd62872, 16'd35913, 16'd63079, 16'd27840, 16'd55803, 16'd7606, 16'd51306, 16'd20664, 16'd64435});
	test_expansion(128'h628c750f7c380d898b10ba53f0b359cd, {16'd38294, 16'd29290, 16'd30148, 16'd19614, 16'd35234, 16'd43458, 16'd52137, 16'd9688, 16'd2394, 16'd16703, 16'd36647, 16'd19050, 16'd10334, 16'd30637, 16'd57360, 16'd21580, 16'd34255, 16'd33588, 16'd25218, 16'd2154, 16'd56706, 16'd8657, 16'd41240, 16'd60840, 16'd17406, 16'd7067});
	test_expansion(128'ha5ee2a91401ae36a98f1a2cdfac5cde1, {16'd30431, 16'd28597, 16'd61484, 16'd26076, 16'd15849, 16'd29014, 16'd60120, 16'd57020, 16'd41087, 16'd7824, 16'd31637, 16'd46306, 16'd10120, 16'd33186, 16'd1684, 16'd35916, 16'd19918, 16'd60499, 16'd53581, 16'd64919, 16'd25774, 16'd233, 16'd29118, 16'd64050, 16'd47164, 16'd11428});
	test_expansion(128'h196cfe8571e2b9ead1c52889066f4d11, {16'd60171, 16'd48244, 16'd16856, 16'd41904, 16'd25173, 16'd13878, 16'd355, 16'd17477, 16'd4045, 16'd27902, 16'd55278, 16'd45542, 16'd1697, 16'd38105, 16'd3793, 16'd53495, 16'd45975, 16'd13654, 16'd1503, 16'd35080, 16'd36328, 16'd5819, 16'd38184, 16'd13460, 16'd13556, 16'd1122});
	test_expansion(128'hea11d821edad6040e7f060cb918b4b9e, {16'd55291, 16'd38022, 16'd7095, 16'd19559, 16'd11150, 16'd4947, 16'd52406, 16'd60203, 16'd45015, 16'd36997, 16'd28760, 16'd5013, 16'd3257, 16'd3675, 16'd30296, 16'd29098, 16'd49468, 16'd38378, 16'd60141, 16'd26537, 16'd40532, 16'd48978, 16'd5138, 16'd49467, 16'd62689, 16'd64907});
	test_expansion(128'h75caecb5c3110242714a5f5eed75a6ab, {16'd32426, 16'd50502, 16'd36664, 16'd187, 16'd42813, 16'd39, 16'd56869, 16'd9872, 16'd12078, 16'd30698, 16'd38792, 16'd54781, 16'd17593, 16'd41075, 16'd29736, 16'd18969, 16'd57952, 16'd18608, 16'd61319, 16'd441, 16'd17669, 16'd35017, 16'd56583, 16'd18919, 16'd55143, 16'd39747});
	test_expansion(128'h645b395ad9022ebef13d7644d470d10b, {16'd2441, 16'd3961, 16'd17957, 16'd3660, 16'd38832, 16'd18288, 16'd20771, 16'd45500, 16'd32361, 16'd14245, 16'd15528, 16'd12588, 16'd24772, 16'd55158, 16'd15276, 16'd64203, 16'd26120, 16'd48600, 16'd53983, 16'd27078, 16'd34359, 16'd29443, 16'd44851, 16'd4536, 16'd8949, 16'd37485});
	test_expansion(128'he1acae5784f90c96dea89c9080c33e0f, {16'd3798, 16'd14330, 16'd21946, 16'd12369, 16'd33180, 16'd45149, 16'd32592, 16'd47619, 16'd57240, 16'd31482, 16'd44278, 16'd45518, 16'd5281, 16'd53865, 16'd65058, 16'd54672, 16'd64844, 16'd23646, 16'd54033, 16'd12008, 16'd23906, 16'd36732, 16'd13332, 16'd23588, 16'd13469, 16'd20966});
	test_expansion(128'h6805979b5365e5c1322dccead9d93565, {16'd14515, 16'd40653, 16'd52654, 16'd1734, 16'd17137, 16'd48668, 16'd26841, 16'd34415, 16'd46071, 16'd56095, 16'd17779, 16'd40444, 16'd12331, 16'd34665, 16'd37540, 16'd17363, 16'd1800, 16'd32515, 16'd35519, 16'd6568, 16'd56928, 16'd11654, 16'd13310, 16'd8591, 16'd3503, 16'd48253});
	test_expansion(128'h6629896b6309aac642c1292f275da188, {16'd25604, 16'd44478, 16'd30249, 16'd5122, 16'd28246, 16'd54479, 16'd1347, 16'd37206, 16'd32685, 16'd10551, 16'd13896, 16'd43725, 16'd63061, 16'd30453, 16'd23569, 16'd46038, 16'd51086, 16'd40379, 16'd2668, 16'd11024, 16'd9079, 16'd16150, 16'd4004, 16'd49793, 16'd27734, 16'd31826});
	test_expansion(128'h325b9cf917b7a8db8082b717ca0ce99b, {16'd8629, 16'd22609, 16'd44558, 16'd58794, 16'd36369, 16'd50868, 16'd64133, 16'd15876, 16'd21082, 16'd29461, 16'd14906, 16'd27906, 16'd15170, 16'd46437, 16'd8599, 16'd20753, 16'd5023, 16'd34826, 16'd64734, 16'd50218, 16'd26499, 16'd44591, 16'd45350, 16'd37222, 16'd25066, 16'd57935});
	test_expansion(128'h8da843a863986ece90d57c8a01aa8282, {16'd1360, 16'd41292, 16'd13415, 16'd28638, 16'd5683, 16'd50687, 16'd44610, 16'd47167, 16'd38752, 16'd63541, 16'd39966, 16'd35127, 16'd59009, 16'd36577, 16'd4547, 16'd64397, 16'd48814, 16'd3711, 16'd1373, 16'd17700, 16'd3868, 16'd60874, 16'd20688, 16'd22979, 16'd58414, 16'd21035});
	test_expansion(128'h5cbcabf52d87f0d6c135ec3978ec7fc9, {16'd60410, 16'd8981, 16'd45899, 16'd3494, 16'd5921, 16'd948, 16'd12964, 16'd43690, 16'd27357, 16'd16440, 16'd14572, 16'd8279, 16'd21212, 16'd23394, 16'd2519, 16'd29873, 16'd56345, 16'd30438, 16'd54633, 16'd50907, 16'd5574, 16'd18760, 16'd40997, 16'd15530, 16'd9380, 16'd48239});
	test_expansion(128'h64a81ebc3016d1510f3189682200ddba, {16'd16722, 16'd57685, 16'd22248, 16'd61691, 16'd8388, 16'd37066, 16'd22171, 16'd35222, 16'd16998, 16'd8616, 16'd28750, 16'd53739, 16'd19299, 16'd51229, 16'd60433, 16'd54679, 16'd703, 16'd59290, 16'd18865, 16'd36833, 16'd22188, 16'd4512, 16'd23581, 16'd29431, 16'd15725, 16'd16958});
	test_expansion(128'h3a14b52f506e5462cd6fbdeaebeae05e, {16'd23468, 16'd18146, 16'd6423, 16'd32740, 16'd11630, 16'd28324, 16'd55415, 16'd14479, 16'd43626, 16'd55238, 16'd5366, 16'd49722, 16'd8528, 16'd14819, 16'd21395, 16'd56626, 16'd40483, 16'd61131, 16'd53130, 16'd19020, 16'd49607, 16'd7441, 16'd19513, 16'd43365, 16'd20836, 16'd11757});
	test_expansion(128'hf07be10658dbe7ce60adedb1241ed17b, {16'd1446, 16'd46064, 16'd50340, 16'd26451, 16'd32683, 16'd2931, 16'd8569, 16'd49419, 16'd61850, 16'd44472, 16'd49384, 16'd36678, 16'd33255, 16'd43109, 16'd13076, 16'd22937, 16'd61941, 16'd58362, 16'd3051, 16'd23561, 16'd46308, 16'd33591, 16'd47042, 16'd59961, 16'd55343, 16'd54611});
	test_expansion(128'h61b491c83c8e33c76456906dc6e5f681, {16'd51124, 16'd55865, 16'd20948, 16'd37731, 16'd31137, 16'd57857, 16'd7685, 16'd57610, 16'd32428, 16'd57174, 16'd17708, 16'd31003, 16'd4086, 16'd2304, 16'd58806, 16'd62235, 16'd38603, 16'd37616, 16'd14166, 16'd16814, 16'd5622, 16'd51929, 16'd28839, 16'd7810, 16'd33175, 16'd46260});
	test_expansion(128'h63604dcf46d9998ca75e2b453a8c3928, {16'd59126, 16'd42785, 16'd45770, 16'd23543, 16'd27090, 16'd42776, 16'd56914, 16'd61731, 16'd37129, 16'd57382, 16'd11780, 16'd54443, 16'd3112, 16'd28912, 16'd55084, 16'd39660, 16'd16077, 16'd20607, 16'd10561, 16'd9464, 16'd3035, 16'd32575, 16'd20990, 16'd38441, 16'd53905, 16'd39707});
	test_expansion(128'he7d2d6f8b482b752c7f0c2d72fe103a3, {16'd12618, 16'd35101, 16'd35363, 16'd12828, 16'd17036, 16'd36171, 16'd9558, 16'd50825, 16'd11988, 16'd54521, 16'd61212, 16'd12790, 16'd51949, 16'd32901, 16'd26484, 16'd25790, 16'd10059, 16'd13351, 16'd10288, 16'd38277, 16'd41985, 16'd49624, 16'd9740, 16'd51457, 16'd34742, 16'd41782});
	test_expansion(128'h05c20ca3646704e238d17326a0f5aaec, {16'd22351, 16'd44726, 16'd28613, 16'd36865, 16'd51371, 16'd41372, 16'd9136, 16'd15715, 16'd31156, 16'd34488, 16'd30513, 16'd26621, 16'd9600, 16'd26644, 16'd40100, 16'd16474, 16'd13760, 16'd15907, 16'd17244, 16'd49886, 16'd17734, 16'd57795, 16'd25167, 16'd730, 16'd13866, 16'd14729});
	test_expansion(128'h81ad1a0344c0b111ff61dfc7bc2dcc25, {16'd36131, 16'd47014, 16'd32468, 16'd28230, 16'd13101, 16'd15057, 16'd38708, 16'd16634, 16'd55108, 16'd47853, 16'd41298, 16'd50209, 16'd2700, 16'd28154, 16'd39953, 16'd56245, 16'd16889, 16'd60303, 16'd9785, 16'd43995, 16'd49443, 16'd3230, 16'd43010, 16'd44970, 16'd19534, 16'd23615});
	test_expansion(128'h3e08d17ee57ff9e6589db4e245a3f6d8, {16'd15434, 16'd12857, 16'd55968, 16'd21293, 16'd29942, 16'd49390, 16'd4357, 16'd44349, 16'd16284, 16'd2177, 16'd35070, 16'd4736, 16'd54771, 16'd53171, 16'd49874, 16'd61184, 16'd8985, 16'd60096, 16'd53803, 16'd24831, 16'd65179, 16'd21947, 16'd6551, 16'd42755, 16'd35225, 16'd7274});
	test_expansion(128'h0095ab0c92822054c120741d923126f9, {16'd42318, 16'd63314, 16'd64665, 16'd47228, 16'd30076, 16'd2112, 16'd25807, 16'd62915, 16'd56570, 16'd61009, 16'd39348, 16'd6673, 16'd39821, 16'd35153, 16'd5233, 16'd49358, 16'd1021, 16'd55996, 16'd8827, 16'd37287, 16'd16285, 16'd51411, 16'd5461, 16'd18498, 16'd52571, 16'd39366});
	test_expansion(128'h0c215237161966d9cb884b3ec6e96403, {16'd63801, 16'd27896, 16'd54351, 16'd45167, 16'd10281, 16'd65387, 16'd64101, 16'd18372, 16'd62014, 16'd26337, 16'd5029, 16'd39112, 16'd34397, 16'd38051, 16'd64025, 16'd14110, 16'd50990, 16'd14394, 16'd44398, 16'd53243, 16'd21938, 16'd801, 16'd36202, 16'd49210, 16'd63203, 16'd65306});
	test_expansion(128'h59b452141ee06a6cd968eb302a23cc30, {16'd21347, 16'd33779, 16'd6854, 16'd23982, 16'd49688, 16'd1144, 16'd62060, 16'd42365, 16'd60891, 16'd47793, 16'd55075, 16'd48094, 16'd2098, 16'd10058, 16'd5515, 16'd48999, 16'd60374, 16'd25764, 16'd39355, 16'd65083, 16'd10652, 16'd22890, 16'd28367, 16'd35640, 16'd31711, 16'd43435});
	test_expansion(128'h1a9676351b6b74f7a039181293d9c66a, {16'd34167, 16'd41995, 16'd5988, 16'd10506, 16'd48779, 16'd47637, 16'd15916, 16'd19699, 16'd35827, 16'd40605, 16'd49001, 16'd45837, 16'd32620, 16'd13658, 16'd40378, 16'd2383, 16'd10539, 16'd7815, 16'd28387, 16'd32757, 16'd44398, 16'd44312, 16'd63983, 16'd43143, 16'd64693, 16'd60173});
	test_expansion(128'h2fa748b88d8ca9ae2592385a5610e2dc, {16'd64145, 16'd42353, 16'd12110, 16'd19588, 16'd941, 16'd57052, 16'd10689, 16'd53792, 16'd10288, 16'd24359, 16'd10488, 16'd64144, 16'd40931, 16'd39545, 16'd38073, 16'd13542, 16'd31822, 16'd48430, 16'd49503, 16'd50378, 16'd23842, 16'd43506, 16'd52073, 16'd25646, 16'd55986, 16'd26888});
	test_expansion(128'h9c45976844f2c2aa48fb37193d2d7738, {16'd41371, 16'd30231, 16'd4955, 16'd36672, 16'd30031, 16'd26733, 16'd20486, 16'd52819, 16'd56866, 16'd15841, 16'd50720, 16'd12884, 16'd11666, 16'd39795, 16'd28933, 16'd44202, 16'd17487, 16'd30077, 16'd12539, 16'd293, 16'd45988, 16'd14564, 16'd47471, 16'd25910, 16'd29188, 16'd55075});
	test_expansion(128'heccf54bf7a6e384efd7593f4fac7faf4, {16'd4811, 16'd32071, 16'd57175, 16'd19013, 16'd57764, 16'd9084, 16'd22161, 16'd58258, 16'd20189, 16'd17034, 16'd7336, 16'd60147, 16'd14473, 16'd41535, 16'd36, 16'd4238, 16'd62902, 16'd16973, 16'd51144, 16'd56340, 16'd61193, 16'd20411, 16'd46183, 16'd14819, 16'd16623, 16'd39060});
	test_expansion(128'ha51e070bda2e389442f4e7af7bf46873, {16'd9014, 16'd8805, 16'd46094, 16'd27457, 16'd8597, 16'd42078, 16'd24535, 16'd12149, 16'd59621, 16'd9101, 16'd44351, 16'd26963, 16'd31469, 16'd31626, 16'd14267, 16'd53656, 16'd8262, 16'd45787, 16'd55371, 16'd45269, 16'd20908, 16'd60672, 16'd63152, 16'd9164, 16'd9183, 16'd53688});
	test_expansion(128'h4239f3b17fa8221c716f8f550cc4c549, {16'd37252, 16'd62979, 16'd8288, 16'd13906, 16'd32910, 16'd42390, 16'd11289, 16'd34463, 16'd29638, 16'd51668, 16'd2248, 16'd37795, 16'd58409, 16'd7503, 16'd6678, 16'd35414, 16'd34735, 16'd56363, 16'd38683, 16'd58542, 16'd34456, 16'd61686, 16'd23001, 16'd46824, 16'd43003, 16'd46962});
	test_expansion(128'ha34a519e212fb85ffd2673e0ec4a99e5, {16'd60588, 16'd48316, 16'd44210, 16'd54798, 16'd35036, 16'd19250, 16'd47089, 16'd60692, 16'd41582, 16'd48000, 16'd42839, 16'd42359, 16'd23205, 16'd57726, 16'd23125, 16'd38325, 16'd49812, 16'd34233, 16'd45427, 16'd22013, 16'd25336, 16'd24071, 16'd27695, 16'd56924, 16'd9514, 16'd14489});
	test_expansion(128'hddc17405cb19b3524c2f7965606c8e50, {16'd63964, 16'd6850, 16'd10956, 16'd34898, 16'd15330, 16'd50432, 16'd40159, 16'd54522, 16'd13274, 16'd7315, 16'd50206, 16'd56190, 16'd46015, 16'd19574, 16'd3315, 16'd52849, 16'd54494, 16'd54219, 16'd7846, 16'd54733, 16'd44896, 16'd32040, 16'd63678, 16'd2505, 16'd64902, 16'd10014});
	test_expansion(128'h59097b73b76e081c9ac5ecde00c8e2fb, {16'd42181, 16'd44856, 16'd43082, 16'd27083, 16'd6584, 16'd19174, 16'd31569, 16'd55917, 16'd31238, 16'd20607, 16'd78, 16'd10479, 16'd38422, 16'd20030, 16'd43877, 16'd13865, 16'd60820, 16'd52844, 16'd41646, 16'd28258, 16'd52623, 16'd19140, 16'd32195, 16'd42766, 16'd8898, 16'd41260});
	test_expansion(128'h644af47b661784bffe95f88cd8971471, {16'd49551, 16'd34257, 16'd31275, 16'd27340, 16'd3387, 16'd47960, 16'd63162, 16'd5830, 16'd50589, 16'd44669, 16'd52941, 16'd26212, 16'd19208, 16'd45263, 16'd21736, 16'd64789, 16'd62680, 16'd47744, 16'd44576, 16'd29269, 16'd3334, 16'd45971, 16'd57228, 16'd48729, 16'd58574, 16'd38262});
	test_expansion(128'he1f6b43f175dc2bb646b1b18dee90708, {16'd49652, 16'd13143, 16'd57110, 16'd22700, 16'd35777, 16'd62583, 16'd8797, 16'd17560, 16'd10570, 16'd14045, 16'd62105, 16'd52852, 16'd58960, 16'd10483, 16'd24559, 16'd38481, 16'd6273, 16'd6322, 16'd13179, 16'd61229, 16'd43833, 16'd60526, 16'd62013, 16'd63527, 16'd39192, 16'd22446});
	test_expansion(128'hc12005fb5732865d1350c5ceb70b224b, {16'd41960, 16'd40535, 16'd42419, 16'd37833, 16'd36709, 16'd18806, 16'd32461, 16'd43996, 16'd6487, 16'd54470, 16'd9181, 16'd51284, 16'd30823, 16'd6169, 16'd34271, 16'd42281, 16'd22245, 16'd4522, 16'd60440, 16'd22556, 16'd19344, 16'd50274, 16'd45581, 16'd16797, 16'd5495, 16'd51441});
	test_expansion(128'h4ce68ce0ce0141dbc3b2b12a17e38833, {16'd7911, 16'd34706, 16'd18972, 16'd55940, 16'd12627, 16'd38653, 16'd60897, 16'd52160, 16'd29502, 16'd36470, 16'd32097, 16'd22797, 16'd4455, 16'd48995, 16'd48685, 16'd45266, 16'd19037, 16'd10384, 16'd22598, 16'd35529, 16'd47681, 16'd11095, 16'd3077, 16'd59774, 16'd32500, 16'd51085});
	test_expansion(128'h6ebee7793a19ca096569c55f28896704, {16'd6765, 16'd2216, 16'd40667, 16'd9258, 16'd46782, 16'd43468, 16'd5964, 16'd28310, 16'd5826, 16'd27379, 16'd41383, 16'd64445, 16'd47327, 16'd46237, 16'd10269, 16'd22756, 16'd24395, 16'd11505, 16'd36989, 16'd8596, 16'd39994, 16'd39256, 16'd11374, 16'd58935, 16'd58236, 16'd36});
	test_expansion(128'h7c9755380aae084cd62288799d233cb2, {16'd13484, 16'd48743, 16'd41596, 16'd38143, 16'd19110, 16'd27867, 16'd19580, 16'd15328, 16'd61294, 16'd23289, 16'd31156, 16'd19493, 16'd27303, 16'd24518, 16'd39633, 16'd6200, 16'd50775, 16'd57769, 16'd1547, 16'd50134, 16'd59911, 16'd25877, 16'd17547, 16'd48168, 16'd41800, 16'd48291});
	test_expansion(128'h88e6c77653d306a7f0aa4e35ea6619ef, {16'd12850, 16'd33751, 16'd23596, 16'd12332, 16'd25482, 16'd6326, 16'd7077, 16'd19872, 16'd26743, 16'd52106, 16'd50490, 16'd23814, 16'd41767, 16'd31347, 16'd64142, 16'd13857, 16'd4471, 16'd3169, 16'd60603, 16'd6855, 16'd9475, 16'd2675, 16'd26191, 16'd26214, 16'd52026, 16'd4050});
	test_expansion(128'h449fe09987f8c44f6bdcd2420bf9a545, {16'd59883, 16'd52627, 16'd24814, 16'd60419, 16'd10092, 16'd59839, 16'd19610, 16'd6549, 16'd43039, 16'd57866, 16'd53737, 16'd5946, 16'd32029, 16'd35309, 16'd30910, 16'd45814, 16'd23750, 16'd26116, 16'd61766, 16'd12940, 16'd8183, 16'd49360, 16'd41906, 16'd15389, 16'd16460, 16'd8847});
	test_expansion(128'h485f3b066b01e11003a72f548d849d75, {16'd501, 16'd2066, 16'd12026, 16'd53050, 16'd43460, 16'd21195, 16'd45103, 16'd3137, 16'd38611, 16'd44458, 16'd7345, 16'd30515, 16'd47391, 16'd23382, 16'd28865, 16'd4059, 16'd19505, 16'd7677, 16'd30884, 16'd18521, 16'd36992, 16'd41617, 16'd39479, 16'd598, 16'd6999, 16'd30569});
	test_expansion(128'h31c2114493d7d38e80e49bd61ca5590e, {16'd15268, 16'd22229, 16'd8758, 16'd34020, 16'd57188, 16'd7044, 16'd36027, 16'd57725, 16'd23580, 16'd18406, 16'd10368, 16'd32598, 16'd59437, 16'd34192, 16'd45253, 16'd19953, 16'd46470, 16'd23320, 16'd45069, 16'd59137, 16'd45656, 16'd12391, 16'd29210, 16'd35445, 16'd6567, 16'd64574});
	test_expansion(128'h95d9631b1d728a683edd0bb5cfdfdc59, {16'd51472, 16'd13138, 16'd33339, 16'd57225, 16'd41776, 16'd20890, 16'd59881, 16'd44416, 16'd11663, 16'd49501, 16'd44564, 16'd23007, 16'd61765, 16'd34088, 16'd54739, 16'd46544, 16'd4472, 16'd59095, 16'd25447, 16'd19997, 16'd53167, 16'd7061, 16'd15986, 16'd32616, 16'd2817, 16'd14900});
	test_expansion(128'h4c952967017d2629cee039ffa2be9b9b, {16'd10008, 16'd43260, 16'd29966, 16'd41690, 16'd11225, 16'd28962, 16'd60583, 16'd1601, 16'd17839, 16'd17437, 16'd1574, 16'd5799, 16'd1458, 16'd45216, 16'd11486, 16'd42782, 16'd19485, 16'd36716, 16'd50836, 16'd13478, 16'd35763, 16'd26402, 16'd1483, 16'd52818, 16'd64140, 16'd27589});
	test_expansion(128'h7a24dd397564e712d3820d09643c8244, {16'd17434, 16'd28166, 16'd8307, 16'd22620, 16'd64428, 16'd42036, 16'd13345, 16'd2803, 16'd53188, 16'd37170, 16'd40828, 16'd15785, 16'd5048, 16'd22674, 16'd60431, 16'd36669, 16'd43253, 16'd17555, 16'd34370, 16'd17271, 16'd62936, 16'd22356, 16'd63241, 16'd27167, 16'd37571, 16'd14237});
	test_expansion(128'h0403b0a77784ae4e579d1434f2ad3087, {16'd39263, 16'd25388, 16'd65520, 16'd1068, 16'd50417, 16'd54121, 16'd55247, 16'd56457, 16'd10673, 16'd58129, 16'd11036, 16'd64437, 16'd47041, 16'd32991, 16'd35088, 16'd57465, 16'd28596, 16'd27791, 16'd52137, 16'd62028, 16'd22286, 16'd8575, 16'd57486, 16'd32305, 16'd55060, 16'd17590});
	test_expansion(128'hf22d74aedc617fa49c748409d5d4211e, {16'd385, 16'd4944, 16'd33482, 16'd32034, 16'd35987, 16'd35450, 16'd31903, 16'd16657, 16'd8096, 16'd49096, 16'd8845, 16'd42598, 16'd10601, 16'd9370, 16'd24601, 16'd51040, 16'd25634, 16'd24587, 16'd8140, 16'd21168, 16'd26414, 16'd31335, 16'd12721, 16'd18985, 16'd9027, 16'd20697});
	test_expansion(128'h2778cd514477823f6fb4019921f5db29, {16'd55458, 16'd32533, 16'd10846, 16'd11349, 16'd48123, 16'd59443, 16'd43476, 16'd49247, 16'd1293, 16'd9447, 16'd13317, 16'd40736, 16'd2471, 16'd30944, 16'd49137, 16'd57113, 16'd34312, 16'd30560, 16'd41164, 16'd51738, 16'd31583, 16'd4154, 16'd14330, 16'd43331, 16'd26126, 16'd22872});
	test_expansion(128'h441daab4cfb3ab560f3c7da37a686d14, {16'd54320, 16'd51578, 16'd19842, 16'd37176, 16'd3205, 16'd44380, 16'd44475, 16'd19302, 16'd57996, 16'd16162, 16'd60154, 16'd32911, 16'd18530, 16'd11565, 16'd18637, 16'd11695, 16'd10251, 16'd7144, 16'd40301, 16'd32490, 16'd58189, 16'd46149, 16'd63012, 16'd63895, 16'd36690, 16'd51489});
	test_expansion(128'h96a2f7015804443e468b272f76b7e712, {16'd60465, 16'd53598, 16'd50199, 16'd22612, 16'd64426, 16'd15039, 16'd22787, 16'd35860, 16'd55520, 16'd63594, 16'd61760, 16'd40605, 16'd16397, 16'd28472, 16'd36594, 16'd56512, 16'd13149, 16'd15995, 16'd11327, 16'd764, 16'd18782, 16'd61804, 16'd51023, 16'd63060, 16'd15240, 16'd64499});
	test_expansion(128'h9e2f39e010d8545acd9bfd73d9a7c66e, {16'd44296, 16'd62310, 16'd8659, 16'd39341, 16'd38956, 16'd11852, 16'd56593, 16'd53622, 16'd49020, 16'd63497, 16'd34523, 16'd18083, 16'd63574, 16'd63250, 16'd46097, 16'd2305, 16'd973, 16'd64419, 16'd33508, 16'd2987, 16'd54112, 16'd5414, 16'd65378, 16'd42932, 16'd12600, 16'd33608});
	test_expansion(128'h643d4afd9fc32a8bb755efb425aa4f18, {16'd45876, 16'd22232, 16'd7236, 16'd15299, 16'd25409, 16'd7907, 16'd5152, 16'd24820, 16'd18370, 16'd38402, 16'd12934, 16'd57671, 16'd20271, 16'd36269, 16'd51468, 16'd23962, 16'd26881, 16'd14118, 16'd3774, 16'd25555, 16'd14873, 16'd18135, 16'd18212, 16'd51426, 16'd13454, 16'd46301});
	test_expansion(128'h48973791bc7827b79e394fa4afcfa259, {16'd4719, 16'd48192, 16'd47523, 16'd7497, 16'd27952, 16'd64685, 16'd13365, 16'd50338, 16'd21963, 16'd32592, 16'd15665, 16'd37588, 16'd30500, 16'd7326, 16'd14599, 16'd44560, 16'd57981, 16'd41492, 16'd41988, 16'd44883, 16'd1806, 16'd47498, 16'd56095, 16'd39113, 16'd49398, 16'd9523});
	test_expansion(128'hd50c21c106f557c2467a886e5d2bd306, {16'd37689, 16'd12989, 16'd49076, 16'd36167, 16'd25078, 16'd38851, 16'd57259, 16'd53106, 16'd33372, 16'd55663, 16'd27286, 16'd36369, 16'd11664, 16'd48881, 16'd24829, 16'd31148, 16'd42949, 16'd30656, 16'd24852, 16'd37176, 16'd61964, 16'd61820, 16'd60521, 16'd17048, 16'd22005, 16'd51538});
	test_expansion(128'h16cc92a669fe737d25eb0dc79c7cdb4b, {16'd19293, 16'd35431, 16'd28093, 16'd22721, 16'd58166, 16'd49362, 16'd4451, 16'd5954, 16'd25626, 16'd29468, 16'd40458, 16'd17892, 16'd34984, 16'd39683, 16'd22594, 16'd26769, 16'd14085, 16'd42261, 16'd63274, 16'd57025, 16'd26044, 16'd58093, 16'd14984, 16'd31823, 16'd5633, 16'd16738});
	test_expansion(128'h914c3bb00a258c49474ec84baa5feb52, {16'd32453, 16'd57950, 16'd22813, 16'd47667, 16'd53387, 16'd680, 16'd65444, 16'd34721, 16'd46810, 16'd26994, 16'd25016, 16'd46497, 16'd61877, 16'd26762, 16'd44738, 16'd23998, 16'd56356, 16'd12057, 16'd3441, 16'd57275, 16'd17896, 16'd52635, 16'd24327, 16'd62420, 16'd34165, 16'd17387});
	test_expansion(128'h3f531ddc6c131af3f2a47875deef083d, {16'd36447, 16'd42953, 16'd30659, 16'd49675, 16'd44002, 16'd47593, 16'd10675, 16'd8047, 16'd14801, 16'd22971, 16'd55914, 16'd41758, 16'd16259, 16'd55158, 16'd21757, 16'd35516, 16'd54082, 16'd61232, 16'd24759, 16'd65432, 16'd18657, 16'd19484, 16'd32494, 16'd25774, 16'd61044, 16'd11591});
	test_expansion(128'h0a970b3b91aafee8e97c11a49505fe62, {16'd11616, 16'd63180, 16'd30989, 16'd58544, 16'd37498, 16'd20899, 16'd61600, 16'd51336, 16'd53973, 16'd6330, 16'd5108, 16'd63428, 16'd46044, 16'd64677, 16'd45661, 16'd6293, 16'd3473, 16'd15503, 16'd38848, 16'd50597, 16'd20792, 16'd6856, 16'd4501, 16'd15707, 16'd22406, 16'd33617});
	test_expansion(128'hd280704bb7f8e17f31952c60ca66a574, {16'd29030, 16'd25001, 16'd32544, 16'd52420, 16'd56314, 16'd25072, 16'd12003, 16'd59839, 16'd46714, 16'd3100, 16'd17326, 16'd50709, 16'd14115, 16'd42669, 16'd2628, 16'd26736, 16'd1551, 16'd5393, 16'd6284, 16'd614, 16'd39771, 16'd60472, 16'd15846, 16'd7891, 16'd32633, 16'd21346});
	test_expansion(128'h0e68a19b3237df3bd2e421cf37461267, {16'd52556, 16'd10093, 16'd9037, 16'd55487, 16'd34454, 16'd3727, 16'd9501, 16'd58696, 16'd64835, 16'd36168, 16'd485, 16'd45109, 16'd1492, 16'd26561, 16'd18191, 16'd26848, 16'd46343, 16'd51059, 16'd64252, 16'd52119, 16'd30295, 16'd38591, 16'd7916, 16'd64936, 16'd48173, 16'd46043});
	test_expansion(128'h07905dbc80e18dcf404991c2c1183201, {16'd17441, 16'd22847, 16'd5211, 16'd60641, 16'd19534, 16'd19251, 16'd26907, 16'd55709, 16'd23484, 16'd40809, 16'd13490, 16'd65197, 16'd5082, 16'd10093, 16'd16453, 16'd46096, 16'd21756, 16'd1228, 16'd54118, 16'd50445, 16'd41240, 16'd37705, 16'd11394, 16'd6405, 16'd26578, 16'd12424});
	test_expansion(128'he970ef5fc48be9b946e048b91bf6442c, {16'd908, 16'd63453, 16'd59253, 16'd14368, 16'd31314, 16'd523, 16'd44193, 16'd50684, 16'd21723, 16'd6639, 16'd50712, 16'd13870, 16'd59064, 16'd52324, 16'd56559, 16'd61145, 16'd14810, 16'd1535, 16'd54500, 16'd58486, 16'd22875, 16'd20212, 16'd41854, 16'd29556, 16'd55510, 16'd6609});
	test_expansion(128'h0fadf4dab96027710f16e04aeb7bb44a, {16'd45749, 16'd26804, 16'd11059, 16'd52757, 16'd2197, 16'd45086, 16'd30931, 16'd28072, 16'd63201, 16'd8471, 16'd2994, 16'd900, 16'd28020, 16'd45885, 16'd6435, 16'd47923, 16'd8564, 16'd32442, 16'd45109, 16'd54794, 16'd20296, 16'd50926, 16'd46473, 16'd47252, 16'd40470, 16'd2951});
	test_expansion(128'h7d05334229e0a53dee00738198471a76, {16'd45555, 16'd62224, 16'd20782, 16'd24088, 16'd4517, 16'd45390, 16'd52944, 16'd11600, 16'd17676, 16'd30677, 16'd31741, 16'd41673, 16'd38149, 16'd7998, 16'd21273, 16'd13449, 16'd63038, 16'd23445, 16'd43252, 16'd36540, 16'd2309, 16'd35839, 16'd38610, 16'd29825, 16'd54650, 16'd40878});
	test_expansion(128'hb397ae5ea37d92fa97097a91a212ba76, {16'd3559, 16'd38369, 16'd31883, 16'd38221, 16'd32413, 16'd40781, 16'd11852, 16'd28769, 16'd63298, 16'd28039, 16'd54451, 16'd24690, 16'd63382, 16'd34997, 16'd7467, 16'd4526, 16'd50479, 16'd12060, 16'd14898, 16'd11136, 16'd58159, 16'd39002, 16'd60457, 16'd5875, 16'd55419, 16'd4});
	test_expansion(128'h88fbd8d2158619e37e480537ad5d5655, {16'd33960, 16'd10279, 16'd41908, 16'd17311, 16'd43636, 16'd17787, 16'd10767, 16'd1327, 16'd9806, 16'd52180, 16'd15571, 16'd53068, 16'd40136, 16'd62648, 16'd46908, 16'd21025, 16'd64323, 16'd3432, 16'd20981, 16'd57103, 16'd58480, 16'd64917, 16'd34587, 16'd50225, 16'd47280, 16'd29920});
	test_expansion(128'h19c562342fa9dafb546f97fc56e0cd36, {16'd28159, 16'd49135, 16'd51275, 16'd53571, 16'd8828, 16'd37504, 16'd43102, 16'd65289, 16'd36720, 16'd15728, 16'd14663, 16'd25927, 16'd20428, 16'd64, 16'd27953, 16'd13465, 16'd29750, 16'd56543, 16'd6131, 16'd49756, 16'd50934, 16'd16736, 16'd63219, 16'd28695, 16'd18491, 16'd31980});
	test_expansion(128'hc99296839d7bb5dd9082c2cea5be341e, {16'd53385, 16'd26497, 16'd50197, 16'd27733, 16'd24419, 16'd41718, 16'd11012, 16'd63296, 16'd49438, 16'd25273, 16'd21354, 16'd33195, 16'd6501, 16'd36053, 16'd62150, 16'd22916, 16'd25233, 16'd59937, 16'd60301, 16'd21342, 16'd28722, 16'd29653, 16'd23566, 16'd31819, 16'd37707, 16'd30441});
	test_expansion(128'hd7af8340eb91031a1eab6cf1419f9b51, {16'd4120, 16'd33579, 16'd7100, 16'd60927, 16'd16374, 16'd32803, 16'd7864, 16'd57612, 16'd31958, 16'd49694, 16'd20179, 16'd28729, 16'd11048, 16'd8481, 16'd18716, 16'd15515, 16'd38908, 16'd38837, 16'd51908, 16'd45095, 16'd6371, 16'd15027, 16'd24576, 16'd16208, 16'd22069, 16'd62534});
	test_expansion(128'hf924bb9f0fe0d362b6513a0196f18b6b, {16'd36403, 16'd31901, 16'd40007, 16'd65014, 16'd11975, 16'd33916, 16'd35206, 16'd22440, 16'd20903, 16'd14519, 16'd10516, 16'd46334, 16'd21484, 16'd31855, 16'd24952, 16'd31077, 16'd21019, 16'd31514, 16'd44640, 16'd9991, 16'd16859, 16'd46419, 16'd42677, 16'd53042, 16'd48399, 16'd59694});
	test_expansion(128'h97b13f6914b0bf6fe899c6514dc227e7, {16'd34374, 16'd34520, 16'd40098, 16'd25809, 16'd44743, 16'd23258, 16'd31491, 16'd37725, 16'd52037, 16'd11290, 16'd61605, 16'd53384, 16'd38247, 16'd33919, 16'd57827, 16'd37116, 16'd56246, 16'd20840, 16'd53085, 16'd11938, 16'd18949, 16'd53063, 16'd13942, 16'd41805, 16'd52873, 16'd41722});
	test_expansion(128'h58a7a55ad6b83b309ca0b76704684eea, {16'd7032, 16'd27569, 16'd7306, 16'd46835, 16'd29285, 16'd35487, 16'd36166, 16'd4995, 16'd50208, 16'd63535, 16'd51947, 16'd18762, 16'd53710, 16'd35319, 16'd14232, 16'd1223, 16'd61345, 16'd4981, 16'd16620, 16'd16837, 16'd29304, 16'd50687, 16'd21730, 16'd2899, 16'd50442, 16'd65465});
	test_expansion(128'h8ed9ab1e768483e7bd294d8c845bba90, {16'd30564, 16'd13323, 16'd58481, 16'd64482, 16'd37313, 16'd7752, 16'd53378, 16'd60143, 16'd24209, 16'd2055, 16'd52777, 16'd1611, 16'd14428, 16'd38930, 16'd287, 16'd16981, 16'd11052, 16'd60841, 16'd35398, 16'd31456, 16'd22526, 16'd1191, 16'd59920, 16'd61954, 16'd12529, 16'd29844});
	test_expansion(128'h8fdfbb81d23b96c08d94c09389d597f6, {16'd62808, 16'd24737, 16'd44339, 16'd33837, 16'd15478, 16'd19563, 16'd32606, 16'd37479, 16'd48444, 16'd17884, 16'd24812, 16'd41133, 16'd36243, 16'd45785, 16'd6349, 16'd23102, 16'd33974, 16'd61149, 16'd48517, 16'd44282, 16'd43165, 16'd32344, 16'd60181, 16'd27497, 16'd20352, 16'd22496});
	test_expansion(128'h03ca898e61ea98c803bda66827940f20, {16'd38078, 16'd35636, 16'd7265, 16'd33743, 16'd3692, 16'd60361, 16'd29183, 16'd59435, 16'd20491, 16'd14842, 16'd40731, 16'd14920, 16'd64473, 16'd10195, 16'd27414, 16'd50423, 16'd24953, 16'd16117, 16'd29929, 16'd33178, 16'd9661, 16'd17334, 16'd57507, 16'd52258, 16'd37006, 16'd61524});
	test_expansion(128'hdb2f225e047fbf4c6fdf8194f35c41e5, {16'd23656, 16'd47817, 16'd55284, 16'd54388, 16'd50733, 16'd9679, 16'd44103, 16'd23649, 16'd53476, 16'd64518, 16'd55436, 16'd33208, 16'd55456, 16'd39822, 16'd31240, 16'd40829, 16'd50715, 16'd42473, 16'd42450, 16'd7813, 16'd15763, 16'd15605, 16'd62149, 16'd7550, 16'd37271, 16'd56980});
	test_expansion(128'he2ec5c9556d335bc5b4fde379a4fef50, {16'd62121, 16'd7849, 16'd45296, 16'd51795, 16'd43467, 16'd12822, 16'd5179, 16'd57528, 16'd36115, 16'd19817, 16'd26688, 16'd37304, 16'd6654, 16'd54998, 16'd12020, 16'd35493, 16'd52849, 16'd14096, 16'd10278, 16'd6119, 16'd46694, 16'd53499, 16'd61756, 16'd47956, 16'd28432, 16'd54260});
	test_expansion(128'h9e948ceb92435a8d3aa3ac91a07b294e, {16'd5344, 16'd5439, 16'd57544, 16'd9831, 16'd38495, 16'd11780, 16'd47618, 16'd5201, 16'd48299, 16'd842, 16'd19441, 16'd52793, 16'd22060, 16'd21047, 16'd56153, 16'd63386, 16'd28542, 16'd35998, 16'd17775, 16'd8127, 16'd52614, 16'd55708, 16'd31098, 16'd64910, 16'd27842, 16'd11286});
	test_expansion(128'h5bfd78a28fb5baa32173a5eee7b0a5b0, {16'd10568, 16'd46899, 16'd52769, 16'd40487, 16'd59914, 16'd25498, 16'd48294, 16'd41875, 16'd52401, 16'd35890, 16'd57316, 16'd58947, 16'd16752, 16'd48570, 16'd58837, 16'd21229, 16'd15766, 16'd27064, 16'd3700, 16'd53963, 16'd10138, 16'd62271, 16'd50594, 16'd2196, 16'd22016, 16'd32899});
	test_expansion(128'h5ac3e7dce3973ca5257a026df705a40a, {16'd60516, 16'd30217, 16'd8570, 16'd10997, 16'd64842, 16'd15980, 16'd23985, 16'd2399, 16'd58347, 16'd27026, 16'd37028, 16'd9202, 16'd63109, 16'd472, 16'd10210, 16'd10020, 16'd35225, 16'd20415, 16'd26800, 16'd18566, 16'd53940, 16'd59884, 16'd37958, 16'd31953, 16'd63098, 16'd18695});
	test_expansion(128'h865f042755ece73b87c0a1b964e9af82, {16'd679, 16'd424, 16'd18969, 16'd9652, 16'd29792, 16'd38207, 16'd9885, 16'd7792, 16'd12189, 16'd51249, 16'd27377, 16'd28785, 16'd49518, 16'd48429, 16'd54236, 16'd50169, 16'd18560, 16'd3193, 16'd25368, 16'd17127, 16'd26294, 16'd55136, 16'd48837, 16'd40287, 16'd7512, 16'd52517});
	test_expansion(128'hd5db5eceb018befd831efaeb3971c7fe, {16'd10832, 16'd60098, 16'd62671, 16'd44566, 16'd35799, 16'd50684, 16'd56527, 16'd31944, 16'd2462, 16'd7489, 16'd4734, 16'd45978, 16'd28055, 16'd10564, 16'd40426, 16'd21522, 16'd19330, 16'd6530, 16'd49612, 16'd55539, 16'd10001, 16'd1297, 16'd15783, 16'd11522, 16'd10714, 16'd23638});
	test_expansion(128'h9ca79556f63c42691212c20f17565802, {16'd32, 16'd8788, 16'd13968, 16'd60514, 16'd46205, 16'd18678, 16'd17186, 16'd47626, 16'd51508, 16'd7737, 16'd60715, 16'd17232, 16'd36319, 16'd47253, 16'd43023, 16'd51614, 16'd42529, 16'd64484, 16'd37429, 16'd48122, 16'd20164, 16'd21473, 16'd41422, 16'd19495, 16'd736, 16'd55596});
	test_expansion(128'h21689e84a7122b4f31a203e5edfa3b34, {16'd12770, 16'd24761, 16'd12385, 16'd28976, 16'd16816, 16'd30104, 16'd22580, 16'd15695, 16'd25599, 16'd27001, 16'd12236, 16'd28452, 16'd7648, 16'd3945, 16'd59777, 16'd13898, 16'd10582, 16'd23089, 16'd28795, 16'd46962, 16'd61529, 16'd24075, 16'd13220, 16'd42827, 16'd7953, 16'd25115});
	test_expansion(128'h6c60ab7d0cb28ed5f204155edab9ac3e, {16'd25084, 16'd21127, 16'd62457, 16'd43130, 16'd51242, 16'd57751, 16'd45523, 16'd9305, 16'd23656, 16'd60895, 16'd25573, 16'd54597, 16'd52610, 16'd56022, 16'd10904, 16'd304, 16'd43163, 16'd54601, 16'd53365, 16'd4498, 16'd60609, 16'd10322, 16'd1049, 16'd29757, 16'd28795, 16'd37060});
	test_expansion(128'h50356b82911216abfd76487cd273f438, {16'd63913, 16'd8816, 16'd27693, 16'd19891, 16'd14270, 16'd57469, 16'd42355, 16'd25165, 16'd46960, 16'd30500, 16'd64160, 16'd28731, 16'd58370, 16'd23140, 16'd51869, 16'd64801, 16'd6656, 16'd32813, 16'd24598, 16'd49923, 16'd1557, 16'd48527, 16'd9998, 16'd56245, 16'd7524, 16'd44041});
	test_expansion(128'hff1d0a897b512a2c9d23deb535e7c2d1, {16'd35218, 16'd51104, 16'd31527, 16'd54560, 16'd37282, 16'd52768, 16'd6968, 16'd41089, 16'd3124, 16'd63212, 16'd31637, 16'd3054, 16'd32425, 16'd40, 16'd2268, 16'd58719, 16'd31908, 16'd7646, 16'd48684, 16'd35930, 16'd41209, 16'd263, 16'd15514, 16'd25332, 16'd56472, 16'd49173});
	test_expansion(128'he2732ba75881c198c3d1f16bf73b372d, {16'd17458, 16'd24728, 16'd60661, 16'd9917, 16'd65154, 16'd49557, 16'd20171, 16'd36660, 16'd28301, 16'd10307, 16'd5828, 16'd4795, 16'd29289, 16'd64983, 16'd36033, 16'd63161, 16'd17834, 16'd54957, 16'd24139, 16'd35067, 16'd50413, 16'd59912, 16'd34694, 16'd41097, 16'd21037, 16'd23155});
	test_expansion(128'h0172fee5fc0a0292a84c8649df8f39d7, {16'd18064, 16'd13483, 16'd42906, 16'd54711, 16'd22272, 16'd52080, 16'd57268, 16'd46289, 16'd29317, 16'd48893, 16'd49618, 16'd26645, 16'd16342, 16'd25360, 16'd7182, 16'd15645, 16'd9821, 16'd45983, 16'd4355, 16'd60943, 16'd58819, 16'd10158, 16'd18008, 16'd49387, 16'd419, 16'd44471});
	test_expansion(128'h1929dca882e604843d1e9a2ccee18db0, {16'd49610, 16'd4098, 16'd5635, 16'd24248, 16'd61911, 16'd15120, 16'd37762, 16'd18199, 16'd60606, 16'd13150, 16'd56846, 16'd15329, 16'd52680, 16'd11364, 16'd28992, 16'd37331, 16'd15707, 16'd59257, 16'd23570, 16'd1420, 16'd3210, 16'd53034, 16'd46730, 16'd40198, 16'd19861, 16'd31885});
	test_expansion(128'hf1cf9001c4c9e66308efa2b774acff89, {16'd19376, 16'd58044, 16'd46973, 16'd35366, 16'd6588, 16'd33656, 16'd455, 16'd16618, 16'd14357, 16'd12789, 16'd14618, 16'd40063, 16'd49439, 16'd59942, 16'd26741, 16'd37453, 16'd31242, 16'd18847, 16'd31691, 16'd17076, 16'd30553, 16'd9717, 16'd30901, 16'd55971, 16'd34572, 16'd5258});
	test_expansion(128'h6cea44999d3c30c05cad74c6aa04b1ce, {16'd20330, 16'd10157, 16'd32905, 16'd16563, 16'd59336, 16'd8539, 16'd48183, 16'd8895, 16'd11793, 16'd57219, 16'd3223, 16'd32372, 16'd32086, 16'd35460, 16'd15264, 16'd7343, 16'd3952, 16'd53548, 16'd58608, 16'd55298, 16'd54546, 16'd47429, 16'd12808, 16'd43947, 16'd60817, 16'd34477});
	test_expansion(128'hd2c30120867d5f7506ffbbe3b89edb18, {16'd52626, 16'd23163, 16'd36379, 16'd15170, 16'd22402, 16'd43931, 16'd5311, 16'd34740, 16'd18213, 16'd58537, 16'd43194, 16'd41020, 16'd26981, 16'd27613, 16'd47715, 16'd15118, 16'd17106, 16'd31614, 16'd9074, 16'd53898, 16'd14324, 16'd6897, 16'd65110, 16'd2303, 16'd10016, 16'd20455});
	test_expansion(128'he3b97fea46b8f21ebf46b1b3c0a913bb, {16'd37742, 16'd9000, 16'd193, 16'd15367, 16'd17517, 16'd46371, 16'd19525, 16'd40720, 16'd45892, 16'd29159, 16'd24053, 16'd56789, 16'd50880, 16'd30589, 16'd15240, 16'd11439, 16'd28826, 16'd5787, 16'd52539, 16'd35651, 16'd749, 16'd194, 16'd45284, 16'd41485, 16'd27886, 16'd23967});
	test_expansion(128'h07fc338dc14f7b499fcca7115b7f7413, {16'd25334, 16'd21964, 16'd20189, 16'd11743, 16'd27096, 16'd60979, 16'd46700, 16'd9389, 16'd47127, 16'd42755, 16'd20163, 16'd46173, 16'd59360, 16'd17249, 16'd46282, 16'd25527, 16'd54607, 16'd43346, 16'd47347, 16'd6529, 16'd50572, 16'd4426, 16'd17377, 16'd12022, 16'd12385, 16'd31280});
	test_expansion(128'h60de7945317e42d1ffe7a2c45189069f, {16'd21673, 16'd20302, 16'd24189, 16'd58549, 16'd28917, 16'd39385, 16'd36450, 16'd39404, 16'd4639, 16'd5295, 16'd63914, 16'd65116, 16'd31795, 16'd48300, 16'd41121, 16'd42493, 16'd31124, 16'd63311, 16'd40259, 16'd51141, 16'd24425, 16'd6438, 16'd60995, 16'd27159, 16'd41188, 16'd45148});
	test_expansion(128'hb5a92011bf8b37916d28100fd912f612, {16'd33894, 16'd3463, 16'd862, 16'd45875, 16'd26073, 16'd6587, 16'd57348, 16'd31431, 16'd1287, 16'd2557, 16'd41204, 16'd26414, 16'd10005, 16'd8563, 16'd49934, 16'd60511, 16'd14760, 16'd9870, 16'd10043, 16'd54876, 16'd1262, 16'd23880, 16'd28492, 16'd53475, 16'd48617, 16'd24835});
	test_expansion(128'h6f5fe97053accaf2ddddaf0ba80256d0, {16'd30173, 16'd47423, 16'd38955, 16'd2589, 16'd16212, 16'd39084, 16'd7584, 16'd19642, 16'd9154, 16'd3139, 16'd20456, 16'd65410, 16'd27414, 16'd34385, 16'd5392, 16'd5571, 16'd40993, 16'd22520, 16'd55150, 16'd27155, 16'd50914, 16'd21208, 16'd24142, 16'd27413, 16'd21378, 16'd48239});
	test_expansion(128'h2206a0a6ee8ab9a11165709640b6db5b, {16'd53427, 16'd25456, 16'd48819, 16'd45202, 16'd27244, 16'd49368, 16'd31901, 16'd10877, 16'd53245, 16'd27778, 16'd39168, 16'd23772, 16'd5118, 16'd32634, 16'd46778, 16'd17877, 16'd38079, 16'd53104, 16'd3944, 16'd53145, 16'd47630, 16'd2818, 16'd54259, 16'd19983, 16'd61706, 16'd29833});
	test_expansion(128'ha254665383c6a58ebbe1e2feffd3a317, {16'd574, 16'd6073, 16'd61987, 16'd56694, 16'd14877, 16'd9310, 16'd54745, 16'd1525, 16'd60458, 16'd46918, 16'd23014, 16'd42895, 16'd35898, 16'd4443, 16'd30298, 16'd4959, 16'd58293, 16'd59600, 16'd19565, 16'd42678, 16'd29694, 16'd13773, 16'd61646, 16'd32702, 16'd49550, 16'd54172});
	test_expansion(128'hd7f7ce395f6d58dff5cfc86d73ceca2c, {16'd65384, 16'd46429, 16'd40280, 16'd10587, 16'd38992, 16'd13960, 16'd25996, 16'd35835, 16'd22149, 16'd29512, 16'd1510, 16'd34955, 16'd43816, 16'd3775, 16'd56131, 16'd39881, 16'd29150, 16'd8744, 16'd6987, 16'd40492, 16'd16255, 16'd45384, 16'd53354, 16'd34412, 16'd20120, 16'd48512});
	test_expansion(128'hcd5f79fb5b31114a6fb4524193be67d8, {16'd11636, 16'd55351, 16'd11557, 16'd15930, 16'd4138, 16'd46548, 16'd47920, 16'd11923, 16'd46603, 16'd10008, 16'd48982, 16'd55032, 16'd64953, 16'd53257, 16'd54022, 16'd38587, 16'd42383, 16'd51236, 16'd32119, 16'd4634, 16'd22441, 16'd44819, 16'd43142, 16'd22836, 16'd65002, 16'd42726});
	test_expansion(128'hc840f1d1f915251c9ed72d20f096c8d1, {16'd18581, 16'd10505, 16'd48513, 16'd31315, 16'd35263, 16'd5325, 16'd51318, 16'd59285, 16'd9149, 16'd56042, 16'd40019, 16'd13880, 16'd46909, 16'd4964, 16'd28690, 16'd25227, 16'd26790, 16'd26295, 16'd56355, 16'd22307, 16'd44057, 16'd7685, 16'd25595, 16'd26191, 16'd27373, 16'd52609});
	test_expansion(128'hdcaa20e09e823996f5abe31c3471bd38, {16'd16885, 16'd62296, 16'd7166, 16'd14755, 16'd61525, 16'd23189, 16'd10546, 16'd59666, 16'd55859, 16'd56691, 16'd20940, 16'd11517, 16'd21498, 16'd48520, 16'd31183, 16'd51683, 16'd32153, 16'd3089, 16'd20145, 16'd6000, 16'd49045, 16'd8402, 16'd31715, 16'd51559, 16'd14570, 16'd42396});
	test_expansion(128'h6d2addb1b2f31ec0a0824f4cdfd7aa95, {16'd61964, 16'd35409, 16'd22495, 16'd5388, 16'd21583, 16'd52624, 16'd17390, 16'd12308, 16'd48031, 16'd16602, 16'd27899, 16'd57922, 16'd24067, 16'd37110, 16'd54183, 16'd58683, 16'd35508, 16'd14760, 16'd41338, 16'd6931, 16'd35738, 16'd28739, 16'd26141, 16'd54137, 16'd60550, 16'd11871});
	test_expansion(128'h6bd6e391c5d94d334a4961cf25d2d63a, {16'd34610, 16'd59718, 16'd45194, 16'd6908, 16'd32651, 16'd18740, 16'd8527, 16'd54330, 16'd38882, 16'd32879, 16'd18061, 16'd51443, 16'd5169, 16'd23996, 16'd64274, 16'd60830, 16'd11039, 16'd63558, 16'd23558, 16'd55778, 16'd16265, 16'd57681, 16'd3124, 16'd42481, 16'd5945, 16'd37406});
	test_expansion(128'h0dd19c74f94e8cfa6c6a5352c61b3cfc, {16'd38574, 16'd17637, 16'd17522, 16'd7703, 16'd33456, 16'd18672, 16'd59336, 16'd32841, 16'd61460, 16'd61292, 16'd13858, 16'd13192, 16'd41813, 16'd7630, 16'd46034, 16'd56581, 16'd4423, 16'd23923, 16'd28605, 16'd43784, 16'd1008, 16'd58450, 16'd1966, 16'd38677, 16'd63510, 16'd26378});
	test_expansion(128'he2262ba2898c9866beb81562a1b138c3, {16'd47459, 16'd6750, 16'd59795, 16'd32619, 16'd47260, 16'd33941, 16'd14945, 16'd30563, 16'd25709, 16'd35354, 16'd47031, 16'd60143, 16'd38896, 16'd50508, 16'd31677, 16'd59724, 16'd14859, 16'd5873, 16'd18545, 16'd54418, 16'd3632, 16'd24368, 16'd50908, 16'd59749, 16'd5479, 16'd2192});
	test_expansion(128'ha7f7a4539ca275ae92132b0e3fed2138, {16'd9889, 16'd7813, 16'd20784, 16'd59854, 16'd28458, 16'd47230, 16'd2995, 16'd54699, 16'd48759, 16'd31782, 16'd5740, 16'd40536, 16'd16463, 16'd2919, 16'd57838, 16'd41043, 16'd6141, 16'd44478, 16'd46874, 16'd16597, 16'd24320, 16'd64117, 16'd20909, 16'd62279, 16'd17051, 16'd14904});
	test_expansion(128'h55b385e503b6f41f93f387a29d2be140, {16'd10675, 16'd57718, 16'd20598, 16'd16602, 16'd41786, 16'd9166, 16'd46326, 16'd15893, 16'd9396, 16'd48475, 16'd6947, 16'd63082, 16'd13215, 16'd26692, 16'd11942, 16'd29013, 16'd65163, 16'd8439, 16'd53364, 16'd32641, 16'd53756, 16'd23614, 16'd41131, 16'd4719, 16'd2073, 16'd60298});
	test_expansion(128'hcfb2ff5700cf83562cb732559b92abdd, {16'd64834, 16'd5353, 16'd57927, 16'd32087, 16'd46953, 16'd59932, 16'd4349, 16'd422, 16'd61926, 16'd15836, 16'd58843, 16'd42272, 16'd50379, 16'd13409, 16'd56633, 16'd63634, 16'd14855, 16'd17332, 16'd59094, 16'd62968, 16'd41685, 16'd40818, 16'd6140, 16'd11356, 16'd23442, 16'd35916});
	test_expansion(128'h326da6b309799a8a377d2e6fd433ebdd, {16'd44389, 16'd57108, 16'd24597, 16'd61444, 16'd59197, 16'd34922, 16'd65170, 16'd7197, 16'd51772, 16'd31566, 16'd16337, 16'd46289, 16'd484, 16'd15048, 16'd15054, 16'd48237, 16'd978, 16'd24147, 16'd34029, 16'd21414, 16'd36067, 16'd43431, 16'd29781, 16'd51263, 16'd31330, 16'd10340});
	test_expansion(128'h9a2f383b34a6003972ab7e9b49cb30ac, {16'd40642, 16'd24679, 16'd13711, 16'd4288, 16'd735, 16'd33082, 16'd6492, 16'd24543, 16'd27129, 16'd6963, 16'd19364, 16'd10807, 16'd53224, 16'd36400, 16'd27568, 16'd33450, 16'd38622, 16'd18846, 16'd60580, 16'd52916, 16'd28961, 16'd21705, 16'd25685, 16'd38745, 16'd49601, 16'd14599});
	test_expansion(128'h2993739a577cb0749dfbd08def586136, {16'd42066, 16'd43485, 16'd26410, 16'd43880, 16'd25944, 16'd54938, 16'd32693, 16'd23717, 16'd50590, 16'd49485, 16'd48443, 16'd30034, 16'd44208, 16'd43996, 16'd7491, 16'd10909, 16'd40330, 16'd63808, 16'd55430, 16'd22414, 16'd24280, 16'd4482, 16'd37560, 16'd50242, 16'd10006, 16'd51051});
	test_expansion(128'h2b74e53aa3d9cd75af48c35d7918efb9, {16'd41207, 16'd44490, 16'd5499, 16'd56365, 16'd2009, 16'd58970, 16'd44798, 16'd6465, 16'd54959, 16'd18084, 16'd36121, 16'd58477, 16'd3036, 16'd63372, 16'd25768, 16'd28617, 16'd60429, 16'd9441, 16'd44956, 16'd14116, 16'd6699, 16'd11581, 16'd4899, 16'd3767, 16'd25742, 16'd11567});
	test_expansion(128'h50312f587b9dd1d70ab79c760275508e, {16'd17737, 16'd10646, 16'd61265, 16'd60736, 16'd1273, 16'd2207, 16'd14729, 16'd10536, 16'd51898, 16'd52003, 16'd42540, 16'd62307, 16'd4163, 16'd52133, 16'd57701, 16'd48928, 16'd38189, 16'd28541, 16'd31832, 16'd1713, 16'd28170, 16'd4352, 16'd30587, 16'd19392, 16'd31038, 16'd60373});
	test_expansion(128'h62aca92ef302f77fe6476b33a52abb40, {16'd5205, 16'd63334, 16'd65246, 16'd51582, 16'd61868, 16'd26317, 16'd39208, 16'd42268, 16'd18254, 16'd58493, 16'd6584, 16'd1638, 16'd35765, 16'd39913, 16'd3097, 16'd52738, 16'd6590, 16'd43394, 16'd15229, 16'd47263, 16'd63614, 16'd12398, 16'd649, 16'd40955, 16'd52714, 16'd55109});
	test_expansion(128'h393320649fe58b683c51c480fd1e9e84, {16'd57019, 16'd55159, 16'd724, 16'd30165, 16'd39442, 16'd48231, 16'd33502, 16'd49394, 16'd59256, 16'd23524, 16'd46062, 16'd55285, 16'd15228, 16'd37429, 16'd34104, 16'd61259, 16'd62225, 16'd36653, 16'd52168, 16'd36886, 16'd543, 16'd31269, 16'd24371, 16'd44838, 16'd8197, 16'd21105});
	test_expansion(128'hfd88bc6bce2bbc9be2901c67ab62b5c8, {16'd26350, 16'd65329, 16'd19587, 16'd41540, 16'd2110, 16'd51272, 16'd52792, 16'd63720, 16'd20750, 16'd31557, 16'd56979, 16'd65277, 16'd46450, 16'd57568, 16'd21985, 16'd63925, 16'd2660, 16'd27916, 16'd18822, 16'd27183, 16'd38016, 16'd28996, 16'd58692, 16'd6768, 16'd7645, 16'd32862});
	test_expansion(128'ha2d5a3af2b93da424e82408961ea17a4, {16'd63817, 16'd24668, 16'd44874, 16'd64161, 16'd50792, 16'd62155, 16'd743, 16'd57543, 16'd3983, 16'd35169, 16'd229, 16'd34125, 16'd39707, 16'd60985, 16'd24831, 16'd24423, 16'd43193, 16'd50236, 16'd12285, 16'd47085, 16'd21800, 16'd8070, 16'd33443, 16'd25744, 16'd51419, 16'd14404});
	test_expansion(128'h6fbaedecb62b5663ea64c5317c55ea7f, {16'd50219, 16'd3390, 16'd65390, 16'd58209, 16'd28489, 16'd60174, 16'd3554, 16'd16161, 16'd15627, 16'd29172, 16'd41263, 16'd35576, 16'd15933, 16'd56977, 16'd21494, 16'd26062, 16'd65340, 16'd16308, 16'd43722, 16'd3147, 16'd30550, 16'd14286, 16'd30163, 16'd19879, 16'd27677, 16'd27162});
	test_expansion(128'h9734bb88d9cd7a215c732dc231ceb31c, {16'd11855, 16'd18698, 16'd50812, 16'd40129, 16'd37891, 16'd49229, 16'd56941, 16'd60601, 16'd43058, 16'd43243, 16'd63657, 16'd37823, 16'd52050, 16'd52240, 16'd43881, 16'd53872, 16'd41523, 16'd630, 16'd56606, 16'd53839, 16'd13805, 16'd7039, 16'd51220, 16'd10663, 16'd53661, 16'd21361});
	test_expansion(128'ha4dbfe37bbf4c3736af0d79a963220af, {16'd25061, 16'd18097, 16'd62174, 16'd2802, 16'd44568, 16'd6142, 16'd44836, 16'd28579, 16'd16395, 16'd31034, 16'd60125, 16'd54531, 16'd52511, 16'd58997, 16'd50436, 16'd2569, 16'd64630, 16'd35270, 16'd31930, 16'd19018, 16'd1458, 16'd52487, 16'd521, 16'd23835, 16'd28280, 16'd24892});
	test_expansion(128'hd896bf05fdc3d781f9911c886be51a87, {16'd21246, 16'd46835, 16'd64866, 16'd57377, 16'd25386, 16'd29735, 16'd58487, 16'd46542, 16'd3314, 16'd2665, 16'd28365, 16'd28094, 16'd60438, 16'd1446, 16'd2796, 16'd17769, 16'd36478, 16'd36012, 16'd46959, 16'd529, 16'd29713, 16'd47296, 16'd7684, 16'd42787, 16'd7317, 16'd62725});
	test_expansion(128'h73c052b2c9a5aed8d5fc91e48408caac, {16'd5221, 16'd53519, 16'd21702, 16'd42113, 16'd13921, 16'd56553, 16'd14166, 16'd61301, 16'd32725, 16'd21818, 16'd13745, 16'd13360, 16'd37379, 16'd57529, 16'd25756, 16'd8888, 16'd65065, 16'd32786, 16'd10190, 16'd50458, 16'd21654, 16'd63106, 16'd19865, 16'd44836, 16'd25326, 16'd6417});
	test_expansion(128'h47a3eacb8d4e8fb2d4b2c6aaff2670c0, {16'd27058, 16'd39202, 16'd45761, 16'd4813, 16'd10843, 16'd21965, 16'd41924, 16'd54801, 16'd42269, 16'd42471, 16'd50693, 16'd32021, 16'd21748, 16'd59189, 16'd58551, 16'd23649, 16'd13731, 16'd44112, 16'd60686, 16'd13797, 16'd2334, 16'd49343, 16'd61072, 16'd55949, 16'd49680, 16'd43579});
	test_expansion(128'hfa156ceb63ae42cbf09e3c1101531a34, {16'd53706, 16'd23531, 16'd42270, 16'd27167, 16'd4209, 16'd42088, 16'd27221, 16'd63636, 16'd33808, 16'd49424, 16'd20733, 16'd6703, 16'd64081, 16'd40415, 16'd60194, 16'd22485, 16'd20494, 16'd63331, 16'd18506, 16'd21767, 16'd61934, 16'd40904, 16'd29625, 16'd20929, 16'd14436, 16'd57177});
	test_expansion(128'h932bfb779d92783f8de0c6d57aaa8cff, {16'd49086, 16'd41950, 16'd47870, 16'd19528, 16'd12233, 16'd8433, 16'd24163, 16'd22973, 16'd34056, 16'd49472, 16'd35214, 16'd27608, 16'd52023, 16'd5648, 16'd50666, 16'd36695, 16'd22386, 16'd60391, 16'd25263, 16'd41772, 16'd20184, 16'd28545, 16'd33879, 16'd10315, 16'd36163, 16'd4296});
	test_expansion(128'hbfd59e53893743591f3fffc3a587d1dd, {16'd51516, 16'd21173, 16'd29932, 16'd8098, 16'd50156, 16'd44269, 16'd37470, 16'd31641, 16'd61145, 16'd61617, 16'd6500, 16'd26120, 16'd25577, 16'd50463, 16'd54242, 16'd38771, 16'd61191, 16'd35204, 16'd57824, 16'd59344, 16'd34971, 16'd29313, 16'd45776, 16'd25080, 16'd22374, 16'd60169});
	test_expansion(128'h01615bb5a1d92d81b8e226b2c5c86c98, {16'd1164, 16'd49232, 16'd51025, 16'd26995, 16'd5528, 16'd12051, 16'd54427, 16'd29683, 16'd37229, 16'd19042, 16'd35525, 16'd4504, 16'd53404, 16'd47376, 16'd60163, 16'd12013, 16'd11083, 16'd7872, 16'd6300, 16'd55230, 16'd60479, 16'd42600, 16'd2475, 16'd27694, 16'd4926, 16'd28702});
	test_expansion(128'h377f7bbea7b6a5cd036834030eefef47, {16'd7000, 16'd4571, 16'd37114, 16'd5128, 16'd17094, 16'd15585, 16'd30685, 16'd55175, 16'd12056, 16'd29629, 16'd1874, 16'd42035, 16'd34465, 16'd40342, 16'd51785, 16'd13168, 16'd58416, 16'd54025, 16'd47664, 16'd63153, 16'd13236, 16'd63232, 16'd10536, 16'd22912, 16'd48367, 16'd39568});
	test_expansion(128'h14137c97d8d12f6bf8f6a7d7d2cd7b38, {16'd17799, 16'd58290, 16'd54368, 16'd32647, 16'd5812, 16'd13006, 16'd36539, 16'd39429, 16'd48290, 16'd19416, 16'd18450, 16'd25233, 16'd5367, 16'd21777, 16'd59575, 16'd12617, 16'd11682, 16'd17739, 16'd60006, 16'd7191, 16'd58285, 16'd54, 16'd3951, 16'd16841, 16'd29475, 16'd8587});
	test_expansion(128'h6e9f567f79a81909be8bb5eec11a929f, {16'd57267, 16'd45663, 16'd25100, 16'd24514, 16'd9360, 16'd5742, 16'd20943, 16'd38069, 16'd939, 16'd8072, 16'd2811, 16'd25142, 16'd21544, 16'd63452, 16'd18916, 16'd61766, 16'd30243, 16'd49043, 16'd34305, 16'd10230, 16'd25490, 16'd8735, 16'd19875, 16'd17015, 16'd14569, 16'd1777});
	test_expansion(128'h227533437f0cc372674e6976f78c9baf, {16'd25016, 16'd27345, 16'd30258, 16'd29656, 16'd60625, 16'd20595, 16'd52708, 16'd18288, 16'd23965, 16'd49080, 16'd51137, 16'd56280, 16'd9839, 16'd8005, 16'd54696, 16'd32675, 16'd54338, 16'd63285, 16'd60641, 16'd11577, 16'd1610, 16'd27053, 16'd45147, 16'd20751, 16'd58464, 16'd53163});
	test_expansion(128'h28b37c66abfbf6cf88c25885126b8ea5, {16'd12950, 16'd54177, 16'd11090, 16'd6513, 16'd10670, 16'd31499, 16'd36229, 16'd58705, 16'd15964, 16'd57193, 16'd57101, 16'd38447, 16'd9182, 16'd2640, 16'd53780, 16'd30021, 16'd60520, 16'd53123, 16'd52305, 16'd12498, 16'd49231, 16'd23795, 16'd49798, 16'd3532, 16'd64888, 16'd47143});
	test_expansion(128'ha5fec3956f5fbec20b7a0ef3deb8cffe, {16'd8574, 16'd54596, 16'd7411, 16'd5382, 16'd13718, 16'd38936, 16'd3932, 16'd32012, 16'd36885, 16'd58941, 16'd29590, 16'd17475, 16'd823, 16'd11073, 16'd54084, 16'd6887, 16'd27050, 16'd21001, 16'd24113, 16'd57718, 16'd56427, 16'd10472, 16'd21375, 16'd7305, 16'd20313, 16'd3695});
	test_expansion(128'he08997e439dd34cec0060090df2180ab, {16'd60298, 16'd8556, 16'd56067, 16'd1644, 16'd34668, 16'd4389, 16'd47663, 16'd27902, 16'd57683, 16'd24328, 16'd13863, 16'd27833, 16'd43078, 16'd36596, 16'd4676, 16'd63410, 16'd24441, 16'd53238, 16'd37493, 16'd59681, 16'd5964, 16'd3996, 16'd60606, 16'd53387, 16'd40092, 16'd34056});
	test_expansion(128'hc51d370e2783e14cf66b4d3318175915, {16'd34116, 16'd28348, 16'd9637, 16'd28139, 16'd28424, 16'd30700, 16'd23923, 16'd16975, 16'd53747, 16'd50935, 16'd58441, 16'd13980, 16'd8295, 16'd1512, 16'd2294, 16'd15948, 16'd48470, 16'd40172, 16'd999, 16'd36695, 16'd10490, 16'd1490, 16'd59470, 16'd16779, 16'd6312, 16'd8360});
	test_expansion(128'h1d8dfa11c6aaaf64aa7cfe9fd8715f0c, {16'd10330, 16'd38558, 16'd48517, 16'd6753, 16'd1592, 16'd47814, 16'd63586, 16'd42765, 16'd47981, 16'd8076, 16'd31286, 16'd53145, 16'd47864, 16'd22519, 16'd7354, 16'd10562, 16'd454, 16'd10565, 16'd57780, 16'd28631, 16'd23695, 16'd28078, 16'd53902, 16'd54260, 16'd52049, 16'd45402});
	test_expansion(128'h77df919b895297e36286bc68ffbf00b3, {16'd6368, 16'd7446, 16'd59877, 16'd50242, 16'd30582, 16'd35011, 16'd36893, 16'd49760, 16'd64506, 16'd11294, 16'd7559, 16'd45230, 16'd29612, 16'd3799, 16'd39648, 16'd19152, 16'd13096, 16'd24841, 16'd24926, 16'd53691, 16'd58904, 16'd31205, 16'd943, 16'd52906, 16'd24287, 16'd18025});
	test_expansion(128'h241b404984ede2b5eaa77c2f62a1dccf, {16'd12297, 16'd52307, 16'd30437, 16'd61160, 16'd50717, 16'd25770, 16'd30399, 16'd28217, 16'd34830, 16'd28493, 16'd11535, 16'd62858, 16'd4113, 16'd65137, 16'd60271, 16'd43635, 16'd41138, 16'd52565, 16'd5219, 16'd38207, 16'd54240, 16'd12879, 16'd35023, 16'd26348, 16'd741, 16'd3892});
	test_expansion(128'h9989222e8d49db7a32e6805dd84cccfb, {16'd19188, 16'd4498, 16'd26350, 16'd55374, 16'd59243, 16'd3449, 16'd54674, 16'd58957, 16'd43643, 16'd8414, 16'd44165, 16'd1512, 16'd7550, 16'd43845, 16'd46058, 16'd50533, 16'd65252, 16'd31112, 16'd48906, 16'd58292, 16'd34461, 16'd63102, 16'd53759, 16'd46728, 16'd15523, 16'd47278});
	test_expansion(128'hb8c9a2700e2e6592fd574dff542a7527, {16'd14498, 16'd44295, 16'd24660, 16'd48250, 16'd48841, 16'd57493, 16'd4543, 16'd37710, 16'd57856, 16'd38083, 16'd2015, 16'd34936, 16'd50511, 16'd36504, 16'd34820, 16'd39730, 16'd25161, 16'd16115, 16'd47901, 16'd37790, 16'd39905, 16'd12798, 16'd33953, 16'd35663, 16'd39553, 16'd9151});
	test_expansion(128'h8fc7d09dad6ee7fa362803069b4bde8f, {16'd63383, 16'd33033, 16'd31061, 16'd12569, 16'd28996, 16'd40759, 16'd30629, 16'd6781, 16'd8799, 16'd35757, 16'd53792, 16'd36797, 16'd25139, 16'd20617, 16'd37729, 16'd30213, 16'd59086, 16'd19084, 16'd63681, 16'd21308, 16'd37711, 16'd49748, 16'd49241, 16'd40873, 16'd18096, 16'd24476});
	test_expansion(128'h681fa42e5adabcf4d93de9ffd6289fe4, {16'd14361, 16'd53896, 16'd16933, 16'd32723, 16'd36361, 16'd47912, 16'd64965, 16'd61441, 16'd60359, 16'd4742, 16'd1826, 16'd13517, 16'd22861, 16'd32176, 16'd58651, 16'd18801, 16'd5929, 16'd28055, 16'd43563, 16'd23953, 16'd55853, 16'd22334, 16'd34116, 16'd60394, 16'd62561, 16'd26710});
	test_expansion(128'h555484d3f2834e8c2435d03156ba52d1, {16'd46631, 16'd36168, 16'd3416, 16'd55151, 16'd58205, 16'd5415, 16'd62493, 16'd46992, 16'd17805, 16'd48016, 16'd14090, 16'd23855, 16'd54832, 16'd6556, 16'd49150, 16'd63261, 16'd32888, 16'd21880, 16'd57761, 16'd41647, 16'd24377, 16'd27870, 16'd13477, 16'd1119, 16'd18456, 16'd51291});
	test_expansion(128'h017f5e8f7391323e85c98d2caad19034, {16'd34189, 16'd3057, 16'd45038, 16'd6825, 16'd43669, 16'd34596, 16'd337, 16'd17921, 16'd26713, 16'd25016, 16'd32722, 16'd65377, 16'd18590, 16'd40610, 16'd20057, 16'd16292, 16'd43401, 16'd56929, 16'd17326, 16'd14154, 16'd55502, 16'd15307, 16'd58958, 16'd57682, 16'd26403, 16'd26133});
	test_expansion(128'h7af02a0d6ab6c985e286ff2369f92ccc, {16'd5157, 16'd18662, 16'd11299, 16'd64039, 16'd39468, 16'd32042, 16'd36704, 16'd59265, 16'd17475, 16'd15819, 16'd65271, 16'd64681, 16'd13954, 16'd25583, 16'd29649, 16'd51841, 16'd31533, 16'd363, 16'd56398, 16'd42652, 16'd53198, 16'd38626, 16'd26904, 16'd12271, 16'd62775, 16'd50597});
	test_expansion(128'h79cec258902b2b01b393bfa54f336256, {16'd19873, 16'd35888, 16'd20929, 16'd4356, 16'd17434, 16'd33715, 16'd18072, 16'd18800, 16'd59486, 16'd39023, 16'd1708, 16'd54622, 16'd62495, 16'd906, 16'd52937, 16'd1023, 16'd1012, 16'd34755, 16'd43004, 16'd7761, 16'd32320, 16'd43172, 16'd26736, 16'd58257, 16'd38659, 16'd18220});
	test_expansion(128'h037d3c72cb1398b1423a348b78def4f1, {16'd31531, 16'd38574, 16'd53878, 16'd16659, 16'd5199, 16'd23148, 16'd56893, 16'd1868, 16'd46794, 16'd14268, 16'd8654, 16'd31890, 16'd2730, 16'd57195, 16'd6432, 16'd57821, 16'd59614, 16'd17838, 16'd22719, 16'd43174, 16'd44009, 16'd1052, 16'd42331, 16'd56575, 16'd51629, 16'd50481});
	test_expansion(128'h31026f9beb5856ef5effbf55def08de0, {16'd27315, 16'd23205, 16'd40883, 16'd14780, 16'd58041, 16'd20922, 16'd60777, 16'd20253, 16'd62442, 16'd49067, 16'd50681, 16'd17400, 16'd9907, 16'd6945, 16'd54836, 16'd24635, 16'd10572, 16'd61721, 16'd19472, 16'd8013, 16'd31691, 16'd12683, 16'd56918, 16'd28586, 16'd1577, 16'd27536});
	test_expansion(128'h1e69175fc95b971e405044e26a3aac19, {16'd366, 16'd1022, 16'd11761, 16'd5410, 16'd40913, 16'd47970, 16'd28147, 16'd60878, 16'd35353, 16'd4614, 16'd58485, 16'd12930, 16'd24276, 16'd44941, 16'd15865, 16'd39112, 16'd32211, 16'd4214, 16'd8587, 16'd35376, 16'd60722, 16'd25046, 16'd39715, 16'd7316, 16'd21066, 16'd13274});
	test_expansion(128'he714d2d5e443d943ad8f2a345b87ef72, {16'd849, 16'd40443, 16'd9757, 16'd51079, 16'd36280, 16'd64754, 16'd18016, 16'd21798, 16'd34612, 16'd28293, 16'd41661, 16'd57843, 16'd57116, 16'd30914, 16'd29192, 16'd14945, 16'd51742, 16'd40679, 16'd29780, 16'd1583, 16'd40217, 16'd3170, 16'd59324, 16'd39576, 16'd11048, 16'd14169});
	test_expansion(128'h2ade9be294b48418fe67ffcdf68243f7, {16'd35971, 16'd4531, 16'd10364, 16'd26275, 16'd30090, 16'd4617, 16'd52155, 16'd13610, 16'd5443, 16'd32920, 16'd28846, 16'd33018, 16'd63226, 16'd28492, 16'd59360, 16'd44745, 16'd62682, 16'd52999, 16'd931, 16'd10765, 16'd14788, 16'd60980, 16'd22929, 16'd57870, 16'd5989, 16'd12918});
	test_expansion(128'hf9991af1490baecc49764f540c60cacf, {16'd46944, 16'd25485, 16'd32008, 16'd28436, 16'd18248, 16'd16979, 16'd17088, 16'd37654, 16'd51425, 16'd19958, 16'd39183, 16'd48466, 16'd64640, 16'd47848, 16'd53533, 16'd62847, 16'd19793, 16'd28713, 16'd58457, 16'd32752, 16'd64084, 16'd54102, 16'd20736, 16'd41578, 16'd26697, 16'd62231});
	test_expansion(128'h12c8ed61809e29489c046cf0f7f3d3c5, {16'd3540, 16'd54908, 16'd41417, 16'd47389, 16'd22818, 16'd50682, 16'd40962, 16'd37189, 16'd6534, 16'd39143, 16'd39451, 16'd50301, 16'd10116, 16'd31002, 16'd49682, 16'd11791, 16'd4127, 16'd64833, 16'd48435, 16'd57703, 16'd55301, 16'd20467, 16'd53451, 16'd50449, 16'd13728, 16'd3037});
	test_expansion(128'hf53b2f446459c3919b9ff4cf3e9595e8, {16'd54199, 16'd46462, 16'd20123, 16'd44860, 16'd46169, 16'd35686, 16'd22286, 16'd39820, 16'd55534, 16'd58389, 16'd58690, 16'd1237, 16'd16389, 16'd45822, 16'd12406, 16'd7481, 16'd64131, 16'd62595, 16'd55605, 16'd16005, 16'd37679, 16'd48766, 16'd45443, 16'd35278, 16'd37294, 16'd41672});
	test_expansion(128'hb4d2cb6259b2a2d8814e8ac1ef4c9454, {16'd51970, 16'd61912, 16'd26422, 16'd34792, 16'd47664, 16'd58453, 16'd35625, 16'd40431, 16'd38736, 16'd54144, 16'd47135, 16'd47042, 16'd11292, 16'd47815, 16'd20012, 16'd58850, 16'd21441, 16'd47621, 16'd33593, 16'd43015, 16'd22529, 16'd55549, 16'd62786, 16'd11842, 16'd54386, 16'd8670});
	test_expansion(128'h9517372ee9f0a7a83bf40abbfa8cc184, {16'd52026, 16'd53558, 16'd61471, 16'd37901, 16'd62833, 16'd35492, 16'd19906, 16'd1683, 16'd28139, 16'd26789, 16'd21537, 16'd64392, 16'd26260, 16'd3299, 16'd46239, 16'd21805, 16'd16156, 16'd11486, 16'd30081, 16'd16421, 16'd35201, 16'd61954, 16'd49610, 16'd57625, 16'd5754, 16'd54290});
	test_expansion(128'h4d80ac3a4d2a1fbd0640c04d0f88fca8, {16'd15357, 16'd6429, 16'd14027, 16'd14483, 16'd18393, 16'd29528, 16'd19953, 16'd4912, 16'd21965, 16'd51626, 16'd58034, 16'd60899, 16'd60963, 16'd45186, 16'd24529, 16'd34822, 16'd31236, 16'd25949, 16'd14441, 16'd49366, 16'd16971, 16'd46382, 16'd13277, 16'd11285, 16'd21518, 16'd14820});
	test_expansion(128'he62c6449c2994d0e6ac86606f6a3fffa, {16'd62500, 16'd12377, 16'd41998, 16'd16597, 16'd48175, 16'd29723, 16'd8291, 16'd45373, 16'd34537, 16'd60436, 16'd10085, 16'd30426, 16'd43050, 16'd46373, 16'd3704, 16'd57904, 16'd65023, 16'd9169, 16'd58857, 16'd37953, 16'd17696, 16'd15236, 16'd21341, 16'd24179, 16'd63900, 16'd60697});
	test_expansion(128'h520670a5f79fbc7e450be58c5bf28d1a, {16'd28697, 16'd13403, 16'd64493, 16'd44285, 16'd11614, 16'd48991, 16'd40102, 16'd52384, 16'd18596, 16'd11506, 16'd62979, 16'd6836, 16'd46729, 16'd64197, 16'd4766, 16'd28389, 16'd25490, 16'd58726, 16'd60732, 16'd47214, 16'd39366, 16'd22185, 16'd61497, 16'd33480, 16'd41518, 16'd63340});
	test_expansion(128'hcd7e544ce8452ded47ab40d2ddda8541, {16'd34657, 16'd58628, 16'd12138, 16'd63448, 16'd41269, 16'd54873, 16'd3704, 16'd13934, 16'd14561, 16'd45910, 16'd14388, 16'd55400, 16'd54436, 16'd27277, 16'd62346, 16'd18499, 16'd13555, 16'd28521, 16'd18348, 16'd55707, 16'd52777, 16'd16530, 16'd37405, 16'd59273, 16'd24197, 16'd5179});
	test_expansion(128'hd3b31f32f0663024bac4d910abfdb2a7, {16'd22695, 16'd16006, 16'd12202, 16'd61294, 16'd45863, 16'd3215, 16'd14049, 16'd61653, 16'd48398, 16'd2242, 16'd49600, 16'd18713, 16'd51426, 16'd3438, 16'd11393, 16'd48542, 16'd7259, 16'd61330, 16'd28236, 16'd42774, 16'd19491, 16'd8408, 16'd1005, 16'd2785, 16'd10343, 16'd44642});
	test_expansion(128'h8b4814398f52b91baaa9acf282532130, {16'd39292, 16'd8825, 16'd48345, 16'd41517, 16'd60511, 16'd32644, 16'd23553, 16'd60385, 16'd28583, 16'd15780, 16'd7127, 16'd22001, 16'd674, 16'd16598, 16'd62211, 16'd16985, 16'd31123, 16'd5624, 16'd31972, 16'd50285, 16'd4861, 16'd56431, 16'd35511, 16'd32035, 16'd1753, 16'd33720});
	test_expansion(128'h9a8d025c5c365bd4a6edd9ee8dfa0bb8, {16'd51489, 16'd46572, 16'd36223, 16'd39992, 16'd36088, 16'd30462, 16'd44325, 16'd63047, 16'd31301, 16'd10578, 16'd37766, 16'd42718, 16'd65444, 16'd27023, 16'd16408, 16'd15225, 16'd40511, 16'd56644, 16'd21527, 16'd48248, 16'd54908, 16'd30371, 16'd40635, 16'd4316, 16'd64765, 16'd31345});
	test_expansion(128'h2603060d2ca9db9d5372bf957edee89c, {16'd26251, 16'd6615, 16'd36993, 16'd46280, 16'd2905, 16'd17040, 16'd40713, 16'd32061, 16'd43747, 16'd27602, 16'd4499, 16'd8493, 16'd51413, 16'd23850, 16'd32468, 16'd58149, 16'd6442, 16'd23422, 16'd41937, 16'd8004, 16'd59266, 16'd17047, 16'd44546, 16'd28393, 16'd50099, 16'd37524});
	test_expansion(128'hc1cfe6c5f41f6e985e2283fdfabbb682, {16'd55404, 16'd21836, 16'd28456, 16'd35113, 16'd14260, 16'd56414, 16'd29535, 16'd47670, 16'd36977, 16'd15701, 16'd36095, 16'd64466, 16'd48612, 16'd37144, 16'd26479, 16'd37821, 16'd26625, 16'd53541, 16'd58943, 16'd30533, 16'd25813, 16'd6849, 16'd5381, 16'd52051, 16'd54408, 16'd5608});
	test_expansion(128'hf23513fc3b914e241d3873d8eca3d889, {16'd51023, 16'd60089, 16'd39376, 16'd63877, 16'd13985, 16'd39174, 16'd28185, 16'd25476, 16'd47868, 16'd20608, 16'd22555, 16'd7471, 16'd7605, 16'd355, 16'd6483, 16'd5037, 16'd854, 16'd19702, 16'd52592, 16'd14314, 16'd29114, 16'd45212, 16'd4694, 16'd36918, 16'd17195, 16'd22109});
	test_expansion(128'h4328b147d6c3235733f2ac8733bc1996, {16'd29141, 16'd47175, 16'd57563, 16'd39174, 16'd55359, 16'd967, 16'd15645, 16'd16964, 16'd39838, 16'd51853, 16'd40064, 16'd9641, 16'd22581, 16'd31979, 16'd16147, 16'd22716, 16'd93, 16'd23697, 16'd53525, 16'd42364, 16'd9841, 16'd21986, 16'd47502, 16'd6415, 16'd54231, 16'd20364});
	test_expansion(128'h2eb169269672e62d260b44a79ab74060, {16'd13207, 16'd34211, 16'd33678, 16'd29270, 16'd4987, 16'd41124, 16'd34787, 16'd57990, 16'd37960, 16'd22397, 16'd62044, 16'd13020, 16'd29014, 16'd52630, 16'd45292, 16'd59598, 16'd6994, 16'd58004, 16'd60005, 16'd14909, 16'd22135, 16'd62193, 16'd2656, 16'd17589, 16'd62534, 16'd54090});
	test_expansion(128'h7b2e04d2f721b7b6b8ed04f0905576ca, {16'd52843, 16'd18423, 16'd17606, 16'd54252, 16'd57804, 16'd45895, 16'd56584, 16'd41704, 16'd24148, 16'd18097, 16'd17406, 16'd64977, 16'd46209, 16'd942, 16'd5976, 16'd53880, 16'd49841, 16'd38772, 16'd17201, 16'd24010, 16'd14853, 16'd18483, 16'd19948, 16'd44167, 16'd40430, 16'd17485});
	test_expansion(128'h6562dff7fdb9ddcc4c371c7e48900912, {16'd27296, 16'd40909, 16'd58089, 16'd51336, 16'd23107, 16'd27983, 16'd47858, 16'd47755, 16'd22419, 16'd29131, 16'd41064, 16'd24068, 16'd51558, 16'd52851, 16'd47102, 16'd48148, 16'd11341, 16'd36010, 16'd51783, 16'd561, 16'd8281, 16'd2769, 16'd3465, 16'd21468, 16'd10381, 16'd47910});
	test_expansion(128'h3c8eca87792ddedeaf566862e0025081, {16'd20512, 16'd3904, 16'd6039, 16'd4283, 16'd47244, 16'd50800, 16'd18565, 16'd60144, 16'd12848, 16'd65535, 16'd47396, 16'd39074, 16'd47262, 16'd30160, 16'd30535, 16'd55601, 16'd13524, 16'd58401, 16'd64182, 16'd50335, 16'd49022, 16'd33894, 16'd48236, 16'd18723, 16'd9351, 16'd22033});
	test_expansion(128'h9a199364144a622edf7edcce2c768528, {16'd5094, 16'd12377, 16'd19678, 16'd28450, 16'd37802, 16'd23336, 16'd37732, 16'd59032, 16'd55626, 16'd29855, 16'd13835, 16'd48483, 16'd15182, 16'd37064, 16'd24524, 16'd7660, 16'd24299, 16'd28054, 16'd50156, 16'd48775, 16'd16260, 16'd34919, 16'd1207, 16'd23367, 16'd22775, 16'd44824});
	test_expansion(128'h112f52c345e1a8d415b9d4e78149d63a, {16'd2029, 16'd29030, 16'd27427, 16'd2253, 16'd35782, 16'd54382, 16'd21457, 16'd54258, 16'd28624, 16'd676, 16'd34344, 16'd53284, 16'd23538, 16'd50872, 16'd18840, 16'd35937, 16'd12537, 16'd62261, 16'd44494, 16'd22042, 16'd44623, 16'd58059, 16'd20740, 16'd54362, 16'd36890, 16'd59461});
	test_expansion(128'h73d3dc64cadc1b87b2127cd9a70721ee, {16'd791, 16'd38548, 16'd28995, 16'd6259, 16'd65013, 16'd56633, 16'd2910, 16'd22374, 16'd32810, 16'd38670, 16'd63152, 16'd33230, 16'd1111, 16'd45034, 16'd16372, 16'd12089, 16'd26908, 16'd34959, 16'd31759, 16'd2649, 16'd24209, 16'd49654, 16'd33501, 16'd58014, 16'd18558, 16'd43215});
	test_expansion(128'h1cb807d047284e4c2ba7c55e20c9f498, {16'd48025, 16'd21779, 16'd62561, 16'd18752, 16'd1991, 16'd40574, 16'd3581, 16'd16817, 16'd46310, 16'd50148, 16'd49588, 16'd52887, 16'd6702, 16'd51103, 16'd29205, 16'd4280, 16'd55521, 16'd44833, 16'd40870, 16'd42464, 16'd35823, 16'd59704, 16'd4133, 16'd7583, 16'd59924, 16'd27150});
	test_expansion(128'h7bcb52d7a48b35645599eb2b9c34b534, {16'd61565, 16'd46721, 16'd1040, 16'd57274, 16'd49619, 16'd7480, 16'd22165, 16'd22914, 16'd61906, 16'd6025, 16'd53317, 16'd57246, 16'd23232, 16'd45412, 16'd8526, 16'd18946, 16'd36072, 16'd18251, 16'd3640, 16'd17221, 16'd48835, 16'd61011, 16'd59927, 16'd30007, 16'd6585, 16'd34175});
	test_expansion(128'h9852e9f32a6b4a49f3ba21a9b8dff2ec, {16'd58482, 16'd48373, 16'd41371, 16'd54941, 16'd2176, 16'd24994, 16'd13429, 16'd31220, 16'd64041, 16'd20025, 16'd312, 16'd16995, 16'd43478, 16'd53082, 16'd39650, 16'd34896, 16'd23731, 16'd62735, 16'd1868, 16'd18346, 16'd40628, 16'd49121, 16'd63679, 16'd38752, 16'd42914, 16'd34321});
	test_expansion(128'ha61501b0e54d2eb876715a36c52d1071, {16'd12238, 16'd21160, 16'd8800, 16'd29507, 16'd12815, 16'd17882, 16'd25290, 16'd17021, 16'd10308, 16'd27957, 16'd46304, 16'd50086, 16'd39933, 16'd44670, 16'd3706, 16'd27467, 16'd59660, 16'd10040, 16'd6711, 16'd25237, 16'd17364, 16'd52158, 16'd63480, 16'd16377, 16'd22792, 16'd54604});
	test_expansion(128'h79d5b7c0ce0b004a2f303e3077210b50, {16'd63521, 16'd17662, 16'd50698, 16'd24695, 16'd6760, 16'd35572, 16'd14993, 16'd53526, 16'd13402, 16'd12185, 16'd23325, 16'd33710, 16'd30781, 16'd4339, 16'd30323, 16'd23523, 16'd61912, 16'd60021, 16'd16287, 16'd28297, 16'd46605, 16'd52932, 16'd259, 16'd61549, 16'd3167, 16'd34141});
	test_expansion(128'h598269ebb12fcb24c0daaecc72069b82, {16'd32034, 16'd58525, 16'd63464, 16'd55775, 16'd10664, 16'd30884, 16'd18059, 16'd20704, 16'd33394, 16'd8926, 16'd63686, 16'd2578, 16'd46191, 16'd11726, 16'd63184, 16'd26544, 16'd32974, 16'd36017, 16'd16746, 16'd653, 16'd10772, 16'd60917, 16'd64652, 16'd47235, 16'd34525, 16'd51362});
	test_expansion(128'h821b3d6cf36f4f0afcc1b704a7518bd4, {16'd36825, 16'd36237, 16'd2635, 16'd2561, 16'd28254, 16'd6955, 16'd10030, 16'd13343, 16'd37802, 16'd42758, 16'd64395, 16'd6543, 16'd6101, 16'd31290, 16'd52683, 16'd32058, 16'd17344, 16'd49784, 16'd61925, 16'd18861, 16'd16199, 16'd11621, 16'd58741, 16'd20044, 16'd3852, 16'd30108});
	test_expansion(128'ha4dd4103c32f0d0926ffcf44f3a8127b, {16'd26901, 16'd1261, 16'd65358, 16'd61281, 16'd21798, 16'd13823, 16'd10677, 16'd51860, 16'd41667, 16'd4709, 16'd25369, 16'd300, 16'd43946, 16'd15109, 16'd13342, 16'd12054, 16'd45337, 16'd19113, 16'd56691, 16'd15452, 16'd2427, 16'd31752, 16'd27694, 16'd4397, 16'd52322, 16'd36637});
	test_expansion(128'h9fcea1e5a8f65463cd548124d96db926, {16'd16550, 16'd1382, 16'd23401, 16'd29170, 16'd34395, 16'd53518, 16'd55410, 16'd41421, 16'd42638, 16'd40140, 16'd18038, 16'd18794, 16'd57437, 16'd10799, 16'd3654, 16'd28771, 16'd56754, 16'd64836, 16'd60769, 16'd63616, 16'd9357, 16'd44885, 16'd7597, 16'd63313, 16'd8164, 16'd13183});
	test_expansion(128'h7b7fd1c8f7fcf04fcf83aa671d635d0e, {16'd21619, 16'd60512, 16'd17788, 16'd13995, 16'd49053, 16'd29655, 16'd25849, 16'd54608, 16'd46703, 16'd24847, 16'd10731, 16'd55752, 16'd55330, 16'd30984, 16'd48327, 16'd61487, 16'd12595, 16'd42323, 16'd60773, 16'd46454, 16'd8550, 16'd55194, 16'd14241, 16'd34728, 16'd26910, 16'd48454});
	test_expansion(128'ha3c90f8785f15c640778a35030c3dc88, {16'd1820, 16'd33208, 16'd1292, 16'd17116, 16'd51442, 16'd37923, 16'd53481, 16'd37496, 16'd29974, 16'd43991, 16'd30275, 16'd4007, 16'd51960, 16'd3742, 16'd31119, 16'd41116, 16'd17759, 16'd19917, 16'd13215, 16'd30308, 16'd34269, 16'd57583, 16'd29901, 16'd36824, 16'd40366, 16'd30108});
	test_expansion(128'h2d5f258ff4381f45df7253536a1a0fc8, {16'd53018, 16'd60035, 16'd36123, 16'd6623, 16'd20916, 16'd54487, 16'd58839, 16'd33188, 16'd32785, 16'd22080, 16'd13987, 16'd60229, 16'd43141, 16'd26654, 16'd26228, 16'd61404, 16'd56237, 16'd10242, 16'd57037, 16'd34023, 16'd20059, 16'd12265, 16'd24074, 16'd51211, 16'd10586, 16'd5213});
	test_expansion(128'hed976210677db10ca327b06cb0146c4f, {16'd33562, 16'd57138, 16'd3730, 16'd61427, 16'd44503, 16'd8579, 16'd26431, 16'd49780, 16'd40613, 16'd53420, 16'd32694, 16'd29880, 16'd57680, 16'd60916, 16'd60027, 16'd34669, 16'd57872, 16'd26033, 16'd34720, 16'd33156, 16'd59923, 16'd24536, 16'd2972, 16'd60561, 16'd25895, 16'd35945});
	test_expansion(128'hb91f8761219dd44f78572757fdf1b4ad, {16'd32494, 16'd46435, 16'd24779, 16'd32630, 16'd39903, 16'd10569, 16'd34446, 16'd41652, 16'd28403, 16'd37572, 16'd60414, 16'd31553, 16'd17367, 16'd31549, 16'd41669, 16'd28203, 16'd21964, 16'd23983, 16'd35152, 16'd45594, 16'd24955, 16'd56461, 16'd27213, 16'd41507, 16'd10663, 16'd13281});
	test_expansion(128'hee285c4a00f05793e020f9f0728b369f, {16'd17614, 16'd23997, 16'd12871, 16'd11467, 16'd16673, 16'd13145, 16'd44431, 16'd28740, 16'd46612, 16'd58425, 16'd60485, 16'd49644, 16'd12452, 16'd34020, 16'd59211, 16'd1136, 16'd22576, 16'd44210, 16'd51764, 16'd9707, 16'd34859, 16'd22596, 16'd24934, 16'd17396, 16'd28095, 16'd46283});
	test_expansion(128'h88a4d530624691d3bb99f19d7b714b22, {16'd22034, 16'd37267, 16'd54826, 16'd23398, 16'd14192, 16'd1615, 16'd30013, 16'd3007, 16'd57164, 16'd22691, 16'd63308, 16'd25979, 16'd32352, 16'd36503, 16'd12658, 16'd32270, 16'd19517, 16'd6833, 16'd51888, 16'd7740, 16'd19667, 16'd20883, 16'd21826, 16'd3502, 16'd26570, 16'd49385});
	test_expansion(128'h99c958aed1df724993cea3a7187957e4, {16'd16886, 16'd37030, 16'd48263, 16'd8729, 16'd59694, 16'd1117, 16'd41519, 16'd46301, 16'd64509, 16'd16618, 16'd14446, 16'd18623, 16'd57032, 16'd14058, 16'd34309, 16'd39678, 16'd54985, 16'd62613, 16'd63233, 16'd46952, 16'd11874, 16'd53863, 16'd64927, 16'd59402, 16'd40671, 16'd38258});
	test_expansion(128'h697d0c087b7780cbfa06d4ee4c43183a, {16'd3547, 16'd1771, 16'd57778, 16'd11285, 16'd31423, 16'd20711, 16'd58334, 16'd14873, 16'd4388, 16'd11696, 16'd6476, 16'd16177, 16'd11090, 16'd62478, 16'd27997, 16'd5850, 16'd232, 16'd46901, 16'd36955, 16'd32455, 16'd64889, 16'd10823, 16'd34586, 16'd18040, 16'd63561, 16'd21662});
	test_expansion(128'he4502d919d1ae4c25af2fdf140738ee7, {16'd28406, 16'd8655, 16'd39983, 16'd32395, 16'd50757, 16'd15060, 16'd46795, 16'd44474, 16'd12446, 16'd52113, 16'd46851, 16'd8770, 16'd39829, 16'd40522, 16'd18580, 16'd17467, 16'd50261, 16'd23960, 16'd43810, 16'd33571, 16'd39800, 16'd39526, 16'd34328, 16'd23015, 16'd60240, 16'd1132});
	test_expansion(128'h0e55923cf5132e9981a8f7a62e2103c8, {16'd27719, 16'd49625, 16'd39623, 16'd20792, 16'd3115, 16'd38289, 16'd32539, 16'd35865, 16'd8879, 16'd60635, 16'd15597, 16'd21885, 16'd61179, 16'd54646, 16'd59499, 16'd12158, 16'd17595, 16'd55851, 16'd50256, 16'd20108, 16'd16122, 16'd10348, 16'd12641, 16'd31412, 16'd28280, 16'd24468});
	test_expansion(128'ha1abd47ff2937655fc8eacf355ff613e, {16'd13179, 16'd22409, 16'd9001, 16'd19112, 16'd64727, 16'd1820, 16'd59949, 16'd27334, 16'd65255, 16'd18767, 16'd10252, 16'd63580, 16'd27851, 16'd25942, 16'd32516, 16'd37068, 16'd33897, 16'd27930, 16'd57876, 16'd40720, 16'd49877, 16'd50917, 16'd13513, 16'd299, 16'd3967, 16'd64759});
	test_expansion(128'h0b2728ed141b58a869dcf2686ee60751, {16'd14821, 16'd28399, 16'd63776, 16'd7996, 16'd47715, 16'd20073, 16'd48345, 16'd42555, 16'd9761, 16'd11110, 16'd1214, 16'd61138, 16'd20366, 16'd22877, 16'd33696, 16'd51883, 16'd11638, 16'd3607, 16'd7433, 16'd55317, 16'd46680, 16'd4326, 16'd6276, 16'd18975, 16'd14305, 16'd57231});
	test_expansion(128'h7fa50c2bdf6daa510c347e4e37f7c65e, {16'd3834, 16'd22630, 16'd44253, 16'd62587, 16'd32880, 16'd35569, 16'd28153, 16'd43455, 16'd34536, 16'd20588, 16'd35906, 16'd2348, 16'd54250, 16'd61554, 16'd54135, 16'd7773, 16'd1562, 16'd7863, 16'd56792, 16'd5115, 16'd19734, 16'd49207, 16'd63780, 16'd48957, 16'd44073, 16'd17729});
	test_expansion(128'h0b1effbe9098c203a9aee73217cf00b8, {16'd14417, 16'd35735, 16'd11227, 16'd12714, 16'd60988, 16'd19359, 16'd6541, 16'd29189, 16'd26305, 16'd9909, 16'd57433, 16'd55421, 16'd9383, 16'd53268, 16'd2029, 16'd17056, 16'd2028, 16'd38061, 16'd17388, 16'd5629, 16'd63609, 16'd16304, 16'd27718, 16'd26620, 16'd21891, 16'd29190});
	test_expansion(128'hb9b220680c01311d297cb499105b9928, {16'd14901, 16'd31617, 16'd22123, 16'd64894, 16'd55166, 16'd43108, 16'd10487, 16'd44606, 16'd657, 16'd52995, 16'd12073, 16'd36024, 16'd36831, 16'd29390, 16'd11957, 16'd54840, 16'd14803, 16'd14539, 16'd60137, 16'd55322, 16'd64098, 16'd9371, 16'd23795, 16'd19372, 16'd21161, 16'd41287});
	test_expansion(128'h7ec45a286f3050e1f667798b58be1114, {16'd54817, 16'd33620, 16'd7200, 16'd46493, 16'd14370, 16'd23461, 16'd9797, 16'd35802, 16'd21693, 16'd39794, 16'd57177, 16'd19668, 16'd56686, 16'd4054, 16'd46781, 16'd32547, 16'd1201, 16'd33200, 16'd29326, 16'd13545, 16'd47967, 16'd60569, 16'd59039, 16'd22163, 16'd35286, 16'd44941});
	test_expansion(128'h5bb90d7c4c5e753db29ee9e9cc9b243e, {16'd57255, 16'd24164, 16'd57207, 16'd59113, 16'd41810, 16'd64188, 16'd16617, 16'd34370, 16'd32960, 16'd52793, 16'd15873, 16'd23086, 16'd63946, 16'd19986, 16'd52254, 16'd9298, 16'd30039, 16'd37742, 16'd34224, 16'd50424, 16'd62845, 16'd57912, 16'd23561, 16'd8689, 16'd61952, 16'd32988});
	test_expansion(128'h2c2e794d37dd63e31da972344e5b9de1, {16'd22807, 16'd28750, 16'd9548, 16'd22802, 16'd6747, 16'd50310, 16'd26991, 16'd61777, 16'd59388, 16'd2958, 16'd58081, 16'd39825, 16'd1380, 16'd12708, 16'd61111, 16'd4367, 16'd61354, 16'd11621, 16'd58741, 16'd29011, 16'd33048, 16'd49768, 16'd54062, 16'd33119, 16'd29618, 16'd54397});
	test_expansion(128'he71e01fd3de3ae51102a18681543d538, {16'd34684, 16'd4690, 16'd64732, 16'd8522, 16'd18150, 16'd3489, 16'd37890, 16'd28339, 16'd20815, 16'd4435, 16'd24745, 16'd4541, 16'd24566, 16'd35565, 16'd53287, 16'd34587, 16'd11449, 16'd1585, 16'd4822, 16'd18153, 16'd2693, 16'd25255, 16'd35260, 16'd52076, 16'd15617, 16'd18452});
	test_expansion(128'h69b479e89b5d637f05e2a3f0558dbd50, {16'd56171, 16'd45920, 16'd31219, 16'd54042, 16'd28857, 16'd57316, 16'd2203, 16'd53435, 16'd48775, 16'd55521, 16'd63239, 16'd13341, 16'd11805, 16'd40545, 16'd57322, 16'd8234, 16'd4735, 16'd17527, 16'd59346, 16'd29058, 16'd12249, 16'd716, 16'd53417, 16'd44193, 16'd63760, 16'd39080});
	test_expansion(128'h287b3d54403b1f83b48f2f92c0a4b8be, {16'd40346, 16'd64712, 16'd33383, 16'd14538, 16'd19763, 16'd47176, 16'd45148, 16'd43985, 16'd64406, 16'd44623, 16'd18794, 16'd26491, 16'd23792, 16'd12870, 16'd45364, 16'd63229, 16'd34283, 16'd34826, 16'd61874, 16'd27723, 16'd35836, 16'd62075, 16'd2384, 16'd8106, 16'd59603, 16'd22949});
	test_expansion(128'h8c952fbda1724aa8ebf1376453a175ce, {16'd65027, 16'd48713, 16'd12500, 16'd37126, 16'd14930, 16'd63140, 16'd3784, 16'd58479, 16'd61298, 16'd8130, 16'd53285, 16'd37957, 16'd8242, 16'd5667, 16'd14052, 16'd58212, 16'd17199, 16'd18271, 16'd32612, 16'd33875, 16'd15275, 16'd1835, 16'd34956, 16'd434, 16'd16667, 16'd28421});
	test_expansion(128'h452e9740a0d9c6b6326a4231c71a38a4, {16'd6483, 16'd54012, 16'd27892, 16'd26926, 16'd46166, 16'd12269, 16'd3395, 16'd2929, 16'd37909, 16'd27993, 16'd55991, 16'd56038, 16'd57301, 16'd39324, 16'd14040, 16'd34106, 16'd11437, 16'd18584, 16'd40284, 16'd30847, 16'd60164, 16'd2807, 16'd1541, 16'd38692, 16'd35993, 16'd64829});
	test_expansion(128'h61e88094b03345094b18a286f1848f3a, {16'd24118, 16'd38978, 16'd46566, 16'd16602, 16'd57198, 16'd11369, 16'd39376, 16'd12644, 16'd14337, 16'd11939, 16'd6146, 16'd20004, 16'd52028, 16'd16159, 16'd52068, 16'd12492, 16'd61852, 16'd49180, 16'd4334, 16'd45843, 16'd8715, 16'd30610, 16'd8324, 16'd54277, 16'd10472, 16'd25475});
	test_expansion(128'h7143a346a1430e1044529849d829ad8a, {16'd38222, 16'd30547, 16'd5916, 16'd2222, 16'd44718, 16'd25933, 16'd39827, 16'd53892, 16'd38699, 16'd30054, 16'd49639, 16'd26916, 16'd9219, 16'd52549, 16'd18835, 16'd35334, 16'd50376, 16'd33481, 16'd5008, 16'd53099, 16'd49635, 16'd53554, 16'd963, 16'd60733, 16'd2388, 16'd51408});
	test_expansion(128'h352ac78b80fc811fc29fa7651b34aa29, {16'd15302, 16'd29466, 16'd1084, 16'd19718, 16'd38561, 16'd52231, 16'd10706, 16'd7887, 16'd23136, 16'd29027, 16'd23994, 16'd35725, 16'd59363, 16'd58488, 16'd25052, 16'd44073, 16'd30551, 16'd34201, 16'd27543, 16'd14524, 16'd43143, 16'd57844, 16'd56555, 16'd14567, 16'd38119, 16'd42703});
	test_expansion(128'hce78b37548bb9eb3ac415aca0123afb1, {16'd12162, 16'd61932, 16'd16659, 16'd14862, 16'd4395, 16'd30847, 16'd2790, 16'd16258, 16'd36757, 16'd48629, 16'd39104, 16'd65231, 16'd49923, 16'd7415, 16'd11142, 16'd29396, 16'd37451, 16'd9470, 16'd54756, 16'd51030, 16'd24661, 16'd15565, 16'd49919, 16'd3651, 16'd24127, 16'd2732});
	test_expansion(128'hc795278ea501f3230a350aa067651f77, {16'd47239, 16'd4709, 16'd11729, 16'd49776, 16'd20655, 16'd9052, 16'd22119, 16'd4134, 16'd10497, 16'd27738, 16'd58805, 16'd12718, 16'd60676, 16'd34714, 16'd56390, 16'd61737, 16'd61725, 16'd13389, 16'd760, 16'd53384, 16'd17178, 16'd30124, 16'd20123, 16'd8705, 16'd24430, 16'd56869});
	test_expansion(128'h6f89a691a6265ec83e054f5df59cff2d, {16'd8493, 16'd25892, 16'd49418, 16'd8571, 16'd38155, 16'd54649, 16'd43843, 16'd10349, 16'd3047, 16'd25579, 16'd41634, 16'd61636, 16'd58381, 16'd5998, 16'd15835, 16'd6229, 16'd26506, 16'd13762, 16'd62659, 16'd691, 16'd39401, 16'd37942, 16'd47943, 16'd38831, 16'd56133, 16'd1380});
	test_expansion(128'h254e80f22152ba9a14b1a132b920edf8, {16'd50204, 16'd13893, 16'd9845, 16'd14145, 16'd1335, 16'd54791, 16'd35557, 16'd22936, 16'd62470, 16'd26685, 16'd11663, 16'd63253, 16'd34151, 16'd47991, 16'd44653, 16'd5984, 16'd44940, 16'd18764, 16'd6059, 16'd32447, 16'd44854, 16'd25786, 16'd54516, 16'd21680, 16'd4866, 16'd12506});
	test_expansion(128'h1c77e015b84a03f217f4819944e40b87, {16'd30457, 16'd5433, 16'd10266, 16'd10860, 16'd23575, 16'd9782, 16'd33764, 16'd26855, 16'd48839, 16'd60733, 16'd37562, 16'd44471, 16'd30514, 16'd51986, 16'd34233, 16'd1891, 16'd23183, 16'd19097, 16'd13109, 16'd65369, 16'd7430, 16'd26953, 16'd62194, 16'd13660, 16'd65507, 16'd55499});
	test_expansion(128'h8819c3baee829db227c70008bb6ee3fc, {16'd10492, 16'd41404, 16'd16976, 16'd30098, 16'd9207, 16'd58388, 16'd23102, 16'd61870, 16'd9693, 16'd52535, 16'd32493, 16'd24461, 16'd56623, 16'd49583, 16'd44700, 16'd23598, 16'd58267, 16'd46607, 16'd53389, 16'd9918, 16'd60522, 16'd8754, 16'd44232, 16'd10604, 16'd23481, 16'd33255});
	test_expansion(128'ha0cbea0ffe185e5165b66e47c7bf32e2, {16'd17595, 16'd2604, 16'd30795, 16'd57488, 16'd36686, 16'd20748, 16'd56936, 16'd31870, 16'd34672, 16'd19769, 16'd64390, 16'd11445, 16'd5860, 16'd51913, 16'd56112, 16'd50581, 16'd50959, 16'd55733, 16'd45100, 16'd56778, 16'd44362, 16'd50980, 16'd56408, 16'd3961, 16'd20221, 16'd44344});
	test_expansion(128'h6269cf0a8edf7902674528d895771271, {16'd13285, 16'd11481, 16'd8620, 16'd13290, 16'd23302, 16'd54455, 16'd32808, 16'd22374, 16'd19898, 16'd49899, 16'd8831, 16'd49831, 16'd16302, 16'd33835, 16'd27001, 16'd6472, 16'd63663, 16'd9099, 16'd28704, 16'd63105, 16'd13771, 16'd19435, 16'd55074, 16'd15565, 16'd31921, 16'd48800});
	test_expansion(128'h2b6ae8ca8973371d27e572c9992f1675, {16'd48242, 16'd8348, 16'd28139, 16'd13535, 16'd54324, 16'd23438, 16'd48401, 16'd39102, 16'd55121, 16'd35672, 16'd64474, 16'd3812, 16'd55490, 16'd55690, 16'd51871, 16'd35582, 16'd49791, 16'd39165, 16'd39917, 16'd14818, 16'd36532, 16'd7235, 16'd51365, 16'd54176, 16'd37823, 16'd43989});
	test_expansion(128'h6c709ce79fe810ba4c0cbcb9c71f503a, {16'd25600, 16'd1473, 16'd19344, 16'd11833, 16'd31707, 16'd590, 16'd54057, 16'd62864, 16'd20454, 16'd21732, 16'd37792, 16'd16762, 16'd45531, 16'd38525, 16'd57392, 16'd28096, 16'd61565, 16'd29779, 16'd532, 16'd24353, 16'd36158, 16'd36017, 16'd29204, 16'd8845, 16'd54513, 16'd32511});
	test_expansion(128'h430669e10f9e9f366f90ececb02debac, {16'd43224, 16'd16181, 16'd25885, 16'd13128, 16'd29176, 16'd46851, 16'd62036, 16'd53912, 16'd39484, 16'd39277, 16'd11431, 16'd40601, 16'd282, 16'd27409, 16'd51260, 16'd23808, 16'd64601, 16'd48332, 16'd21997, 16'd34224, 16'd14841, 16'd44825, 16'd2075, 16'd52928, 16'd53986, 16'd12464});
	test_expansion(128'he2045e07012d33f84677d1f3e5a843c4, {16'd31381, 16'd20401, 16'd53780, 16'd29739, 16'd978, 16'd43201, 16'd55950, 16'd41418, 16'd51758, 16'd55078, 16'd56398, 16'd41011, 16'd11495, 16'd20442, 16'd17554, 16'd54321, 16'd64092, 16'd876, 16'd31872, 16'd52224, 16'd29397, 16'd17010, 16'd60911, 16'd42928, 16'd6594, 16'd64165});
	test_expansion(128'hec2ed10f9c4ebad4cf43dc8191e6b765, {16'd34179, 16'd61049, 16'd59817, 16'd4970, 16'd55930, 16'd41715, 16'd26501, 16'd21993, 16'd2349, 16'd1658, 16'd41601, 16'd1806, 16'd13728, 16'd13572, 16'd55818, 16'd55045, 16'd12755, 16'd35271, 16'd55580, 16'd55368, 16'd13851, 16'd31787, 16'd54151, 16'd51621, 16'd45269, 16'd60217});
	test_expansion(128'hd19426766162b3ebada037ee067a8542, {16'd59989, 16'd15697, 16'd30816, 16'd52896, 16'd1683, 16'd35386, 16'd47521, 16'd12750, 16'd30193, 16'd23547, 16'd4055, 16'd37233, 16'd15763, 16'd5070, 16'd57613, 16'd46204, 16'd33771, 16'd48386, 16'd57951, 16'd25874, 16'd36071, 16'd14579, 16'd64549, 16'd47629, 16'd52490, 16'd31223});
	test_expansion(128'hf22add661642865abaa03ae8aeaf5f60, {16'd8752, 16'd4206, 16'd25837, 16'd10044, 16'd52977, 16'd8253, 16'd34433, 16'd34513, 16'd3690, 16'd30141, 16'd24811, 16'd54716, 16'd22736, 16'd51792, 16'd57741, 16'd24530, 16'd62875, 16'd18801, 16'd64170, 16'd37955, 16'd27966, 16'd16914, 16'd52389, 16'd45364, 16'd54854, 16'd23763});
	test_expansion(128'haaeb8a08e202ea54635a0c4b5be7535c, {16'd16975, 16'd10561, 16'd51026, 16'd35099, 16'd29153, 16'd18361, 16'd32727, 16'd48878, 16'd29391, 16'd39849, 16'd19582, 16'd20030, 16'd36274, 16'd30938, 16'd48215, 16'd56777, 16'd49003, 16'd59684, 16'd33008, 16'd49010, 16'd11477, 16'd33455, 16'd64949, 16'd12968, 16'd6851, 16'd10014});
	test_expansion(128'h0c64a1f07fcd730183c94bb8c596fa5f, {16'd14196, 16'd49076, 16'd30160, 16'd35758, 16'd36953, 16'd3550, 16'd49488, 16'd56219, 16'd31979, 16'd32211, 16'd31452, 16'd29172, 16'd15253, 16'd42664, 16'd31058, 16'd6533, 16'd13361, 16'd49877, 16'd40564, 16'd44980, 16'd35787, 16'd59014, 16'd13760, 16'd63108, 16'd7696, 16'd12434});
	test_expansion(128'h39dcd938089c2dd414c69e3fa19f0f2f, {16'd49455, 16'd62548, 16'd32585, 16'd14081, 16'd30746, 16'd47384, 16'd58373, 16'd11274, 16'd11960, 16'd31951, 16'd10365, 16'd30024, 16'd48671, 16'd23400, 16'd2004, 16'd11750, 16'd30790, 16'd27314, 16'd23825, 16'd18535, 16'd28066, 16'd51106, 16'd44487, 16'd11923, 16'd11248, 16'd32475});
	test_expansion(128'h69fb0835598f1e41bea63cbbad8e7aee, {16'd56091, 16'd16407, 16'd30017, 16'd43266, 16'd33026, 16'd2382, 16'd11411, 16'd15285, 16'd5186, 16'd33069, 16'd50654, 16'd23752, 16'd17362, 16'd734, 16'd18415, 16'd30894, 16'd28372, 16'd28529, 16'd39117, 16'd57318, 16'd55530, 16'd53006, 16'd47492, 16'd44859, 16'd42342, 16'd46857});
	test_expansion(128'hb198d9725a6ae0af05ed4b51c62633a8, {16'd17929, 16'd25536, 16'd29583, 16'd19481, 16'd46875, 16'd6274, 16'd56074, 16'd62661, 16'd49802, 16'd62285, 16'd23738, 16'd63539, 16'd12813, 16'd43546, 16'd24184, 16'd6266, 16'd16640, 16'd45935, 16'd49687, 16'd5129, 16'd4447, 16'd12914, 16'd45775, 16'd33838, 16'd56490, 16'd6470});
	test_expansion(128'he27b7560a9ed2378bce6481cf806eebf, {16'd50547, 16'd12561, 16'd26964, 16'd29719, 16'd53808, 16'd46559, 16'd28246, 16'd3522, 16'd6741, 16'd14173, 16'd32818, 16'd10131, 16'd1111, 16'd65242, 16'd64836, 16'd29010, 16'd20862, 16'd47974, 16'd27778, 16'd52406, 16'd8865, 16'd38111, 16'd49841, 16'd19044, 16'd28155, 16'd61863});
	test_expansion(128'hd8d7867a54e9355752add3effe98dcd1, {16'd25495, 16'd1935, 16'd81, 16'd45351, 16'd58645, 16'd29213, 16'd27145, 16'd12049, 16'd35505, 16'd38866, 16'd36361, 16'd37593, 16'd21287, 16'd14720, 16'd58791, 16'd32494, 16'd62987, 16'd15710, 16'd26341, 16'd29515, 16'd42432, 16'd7735, 16'd9154, 16'd38202, 16'd35722, 16'd14986});
	test_expansion(128'hec49961dbc38fa0d0dc07c2d16f3a31e, {16'd7934, 16'd47832, 16'd56168, 16'd27287, 16'd20538, 16'd62802, 16'd30245, 16'd30361, 16'd48447, 16'd5917, 16'd65284, 16'd27587, 16'd43311, 16'd30629, 16'd24792, 16'd23332, 16'd28710, 16'd46068, 16'd44440, 16'd12467, 16'd38407, 16'd3887, 16'd26258, 16'd33000, 16'd35409, 16'd55245});
	test_expansion(128'he88ccf7c2404bb23e4bf6d0a6c0b362f, {16'd62487, 16'd51072, 16'd20275, 16'd42475, 16'd27916, 16'd44020, 16'd52589, 16'd24735, 16'd64946, 16'd52654, 16'd46801, 16'd4166, 16'd39523, 16'd50548, 16'd38886, 16'd64764, 16'd7942, 16'd35108, 16'd60174, 16'd50440, 16'd30650, 16'd22886, 16'd12019, 16'd33116, 16'd61783, 16'd18299});
	test_expansion(128'h02fc35641d7f640343747c893247cb88, {16'd61449, 16'd17856, 16'd40872, 16'd59196, 16'd15884, 16'd22457, 16'd52574, 16'd62920, 16'd28376, 16'd51187, 16'd48448, 16'd58072, 16'd10141, 16'd12112, 16'd57910, 16'd23789, 16'd42921, 16'd14057, 16'd25554, 16'd24318, 16'd4326, 16'd59856, 16'd25623, 16'd46051, 16'd16955, 16'd32043});
	test_expansion(128'h92113994745a341d146c868353f95b67, {16'd44902, 16'd60259, 16'd45835, 16'd38085, 16'd5759, 16'd22040, 16'd14057, 16'd671, 16'd56300, 16'd18166, 16'd20853, 16'd62915, 16'd11223, 16'd21892, 16'd50769, 16'd54121, 16'd3478, 16'd914, 16'd58758, 16'd56965, 16'd780, 16'd4259, 16'd27695, 16'd38955, 16'd35055, 16'd15443});
	test_expansion(128'h9c2cb1dd4b04c17219fa30542c2bf960, {16'd14304, 16'd21790, 16'd58149, 16'd11713, 16'd45880, 16'd62500, 16'd53009, 16'd6732, 16'd28174, 16'd48210, 16'd32538, 16'd40835, 16'd36346, 16'd54990, 16'd9511, 16'd28546, 16'd60535, 16'd35830, 16'd17856, 16'd63460, 16'd37374, 16'd17628, 16'd11201, 16'd25556, 16'd55400, 16'd32007});
	test_expansion(128'h714ae7a18db2511c2f6282b913e51b80, {16'd39761, 16'd30711, 16'd31231, 16'd20998, 16'd55821, 16'd42243, 16'd36299, 16'd29178, 16'd25610, 16'd23443, 16'd37261, 16'd30274, 16'd18889, 16'd56538, 16'd38080, 16'd44697, 16'd48085, 16'd55664, 16'd7213, 16'd2941, 16'd64826, 16'd53554, 16'd63386, 16'd2985, 16'd64007, 16'd18223});
	test_expansion(128'hf3da634ce57f0b40656a2a18b0916d8d, {16'd37683, 16'd1052, 16'd35233, 16'd17382, 16'd7126, 16'd40518, 16'd27407, 16'd8968, 16'd22370, 16'd9655, 16'd60410, 16'd38780, 16'd1621, 16'd15443, 16'd61043, 16'd6036, 16'd6976, 16'd16851, 16'd25026, 16'd60499, 16'd42603, 16'd6709, 16'd6198, 16'd1377, 16'd38870, 16'd25764});
	test_expansion(128'h76630b250b80ae3acefd2ad447bbc0ff, {16'd38709, 16'd21880, 16'd7990, 16'd63770, 16'd27558, 16'd22745, 16'd45734, 16'd44591, 16'd6939, 16'd12700, 16'd20676, 16'd28190, 16'd20784, 16'd39803, 16'd3443, 16'd47624, 16'd46293, 16'd62600, 16'd20171, 16'd20767, 16'd53147, 16'd47511, 16'd56254, 16'd47011, 16'd46751, 16'd3248});
	test_expansion(128'he4c2d09187dcacf16c6d754d98434640, {16'd20666, 16'd36852, 16'd20549, 16'd35212, 16'd55959, 16'd19488, 16'd59923, 16'd20532, 16'd49568, 16'd9809, 16'd53414, 16'd3377, 16'd60172, 16'd60791, 16'd2098, 16'd62849, 16'd5569, 16'd23440, 16'd36956, 16'd3188, 16'd53764, 16'd27329, 16'd53890, 16'd60476, 16'd63301, 16'd32025});
	test_expansion(128'h5c4271339a23d406e37998b6580faf77, {16'd21735, 16'd5810, 16'd49312, 16'd59770, 16'd38901, 16'd24291, 16'd50923, 16'd1399, 16'd35091, 16'd27038, 16'd26319, 16'd57950, 16'd14595, 16'd51571, 16'd4845, 16'd19572, 16'd60231, 16'd56812, 16'd57, 16'd60128, 16'd7894, 16'd39582, 16'd48172, 16'd13756, 16'd60429, 16'd8518});
	test_expansion(128'h93289144a9cd071aa7243efe8e51a755, {16'd41430, 16'd36122, 16'd59461, 16'd12280, 16'd40009, 16'd9882, 16'd33605, 16'd54004, 16'd64190, 16'd10053, 16'd23458, 16'd21897, 16'd13124, 16'd12912, 16'd29997, 16'd13022, 16'd8001, 16'd46029, 16'd36276, 16'd19359, 16'd16530, 16'd43078, 16'd13541, 16'd53749, 16'd27887, 16'd61635});
	test_expansion(128'hf5b791273b49486046c9a83bdf00a697, {16'd57749, 16'd13366, 16'd17482, 16'd26077, 16'd15287, 16'd60819, 16'd53890, 16'd9672, 16'd49421, 16'd54529, 16'd18348, 16'd65215, 16'd32161, 16'd21159, 16'd16963, 16'd13369, 16'd52138, 16'd29325, 16'd9412, 16'd34971, 16'd56308, 16'd53611, 16'd57824, 16'd60552, 16'd17105, 16'd3545});
	test_expansion(128'h952ead865e5fd179b39bacd9ac5c9dc3, {16'd41692, 16'd46595, 16'd59658, 16'd27425, 16'd39542, 16'd59197, 16'd22462, 16'd24794, 16'd54007, 16'd52051, 16'd37489, 16'd56675, 16'd35712, 16'd57124, 16'd1834, 16'd32456, 16'd37587, 16'd32273, 16'd4799, 16'd3209, 16'd13043, 16'd52612, 16'd21734, 16'd42821, 16'd14328, 16'd20727});
	test_expansion(128'hff00cb4e46916fa6ca7c788478250332, {16'd22083, 16'd63441, 16'd30488, 16'd42915, 16'd60478, 16'd21132, 16'd13189, 16'd25321, 16'd15077, 16'd411, 16'd17196, 16'd49533, 16'd7137, 16'd65054, 16'd8009, 16'd18257, 16'd39521, 16'd10386, 16'd6256, 16'd20907, 16'd4153, 16'd65456, 16'd54150, 16'd45400, 16'd8335, 16'd49961});
	test_expansion(128'h1bac9f29d2fdbac94e2e6f4aedac2029, {16'd4750, 16'd1185, 16'd31814, 16'd54231, 16'd20384, 16'd55344, 16'd37130, 16'd63193, 16'd24051, 16'd42934, 16'd7050, 16'd17763, 16'd40196, 16'd41594, 16'd358, 16'd33426, 16'd13860, 16'd42337, 16'd47122, 16'd20981, 16'd10495, 16'd29057, 16'd50623, 16'd32552, 16'd51133, 16'd34483});
	test_expansion(128'hc637367f2b5b9cc44e2cd5e280addb6f, {16'd5559, 16'd9171, 16'd33256, 16'd4390, 16'd38334, 16'd19142, 16'd45375, 16'd45295, 16'd10930, 16'd39641, 16'd55294, 16'd44786, 16'd986, 16'd25389, 16'd51655, 16'd63827, 16'd32819, 16'd44060, 16'd64416, 16'd36956, 16'd22407, 16'd45319, 16'd48074, 16'd30102, 16'd17463, 16'd36323});
	test_expansion(128'hb2b00e2281b5c04f23598e1004eea948, {16'd52755, 16'd60405, 16'd8659, 16'd32116, 16'd19669, 16'd63652, 16'd15613, 16'd14837, 16'd10943, 16'd35462, 16'd56726, 16'd45370, 16'd18643, 16'd8556, 16'd52819, 16'd32457, 16'd27260, 16'd56113, 16'd32664, 16'd39034, 16'd2271, 16'd64102, 16'd43779, 16'd11234, 16'd30942, 16'd31365});
	test_expansion(128'h58e46ceab6ffaf1fbe12f0a65daaccd9, {16'd3525, 16'd27859, 16'd50366, 16'd35225, 16'd41765, 16'd37717, 16'd1736, 16'd62718, 16'd7086, 16'd15890, 16'd19150, 16'd48243, 16'd37797, 16'd33428, 16'd57776, 16'd7196, 16'd18773, 16'd54573, 16'd49732, 16'd23998, 16'd63186, 16'd47035, 16'd52455, 16'd25279, 16'd54945, 16'd15953});
	test_expansion(128'h68a2d6f2c8ad3a3ee0765a120f04aa93, {16'd59939, 16'd25474, 16'd26683, 16'd46797, 16'd49750, 16'd61005, 16'd64391, 16'd35196, 16'd55999, 16'd39142, 16'd10901, 16'd7763, 16'd4543, 16'd30899, 16'd28363, 16'd10821, 16'd9942, 16'd2123, 16'd18765, 16'd20573, 16'd28749, 16'd12240, 16'd46394, 16'd19797, 16'd60635, 16'd61466});
	test_expansion(128'h9732f00ef8630c8375a1408a4d36da11, {16'd48478, 16'd41936, 16'd22045, 16'd64603, 16'd17515, 16'd52249, 16'd15759, 16'd44866, 16'd9056, 16'd33705, 16'd26748, 16'd28777, 16'd43901, 16'd39572, 16'd5157, 16'd59891, 16'd57406, 16'd41096, 16'd35646, 16'd50343, 16'd30517, 16'd32730, 16'd16768, 16'd64898, 16'd40014, 16'd7294});
	test_expansion(128'hc2dd01be2b4fb7d0f2b9c78d7b378bb3, {16'd59357, 16'd29415, 16'd2665, 16'd27441, 16'd47125, 16'd11721, 16'd12476, 16'd10991, 16'd8922, 16'd57713, 16'd5364, 16'd48229, 16'd63546, 16'd22863, 16'd38489, 16'd7102, 16'd29429, 16'd50501, 16'd53583, 16'd31741, 16'd32793, 16'd33392, 16'd64421, 16'd56118, 16'd27378, 16'd32538});
	test_expansion(128'hbf02718665ec0aeb640004c9b25c76e5, {16'd24151, 16'd49416, 16'd15897, 16'd8684, 16'd19960, 16'd48326, 16'd49733, 16'd8896, 16'd56607, 16'd37513, 16'd16953, 16'd12397, 16'd44648, 16'd58978, 16'd33181, 16'd51669, 16'd42977, 16'd26152, 16'd61302, 16'd42584, 16'd65048, 16'd48364, 16'd13583, 16'd43402, 16'd53531, 16'd63381});
	test_expansion(128'h893a80a553066ac6def9adc60164a6c2, {16'd43377, 16'd57848, 16'd54695, 16'd33127, 16'd9417, 16'd38228, 16'd7860, 16'd9232, 16'd9444, 16'd12082, 16'd34031, 16'd28705, 16'd3089, 16'd48945, 16'd49849, 16'd55712, 16'd60904, 16'd47241, 16'd36998, 16'd22153, 16'd5842, 16'd40662, 16'd42119, 16'd40995, 16'd5484, 16'd16502});
	test_expansion(128'ha96b24db079530f538fe7f856c0063da, {16'd30100, 16'd62948, 16'd65052, 16'd36711, 16'd43777, 16'd17239, 16'd17479, 16'd39011, 16'd11131, 16'd3499, 16'd9458, 16'd13530, 16'd13655, 16'd11978, 16'd38822, 16'd45393, 16'd3041, 16'd3050, 16'd38555, 16'd45819, 16'd35844, 16'd36806, 16'd29011, 16'd51430, 16'd3705, 16'd62291});
	test_expansion(128'h1e6d4e5f2248aaa44e32d12249f6456f, {16'd40307, 16'd45429, 16'd54222, 16'd32832, 16'd35253, 16'd39592, 16'd6774, 16'd42558, 16'd4342, 16'd38550, 16'd50887, 16'd20742, 16'd34995, 16'd24997, 16'd39411, 16'd34476, 16'd62671, 16'd58102, 16'd2858, 16'd9524, 16'd9919, 16'd28409, 16'd6567, 16'd22793, 16'd26199, 16'd22327});
	test_expansion(128'h893e1b8628210fe18e0ce0702e156677, {16'd48261, 16'd53721, 16'd4379, 16'd15962, 16'd25660, 16'd25510, 16'd7970, 16'd45879, 16'd23412, 16'd12042, 16'd7540, 16'd51700, 16'd4359, 16'd3376, 16'd2395, 16'd45658, 16'd13746, 16'd46212, 16'd55178, 16'd56607, 16'd60662, 16'd23408, 16'd57274, 16'd6457, 16'd37992, 16'd23844});
	test_expansion(128'hf407a579ef6842c5f8acac88ca872bd5, {16'd5104, 16'd64587, 16'd65414, 16'd15254, 16'd44641, 16'd14389, 16'd4407, 16'd23163, 16'd9953, 16'd33236, 16'd32776, 16'd39721, 16'd41738, 16'd7335, 16'd33542, 16'd6846, 16'd44382, 16'd3418, 16'd63700, 16'd61248, 16'd49902, 16'd56605, 16'd62886, 16'd34484, 16'd65418, 16'd60326});
	test_expansion(128'hc2908a7d49da4fa4ba4c6518f6243fb2, {16'd16226, 16'd43252, 16'd62758, 16'd27510, 16'd18753, 16'd34649, 16'd22783, 16'd60288, 16'd65472, 16'd4246, 16'd54914, 16'd24654, 16'd19242, 16'd51667, 16'd37875, 16'd65520, 16'd28473, 16'd55143, 16'd21504, 16'd45101, 16'd40273, 16'd5600, 16'd46372, 16'd64896, 16'd39859, 16'd16752});
	test_expansion(128'h554bdd0831e189e6b29bb0e6a3d302ca, {16'd60012, 16'd39583, 16'd8602, 16'd64294, 16'd25661, 16'd47259, 16'd1934, 16'd52507, 16'd43922, 16'd59698, 16'd31671, 16'd62141, 16'd48638, 16'd16862, 16'd62613, 16'd57478, 16'd41328, 16'd9748, 16'd46395, 16'd7092, 16'd6547, 16'd14236, 16'd4070, 16'd64388, 16'd4890, 16'd46647});
	test_expansion(128'h2dc3ddcebc25fc1fbc96bd22fd6b496a, {16'd18295, 16'd49122, 16'd7394, 16'd29421, 16'd41957, 16'd60124, 16'd37592, 16'd11679, 16'd65515, 16'd18039, 16'd43122, 16'd11828, 16'd9133, 16'd34992, 16'd7084, 16'd37116, 16'd1799, 16'd60645, 16'd13461, 16'd12620, 16'd60671, 16'd36703, 16'd29884, 16'd15783, 16'd46951, 16'd60281});
	test_expansion(128'hc8a1926aa903ea9209c8ebccc12c38f1, {16'd32503, 16'd47386, 16'd20275, 16'd55659, 16'd9677, 16'd49335, 16'd25336, 16'd4627, 16'd10477, 16'd64922, 16'd33690, 16'd25084, 16'd36432, 16'd49566, 16'd38110, 16'd891, 16'd18205, 16'd46680, 16'd19486, 16'd36337, 16'd28511, 16'd37786, 16'd8011, 16'd39737, 16'd17736, 16'd55485});
	test_expansion(128'h1243364d570756633f0b50ea7fbc05f8, {16'd24559, 16'd10105, 16'd24360, 16'd43469, 16'd42020, 16'd60159, 16'd1811, 16'd5609, 16'd43743, 16'd21583, 16'd42621, 16'd21063, 16'd52827, 16'd55816, 16'd1112, 16'd41968, 16'd62336, 16'd19819, 16'd13332, 16'd15868, 16'd43601, 16'd44793, 16'd3085, 16'd33658, 16'd13271, 16'd36791});
	test_expansion(128'hbdda9789a595045630372f7613bcd440, {16'd27681, 16'd44278, 16'd8761, 16'd49622, 16'd22951, 16'd48861, 16'd63590, 16'd63086, 16'd57861, 16'd10535, 16'd7312, 16'd8743, 16'd26460, 16'd21633, 16'd26267, 16'd52524, 16'd34586, 16'd47338, 16'd43817, 16'd2213, 16'd19298, 16'd36392, 16'd46263, 16'd12422, 16'd34490, 16'd32941});
	test_expansion(128'hd06d39d2ffef977fa6cdc524cabc0695, {16'd22617, 16'd33790, 16'd62819, 16'd49279, 16'd31211, 16'd24179, 16'd53409, 16'd1886, 16'd7813, 16'd39565, 16'd62204, 16'd29625, 16'd17872, 16'd951, 16'd55547, 16'd6808, 16'd23442, 16'd26784, 16'd3421, 16'd6523, 16'd37911, 16'd45510, 16'd55048, 16'd10684, 16'd48525, 16'd27878});
	test_expansion(128'h8225adc76b27852f1e9d7f61449f90b1, {16'd56536, 16'd25232, 16'd14089, 16'd15220, 16'd17448, 16'd44143, 16'd19547, 16'd3534, 16'd60819, 16'd25195, 16'd63143, 16'd509, 16'd14754, 16'd40985, 16'd37483, 16'd61773, 16'd12528, 16'd53756, 16'd24816, 16'd41506, 16'd52607, 16'd32897, 16'd23175, 16'd64817, 16'd45603, 16'd59010});
	test_expansion(128'h39e3ab8d226054d4d8d3e5882d48c2d6, {16'd37532, 16'd45771, 16'd48849, 16'd21338, 16'd13867, 16'd57252, 16'd20473, 16'd38634, 16'd17876, 16'd9659, 16'd4841, 16'd35439, 16'd57052, 16'd50073, 16'd27861, 16'd12543, 16'd1354, 16'd29144, 16'd16782, 16'd9355, 16'd53059, 16'd44145, 16'd11810, 16'd24173, 16'd43497, 16'd65036});
	test_expansion(128'ha2427cb43924d40f3672cf1d952231fc, {16'd48412, 16'd57629, 16'd36132, 16'd47121, 16'd28640, 16'd48321, 16'd46061, 16'd61897, 16'd9578, 16'd22875, 16'd55845, 16'd33380, 16'd31579, 16'd54530, 16'd4702, 16'd51423, 16'd60097, 16'd3169, 16'd9185, 16'd53069, 16'd54601, 16'd50907, 16'd5779, 16'd21990, 16'd6134, 16'd53366});
	test_expansion(128'h83652a2d6b321ed76e8f33457e966607, {16'd37041, 16'd6581, 16'd55696, 16'd60311, 16'd22348, 16'd30905, 16'd20976, 16'd53175, 16'd50519, 16'd17145, 16'd65505, 16'd42755, 16'd49744, 16'd59279, 16'd15043, 16'd21966, 16'd49940, 16'd51760, 16'd19052, 16'd14998, 16'd34150, 16'd24227, 16'd39831, 16'd1314, 16'd1901, 16'd5396});
	test_expansion(128'h0fff2ee30a3138d7284a4309334f1f57, {16'd12103, 16'd63638, 16'd1300, 16'd60007, 16'd48488, 16'd32470, 16'd54456, 16'd50993, 16'd48620, 16'd64193, 16'd17400, 16'd29771, 16'd5453, 16'd44954, 16'd55491, 16'd40982, 16'd41992, 16'd47076, 16'd31145, 16'd9458, 16'd49976, 16'd24521, 16'd17261, 16'd61011, 16'd10445, 16'd33046});
	test_expansion(128'h9dfef86882dba25f0f95fbdbde064786, {16'd47675, 16'd49494, 16'd28205, 16'd40375, 16'd3658, 16'd56541, 16'd39790, 16'd55563, 16'd23862, 16'd3949, 16'd4851, 16'd7435, 16'd47211, 16'd51072, 16'd16410, 16'd17183, 16'd44533, 16'd27311, 16'd51686, 16'd53157, 16'd32378, 16'd52466, 16'd39950, 16'd51354, 16'd44302, 16'd33437});
	test_expansion(128'h2fc4863155809209b9a000bdfa5faebd, {16'd64288, 16'd38969, 16'd39971, 16'd27637, 16'd21033, 16'd27910, 16'd60497, 16'd25718, 16'd20959, 16'd38, 16'd32089, 16'd54900, 16'd44520, 16'd32284, 16'd42350, 16'd18736, 16'd47424, 16'd4377, 16'd33096, 16'd18275, 16'd53992, 16'd22708, 16'd16219, 16'd21924, 16'd22516, 16'd17919});
	test_expansion(128'h31485de4167155aa53d4a234fc36c9b6, {16'd60498, 16'd14452, 16'd36438, 16'd34763, 16'd2817, 16'd32851, 16'd43704, 16'd36042, 16'd36643, 16'd36074, 16'd2198, 16'd38188, 16'd53434, 16'd24977, 16'd8416, 16'd26890, 16'd42975, 16'd8507, 16'd26271, 16'd23752, 16'd49947, 16'd54178, 16'd17525, 16'd1926, 16'd47034, 16'd12236});
	test_expansion(128'h93600fd502985d1142092133e73f29f0, {16'd20326, 16'd26426, 16'd34004, 16'd32305, 16'd42446, 16'd28509, 16'd20105, 16'd56871, 16'd33411, 16'd59701, 16'd20677, 16'd24190, 16'd9447, 16'd43781, 16'd41282, 16'd34043, 16'd44964, 16'd57589, 16'd13574, 16'd1751, 16'd3316, 16'd54616, 16'd21637, 16'd62999, 16'd37008, 16'd7729});
	test_expansion(128'h72137d60115b5eabd2c0c38a3d46dda8, {16'd49444, 16'd45636, 16'd6453, 16'd64627, 16'd28313, 16'd25759, 16'd28672, 16'd8114, 16'd7663, 16'd13237, 16'd32148, 16'd8959, 16'd40385, 16'd61182, 16'd13335, 16'd23110, 16'd53655, 16'd42044, 16'd25026, 16'd52311, 16'd41101, 16'd19358, 16'd19277, 16'd52112, 16'd62885, 16'd27990});
	test_expansion(128'h07d87cba1b7d7d3b2f90108f4488d97e, {16'd45328, 16'd29317, 16'd56847, 16'd55838, 16'd34156, 16'd54707, 16'd33374, 16'd47062, 16'd26692, 16'd35902, 16'd15626, 16'd25234, 16'd38446, 16'd50593, 16'd44046, 16'd1472, 16'd28354, 16'd38778, 16'd23697, 16'd25516, 16'd11198, 16'd42037, 16'd15126, 16'd19979, 16'd45546, 16'd15185});
	test_expansion(128'h92acaa008694aac3bcde7855c58544ae, {16'd23402, 16'd16238, 16'd57630, 16'd54808, 16'd29694, 16'd63747, 16'd37231, 16'd48781, 16'd1504, 16'd55543, 16'd30919, 16'd62013, 16'd39808, 16'd9540, 16'd47180, 16'd45366, 16'd2046, 16'd44631, 16'd55844, 16'd5978, 16'd29233, 16'd7708, 16'd11807, 16'd62779, 16'd57105, 16'd59744});
	test_expansion(128'h6d9685e84ea52aebfddb0e63a4ead0cd, {16'd10763, 16'd62647, 16'd26847, 16'd14847, 16'd18458, 16'd17675, 16'd18582, 16'd62439, 16'd2444, 16'd55860, 16'd21696, 16'd41166, 16'd46547, 16'd33895, 16'd8445, 16'd9369, 16'd49164, 16'd46521, 16'd55811, 16'd11754, 16'd44680, 16'd58880, 16'd35380, 16'd56435, 16'd44358, 16'd15316});
	test_expansion(128'hccaaf3a3f713d75f6b6ea2a1037cde75, {16'd2278, 16'd39416, 16'd2057, 16'd30895, 16'd32936, 16'd6497, 16'd56147, 16'd54769, 16'd28179, 16'd5436, 16'd18448, 16'd9131, 16'd33287, 16'd38522, 16'd55720, 16'd2528, 16'd32942, 16'd15845, 16'd60509, 16'd45208, 16'd58593, 16'd39190, 16'd45113, 16'd18682, 16'd10289, 16'd10565});
	test_expansion(128'ha5a36b8a26c7dfb7f8066be48ef70c89, {16'd4668, 16'd37566, 16'd23177, 16'd21962, 16'd59634, 16'd4485, 16'd38321, 16'd46381, 16'd10872, 16'd44788, 16'd29748, 16'd41334, 16'd21469, 16'd21057, 16'd58930, 16'd23354, 16'd59299, 16'd41890, 16'd27073, 16'd9364, 16'd54496, 16'd53840, 16'd51039, 16'd51446, 16'd58836, 16'd16267});
	test_expansion(128'h661b947a42db02cc2afb6271fae9ae11, {16'd2457, 16'd63612, 16'd46465, 16'd42436, 16'd19743, 16'd17298, 16'd11003, 16'd64725, 16'd11740, 16'd14822, 16'd49839, 16'd5145, 16'd21737, 16'd27136, 16'd10210, 16'd57067, 16'd46584, 16'd16408, 16'd22847, 16'd32547, 16'd9758, 16'd49674, 16'd27395, 16'd21278, 16'd23456, 16'd3363});
	test_expansion(128'h674783fd349a4767b50c980f195b53dc, {16'd41772, 16'd54736, 16'd13387, 16'd50542, 16'd19835, 16'd61039, 16'd4681, 16'd43551, 16'd47233, 16'd38820, 16'd47978, 16'd32047, 16'd746, 16'd35230, 16'd8471, 16'd33407, 16'd15197, 16'd59444, 16'd15529, 16'd14477, 16'd40857, 16'd48097, 16'd25540, 16'd52534, 16'd9556, 16'd15542});
	test_expansion(128'he9eae751d9406ad5d5abde58fad9ac41, {16'd62015, 16'd35567, 16'd28496, 16'd2005, 16'd9371, 16'd36927, 16'd45211, 16'd10459, 16'd16184, 16'd34731, 16'd40602, 16'd61215, 16'd17000, 16'd14080, 16'd23642, 16'd4740, 16'd62057, 16'd36084, 16'd36780, 16'd22582, 16'd49711, 16'd46200, 16'd10170, 16'd52999, 16'd53732, 16'd33330});
	test_expansion(128'hcfd60c45668e853e52c306d00064f39c, {16'd65128, 16'd57150, 16'd19052, 16'd28206, 16'd30914, 16'd27443, 16'd38085, 16'd39906, 16'd30907, 16'd51799, 16'd49495, 16'd19439, 16'd45709, 16'd31660, 16'd58620, 16'd6218, 16'd60374, 16'd5903, 16'd11355, 16'd47401, 16'd54607, 16'd60978, 16'd13171, 16'd45676, 16'd15826, 16'd4764});
	test_expansion(128'hae6f0e549854d9d1dbcde8a1d9de3ff8, {16'd30225, 16'd49775, 16'd37912, 16'd12454, 16'd35201, 16'd29175, 16'd9104, 16'd29510, 16'd55574, 16'd22629, 16'd57429, 16'd1133, 16'd45987, 16'd60315, 16'd23416, 16'd43800, 16'd16715, 16'd62120, 16'd61048, 16'd8596, 16'd11802, 16'd62673, 16'd20436, 16'd64379, 16'd12999, 16'd60738});
	test_expansion(128'hb4f0f13d411b5baefcc5959a60d4115e, {16'd53547, 16'd64163, 16'd61733, 16'd30559, 16'd8728, 16'd23790, 16'd39755, 16'd26712, 16'd5741, 16'd29329, 16'd9, 16'd10288, 16'd3092, 16'd48857, 16'd45739, 16'd54215, 16'd9371, 16'd42095, 16'd44802, 16'd58741, 16'd58087, 16'd13548, 16'd11337, 16'd41052, 16'd2431, 16'd26509});
	test_expansion(128'he9fc74951ca66606e14cf902b5f22083, {16'd1961, 16'd23596, 16'd35968, 16'd39410, 16'd1841, 16'd7292, 16'd39387, 16'd56255, 16'd28997, 16'd34576, 16'd44357, 16'd25293, 16'd9122, 16'd29831, 16'd56127, 16'd52487, 16'd38534, 16'd14579, 16'd19563, 16'd15180, 16'd16597, 16'd28292, 16'd52561, 16'd16645, 16'd19761, 16'd26438});
	test_expansion(128'h4b7493ed156d1e247552d59eff8f438e, {16'd49290, 16'd30382, 16'd10205, 16'd21205, 16'd29539, 16'd52192, 16'd31437, 16'd3610, 16'd5068, 16'd7805, 16'd6584, 16'd27642, 16'd58151, 16'd18404, 16'd12144, 16'd60311, 16'd34878, 16'd27979, 16'd2447, 16'd20585, 16'd19747, 16'd44425, 16'd56566, 16'd57769, 16'd34463, 16'd54750});
	test_expansion(128'h53b47d961a7e6a59bfbd11b8f5422231, {16'd21994, 16'd16989, 16'd7191, 16'd3823, 16'd6651, 16'd65274, 16'd53859, 16'd35231, 16'd15346, 16'd50210, 16'd14875, 16'd762, 16'd57544, 16'd14026, 16'd12319, 16'd61106, 16'd37802, 16'd44890, 16'd13753, 16'd2391, 16'd13301, 16'd2659, 16'd28564, 16'd38827, 16'd17361, 16'd24843});
	test_expansion(128'he32274e97b03b8db0a36a85ec238758f, {16'd62867, 16'd13564, 16'd35120, 16'd22015, 16'd8248, 16'd10667, 16'd55220, 16'd52576, 16'd35405, 16'd28995, 16'd22260, 16'd48454, 16'd15711, 16'd5522, 16'd16793, 16'd41527, 16'd59340, 16'd13260, 16'd14313, 16'd19865, 16'd7958, 16'd50705, 16'd60818, 16'd9948, 16'd41348, 16'd9970});
	test_expansion(128'ha3e6e2eed2f4126bb42a50264cad1939, {16'd31314, 16'd14675, 16'd22402, 16'd10430, 16'd29681, 16'd61619, 16'd45597, 16'd42316, 16'd3998, 16'd56177, 16'd50077, 16'd23008, 16'd41435, 16'd37709, 16'd42379, 16'd57583, 16'd11630, 16'd56195, 16'd17786, 16'd28613, 16'd46781, 16'd37276, 16'd42136, 16'd5975, 16'd23355, 16'd19655});
	test_expansion(128'h93c6eb8615119ae64c602b496fa91db2, {16'd53167, 16'd15738, 16'd43678, 16'd1671, 16'd49538, 16'd45269, 16'd17068, 16'd2243, 16'd62080, 16'd30564, 16'd11605, 16'd29730, 16'd32080, 16'd51070, 16'd58878, 16'd23965, 16'd39726, 16'd41538, 16'd7478, 16'd33621, 16'd49827, 16'd41672, 16'd25527, 16'd57285, 16'd64638, 16'd26633});
	test_expansion(128'hcf64719b125e6035e5f7dc638092b903, {16'd26412, 16'd39155, 16'd15815, 16'd3572, 16'd6393, 16'd44037, 16'd61261, 16'd53031, 16'd65062, 16'd25937, 16'd33099, 16'd30704, 16'd44822, 16'd59455, 16'd23161, 16'd42844, 16'd51550, 16'd36741, 16'd113, 16'd57847, 16'd58946, 16'd56048, 16'd57352, 16'd17737, 16'd28165, 16'd52478});
	test_expansion(128'h2613cc0da9e0006820743162742e6bbc, {16'd915, 16'd8341, 16'd55835, 16'd38705, 16'd56978, 16'd36976, 16'd3807, 16'd11576, 16'd56188, 16'd11950, 16'd25301, 16'd1717, 16'd8168, 16'd33803, 16'd30199, 16'd11371, 16'd55603, 16'd13987, 16'd32996, 16'd41982, 16'd45260, 16'd17064, 16'd36013, 16'd25100, 16'd46958, 16'd9063});
	test_expansion(128'he94a9e92863cb92dd0c68db84eaee8d9, {16'd43661, 16'd1723, 16'd14548, 16'd43961, 16'd17411, 16'd13520, 16'd10285, 16'd13252, 16'd27633, 16'd32549, 16'd35521, 16'd12154, 16'd46744, 16'd11846, 16'd46173, 16'd37165, 16'd41175, 16'd59445, 16'd34842, 16'd51355, 16'd43576, 16'd35394, 16'd14020, 16'd15889, 16'd10235, 16'd19442});
	test_expansion(128'h33626fb19db9faac3edf03c88cc6e6a3, {16'd44096, 16'd13189, 16'd41223, 16'd42335, 16'd35860, 16'd15838, 16'd61275, 16'd21704, 16'd57758, 16'd28163, 16'd17445, 16'd49726, 16'd29064, 16'd1684, 16'd64125, 16'd46138, 16'd1649, 16'd18021, 16'd18794, 16'd56216, 16'd9428, 16'd27551, 16'd6222, 16'd26878, 16'd58869, 16'd54720});
	test_expansion(128'h6754d6b8275e2aebf191fa44f07e4d67, {16'd60232, 16'd42505, 16'd18848, 16'd44877, 16'd51701, 16'd5231, 16'd5020, 16'd62064, 16'd30995, 16'd56833, 16'd1527, 16'd53996, 16'd52787, 16'd47507, 16'd6668, 16'd65326, 16'd29248, 16'd33399, 16'd9474, 16'd3314, 16'd43112, 16'd54935, 16'd21735, 16'd1296, 16'd25527, 16'd7349});
	test_expansion(128'h7cde219e471c7256fcedba4a897ce7c1, {16'd22747, 16'd48115, 16'd28449, 16'd10737, 16'd9464, 16'd47623, 16'd51314, 16'd21243, 16'd12391, 16'd9689, 16'd57469, 16'd10090, 16'd38815, 16'd29736, 16'd29264, 16'd51208, 16'd54070, 16'd50432, 16'd13855, 16'd17640, 16'd38189, 16'd64067, 16'd26848, 16'd55933, 16'd52371, 16'd40963});
	test_expansion(128'hcfdaefbac4829a164f438b888e66c66e, {16'd52193, 16'd65420, 16'd58643, 16'd6586, 16'd65164, 16'd63432, 16'd60191, 16'd4982, 16'd4495, 16'd45764, 16'd60758, 16'd17076, 16'd23610, 16'd51871, 16'd30000, 16'd55605, 16'd23504, 16'd197, 16'd64690, 16'd56019, 16'd15554, 16'd2775, 16'd35276, 16'd63142, 16'd45889, 16'd46756});
	test_expansion(128'hd3a664349592b7b93a01f67acb02825d, {16'd42814, 16'd6065, 16'd60422, 16'd9719, 16'd4664, 16'd63341, 16'd53420, 16'd9276, 16'd52175, 16'd25124, 16'd7949, 16'd50152, 16'd50316, 16'd41645, 16'd46821, 16'd17803, 16'd37774, 16'd37090, 16'd56145, 16'd19082, 16'd14947, 16'd13959, 16'd4331, 16'd5850, 16'd40117, 16'd61634});
	test_expansion(128'h188deb11bdf6abba5b60de66e336a7d3, {16'd31616, 16'd48819, 16'd20971, 16'd17009, 16'd29502, 16'd3285, 16'd30237, 16'd47748, 16'd16800, 16'd36257, 16'd36940, 16'd31971, 16'd52493, 16'd17412, 16'd24846, 16'd42444, 16'd64522, 16'd8738, 16'd27270, 16'd34419, 16'd65023, 16'd53603, 16'd3232, 16'd19221, 16'd22504, 16'd56217});
	test_expansion(128'hb925865f0c274e0807aa78e6e7045587, {16'd32443, 16'd57712, 16'd15731, 16'd57532, 16'd13779, 16'd26096, 16'd5852, 16'd49470, 16'd18644, 16'd25383, 16'd28328, 16'd2042, 16'd8090, 16'd45788, 16'd63580, 16'd2897, 16'd1094, 16'd50223, 16'd4782, 16'd62079, 16'd59308, 16'd15797, 16'd42033, 16'd62614, 16'd65377, 16'd45800});
	test_expansion(128'h1a1208e685bdc369a8a9e8bdafbcdad2, {16'd59613, 16'd8735, 16'd55722, 16'd45213, 16'd34705, 16'd58228, 16'd51259, 16'd31927, 16'd34910, 16'd19043, 16'd61253, 16'd49090, 16'd38924, 16'd22398, 16'd24569, 16'd37171, 16'd43653, 16'd51338, 16'd7658, 16'd49930, 16'd22442, 16'd60031, 16'd55725, 16'd61549, 16'd62431, 16'd4750});
	test_expansion(128'hedae52ba1621ab70248835ad74241fd4, {16'd39464, 16'd11516, 16'd30441, 16'd21684, 16'd8853, 16'd22366, 16'd41935, 16'd29709, 16'd37524, 16'd46144, 16'd35348, 16'd39112, 16'd11844, 16'd34809, 16'd26491, 16'd64070, 16'd43211, 16'd50656, 16'd30129, 16'd31550, 16'd4292, 16'd28619, 16'd52821, 16'd49655, 16'd4344, 16'd1280});
	test_expansion(128'h86b534bbf06af21c6f12f7890cd14680, {16'd26971, 16'd39054, 16'd43055, 16'd47399, 16'd4851, 16'd53062, 16'd15920, 16'd24045, 16'd18593, 16'd21067, 16'd65140, 16'd38310, 16'd32715, 16'd28745, 16'd1429, 16'd14215, 16'd16000, 16'd21705, 16'd33335, 16'd10977, 16'd51728, 16'd48592, 16'd11617, 16'd26681, 16'd17893, 16'd10365});
	test_expansion(128'h67d451b8d003bc52373d9859da0b8b05, {16'd51484, 16'd44247, 16'd10785, 16'd2216, 16'd17982, 16'd20044, 16'd5674, 16'd26365, 16'd11960, 16'd44441, 16'd56081, 16'd49870, 16'd31692, 16'd25889, 16'd63505, 16'd48958, 16'd16817, 16'd43465, 16'd24108, 16'd45414, 16'd12240, 16'd29061, 16'd42428, 16'd36391, 16'd51717, 16'd3461});
	test_expansion(128'h3b2dbf79b0c88b7da7e6652d8cdc2242, {16'd10146, 16'd24603, 16'd58898, 16'd25180, 16'd40329, 16'd25169, 16'd7217, 16'd38112, 16'd57158, 16'd64686, 16'd35642, 16'd12403, 16'd46584, 16'd56787, 16'd35622, 16'd38994, 16'd8870, 16'd55217, 16'd24087, 16'd16980, 16'd18096, 16'd7472, 16'd24806, 16'd42563, 16'd3350, 16'd34199});
	test_expansion(128'hd28a548f388d105a2b1cfe81cb5d232e, {16'd18305, 16'd53507, 16'd25935, 16'd45112, 16'd2212, 16'd6189, 16'd9432, 16'd41168, 16'd26015, 16'd38667, 16'd16616, 16'd23731, 16'd28438, 16'd42711, 16'd32907, 16'd24655, 16'd54063, 16'd33717, 16'd13336, 16'd14493, 16'd11558, 16'd31165, 16'd46472, 16'd23879, 16'd30255, 16'd51521});
	test_expansion(128'ha5a0e8b89d37299b277899785385eb80, {16'd57463, 16'd22538, 16'd65146, 16'd63189, 16'd57759, 16'd63050, 16'd28657, 16'd7234, 16'd56884, 16'd3949, 16'd42194, 16'd32710, 16'd62243, 16'd44062, 16'd31819, 16'd12883, 16'd17812, 16'd21268, 16'd53401, 16'd7169, 16'd33920, 16'd23151, 16'd42209, 16'd30249, 16'd30684, 16'd63223});
	test_expansion(128'hc43f070d4f8e3c625d9bbd6c0f58a79d, {16'd23323, 16'd52615, 16'd64788, 16'd25899, 16'd20404, 16'd31694, 16'd22133, 16'd33864, 16'd27203, 16'd29302, 16'd34652, 16'd39613, 16'd46468, 16'd7747, 16'd50382, 16'd43373, 16'd44267, 16'd33857, 16'd57383, 16'd62361, 16'd39779, 16'd55442, 16'd50207, 16'd10365, 16'd40204, 16'd245});
	test_expansion(128'hf779a7c21c394d24d6d213bf4f2414e6, {16'd56640, 16'd17002, 16'd65227, 16'd41266, 16'd27139, 16'd49653, 16'd36872, 16'd34365, 16'd18968, 16'd2337, 16'd51714, 16'd44206, 16'd64632, 16'd56562, 16'd26739, 16'd58629, 16'd58655, 16'd29591, 16'd19208, 16'd42259, 16'd28906, 16'd7595, 16'd51163, 16'd24009, 16'd51858, 16'd40305});
	test_expansion(128'h4c80d593e4cd5151666cbbb8fe42bfad, {16'd1559, 16'd23986, 16'd47039, 16'd58395, 16'd25997, 16'd41755, 16'd59041, 16'd46158, 16'd55743, 16'd46425, 16'd33893, 16'd24588, 16'd28021, 16'd13316, 16'd51970, 16'd28652, 16'd59424, 16'd25971, 16'd56122, 16'd4051, 16'd59261, 16'd59130, 16'd51906, 16'd15389, 16'd51858, 16'd56905});
	test_expansion(128'h9bac522511e8e89fca854e1f4992e71e, {16'd65314, 16'd12785, 16'd13231, 16'd29366, 16'd50242, 16'd41771, 16'd54733, 16'd37834, 16'd29995, 16'd1262, 16'd62704, 16'd45477, 16'd2302, 16'd16683, 16'd16241, 16'd59181, 16'd5494, 16'd40049, 16'd23342, 16'd33765, 16'd29574, 16'd4105, 16'd50405, 16'd59633, 16'd40340, 16'd3912});
	test_expansion(128'h1ae560cb249c4b8ed69cdd706d4fd066, {16'd26140, 16'd7151, 16'd33626, 16'd18633, 16'd63011, 16'd62790, 16'd10484, 16'd65471, 16'd53862, 16'd13654, 16'd2385, 16'd33613, 16'd32547, 16'd29563, 16'd10462, 16'd35842, 16'd56493, 16'd4562, 16'd29894, 16'd34690, 16'd61908, 16'd6923, 16'd36963, 16'd28495, 16'd24630, 16'd4683});
	test_expansion(128'ha10175696181677bae51387d017f0d8d, {16'd3786, 16'd33268, 16'd61711, 16'd11088, 16'd38998, 16'd2338, 16'd47886, 16'd35414, 16'd35332, 16'd29863, 16'd5444, 16'd2533, 16'd29262, 16'd59665, 16'd41183, 16'd24893, 16'd30325, 16'd27861, 16'd48812, 16'd37512, 16'd34829, 16'd64949, 16'd52403, 16'd58574, 16'd23842, 16'd58688});
	test_expansion(128'h3274e38aec56cf8e3ee6e8ffb7208878, {16'd22642, 16'd4867, 16'd61346, 16'd37632, 16'd57725, 16'd39798, 16'd5261, 16'd61313, 16'd33459, 16'd41521, 16'd1916, 16'd1697, 16'd46021, 16'd40104, 16'd52318, 16'd53437, 16'd42251, 16'd37469, 16'd20786, 16'd53960, 16'd9125, 16'd43972, 16'd4104, 16'd22720, 16'd50311, 16'd64151});
	test_expansion(128'h36558d05ba1f0b02004413303877c54e, {16'd22645, 16'd55783, 16'd176, 16'd45709, 16'd6555, 16'd43455, 16'd60072, 16'd58447, 16'd31425, 16'd19283, 16'd10714, 16'd34706, 16'd24910, 16'd34256, 16'd21429, 16'd28812, 16'd37589, 16'd56628, 16'd24341, 16'd52696, 16'd18660, 16'd37277, 16'd35789, 16'd35338, 16'd18615, 16'd40104});
	test_expansion(128'h6909ad46fe155a6b17288bbacca10239, {16'd22778, 16'd3617, 16'd29748, 16'd49688, 16'd64626, 16'd60745, 16'd19998, 16'd49597, 16'd4059, 16'd17745, 16'd2724, 16'd59194, 16'd51962, 16'd60831, 16'd19337, 16'd26548, 16'd20443, 16'd35184, 16'd40558, 16'd52795, 16'd5622, 16'd35978, 16'd61698, 16'd62394, 16'd51228, 16'd21198});
	test_expansion(128'hc7c96d208fc001b20b667881371f5756, {16'd42677, 16'd44355, 16'd278, 16'd48705, 16'd35332, 16'd60608, 16'd45536, 16'd65229, 16'd18195, 16'd48356, 16'd38632, 16'd38445, 16'd22822, 16'd8613, 16'd43608, 16'd56189, 16'd58119, 16'd38066, 16'd24164, 16'd31156, 16'd12803, 16'd8018, 16'd46247, 16'd61005, 16'd14422, 16'd1214});
	test_expansion(128'h04ed2d195c9112c83add8dbbc79d6e72, {16'd49815, 16'd35454, 16'd34443, 16'd44252, 16'd51989, 16'd47291, 16'd49811, 16'd58739, 16'd18437, 16'd17532, 16'd48537, 16'd61381, 16'd58395, 16'd12290, 16'd41785, 16'd43789, 16'd48048, 16'd61083, 16'd32737, 16'd16839, 16'd57277, 16'd10233, 16'd401, 16'd7826, 16'd36208, 16'd24857});
	test_expansion(128'h914ca1925c5b9f38f17bc43bf2ba4dda, {16'd47719, 16'd18853, 16'd14402, 16'd59652, 16'd7737, 16'd27253, 16'd40920, 16'd51560, 16'd46079, 16'd63433, 16'd25894, 16'd59814, 16'd20532, 16'd1239, 16'd27804, 16'd36544, 16'd55598, 16'd35901, 16'd13629, 16'd3333, 16'd9033, 16'd24929, 16'd62750, 16'd13894, 16'd28078, 16'd48877});
	test_expansion(128'hdb9dcb94fb67a7d64f1e9b4bf5f99734, {16'd34940, 16'd57411, 16'd49972, 16'd36726, 16'd37986, 16'd50802, 16'd13156, 16'd19772, 16'd51502, 16'd52194, 16'd27432, 16'd12272, 16'd58449, 16'd15395, 16'd11160, 16'd57050, 16'd45589, 16'd28384, 16'd7482, 16'd4204, 16'd17570, 16'd12176, 16'd26839, 16'd13026, 16'd55230, 16'd37752});
	test_expansion(128'h8bf6ca88a6d53cd6a2db7eace9cd8dc2, {16'd39690, 16'd5183, 16'd28308, 16'd8749, 16'd37351, 16'd12123, 16'd12949, 16'd4297, 16'd55770, 16'd43063, 16'd8644, 16'd54403, 16'd45903, 16'd6652, 16'd43837, 16'd21415, 16'd65283, 16'd52920, 16'd17804, 16'd64189, 16'd61304, 16'd40728, 16'd3146, 16'd61973, 16'd25284, 16'd19961});
	test_expansion(128'hea56a7aeade87985372f5624a0adfa6a, {16'd29321, 16'd50643, 16'd1705, 16'd9975, 16'd32244, 16'd51312, 16'd28807, 16'd32523, 16'd10798, 16'd45532, 16'd19434, 16'd57330, 16'd28168, 16'd40226, 16'd59964, 16'd4105, 16'd8295, 16'd41143, 16'd43930, 16'd51754, 16'd57532, 16'd62783, 16'd19777, 16'd52784, 16'd54057, 16'd51363});
	test_expansion(128'h4ccc454569ae8b4bce98784d4c7eea12, {16'd50219, 16'd26255, 16'd27926, 16'd20768, 16'd45051, 16'd43335, 16'd24667, 16'd22554, 16'd40772, 16'd50583, 16'd54812, 16'd29551, 16'd60436, 16'd11346, 16'd23816, 16'd49558, 16'd9224, 16'd54263, 16'd2268, 16'd41863, 16'd29793, 16'd35019, 16'd43700, 16'd49103, 16'd998, 16'd48438});
	test_expansion(128'he99bcac73a2f0e04bb8ee0bf394a8c0e, {16'd48484, 16'd14184, 16'd7525, 16'd19661, 16'd60567, 16'd18711, 16'd49921, 16'd9315, 16'd7046, 16'd50596, 16'd29745, 16'd52319, 16'd55693, 16'd7310, 16'd7559, 16'd22825, 16'd13942, 16'd61538, 16'd21204, 16'd42116, 16'd51748, 16'd29397, 16'd43909, 16'd50259, 16'd53386, 16'd25304});
	test_expansion(128'h12f028c3da59ea7f4912a40f1477a54f, {16'd49292, 16'd7196, 16'd11844, 16'd50175, 16'd56973, 16'd9206, 16'd7479, 16'd47064, 16'd50210, 16'd20388, 16'd59146, 16'd59405, 16'd14929, 16'd47313, 16'd25128, 16'd29067, 16'd61673, 16'd48457, 16'd27020, 16'd41406, 16'd5551, 16'd10888, 16'd8518, 16'd6144, 16'd59408, 16'd11714});
	test_expansion(128'h063c618ad53fb1325a9391fb59e20bfb, {16'd1039, 16'd44012, 16'd56750, 16'd38196, 16'd4504, 16'd23425, 16'd4, 16'd15806, 16'd19085, 16'd2854, 16'd9364, 16'd10229, 16'd59252, 16'd64471, 16'd5642, 16'd54086, 16'd35207, 16'd55458, 16'd32107, 16'd48864, 16'd31551, 16'd58562, 16'd14246, 16'd54157, 16'd64249, 16'd39378});
	test_expansion(128'hff7c14819e1db21ae7fb1c9b2bc594dc, {16'd56281, 16'd4575, 16'd55919, 16'd2624, 16'd59799, 16'd61015, 16'd64409, 16'd18975, 16'd63261, 16'd11184, 16'd9958, 16'd53983, 16'd50728, 16'd29071, 16'd33855, 16'd39280, 16'd15535, 16'd41882, 16'd15417, 16'd50757, 16'd49360, 16'd6149, 16'd12967, 16'd29737, 16'd31915, 16'd7970});
	test_expansion(128'h6c57a839107a674510061d3caf1290ca, {16'd5692, 16'd30130, 16'd6412, 16'd51509, 16'd25489, 16'd45846, 16'd46240, 16'd35043, 16'd24167, 16'd57098, 16'd43106, 16'd24368, 16'd32092, 16'd42455, 16'd54592, 16'd59480, 16'd10507, 16'd4730, 16'd5028, 16'd16027, 16'd264, 16'd52270, 16'd33693, 16'd41682, 16'd61514, 16'd9178});
	test_expansion(128'h882bb3e5c61046c1b3282bf2de802dcb, {16'd64077, 16'd11393, 16'd63041, 16'd359, 16'd22901, 16'd48931, 16'd17388, 16'd22494, 16'd31608, 16'd12516, 16'd64108, 16'd17535, 16'd58109, 16'd12421, 16'd19682, 16'd2067, 16'd24811, 16'd45418, 16'd62244, 16'd61234, 16'd56067, 16'd20167, 16'd9636, 16'd50587, 16'd28228, 16'd44394});
	test_expansion(128'h2dc7ac3fa6d2e0df009a259b0ef996b3, {16'd31718, 16'd34253, 16'd62395, 16'd40338, 16'd1498, 16'd13508, 16'd8620, 16'd10981, 16'd7170, 16'd50705, 16'd33737, 16'd8583, 16'd63020, 16'd62713, 16'd16207, 16'd25482, 16'd49072, 16'd24293, 16'd38998, 16'd56054, 16'd58034, 16'd592, 16'd28225, 16'd28734, 16'd57948, 16'd44752});
	test_expansion(128'h851d27d076d4e56c25c9ba8baecc4049, {16'd62118, 16'd34724, 16'd28991, 16'd43637, 16'd54190, 16'd27836, 16'd35106, 16'd28589, 16'd23188, 16'd55, 16'd50675, 16'd35121, 16'd39668, 16'd29290, 16'd32356, 16'd31364, 16'd49153, 16'd52839, 16'd49112, 16'd34207, 16'd44193, 16'd37302, 16'd25795, 16'd58384, 16'd53664, 16'd58541});
	test_expansion(128'h626c9d63b59495c62bb044cadb53af87, {16'd39052, 16'd31653, 16'd52226, 16'd36122, 16'd64217, 16'd14606, 16'd21838, 16'd32605, 16'd49634, 16'd43545, 16'd39202, 16'd57190, 16'd51160, 16'd45690, 16'd41996, 16'd11124, 16'd54527, 16'd52853, 16'd19640, 16'd5687, 16'd53170, 16'd3446, 16'd48696, 16'd56372, 16'd39669, 16'd44231});
	test_expansion(128'h0a3c49b630088335d01ecd84bfd74d73, {16'd3975, 16'd9693, 16'd24593, 16'd5509, 16'd20451, 16'd37056, 16'd47242, 16'd22693, 16'd12358, 16'd7919, 16'd61538, 16'd45551, 16'd5630, 16'd7174, 16'd54198, 16'd11515, 16'd28772, 16'd22808, 16'd19082, 16'd56392, 16'd40454, 16'd42191, 16'd46157, 16'd8481, 16'd48915, 16'd39074});
	test_expansion(128'he5f23d4ecefa0be443e7ea8f23d69601, {16'd40357, 16'd32384, 16'd63650, 16'd30514, 16'd24459, 16'd16995, 16'd64298, 16'd21062, 16'd6550, 16'd22715, 16'd46471, 16'd44254, 16'd40671, 16'd21726, 16'd60621, 16'd3315, 16'd43858, 16'd54771, 16'd8096, 16'd8564, 16'd13327, 16'd10309, 16'd46122, 16'd62445, 16'd6846, 16'd30610});
	test_expansion(128'h06f0b18baf47a5fb1622cc197af66c5e, {16'd10636, 16'd60721, 16'd1643, 16'd60735, 16'd38215, 16'd61427, 16'd34865, 16'd27255, 16'd10764, 16'd21811, 16'd32065, 16'd58638, 16'd14247, 16'd33869, 16'd51328, 16'd52669, 16'd58557, 16'd33632, 16'd56124, 16'd34834, 16'd17241, 16'd39891, 16'd33829, 16'd29411, 16'd53902, 16'd15484});
	test_expansion(128'h4785d59eed829d2128427bb64c06361e, {16'd59731, 16'd37825, 16'd17363, 16'd65130, 16'd38006, 16'd21451, 16'd57699, 16'd7438, 16'd61080, 16'd24984, 16'd55763, 16'd32964, 16'd44911, 16'd40553, 16'd2107, 16'd6141, 16'd37842, 16'd52647, 16'd56485, 16'd15758, 16'd22945, 16'd65269, 16'd35228, 16'd62428, 16'd62079, 16'd57304});
	test_expansion(128'h35d2380d5bb0e014c949e0035860a2e3, {16'd21303, 16'd57566, 16'd30776, 16'd19296, 16'd26754, 16'd61634, 16'd43856, 16'd14890, 16'd40627, 16'd37268, 16'd46243, 16'd64140, 16'd47708, 16'd44125, 16'd1604, 16'd40729, 16'd7204, 16'd24343, 16'd61597, 16'd56083, 16'd3381, 16'd18270, 16'd27063, 16'd61705, 16'd17598, 16'd27552});
	test_expansion(128'hde221a5ea22a0af40b08c1ce1df04ddc, {16'd42939, 16'd31608, 16'd39678, 16'd26989, 16'd47357, 16'd19644, 16'd42003, 16'd19252, 16'd42204, 16'd10751, 16'd3262, 16'd56565, 16'd30844, 16'd41037, 16'd56576, 16'd18089, 16'd57085, 16'd10622, 16'd60821, 16'd47316, 16'd7324, 16'd51453, 16'd22994, 16'd19385, 16'd7316, 16'd9567});
	test_expansion(128'h3209e318a968482bc71cb660eb4b4f01, {16'd29736, 16'd64444, 16'd39703, 16'd52036, 16'd59944, 16'd131, 16'd47928, 16'd43926, 16'd11097, 16'd23096, 16'd21370, 16'd15459, 16'd63783, 16'd23850, 16'd9234, 16'd11955, 16'd14709, 16'd21730, 16'd16306, 16'd49376, 16'd40051, 16'd44480, 16'd7939, 16'd56050, 16'd47417, 16'd44644});
	test_expansion(128'h387c16557dffb931637c03670a339611, {16'd45719, 16'd54189, 16'd61676, 16'd45945, 16'd55387, 16'd8171, 16'd18894, 16'd54449, 16'd25292, 16'd33135, 16'd58054, 16'd29631, 16'd26186, 16'd31168, 16'd12770, 16'd21659, 16'd23020, 16'd16793, 16'd361, 16'd63413, 16'd47362, 16'd3277, 16'd21730, 16'd47538, 16'd63938, 16'd59114});
	test_expansion(128'h7164492596ed786eb05e9652c0168558, {16'd61369, 16'd60791, 16'd23111, 16'd44915, 16'd13356, 16'd18350, 16'd35747, 16'd60018, 16'd51712, 16'd21363, 16'd9878, 16'd14794, 16'd38697, 16'd59982, 16'd61837, 16'd29843, 16'd12530, 16'd58103, 16'd4197, 16'd30422, 16'd10312, 16'd63745, 16'd46663, 16'd14499, 16'd24682, 16'd31550});
	test_expansion(128'h1e2ccd7ae650fedf45e58915c3712f71, {16'd4224, 16'd35552, 16'd65040, 16'd39459, 16'd23087, 16'd16198, 16'd57692, 16'd63384, 16'd11070, 16'd6177, 16'd5223, 16'd35142, 16'd57645, 16'd7351, 16'd57296, 16'd9830, 16'd43010, 16'd12252, 16'd46613, 16'd36210, 16'd49296, 16'd42791, 16'd49760, 16'd19995, 16'd56732, 16'd10358});
	test_expansion(128'hab3dfa445f6fd5bd63b27813e0a8a64a, {16'd60092, 16'd50425, 16'd9918, 16'd13123, 16'd32893, 16'd41120, 16'd38, 16'd43447, 16'd61551, 16'd18053, 16'd56499, 16'd60329, 16'd51068, 16'd48940, 16'd61492, 16'd57653, 16'd580, 16'd11405, 16'd10890, 16'd52969, 16'd26088, 16'd57311, 16'd47103, 16'd32161, 16'd55869, 16'd29006});
	test_expansion(128'he39132403a906922b3acd49e7b409a3a, {16'd52750, 16'd28349, 16'd53829, 16'd65278, 16'd36456, 16'd4318, 16'd9560, 16'd5296, 16'd56922, 16'd50493, 16'd19744, 16'd35807, 16'd56523, 16'd13006, 16'd6390, 16'd65473, 16'd45127, 16'd33880, 16'd15734, 16'd63858, 16'd22299, 16'd6650, 16'd59655, 16'd12785, 16'd29913, 16'd50754});
	test_expansion(128'ha2720b2d3a66f8d2fd7916e3b3e9bd32, {16'd46342, 16'd64910, 16'd43720, 16'd22548, 16'd55445, 16'd36551, 16'd3771, 16'd65022, 16'd45080, 16'd29931, 16'd51724, 16'd18221, 16'd14674, 16'd52224, 16'd47047, 16'd37145, 16'd49579, 16'd42103, 16'd47814, 16'd29430, 16'd34021, 16'd19919, 16'd31532, 16'd5628, 16'd27814, 16'd16110});
	test_expansion(128'h110a4a8d9476faf305caf613808fa149, {16'd8914, 16'd46798, 16'd59590, 16'd49891, 16'd28696, 16'd11706, 16'd31372, 16'd29458, 16'd21821, 16'd18167, 16'd22759, 16'd60836, 16'd48111, 16'd28330, 16'd396, 16'd39972, 16'd30657, 16'd764, 16'd16973, 16'd24356, 16'd3408, 16'd32042, 16'd17304, 16'd43121, 16'd39700, 16'd1234});
	test_expansion(128'hd87b7f642574a3ea9e6b01ec3986f8ad, {16'd40089, 16'd21020, 16'd25258, 16'd53821, 16'd45226, 16'd46628, 16'd64646, 16'd1348, 16'd28130, 16'd9710, 16'd34321, 16'd37307, 16'd13383, 16'd6259, 16'd17481, 16'd40289, 16'd42594, 16'd34207, 16'd51382, 16'd2725, 16'd39295, 16'd3913, 16'd62391, 16'd33529, 16'd23281, 16'd38461});
	test_expansion(128'hede8e634fe07580dabe1aec25803eaba, {16'd9789, 16'd51104, 16'd32758, 16'd46237, 16'd28909, 16'd25494, 16'd47209, 16'd46513, 16'd16734, 16'd9566, 16'd52657, 16'd23162, 16'd59520, 16'd40754, 16'd9400, 16'd48540, 16'd5091, 16'd23944, 16'd13921, 16'd10448, 16'd14681, 16'd2755, 16'd32896, 16'd42924, 16'd26370, 16'd15926});
	test_expansion(128'h9550e52ff87d12d44ceae8c2e6d342db, {16'd31757, 16'd41380, 16'd28710, 16'd3187, 16'd36765, 16'd54300, 16'd8673, 16'd4594, 16'd11365, 16'd61539, 16'd43371, 16'd27491, 16'd20903, 16'd51082, 16'd2811, 16'd43893, 16'd61489, 16'd36653, 16'd58509, 16'd54778, 16'd30154, 16'd26667, 16'd52142, 16'd43277, 16'd12237, 16'd13871});
	test_expansion(128'h674a2ab869213f278821b55812daf287, {16'd63923, 16'd24833, 16'd54460, 16'd8340, 16'd458, 16'd45483, 16'd37508, 16'd11081, 16'd39376, 16'd2203, 16'd11679, 16'd34985, 16'd34587, 16'd11692, 16'd48748, 16'd30953, 16'd1859, 16'd1640, 16'd9027, 16'd50519, 16'd24591, 16'd35471, 16'd3282, 16'd49712, 16'd9936, 16'd31883});
	test_expansion(128'h1444e520185f462e4f10c2703515d943, {16'd4187, 16'd17601, 16'd5666, 16'd62058, 16'd46854, 16'd52601, 16'd18581, 16'd47336, 16'd64968, 16'd9320, 16'd44874, 16'd11507, 16'd59793, 16'd29947, 16'd58241, 16'd20806, 16'd33675, 16'd64627, 16'd39750, 16'd45011, 16'd60876, 16'd721, 16'd49292, 16'd14406, 16'd11347, 16'd32928});
	test_expansion(128'h57f42572d6aaad2fdd84aac49d74362b, {16'd22509, 16'd7471, 16'd37142, 16'd27653, 16'd5176, 16'd22709, 16'd32107, 16'd37731, 16'd29705, 16'd15318, 16'd40272, 16'd26214, 16'd6913, 16'd29443, 16'd32649, 16'd41573, 16'd37572, 16'd17965, 16'd6406, 16'd9936, 16'd59718, 16'd41937, 16'd9660, 16'd56680, 16'd12627, 16'd23958});
	test_expansion(128'h5420c46725fa7c70309a62ca7195c353, {16'd32774, 16'd57327, 16'd45236, 16'd54343, 16'd17809, 16'd19996, 16'd570, 16'd37106, 16'd60133, 16'd18129, 16'd11066, 16'd22448, 16'd48013, 16'd17604, 16'd43910, 16'd39092, 16'd37598, 16'd7279, 16'd2031, 16'd23530, 16'd58162, 16'd56947, 16'd13846, 16'd7894, 16'd4306, 16'd13009});
	test_expansion(128'h7530c52f4057e3c1da1f14619482f75f, {16'd7176, 16'd22720, 16'd49073, 16'd409, 16'd27253, 16'd50711, 16'd37985, 16'd11486, 16'd22156, 16'd8054, 16'd5056, 16'd3024, 16'd17036, 16'd62296, 16'd36002, 16'd43554, 16'd4163, 16'd45659, 16'd55159, 16'd32593, 16'd51763, 16'd6879, 16'd40352, 16'd30583, 16'd9774, 16'd57232});
	test_expansion(128'hac60e37154c938fb856b174fa5b5eae1, {16'd17225, 16'd62764, 16'd61034, 16'd21559, 16'd8293, 16'd24019, 16'd27388, 16'd15617, 16'd14685, 16'd24551, 16'd8702, 16'd53113, 16'd53574, 16'd21602, 16'd64699, 16'd797, 16'd48929, 16'd4281, 16'd13788, 16'd42803, 16'd47776, 16'd37051, 16'd33249, 16'd56109, 16'd29143, 16'd46784});
	test_expansion(128'he3022716a4c48e338a692550f54aa850, {16'd8880, 16'd38352, 16'd21893, 16'd11499, 16'd31778, 16'd55966, 16'd9706, 16'd40501, 16'd26753, 16'd20456, 16'd34471, 16'd34774, 16'd27327, 16'd60523, 16'd51223, 16'd54933, 16'd33342, 16'd1636, 16'd5966, 16'd6519, 16'd25534, 16'd40924, 16'd40250, 16'd63404, 16'd17970, 16'd1413});
	test_expansion(128'h4c900213c65c78a9ba0ee00086f5edd1, {16'd34013, 16'd53619, 16'd19812, 16'd3441, 16'd582, 16'd46902, 16'd35197, 16'd17863, 16'd5761, 16'd656, 16'd49576, 16'd58231, 16'd5410, 16'd23137, 16'd7332, 16'd21216, 16'd53598, 16'd3842, 16'd37684, 16'd14985, 16'd35973, 16'd18828, 16'd12652, 16'd24549, 16'd32608, 16'd61934});
	test_expansion(128'h8223f24a436e850f77aa4f63599f06be, {16'd33593, 16'd49371, 16'd32110, 16'd7213, 16'd61382, 16'd427, 16'd16932, 16'd13195, 16'd16229, 16'd30006, 16'd34074, 16'd17291, 16'd3887, 16'd10285, 16'd22455, 16'd25120, 16'd55518, 16'd54339, 16'd59174, 16'd46506, 16'd62185, 16'd7976, 16'd60489, 16'd2975, 16'd26108, 16'd32269});
	test_expansion(128'hecc8953d7a55b95341dce9aba3fbca1c, {16'd888, 16'd28077, 16'd38324, 16'd60455, 16'd54999, 16'd39419, 16'd51616, 16'd36825, 16'd51294, 16'd64959, 16'd40030, 16'd65520, 16'd6648, 16'd14706, 16'd29101, 16'd33376, 16'd21034, 16'd63701, 16'd10656, 16'd34375, 16'd42619, 16'd36141, 16'd2627, 16'd60070, 16'd9662, 16'd18168});
	test_expansion(128'h16cb4a46544d015fe652a5f7e1bc62c0, {16'd11356, 16'd33316, 16'd34380, 16'd1323, 16'd63890, 16'd29995, 16'd44349, 16'd62659, 16'd45034, 16'd10191, 16'd14356, 16'd26888, 16'd10052, 16'd33060, 16'd40689, 16'd63148, 16'd24343, 16'd1488, 16'd31748, 16'd2365, 16'd27097, 16'd8946, 16'd51733, 16'd13017, 16'd31713, 16'd25766});
	test_expansion(128'hee3540382c40f1957c7ac06e99a26dbc, {16'd53405, 16'd17267, 16'd18367, 16'd20633, 16'd39755, 16'd6938, 16'd6125, 16'd21547, 16'd64866, 16'd6679, 16'd18222, 16'd26631, 16'd7824, 16'd36573, 16'd25112, 16'd63425, 16'd8608, 16'd4570, 16'd16698, 16'd25088, 16'd751, 16'd15423, 16'd7439, 16'd16545, 16'd54364, 16'd39143});
	test_expansion(128'h12a47fdd0f57cb06ca7518f693854927, {16'd61594, 16'd36132, 16'd65428, 16'd55693, 16'd65405, 16'd28178, 16'd27832, 16'd23325, 16'd28556, 16'd39167, 16'd1694, 16'd36333, 16'd17775, 16'd55452, 16'd19259, 16'd42589, 16'd6515, 16'd62845, 16'd21323, 16'd1198, 16'd63761, 16'd21832, 16'd18331, 16'd1251, 16'd1748, 16'd7913});
	test_expansion(128'he7e7a51f611d62be39c7492f05fba54a, {16'd11516, 16'd379, 16'd37292, 16'd1426, 16'd59150, 16'd56157, 16'd37888, 16'd24747, 16'd62536, 16'd7963, 16'd30325, 16'd16523, 16'd24985, 16'd12233, 16'd40793, 16'd46853, 16'd37163, 16'd39857, 16'd32340, 16'd32931, 16'd708, 16'd28879, 16'd61747, 16'd9991, 16'd42834, 16'd13672});
	test_expansion(128'h2a75aa3726fff08cf322cd76891b69b0, {16'd57565, 16'd25713, 16'd5970, 16'd36870, 16'd49058, 16'd27176, 16'd54488, 16'd39996, 16'd110, 16'd29136, 16'd1655, 16'd46025, 16'd38919, 16'd15906, 16'd53654, 16'd13116, 16'd25123, 16'd5539, 16'd65007, 16'd18622, 16'd26955, 16'd19852, 16'd31920, 16'd23150, 16'd21033, 16'd5389});
	test_expansion(128'h9cc5b668c6693453e5d56deb04febf05, {16'd13193, 16'd45840, 16'd28767, 16'd6416, 16'd49044, 16'd42980, 16'd33826, 16'd56174, 16'd45293, 16'd35413, 16'd54326, 16'd45744, 16'd22090, 16'd32083, 16'd61817, 16'd18323, 16'd50107, 16'd60170, 16'd45048, 16'd6416, 16'd26658, 16'd23137, 16'd4542, 16'd24072, 16'd41106, 16'd196});
	test_expansion(128'h3004aecce3df4d5202ee160a04c13559, {16'd42168, 16'd58367, 16'd49507, 16'd3382, 16'd58585, 16'd12172, 16'd51402, 16'd7639, 16'd9083, 16'd49683, 16'd15553, 16'd20047, 16'd47017, 16'd53057, 16'd4048, 16'd12649, 16'd21037, 16'd8388, 16'd17585, 16'd18578, 16'd45986, 16'd13959, 16'd37606, 16'd14307, 16'd29878, 16'd18265});
	test_expansion(128'h4c79055c0e0718d9b9d1251bdda89736, {16'd45073, 16'd43838, 16'd35376, 16'd6785, 16'd16012, 16'd50811, 16'd26331, 16'd41398, 16'd49595, 16'd41323, 16'd56173, 16'd52010, 16'd12453, 16'd29960, 16'd42755, 16'd21230, 16'd14614, 16'd47753, 16'd26305, 16'd33392, 16'd1534, 16'd51151, 16'd14010, 16'd29158, 16'd31106, 16'd31448});
	test_expansion(128'hc6ecdea46aeecba6fcc551a2a1d06511, {16'd1635, 16'd10012, 16'd16880, 16'd17132, 16'd59297, 16'd52552, 16'd63363, 16'd1531, 16'd32289, 16'd34241, 16'd57051, 16'd6228, 16'd4322, 16'd33695, 16'd50141, 16'd13947, 16'd30694, 16'd38009, 16'd58185, 16'd32161, 16'd10409, 16'd46939, 16'd38450, 16'd17063, 16'd57230, 16'd383});
	test_expansion(128'h15f18bf4b46ed1d9f2fcaaa50e0629d2, {16'd43189, 16'd57861, 16'd38659, 16'd61779, 16'd6332, 16'd53471, 16'd17958, 16'd48038, 16'd9772, 16'd5814, 16'd5674, 16'd48021, 16'd23627, 16'd32389, 16'd27237, 16'd63949, 16'd53556, 16'd13787, 16'd27681, 16'd14257, 16'd20715, 16'd13514, 16'd64082, 16'd30481, 16'd52899, 16'd35221});
	test_expansion(128'h0b7e79fbc10510f778085567d5c386df, {16'd2546, 16'd14868, 16'd24701, 16'd41422, 16'd55298, 16'd53834, 16'd58153, 16'd11185, 16'd53060, 16'd49032, 16'd61802, 16'd10027, 16'd54377, 16'd49068, 16'd62056, 16'd36263, 16'd9070, 16'd15366, 16'd18007, 16'd20277, 16'd21409, 16'd13850, 16'd4424, 16'd24839, 16'd7252, 16'd29104});
	test_expansion(128'he199236854619844e1978713e9b55a4b, {16'd27205, 16'd62250, 16'd10486, 16'd16925, 16'd63547, 16'd4329, 16'd45908, 16'd11521, 16'd55086, 16'd54036, 16'd16309, 16'd27415, 16'd59549, 16'd10385, 16'd7273, 16'd58198, 16'd37737, 16'd53854, 16'd35250, 16'd6462, 16'd29050, 16'd2475, 16'd11607, 16'd31711, 16'd23648, 16'd49346});
	test_expansion(128'hbd3c8d6fffe8dd7b256cd042ff543fc2, {16'd4451, 16'd48656, 16'd47641, 16'd3794, 16'd13516, 16'd46438, 16'd12029, 16'd6098, 16'd59149, 16'd18172, 16'd48444, 16'd49545, 16'd1647, 16'd53255, 16'd35005, 16'd19589, 16'd21801, 16'd54156, 16'd43553, 16'd57844, 16'd31744, 16'd37404, 16'd34765, 16'd62237, 16'd31142, 16'd5740});
	test_expansion(128'h9beba1c81e347a6a191cd089c1d7bc95, {16'd4178, 16'd11058, 16'd49556, 16'd55771, 16'd46782, 16'd2016, 16'd51092, 16'd33514, 16'd16371, 16'd41380, 16'd52639, 16'd2698, 16'd53509, 16'd44296, 16'd37526, 16'd65045, 16'd9745, 16'd60804, 16'd17698, 16'd29725, 16'd54752, 16'd23088, 16'd53943, 16'd22592, 16'd34262, 16'd55059});
	test_expansion(128'h988c166a2994a578a956c00cd9bf9416, {16'd63486, 16'd15155, 16'd15158, 16'd30391, 16'd35572, 16'd763, 16'd24564, 16'd41330, 16'd64677, 16'd65073, 16'd32942, 16'd54784, 16'd62675, 16'd60680, 16'd28687, 16'd59147, 16'd22195, 16'd14474, 16'd73, 16'd9450, 16'd5553, 16'd21651, 16'd19840, 16'd2149, 16'd31600, 16'd8036});
	test_expansion(128'h15e51ef50bc790bd79480de2cc7133c1, {16'd44645, 16'd43082, 16'd34807, 16'd19709, 16'd40324, 16'd40694, 16'd50546, 16'd59591, 16'd9594, 16'd8182, 16'd18562, 16'd58652, 16'd25689, 16'd23113, 16'd62813, 16'd11065, 16'd41393, 16'd10001, 16'd7706, 16'd31405, 16'd6672, 16'd35707, 16'd6151, 16'd52179, 16'd18647, 16'd15228});
	test_expansion(128'hbe729edeaa95774876ee534c4e9a42e7, {16'd4930, 16'd28641, 16'd8950, 16'd11665, 16'd10612, 16'd54940, 16'd33423, 16'd40185, 16'd64887, 16'd56980, 16'd51981, 16'd52968, 16'd26237, 16'd19072, 16'd35059, 16'd9840, 16'd3441, 16'd9747, 16'd7506, 16'd9848, 16'd28214, 16'd57492, 16'd8847, 16'd51651, 16'd45779, 16'd23996});
	test_expansion(128'h49ca1969fb7cac4f0aa21170a5214c1e, {16'd290, 16'd4930, 16'd38282, 16'd20422, 16'd17144, 16'd43652, 16'd32583, 16'd41304, 16'd46320, 16'd57455, 16'd50413, 16'd30677, 16'd48743, 16'd60985, 16'd47169, 16'd63593, 16'd26736, 16'd53070, 16'd27603, 16'd21377, 16'd6181, 16'd35503, 16'd23541, 16'd62227, 16'd61161, 16'd8756});
	test_expansion(128'h68ef7fd426507033ef44a0b457bdba8d, {16'd5418, 16'd57929, 16'd27089, 16'd33592, 16'd27063, 16'd63661, 16'd9106, 16'd27530, 16'd56249, 16'd49782, 16'd39356, 16'd33718, 16'd18758, 16'd35762, 16'd45093, 16'd1722, 16'd41931, 16'd39627, 16'd52240, 16'd17252, 16'd23180, 16'd22631, 16'd41431, 16'd36480, 16'd58581, 16'd62326});
	test_expansion(128'hb8953e0085e96671abb5e2bf66deb38d, {16'd4430, 16'd20812, 16'd27296, 16'd15839, 16'd61408, 16'd7622, 16'd5784, 16'd24201, 16'd55188, 16'd57493, 16'd42316, 16'd13027, 16'd45128, 16'd2296, 16'd30446, 16'd18912, 16'd43392, 16'd44932, 16'd816, 16'd8783, 16'd54365, 16'd62419, 16'd53941, 16'd31904, 16'd55424, 16'd54592});
	test_expansion(128'h1cbb4cef090abd2b9af9243ffbfd4aaa, {16'd4314, 16'd31006, 16'd12703, 16'd11399, 16'd2262, 16'd17387, 16'd57605, 16'd24405, 16'd12626, 16'd43311, 16'd26314, 16'd55650, 16'd21602, 16'd162, 16'd42465, 16'd46141, 16'd19501, 16'd45126, 16'd54436, 16'd21913, 16'd45326, 16'd9516, 16'd20701, 16'd54283, 16'd39574, 16'd58792});
	test_expansion(128'h8b9f3a0e47ff6c1a394aa4310dff8b84, {16'd62719, 16'd29991, 16'd16398, 16'd1511, 16'd36229, 16'd64664, 16'd53334, 16'd34954, 16'd27677, 16'd52218, 16'd29543, 16'd53400, 16'd9821, 16'd25768, 16'd45836, 16'd19747, 16'd51379, 16'd43964, 16'd6939, 16'd10547, 16'd55896, 16'd45132, 16'd45557, 16'd24566, 16'd54368, 16'd39364});
	test_expansion(128'hdcdf70afb82b83ebb6b8f33140db5d12, {16'd46226, 16'd65, 16'd46481, 16'd63806, 16'd57156, 16'd19925, 16'd51528, 16'd29236, 16'd62167, 16'd3170, 16'd57791, 16'd43955, 16'd22790, 16'd27074, 16'd53379, 16'd3091, 16'd8761, 16'd37976, 16'd58401, 16'd6739, 16'd65137, 16'd33080, 16'd60645, 16'd11448, 16'd5440, 16'd22722});
	test_expansion(128'h63dfb58013878fa42209a58b2726fe3b, {16'd5967, 16'd16447, 16'd10307, 16'd18013, 16'd56071, 16'd61048, 16'd56944, 16'd37619, 16'd46728, 16'd62296, 16'd2314, 16'd32172, 16'd26665, 16'd46805, 16'd32085, 16'd26263, 16'd56476, 16'd42593, 16'd61502, 16'd30525, 16'd4717, 16'd38184, 16'd48406, 16'd9880, 16'd41672, 16'd7253});
	test_expansion(128'hc630cd988eb1039e426471231029f9c6, {16'd4578, 16'd64593, 16'd33578, 16'd22864, 16'd11512, 16'd13013, 16'd32551, 16'd42165, 16'd54005, 16'd4919, 16'd7233, 16'd22338, 16'd28011, 16'd38881, 16'd61840, 16'd39191, 16'd50579, 16'd57075, 16'd40748, 16'd15293, 16'd34161, 16'd43820, 16'd27102, 16'd44647, 16'd26875, 16'd40167});
	test_expansion(128'hb36bdd6e877f407933aefd5958cba4be, {16'd26023, 16'd28614, 16'd42328, 16'd48013, 16'd47948, 16'd4839, 16'd61013, 16'd8696, 16'd22126, 16'd3156, 16'd28884, 16'd38535, 16'd48764, 16'd2624, 16'd49649, 16'd58130, 16'd28018, 16'd48182, 16'd57322, 16'd55600, 16'd2332, 16'd13186, 16'd8158, 16'd12282, 16'd49192, 16'd41842});
	test_expansion(128'h3ff5d223e7cfcecb36477053fca4f70c, {16'd46540, 16'd37092, 16'd22126, 16'd46930, 16'd40523, 16'd18294, 16'd25272, 16'd62655, 16'd14410, 16'd45125, 16'd11733, 16'd25679, 16'd62259, 16'd53226, 16'd271, 16'd47366, 16'd11395, 16'd12252, 16'd23658, 16'd55468, 16'd31940, 16'd58932, 16'd48225, 16'd18282, 16'd1488, 16'd19948});
	test_expansion(128'h6a6f537441c6d30fb8f48f737e9593ed, {16'd59370, 16'd64588, 16'd49062, 16'd61842, 16'd38843, 16'd53865, 16'd63137, 16'd8416, 16'd23373, 16'd4093, 16'd5042, 16'd785, 16'd9079, 16'd40801, 16'd56383, 16'd22198, 16'd58137, 16'd9790, 16'd48033, 16'd2239, 16'd53995, 16'd65481, 16'd7284, 16'd47086, 16'd902, 16'd21612});
	test_expansion(128'h45d63da5aa03848ebd711b6d503d54c7, {16'd4340, 16'd21960, 16'd58836, 16'd8938, 16'd49741, 16'd63499, 16'd9926, 16'd57698, 16'd39331, 16'd32898, 16'd51030, 16'd64315, 16'd61191, 16'd28131, 16'd47668, 16'd17222, 16'd35114, 16'd40872, 16'd18683, 16'd53987, 16'd39928, 16'd58704, 16'd60803, 16'd20769, 16'd59214, 16'd45401});
	test_expansion(128'h6607a9830172d91c21c0fe1fac2a8fd9, {16'd44706, 16'd10277, 16'd2894, 16'd48698, 16'd54052, 16'd64742, 16'd57636, 16'd58352, 16'd20759, 16'd19650, 16'd48904, 16'd7245, 16'd54960, 16'd44689, 16'd46142, 16'd49427, 16'd60962, 16'd30521, 16'd46490, 16'd1163, 16'd55772, 16'd12301, 16'd2357, 16'd45097, 16'd37978, 16'd7993});
	test_expansion(128'hb9a457dc9c8673da92ae535ac6806578, {16'd19329, 16'd31238, 16'd38539, 16'd53493, 16'd54623, 16'd36491, 16'd59881, 16'd14000, 16'd16766, 16'd6233, 16'd65119, 16'd50472, 16'd43873, 16'd13411, 16'd63829, 16'd61070, 16'd52925, 16'd61690, 16'd43165, 16'd27772, 16'd58161, 16'd56988, 16'd27731, 16'd24006, 16'd18741, 16'd19279});
	test_expansion(128'hf4552d45ad58a38716ed54666411040c, {16'd32648, 16'd48468, 16'd22188, 16'd25411, 16'd7208, 16'd4656, 16'd34930, 16'd26641, 16'd18860, 16'd40725, 16'd61691, 16'd65498, 16'd23555, 16'd19995, 16'd2061, 16'd60034, 16'd60508, 16'd44809, 16'd52314, 16'd30498, 16'd31771, 16'd5501, 16'd43309, 16'd16788, 16'd39396, 16'd37182});
	test_expansion(128'h3af6a563554434c7ecb3f5d8dcbf0113, {16'd15524, 16'd13045, 16'd2982, 16'd39203, 16'd28292, 16'd9218, 16'd44832, 16'd20413, 16'd50303, 16'd8177, 16'd23635, 16'd41159, 16'd20771, 16'd51148, 16'd62226, 16'd58160, 16'd55682, 16'd47281, 16'd17533, 16'd30019, 16'd27966, 16'd49241, 16'd38425, 16'd50834, 16'd19499, 16'd4848});
	test_expansion(128'haad9973e8c33cf808da26e9bb002c8da, {16'd7050, 16'd19555, 16'd65462, 16'd37616, 16'd50124, 16'd59242, 16'd57669, 16'd5414, 16'd46218, 16'd64958, 16'd56881, 16'd64894, 16'd651, 16'd65434, 16'd18441, 16'd50948, 16'd35310, 16'd5817, 16'd34477, 16'd4547, 16'd4996, 16'd57181, 16'd31739, 16'd10508, 16'd9189, 16'd62290});
	test_expansion(128'hc782a408766eb80d06e4a0aa15a2f917, {16'd27580, 16'd51740, 16'd56603, 16'd24321, 16'd33647, 16'd56863, 16'd55078, 16'd65288, 16'd58869, 16'd23675, 16'd31852, 16'd33715, 16'd54741, 16'd27266, 16'd25791, 16'd33313, 16'd64715, 16'd24128, 16'd49523, 16'd42524, 16'd52744, 16'd24796, 16'd328, 16'd27506, 16'd62913, 16'd6297});
	test_expansion(128'h7e18df2c3d0c8d1b94944822a5336b78, {16'd26419, 16'd2334, 16'd57191, 16'd912, 16'd22443, 16'd1745, 16'd64414, 16'd53177, 16'd48502, 16'd9962, 16'd19393, 16'd23591, 16'd12680, 16'd30474, 16'd22509, 16'd47215, 16'd18224, 16'd51896, 16'd65094, 16'd51135, 16'd31456, 16'd17352, 16'd29173, 16'd58184, 16'd11777, 16'd22344});
	test_expansion(128'h4054185854d83cf78e7ae30af61deada, {16'd417, 16'd52023, 16'd29188, 16'd15714, 16'd31597, 16'd48596, 16'd43790, 16'd44648, 16'd59520, 16'd17052, 16'd35753, 16'd5759, 16'd19781, 16'd41066, 16'd27601, 16'd62002, 16'd54596, 16'd58927, 16'd43713, 16'd45998, 16'd62934, 16'd12738, 16'd41921, 16'd5360, 16'd13436, 16'd42469});
	test_expansion(128'h7fb6768e6a1fc90bf19dca6724371a77, {16'd54470, 16'd57463, 16'd14998, 16'd58519, 16'd5952, 16'd60323, 16'd24547, 16'd19700, 16'd6397, 16'd8558, 16'd20805, 16'd23970, 16'd6476, 16'd38765, 16'd37113, 16'd33298, 16'd22255, 16'd29977, 16'd11370, 16'd5640, 16'd2553, 16'd64618, 16'd56722, 16'd42119, 16'd32802, 16'd12788});
	test_expansion(128'h6cd4a6dc3e17c733b8bd3ffdc1d7e584, {16'd3879, 16'd30125, 16'd43459, 16'd47116, 16'd64566, 16'd22315, 16'd7451, 16'd63552, 16'd9058, 16'd19178, 16'd30958, 16'd38533, 16'd27613, 16'd9404, 16'd49816, 16'd29803, 16'd53538, 16'd7592, 16'd19439, 16'd7319, 16'd16077, 16'd45254, 16'd22570, 16'd15812, 16'd53316, 16'd64386});
	test_expansion(128'hd0cbcb65d0c8d2b815de84afe1929a64, {16'd61278, 16'd43687, 16'd37396, 16'd53792, 16'd31375, 16'd36139, 16'd64235, 16'd1640, 16'd27375, 16'd2075, 16'd18831, 16'd22301, 16'd39520, 16'd26505, 16'd46759, 16'd37942, 16'd51794, 16'd48443, 16'd64157, 16'd40099, 16'd21869, 16'd57670, 16'd38766, 16'd55867, 16'd47008, 16'd38851});
	test_expansion(128'hf2cd45fffd736535b25804ef230b64f3, {16'd9164, 16'd15895, 16'd49227, 16'd55229, 16'd29084, 16'd36918, 16'd56544, 16'd2073, 16'd40258, 16'd32633, 16'd59627, 16'd28677, 16'd1574, 16'd2242, 16'd42970, 16'd24844, 16'd33923, 16'd15020, 16'd39529, 16'd10253, 16'd31137, 16'd30999, 16'd41570, 16'd4689, 16'd11174, 16'd58424});
	test_expansion(128'h49a1ab4196f1fec87ed7fa229f102f35, {16'd44456, 16'd59573, 16'd62103, 16'd8439, 16'd45057, 16'd38944, 16'd30521, 16'd24482, 16'd28465, 16'd40025, 16'd25902, 16'd57879, 16'd19214, 16'd29495, 16'd49019, 16'd33227, 16'd35241, 16'd1495, 16'd18347, 16'd45654, 16'd52613, 16'd10267, 16'd61090, 16'd2538, 16'd48425, 16'd25803});
	test_expansion(128'h0a0fa61d139f24d5418f84496ebb23ce, {16'd9481, 16'd29565, 16'd40230, 16'd49508, 16'd47628, 16'd2261, 16'd61812, 16'd45801, 16'd49336, 16'd13717, 16'd56903, 16'd24516, 16'd42689, 16'd46208, 16'd43905, 16'd37352, 16'd64418, 16'd38750, 16'd11774, 16'd5650, 16'd5365, 16'd11670, 16'd33837, 16'd60059, 16'd17616, 16'd13871});
	test_expansion(128'h773a3e118ecbc75a6d2b33bcdc2a992c, {16'd9047, 16'd38115, 16'd26723, 16'd47908, 16'd54676, 16'd34324, 16'd13665, 16'd19027, 16'd35301, 16'd20982, 16'd53465, 16'd27611, 16'd15609, 16'd12470, 16'd26968, 16'd19625, 16'd25600, 16'd20793, 16'd55271, 16'd29301, 16'd57070, 16'd53910, 16'd39832, 16'd47492, 16'd31204, 16'd20281});
	test_expansion(128'h1692824fccfe0e7688ea2adb70acc2d5, {16'd41826, 16'd44838, 16'd34327, 16'd22480, 16'd10701, 16'd9877, 16'd1143, 16'd17978, 16'd29872, 16'd50750, 16'd28961, 16'd24409, 16'd2978, 16'd51666, 16'd22920, 16'd44181, 16'd24214, 16'd25696, 16'd59526, 16'd65035, 16'd16934, 16'd29210, 16'd61393, 16'd56226, 16'd32017, 16'd22607});
	test_expansion(128'hd20536edeee4084d5c9c4a5ac4923741, {16'd44612, 16'd63152, 16'd20966, 16'd55380, 16'd8175, 16'd63642, 16'd17273, 16'd21822, 16'd28981, 16'd37010, 16'd45626, 16'd63053, 16'd59636, 16'd39780, 16'd24447, 16'd35973, 16'd2642, 16'd57727, 16'd44159, 16'd5799, 16'd11811, 16'd40209, 16'd17603, 16'd27103, 16'd59134, 16'd62785});
	test_expansion(128'hba576d5b05f29180bfff05340f8469a1, {16'd26535, 16'd46040, 16'd60835, 16'd10400, 16'd29466, 16'd52586, 16'd41402, 16'd50731, 16'd62606, 16'd14950, 16'd29015, 16'd43197, 16'd50631, 16'd1365, 16'd11936, 16'd22929, 16'd28472, 16'd22808, 16'd63433, 16'd34959, 16'd19639, 16'd8035, 16'd41970, 16'd61705, 16'd46401, 16'd16521});
	test_expansion(128'hcb3edbf81cb6a5cfd9705bde2f0d2bff, {16'd19183, 16'd50629, 16'd11075, 16'd45820, 16'd9440, 16'd65429, 16'd19491, 16'd25119, 16'd9423, 16'd62253, 16'd13821, 16'd50144, 16'd64457, 16'd17308, 16'd61959, 16'd32056, 16'd53810, 16'd48205, 16'd5001, 16'd39761, 16'd61123, 16'd62518, 16'd39077, 16'd8698, 16'd53755, 16'd14383});
	test_expansion(128'h7b68c0984f4e3d23ba43bbc52bba83bd, {16'd31004, 16'd8541, 16'd45213, 16'd27973, 16'd22957, 16'd52181, 16'd36315, 16'd28421, 16'd21290, 16'd5019, 16'd47968, 16'd25522, 16'd54708, 16'd12868, 16'd42649, 16'd19828, 16'd51716, 16'd11697, 16'd11323, 16'd2505, 16'd944, 16'd58232, 16'd12027, 16'd63480, 16'd22452, 16'd10678});
	test_expansion(128'hab760d4726a339d8c56263cfa6b4a26b, {16'd22853, 16'd48794, 16'd64532, 16'd41066, 16'd26843, 16'd56743, 16'd46674, 16'd34796, 16'd12077, 16'd12837, 16'd16887, 16'd29555, 16'd39454, 16'd58320, 16'd20196, 16'd3324, 16'd40659, 16'd5747, 16'd24535, 16'd11146, 16'd17869, 16'd45286, 16'd32402, 16'd57757, 16'd62156, 16'd38122});
	test_expansion(128'h6997f3dea115a74f952abbd08bfdb6b6, {16'd54476, 16'd1064, 16'd46146, 16'd18821, 16'd52529, 16'd59045, 16'd30904, 16'd2005, 16'd22939, 16'd588, 16'd44620, 16'd15099, 16'd55636, 16'd44121, 16'd9579, 16'd51315, 16'd29538, 16'd22474, 16'd49469, 16'd5659, 16'd22907, 16'd13741, 16'd45652, 16'd32439, 16'd58339, 16'd14990});
	test_expansion(128'he52c84109d1d59bd666ff21c98128dea, {16'd2056, 16'd40570, 16'd59157, 16'd8311, 16'd25611, 16'd36570, 16'd59523, 16'd7377, 16'd43372, 16'd60460, 16'd32665, 16'd24896, 16'd23051, 16'd30023, 16'd12598, 16'd45017, 16'd38744, 16'd32465, 16'd45502, 16'd45042, 16'd15067, 16'd37881, 16'd59141, 16'd549, 16'd14981, 16'd10870});
	test_expansion(128'h79889ad3b5fdf16f0b32b271edcb1703, {16'd64129, 16'd11172, 16'd61765, 16'd35570, 16'd4487, 16'd20787, 16'd928, 16'd25103, 16'd34311, 16'd41072, 16'd16335, 16'd56134, 16'd54397, 16'd61022, 16'd12993, 16'd24363, 16'd55641, 16'd60804, 16'd55385, 16'd60447, 16'd32035, 16'd35420, 16'd49468, 16'd40667, 16'd572, 16'd52034});
	test_expansion(128'h0030f2248a9dbcca43f1c4acb7350663, {16'd48353, 16'd51133, 16'd57464, 16'd6956, 16'd23282, 16'd60040, 16'd52457, 16'd59141, 16'd50656, 16'd15557, 16'd27497, 16'd15005, 16'd50907, 16'd60628, 16'd13676, 16'd60661, 16'd58173, 16'd41734, 16'd653, 16'd19777, 16'd56579, 16'd9400, 16'd44024, 16'd50886, 16'd13860, 16'd9789});
	test_expansion(128'hac123daf2c105421f603c8a9ecfe3d11, {16'd27042, 16'd5407, 16'd51604, 16'd20344, 16'd51767, 16'd36714, 16'd38128, 16'd12563, 16'd4202, 16'd45327, 16'd36954, 16'd51930, 16'd41152, 16'd591, 16'd41430, 16'd7286, 16'd13788, 16'd57894, 16'd47042, 16'd40889, 16'd37317, 16'd34524, 16'd14599, 16'd32395, 16'd11387, 16'd142});
	test_expansion(128'hcd5fbb3d9eca13bb6a1624d18fc29e2f, {16'd53503, 16'd26910, 16'd25216, 16'd24070, 16'd33277, 16'd53647, 16'd56474, 16'd14712, 16'd22178, 16'd64440, 16'd59989, 16'd42333, 16'd7235, 16'd1254, 16'd9028, 16'd56991, 16'd64862, 16'd3052, 16'd27304, 16'd41223, 16'd49532, 16'd30215, 16'd52454, 16'd17661, 16'd21651, 16'd24478});
	test_expansion(128'h7e3b6b0c90ef65c60d474da84eb0fb24, {16'd38434, 16'd58155, 16'd31384, 16'd1495, 16'd17447, 16'd43556, 16'd40562, 16'd34235, 16'd41947, 16'd64597, 16'd7576, 16'd49179, 16'd35059, 16'd168, 16'd24216, 16'd40176, 16'd6644, 16'd31436, 16'd53168, 16'd4030, 16'd56518, 16'd50661, 16'd28847, 16'd8587, 16'd42042, 16'd36165});
	test_expansion(128'hdbb4aba6edfc3d9f9c2f409b9b0b1c98, {16'd17346, 16'd36749, 16'd48706, 16'd50243, 16'd60980, 16'd22653, 16'd52801, 16'd58984, 16'd7296, 16'd26171, 16'd43319, 16'd32711, 16'd16009, 16'd60859, 16'd65006, 16'd5114, 16'd5600, 16'd23261, 16'd59366, 16'd61130, 16'd62496, 16'd21298, 16'd1484, 16'd59560, 16'd24259, 16'd53087});
	test_expansion(128'h4c880cc55bc97430d2c7e2b4d2f96f05, {16'd14839, 16'd25051, 16'd64793, 16'd62699, 16'd61255, 16'd61573, 16'd9126, 16'd7845, 16'd12634, 16'd28827, 16'd37653, 16'd37221, 16'd13819, 16'd7870, 16'd13159, 16'd49849, 16'd25743, 16'd56240, 16'd44481, 16'd4140, 16'd38190, 16'd50659, 16'd43268, 16'd26192, 16'd38442, 16'd12041});
	test_expansion(128'hf13fed3761249fbbe3fdb9385009f7f4, {16'd59198, 16'd13616, 16'd29956, 16'd23583, 16'd47055, 16'd30420, 16'd3685, 16'd9928, 16'd48554, 16'd6643, 16'd31619, 16'd30957, 16'd60284, 16'd47912, 16'd53132, 16'd33982, 16'd50057, 16'd51830, 16'd14376, 16'd65185, 16'd16622, 16'd2901, 16'd30537, 16'd15309, 16'd13732, 16'd33994});
	test_expansion(128'h5067f82796ffd2dc3536969f060146f8, {16'd47139, 16'd15242, 16'd3103, 16'd63961, 16'd30682, 16'd1710, 16'd40017, 16'd22899, 16'd8590, 16'd43948, 16'd46233, 16'd15946, 16'd34135, 16'd30594, 16'd30245, 16'd9729, 16'd40846, 16'd41730, 16'd61030, 16'd4474, 16'd46557, 16'd46883, 16'd61856, 16'd17280, 16'd16397, 16'd62668});
	test_expansion(128'h9a919083de4fef204ad046ea08201107, {16'd51745, 16'd56225, 16'd28201, 16'd44129, 16'd21655, 16'd52511, 16'd25042, 16'd51297, 16'd29880, 16'd7069, 16'd22025, 16'd53000, 16'd37886, 16'd61028, 16'd51643, 16'd33758, 16'd55789, 16'd36534, 16'd49276, 16'd13321, 16'd14882, 16'd29288, 16'd49754, 16'd59140, 16'd53582, 16'd53372});
	test_expansion(128'ha13f9b2bbe3905d08f5ae44551fb0fbc, {16'd57031, 16'd38306, 16'd12224, 16'd32351, 16'd55060, 16'd26025, 16'd50315, 16'd51218, 16'd19794, 16'd55899, 16'd64035, 16'd366, 16'd51765, 16'd63474, 16'd9423, 16'd36000, 16'd47918, 16'd23567, 16'd40555, 16'd49098, 16'd30685, 16'd64917, 16'd46433, 16'd24244, 16'd33899, 16'd8659});
	test_expansion(128'h8a1e7cbb3285b81905278a96fdf62ea3, {16'd18779, 16'd43062, 16'd41319, 16'd29471, 16'd56110, 16'd28217, 16'd64928, 16'd18177, 16'd16398, 16'd26330, 16'd28982, 16'd47495, 16'd57506, 16'd34465, 16'd4386, 16'd13830, 16'd60028, 16'd31626, 16'd35006, 16'd28558, 16'd48852, 16'd6973, 16'd4705, 16'd22523, 16'd41745, 16'd30301});
	test_expansion(128'h779ce036015838aa52cf72561eba9820, {16'd62281, 16'd42541, 16'd32274, 16'd14596, 16'd51883, 16'd61381, 16'd2503, 16'd16309, 16'd59139, 16'd47359, 16'd28398, 16'd12927, 16'd25203, 16'd9510, 16'd7100, 16'd41506, 16'd62906, 16'd35261, 16'd21728, 16'd46123, 16'd40583, 16'd30736, 16'd24545, 16'd22184, 16'd12439, 16'd31400});
	test_expansion(128'h08804e75f805409fb8ed59d1fa6676c3, {16'd24738, 16'd43507, 16'd3560, 16'd65067, 16'd37738, 16'd39, 16'd35916, 16'd36039, 16'd2908, 16'd55382, 16'd46720, 16'd25341, 16'd51469, 16'd37420, 16'd44476, 16'd5462, 16'd11269, 16'd28125, 16'd26610, 16'd34978, 16'd61208, 16'd40159, 16'd17236, 16'd65101, 16'd4335, 16'd35702});
	test_expansion(128'hfafc068cfd4135443c2cdbb2c8a46aa8, {16'd52151, 16'd1459, 16'd47165, 16'd47062, 16'd2677, 16'd4671, 16'd49836, 16'd41464, 16'd60386, 16'd10017, 16'd19602, 16'd40813, 16'd30738, 16'd63281, 16'd50746, 16'd39074, 16'd2714, 16'd64062, 16'd46561, 16'd51393, 16'd32550, 16'd6508, 16'd64355, 16'd38879, 16'd52507, 16'd53776});
	test_expansion(128'h392b612d874f8600d9e9fe1387df48ff, {16'd33627, 16'd57367, 16'd49802, 16'd46809, 16'd40550, 16'd24030, 16'd55438, 16'd54715, 16'd42823, 16'd34047, 16'd28154, 16'd3420, 16'd27490, 16'd3434, 16'd9546, 16'd49826, 16'd41464, 16'd51434, 16'd61397, 16'd24945, 16'd53753, 16'd15787, 16'd7280, 16'd30063, 16'd2400, 16'd9567});
	test_expansion(128'he3d9eb214fb8071ee631342102c73567, {16'd45583, 16'd34329, 16'd10797, 16'd26011, 16'd39441, 16'd53661, 16'd53680, 16'd37179, 16'd8840, 16'd56386, 16'd27007, 16'd24720, 16'd1688, 16'd41215, 16'd59241, 16'd5698, 16'd9606, 16'd62886, 16'd42503, 16'd40203, 16'd4376, 16'd49925, 16'd60729, 16'd21496, 16'd4203, 16'd21236});
	test_expansion(128'h38e05b8d7a2549911b7cdaec44590fe6, {16'd49918, 16'd61413, 16'd46503, 16'd62177, 16'd2856, 16'd54497, 16'd46809, 16'd60688, 16'd65059, 16'd58768, 16'd23954, 16'd54540, 16'd24672, 16'd47554, 16'd53266, 16'd28031, 16'd60400, 16'd18616, 16'd14353, 16'd25399, 16'd11605, 16'd26765, 16'd533, 16'd32409, 16'd30652, 16'd12916});
	test_expansion(128'h7749908e70ab9884f459ab0db60ca760, {16'd34112, 16'd555, 16'd34189, 16'd63622, 16'd4713, 16'd2324, 16'd27173, 16'd24820, 16'd25588, 16'd7719, 16'd63316, 16'd17491, 16'd28360, 16'd8699, 16'd2509, 16'd35289, 16'd52028, 16'd59347, 16'd45386, 16'd52382, 16'd7318, 16'd34475, 16'd59260, 16'd54207, 16'd57120, 16'd617});
	test_expansion(128'h1a25fdb9725a1f34401ddbe9278c0455, {16'd14404, 16'd32785, 16'd17733, 16'd40276, 16'd60558, 16'd49408, 16'd22408, 16'd46111, 16'd61767, 16'd49364, 16'd48148, 16'd3837, 16'd56489, 16'd16296, 16'd31983, 16'd33182, 16'd34393, 16'd48645, 16'd47121, 16'd38502, 16'd33100, 16'd2158, 16'd7581, 16'd36786, 16'd23120, 16'd26808});
	test_expansion(128'h56c79927ff366e46d2e48bc6d9f81f14, {16'd10206, 16'd58994, 16'd26044, 16'd49854, 16'd39296, 16'd41659, 16'd39048, 16'd52880, 16'd50213, 16'd32771, 16'd49094, 16'd22351, 16'd13498, 16'd50475, 16'd13952, 16'd43614, 16'd40002, 16'd50128, 16'd41561, 16'd37327, 16'd12884, 16'd45027, 16'd16039, 16'd31672, 16'd18691, 16'd36767});
	test_expansion(128'h849f0d94886b776ad9c275568cbd715e, {16'd51546, 16'd37506, 16'd60617, 16'd63544, 16'd51412, 16'd45552, 16'd44799, 16'd44702, 16'd28267, 16'd36578, 16'd22597, 16'd51609, 16'd29078, 16'd29893, 16'd12241, 16'd49103, 16'd49225, 16'd39907, 16'd61293, 16'd42104, 16'd45374, 16'd2, 16'd60579, 16'd60649, 16'd52480, 16'd20787});
	test_expansion(128'h09225f6d3ac67925085dd327c3ece826, {16'd46187, 16'd13376, 16'd17601, 16'd57209, 16'd14343, 16'd51344, 16'd17431, 16'd41193, 16'd10082, 16'd32193, 16'd18228, 16'd21347, 16'd50032, 16'd54213, 16'd24720, 16'd21249, 16'd30228, 16'd22777, 16'd41691, 16'd24331, 16'd32768, 16'd24586, 16'd11806, 16'd21895, 16'd10311, 16'd20808});
	test_expansion(128'hb01b43cc26a2b16fd46a3be995dd5659, {16'd33498, 16'd26664, 16'd3504, 16'd28256, 16'd679, 16'd1702, 16'd13634, 16'd63233, 16'd11532, 16'd51562, 16'd63874, 16'd34769, 16'd2503, 16'd56415, 16'd14114, 16'd26506, 16'd26013, 16'd52757, 16'd58189, 16'd45265, 16'd42279, 16'd32870, 16'd44502, 16'd26297, 16'd43830, 16'd17420});
	test_expansion(128'hf4c819bf60d731fd4db7cc0ed152dfe6, {16'd20379, 16'd10227, 16'd25206, 16'd34831, 16'd48382, 16'd49453, 16'd48611, 16'd62145, 16'd39634, 16'd25310, 16'd58937, 16'd41399, 16'd46068, 16'd56423, 16'd2978, 16'd48392, 16'd58385, 16'd29929, 16'd11647, 16'd51534, 16'd39759, 16'd23578, 16'd48292, 16'd3612, 16'd33479, 16'd11126});
	test_expansion(128'hdc2acd92ff67ef01004896c75454a927, {16'd60108, 16'd2798, 16'd44521, 16'd19780, 16'd49468, 16'd57716, 16'd14148, 16'd20415, 16'd27901, 16'd53696, 16'd19634, 16'd50975, 16'd24414, 16'd52752, 16'd2764, 16'd13070, 16'd11460, 16'd50674, 16'd38598, 16'd19522, 16'd62568, 16'd26467, 16'd7318, 16'd44581, 16'd21596, 16'd53645});
	test_expansion(128'hf05d8b0b7c99317f6fb981f7347b2c5c, {16'd52908, 16'd38548, 16'd29527, 16'd56489, 16'd45441, 16'd10565, 16'd36668, 16'd27991, 16'd110, 16'd56311, 16'd53257, 16'd3208, 16'd48789, 16'd29637, 16'd18748, 16'd36017, 16'd64966, 16'd60443, 16'd57169, 16'd15190, 16'd28144, 16'd46412, 16'd17758, 16'd44381, 16'd56790, 16'd4054});
	test_expansion(128'h99187a346bfef66bd76efea0f74d2c87, {16'd31963, 16'd17559, 16'd19154, 16'd14145, 16'd18837, 16'd24234, 16'd6983, 16'd42539, 16'd60417, 16'd34416, 16'd57223, 16'd35534, 16'd714, 16'd24881, 16'd56068, 16'd53201, 16'd10791, 16'd49257, 16'd59168, 16'd34943, 16'd17143, 16'd63362, 16'd8563, 16'd14150, 16'd38351, 16'd58771});
	test_expansion(128'h809676a9e0c2620c800269d8718f29ff, {16'd9594, 16'd16891, 16'd36674, 16'd63778, 16'd10507, 16'd13045, 16'd25234, 16'd58994, 16'd794, 16'd61979, 16'd40766, 16'd30526, 16'd60867, 16'd52237, 16'd63384, 16'd57037, 16'd7087, 16'd1235, 16'd41779, 16'd47164, 16'd58658, 16'd19640, 16'd25739, 16'd22768, 16'd60669, 16'd53933});
	test_expansion(128'h3f08a4acf2d82c7e85477425c0829c34, {16'd28458, 16'd341, 16'd38205, 16'd14129, 16'd28598, 16'd1136, 16'd342, 16'd56491, 16'd46800, 16'd10975, 16'd21748, 16'd47123, 16'd51460, 16'd6562, 16'd18608, 16'd61084, 16'd36946, 16'd30412, 16'd55723, 16'd47741, 16'd53945, 16'd44689, 16'd12260, 16'd62389, 16'd38644, 16'd55701});
	test_expansion(128'h17b59622271fe37870d6db9e777a95d3, {16'd51800, 16'd57596, 16'd51972, 16'd57041, 16'd49478, 16'd9265, 16'd22450, 16'd59947, 16'd34338, 16'd50959, 16'd55168, 16'd30763, 16'd37941, 16'd25925, 16'd45866, 16'd54104, 16'd18883, 16'd50157, 16'd25249, 16'd56815, 16'd6052, 16'd60146, 16'd28144, 16'd9510, 16'd26119, 16'd18842});
	test_expansion(128'h9761d0308d1f5c831bd5f92026a167c8, {16'd29876, 16'd20314, 16'd29637, 16'd53480, 16'd49146, 16'd36247, 16'd29065, 16'd1430, 16'd55338, 16'd61235, 16'd23334, 16'd17979, 16'd30867, 16'd55727, 16'd195, 16'd57919, 16'd57007, 16'd5670, 16'd52515, 16'd24212, 16'd48375, 16'd19117, 16'd28157, 16'd35438, 16'd14309, 16'd41748});
	test_expansion(128'h39ec776cf87b57a005630286107b9c5c, {16'd22383, 16'd4559, 16'd34918, 16'd1565, 16'd24856, 16'd61852, 16'd48563, 16'd2841, 16'd49676, 16'd34235, 16'd27734, 16'd9555, 16'd5522, 16'd62326, 16'd27634, 16'd15500, 16'd59891, 16'd583, 16'd27777, 16'd51469, 16'd57335, 16'd19261, 16'd6148, 16'd1141, 16'd49057, 16'd43711});
	test_expansion(128'h6c66441fe64d7af9a7fad74255d09b67, {16'd29660, 16'd41524, 16'd65128, 16'd13478, 16'd51799, 16'd28470, 16'd10979, 16'd31982, 16'd63167, 16'd39089, 16'd11989, 16'd36539, 16'd45301, 16'd64462, 16'd62570, 16'd43391, 16'd40042, 16'd48128, 16'd9043, 16'd39696, 16'd56343, 16'd27176, 16'd60345, 16'd20956, 16'd17735, 16'd40816});
	test_expansion(128'hbe14d91cc8385cfb6183d121f1be0c21, {16'd50000, 16'd799, 16'd42374, 16'd52914, 16'd29461, 16'd21877, 16'd17204, 16'd40546, 16'd2892, 16'd42073, 16'd7137, 16'd33004, 16'd26983, 16'd36759, 16'd10351, 16'd15446, 16'd5475, 16'd54053, 16'd54876, 16'd3187, 16'd25519, 16'd29427, 16'd25326, 16'd31130, 16'd63049, 16'd26207});
	test_expansion(128'he231e348f8132b9ee675fa7d9a0866a2, {16'd25112, 16'd38991, 16'd27878, 16'd9628, 16'd38561, 16'd17851, 16'd36389, 16'd4572, 16'd11580, 16'd316, 16'd11406, 16'd50086, 16'd42948, 16'd47650, 16'd34831, 16'd61302, 16'd1968, 16'd17629, 16'd30780, 16'd13271, 16'd65105, 16'd41415, 16'd37613, 16'd49619, 16'd34544, 16'd38202});
	test_expansion(128'hcc2019552bb77111e11c7d1dd506b33d, {16'd27813, 16'd56965, 16'd12057, 16'd13985, 16'd35771, 16'd16042, 16'd55841, 16'd10071, 16'd37789, 16'd64676, 16'd24852, 16'd55993, 16'd52393, 16'd5153, 16'd5864, 16'd50860, 16'd46546, 16'd59452, 16'd34443, 16'd44948, 16'd17701, 16'd10071, 16'd40697, 16'd982, 16'd21027, 16'd24117});
	test_expansion(128'he3bcf8c1ef25e466806f5ff125a91433, {16'd45294, 16'd21361, 16'd30893, 16'd47778, 16'd48058, 16'd52138, 16'd31183, 16'd49169, 16'd27073, 16'd51374, 16'd42178, 16'd44169, 16'd21426, 16'd29976, 16'd46848, 16'd45773, 16'd42488, 16'd37472, 16'd14465, 16'd10732, 16'd64894, 16'd53816, 16'd39324, 16'd17914, 16'd36953, 16'd49305});
	test_expansion(128'hf164532c4cf8ac46e33166be593234dd, {16'd28238, 16'd6982, 16'd40143, 16'd27931, 16'd52481, 16'd29273, 16'd60157, 16'd19172, 16'd50254, 16'd5946, 16'd63816, 16'd17964, 16'd40770, 16'd3113, 16'd3543, 16'd7028, 16'd38217, 16'd58652, 16'd39295, 16'd53248, 16'd32195, 16'd36315, 16'd49513, 16'd56906, 16'd26052, 16'd65046});
	test_expansion(128'hfac8b5b014b1b41b6a7c1938dc3aa7c7, {16'd15687, 16'd7884, 16'd13850, 16'd16280, 16'd57827, 16'd18503, 16'd45096, 16'd32299, 16'd24618, 16'd34196, 16'd11509, 16'd23262, 16'd53292, 16'd18677, 16'd28125, 16'd14118, 16'd20566, 16'd21533, 16'd24287, 16'd50979, 16'd58220, 16'd26235, 16'd7566, 16'd33082, 16'd33770, 16'd11812});
	test_expansion(128'h237ffde0fa7405cee385e71cf00dfc35, {16'd12960, 16'd17961, 16'd50128, 16'd43957, 16'd12881, 16'd45286, 16'd63633, 16'd54186, 16'd20716, 16'd3940, 16'd61435, 16'd47, 16'd15531, 16'd36579, 16'd20684, 16'd47147, 16'd7061, 16'd46142, 16'd14472, 16'd40409, 16'd4111, 16'd10984, 16'd35422, 16'd53659, 16'd29018, 16'd51772});
	test_expansion(128'hfc78bfd829a5e007d76473e57b33606c, {16'd26469, 16'd29631, 16'd6683, 16'd32874, 16'd57526, 16'd16548, 16'd60952, 16'd22743, 16'd31945, 16'd62935, 16'd59225, 16'd6607, 16'd2377, 16'd20615, 16'd45010, 16'd1114, 16'd58630, 16'd10792, 16'd39545, 16'd17151, 16'd15113, 16'd112, 16'd40926, 16'd53115, 16'd47947, 16'd53180});
	test_expansion(128'hdfa9e014e1e3623c3c62bcd86a5dea08, {16'd53276, 16'd35724, 16'd13698, 16'd5520, 16'd23219, 16'd46896, 16'd6216, 16'd58917, 16'd6030, 16'd56152, 16'd45914, 16'd1726, 16'd54313, 16'd53037, 16'd32342, 16'd54557, 16'd10707, 16'd616, 16'd40295, 16'd2311, 16'd12682, 16'd57428, 16'd23367, 16'd42040, 16'd6299, 16'd18762});
	test_expansion(128'h16f87a371761ec003a63b2627a6d56cd, {16'd52388, 16'd29859, 16'd14232, 16'd8558, 16'd51457, 16'd11089, 16'd27155, 16'd64947, 16'd1204, 16'd56950, 16'd25093, 16'd19113, 16'd175, 16'd2804, 16'd8189, 16'd305, 16'd53261, 16'd56517, 16'd34696, 16'd63662, 16'd46472, 16'd35894, 16'd7152, 16'd50141, 16'd40297, 16'd32311});
	test_expansion(128'h7284a946225634e9eba6b83e09702047, {16'd61227, 16'd3959, 16'd20694, 16'd11854, 16'd57635, 16'd3883, 16'd49996, 16'd26784, 16'd61878, 16'd40013, 16'd19630, 16'd23118, 16'd47993, 16'd3853, 16'd18543, 16'd25734, 16'd29272, 16'd10889, 16'd42276, 16'd49050, 16'd62220, 16'd65235, 16'd30981, 16'd316, 16'd23613, 16'd54797});
	test_expansion(128'hec51b68df139a8bc830ecd74b6d25094, {16'd9683, 16'd52745, 16'd4363, 16'd8852, 16'd45381, 16'd8435, 16'd4505, 16'd17205, 16'd36271, 16'd13537, 16'd7533, 16'd10095, 16'd65156, 16'd47208, 16'd3545, 16'd58003, 16'd19929, 16'd29797, 16'd23979, 16'd5947, 16'd24848, 16'd41824, 16'd18802, 16'd35636, 16'd57029, 16'd56371});
	test_expansion(128'h416e155ade6c9c896b36ed9137afc34e, {16'd47849, 16'd57526, 16'd51804, 16'd8251, 16'd27303, 16'd37446, 16'd15176, 16'd13315, 16'd44716, 16'd50657, 16'd65069, 16'd21808, 16'd1285, 16'd24150, 16'd56087, 16'd4595, 16'd6654, 16'd41768, 16'd35421, 16'd42996, 16'd62310, 16'd61202, 16'd54041, 16'd23477, 16'd53218, 16'd19499});
	test_expansion(128'h8a54de6115eefaa789c6c72acd800aea, {16'd38968, 16'd30683, 16'd33829, 16'd55427, 16'd35685, 16'd8027, 16'd33981, 16'd32646, 16'd52872, 16'd32481, 16'd41293, 16'd18949, 16'd23354, 16'd11179, 16'd18770, 16'd58586, 16'd38703, 16'd15102, 16'd42327, 16'd64220, 16'd56447, 16'd29257, 16'd17422, 16'd29487, 16'd1642, 16'd51594});
	test_expansion(128'h5cbe06d292a8438de7d849dda02c9699, {16'd24194, 16'd58938, 16'd63600, 16'd54337, 16'd2076, 16'd13554, 16'd49147, 16'd62042, 16'd41330, 16'd30512, 16'd19550, 16'd43899, 16'd28575, 16'd25785, 16'd56092, 16'd43094, 16'd1226, 16'd2189, 16'd1476, 16'd31473, 16'd36236, 16'd47718, 16'd11202, 16'd62280, 16'd16163, 16'd17471});
	test_expansion(128'hed59933c38c3ce819044eb003688fd4b, {16'd61038, 16'd47718, 16'd1982, 16'd60422, 16'd22927, 16'd35714, 16'd62367, 16'd42709, 16'd2369, 16'd48508, 16'd40243, 16'd8492, 16'd19543, 16'd42292, 16'd12693, 16'd13783, 16'd6730, 16'd16437, 16'd62016, 16'd45255, 16'd62112, 16'd2234, 16'd17874, 16'd6433, 16'd3818, 16'd20726});
	test_expansion(128'h235f84bd3b7c7206308745f6f9bbd03f, {16'd30291, 16'd55476, 16'd16775, 16'd24785, 16'd6133, 16'd14214, 16'd5023, 16'd40870, 16'd20532, 16'd6238, 16'd53480, 16'd266, 16'd27110, 16'd56058, 16'd37472, 16'd58363, 16'd12173, 16'd38967, 16'd10720, 16'd36510, 16'd58677, 16'd22530, 16'd8515, 16'd55913, 16'd3167, 16'd3666});
	test_expansion(128'h53bf5330e453ff6d6f5c42f25a465432, {16'd26506, 16'd42469, 16'd4160, 16'd25796, 16'd60877, 16'd18253, 16'd39124, 16'd16514, 16'd40679, 16'd28057, 16'd26562, 16'd11575, 16'd14432, 16'd2878, 16'd37933, 16'd42367, 16'd32607, 16'd15276, 16'd28740, 16'd18239, 16'd51468, 16'd14517, 16'd2970, 16'd50090, 16'd61796, 16'd58098});
	test_expansion(128'h8003ea056eb721506b5db4d37cf70c57, {16'd19160, 16'd40153, 16'd59733, 16'd29003, 16'd55931, 16'd28789, 16'd21913, 16'd11736, 16'd57266, 16'd26794, 16'd26944, 16'd21432, 16'd23599, 16'd62339, 16'd7612, 16'd25446, 16'd65489, 16'd44135, 16'd5974, 16'd33172, 16'd17290, 16'd35957, 16'd26487, 16'd4491, 16'd4570, 16'd8371});
	test_expansion(128'h36d20350331b489ba64bfd30544c4c3b, {16'd3873, 16'd2417, 16'd22846, 16'd50785, 16'd56604, 16'd38575, 16'd45760, 16'd24466, 16'd57140, 16'd4055, 16'd25138, 16'd61310, 16'd35742, 16'd48667, 16'd11131, 16'd33293, 16'd50815, 16'd55534, 16'd9373, 16'd26957, 16'd1054, 16'd10625, 16'd31115, 16'd64043, 16'd2764, 16'd59564});
	test_expansion(128'h61f588e6b53843938aaa29ec11d05165, {16'd10436, 16'd53643, 16'd64147, 16'd10582, 16'd58912, 16'd36036, 16'd14095, 16'd40203, 16'd2549, 16'd61101, 16'd56239, 16'd44768, 16'd43384, 16'd36201, 16'd43795, 16'd31380, 16'd55351, 16'd10809, 16'd9012, 16'd28704, 16'd28873, 16'd38650, 16'd58666, 16'd4156, 16'd37372, 16'd45509});
	test_expansion(128'ha600a8b1a41f7c2fb44889714b22b2d5, {16'd22874, 16'd15911, 16'd34429, 16'd25778, 16'd52111, 16'd19939, 16'd41437, 16'd6421, 16'd12930, 16'd10096, 16'd49704, 16'd26352, 16'd62113, 16'd64754, 16'd280, 16'd55029, 16'd46103, 16'd50328, 16'd4784, 16'd5464, 16'd8766, 16'd32570, 16'd61806, 16'd31360, 16'd7271, 16'd19165});
	test_expansion(128'h37a322e6c1c3ecc5b4ae672230950bed, {16'd11922, 16'd9308, 16'd45119, 16'd8383, 16'd33325, 16'd5189, 16'd6098, 16'd10410, 16'd52830, 16'd383, 16'd13396, 16'd15307, 16'd60248, 16'd34833, 16'd42328, 16'd24243, 16'd3149, 16'd63137, 16'd56711, 16'd1184, 16'd46616, 16'd52727, 16'd51435, 16'd34209, 16'd13780, 16'd29729});
	test_expansion(128'h5afab401a2a2b51274ddaa129b056fa4, {16'd25263, 16'd27913, 16'd58982, 16'd16427, 16'd45689, 16'd31380, 16'd46148, 16'd60868, 16'd12909, 16'd15986, 16'd40061, 16'd13883, 16'd63898, 16'd27224, 16'd32130, 16'd30179, 16'd43853, 16'd23988, 16'd37896, 16'd5921, 16'd15395, 16'd20700, 16'd34005, 16'd35100, 16'd40153, 16'd17200});
	test_expansion(128'h6c2087768ffe4d769e6a743284428332, {16'd44080, 16'd37822, 16'd42055, 16'd4181, 16'd49681, 16'd6689, 16'd42840, 16'd34646, 16'd28914, 16'd49189, 16'd4715, 16'd56577, 16'd34547, 16'd63177, 16'd45578, 16'd23493, 16'd5282, 16'd64550, 16'd689, 16'd61204, 16'd52950, 16'd62575, 16'd50415, 16'd3351, 16'd44933, 16'd63854});
	test_expansion(128'hd23b09087237dd9aa234238b29e07a14, {16'd63801, 16'd56356, 16'd54407, 16'd19482, 16'd602, 16'd25358, 16'd20171, 16'd31661, 16'd54183, 16'd19758, 16'd49430, 16'd829, 16'd33728, 16'd33030, 16'd7821, 16'd14559, 16'd16148, 16'd29778, 16'd37839, 16'd26430, 16'd29604, 16'd38102, 16'd36014, 16'd32383, 16'd19523, 16'd52802});
	test_expansion(128'hf4e8f08c877a6816ce95c79e95c40d85, {16'd22571, 16'd54539, 16'd50480, 16'd8591, 16'd40526, 16'd63279, 16'd62376, 16'd44827, 16'd25642, 16'd59414, 16'd51302, 16'd6802, 16'd4724, 16'd57239, 16'd24141, 16'd9254, 16'd25469, 16'd46797, 16'd39237, 16'd45099, 16'd39860, 16'd37655, 16'd3122, 16'd13157, 16'd39554, 16'd17951});
	test_expansion(128'hca24296edce55e11fc9414e2d4f02261, {16'd5197, 16'd56253, 16'd47357, 16'd4727, 16'd36964, 16'd54611, 16'd47955, 16'd31659, 16'd14181, 16'd36009, 16'd26067, 16'd53915, 16'd25235, 16'd10009, 16'd41589, 16'd11663, 16'd8866, 16'd38339, 16'd34855, 16'd64909, 16'd45001, 16'd15410, 16'd5485, 16'd54777, 16'd26922, 16'd22369});
	test_expansion(128'h6de016c42212ff702dc7781535e11925, {16'd41935, 16'd182, 16'd9805, 16'd33630, 16'd27723, 16'd10709, 16'd17868, 16'd31130, 16'd22449, 16'd14420, 16'd16397, 16'd41016, 16'd45713, 16'd765, 16'd54709, 16'd19636, 16'd28802, 16'd44028, 16'd62746, 16'd54898, 16'd5736, 16'd39895, 16'd60947, 16'd42895, 16'd64066, 16'd6041});
	test_expansion(128'hef6e06802a7ea70e9ac105ffa139ec99, {16'd32995, 16'd26968, 16'd12345, 16'd30591, 16'd60855, 16'd19882, 16'd29302, 16'd16390, 16'd49523, 16'd38979, 16'd9693, 16'd5663, 16'd32734, 16'd65470, 16'd54928, 16'd26638, 16'd26670, 16'd59727, 16'd42759, 16'd50431, 16'd31418, 16'd46482, 16'd41911, 16'd14058, 16'd13060, 16'd58952});
	test_expansion(128'h063940b6830924314ac4e99853799f8b, {16'd30773, 16'd64534, 16'd10984, 16'd51906, 16'd41600, 16'd25624, 16'd54157, 16'd55767, 16'd11061, 16'd22403, 16'd46486, 16'd10017, 16'd41583, 16'd25077, 16'd59871, 16'd36225, 16'd38051, 16'd27076, 16'd6340, 16'd25914, 16'd45049, 16'd47659, 16'd42630, 16'd36245, 16'd21421, 16'd51764});
	test_expansion(128'hc91e3665d7f4f9e07ee9688b47aa62a3, {16'd47888, 16'd2505, 16'd57803, 16'd49522, 16'd38892, 16'd2967, 16'd7486, 16'd4714, 16'd55502, 16'd18739, 16'd3346, 16'd13545, 16'd38801, 16'd3832, 16'd40064, 16'd9655, 16'd31229, 16'd26226, 16'd4429, 16'd38850, 16'd61193, 16'd4781, 16'd42781, 16'd36064, 16'd44707, 16'd46665});
	test_expansion(128'h03617f0e15a59872958ce25b753f10cb, {16'd63000, 16'd23574, 16'd64050, 16'd15185, 16'd3941, 16'd63533, 16'd7049, 16'd21184, 16'd27796, 16'd59857, 16'd3942, 16'd24624, 16'd21305, 16'd19119, 16'd49018, 16'd1856, 16'd12627, 16'd23179, 16'd13268, 16'd54317, 16'd23053, 16'd8732, 16'd54812, 16'd3537, 16'd60750, 16'd47612});
	test_expansion(128'h1e1a4913572842baab45a436bfea7b8e, {16'd54451, 16'd6806, 16'd10849, 16'd18871, 16'd24361, 16'd57052, 16'd18252, 16'd12811, 16'd53707, 16'd14651, 16'd45116, 16'd3049, 16'd48026, 16'd65495, 16'd20447, 16'd55815, 16'd4654, 16'd37903, 16'd14487, 16'd63258, 16'd58956, 16'd29859, 16'd59002, 16'd52471, 16'd2950, 16'd56548});
	test_expansion(128'he4a76d7ecbe6977cd0fd89270e6e498b, {16'd9402, 16'd28776, 16'd34906, 16'd23618, 16'd42914, 16'd59719, 16'd63658, 16'd43396, 16'd19594, 16'd14664, 16'd52811, 16'd19026, 16'd14564, 16'd58360, 16'd43287, 16'd30759, 16'd32878, 16'd33646, 16'd15102, 16'd49956, 16'd32670, 16'd36686, 16'd32871, 16'd22730, 16'd11146, 16'd63423});
	test_expansion(128'hd5819341fdd6b831dad08aa9bddbd734, {16'd60981, 16'd32008, 16'd62954, 16'd45785, 16'd41345, 16'd22037, 16'd3909, 16'd46539, 16'd39413, 16'd3465, 16'd53497, 16'd12470, 16'd16681, 16'd17227, 16'd50699, 16'd40920, 16'd31630, 16'd11178, 16'd15932, 16'd48205, 16'd10612, 16'd61868, 16'd3915, 16'd45571, 16'd38940, 16'd19895});
	test_expansion(128'h9496127b93b19ae0f8e2290ace05e6a6, {16'd30537, 16'd33004, 16'd64827, 16'd42953, 16'd43848, 16'd59061, 16'd55723, 16'd31773, 16'd270, 16'd3961, 16'd57089, 16'd33525, 16'd50888, 16'd58261, 16'd59716, 16'd7696, 16'd44861, 16'd22253, 16'd12522, 16'd15550, 16'd14813, 16'd33127, 16'd17002, 16'd836, 16'd25874, 16'd16925});
	test_expansion(128'hf8134407a7e6a1fa881a3d58a7698f5b, {16'd52385, 16'd35024, 16'd37739, 16'd23588, 16'd30763, 16'd55801, 16'd6643, 16'd59143, 16'd31805, 16'd8505, 16'd18494, 16'd25993, 16'd13294, 16'd47859, 16'd47933, 16'd10383, 16'd24663, 16'd9829, 16'd24774, 16'd28114, 16'd2704, 16'd7850, 16'd59874, 16'd63478, 16'd20806, 16'd18272});
	test_expansion(128'h805ebacd19879abc9e73894ebedcba5a, {16'd16449, 16'd61875, 16'd49992, 16'd31250, 16'd2179, 16'd47433, 16'd48758, 16'd61428, 16'd12206, 16'd61585, 16'd2247, 16'd45451, 16'd37309, 16'd28117, 16'd46497, 16'd48115, 16'd63845, 16'd49613, 16'd53388, 16'd22196, 16'd55204, 16'd3001, 16'd43261, 16'd2769, 16'd63838, 16'd8801});
	test_expansion(128'hdde6a60f2e3223c3fdcb3e79d8c9d9b2, {16'd42984, 16'd42010, 16'd33888, 16'd35146, 16'd42525, 16'd22940, 16'd20220, 16'd37275, 16'd37931, 16'd2971, 16'd38097, 16'd17788, 16'd18740, 16'd53485, 16'd2092, 16'd46186, 16'd56639, 16'd51832, 16'd2993, 16'd57984, 16'd34714, 16'd55993, 16'd55825, 16'd60835, 16'd4647, 16'd38859});
	test_expansion(128'hec577d6676de847f434930710c5d758a, {16'd27067, 16'd37530, 16'd37545, 16'd45623, 16'd32507, 16'd21398, 16'd3787, 16'd37559, 16'd18103, 16'd28070, 16'd6310, 16'd62619, 16'd119, 16'd17202, 16'd46000, 16'd55260, 16'd23494, 16'd5124, 16'd48712, 16'd61478, 16'd11990, 16'd36213, 16'd43644, 16'd13204, 16'd37006, 16'd850});
	test_expansion(128'h11168d27fa56780e8f74a7250235f5b4, {16'd19505, 16'd4360, 16'd43509, 16'd58720, 16'd36865, 16'd6956, 16'd27134, 16'd12951, 16'd51332, 16'd8357, 16'd57051, 16'd16196, 16'd13302, 16'd8903, 16'd58034, 16'd36769, 16'd45294, 16'd3684, 16'd47586, 16'd9163, 16'd32965, 16'd51242, 16'd4696, 16'd3476, 16'd53941, 16'd20876});
	test_expansion(128'h0edf3a6c91369ac11a7632a03ebb9f5f, {16'd23101, 16'd40964, 16'd46229, 16'd45621, 16'd49027, 16'd51226, 16'd11423, 16'd23159, 16'd62796, 16'd62563, 16'd22256, 16'd10020, 16'd17895, 16'd51596, 16'd64705, 16'd57770, 16'd36644, 16'd20564, 16'd40840, 16'd57656, 16'd52788, 16'd32480, 16'd15949, 16'd44795, 16'd61259, 16'd19540});
	test_expansion(128'h97cc9ac5ffce39c3a5734dafa7606776, {16'd50409, 16'd42712, 16'd65034, 16'd1094, 16'd46461, 16'd1532, 16'd51780, 16'd19467, 16'd21400, 16'd47559, 16'd62691, 16'd25802, 16'd25924, 16'd59468, 16'd64404, 16'd53605, 16'd63893, 16'd52762, 16'd2763, 16'd48386, 16'd19065, 16'd3461, 16'd64565, 16'd6761, 16'd25104, 16'd44841});
	test_expansion(128'h751ff22d55670f7d202aa3df45167601, {16'd14510, 16'd52513, 16'd46127, 16'd24596, 16'd6885, 16'd20201, 16'd56371, 16'd10768, 16'd44772, 16'd51875, 16'd26251, 16'd62654, 16'd38251, 16'd47403, 16'd33962, 16'd57629, 16'd5793, 16'd1772, 16'd12412, 16'd27878, 16'd3374, 16'd42372, 16'd59416, 16'd30772, 16'd42737, 16'd5653});
	test_expansion(128'hee79a2a90b97822e0a585b0d063915a7, {16'd43869, 16'd55161, 16'd11380, 16'd29333, 16'd27054, 16'd30170, 16'd831, 16'd56919, 16'd61721, 16'd53902, 16'd26197, 16'd55979, 16'd13339, 16'd14073, 16'd22031, 16'd30332, 16'd32774, 16'd36132, 16'd31786, 16'd36568, 16'd22609, 16'd28037, 16'd33177, 16'd42712, 16'd26561, 16'd9185});
	test_expansion(128'hecc41016517a17fed9fe6b8d1d668318, {16'd57743, 16'd13920, 16'd23036, 16'd42478, 16'd10488, 16'd49970, 16'd41246, 16'd45892, 16'd47699, 16'd20179, 16'd1443, 16'd47564, 16'd50996, 16'd23530, 16'd18599, 16'd21941, 16'd12232, 16'd18366, 16'd18807, 16'd28052, 16'd19400, 16'd30485, 16'd30126, 16'd16834, 16'd2713, 16'd54326});
	test_expansion(128'he4a1ad4d7a749bcc6ee5f7a73a8e2b94, {16'd10503, 16'd3797, 16'd44327, 16'd59980, 16'd58051, 16'd47669, 16'd48290, 16'd9051, 16'd59753, 16'd39049, 16'd55318, 16'd58223, 16'd18817, 16'd48094, 16'd18585, 16'd61970, 16'd61549, 16'd56973, 16'd47456, 16'd61690, 16'd33, 16'd63945, 16'd37456, 16'd1936, 16'd32319, 16'd50382});
	test_expansion(128'hffb96b0ce00cb69cc1c84238604d1640, {16'd54699, 16'd2913, 16'd7031, 16'd53027, 16'd2683, 16'd51059, 16'd10258, 16'd2368, 16'd28720, 16'd62734, 16'd56043, 16'd4913, 16'd56851, 16'd64740, 16'd62898, 16'd7628, 16'd15909, 16'd57723, 16'd11795, 16'd57064, 16'd2110, 16'd12419, 16'd65441, 16'd52464, 16'd5030, 16'd59190});
	test_expansion(128'h07c9f6ce6f02ac76e19438191f902ed1, {16'd31551, 16'd62866, 16'd5582, 16'd12794, 16'd46099, 16'd48622, 16'd37613, 16'd8127, 16'd23986, 16'd26759, 16'd33296, 16'd40664, 16'd53524, 16'd50627, 16'd50189, 16'd32574, 16'd19726, 16'd63114, 16'd51466, 16'd28167, 16'd21169, 16'd26201, 16'd5386, 16'd20181, 16'd16790, 16'd35841});
	test_expansion(128'hfe06895ddc6f192b08d8c94fb61eac84, {16'd31286, 16'd58123, 16'd49476, 16'd447, 16'd10994, 16'd19134, 16'd24423, 16'd45872, 16'd58678, 16'd4445, 16'd27934, 16'd27788, 16'd63291, 16'd63908, 16'd38683, 16'd40162, 16'd11964, 16'd45286, 16'd11861, 16'd38846, 16'd49370, 16'd8119, 16'd59355, 16'd20417, 16'd47749, 16'd32898});
	test_expansion(128'h53ce2ad98fd3c8bd21fc6b1b95d74bfc, {16'd42369, 16'd29318, 16'd2914, 16'd42951, 16'd21973, 16'd10127, 16'd34812, 16'd48978, 16'd51032, 16'd47694, 16'd36123, 16'd47554, 16'd29637, 16'd19258, 16'd24221, 16'd6838, 16'd44339, 16'd39142, 16'd60692, 16'd45727, 16'd53298, 16'd36989, 16'd56949, 16'd48535, 16'd6834, 16'd48048});
	test_expansion(128'h6f787c6a427b9e996d0c83526ffbbd3d, {16'd40995, 16'd62230, 16'd30007, 16'd56717, 16'd49964, 16'd54096, 16'd12649, 16'd63079, 16'd24035, 16'd25581, 16'd26932, 16'd51264, 16'd21122, 16'd48560, 16'd10900, 16'd57226, 16'd33871, 16'd55125, 16'd65347, 16'd13949, 16'd30448, 16'd58782, 16'd4749, 16'd2153, 16'd61846, 16'd59409});
	test_expansion(128'h9a17b2cc8863da6138ba99638b92a1d5, {16'd33608, 16'd46848, 16'd2036, 16'd20415, 16'd39228, 16'd7456, 16'd42401, 16'd34839, 16'd14566, 16'd35269, 16'd30590, 16'd32036, 16'd8279, 16'd20636, 16'd43669, 16'd16277, 16'd60219, 16'd12191, 16'd61033, 16'd10715, 16'd8511, 16'd27250, 16'd35834, 16'd49061, 16'd25649, 16'd55638});
	test_expansion(128'he3a5f7085224b16058fe2caedc67efbf, {16'd25663, 16'd62059, 16'd53263, 16'd3954, 16'd60377, 16'd17360, 16'd33577, 16'd3237, 16'd49164, 16'd18318, 16'd6937, 16'd60662, 16'd14560, 16'd4374, 16'd53440, 16'd59066, 16'd30376, 16'd49365, 16'd65422, 16'd28391, 16'd26429, 16'd2150, 16'd12134, 16'd33994, 16'd13268, 16'd13711});
	test_expansion(128'h4c3613cc93979ab7b01622a4748a1d5c, {16'd56407, 16'd34657, 16'd3272, 16'd24781, 16'd51986, 16'd7607, 16'd9241, 16'd60874, 16'd13156, 16'd41255, 16'd48743, 16'd58663, 16'd10896, 16'd1764, 16'd24511, 16'd60435, 16'd19068, 16'd36545, 16'd50506, 16'd107, 16'd30728, 16'd31604, 16'd8768, 16'd1739, 16'd36263, 16'd26466});
	test_expansion(128'hb716353b6842d4e3de711a21432b8299, {16'd41091, 16'd63703, 16'd58704, 16'd20651, 16'd15971, 16'd60788, 16'd30585, 16'd19853, 16'd63308, 16'd59351, 16'd47721, 16'd17895, 16'd8359, 16'd38333, 16'd18470, 16'd60420, 16'd40116, 16'd7269, 16'd21915, 16'd45132, 16'd11503, 16'd64704, 16'd62940, 16'd65170, 16'd17243, 16'd14992});
	test_expansion(128'hbabed485c98eb29997adb7063e05fd35, {16'd51367, 16'd57629, 16'd58056, 16'd19339, 16'd27586, 16'd24239, 16'd12403, 16'd46676, 16'd37563, 16'd34438, 16'd32224, 16'd1364, 16'd12624, 16'd18622, 16'd40395, 16'd8218, 16'd19532, 16'd57230, 16'd58643, 16'd50006, 16'd15566, 16'd18633, 16'd23424, 16'd7499, 16'd6859, 16'd46563});
	test_expansion(128'ha8bd70a9a22ca4920dfd73579babd29a, {16'd16712, 16'd32794, 16'd38801, 16'd22559, 16'd26072, 16'd35569, 16'd50942, 16'd8344, 16'd33927, 16'd57497, 16'd10377, 16'd41615, 16'd17735, 16'd40906, 16'd18791, 16'd29074, 16'd36816, 16'd37457, 16'd58572, 16'd5290, 16'd34545, 16'd24468, 16'd27634, 16'd25938, 16'd54024, 16'd41302});
	test_expansion(128'ha833023aaa0a42d50e2a01cdda32c642, {16'd55932, 16'd31451, 16'd38625, 16'd3989, 16'd30131, 16'd55901, 16'd29279, 16'd56400, 16'd8963, 16'd63239, 16'd47502, 16'd5285, 16'd22473, 16'd28103, 16'd54433, 16'd36739, 16'd56750, 16'd35634, 16'd26980, 16'd15237, 16'd62695, 16'd10359, 16'd1402, 16'd20668, 16'd15728, 16'd24635});
	test_expansion(128'h770ac624974428caf7d62d315f1c379f, {16'd30752, 16'd38162, 16'd57477, 16'd29129, 16'd10661, 16'd5318, 16'd30580, 16'd59035, 16'd11678, 16'd45447, 16'd28262, 16'd33656, 16'd12336, 16'd37932, 16'd39208, 16'd48971, 16'd36530, 16'd29837, 16'd19891, 16'd39257, 16'd29580, 16'd39730, 16'd23796, 16'd28453, 16'd27239, 16'd29131});
	test_expansion(128'h7f4d7f0113a5f4be789501c0337e5e50, {16'd32436, 16'd59887, 16'd4266, 16'd18213, 16'd59444, 16'd49695, 16'd15130, 16'd10931, 16'd36514, 16'd19569, 16'd46940, 16'd15011, 16'd39862, 16'd24893, 16'd36624, 16'd61610, 16'd44620, 16'd57454, 16'd61901, 16'd26942, 16'd13339, 16'd15440, 16'd55405, 16'd13628, 16'd18943, 16'd22908});
	test_expansion(128'h1fd0839e9b71d6831d23105f56dad4ad, {16'd10326, 16'd51714, 16'd39882, 16'd52304, 16'd30404, 16'd62028, 16'd56392, 16'd61954, 16'd9784, 16'd43636, 16'd15048, 16'd64606, 16'd15349, 16'd52804, 16'd32860, 16'd33872, 16'd50682, 16'd57463, 16'd45235, 16'd9012, 16'd2076, 16'd12504, 16'd48430, 16'd64764, 16'd52152, 16'd25189});
	test_expansion(128'h1d5de91c3b21ce857f23c515214f5ac9, {16'd46223, 16'd44348, 16'd14773, 16'd58440, 16'd16263, 16'd28283, 16'd51215, 16'd20628, 16'd1460, 16'd10575, 16'd42596, 16'd58257, 16'd18696, 16'd50047, 16'd2509, 16'd20667, 16'd45127, 16'd14751, 16'd27021, 16'd41748, 16'd23900, 16'd64636, 16'd63181, 16'd17370, 16'd20377, 16'd6856});
	test_expansion(128'hb38df384eb9197adc93253fb55cbb843, {16'd27861, 16'd11374, 16'd14914, 16'd31623, 16'd46476, 16'd57109, 16'd48010, 16'd51526, 16'd49837, 16'd45815, 16'd23051, 16'd16222, 16'd630, 16'd61822, 16'd9473, 16'd13001, 16'd40540, 16'd53418, 16'd24815, 16'd15516, 16'd39409, 16'd2904, 16'd17, 16'd52998, 16'd59975, 16'd20994});
	test_expansion(128'h702d090b2c043b7502810063e74ce751, {16'd11208, 16'd18782, 16'd30156, 16'd13794, 16'd53485, 16'd64226, 16'd2899, 16'd4030, 16'd23752, 16'd46175, 16'd18230, 16'd43084, 16'd56895, 16'd40531, 16'd2978, 16'd31302, 16'd23112, 16'd8702, 16'd18220, 16'd7643, 16'd58965, 16'd53447, 16'd60024, 16'd45186, 16'd28862, 16'd61199});
	test_expansion(128'h40bbdbcddb8b07ea7b05a07cb856abd6, {16'd37229, 16'd10203, 16'd4225, 16'd27739, 16'd37661, 16'd60646, 16'd44123, 16'd21164, 16'd46311, 16'd18280, 16'd62551, 16'd36538, 16'd54685, 16'd47688, 16'd5520, 16'd40776, 16'd64144, 16'd60872, 16'd29240, 16'd52437, 16'd36740, 16'd46212, 16'd33878, 16'd34958, 16'd20797, 16'd58400});
	test_expansion(128'he2a584c18b951122e7adb74cd2a945b7, {16'd473, 16'd48231, 16'd28951, 16'd40869, 16'd65137, 16'd58578, 16'd61787, 16'd32791, 16'd40902, 16'd27560, 16'd7246, 16'd5635, 16'd1691, 16'd24204, 16'd62045, 16'd21245, 16'd58934, 16'd34763, 16'd54966, 16'd12132, 16'd56123, 16'd27003, 16'd795, 16'd14025, 16'd26749, 16'd40702});
	test_expansion(128'h1e5e2c3da681c7469dfa65516aa21cff, {16'd47324, 16'd13840, 16'd10626, 16'd18439, 16'd21064, 16'd13971, 16'd20469, 16'd21620, 16'd24604, 16'd47565, 16'd35453, 16'd49478, 16'd52024, 16'd31432, 16'd33167, 16'd22582, 16'd4, 16'd34318, 16'd22734, 16'd19313, 16'd39367, 16'd33205, 16'd8142, 16'd41158, 16'd62515, 16'd46170});
	test_expansion(128'h7ca2ec24af3aca4f9f42d4b3fcd2f0fd, {16'd64836, 16'd25034, 16'd44913, 16'd54784, 16'd12315, 16'd54689, 16'd12888, 16'd28859, 16'd21643, 16'd2630, 16'd58983, 16'd35674, 16'd36913, 16'd22901, 16'd35319, 16'd2254, 16'd8582, 16'd60987, 16'd33226, 16'd5252, 16'd24191, 16'd37907, 16'd47100, 16'd35592, 16'd43402, 16'd53368});
	test_expansion(128'h3e126ea357ef57c1eb36f055312c16b1, {16'd3751, 16'd41147, 16'd44656, 16'd43922, 16'd22611, 16'd36866, 16'd15204, 16'd62432, 16'd5768, 16'd64841, 16'd25321, 16'd1080, 16'd57655, 16'd47526, 16'd9649, 16'd22343, 16'd32306, 16'd49726, 16'd63770, 16'd57379, 16'd17910, 16'd46354, 16'd57836, 16'd43499, 16'd21677, 16'd9612});
	test_expansion(128'h5c0dc2d05a886358f0452f5c12eeb31e, {16'd3551, 16'd61524, 16'd26055, 16'd44386, 16'd28227, 16'd48600, 16'd60573, 16'd57733, 16'd43021, 16'd35039, 16'd63017, 16'd48796, 16'd14453, 16'd56578, 16'd20613, 16'd64911, 16'd55868, 16'd49101, 16'd13938, 16'd14853, 16'd5081, 16'd17969, 16'd46023, 16'd24852, 16'd3128, 16'd24385});
	test_expansion(128'h46700475c7a80178137151c047aa2283, {16'd40223, 16'd48795, 16'd48956, 16'd56250, 16'd35883, 16'd3615, 16'd30710, 16'd6695, 16'd42178, 16'd50506, 16'd10916, 16'd9219, 16'd64225, 16'd55479, 16'd35080, 16'd32460, 16'd33485, 16'd53662, 16'd42534, 16'd27796, 16'd43795, 16'd7444, 16'd14666, 16'd19276, 16'd5165, 16'd45334});
	test_expansion(128'he9381037a1324f59df266777fac294fa, {16'd35884, 16'd55314, 16'd35739, 16'd36453, 16'd61424, 16'd23620, 16'd44308, 16'd2915, 16'd30415, 16'd20766, 16'd15824, 16'd48574, 16'd32556, 16'd26267, 16'd41066, 16'd43707, 16'd3630, 16'd43761, 16'd32411, 16'd58214, 16'd30125, 16'd29290, 16'd978, 16'd21553, 16'd31063, 16'd54708});
	test_expansion(128'hf1ff205e1f1d0d2a0b6e6355b6b3efb3, {16'd36503, 16'd50294, 16'd57521, 16'd49535, 16'd59104, 16'd6023, 16'd28152, 16'd8813, 16'd2734, 16'd28305, 16'd14356, 16'd33581, 16'd63253, 16'd16883, 16'd63449, 16'd19686, 16'd44923, 16'd60654, 16'd57344, 16'd13374, 16'd16196, 16'd4361, 16'd23314, 16'd15612, 16'd52883, 16'd19811});
	test_expansion(128'h47ed98f5f6b5a268fb009815048ec211, {16'd21713, 16'd32793, 16'd13626, 16'd63095, 16'd57611, 16'd6892, 16'd50331, 16'd32573, 16'd52923, 16'd14208, 16'd49090, 16'd57967, 16'd1777, 16'd40867, 16'd12621, 16'd15392, 16'd12295, 16'd5680, 16'd45062, 16'd65132, 16'd49530, 16'd50075, 16'd21237, 16'd217, 16'd18534, 16'd2237});
	test_expansion(128'h12f08975bcf90088e5f85d6c22c69a76, {16'd38783, 16'd31951, 16'd35907, 16'd10534, 16'd8238, 16'd43192, 16'd24906, 16'd23718, 16'd33605, 16'd15652, 16'd54616, 16'd9133, 16'd42238, 16'd42797, 16'd54621, 16'd38321, 16'd50978, 16'd19873, 16'd17036, 16'd47145, 16'd55557, 16'd20100, 16'd32061, 16'd25453, 16'd2574, 16'd5886});
	test_expansion(128'h8af8a65af6fa483d4de580fefa3e3a08, {16'd2087, 16'd29109, 16'd63447, 16'd9162, 16'd53159, 16'd25587, 16'd37718, 16'd18802, 16'd41860, 16'd33671, 16'd8416, 16'd2276, 16'd57395, 16'd49205, 16'd14187, 16'd47413, 16'd63840, 16'd63415, 16'd13785, 16'd511, 16'd39192, 16'd20538, 16'd54737, 16'd3272, 16'd28671, 16'd50176});
	test_expansion(128'h388e4e2bc9c332911f2c9f3541a4c659, {16'd15288, 16'd41994, 16'd18067, 16'd36692, 16'd4840, 16'd28125, 16'd54491, 16'd45087, 16'd51121, 16'd56492, 16'd49956, 16'd2051, 16'd61854, 16'd20145, 16'd4861, 16'd1178, 16'd64719, 16'd26861, 16'd27856, 16'd22247, 16'd571, 16'd54412, 16'd54924, 16'd15240, 16'd481, 16'd25733});
	test_expansion(128'h4df8cbb7bbb82efe2c3ff9dc1394256b, {16'd61126, 16'd53635, 16'd5902, 16'd63115, 16'd40652, 16'd21252, 16'd27037, 16'd45198, 16'd62953, 16'd63356, 16'd27937, 16'd50085, 16'd30957, 16'd32187, 16'd16588, 16'd58404, 16'd6828, 16'd58098, 16'd59055, 16'd36612, 16'd683, 16'd34353, 16'd57421, 16'd3325, 16'd33356, 16'd49877});
	test_expansion(128'hb801b21b7647ec0fd00c6732efacb74b, {16'd64803, 16'd64826, 16'd21187, 16'd20307, 16'd64020, 16'd13029, 16'd8058, 16'd4710, 16'd48369, 16'd56153, 16'd40981, 16'd6261, 16'd9226, 16'd56885, 16'd15065, 16'd43086, 16'd13142, 16'd22470, 16'd38403, 16'd56677, 16'd8926, 16'd34194, 16'd13745, 16'd2254, 16'd29889, 16'd19952});
	test_expansion(128'h4b813986bad13697e33f594a28012101, {16'd18872, 16'd32212, 16'd1458, 16'd20777, 16'd21861, 16'd25891, 16'd51054, 16'd25467, 16'd36273, 16'd4591, 16'd7918, 16'd62642, 16'd42379, 16'd35461, 16'd8949, 16'd42441, 16'd32404, 16'd9412, 16'd42732, 16'd50251, 16'd46627, 16'd15552, 16'd33834, 16'd51517, 16'd53950, 16'd21479});
	test_expansion(128'had744a6329ebdab019b89b6ff2aa718f, {16'd64461, 16'd49219, 16'd24887, 16'd16320, 16'd56933, 16'd21588, 16'd64648, 16'd54377, 16'd24951, 16'd46337, 16'd17618, 16'd47062, 16'd16802, 16'd55172, 16'd49838, 16'd8622, 16'd58917, 16'd43687, 16'd33133, 16'd31483, 16'd42011, 16'd12373, 16'd29964, 16'd29254, 16'd46623, 16'd43559});
	test_expansion(128'hba54d02eed4ed81d87e1f1eca124d74e, {16'd44919, 16'd47667, 16'd31213, 16'd37984, 16'd7209, 16'd41109, 16'd49634, 16'd31309, 16'd15379, 16'd18695, 16'd61663, 16'd55175, 16'd33508, 16'd14987, 16'd64447, 16'd59110, 16'd52145, 16'd28022, 16'd56915, 16'd53617, 16'd60577, 16'd48327, 16'd1495, 16'd63958, 16'd19703, 16'd41056});
	test_expansion(128'h4d3c09f232bc08dac6a5a6bb1f11c230, {16'd63305, 16'd5257, 16'd58798, 16'd5948, 16'd42113, 16'd11037, 16'd9636, 16'd24611, 16'd44356, 16'd22679, 16'd27978, 16'd19230, 16'd9527, 16'd53669, 16'd5768, 16'd33912, 16'd27335, 16'd60089, 16'd60930, 16'd63966, 16'd746, 16'd31279, 16'd33454, 16'd21693, 16'd12602, 16'd18840});
	test_expansion(128'h620e12e2108ae8d735060e7441cd597a, {16'd44447, 16'd29582, 16'd50756, 16'd61399, 16'd43360, 16'd42132, 16'd34583, 16'd15859, 16'd51756, 16'd11666, 16'd36859, 16'd22824, 16'd36306, 16'd48071, 16'd32808, 16'd51688, 16'd37195, 16'd61255, 16'd60684, 16'd51632, 16'd9162, 16'd37116, 16'd14943, 16'd38823, 16'd56923, 16'd53813});
	test_expansion(128'h042e844fb7c42671f5ca2e6e8de133d3, {16'd6030, 16'd27795, 16'd49903, 16'd41633, 16'd12067, 16'd57242, 16'd60422, 16'd27803, 16'd45398, 16'd52905, 16'd29941, 16'd32639, 16'd19500, 16'd50635, 16'd46431, 16'd33317, 16'd39636, 16'd62446, 16'd25203, 16'd39776, 16'd13777, 16'd61316, 16'd5249, 16'd18959, 16'd19189, 16'd24595});
	test_expansion(128'hf102396263b44d2bf798db8cd694f7a3, {16'd56021, 16'd15512, 16'd16570, 16'd60707, 16'd21550, 16'd13988, 16'd43640, 16'd32802, 16'd6861, 16'd58490, 16'd37937, 16'd57736, 16'd1748, 16'd5562, 16'd17945, 16'd62478, 16'd41429, 16'd63247, 16'd55831, 16'd6304, 16'd43601, 16'd62508, 16'd16200, 16'd36982, 16'd3634, 16'd61324});
	test_expansion(128'hc3c6075a1d03ae64fcc1b3e426803cb2, {16'd43392, 16'd61342, 16'd42198, 16'd36987, 16'd56813, 16'd57566, 16'd51194, 16'd16377, 16'd44664, 16'd26408, 16'd39605, 16'd43663, 16'd24362, 16'd59968, 16'd59697, 16'd7820, 16'd24901, 16'd8706, 16'd55668, 16'd59753, 16'd58906, 16'd40722, 16'd35294, 16'd14235, 16'd48116, 16'd5480});
	test_expansion(128'hf5490df7a0f4d01935bd74928b8a2835, {16'd13479, 16'd22808, 16'd8061, 16'd42705, 16'd56662, 16'd14256, 16'd3278, 16'd28772, 16'd64080, 16'd6212, 16'd50392, 16'd53505, 16'd52397, 16'd6885, 16'd20932, 16'd26151, 16'd26953, 16'd62671, 16'd26673, 16'd12064, 16'd43026, 16'd53867, 16'd22864, 16'd59838, 16'd18180, 16'd1112});
	test_expansion(128'he59b0614a48ebbc7ba9beb20b1e387bf, {16'd7383, 16'd58326, 16'd34675, 16'd1857, 16'd39690, 16'd54636, 16'd64062, 16'd53358, 16'd59244, 16'd56329, 16'd26433, 16'd35806, 16'd60048, 16'd36094, 16'd16928, 16'd6806, 16'd6494, 16'd36204, 16'd61673, 16'd34807, 16'd38898, 16'd29634, 16'd23848, 16'd15744, 16'd31543, 16'd31741});
	test_expansion(128'h98c5d62077880a7852d33d9892904a58, {16'd61915, 16'd42915, 16'd48913, 16'd57843, 16'd40620, 16'd49762, 16'd43710, 16'd58768, 16'd6233, 16'd32866, 16'd63253, 16'd8284, 16'd40463, 16'd59495, 16'd679, 16'd9538, 16'd60444, 16'd15113, 16'd54317, 16'd30220, 16'd6229, 16'd15050, 16'd22997, 16'd63702, 16'd59167, 16'd64076});
	test_expansion(128'h32c6bf72b018e543863b33f973f34efe, {16'd529, 16'd52843, 16'd11373, 16'd2511, 16'd52896, 16'd34759, 16'd27304, 16'd59848, 16'd21735, 16'd31947, 16'd30245, 16'd37511, 16'd55797, 16'd19327, 16'd36640, 16'd26345, 16'd54715, 16'd52450, 16'd57232, 16'd47321, 16'd59111, 16'd9042, 16'd13781, 16'd53200, 16'd45854, 16'd39853});
	test_expansion(128'h8900e7cd1aef9fd5538dde005c338bce, {16'd36045, 16'd17136, 16'd40600, 16'd21920, 16'd11376, 16'd35555, 16'd34529, 16'd40298, 16'd34551, 16'd8727, 16'd22594, 16'd31389, 16'd2029, 16'd34827, 16'd17167, 16'd14273, 16'd32512, 16'd40198, 16'd2819, 16'd17670, 16'd22527, 16'd4379, 16'd45329, 16'd23452, 16'd63464, 16'd58167});
	test_expansion(128'h131c555508cd586450e1d4df4da83d89, {16'd13591, 16'd55338, 16'd38131, 16'd32096, 16'd45309, 16'd23887, 16'd23984, 16'd56669, 16'd20925, 16'd9682, 16'd57484, 16'd60903, 16'd41279, 16'd17929, 16'd38546, 16'd12900, 16'd34219, 16'd28259, 16'd31666, 16'd28664, 16'd12058, 16'd64150, 16'd52979, 16'd51871, 16'd25222, 16'd50237});
	test_expansion(128'h9ba2bfec4fab2bb1737e1f0fc300087c, {16'd51283, 16'd9868, 16'd4801, 16'd28522, 16'd43796, 16'd17567, 16'd41017, 16'd38281, 16'd13780, 16'd49044, 16'd2574, 16'd35568, 16'd57320, 16'd31057, 16'd52161, 16'd26345, 16'd16278, 16'd40771, 16'd36766, 16'd39406, 16'd46726, 16'd13393, 16'd1325, 16'd37833, 16'd9578, 16'd1293});
	test_expansion(128'h10a80dc1e2c864ce5b6dc3d6e13889b2, {16'd65080, 16'd64764, 16'd44638, 16'd10593, 16'd37547, 16'd54689, 16'd59724, 16'd28615, 16'd55028, 16'd62855, 16'd12068, 16'd49747, 16'd39952, 16'd2611, 16'd15630, 16'd51761, 16'd50967, 16'd45617, 16'd10818, 16'd16101, 16'd41691, 16'd58686, 16'd40007, 16'd38332, 16'd40402, 16'd56301});
	test_expansion(128'hda2fbc3eb478c8ca334e6c14c499c4b5, {16'd49551, 16'd5450, 16'd50476, 16'd5180, 16'd28997, 16'd49530, 16'd15513, 16'd39828, 16'd30626, 16'd61205, 16'd57663, 16'd42751, 16'd9577, 16'd24534, 16'd65224, 16'd25673, 16'd49585, 16'd42946, 16'd45702, 16'd28185, 16'd355, 16'd2631, 16'd23413, 16'd28797, 16'd24056, 16'd6046});
	test_expansion(128'ha06a165c1a154772fd73f4fa90e713be, {16'd6159, 16'd14425, 16'd38434, 16'd8, 16'd61666, 16'd64346, 16'd15431, 16'd13977, 16'd16322, 16'd42752, 16'd46386, 16'd43905, 16'd31215, 16'd40554, 16'd40956, 16'd26846, 16'd38473, 16'd32485, 16'd6009, 16'd19997, 16'd50080, 16'd25846, 16'd31834, 16'd32667, 16'd33472, 16'd3161});
	test_expansion(128'h05441bc4fc0c29108e79038555026721, {16'd42684, 16'd52086, 16'd64365, 16'd34368, 16'd52867, 16'd3581, 16'd24660, 16'd53872, 16'd38077, 16'd13698, 16'd39874, 16'd16385, 16'd21235, 16'd41099, 16'd64902, 16'd24263, 16'd10506, 16'd47163, 16'd55104, 16'd31720, 16'd34696, 16'd19064, 16'd63313, 16'd9981, 16'd1667, 16'd17125});
	test_expansion(128'h67117feca4ab584f666dbb153db26daf, {16'd52318, 16'd17308, 16'd35119, 16'd21359, 16'd39257, 16'd35416, 16'd6176, 16'd6062, 16'd49427, 16'd5460, 16'd59683, 16'd5277, 16'd29939, 16'd37494, 16'd30057, 16'd62690, 16'd45027, 16'd24165, 16'd29459, 16'd10928, 16'd38368, 16'd64958, 16'd44412, 16'd1520, 16'd43508, 16'd64085});
	test_expansion(128'h35a0587347d2aeec626f7ad74bb589e2, {16'd52502, 16'd10919, 16'd13817, 16'd39597, 16'd22356, 16'd34771, 16'd35715, 16'd63024, 16'd29688, 16'd38682, 16'd29145, 16'd48460, 16'd1676, 16'd51515, 16'd64446, 16'd4756, 16'd10288, 16'd27120, 16'd10137, 16'd40821, 16'd28045, 16'd20274, 16'd15174, 16'd21211, 16'd32571, 16'd22942});
	test_expansion(128'h7c841f0ed8696dc961694a9dec1fd4e0, {16'd29383, 16'd58125, 16'd30569, 16'd2156, 16'd52825, 16'd18547, 16'd52428, 16'd50490, 16'd748, 16'd53877, 16'd54727, 16'd2203, 16'd45458, 16'd47912, 16'd40036, 16'd45575, 16'd18421, 16'd41327, 16'd61816, 16'd52909, 16'd46576, 16'd19233, 16'd369, 16'd3143, 16'd21019, 16'd39538});
	test_expansion(128'hf88e530fe1bba23b6a9a044fe84366f1, {16'd7393, 16'd49846, 16'd45598, 16'd26127, 16'd46547, 16'd25819, 16'd53188, 16'd12977, 16'd24669, 16'd19310, 16'd29349, 16'd57416, 16'd2804, 16'd15, 16'd40738, 16'd63789, 16'd43914, 16'd53180, 16'd7055, 16'd14097, 16'd28859, 16'd1300, 16'd16389, 16'd36072, 16'd58482, 16'd33321});
	test_expansion(128'hb46226897a57ff638e9ad3688d7cf192, {16'd10747, 16'd61175, 16'd25954, 16'd27974, 16'd38298, 16'd15727, 16'd2424, 16'd37887, 16'd58526, 16'd25680, 16'd38334, 16'd56407, 16'd23201, 16'd18584, 16'd22433, 16'd61855, 16'd23094, 16'd32170, 16'd44203, 16'd51273, 16'd44669, 16'd14998, 16'd30791, 16'd49413, 16'd61043, 16'd40283});
	test_expansion(128'h597dc7462de189719ae48b51cf6afbb9, {16'd52311, 16'd58827, 16'd3577, 16'd9427, 16'd51063, 16'd53376, 16'd42477, 16'd8548, 16'd2509, 16'd41737, 16'd45085, 16'd27788, 16'd5363, 16'd44279, 16'd25781, 16'd6677, 16'd41628, 16'd25071, 16'd18123, 16'd59420, 16'd22468, 16'd18113, 16'd10844, 16'd48376, 16'd50113, 16'd39867});
	test_expansion(128'h4393cb4e25f728be6de41db7202a19e2, {16'd11836, 16'd63064, 16'd18882, 16'd8233, 16'd63111, 16'd29586, 16'd5024, 16'd37370, 16'd14348, 16'd13088, 16'd25122, 16'd55835, 16'd3718, 16'd33315, 16'd20294, 16'd12344, 16'd33850, 16'd14288, 16'd14353, 16'd18055, 16'd17419, 16'd50965, 16'd23944, 16'd14109, 16'd54779, 16'd63477});
	test_expansion(128'h1cfdf93ac38cd81a343a9cb6add8ccb4, {16'd2081, 16'd3041, 16'd62354, 16'd51493, 16'd56794, 16'd60888, 16'd19462, 16'd19757, 16'd28176, 16'd62100, 16'd41827, 16'd32425, 16'd11639, 16'd43357, 16'd3038, 16'd421, 16'd62771, 16'd4320, 16'd17627, 16'd44287, 16'd54913, 16'd58611, 16'd1286, 16'd60838, 16'd55416, 16'd6472});
	test_expansion(128'h6271c8cd5d79ce73bfb6ec1d89538994, {16'd4027, 16'd60745, 16'd36038, 16'd12165, 16'd15647, 16'd65011, 16'd8940, 16'd53674, 16'd4757, 16'd8798, 16'd1056, 16'd42289, 16'd22775, 16'd36956, 16'd15370, 16'd8929, 16'd54292, 16'd29127, 16'd13798, 16'd5751, 16'd54948, 16'd33482, 16'd3, 16'd13036, 16'd39734, 16'd7837});
	test_expansion(128'hf87ee789a94c8fdc3879a9dc90feafd2, {16'd51117, 16'd15651, 16'd16026, 16'd34267, 16'd51114, 16'd49883, 16'd42212, 16'd17211, 16'd1123, 16'd48479, 16'd26107, 16'd57736, 16'd37272, 16'd21062, 16'd65310, 16'd29618, 16'd65137, 16'd14926, 16'd52048, 16'd3736, 16'd12475, 16'd55795, 16'd24613, 16'd52243, 16'd34232, 16'd36022});
	test_expansion(128'hd0b56a4c7b0d4053883c576038406cdf, {16'd5512, 16'd6055, 16'd18525, 16'd54966, 16'd3622, 16'd24480, 16'd24901, 16'd42869, 16'd11447, 16'd45529, 16'd49835, 16'd31189, 16'd44447, 16'd48065, 16'd14751, 16'd3379, 16'd52722, 16'd20323, 16'd24162, 16'd14462, 16'd48007, 16'd44901, 16'd3226, 16'd6925, 16'd60125, 16'd57212});
	test_expansion(128'hf50ccf6e9153064c84ab4ea83d189ff9, {16'd26670, 16'd30830, 16'd46925, 16'd43152, 16'd45291, 16'd26585, 16'd49913, 16'd54827, 16'd51203, 16'd27609, 16'd31213, 16'd42908, 16'd63979, 16'd50687, 16'd18907, 16'd27731, 16'd6705, 16'd36959, 16'd55, 16'd46688, 16'd33472, 16'd51544, 16'd21170, 16'd25236, 16'd64202, 16'd8384});
	test_expansion(128'h8fc346504997c59c6d58b6d6d8c499e0, {16'd7486, 16'd259, 16'd49123, 16'd33706, 16'd35075, 16'd53597, 16'd4285, 16'd13332, 16'd63920, 16'd16176, 16'd10621, 16'd62500, 16'd18752, 16'd61257, 16'd34635, 16'd62342, 16'd48553, 16'd21285, 16'd2329, 16'd33119, 16'd25840, 16'd54725, 16'd55088, 16'd8984, 16'd294, 16'd48731});
	test_expansion(128'h4e6ecacc2fb1c21dd56a47a390bd4b4d, {16'd14235, 16'd11538, 16'd1079, 16'd30058, 16'd14261, 16'd6754, 16'd54672, 16'd63011, 16'd31428, 16'd20371, 16'd63516, 16'd41005, 16'd42728, 16'd26754, 16'd30493, 16'd8271, 16'd29960, 16'd57650, 16'd18094, 16'd55985, 16'd51330, 16'd36672, 16'd62, 16'd15244, 16'd55968, 16'd51783});
	test_expansion(128'ha9e93f9f9aec4a3a40c4e0e15b693052, {16'd57117, 16'd23091, 16'd44035, 16'd57126, 16'd20889, 16'd18288, 16'd3031, 16'd42039, 16'd20830, 16'd42931, 16'd37094, 16'd58467, 16'd17142, 16'd60966, 16'd28888, 16'd17397, 16'd12933, 16'd32196, 16'd57094, 16'd29997, 16'd63011, 16'd38862, 16'd54885, 16'd35532, 16'd1951, 16'd60801});
	test_expansion(128'h22616078f277cab3443778707e112e60, {16'd21604, 16'd18401, 16'd33127, 16'd10072, 16'd44679, 16'd57799, 16'd18510, 16'd35887, 16'd6120, 16'd10331, 16'd1706, 16'd8084, 16'd30712, 16'd31917, 16'd12878, 16'd8429, 16'd38395, 16'd8308, 16'd17772, 16'd57238, 16'd13986, 16'd34214, 16'd56508, 16'd19954, 16'd8111, 16'd8017});
	test_expansion(128'h4b474d0db9ff6db52ece405356460b82, {16'd25520, 16'd8315, 16'd2035, 16'd50018, 16'd3871, 16'd33742, 16'd57947, 16'd20151, 16'd37126, 16'd35585, 16'd1586, 16'd536, 16'd13897, 16'd24606, 16'd6077, 16'd17479, 16'd30220, 16'd4038, 16'd43563, 16'd19749, 16'd49450, 16'd57496, 16'd16866, 16'd15773, 16'd28849, 16'd10645});
	test_expansion(128'hd7da18f9b180c34f97b4be3d28f3f863, {16'd16837, 16'd58334, 16'd45747, 16'd36972, 16'd21128, 16'd2780, 16'd34121, 16'd35200, 16'd8062, 16'd10888, 16'd50575, 16'd25621, 16'd40511, 16'd40827, 16'd56195, 16'd600, 16'd49067, 16'd23419, 16'd48019, 16'd34073, 16'd35071, 16'd16961, 16'd56049, 16'd23587, 16'd28561, 16'd3155});
	test_expansion(128'h85d6cb4ac2ce5c86dbf8be3145c6110f, {16'd40029, 16'd44730, 16'd14169, 16'd646, 16'd17950, 16'd57145, 16'd7664, 16'd62290, 16'd30141, 16'd7879, 16'd258, 16'd64668, 16'd63571, 16'd52380, 16'd6356, 16'd36447, 16'd15218, 16'd56672, 16'd11151, 16'd62282, 16'd53710, 16'd42199, 16'd35105, 16'd60528, 16'd58758, 16'd1471});
	test_expansion(128'h806c53ab137a790b0cdff94235ff4f15, {16'd14053, 16'd52770, 16'd31012, 16'd64563, 16'd23569, 16'd45407, 16'd53768, 16'd33670, 16'd7083, 16'd18853, 16'd45855, 16'd18181, 16'd36574, 16'd54790, 16'd23962, 16'd24917, 16'd39907, 16'd55365, 16'd29065, 16'd47768, 16'd21017, 16'd5776, 16'd64869, 16'd55860, 16'd29702, 16'd51432});
	test_expansion(128'h6f685f5661d161c4b0e6a76492555053, {16'd46260, 16'd3744, 16'd34730, 16'd20068, 16'd26919, 16'd42991, 16'd6999, 16'd62367, 16'd22618, 16'd3596, 16'd7279, 16'd53611, 16'd58638, 16'd19998, 16'd11433, 16'd40283, 16'd22837, 16'd16558, 16'd15580, 16'd56116, 16'd44299, 16'd4362, 16'd26146, 16'd45974, 16'd831, 16'd49987});
	test_expansion(128'h738ff437b763a3f18417b75567dd88da, {16'd22789, 16'd5430, 16'd43050, 16'd44675, 16'd535, 16'd36989, 16'd45651, 16'd38960, 16'd63152, 16'd30938, 16'd11794, 16'd9690, 16'd61395, 16'd22657, 16'd61469, 16'd46799, 16'd16686, 16'd43629, 16'd47222, 16'd18752, 16'd1078, 16'd37455, 16'd51709, 16'd24495, 16'd33367, 16'd3109});
	test_expansion(128'h7b4380d2a38349a22b6e6e77ad7aead6, {16'd58909, 16'd49467, 16'd46221, 16'd52766, 16'd11441, 16'd29643, 16'd5953, 16'd49473, 16'd32132, 16'd18272, 16'd6104, 16'd49565, 16'd60468, 16'd868, 16'd41867, 16'd51994, 16'd52791, 16'd62849, 16'd39899, 16'd14055, 16'd15155, 16'd60153, 16'd25087, 16'd6529, 16'd58816, 16'd40158});
	test_expansion(128'h77f1f34fac876f87eac526da29c207de, {16'd23519, 16'd12754, 16'd47177, 16'd36964, 16'd39255, 16'd57304, 16'd23958, 16'd60556, 16'd46564, 16'd64473, 16'd41446, 16'd37427, 16'd55365, 16'd17764, 16'd44555, 16'd26199, 16'd61076, 16'd52500, 16'd6267, 16'd62415, 16'd45463, 16'd32941, 16'd34621, 16'd40271, 16'd49560, 16'd13253});
	test_expansion(128'hcf9502dee324c42658a8cfc32bf7fa38, {16'd10927, 16'd57023, 16'd52096, 16'd12161, 16'd25507, 16'd29958, 16'd56091, 16'd59737, 16'd15831, 16'd26345, 16'd37459, 16'd16726, 16'd10128, 16'd17788, 16'd46012, 16'd14154, 16'd9159, 16'd60637, 16'd11269, 16'd11616, 16'd32430, 16'd37320, 16'd42454, 16'd13972, 16'd57917, 16'd7441});
	test_expansion(128'h72bbb25ffcb34a13c2a6cb8f9245f37c, {16'd52793, 16'd33249, 16'd21526, 16'd9948, 16'd24698, 16'd48239, 16'd48699, 16'd33340, 16'd58592, 16'd44007, 16'd49838, 16'd52748, 16'd9083, 16'd5387, 16'd11824, 16'd33600, 16'd53891, 16'd27551, 16'd63977, 16'd20226, 16'd30289, 16'd44266, 16'd7456, 16'd60722, 16'd51254, 16'd3866});
	test_expansion(128'h5d33f8dae95c3c0792d06936a6dd4227, {16'd6838, 16'd37778, 16'd19227, 16'd38007, 16'd36836, 16'd56928, 16'd6528, 16'd56047, 16'd878, 16'd64754, 16'd3437, 16'd41763, 16'd9399, 16'd24591, 16'd58586, 16'd20332, 16'd4288, 16'd65495, 16'd65018, 16'd33973, 16'd29725, 16'd64047, 16'd22638, 16'd37399, 16'd33522, 16'd53019});
	test_expansion(128'hbb0858aa9a845e554eb89da3a20e19a0, {16'd30604, 16'd23545, 16'd15684, 16'd2259, 16'd64710, 16'd8892, 16'd32532, 16'd27919, 16'd63100, 16'd35966, 16'd18586, 16'd30982, 16'd48937, 16'd62837, 16'd27083, 16'd56198, 16'd46317, 16'd8132, 16'd25257, 16'd37154, 16'd6655, 16'd15078, 16'd9111, 16'd10187, 16'd56671, 16'd33705});
	test_expansion(128'h928b9516a1a7e635802cd633ecf2f795, {16'd15901, 16'd46342, 16'd30926, 16'd54165, 16'd26995, 16'd38646, 16'd52986, 16'd61514, 16'd4330, 16'd40130, 16'd40466, 16'd33167, 16'd17041, 16'd3070, 16'd52353, 16'd6697, 16'd46933, 16'd22284, 16'd58686, 16'd17672, 16'd33491, 16'd23166, 16'd6252, 16'd28731, 16'd28859, 16'd52428});
	test_expansion(128'h745931155273e33ef13064c87b2a4aa4, {16'd34907, 16'd63976, 16'd9570, 16'd27337, 16'd38755, 16'd64380, 16'd16500, 16'd29515, 16'd25396, 16'd58169, 16'd39144, 16'd18241, 16'd62110, 16'd29067, 16'd64012, 16'd20654, 16'd37803, 16'd2943, 16'd33972, 16'd43541, 16'd2359, 16'd19070, 16'd46883, 16'd18727, 16'd37492, 16'd16955});
	test_expansion(128'h4501099af0826379475a02adb9bfba21, {16'd22611, 16'd24351, 16'd21995, 16'd23946, 16'd29892, 16'd33339, 16'd28473, 16'd4457, 16'd5053, 16'd44903, 16'd62574, 16'd33050, 16'd9911, 16'd58297, 16'd61451, 16'd12973, 16'd12741, 16'd60592, 16'd47219, 16'd27888, 16'd52984, 16'd20341, 16'd45071, 16'd63041, 16'd21989, 16'd39142});
	test_expansion(128'h3eff18c98b8a681797767b0334f1bf8b, {16'd9565, 16'd11883, 16'd18675, 16'd7901, 16'd50502, 16'd44982, 16'd29508, 16'd26265, 16'd10355, 16'd53861, 16'd9864, 16'd63808, 16'd6196, 16'd57079, 16'd19607, 16'd27340, 16'd45775, 16'd48202, 16'd28882, 16'd9675, 16'd21062, 16'd51501, 16'd54861, 16'd4735, 16'd26701, 16'd19882});
	test_expansion(128'h47e93928c199acc272b133875b8d0184, {16'd23907, 16'd46706, 16'd40669, 16'd40210, 16'd60232, 16'd43665, 16'd12232, 16'd56955, 16'd46878, 16'd11688, 16'd43715, 16'd41014, 16'd61583, 16'd58623, 16'd20874, 16'd53688, 16'd6920, 16'd36964, 16'd4468, 16'd29542, 16'd42989, 16'd22211, 16'd14761, 16'd5709, 16'd8182, 16'd1938});
	test_expansion(128'hbb6ba26cb2bdb9e8ed0da4697db92fa1, {16'd8652, 16'd6389, 16'd40818, 16'd21124, 16'd52950, 16'd62477, 16'd11939, 16'd41233, 16'd25674, 16'd29998, 16'd54030, 16'd63015, 16'd42625, 16'd48910, 16'd35377, 16'd7391, 16'd31834, 16'd52423, 16'd39248, 16'd27083, 16'd48579, 16'd30322, 16'd44416, 16'd24685, 16'd38362, 16'd45705});
	test_expansion(128'h6d5744a07cc9b26908abace2eaad104f, {16'd34178, 16'd21400, 16'd52585, 16'd6817, 16'd22077, 16'd57377, 16'd29641, 16'd17531, 16'd62776, 16'd17255, 16'd36497, 16'd8501, 16'd4788, 16'd15548, 16'd1943, 16'd4597, 16'd8436, 16'd46547, 16'd42791, 16'd58114, 16'd31884, 16'd26948, 16'd56278, 16'd11954, 16'd23534, 16'd5833});
	test_expansion(128'h6c1b736efffcb9aff6b313d5bf48ed09, {16'd64649, 16'd23348, 16'd35094, 16'd44097, 16'd38213, 16'd48946, 16'd4376, 16'd5875, 16'd33717, 16'd4414, 16'd18811, 16'd64182, 16'd52477, 16'd30925, 16'd51732, 16'd28018, 16'd54342, 16'd23130, 16'd33319, 16'd34970, 16'd60793, 16'd54140, 16'd64051, 16'd32504, 16'd53071, 16'd57382});
	test_expansion(128'h3b4615bc7904c1210475f321442262c7, {16'd15389, 16'd26269, 16'd3293, 16'd5632, 16'd4346, 16'd20809, 16'd48698, 16'd32471, 16'd25472, 16'd63599, 16'd13909, 16'd20599, 16'd19282, 16'd47487, 16'd28008, 16'd43697, 16'd53525, 16'd48889, 16'd31659, 16'd18105, 16'd42285, 16'd37634, 16'd48898, 16'd22789, 16'd63505, 16'd34141});
	test_expansion(128'h214fe883574b0569c749ff373a08a11f, {16'd16970, 16'd35213, 16'd48437, 16'd6728, 16'd48665, 16'd37973, 16'd42040, 16'd58561, 16'd2649, 16'd26182, 16'd11450, 16'd49576, 16'd58308, 16'd55955, 16'd8219, 16'd57749, 16'd11888, 16'd11051, 16'd60837, 16'd3124, 16'd9716, 16'd15150, 16'd11155, 16'd38230, 16'd35762, 16'd36766});
	test_expansion(128'h53c3d9a77f6d17ee9d8003c2771df22e, {16'd8251, 16'd43521, 16'd61653, 16'd10436, 16'd47431, 16'd48428, 16'd55218, 16'd59527, 16'd38024, 16'd45813, 16'd33323, 16'd46848, 16'd57567, 16'd25981, 16'd1775, 16'd23109, 16'd53715, 16'd31373, 16'd16864, 16'd12054, 16'd44237, 16'd3835, 16'd23094, 16'd7876, 16'd23824, 16'd20070});
	test_expansion(128'hbca6f2bb28a52f1c635208c372ed49aa, {16'd29490, 16'd15703, 16'd44111, 16'd49610, 16'd40859, 16'd33846, 16'd42820, 16'd23630, 16'd3352, 16'd7205, 16'd64768, 16'd9842, 16'd18455, 16'd35729, 16'd32121, 16'd63029, 16'd37211, 16'd31127, 16'd6913, 16'd23672, 16'd8653, 16'd16206, 16'd33095, 16'd11127, 16'd47592, 16'd32239});
	test_expansion(128'hbe6788f1e957111f0a42877a051de12b, {16'd24415, 16'd25392, 16'd58803, 16'd16521, 16'd46123, 16'd60033, 16'd13897, 16'd411, 16'd34121, 16'd65198, 16'd59410, 16'd4987, 16'd35631, 16'd63153, 16'd49502, 16'd14523, 16'd30328, 16'd58178, 16'd40695, 16'd37704, 16'd58828, 16'd33888, 16'd8245, 16'd7031, 16'd2645, 16'd56539});
	test_expansion(128'h81b68bd42ba23d894eae361fdbf55fa9, {16'd5978, 16'd44637, 16'd25048, 16'd35906, 16'd49575, 16'd16122, 16'd37745, 16'd58671, 16'd1779, 16'd42843, 16'd501, 16'd42281, 16'd62357, 16'd24691, 16'd35269, 16'd61874, 16'd55660, 16'd18679, 16'd36606, 16'd3194, 16'd7537, 16'd30396, 16'd5256, 16'd22722, 16'd53714, 16'd2298});
	test_expansion(128'h2c43dbfc01606ef67c9879b4bd4d067d, {16'd64902, 16'd22021, 16'd5046, 16'd36787, 16'd42722, 16'd58943, 16'd39285, 16'd25038, 16'd23170, 16'd1349, 16'd44252, 16'd39743, 16'd9917, 16'd47790, 16'd26245, 16'd5639, 16'd17362, 16'd17492, 16'd52457, 16'd64415, 16'd14738, 16'd32834, 16'd33201, 16'd30536, 16'd12635, 16'd25372});
	test_expansion(128'h0f24ea37d5095eee4a42621567618228, {16'd55321, 16'd64807, 16'd9620, 16'd53736, 16'd11793, 16'd56706, 16'd52092, 16'd25197, 16'd34581, 16'd16593, 16'd53721, 16'd16524, 16'd31094, 16'd15048, 16'd21478, 16'd41784, 16'd44547, 16'd8737, 16'd14932, 16'd55664, 16'd25051, 16'd16225, 16'd24383, 16'd55252, 16'd49304, 16'd65324});
	test_expansion(128'h85bebfe54805a070662e241d8c957ca4, {16'd19858, 16'd50097, 16'd63732, 16'd18892, 16'd39588, 16'd62257, 16'd59565, 16'd6613, 16'd35947, 16'd52095, 16'd32860, 16'd63899, 16'd59653, 16'd29385, 16'd48838, 16'd35623, 16'd63485, 16'd46745, 16'd53194, 16'd47044, 16'd56552, 16'd25199, 16'd42277, 16'd26429, 16'd31404, 16'd58301});
	test_expansion(128'h875998ac8c79d7fdc661970dc0a391ec, {16'd10240, 16'd48823, 16'd39965, 16'd54198, 16'd11721, 16'd41401, 16'd40818, 16'd45072, 16'd12988, 16'd22342, 16'd28086, 16'd27119, 16'd47875, 16'd18151, 16'd29063, 16'd36880, 16'd64453, 16'd29706, 16'd64068, 16'd9997, 16'd37309, 16'd16672, 16'd17130, 16'd12666, 16'd55178, 16'd13576});
	test_expansion(128'hadaeb3a5a463ab3a3ef55955ca424d62, {16'd36724, 16'd37769, 16'd39863, 16'd16110, 16'd3224, 16'd37848, 16'd17623, 16'd25310, 16'd62659, 16'd1729, 16'd54376, 16'd29616, 16'd46064, 16'd23921, 16'd57679, 16'd58458, 16'd2670, 16'd34880, 16'd49871, 16'd57970, 16'd52313, 16'd650, 16'd64906, 16'd1198, 16'd53051, 16'd9023});
	test_expansion(128'h67b74f387a07f1a7aa5009952ed3f2d0, {16'd54429, 16'd31289, 16'd43590, 16'd15338, 16'd44010, 16'd24304, 16'd16013, 16'd45775, 16'd18255, 16'd22905, 16'd1932, 16'd39900, 16'd51521, 16'd49080, 16'd36646, 16'd38101, 16'd25515, 16'd5623, 16'd5133, 16'd40069, 16'd20838, 16'd42353, 16'd28678, 16'd52573, 16'd55098, 16'd11004});
	test_expansion(128'h5b147493b237c8c6b8503c565f5914dd, {16'd40287, 16'd22492, 16'd44242, 16'd12870, 16'd14047, 16'd46751, 16'd6330, 16'd10013, 16'd42715, 16'd26097, 16'd63424, 16'd39968, 16'd43420, 16'd35377, 16'd15396, 16'd16218, 16'd57897, 16'd59287, 16'd8197, 16'd46392, 16'd16853, 16'd7316, 16'd8319, 16'd19967, 16'd12434, 16'd17723});
	test_expansion(128'h939a18942874f43f6b74388f604f7bfb, {16'd45310, 16'd40313, 16'd20851, 16'd63609, 16'd9687, 16'd52835, 16'd42584, 16'd31473, 16'd53979, 16'd3135, 16'd51097, 16'd34837, 16'd3850, 16'd63560, 16'd58388, 16'd5426, 16'd27179, 16'd44840, 16'd7843, 16'd57094, 16'd30592, 16'd62965, 16'd18186, 16'd34253, 16'd3044, 16'd40174});
	test_expansion(128'hd84631296ad145aede2e7c9f6a086c05, {16'd58835, 16'd25403, 16'd55654, 16'd30440, 16'd44120, 16'd59258, 16'd29478, 16'd34182, 16'd13084, 16'd22813, 16'd49225, 16'd22531, 16'd65455, 16'd21701, 16'd24197, 16'd22584, 16'd31896, 16'd39958, 16'd46416, 16'd52839, 16'd14059, 16'd14514, 16'd60599, 16'd34374, 16'd58796, 16'd53629});
	test_expansion(128'hf3210e1feb4d604e84c94d4788c3fa2b, {16'd24609, 16'd58507, 16'd16661, 16'd12628, 16'd30027, 16'd26882, 16'd59112, 16'd14457, 16'd6594, 16'd35668, 16'd61775, 16'd9363, 16'd34204, 16'd11632, 16'd14872, 16'd40001, 16'd24778, 16'd36872, 16'd20131, 16'd59319, 16'd2009, 16'd10874, 16'd59114, 16'd17596, 16'd53684, 16'd4537});
	test_expansion(128'h21f2222de38b8b0af6e8c9a8909e3e45, {16'd45620, 16'd27022, 16'd62020, 16'd37672, 16'd4948, 16'd17193, 16'd49975, 16'd26565, 16'd64343, 16'd53277, 16'd40202, 16'd30865, 16'd48928, 16'd64389, 16'd6996, 16'd54119, 16'd3117, 16'd48982, 16'd32887, 16'd25495, 16'd12601, 16'd43403, 16'd81, 16'd28731, 16'd3654, 16'd48531});
	test_expansion(128'h0e3daf60f811d060ca91ae9a38aafee7, {16'd16247, 16'd58399, 16'd52982, 16'd18335, 16'd795, 16'd11296, 16'd48535, 16'd2582, 16'd11076, 16'd59487, 16'd7046, 16'd7518, 16'd56108, 16'd17430, 16'd20145, 16'd29333, 16'd60869, 16'd26619, 16'd9892, 16'd20245, 16'd6308, 16'd60962, 16'd10062, 16'd65160, 16'd19592, 16'd22930});
	test_expansion(128'hd72c4da7acc9d2c29bc1b7025a51c7fe, {16'd4470, 16'd36966, 16'd39456, 16'd18188, 16'd45628, 16'd44789, 16'd38028, 16'd34728, 16'd31560, 16'd62524, 16'd30741, 16'd41644, 16'd26118, 16'd58089, 16'd44921, 16'd8736, 16'd55771, 16'd41161, 16'd22226, 16'd17523, 16'd51235, 16'd27137, 16'd8025, 16'd39628, 16'd13044, 16'd41932});
	test_expansion(128'h7e86f1f12f2ecac7f896f64ffad5984a, {16'd19111, 16'd12397, 16'd49120, 16'd41363, 16'd1005, 16'd22599, 16'd42701, 16'd44160, 16'd57663, 16'd12449, 16'd10631, 16'd34961, 16'd65405, 16'd6488, 16'd55115, 16'd19761, 16'd27542, 16'd22086, 16'd15168, 16'd48087, 16'd31553, 16'd5182, 16'd52237, 16'd12025, 16'd27464, 16'd47290});
	test_expansion(128'hdde3204a135ee126b6cbf043c6fde49c, {16'd21478, 16'd23790, 16'd9794, 16'd7220, 16'd16895, 16'd50704, 16'd54130, 16'd34190, 16'd9977, 16'd26141, 16'd43502, 16'd33038, 16'd56471, 16'd22298, 16'd33746, 16'd36131, 16'd17443, 16'd63794, 16'd20182, 16'd13045, 16'd353, 16'd4771, 16'd44752, 16'd46120, 16'd18151, 16'd58172});
	test_expansion(128'h8423f762395b492701e5615131139e2b, {16'd61497, 16'd56735, 16'd35456, 16'd37555, 16'd55313, 16'd37620, 16'd16467, 16'd837, 16'd52421, 16'd3354, 16'd37282, 16'd1808, 16'd21376, 16'd39850, 16'd9757, 16'd36340, 16'd25193, 16'd53979, 16'd54717, 16'd15028, 16'd53222, 16'd26835, 16'd25332, 16'd32053, 16'd16729, 16'd52104});
	test_expansion(128'h9c40656435f2daa8e6902ca2fc29062b, {16'd2580, 16'd43510, 16'd61666, 16'd43185, 16'd44598, 16'd52715, 16'd4103, 16'd6580, 16'd30308, 16'd62988, 16'd705, 16'd39865, 16'd50220, 16'd42513, 16'd48558, 16'd20567, 16'd12249, 16'd50516, 16'd24731, 16'd19587, 16'd49437, 16'd31102, 16'd15869, 16'd9816, 16'd63532, 16'd6086});
	test_expansion(128'hbe8463ea5048cb22890980d4ae694f28, {16'd30508, 16'd5431, 16'd45005, 16'd19538, 16'd7946, 16'd4359, 16'd10923, 16'd27360, 16'd16284, 16'd33267, 16'd41894, 16'd55984, 16'd29101, 16'd42526, 16'd1847, 16'd24818, 16'd40106, 16'd13424, 16'd5542, 16'd51606, 16'd39174, 16'd25474, 16'd9744, 16'd28980, 16'd17169, 16'd47753});
	test_expansion(128'h55799280d2dbaf938dad3df4f98e338a, {16'd7510, 16'd57685, 16'd23685, 16'd4703, 16'd22123, 16'd42843, 16'd53850, 16'd2890, 16'd51444, 16'd13461, 16'd21900, 16'd31858, 16'd46968, 16'd61496, 16'd31333, 16'd55581, 16'd16105, 16'd38171, 16'd11092, 16'd40650, 16'd44892, 16'd11705, 16'd62280, 16'd51207, 16'd12892, 16'd14752});
	test_expansion(128'h3a992a6313ce21b6412ca8992c29e3a8, {16'd32882, 16'd41230, 16'd7451, 16'd47263, 16'd40913, 16'd37111, 16'd25316, 16'd10724, 16'd44504, 16'd26876, 16'd34835, 16'd48537, 16'd40060, 16'd46184, 16'd51597, 16'd28453, 16'd50896, 16'd16879, 16'd24100, 16'd42891, 16'd31541, 16'd111, 16'd17265, 16'd24817, 16'd41989, 16'd47177});
	test_expansion(128'hd63a60eb95bee214f01707ec77c5cad2, {16'd40458, 16'd55375, 16'd12760, 16'd59648, 16'd20859, 16'd53360, 16'd54053, 16'd14756, 16'd65189, 16'd28446, 16'd32067, 16'd48097, 16'd17322, 16'd34028, 16'd8785, 16'd28361, 16'd52217, 16'd19764, 16'd4150, 16'd9691, 16'd12888, 16'd7531, 16'd33769, 16'd31252, 16'd24063, 16'd24795});
	test_expansion(128'h498569ad6ccf90b7f923a6edcf9e00ab, {16'd55381, 16'd50769, 16'd31740, 16'd22778, 16'd26991, 16'd29092, 16'd12483, 16'd25403, 16'd46185, 16'd48024, 16'd634, 16'd54156, 16'd63439, 16'd4662, 16'd62188, 16'd57134, 16'd29185, 16'd48129, 16'd35100, 16'd64059, 16'd41120, 16'd61013, 16'd14340, 16'd39552, 16'd51930, 16'd17327});
	test_expansion(128'h48f4418bfda1256513149afb76213a29, {16'd53488, 16'd37791, 16'd33359, 16'd27378, 16'd43881, 16'd57836, 16'd25451, 16'd61575, 16'd56585, 16'd19365, 16'd63784, 16'd8188, 16'd949, 16'd51346, 16'd39723, 16'd48735, 16'd51473, 16'd58071, 16'd34908, 16'd27400, 16'd22562, 16'd25415, 16'd43878, 16'd50555, 16'd46681, 16'd63198});
	test_expansion(128'h15b0dbc3a361c5b40d1c6c5477b3a103, {16'd16338, 16'd47810, 16'd52351, 16'd20243, 16'd48360, 16'd11390, 16'd35683, 16'd24942, 16'd28156, 16'd29611, 16'd59349, 16'd3499, 16'd20634, 16'd62731, 16'd17941, 16'd4693, 16'd12499, 16'd58119, 16'd3352, 16'd4978, 16'd51860, 16'd58352, 16'd31096, 16'd14246, 16'd3401, 16'd53946});
	test_expansion(128'h0ae3d21af86cc163df9dfd16d2170d89, {16'd49366, 16'd18890, 16'd38559, 16'd21269, 16'd29698, 16'd14144, 16'd64705, 16'd5953, 16'd55117, 16'd7985, 16'd3181, 16'd27972, 16'd65273, 16'd50556, 16'd52314, 16'd30455, 16'd40340, 16'd28906, 16'd50961, 16'd22062, 16'd43669, 16'd45159, 16'd15500, 16'd36199, 16'd53255, 16'd65024});
	test_expansion(128'hab30715e1f7fb55ab479253d2af907e2, {16'd62110, 16'd55791, 16'd33486, 16'd2065, 16'd23862, 16'd19074, 16'd40641, 16'd39157, 16'd30757, 16'd25150, 16'd13015, 16'd53389, 16'd57062, 16'd17492, 16'd63141, 16'd42834, 16'd53207, 16'd43398, 16'd63896, 16'd28164, 16'd54260, 16'd46544, 16'd15200, 16'd3889, 16'd42447, 16'd14914});
	test_expansion(128'h9573769b873485fda9b24ccdf54babdd, {16'd32427, 16'd17326, 16'd10598, 16'd21476, 16'd22163, 16'd21099, 16'd27378, 16'd48096, 16'd57703, 16'd43525, 16'd53559, 16'd17292, 16'd8591, 16'd51502, 16'd26404, 16'd52139, 16'd33401, 16'd46345, 16'd55449, 16'd62605, 16'd62516, 16'd38323, 16'd43530, 16'd37208, 16'd23666, 16'd35516});
	test_expansion(128'h9b8538df49af3d2d825d017a6286664f, {16'd49562, 16'd254, 16'd58756, 16'd59161, 16'd49324, 16'd12645, 16'd25770, 16'd48189, 16'd34490, 16'd54764, 16'd65455, 16'd61162, 16'd24318, 16'd61453, 16'd19092, 16'd63429, 16'd41589, 16'd22783, 16'd39051, 16'd7422, 16'd14676, 16'd34667, 16'd28571, 16'd643, 16'd54886, 16'd40150});
	test_expansion(128'h039e05a8c7204cee747eab026a46a10e, {16'd1181, 16'd2321, 16'd20271, 16'd8206, 16'd39778, 16'd50508, 16'd16434, 16'd34067, 16'd9030, 16'd31545, 16'd30292, 16'd57386, 16'd40925, 16'd13075, 16'd36663, 16'd40567, 16'd38395, 16'd21477, 16'd43699, 16'd59139, 16'd18256, 16'd52274, 16'd2446, 16'd8226, 16'd30070, 16'd60944});
	test_expansion(128'h8cdcd4fe4e52c7218c9366cdf4540d92, {16'd24003, 16'd50257, 16'd4392, 16'd58593, 16'd35504, 16'd29825, 16'd48639, 16'd56193, 16'd36565, 16'd34395, 16'd14886, 16'd8703, 16'd24986, 16'd26649, 16'd11056, 16'd819, 16'd31413, 16'd19275, 16'd57307, 16'd12104, 16'd37270, 16'd26510, 16'd19076, 16'd59837, 16'd30561, 16'd5304});
	test_expansion(128'hcf09677fcd6fbb4b69550361dad31928, {16'd3581, 16'd49471, 16'd49984, 16'd25928, 16'd46844, 16'd56579, 16'd7347, 16'd53455, 16'd6170, 16'd43110, 16'd58880, 16'd27274, 16'd46135, 16'd38780, 16'd59003, 16'd6325, 16'd48395, 16'd10381, 16'd22031, 16'd18958, 16'd4055, 16'd23129, 16'd20852, 16'd30220, 16'd62268, 16'd16844});
	test_expansion(128'h3ac043ed778eca3e14ad3de8d6df8988, {16'd48185, 16'd19887, 16'd12553, 16'd14287, 16'd17336, 16'd11987, 16'd22403, 16'd44268, 16'd1874, 16'd38993, 16'd36344, 16'd58720, 16'd43196, 16'd14846, 16'd13915, 16'd21580, 16'd43078, 16'd44430, 16'd41908, 16'd26644, 16'd56544, 16'd17968, 16'd62407, 16'd29851, 16'd10182, 16'd35459});
	test_expansion(128'h002b659f7f349af935c2c34815883298, {16'd36711, 16'd61045, 16'd13916, 16'd28636, 16'd63537, 16'd27225, 16'd24962, 16'd5059, 16'd38915, 16'd30974, 16'd52269, 16'd61608, 16'd25247, 16'd17900, 16'd65436, 16'd59460, 16'd10222, 16'd59499, 16'd4631, 16'd52854, 16'd29166, 16'd25397, 16'd56543, 16'd18649, 16'd206, 16'd4769});
	test_expansion(128'hbd6c65b5ca7ea8d5e81a26640747b368, {16'd21073, 16'd7652, 16'd1681, 16'd65106, 16'd26643, 16'd45947, 16'd13033, 16'd17072, 16'd3202, 16'd47818, 16'd55110, 16'd48951, 16'd6779, 16'd63361, 16'd2936, 16'd54932, 16'd28143, 16'd50361, 16'd19662, 16'd10696, 16'd2286, 16'd378, 16'd1633, 16'd13299, 16'd21313, 16'd988});
	test_expansion(128'h3574a255dc317c6a5a2e12f034bae93b, {16'd49537, 16'd54868, 16'd15756, 16'd60681, 16'd877, 16'd28672, 16'd45627, 16'd30164, 16'd26515, 16'd30329, 16'd29311, 16'd7547, 16'd24165, 16'd18856, 16'd27060, 16'd52320, 16'd55646, 16'd30424, 16'd1357, 16'd62697, 16'd7825, 16'd11153, 16'd11002, 16'd59205, 16'd53832, 16'd1059});
	test_expansion(128'h3bdb43e57893cc85812717330fd8417f, {16'd19786, 16'd16317, 16'd19885, 16'd27744, 16'd26425, 16'd45021, 16'd26060, 16'd33243, 16'd54864, 16'd50151, 16'd1227, 16'd28363, 16'd5420, 16'd36380, 16'd962, 16'd39443, 16'd38697, 16'd52271, 16'd61421, 16'd44221, 16'd15512, 16'd32286, 16'd9824, 16'd17366, 16'd31822, 16'd42201});
	test_expansion(128'h3d82397f83db5d37173faace34de96c8, {16'd14681, 16'd5344, 16'd19880, 16'd46419, 16'd11407, 16'd283, 16'd51949, 16'd53282, 16'd20411, 16'd5050, 16'd2504, 16'd4704, 16'd20993, 16'd44709, 16'd18133, 16'd25392, 16'd34235, 16'd49364, 16'd53599, 16'd58281, 16'd47103, 16'd8841, 16'd32023, 16'd31233, 16'd30672, 16'd8321});
	test_expansion(128'he6c34fabc2b1ee09f4010d3320b73ad2, {16'd39998, 16'd12793, 16'd55739, 16'd49432, 16'd27324, 16'd1350, 16'd24228, 16'd61884, 16'd27579, 16'd21157, 16'd58133, 16'd38284, 16'd2479, 16'd31489, 16'd6154, 16'd59227, 16'd11167, 16'd28727, 16'd56584, 16'd46957, 16'd21437, 16'd1686, 16'd61319, 16'd55815, 16'd52820, 16'd50349});
	test_expansion(128'h97fb4f7932ed506355fb2c42877f5a39, {16'd58488, 16'd53057, 16'd14628, 16'd17662, 16'd52115, 16'd57461, 16'd11058, 16'd19420, 16'd18802, 16'd52553, 16'd35207, 16'd51871, 16'd25840, 16'd13584, 16'd39086, 16'd47642, 16'd48079, 16'd53773, 16'd18919, 16'd24513, 16'd51787, 16'd8162, 16'd15640, 16'd36017, 16'd64247, 16'd22674});
	test_expansion(128'h0c46eef34e2a8703839c65884b3c3654, {16'd12641, 16'd35505, 16'd187, 16'd54587, 16'd28955, 16'd47949, 16'd37618, 16'd16246, 16'd18320, 16'd31143, 16'd56262, 16'd15239, 16'd60160, 16'd58869, 16'd42495, 16'd33949, 16'd28818, 16'd56694, 16'd50303, 16'd8012, 16'd56325, 16'd11767, 16'd11159, 16'd45232, 16'd26498, 16'd32038});
	test_expansion(128'h21b1b61550e13b616c0d7e10e4d9bb4e, {16'd36014, 16'd48644, 16'd40825, 16'd43891, 16'd11223, 16'd58838, 16'd28874, 16'd61846, 16'd47091, 16'd56072, 16'd37015, 16'd59035, 16'd36906, 16'd57684, 16'd25012, 16'd29077, 16'd36943, 16'd12627, 16'd35076, 16'd61005, 16'd13673, 16'd12963, 16'd63703, 16'd33731, 16'd16570, 16'd30836});
	test_expansion(128'hc7f484fe1450134a91feb8940668e620, {16'd28153, 16'd43607, 16'd50628, 16'd36229, 16'd49342, 16'd18526, 16'd35907, 16'd44933, 16'd61986, 16'd64740, 16'd29345, 16'd30022, 16'd52919, 16'd41115, 16'd38671, 16'd26464, 16'd4217, 16'd5414, 16'd55088, 16'd55084, 16'd37902, 16'd35658, 16'd22606, 16'd17001, 16'd12761, 16'd45261});
	test_expansion(128'hdd3346b69d703a297d815bcc9a64518b, {16'd27196, 16'd8951, 16'd54676, 16'd17965, 16'd6422, 16'd48771, 16'd35704, 16'd36523, 16'd14091, 16'd6879, 16'd46693, 16'd21978, 16'd27307, 16'd54781, 16'd22200, 16'd63460, 16'd15383, 16'd32527, 16'd55759, 16'd57814, 16'd53387, 16'd7984, 16'd34492, 16'd48141, 16'd8344, 16'd41955});
	test_expansion(128'ha3f3e9cc376ae0eafff3080a756a05ed, {16'd60350, 16'd30919, 16'd20061, 16'd41411, 16'd21422, 16'd1815, 16'd14043, 16'd44161, 16'd39348, 16'd4241, 16'd61601, 16'd34404, 16'd39250, 16'd14366, 16'd23763, 16'd49324, 16'd12675, 16'd51195, 16'd27291, 16'd40595, 16'd3590, 16'd45496, 16'd59314, 16'd35134, 16'd35607, 16'd58897});
	test_expansion(128'he25f46db1632a2bb72e9823c4ee168d2, {16'd27552, 16'd43278, 16'd48413, 16'd62419, 16'd6635, 16'd37187, 16'd27445, 16'd12929, 16'd55103, 16'd43557, 16'd956, 16'd35673, 16'd5278, 16'd154, 16'd36646, 16'd63851, 16'd31407, 16'd23398, 16'd7133, 16'd6104, 16'd35781, 16'd51454, 16'd63910, 16'd58945, 16'd25076, 16'd13426});
	test_expansion(128'hf84f11d14b6d73eb938b1fc56d0bd058, {16'd63776, 16'd51834, 16'd18976, 16'd7266, 16'd26766, 16'd17281, 16'd11956, 16'd41498, 16'd17916, 16'd17437, 16'd51189, 16'd52376, 16'd64647, 16'd5167, 16'd1736, 16'd18274, 16'd61254, 16'd59729, 16'd36179, 16'd26397, 16'd16474, 16'd36539, 16'd31768, 16'd28453, 16'd24194, 16'd12301});
	test_expansion(128'hc66c221587cf75adbf8ca2b274b3350a, {16'd25422, 16'd58443, 16'd51918, 16'd62780, 16'd28036, 16'd11492, 16'd51604, 16'd54103, 16'd43548, 16'd28040, 16'd6809, 16'd20617, 16'd50920, 16'd25704, 16'd16323, 16'd55859, 16'd45061, 16'd53114, 16'd49767, 16'd18823, 16'd13775, 16'd13338, 16'd3146, 16'd22174, 16'd15749, 16'd8968});
	test_expansion(128'h1f304bcf1e1c308532ad4f2278d31cf4, {16'd30338, 16'd56077, 16'd10971, 16'd65127, 16'd27452, 16'd22073, 16'd38129, 16'd18982, 16'd8348, 16'd61507, 16'd3064, 16'd41650, 16'd7514, 16'd7, 16'd12085, 16'd28883, 16'd51684, 16'd61106, 16'd3081, 16'd30721, 16'd1492, 16'd8536, 16'd62235, 16'd55213, 16'd21264, 16'd12115});
	test_expansion(128'h09e5169630c35e55b4416b49da1e46dc, {16'd37787, 16'd61558, 16'd49288, 16'd50793, 16'd60260, 16'd356, 16'd19225, 16'd35560, 16'd58344, 16'd59001, 16'd41399, 16'd34572, 16'd27898, 16'd63165, 16'd10906, 16'd64612, 16'd19881, 16'd55569, 16'd59052, 16'd14863, 16'd40336, 16'd10591, 16'd39836, 16'd61947, 16'd19616, 16'd10207});
	test_expansion(128'ha43bd9db3a5b8b6cd159e978185cea16, {16'd13659, 16'd18066, 16'd46550, 16'd18505, 16'd42539, 16'd51122, 16'd7418, 16'd25152, 16'd49142, 16'd7580, 16'd55761, 16'd12051, 16'd41355, 16'd57952, 16'd40390, 16'd43795, 16'd35804, 16'd41416, 16'd34546, 16'd13230, 16'd46148, 16'd21481, 16'd42638, 16'd46506, 16'd47124, 16'd63343});
	test_expansion(128'h0149411cddb9235f76ba508f683b1f06, {16'd62091, 16'd51010, 16'd974, 16'd31623, 16'd51653, 16'd29646, 16'd34982, 16'd30863, 16'd17540, 16'd31636, 16'd62311, 16'd16855, 16'd20821, 16'd44089, 16'd29661, 16'd64402, 16'd30607, 16'd51326, 16'd13731, 16'd25432, 16'd58783, 16'd36561, 16'd9750, 16'd3114, 16'd56773, 16'd32808});
	test_expansion(128'h5c4940f59452b3737356930517ff436e, {16'd11569, 16'd43213, 16'd26637, 16'd53710, 16'd25097, 16'd7063, 16'd25181, 16'd62014, 16'd24075, 16'd6176, 16'd31598, 16'd21983, 16'd19327, 16'd42349, 16'd33630, 16'd20990, 16'd30215, 16'd17672, 16'd3522, 16'd3240, 16'd54013, 16'd65124, 16'd19397, 16'd3955, 16'd12193, 16'd60434});
	test_expansion(128'h78a6c3b930dbc5be425216b6dc317587, {16'd22483, 16'd21008, 16'd41572, 16'd24787, 16'd41137, 16'd45679, 16'd52752, 16'd19054, 16'd33570, 16'd62834, 16'd58691, 16'd422, 16'd51729, 16'd43365, 16'd16798, 16'd41243, 16'd25754, 16'd7757, 16'd50492, 16'd22081, 16'd11629, 16'd62466, 16'd2536, 16'd15312, 16'd48265, 16'd42084});
	test_expansion(128'h8f5e4136cc10c8bb020c21270b020058, {16'd21060, 16'd4794, 16'd44346, 16'd12321, 16'd33170, 16'd26842, 16'd52861, 16'd44357, 16'd38903, 16'd15479, 16'd60525, 16'd29013, 16'd34029, 16'd34640, 16'd64886, 16'd31843, 16'd27451, 16'd1841, 16'd36542, 16'd33498, 16'd7065, 16'd43652, 16'd26353, 16'd7015, 16'd22616, 16'd10004});
	test_expansion(128'he1b74d9c670a28c104416f6c1972df68, {16'd37689, 16'd42742, 16'd24248, 16'd5441, 16'd30917, 16'd64727, 16'd24448, 16'd39085, 16'd41302, 16'd49238, 16'd43722, 16'd44088, 16'd9108, 16'd33279, 16'd42056, 16'd3288, 16'd17190, 16'd34294, 16'd6480, 16'd47544, 16'd36605, 16'd1169, 16'd62065, 16'd25458, 16'd37560, 16'd28649});
	test_expansion(128'hc4a4587b5de11e86ab10c47f9bae94cf, {16'd36257, 16'd7276, 16'd27788, 16'd26337, 16'd26654, 16'd35369, 16'd34022, 16'd6680, 16'd36192, 16'd38611, 16'd4970, 16'd16753, 16'd10586, 16'd9796, 16'd21648, 16'd51634, 16'd9625, 16'd46689, 16'd32861, 16'd50219, 16'd1666, 16'd16726, 16'd48496, 16'd59642, 16'd23210, 16'd26069});
	test_expansion(128'h1ddb8d0bfd864cc869a4e18a9695aa12, {16'd29995, 16'd39254, 16'd8737, 16'd14146, 16'd36730, 16'd6396, 16'd19347, 16'd38780, 16'd11494, 16'd26347, 16'd45039, 16'd52458, 16'd10477, 16'd28311, 16'd4323, 16'd45349, 16'd38640, 16'd15938, 16'd56392, 16'd47461, 16'd19462, 16'd47065, 16'd55963, 16'd43902, 16'd53955, 16'd63202});
	test_expansion(128'h8eddffcf7419aa54f9700fdfe549e35e, {16'd47171, 16'd48552, 16'd18125, 16'd59435, 16'd58135, 16'd35380, 16'd1730, 16'd32675, 16'd50915, 16'd23675, 16'd10525, 16'd62002, 16'd34299, 16'd20004, 16'd35491, 16'd17614, 16'd46448, 16'd38347, 16'd61782, 16'd47620, 16'd18184, 16'd19915, 16'd33531, 16'd47432, 16'd52903, 16'd35377});
	test_expansion(128'h11ed90971612ae7669cbd4289a21ed38, {16'd21004, 16'd10805, 16'd3514, 16'd421, 16'd8812, 16'd46411, 16'd23417, 16'd27711, 16'd39462, 16'd14093, 16'd58653, 16'd44515, 16'd63749, 16'd41554, 16'd40283, 16'd26293, 16'd28371, 16'd42921, 16'd24748, 16'd56297, 16'd46719, 16'd13569, 16'd49349, 16'd36473, 16'd63249, 16'd60658});
	test_expansion(128'h04296efcf1fe260e1188d170e684a83a, {16'd18813, 16'd41759, 16'd25586, 16'd60861, 16'd25976, 16'd55233, 16'd4792, 16'd31781, 16'd15563, 16'd17879, 16'd56421, 16'd28086, 16'd35958, 16'd47608, 16'd56089, 16'd10559, 16'd17428, 16'd59192, 16'd64541, 16'd389, 16'd61356, 16'd41784, 16'd55106, 16'd35347, 16'd58403, 16'd59555});
	test_expansion(128'h9868c2dbc5cabc3cdfa27b3278f59a98, {16'd29906, 16'd9577, 16'd22192, 16'd32173, 16'd44021, 16'd58052, 16'd53925, 16'd12782, 16'd47811, 16'd14788, 16'd6637, 16'd14343, 16'd48564, 16'd33890, 16'd9186, 16'd11069, 16'd30191, 16'd11344, 16'd7475, 16'd61389, 16'd28250, 16'd18490, 16'd19687, 16'd61030, 16'd31023, 16'd24266});
	test_expansion(128'hb6eec0c4ac21ae0c8a05dfb0b0e2fc99, {16'd56362, 16'd29072, 16'd16473, 16'd21970, 16'd45139, 16'd65428, 16'd22156, 16'd40412, 16'd16762, 16'd41801, 16'd11999, 16'd50871, 16'd2479, 16'd51560, 16'd48225, 16'd9792, 16'd27923, 16'd57216, 16'd1881, 16'd27892, 16'd7249, 16'd36892, 16'd22652, 16'd473, 16'd34899, 16'd12362});
	test_expansion(128'h7c3ae4b0c58ab6d8b6a9ce37a829fc95, {16'd45715, 16'd36917, 16'd27974, 16'd50536, 16'd31799, 16'd33796, 16'd10400, 16'd58289, 16'd62516, 16'd23085, 16'd24683, 16'd20439, 16'd34149, 16'd43542, 16'd27802, 16'd28238, 16'd60863, 16'd2102, 16'd62410, 16'd49125, 16'd33105, 16'd13029, 16'd2602, 16'd12888, 16'd29268, 16'd51092});
	test_expansion(128'h218b562d76c4be999b19e29205c6f0da, {16'd40387, 16'd13236, 16'd41527, 16'd22746, 16'd1658, 16'd59044, 16'd18667, 16'd13056, 16'd59870, 16'd65348, 16'd7267, 16'd50583, 16'd48575, 16'd30954, 16'd4180, 16'd15791, 16'd22505, 16'd48334, 16'd16721, 16'd62473, 16'd24480, 16'd41293, 16'd46886, 16'd40466, 16'd19130, 16'd58864});
	test_expansion(128'h832a5163fc99fad802ce144393bb9293, {16'd36957, 16'd61838, 16'd4842, 16'd59428, 16'd15358, 16'd46219, 16'd13651, 16'd9619, 16'd39871, 16'd53875, 16'd57291, 16'd32324, 16'd11122, 16'd64252, 16'd44786, 16'd43047, 16'd31887, 16'd50117, 16'd13950, 16'd54460, 16'd43953, 16'd44748, 16'd29600, 16'd36392, 16'd52783, 16'd6019});
	test_expansion(128'h02b40bea34775d817926b2c75ed7d390, {16'd63650, 16'd21284, 16'd54117, 16'd2347, 16'd36580, 16'd751, 16'd61848, 16'd59917, 16'd9173, 16'd25403, 16'd45214, 16'd25299, 16'd56189, 16'd12622, 16'd17424, 16'd6415, 16'd1450, 16'd54420, 16'd10250, 16'd22549, 16'd19750, 16'd26929, 16'd16574, 16'd13618, 16'd12241, 16'd49650});
	test_expansion(128'h5269b5aa460536b7b9b5d6df36b5496f, {16'd22699, 16'd18459, 16'd4754, 16'd52092, 16'd26156, 16'd63697, 16'd12017, 16'd24084, 16'd49798, 16'd58169, 16'd43377, 16'd27187, 16'd55687, 16'd3611, 16'd48818, 16'd61599, 16'd25951, 16'd16300, 16'd9304, 16'd34644, 16'd46093, 16'd47860, 16'd29980, 16'd59648, 16'd46427, 16'd23842});
	test_expansion(128'h38cf3f23f4e842ec348ab0ba492ec124, {16'd8614, 16'd61258, 16'd42101, 16'd8596, 16'd7234, 16'd24855, 16'd20024, 16'd12791, 16'd19658, 16'd47110, 16'd51518, 16'd49698, 16'd17943, 16'd35340, 16'd65485, 16'd25335, 16'd16098, 16'd57268, 16'd52275, 16'd8345, 16'd63419, 16'd38242, 16'd56431, 16'd49944, 16'd38154, 16'd44768});
	test_expansion(128'h9d687bc7770b45ae1184516b0d2edbc6, {16'd26435, 16'd44289, 16'd21866, 16'd24278, 16'd60286, 16'd62122, 16'd8118, 16'd34001, 16'd395, 16'd46508, 16'd53670, 16'd25719, 16'd50787, 16'd38691, 16'd25389, 16'd485, 16'd62431, 16'd30054, 16'd7477, 16'd4085, 16'd20032, 16'd9363, 16'd11586, 16'd64777, 16'd60095, 16'd28561});
	test_expansion(128'h0cd64af93cc4ca919ee01d5611fd50ac, {16'd53414, 16'd18441, 16'd22440, 16'd40321, 16'd33828, 16'd2819, 16'd6772, 16'd16078, 16'd64106, 16'd62618, 16'd39030, 16'd28691, 16'd13502, 16'd52494, 16'd11563, 16'd4288, 16'd21321, 16'd36075, 16'd285, 16'd33742, 16'd24680, 16'd58630, 16'd50643, 16'd30091, 16'd45236, 16'd41604});
	test_expansion(128'h2d36148fedbd8ddb8b19bab4f3116814, {16'd34678, 16'd20107, 16'd14369, 16'd16660, 16'd1446, 16'd50494, 16'd21932, 16'd38937, 16'd39246, 16'd24249, 16'd5565, 16'd50733, 16'd28963, 16'd7462, 16'd1639, 16'd20116, 16'd38805, 16'd6143, 16'd64745, 16'd36032, 16'd11760, 16'd16054, 16'd21417, 16'd28284, 16'd63812, 16'd20243});
	test_expansion(128'hd9a09d0a48d175b0459059d3e903978b, {16'd44315, 16'd14277, 16'd25212, 16'd31266, 16'd20868, 16'd63251, 16'd19090, 16'd37368, 16'd27281, 16'd7742, 16'd59662, 16'd60215, 16'd15797, 16'd28448, 16'd1912, 16'd464, 16'd4534, 16'd32097, 16'd61561, 16'd55673, 16'd58330, 16'd43708, 16'd27457, 16'd1081, 16'd50454, 16'd11496});
	test_expansion(128'h2cb74acb5c70b8068b26670312074b10, {16'd2873, 16'd47242, 16'd17414, 16'd48292, 16'd22599, 16'd26279, 16'd2983, 16'd12802, 16'd30335, 16'd53216, 16'd46478, 16'd55407, 16'd53882, 16'd25788, 16'd53610, 16'd31351, 16'd59119, 16'd27879, 16'd40301, 16'd2178, 16'd65189, 16'd36434, 16'd25360, 16'd62721, 16'd59036, 16'd17837});
	test_expansion(128'h45d5b7a60814245e4510a01453ffef22, {16'd6543, 16'd37675, 16'd22862, 16'd22697, 16'd16056, 16'd52533, 16'd41358, 16'd11350, 16'd50258, 16'd1899, 16'd12725, 16'd36955, 16'd60022, 16'd11481, 16'd15480, 16'd41274, 16'd28724, 16'd61330, 16'd33600, 16'd25009, 16'd27555, 16'd31834, 16'd49626, 16'd17899, 16'd42143, 16'd22203});
	test_expansion(128'he5f36cbb03806063e1a0ce1694c5bd00, {16'd41989, 16'd65477, 16'd37210, 16'd60333, 16'd2913, 16'd11812, 16'd14430, 16'd6197, 16'd14605, 16'd20641, 16'd58857, 16'd23013, 16'd9189, 16'd44618, 16'd54990, 16'd27724, 16'd18421, 16'd45843, 16'd49024, 16'd51389, 16'd8158, 16'd59398, 16'd47415, 16'd2180, 16'd63991, 16'd40882});
	test_expansion(128'he56e355f254890b3e5448468be105c47, {16'd13759, 16'd59548, 16'd23765, 16'd27991, 16'd56054, 16'd30126, 16'd25136, 16'd39209, 16'd60949, 16'd22101, 16'd28503, 16'd17883, 16'd42905, 16'd635, 16'd22081, 16'd45213, 16'd55202, 16'd16556, 16'd46485, 16'd21183, 16'd42745, 16'd51805, 16'd15615, 16'd31835, 16'd54561, 16'd56312});
	test_expansion(128'h9158cb594819f6b334414300e0d02a1d, {16'd19023, 16'd59624, 16'd45193, 16'd26175, 16'd54934, 16'd54627, 16'd46444, 16'd46887, 16'd29696, 16'd41183, 16'd40451, 16'd10927, 16'd26242, 16'd62299, 16'd37459, 16'd24142, 16'd38272, 16'd7620, 16'd1032, 16'd41407, 16'd1424, 16'd55907, 16'd12376, 16'd48292, 16'd46194, 16'd45402});
	test_expansion(128'h77d0842ed6f719ee3a00e28e749e7ace, {16'd58076, 16'd16705, 16'd873, 16'd53833, 16'd53109, 16'd58015, 16'd25198, 16'd62930, 16'd35792, 16'd62684, 16'd61321, 16'd1842, 16'd53285, 16'd21018, 16'd36187, 16'd24464, 16'd1319, 16'd24018, 16'd12441, 16'd7289, 16'd52759, 16'd9813, 16'd40773, 16'd53327, 16'd59370, 16'd60423});
	test_expansion(128'had0aec1fff75a35158d67c5103f4e465, {16'd3521, 16'd3440, 16'd12326, 16'd52014, 16'd29426, 16'd2077, 16'd49110, 16'd43494, 16'd22121, 16'd28668, 16'd61005, 16'd23961, 16'd41209, 16'd60360, 16'd29915, 16'd54571, 16'd47496, 16'd18361, 16'd37270, 16'd60135, 16'd43265, 16'd41, 16'd39249, 16'd19587, 16'd25948, 16'd3396});
	test_expansion(128'h9faac317b4878ef4d905b55e390021e5, {16'd16384, 16'd42861, 16'd25178, 16'd34421, 16'd48969, 16'd14421, 16'd5428, 16'd60425, 16'd19655, 16'd13942, 16'd54591, 16'd31192, 16'd8590, 16'd57528, 16'd8179, 16'd19428, 16'd64137, 16'd34893, 16'd28225, 16'd13117, 16'd13027, 16'd45843, 16'd64612, 16'd10668, 16'd1378, 16'd40205});
	test_expansion(128'hd9cdfd3d86b9e1ce662c6c8de6bd68bb, {16'd6261, 16'd3576, 16'd32870, 16'd45370, 16'd20059, 16'd6974, 16'd7199, 16'd2605, 16'd18245, 16'd6253, 16'd27704, 16'd61613, 16'd34805, 16'd36445, 16'd39833, 16'd24847, 16'd50890, 16'd30789, 16'd3147, 16'd49166, 16'd56521, 16'd16083, 16'd23424, 16'd52911, 16'd42349, 16'd49237});
	test_expansion(128'he1e578c51a41de4b336544803fb9d403, {16'd22073, 16'd58409, 16'd12879, 16'd52552, 16'd61500, 16'd19569, 16'd6004, 16'd10899, 16'd27618, 16'd56637, 16'd3627, 16'd25874, 16'd57412, 16'd26580, 16'd32478, 16'd25603, 16'd41911, 16'd55056, 16'd19411, 16'd15428, 16'd2393, 16'd48013, 16'd47341, 16'd52436, 16'd41869, 16'd17818});
	test_expansion(128'h2e17974552a0dc513aae6ccb0b896292, {16'd44980, 16'd29575, 16'd44639, 16'd46695, 16'd58695, 16'd10501, 16'd48467, 16'd51841, 16'd22590, 16'd57531, 16'd37578, 16'd6349, 16'd43562, 16'd29699, 16'd54173, 16'd42810, 16'd38204, 16'd50132, 16'd58444, 16'd44638, 16'd37881, 16'd47453, 16'd40753, 16'd3758, 16'd52380, 16'd36628});
	test_expansion(128'h390f0040a8922c829b3b0282dca17168, {16'd34190, 16'd64722, 16'd64255, 16'd11372, 16'd51475, 16'd49878, 16'd65111, 16'd18812, 16'd59302, 16'd3241, 16'd21557, 16'd209, 16'd29395, 16'd52070, 16'd54443, 16'd61347, 16'd57406, 16'd29860, 16'd47236, 16'd58209, 16'd8181, 16'd41363, 16'd9919, 16'd36538, 16'd17935, 16'd19127});
	test_expansion(128'h1ac741d6d29d906e73c1e49cafbfd6ac, {16'd31577, 16'd23339, 16'd5252, 16'd49846, 16'd63536, 16'd46383, 16'd11173, 16'd35319, 16'd29327, 16'd5501, 16'd12189, 16'd5189, 16'd60835, 16'd6448, 16'd15114, 16'd17574, 16'd42927, 16'd21882, 16'd63428, 16'd1459, 16'd22775, 16'd15021, 16'd32878, 16'd41910, 16'd18677, 16'd38046});
	test_expansion(128'h5cfd34237da139f3ae1e4909799e826d, {16'd51449, 16'd49468, 16'd51451, 16'd64237, 16'd52700, 16'd7028, 16'd17542, 16'd37101, 16'd42509, 16'd21611, 16'd28908, 16'd11930, 16'd64415, 16'd11620, 16'd26733, 16'd11244, 16'd62181, 16'd26570, 16'd42468, 16'd1757, 16'd11256, 16'd58395, 16'd22358, 16'd47514, 16'd32326, 16'd49481});
	test_expansion(128'hcce6d11886107663723cbba58095f7fa, {16'd50475, 16'd9747, 16'd15721, 16'd30000, 16'd18271, 16'd5661, 16'd11979, 16'd50244, 16'd47163, 16'd20263, 16'd17190, 16'd32252, 16'd39023, 16'd49568, 16'd30788, 16'd31830, 16'd31826, 16'd9225, 16'd11418, 16'd22993, 16'd49248, 16'd28166, 16'd53602, 16'd61937, 16'd9325, 16'd25509});
	test_expansion(128'h13f9572ee65cf61499a626e35855ed92, {16'd10789, 16'd40693, 16'd39088, 16'd34658, 16'd52390, 16'd65004, 16'd6542, 16'd25183, 16'd16122, 16'd6266, 16'd10666, 16'd59437, 16'd25811, 16'd54435, 16'd23493, 16'd55246, 16'd15506, 16'd26666, 16'd16819, 16'd5875, 16'd4744, 16'd63692, 16'd33168, 16'd63753, 16'd22744, 16'd58760});
	test_expansion(128'h68a7d6ea24e7310b8deac7c7770022b6, {16'd48575, 16'd4905, 16'd9210, 16'd4609, 16'd47295, 16'd44301, 16'd4944, 16'd45416, 16'd55103, 16'd23608, 16'd24864, 16'd55521, 16'd7258, 16'd12894, 16'd63391, 16'd62471, 16'd35945, 16'd26654, 16'd22605, 16'd22016, 16'd55019, 16'd62119, 16'd11603, 16'd58364, 16'd10663, 16'd12447});
	test_expansion(128'h08f02ae0726d11b865a2c022f039da93, {16'd19073, 16'd5625, 16'd19150, 16'd18802, 16'd15538, 16'd16297, 16'd50489, 16'd48107, 16'd46943, 16'd58679, 16'd34822, 16'd36193, 16'd41993, 16'd19111, 16'd31143, 16'd50045, 16'd27147, 16'd21, 16'd55498, 16'd31231, 16'd39690, 16'd48175, 16'd51668, 16'd19778, 16'd46436, 16'd61358});
	test_expansion(128'hfa3a2d4f0ac2cea45e280265fd938cc0, {16'd61876, 16'd55848, 16'd35636, 16'd37627, 16'd33693, 16'd278, 16'd28494, 16'd11917, 16'd5975, 16'd19608, 16'd61586, 16'd10767, 16'd5735, 16'd49993, 16'd44151, 16'd4021, 16'd1269, 16'd44650, 16'd2262, 16'd27618, 16'd22041, 16'd24163, 16'd14529, 16'd36570, 16'd15296, 16'd52785});
	test_expansion(128'h6d075ea35d38c5df5b14e5e9b1c5b4b1, {16'd49501, 16'd24518, 16'd39209, 16'd47098, 16'd12436, 16'd12497, 16'd61865, 16'd53574, 16'd33164, 16'd32007, 16'd1645, 16'd17674, 16'd49170, 16'd47292, 16'd37188, 16'd54232, 16'd61165, 16'd64846, 16'd47142, 16'd41543, 16'd22810, 16'd43277, 16'd60212, 16'd53851, 16'd2664, 16'd39148});
	test_expansion(128'haae122025530f263e9005c99f6183650, {16'd46173, 16'd9514, 16'd23077, 16'd56162, 16'd5329, 16'd61168, 16'd37736, 16'd13356, 16'd55622, 16'd59269, 16'd43003, 16'd5250, 16'd6396, 16'd34787, 16'd6561, 16'd28884, 16'd3521, 16'd2592, 16'd6025, 16'd4525, 16'd12066, 16'd28462, 16'd20147, 16'd25732, 16'd6908, 16'd32808});
	test_expansion(128'h7f672e15e426b172882a913a51c6e45e, {16'd6112, 16'd47783, 16'd6643, 16'd26409, 16'd24533, 16'd5195, 16'd16321, 16'd39679, 16'd58074, 16'd2545, 16'd57719, 16'd44565, 16'd39129, 16'd25065, 16'd43891, 16'd8618, 16'd9109, 16'd11681, 16'd44321, 16'd31823, 16'd33590, 16'd56091, 16'd11434, 16'd63471, 16'd2583, 16'd25817});
	test_expansion(128'h077fcaeda636aa4eeab1f8548064e2b5, {16'd23280, 16'd58394, 16'd12226, 16'd18403, 16'd17583, 16'd46764, 16'd35188, 16'd44047, 16'd19145, 16'd5327, 16'd40027, 16'd49415, 16'd28175, 16'd9819, 16'd14351, 16'd25707, 16'd43767, 16'd34185, 16'd49161, 16'd17636, 16'd24980, 16'd8927, 16'd13730, 16'd21355, 16'd4229, 16'd56869});
	test_expansion(128'hd401bb9d4c0caf0e90ae722f648f2b8f, {16'd41975, 16'd62915, 16'd26861, 16'd46968, 16'd24578, 16'd20017, 16'd28526, 16'd46535, 16'd24374, 16'd26366, 16'd49861, 16'd26529, 16'd61073, 16'd40670, 16'd16130, 16'd674, 16'd46659, 16'd9195, 16'd52335, 16'd35609, 16'd42967, 16'd33241, 16'd19853, 16'd34071, 16'd15511, 16'd14090});
	test_expansion(128'h35ef228a95f498c73c110719900e0eeb, {16'd10919, 16'd57710, 16'd24941, 16'd14510, 16'd51129, 16'd3887, 16'd4877, 16'd3652, 16'd4011, 16'd41319, 16'd39029, 16'd6913, 16'd11945, 16'd35064, 16'd58382, 16'd41375, 16'd14279, 16'd32884, 16'd58959, 16'd42904, 16'd32171, 16'd41744, 16'd30582, 16'd22487, 16'd17156, 16'd13388});
	test_expansion(128'h24c65f315d23dd2da5fe6dd341ac3684, {16'd44846, 16'd54239, 16'd51120, 16'd61750, 16'd58552, 16'd12073, 16'd58860, 16'd10218, 16'd34362, 16'd11618, 16'd43276, 16'd8199, 16'd10783, 16'd50413, 16'd39361, 16'd60590, 16'd10434, 16'd911, 16'd61387, 16'd52195, 16'd21099, 16'd37121, 16'd38474, 16'd16087, 16'd57857, 16'd1862});
	test_expansion(128'he95626f71db7a2a8a22a5424209f7273, {16'd9313, 16'd52640, 16'd39411, 16'd20820, 16'd15887, 16'd64714, 16'd17143, 16'd3068, 16'd34356, 16'd53841, 16'd28217, 16'd23929, 16'd20079, 16'd64533, 16'd5175, 16'd60966, 16'd53915, 16'd32775, 16'd14427, 16'd43172, 16'd55393, 16'd38048, 16'd52091, 16'd9361, 16'd1537, 16'd54173});
	test_expansion(128'hfd5488428acbb5298e2221dd3d4de7b7, {16'd22078, 16'd13583, 16'd24819, 16'd33814, 16'd57575, 16'd9737, 16'd42655, 16'd27723, 16'd22439, 16'd50351, 16'd3241, 16'd19923, 16'd32838, 16'd20707, 16'd29172, 16'd50644, 16'd38482, 16'd55861, 16'd5787, 16'd6986, 16'd19919, 16'd28789, 16'd19904, 16'd20897, 16'd53136, 16'd14791});
	test_expansion(128'ha7f87906522746ecfa2bb362d91ffed3, {16'd13934, 16'd21014, 16'd22142, 16'd41362, 16'd12940, 16'd36201, 16'd56642, 16'd19129, 16'd49163, 16'd20275, 16'd1333, 16'd6829, 16'd51416, 16'd17144, 16'd15, 16'd56246, 16'd48357, 16'd32913, 16'd38283, 16'd41648, 16'd7351, 16'd4048, 16'd42118, 16'd48059, 16'd44547, 16'd36491});
	test_expansion(128'h171c6802957c9f8e3163d3006076ab03, {16'd12620, 16'd31996, 16'd37138, 16'd18582, 16'd6744, 16'd52378, 16'd48725, 16'd6038, 16'd55373, 16'd62714, 16'd59562, 16'd34409, 16'd39191, 16'd38316, 16'd64131, 16'd62390, 16'd44355, 16'd30543, 16'd63924, 16'd50018, 16'd33183, 16'd38223, 16'd51766, 16'd667, 16'd37179, 16'd15796});
	test_expansion(128'h5c045e0d2d408909f46323221f847bd4, {16'd11976, 16'd45088, 16'd54526, 16'd3149, 16'd57167, 16'd45245, 16'd21723, 16'd29933, 16'd61628, 16'd42271, 16'd23491, 16'd25618, 16'd11523, 16'd14380, 16'd57032, 16'd59447, 16'd50469, 16'd12371, 16'd1290, 16'd7799, 16'd2126, 16'd10403, 16'd19279, 16'd10937, 16'd14842, 16'd22434});
	test_expansion(128'hc59f5feb5838f38c77cbd824570bb7d8, {16'd59872, 16'd13618, 16'd51396, 16'd18964, 16'd64693, 16'd41086, 16'd32766, 16'd13807, 16'd32266, 16'd52140, 16'd54702, 16'd41600, 16'd3286, 16'd30179, 16'd9777, 16'd2830, 16'd26993, 16'd42949, 16'd4374, 16'd4606, 16'd51506, 16'd45020, 16'd27628, 16'd37703, 16'd28887, 16'd42636});
	test_expansion(128'h4b48c8a12f8d740cdd78d12cccb38967, {16'd53228, 16'd17436, 16'd17909, 16'd54457, 16'd17117, 16'd27669, 16'd62236, 16'd33659, 16'd42429, 16'd3195, 16'd36258, 16'd10635, 16'd54082, 16'd14525, 16'd43780, 16'd26623, 16'd42545, 16'd22763, 16'd42558, 16'd44368, 16'd7840, 16'd44247, 16'd20504, 16'd24376, 16'd30684, 16'd12006});
	test_expansion(128'h1431606cc4877c1e6d1bb566fe06f1ef, {16'd36707, 16'd11379, 16'd3289, 16'd17883, 16'd53632, 16'd6715, 16'd48772, 16'd47745, 16'd47053, 16'd807, 16'd27869, 16'd6835, 16'd25575, 16'd16972, 16'd61129, 16'd14944, 16'd8179, 16'd45766, 16'd20678, 16'd18883, 16'd48223, 16'd46625, 16'd28273, 16'd36831, 16'd15223, 16'd63765});
	test_expansion(128'h804fe8cd0e77e41eb6887c30d9bfbd4f, {16'd14446, 16'd63067, 16'd32240, 16'd12373, 16'd24821, 16'd50141, 16'd28896, 16'd10878, 16'd41276, 16'd16156, 16'd12677, 16'd23725, 16'd26672, 16'd28458, 16'd44976, 16'd37766, 16'd7646, 16'd18269, 16'd42107, 16'd7454, 16'd36131, 16'd11336, 16'd22345, 16'd20419, 16'd14024, 16'd1817});
	test_expansion(128'hb78f67638091907e325431bf2ce6db42, {16'd37456, 16'd45678, 16'd51399, 16'd62258, 16'd45340, 16'd48927, 16'd43857, 16'd45824, 16'd36777, 16'd24641, 16'd47564, 16'd65501, 16'd27154, 16'd27711, 16'd42058, 16'd41377, 16'd34716, 16'd52798, 16'd17069, 16'd4190, 16'd47809, 16'd12328, 16'd28154, 16'd576, 16'd35209, 16'd60005});
	test_expansion(128'h61ce0444bc04a1fab2327568facfe39f, {16'd22081, 16'd64865, 16'd1255, 16'd26423, 16'd59480, 16'd34757, 16'd37352, 16'd20652, 16'd35255, 16'd48924, 16'd37497, 16'd1292, 16'd26418, 16'd34712, 16'd3224, 16'd7058, 16'd32566, 16'd55772, 16'd37792, 16'd65433, 16'd21154, 16'd62969, 16'd44701, 16'd35996, 16'd9358, 16'd64986});
	test_expansion(128'h5e7febc958314840784500e6596bd48d, {16'd9162, 16'd12858, 16'd63225, 16'd29682, 16'd3055, 16'd49598, 16'd20484, 16'd34550, 16'd2772, 16'd51329, 16'd20702, 16'd12998, 16'd32671, 16'd34571, 16'd58226, 16'd42242, 16'd39490, 16'd40641, 16'd36133, 16'd25883, 16'd48690, 16'd1945, 16'd29835, 16'd26209, 16'd17148, 16'd17231});
	test_expansion(128'h51616c02a929faa062c7da4a47036f7f, {16'd36752, 16'd45064, 16'd54785, 16'd57560, 16'd16923, 16'd32617, 16'd65473, 16'd38680, 16'd42444, 16'd61094, 16'd12276, 16'd25004, 16'd17500, 16'd31054, 16'd26840, 16'd53446, 16'd8091, 16'd50732, 16'd63471, 16'd12315, 16'd6109, 16'd8001, 16'd3587, 16'd41903, 16'd26587, 16'd13025});
	test_expansion(128'hf4a14b3e71f5d3fe6b40ad5a18858293, {16'd4498, 16'd64103, 16'd21004, 16'd60480, 16'd13523, 16'd40856, 16'd59337, 16'd21060, 16'd3315, 16'd34139, 16'd59708, 16'd42235, 16'd33242, 16'd17669, 16'd4678, 16'd34879, 16'd39170, 16'd40254, 16'd20378, 16'd46338, 16'd64615, 16'd10778, 16'd54420, 16'd14207, 16'd11886, 16'd11998});
	test_expansion(128'hc8620c0ce1c7ef8d8785ca2b3e007aec, {16'd30949, 16'd23251, 16'd39206, 16'd15490, 16'd55471, 16'd29853, 16'd35549, 16'd29227, 16'd5100, 16'd21520, 16'd37605, 16'd53305, 16'd49257, 16'd65061, 16'd23777, 16'd56681, 16'd58859, 16'd9915, 16'd33727, 16'd15286, 16'd1159, 16'd50963, 16'd25997, 16'd59395, 16'd2100, 16'd42261});
	test_expansion(128'hed5b1bcc24a97f13ce38d923ea35ec33, {16'd10248, 16'd9698, 16'd57286, 16'd31039, 16'd2637, 16'd6745, 16'd7517, 16'd58159, 16'd31157, 16'd28570, 16'd57306, 16'd23820, 16'd41061, 16'd52763, 16'd45890, 16'd58869, 16'd9877, 16'd44529, 16'd31104, 16'd15163, 16'd41060, 16'd47667, 16'd54614, 16'd14710, 16'd34850, 16'd54823});
	test_expansion(128'h764d0f50da0044d14c256a34b96c8fa7, {16'd45165, 16'd9255, 16'd62561, 16'd55546, 16'd9900, 16'd20454, 16'd56181, 16'd3563, 16'd62270, 16'd62911, 16'd56619, 16'd5093, 16'd37663, 16'd1177, 16'd3377, 16'd27879, 16'd31252, 16'd16326, 16'd30556, 16'd49229, 16'd7510, 16'd38134, 16'd169, 16'd23396, 16'd35764, 16'd24952});
	test_expansion(128'hd92cdd88edbe7c71164002722d58dbb2, {16'd30174, 16'd14484, 16'd47884, 16'd27724, 16'd63960, 16'd38223, 16'd46221, 16'd37813, 16'd59651, 16'd34019, 16'd875, 16'd4117, 16'd32619, 16'd1543, 16'd55565, 16'd49481, 16'd57093, 16'd35426, 16'd62769, 16'd5415, 16'd24644, 16'd43991, 16'd47227, 16'd4598, 16'd37184, 16'd31988});
	test_expansion(128'h60a17f847b9b275ab9f6a42c484cd959, {16'd13717, 16'd44107, 16'd60198, 16'd55785, 16'd22008, 16'd33087, 16'd54311, 16'd48032, 16'd22273, 16'd17742, 16'd16800, 16'd63153, 16'd19250, 16'd17736, 16'd46035, 16'd18776, 16'd34984, 16'd21472, 16'd29600, 16'd2389, 16'd5311, 16'd15162, 16'd20783, 16'd59559, 16'd43433, 16'd20268});
	test_expansion(128'h39a0211a94b9970dac6eed8926b403bf, {16'd16285, 16'd58865, 16'd63296, 16'd11019, 16'd22306, 16'd28833, 16'd38297, 16'd57274, 16'd42623, 16'd17493, 16'd50229, 16'd28274, 16'd39658, 16'd47980, 16'd52233, 16'd53298, 16'd9184, 16'd26617, 16'd61502, 16'd38694, 16'd10030, 16'd51013, 16'd12397, 16'd34098, 16'd46717, 16'd19399});
	test_expansion(128'hca63eecbc4e98134dab69dfd38ae5c10, {16'd47773, 16'd26421, 16'd2570, 16'd33962, 16'd7416, 16'd35053, 16'd13475, 16'd46368, 16'd62605, 16'd20954, 16'd5997, 16'd39468, 16'd39035, 16'd33863, 16'd60962, 16'd61829, 16'd49114, 16'd18658, 16'd8026, 16'd52198, 16'd18642, 16'd2031, 16'd43583, 16'd31614, 16'd10006, 16'd5040});
	test_expansion(128'hb5bb7753c7168958d9cf8a32954a242a, {16'd45117, 16'd45556, 16'd30983, 16'd9887, 16'd58727, 16'd24629, 16'd6996, 16'd40065, 16'd39820, 16'd31608, 16'd23808, 16'd50678, 16'd14267, 16'd63809, 16'd40193, 16'd40471, 16'd36354, 16'd47830, 16'd14095, 16'd47394, 16'd49075, 16'd51317, 16'd40697, 16'd12687, 16'd37082, 16'd46869});
	test_expansion(128'hf83db4763b2856192b90e6b21e85f113, {16'd1739, 16'd53110, 16'd27088, 16'd6642, 16'd16660, 16'd42866, 16'd19497, 16'd9690, 16'd7421, 16'd53040, 16'd10491, 16'd32226, 16'd19784, 16'd10642, 16'd25313, 16'd44292, 16'd48286, 16'd28855, 16'd23369, 16'd3651, 16'd4721, 16'd49922, 16'd38337, 16'd62556, 16'd51302, 16'd29226});
	test_expansion(128'h249a7bfdc24a3d0cb3e0a83632718074, {16'd47287, 16'd869, 16'd40612, 16'd458, 16'd31642, 16'd60944, 16'd2982, 16'd57053, 16'd1013, 16'd21677, 16'd447, 16'd57028, 16'd23738, 16'd54070, 16'd41164, 16'd25876, 16'd35442, 16'd63232, 16'd22233, 16'd14392, 16'd46683, 16'd17560, 16'd11887, 16'd17569, 16'd31970, 16'd4669});
	test_expansion(128'h79271bf0fbf140ad30bddcc1a1a8eae9, {16'd59045, 16'd29390, 16'd35282, 16'd59624, 16'd48909, 16'd19992, 16'd37698, 16'd4515, 16'd45123, 16'd64998, 16'd45912, 16'd51866, 16'd34779, 16'd4058, 16'd26906, 16'd12706, 16'd16593, 16'd13945, 16'd55853, 16'd4742, 16'd21404, 16'd61665, 16'd11188, 16'd39890, 16'd39288, 16'd48940});
	test_expansion(128'hc45dd66e82ac7ee40b737f05037ec2fb, {16'd37585, 16'd27131, 16'd42951, 16'd49457, 16'd41548, 16'd57238, 16'd28446, 16'd59179, 16'd19957, 16'd56406, 16'd51839, 16'd30794, 16'd27206, 16'd14715, 16'd37899, 16'd56789, 16'd47473, 16'd46891, 16'd36267, 16'd31528, 16'd33927, 16'd60029, 16'd50522, 16'd14104, 16'd25854, 16'd33854});
	test_expansion(128'h4587276dfc5cf7e1f6a390ee0e3ae40d, {16'd52473, 16'd56582, 16'd37204, 16'd63430, 16'd29755, 16'd10070, 16'd39930, 16'd16866, 16'd24738, 16'd23664, 16'd7689, 16'd24230, 16'd53112, 16'd25606, 16'd61853, 16'd62982, 16'd58056, 16'd65464, 16'd54164, 16'd15022, 16'd10087, 16'd57308, 16'd46300, 16'd3557, 16'd60700, 16'd11751});
	test_expansion(128'h01507e5d578ec0114f13e5df9a782d47, {16'd51382, 16'd29362, 16'd23081, 16'd10512, 16'd37256, 16'd11218, 16'd7647, 16'd3560, 16'd9185, 16'd61126, 16'd31216, 16'd64821, 16'd41868, 16'd9235, 16'd7956, 16'd52694, 16'd29843, 16'd5928, 16'd62063, 16'd14320, 16'd31518, 16'd55737, 16'd59874, 16'd45489, 16'd42952, 16'd6904});
	test_expansion(128'h0b3df55e4fecfcf8158b4bfe492ad86d, {16'd40418, 16'd45098, 16'd50016, 16'd35667, 16'd51471, 16'd11425, 16'd21155, 16'd5528, 16'd40137, 16'd39794, 16'd7544, 16'd49208, 16'd29174, 16'd2702, 16'd6836, 16'd2387, 16'd21570, 16'd50240, 16'd27742, 16'd12499, 16'd15623, 16'd6528, 16'd10606, 16'd14408, 16'd11389, 16'd18139});
	test_expansion(128'h980a577c5767f67c30721132cdc3ebb0, {16'd38723, 16'd6520, 16'd36231, 16'd15204, 16'd13620, 16'd55497, 16'd53145, 16'd52741, 16'd10791, 16'd19060, 16'd14005, 16'd42114, 16'd3431, 16'd29804, 16'd39412, 16'd31173, 16'd40237, 16'd60004, 16'd52925, 16'd20288, 16'd18152, 16'd6535, 16'd12186, 16'd53083, 16'd3058, 16'd14024});
	test_expansion(128'hf9b6048a8043713b3624998be4e91869, {16'd54865, 16'd49433, 16'd12747, 16'd1248, 16'd57140, 16'd24073, 16'd8657, 16'd10521, 16'd39616, 16'd45321, 16'd12061, 16'd27713, 16'd28830, 16'd64984, 16'd51015, 16'd62309, 16'd20836, 16'd35980, 16'd46265, 16'd13705, 16'd35495, 16'd19554, 16'd45446, 16'd39979, 16'd49833, 16'd57284});
	test_expansion(128'hcf8fdd86abd5dcd0fb286710620fa32a, {16'd12833, 16'd46743, 16'd60442, 16'd15749, 16'd34639, 16'd27487, 16'd58214, 16'd43447, 16'd18639, 16'd2896, 16'd9734, 16'd23095, 16'd14593, 16'd32387, 16'd22450, 16'd62767, 16'd9672, 16'd40075, 16'd58352, 16'd23808, 16'd61443, 16'd7458, 16'd52838, 16'd1063, 16'd29989, 16'd15109});
	test_expansion(128'h6b852daebfbef7cbbe2fecedc96b4189, {16'd47134, 16'd47371, 16'd40253, 16'd30725, 16'd64830, 16'd56768, 16'd17740, 16'd63311, 16'd60254, 16'd51123, 16'd28948, 16'd21275, 16'd57562, 16'd4695, 16'd11230, 16'd41703, 16'd13953, 16'd54708, 16'd4515, 16'd56067, 16'd24797, 16'd57980, 16'd57659, 16'd11118, 16'd62620, 16'd49035});
	test_expansion(128'h4188de16262ad1c73bd030a631e37736, {16'd31039, 16'd15046, 16'd21616, 16'd58096, 16'd62912, 16'd63802, 16'd43758, 16'd6149, 16'd48356, 16'd19918, 16'd56364, 16'd10791, 16'd23465, 16'd32002, 16'd50652, 16'd37883, 16'd57559, 16'd2842, 16'd785, 16'd35590, 16'd45124, 16'd558, 16'd41240, 16'd257, 16'd7576, 16'd61109});
	test_expansion(128'hafc9db831a5da2fb6e94475b37e5b50c, {16'd568, 16'd14404, 16'd13691, 16'd64711, 16'd57910, 16'd38028, 16'd25417, 16'd35725, 16'd23120, 16'd55685, 16'd58494, 16'd31493, 16'd40319, 16'd47765, 16'd53519, 16'd51005, 16'd20978, 16'd10717, 16'd64106, 16'd43849, 16'd52104, 16'd60340, 16'd14024, 16'd7167, 16'd52290, 16'd1822});
	test_expansion(128'h9e7e5eb94b39313d59380e43ec43dc43, {16'd7476, 16'd15229, 16'd329, 16'd3822, 16'd21896, 16'd64279, 16'd38917, 16'd41191, 16'd39650, 16'd52902, 16'd59323, 16'd41925, 16'd53177, 16'd19135, 16'd46983, 16'd2755, 16'd57840, 16'd4632, 16'd39151, 16'd62, 16'd3988, 16'd11522, 16'd38664, 16'd39577, 16'd27197, 16'd60811});
	test_expansion(128'h0843520211592a5c26d32900fcc7f49f, {16'd23705, 16'd15713, 16'd47009, 16'd49622, 16'd8490, 16'd51289, 16'd52033, 16'd34112, 16'd471, 16'd12714, 16'd49036, 16'd19631, 16'd5054, 16'd10249, 16'd31779, 16'd3646, 16'd9457, 16'd28890, 16'd53057, 16'd48081, 16'd16705, 16'd5101, 16'd20782, 16'd20953, 16'd23352, 16'd14324});
	test_expansion(128'h1ab8fc39ebdc9992fb5977e9f73a1609, {16'd17030, 16'd25246, 16'd39736, 16'd60682, 16'd34442, 16'd1958, 16'd17148, 16'd16058, 16'd39545, 16'd36723, 16'd20673, 16'd28635, 16'd58639, 16'd56095, 16'd58191, 16'd54679, 16'd44545, 16'd62513, 16'd14030, 16'd60687, 16'd59902, 16'd23619, 16'd44148, 16'd41346, 16'd52232, 16'd49287});
	test_expansion(128'h5ed16fe3df656f11ed41ed920a9585bb, {16'd62989, 16'd32010, 16'd5428, 16'd38523, 16'd40966, 16'd38342, 16'd3855, 16'd3499, 16'd56730, 16'd25760, 16'd35924, 16'd58057, 16'd33554, 16'd22347, 16'd42536, 16'd33774, 16'd15167, 16'd32821, 16'd16536, 16'd61083, 16'd14451, 16'd47088, 16'd40349, 16'd53735, 16'd45133, 16'd21624});
	test_expansion(128'h6f5580a246dcfd5cdf132844025aff07, {16'd50496, 16'd34503, 16'd45961, 16'd15245, 16'd59721, 16'd14767, 16'd31107, 16'd37875, 16'd50689, 16'd29393, 16'd36914, 16'd5113, 16'd20790, 16'd22561, 16'd18718, 16'd3142, 16'd7354, 16'd31619, 16'd7215, 16'd48329, 16'd44821, 16'd4822, 16'd14459, 16'd28167, 16'd50038, 16'd7020});
	test_expansion(128'hf81a6c9d22a4ba543f62966d22eaa798, {16'd41813, 16'd35322, 16'd49105, 16'd24690, 16'd26641, 16'd60565, 16'd43949, 16'd17243, 16'd29235, 16'd26675, 16'd42534, 16'd5523, 16'd57653, 16'd54937, 16'd40318, 16'd11361, 16'd13138, 16'd35666, 16'd42997, 16'd17660, 16'd49824, 16'd65052, 16'd35529, 16'd3562, 16'd38416, 16'd23186});
	test_expansion(128'hda1ca34d11616540250bafdaa2c0d234, {16'd41429, 16'd4727, 16'd57044, 16'd48635, 16'd4437, 16'd60764, 16'd47524, 16'd31215, 16'd9792, 16'd13667, 16'd40101, 16'd47249, 16'd15151, 16'd37588, 16'd675, 16'd55526, 16'd60723, 16'd30228, 16'd12687, 16'd17897, 16'd10340, 16'd16726, 16'd51536, 16'd58937, 16'd51322, 16'd29301});
	test_expansion(128'h0aae02cbb5b8561953d9bcff1a43445a, {16'd2089, 16'd27932, 16'd47398, 16'd4504, 16'd51116, 16'd60643, 16'd37352, 16'd20889, 16'd39484, 16'd39579, 16'd54713, 16'd20192, 16'd61143, 16'd49599, 16'd7071, 16'd3432, 16'd46612, 16'd27830, 16'd42190, 16'd16443, 16'd17272, 16'd29064, 16'd6984, 16'd17439, 16'd54840, 16'd18165});
	test_expansion(128'hae5c817fd1b0925caecb7a1ea3bbdf94, {16'd19561, 16'd50571, 16'd17172, 16'd29612, 16'd53205, 16'd58403, 16'd1273, 16'd10365, 16'd12679, 16'd18947, 16'd53207, 16'd23920, 16'd28136, 16'd39433, 16'd48477, 16'd664, 16'd4662, 16'd43818, 16'd34059, 16'd34876, 16'd38044, 16'd12372, 16'd34490, 16'd1119, 16'd24239, 16'd12849});
	test_expansion(128'ha1ac4e4828aa9b691e2d0339d7cf7284, {16'd12281, 16'd16665, 16'd10497, 16'd31010, 16'd7632, 16'd10010, 16'd28429, 16'd26540, 16'd20649, 16'd47001, 16'd22731, 16'd35297, 16'd39578, 16'd49824, 16'd45659, 16'd13157, 16'd60650, 16'd20520, 16'd8502, 16'd53924, 16'd64760, 16'd39893, 16'd9441, 16'd15897, 16'd40586, 16'd21005});
	test_expansion(128'hfe253f97ca19ca6083028efdcf05790a, {16'd24213, 16'd5874, 16'd60802, 16'd3385, 16'd56108, 16'd11650, 16'd56577, 16'd17073, 16'd25452, 16'd30299, 16'd26892, 16'd49415, 16'd5223, 16'd58866, 16'd20275, 16'd14867, 16'd21757, 16'd27649, 16'd14801, 16'd52988, 16'd14651, 16'd10912, 16'd4433, 16'd57754, 16'd61351, 16'd63890});
	test_expansion(128'hb245e58fe504d70bc8b8b02bc3c73383, {16'd27576, 16'd63451, 16'd28522, 16'd27845, 16'd24301, 16'd10746, 16'd36621, 16'd8210, 16'd64301, 16'd8058, 16'd53214, 16'd3994, 16'd64458, 16'd37535, 16'd63494, 16'd51689, 16'd45313, 16'd56334, 16'd60239, 16'd19956, 16'd57272, 16'd4243, 16'd61822, 16'd48164, 16'd5911, 16'd52092});
	test_expansion(128'h6b280e93eea1bced901fe75915b5359f, {16'd17661, 16'd22608, 16'd65226, 16'd61450, 16'd38117, 16'd44845, 16'd17053, 16'd9112, 16'd17855, 16'd7659, 16'd3271, 16'd53657, 16'd55907, 16'd3131, 16'd18258, 16'd37162, 16'd65050, 16'd37710, 16'd14724, 16'd54059, 16'd32863, 16'd57410, 16'd10492, 16'd18065, 16'd10309, 16'd3554});
	test_expansion(128'h3f6cde82615880ffbb9cd42719e3d02d, {16'd48368, 16'd19834, 16'd47881, 16'd27668, 16'd57032, 16'd9020, 16'd6984, 16'd10101, 16'd35564, 16'd16459, 16'd30864, 16'd51105, 16'd23339, 16'd33073, 16'd22909, 16'd60363, 16'd24216, 16'd2826, 16'd43350, 16'd36100, 16'd7117, 16'd53529, 16'd32043, 16'd45681, 16'd51887, 16'd40548});
	test_expansion(128'hea305f9b251055dd68b25ad6a981d616, {16'd16779, 16'd53787, 16'd27962, 16'd16811, 16'd61452, 16'd8954, 16'd58880, 16'd41802, 16'd27094, 16'd20030, 16'd18623, 16'd13732, 16'd31672, 16'd60583, 16'd921, 16'd14067, 16'd41178, 16'd23899, 16'd49291, 16'd26001, 16'd64896, 16'd810, 16'd1551, 16'd40562, 16'd18007, 16'd25749});
	test_expansion(128'hbc51c58addccfbe8b0ee36b6c9891b29, {16'd33765, 16'd2865, 16'd51084, 16'd15608, 16'd13606, 16'd61063, 16'd8770, 16'd8764, 16'd4729, 16'd46735, 16'd33894, 16'd47266, 16'd21470, 16'd33495, 16'd5700, 16'd33229, 16'd30429, 16'd33899, 16'd12041, 16'd44013, 16'd25956, 16'd14466, 16'd18656, 16'd60677, 16'd33693, 16'd12442});
	test_expansion(128'h1ea5a9cc78669cc36189815d4e3e157f, {16'd24345, 16'd64089, 16'd48838, 16'd64464, 16'd63571, 16'd26322, 16'd37841, 16'd2213, 16'd58349, 16'd46015, 16'd61256, 16'd39861, 16'd439, 16'd39971, 16'd15111, 16'd54593, 16'd49575, 16'd41971, 16'd46506, 16'd47039, 16'd34035, 16'd29257, 16'd36452, 16'd47597, 16'd49742, 16'd29598});
	test_expansion(128'h9a286ec4103eaae7a2af1b62222108cc, {16'd50567, 16'd6360, 16'd7457, 16'd48956, 16'd48855, 16'd53738, 16'd24278, 16'd20456, 16'd52113, 16'd26877, 16'd33390, 16'd63882, 16'd15861, 16'd47169, 16'd64422, 16'd52314, 16'd7676, 16'd33186, 16'd47591, 16'd22445, 16'd59605, 16'd4349, 16'd33848, 16'd1570, 16'd55587, 16'd25173});
	test_expansion(128'hb6cac1acd337808adbedc380708d27bc, {16'd10668, 16'd61291, 16'd60768, 16'd41653, 16'd49482, 16'd44920, 16'd8003, 16'd41686, 16'd18349, 16'd39903, 16'd5337, 16'd19748, 16'd3857, 16'd52301, 16'd35654, 16'd17102, 16'd51426, 16'd11270, 16'd42355, 16'd30648, 16'd2732, 16'd14713, 16'd4162, 16'd13610, 16'd28425, 16'd14216});
	test_expansion(128'h48765c3b3e043032ad87233238b8f111, {16'd16780, 16'd39883, 16'd62994, 16'd26371, 16'd3763, 16'd46270, 16'd14473, 16'd8188, 16'd56980, 16'd40968, 16'd49785, 16'd8054, 16'd14992, 16'd53741, 16'd28401, 16'd3130, 16'd5630, 16'd40136, 16'd48189, 16'd3231, 16'd59560, 16'd30732, 16'd54820, 16'd16499, 16'd60413, 16'd51320});
	test_expansion(128'haf8634bef6c8e9abd906ec34214b5457, {16'd15320, 16'd48932, 16'd25213, 16'd3729, 16'd36563, 16'd20638, 16'd4535, 16'd29642, 16'd35232, 16'd29453, 16'd254, 16'd46063, 16'd42167, 16'd37016, 16'd48093, 16'd46593, 16'd59463, 16'd35813, 16'd31209, 16'd37005, 16'd7223, 16'd64349, 16'd53546, 16'd52131, 16'd34755, 16'd64536});
	test_expansion(128'hed842f340fe87a55c259172781ef49fa, {16'd5098, 16'd27360, 16'd59650, 16'd51408, 16'd27979, 16'd60406, 16'd56355, 16'd36167, 16'd4021, 16'd11560, 16'd4149, 16'd6303, 16'd17947, 16'd31074, 16'd6446, 16'd30857, 16'd27545, 16'd24856, 16'd49568, 16'd60340, 16'd41099, 16'd22461, 16'd45719, 16'd19885, 16'd56013, 16'd14168});
	test_expansion(128'hd46ab6df59d8fae9f43dce2bf69fc40c, {16'd54296, 16'd38090, 16'd16450, 16'd9831, 16'd12446, 16'd20246, 16'd52551, 16'd43586, 16'd33079, 16'd13360, 16'd2030, 16'd52308, 16'd9158, 16'd1281, 16'd48345, 16'd6107, 16'd39906, 16'd4105, 16'd39589, 16'd5634, 16'd3328, 16'd34863, 16'd48873, 16'd29263, 16'd52414, 16'd56728});
	test_expansion(128'hbe1ad29872ed8d7e274123e262aff57d, {16'd26931, 16'd18993, 16'd30366, 16'd12994, 16'd31811, 16'd35994, 16'd16436, 16'd45696, 16'd6849, 16'd10409, 16'd46316, 16'd58454, 16'd29811, 16'd29973, 16'd65439, 16'd12076, 16'd18546, 16'd35832, 16'd23443, 16'd56062, 16'd25629, 16'd26518, 16'd25668, 16'd19716, 16'd4984, 16'd3652});
	test_expansion(128'hba97bf1b2ab9f84956373e72f65c4581, {16'd21157, 16'd59303, 16'd62182, 16'd51877, 16'd18742, 16'd1498, 16'd15004, 16'd51965, 16'd34983, 16'd8683, 16'd63386, 16'd58884, 16'd5117, 16'd21025, 16'd29345, 16'd1111, 16'd47375, 16'd64291, 16'd2192, 16'd43054, 16'd60809, 16'd31865, 16'd13006, 16'd39432, 16'd49107, 16'd55135});
	test_expansion(128'hede10eacd5cc3b509914a8f59cf6ee9e, {16'd13613, 16'd294, 16'd9660, 16'd24689, 16'd56909, 16'd58640, 16'd15143, 16'd33066, 16'd46600, 16'd48985, 16'd14466, 16'd11706, 16'd53494, 16'd18873, 16'd40554, 16'd17383, 16'd15837, 16'd38590, 16'd25445, 16'd19307, 16'd53907, 16'd28809, 16'd55178, 16'd49357, 16'd47670, 16'd5130});
	test_expansion(128'h4d08dfa4853373817576cca9cf0bc7ae, {16'd47990, 16'd54678, 16'd7488, 16'd30118, 16'd50987, 16'd58525, 16'd13834, 16'd3299, 16'd40502, 16'd46997, 16'd36318, 16'd43697, 16'd63787, 16'd57482, 16'd18074, 16'd43669, 16'd49802, 16'd25007, 16'd3372, 16'd52371, 16'd7924, 16'd40228, 16'd60789, 16'd24395, 16'd6855, 16'd4290});
	test_expansion(128'h4541983daa475dd18ccdcb6c55666619, {16'd15776, 16'd883, 16'd46708, 16'd34572, 16'd43950, 16'd27588, 16'd40596, 16'd63737, 16'd61115, 16'd19452, 16'd49128, 16'd60748, 16'd6935, 16'd7266, 16'd11586, 16'd33882, 16'd35560, 16'd44653, 16'd32428, 16'd15527, 16'd9578, 16'd60810, 16'd40179, 16'd19200, 16'd53418, 16'd22435});
	test_expansion(128'ha4b5af37cc69c24778dd255bac601159, {16'd53788, 16'd53074, 16'd62533, 16'd21668, 16'd56385, 16'd62805, 16'd35694, 16'd24513, 16'd25757, 16'd24957, 16'd35153, 16'd31344, 16'd18268, 16'd6171, 16'd61238, 16'd55576, 16'd1852, 16'd57606, 16'd58737, 16'd55841, 16'd18262, 16'd53304, 16'd28722, 16'd60536, 16'd56985, 16'd29396});
	test_expansion(128'h80226cfd4fa1b6798d02e58e2ef203b6, {16'd7321, 16'd44338, 16'd9374, 16'd43064, 16'd7059, 16'd17579, 16'd25398, 16'd49686, 16'd42506, 16'd14942, 16'd55209, 16'd9575, 16'd53869, 16'd49578, 16'd37507, 16'd51496, 16'd38954, 16'd5831, 16'd25569, 16'd38968, 16'd29912, 16'd24238, 16'd49985, 16'd28568, 16'd6093, 16'd49751});
	test_expansion(128'h4aa132226ad84f2a03fc9de9e4bf0969, {16'd43574, 16'd36135, 16'd5526, 16'd12012, 16'd20226, 16'd30542, 16'd12044, 16'd45350, 16'd63613, 16'd9279, 16'd19889, 16'd45046, 16'd58923, 16'd51439, 16'd10512, 16'd44456, 16'd7511, 16'd61608, 16'd27836, 16'd29879, 16'd21450, 16'd10185, 16'd8951, 16'd26160, 16'd57946, 16'd37047});
	test_expansion(128'h669b060136d70c07e030fa75e07c6484, {16'd41929, 16'd16833, 16'd25536, 16'd55436, 16'd45156, 16'd39601, 16'd31672, 16'd6026, 16'd6799, 16'd57769, 16'd1863, 16'd16662, 16'd48937, 16'd5696, 16'd22876, 16'd56172, 16'd64889, 16'd1724, 16'd26026, 16'd46337, 16'd13360, 16'd61941, 16'd28411, 16'd825, 16'd56362, 16'd45115});
	test_expansion(128'he2c2f7ba4af67775c79944bfa33b7357, {16'd30593, 16'd20090, 16'd16731, 16'd12729, 16'd4318, 16'd59192, 16'd22413, 16'd42399, 16'd43856, 16'd19980, 16'd55497, 16'd49092, 16'd52430, 16'd30435, 16'd44760, 16'd27087, 16'd63662, 16'd30989, 16'd35522, 16'd58545, 16'd13854, 16'd11774, 16'd16403, 16'd33685, 16'd33243, 16'd60174});
	test_expansion(128'h25c72691bdabf3838d789f6ef5280afe, {16'd45632, 16'd28538, 16'd22570, 16'd38425, 16'd49698, 16'd27586, 16'd50167, 16'd44121, 16'd6074, 16'd33788, 16'd15718, 16'd63443, 16'd4590, 16'd14246, 16'd24578, 16'd5093, 16'd24346, 16'd12551, 16'd10692, 16'd7966, 16'd57182, 16'd46770, 16'd14269, 16'd37032, 16'd35015, 16'd60733});
	test_expansion(128'h6ba83eb191d43ce65a76dfdc91e8ae5c, {16'd54261, 16'd43727, 16'd33326, 16'd24825, 16'd23273, 16'd15934, 16'd63351, 16'd50897, 16'd32629, 16'd11433, 16'd13902, 16'd41578, 16'd17127, 16'd39100, 16'd45451, 16'd49187, 16'd47929, 16'd50845, 16'd57551, 16'd63661, 16'd41683, 16'd9475, 16'd28954, 16'd11186, 16'd50424, 16'd18525});
	test_expansion(128'hb981087815ed93dbaf92eb3656657632, {16'd25590, 16'd59669, 16'd279, 16'd20263, 16'd2870, 16'd56336, 16'd32062, 16'd62275, 16'd58507, 16'd41520, 16'd20901, 16'd13864, 16'd44107, 16'd15731, 16'd42472, 16'd1803, 16'd8877, 16'd7394, 16'd61173, 16'd59061, 16'd10138, 16'd3158, 16'd56716, 16'd45969, 16'd7080, 16'd5003});
	test_expansion(128'h24d4a2567cc5acffbe2af6fda985b826, {16'd30360, 16'd7431, 16'd18698, 16'd24454, 16'd30283, 16'd7252, 16'd19089, 16'd25849, 16'd27019, 16'd39604, 16'd41705, 16'd678, 16'd51322, 16'd26460, 16'd62582, 16'd56719, 16'd38931, 16'd12612, 16'd4637, 16'd13139, 16'd24827, 16'd54509, 16'd2765, 16'd35142, 16'd25968, 16'd56694});
	test_expansion(128'h799e297b27518a58cae2141991113f35, {16'd27734, 16'd18313, 16'd34365, 16'd14909, 16'd30991, 16'd16046, 16'd11484, 16'd42450, 16'd28960, 16'd17082, 16'd17725, 16'd19072, 16'd27692, 16'd57847, 16'd26660, 16'd48933, 16'd46744, 16'd48898, 16'd32876, 16'd53150, 16'd33654, 16'd17690, 16'd25245, 16'd3927, 16'd2312, 16'd57862});
	test_expansion(128'hf48a084bb3bd6052672bf311ade3ae75, {16'd20081, 16'd28851, 16'd65166, 16'd46754, 16'd4542, 16'd29153, 16'd41168, 16'd26547, 16'd39116, 16'd23837, 16'd28549, 16'd21721, 16'd41875, 16'd55872, 16'd6546, 16'd30639, 16'd25571, 16'd26721, 16'd24503, 16'd2006, 16'd57090, 16'd50821, 16'd47811, 16'd22718, 16'd6693, 16'd41429});
	test_expansion(128'h5aa38fd30fc73352debc5d35f3e958e8, {16'd39936, 16'd8260, 16'd56238, 16'd58603, 16'd15345, 16'd49367, 16'd54889, 16'd51669, 16'd32032, 16'd29284, 16'd15749, 16'd51914, 16'd48239, 16'd55609, 16'd48253, 16'd15078, 16'd65312, 16'd45249, 16'd2384, 16'd63376, 16'd13426, 16'd27184, 16'd4472, 16'd52839, 16'd6656, 16'd29372});
	test_expansion(128'h3cc2b945889201d066d81f14baf56be7, {16'd57429, 16'd31775, 16'd25619, 16'd8294, 16'd25736, 16'd48386, 16'd18862, 16'd21385, 16'd28281, 16'd39101, 16'd55567, 16'd62146, 16'd12418, 16'd19758, 16'd11534, 16'd52674, 16'd2335, 16'd33273, 16'd914, 16'd53860, 16'd9001, 16'd2500, 16'd33494, 16'd1416, 16'd51753, 16'd3412});
	test_expansion(128'h624297ce7ee8f552a51049a468630be6, {16'd15800, 16'd26933, 16'd47280, 16'd22721, 16'd20330, 16'd18092, 16'd50019, 16'd14887, 16'd38841, 16'd47458, 16'd53079, 16'd23296, 16'd50838, 16'd31553, 16'd38564, 16'd28103, 16'd50081, 16'd58791, 16'd8282, 16'd47137, 16'd59302, 16'd56296, 16'd51351, 16'd15278, 16'd62868, 16'd12343});
	test_expansion(128'h1415ffad4a5a31f0b63c96471f5fda14, {16'd61857, 16'd49884, 16'd57732, 16'd34785, 16'd8374, 16'd44901, 16'd35309, 16'd51119, 16'd55701, 16'd25950, 16'd23234, 16'd40510, 16'd17842, 16'd29204, 16'd30757, 16'd50177, 16'd10303, 16'd21392, 16'd28921, 16'd63448, 16'd7429, 16'd38286, 16'd31042, 16'd4950, 16'd31283, 16'd37477});
	test_expansion(128'h7d2893eb8c2400e58f611bfe4188c296, {16'd31058, 16'd60942, 16'd61870, 16'd34421, 16'd39735, 16'd40448, 16'd64172, 16'd22843, 16'd41195, 16'd24135, 16'd59961, 16'd3266, 16'd15224, 16'd60722, 16'd844, 16'd5507, 16'd31935, 16'd30750, 16'd474, 16'd14049, 16'd43266, 16'd30306, 16'd45318, 16'd4944, 16'd53252, 16'd3917});
	test_expansion(128'hd5969f9e2d1f49b7afe533e372a9344c, {16'd64429, 16'd51533, 16'd36773, 16'd49669, 16'd11038, 16'd8946, 16'd15403, 16'd56520, 16'd33981, 16'd25785, 16'd59393, 16'd64336, 16'd33640, 16'd23207, 16'd23613, 16'd20303, 16'd42589, 16'd55726, 16'd49285, 16'd16192, 16'd33720, 16'd40531, 16'd45525, 16'd30880, 16'd16436, 16'd19934});
	test_expansion(128'hcffab165d7d83ec6d957d7245ebf2af5, {16'd41468, 16'd37919, 16'd25124, 16'd38314, 16'd44811, 16'd43496, 16'd56518, 16'd56297, 16'd12149, 16'd50544, 16'd8090, 16'd29065, 16'd62368, 16'd16140, 16'd23977, 16'd27576, 16'd49564, 16'd40984, 16'd59460, 16'd10444, 16'd24371, 16'd8294, 16'd758, 16'd5019, 16'd57848, 16'd41333});
	test_expansion(128'h3646d4aaa691651f57129b11052a5410, {16'd18788, 16'd65403, 16'd22663, 16'd46756, 16'd9336, 16'd58358, 16'd11688, 16'd46357, 16'd22601, 16'd53149, 16'd27526, 16'd37597, 16'd24537, 16'd7725, 16'd16018, 16'd29172, 16'd54279, 16'd8527, 16'd48369, 16'd59503, 16'd32904, 16'd6048, 16'd63618, 16'd4182, 16'd33523, 16'd15066});
	test_expansion(128'hf7a3e0bed09c7ea3bcdfe1ab85d688b3, {16'd2278, 16'd26789, 16'd35935, 16'd52353, 16'd21952, 16'd11130, 16'd41228, 16'd55619, 16'd10502, 16'd46657, 16'd48199, 16'd28678, 16'd56342, 16'd52641, 16'd32802, 16'd44048, 16'd26714, 16'd21227, 16'd26912, 16'd20402, 16'd40125, 16'd13951, 16'd23587, 16'd34140, 16'd41459, 16'd40307});
	test_expansion(128'h25bf2b236969c55b4f0538f9ec7cce91, {16'd22326, 16'd54376, 16'd18261, 16'd26091, 16'd43981, 16'd65410, 16'd50280, 16'd4396, 16'd49481, 16'd4759, 16'd4390, 16'd35379, 16'd24875, 16'd16760, 16'd55507, 16'd48560, 16'd9382, 16'd29, 16'd47179, 16'd55789, 16'd42659, 16'd53768, 16'd65402, 16'd11256, 16'd41447, 16'd14459});
	test_expansion(128'h33d8dc5b6c144caf96229ef3151a5f07, {16'd11710, 16'd55445, 16'd25324, 16'd33352, 16'd52854, 16'd1812, 16'd30846, 16'd34645, 16'd58311, 16'd22595, 16'd24490, 16'd62207, 16'd35504, 16'd20058, 16'd5969, 16'd24318, 16'd57903, 16'd6492, 16'd7976, 16'd23437, 16'd27383, 16'd17379, 16'd61573, 16'd10327, 16'd10856, 16'd38923});
	test_expansion(128'hb8778921fc581d467324be57cf41dafc, {16'd61728, 16'd46203, 16'd25082, 16'd43942, 16'd25142, 16'd38749, 16'd12561, 16'd11881, 16'd65196, 16'd51636, 16'd36675, 16'd46950, 16'd27833, 16'd56348, 16'd51432, 16'd36322, 16'd47673, 16'd37732, 16'd63436, 16'd10665, 16'd58322, 16'd14023, 16'd63096, 16'd12140, 16'd12646, 16'd41137});
	test_expansion(128'hb60f625d1b3c7f100fe7fb817d1f0382, {16'd42888, 16'd26212, 16'd7621, 16'd1067, 16'd59673, 16'd11950, 16'd50857, 16'd16299, 16'd53329, 16'd6141, 16'd56851, 16'd22310, 16'd27136, 16'd27584, 16'd23486, 16'd15440, 16'd63321, 16'd45937, 16'd38340, 16'd64962, 16'd53286, 16'd61166, 16'd5314, 16'd4585, 16'd41615, 16'd49882});
	test_expansion(128'h3719fe9a96bb59f6b89cd7c5981f046b, {16'd19507, 16'd65446, 16'd7651, 16'd2307, 16'd47565, 16'd33297, 16'd14099, 16'd43366, 16'd64393, 16'd6928, 16'd20042, 16'd33992, 16'd41102, 16'd8541, 16'd45072, 16'd1701, 16'd36244, 16'd37334, 16'd7312, 16'd26045, 16'd19166, 16'd37762, 16'd36571, 16'd55086, 16'd9958, 16'd22020});
	test_expansion(128'hb8d84b5a5019847a0acd984b401268d7, {16'd56639, 16'd31449, 16'd17196, 16'd54791, 16'd31827, 16'd49998, 16'd38420, 16'd64905, 16'd60946, 16'd13993, 16'd11336, 16'd33654, 16'd32606, 16'd30879, 16'd2333, 16'd4889, 16'd59675, 16'd46235, 16'd21023, 16'd56170, 16'd29668, 16'd30991, 16'd60416, 16'd7918, 16'd8164, 16'd57737});
	test_expansion(128'h82e15658358b7d056da8fe7ce66e2d7f, {16'd2925, 16'd29937, 16'd36562, 16'd35421, 16'd24562, 16'd34198, 16'd16363, 16'd51130, 16'd34785, 16'd48262, 16'd27810, 16'd17842, 16'd35492, 16'd22689, 16'd39910, 16'd17462, 16'd58127, 16'd38451, 16'd4119, 16'd23637, 16'd38164, 16'd2594, 16'd23538, 16'd58825, 16'd30326, 16'd4776});
	test_expansion(128'h5ec961c9598fc1819c05b981d48abbd4, {16'd18239, 16'd47787, 16'd57243, 16'd57322, 16'd723, 16'd21105, 16'd46430, 16'd43859, 16'd58231, 16'd15420, 16'd32889, 16'd23311, 16'd11349, 16'd60177, 16'd48696, 16'd48580, 16'd45154, 16'd40210, 16'd37074, 16'd7827, 16'd53976, 16'd26602, 16'd41448, 16'd52997, 16'd61872, 16'd24722});
	test_expansion(128'h13ec6e8738c779c208032c8eb97c22dd, {16'd4555, 16'd48768, 16'd33715, 16'd14983, 16'd2211, 16'd46801, 16'd5165, 16'd65448, 16'd57581, 16'd3459, 16'd7762, 16'd13655, 16'd13801, 16'd28167, 16'd11150, 16'd52347, 16'd46231, 16'd4149, 16'd36035, 16'd26137, 16'd63490, 16'd13923, 16'd22299, 16'd609, 16'd58234, 16'd5628});
	test_expansion(128'h2694b332d741959632db0330cbc296fe, {16'd11967, 16'd31570, 16'd13160, 16'd56776, 16'd36753, 16'd7211, 16'd47812, 16'd50509, 16'd52251, 16'd50313, 16'd18873, 16'd4988, 16'd36831, 16'd5915, 16'd45564, 16'd47724, 16'd16247, 16'd5874, 16'd7555, 16'd56696, 16'd48874, 16'd29214, 16'd22106, 16'd31022, 16'd56057, 16'd65150});
	test_expansion(128'h2dfa4c807fa3b4be26e3f57af978f635, {16'd8471, 16'd7167, 16'd28409, 16'd50456, 16'd4856, 16'd64309, 16'd45170, 16'd23026, 16'd22869, 16'd52763, 16'd62006, 16'd23051, 16'd29977, 16'd1159, 16'd34328, 16'd29578, 16'd20892, 16'd59837, 16'd32438, 16'd10956, 16'd53436, 16'd10362, 16'd50070, 16'd53852, 16'd27374, 16'd63926});
	test_expansion(128'h3c0641f180746aeaff520cf64ed7242d, {16'd49379, 16'd3459, 16'd30745, 16'd15955, 16'd55033, 16'd17776, 16'd5369, 16'd41859, 16'd17416, 16'd26747, 16'd24681, 16'd58786, 16'd10116, 16'd14119, 16'd53492, 16'd36633, 16'd63814, 16'd37571, 16'd57993, 16'd2189, 16'd51918, 16'd47308, 16'd44795, 16'd48609, 16'd3034, 16'd64990});
	test_expansion(128'h310b91938554e5f381465fb4ab3cd36d, {16'd59172, 16'd16758, 16'd11483, 16'd21822, 16'd11414, 16'd14903, 16'd23022, 16'd64858, 16'd41897, 16'd21047, 16'd65244, 16'd38906, 16'd16572, 16'd2015, 16'd11155, 16'd60765, 16'd14207, 16'd26253, 16'd30075, 16'd53864, 16'd12817, 16'd3603, 16'd11046, 16'd50341, 16'd35581, 16'd40034});
	test_expansion(128'hb55a66a53c862dfdf611ef635e1d67ef, {16'd19561, 16'd51252, 16'd53964, 16'd1827, 16'd42447, 16'd35574, 16'd12002, 16'd49807, 16'd58839, 16'd62751, 16'd3068, 16'd20040, 16'd63236, 16'd995, 16'd39208, 16'd40043, 16'd46308, 16'd29086, 16'd33624, 16'd58047, 16'd63906, 16'd15706, 16'd55539, 16'd29058, 16'd11147, 16'd61745});
	test_expansion(128'hc916781a53dcf722462dce9d55dfbbcf, {16'd62769, 16'd3221, 16'd11243, 16'd33298, 16'd17503, 16'd37374, 16'd27504, 16'd58269, 16'd34730, 16'd28142, 16'd56765, 16'd49839, 16'd4852, 16'd11551, 16'd35527, 16'd21545, 16'd51343, 16'd7710, 16'd49136, 16'd8052, 16'd43210, 16'd35418, 16'd26416, 16'd62304, 16'd22802, 16'd34984});
	test_expansion(128'hfd574e6ec57ea446c471a2cfcb223c96, {16'd31526, 16'd47382, 16'd30795, 16'd23517, 16'd21173, 16'd44809, 16'd48952, 16'd16287, 16'd56526, 16'd42262, 16'd1417, 16'd52851, 16'd7334, 16'd24634, 16'd63103, 16'd13347, 16'd10535, 16'd39594, 16'd34123, 16'd28868, 16'd47230, 16'd33518, 16'd23936, 16'd65369, 16'd6082, 16'd53402});
	test_expansion(128'hc1f8a99cb869947c75c2951784bb7475, {16'd43999, 16'd19259, 16'd34761, 16'd58772, 16'd16995, 16'd36159, 16'd28639, 16'd47933, 16'd52151, 16'd42704, 16'd46940, 16'd37560, 16'd18515, 16'd11739, 16'd17170, 16'd39941, 16'd49420, 16'd9893, 16'd15505, 16'd44421, 16'd18032, 16'd48439, 16'd60370, 16'd2405, 16'd7008, 16'd55555});
	test_expansion(128'hbb9b36533d39699c43ef90ef23c0c802, {16'd61121, 16'd50226, 16'd58717, 16'd4527, 16'd15007, 16'd31043, 16'd38215, 16'd13229, 16'd47516, 16'd48548, 16'd9648, 16'd45760, 16'd6782, 16'd55789, 16'd14624, 16'd63936, 16'd4576, 16'd64489, 16'd43073, 16'd32894, 16'd4604, 16'd16506, 16'd44004, 16'd33104, 16'd24822, 16'd6433});
	test_expansion(128'h867c5b1198e933eb267ad9a06c269cfa, {16'd60078, 16'd48234, 16'd30978, 16'd20916, 16'd46648, 16'd38293, 16'd4724, 16'd17199, 16'd52655, 16'd44714, 16'd8151, 16'd38208, 16'd25883, 16'd45346, 16'd16166, 16'd55230, 16'd40344, 16'd64254, 16'd27802, 16'd1144, 16'd5273, 16'd458, 16'd15605, 16'd39091, 16'd6613, 16'd64088});
	test_expansion(128'heca3d32b98d1ca1879c404228ca534b5, {16'd42147, 16'd29922, 16'd12219, 16'd49127, 16'd55843, 16'd4857, 16'd21074, 16'd56127, 16'd5360, 16'd64991, 16'd57758, 16'd24778, 16'd36642, 16'd47004, 16'd48889, 16'd20853, 16'd64089, 16'd64510, 16'd32732, 16'd11440, 16'd43865, 16'd59911, 16'd59794, 16'd40419, 16'd35798, 16'd63181});
	test_expansion(128'hae993befa94eba236df2f74fec177dd4, {16'd19166, 16'd45283, 16'd21688, 16'd37269, 16'd22536, 16'd35764, 16'd27158, 16'd36635, 16'd51030, 16'd61823, 16'd47317, 16'd12040, 16'd21191, 16'd42598, 16'd21550, 16'd54148, 16'd3996, 16'd44881, 16'd53611, 16'd47001, 16'd51927, 16'd12629, 16'd44785, 16'd38597, 16'd32118, 16'd5808});
	test_expansion(128'hf2abb4d03f779f128bbe1799d956e739, {16'd55849, 16'd38376, 16'd139, 16'd6932, 16'd19567, 16'd37511, 16'd906, 16'd10772, 16'd32122, 16'd40168, 16'd3644, 16'd61766, 16'd29823, 16'd14741, 16'd32671, 16'd64950, 16'd37045, 16'd8951, 16'd45747, 16'd35503, 16'd56672, 16'd62208, 16'd57854, 16'd31563, 16'd23643, 16'd2666});
	test_expansion(128'he05d57280510ad5c5ba16f8bde864888, {16'd19652, 16'd5876, 16'd36116, 16'd56395, 16'd40031, 16'd48784, 16'd17315, 16'd25102, 16'd5027, 16'd31286, 16'd12738, 16'd11523, 16'd1969, 16'd48232, 16'd42234, 16'd56668, 16'd58233, 16'd27661, 16'd26145, 16'd64897, 16'd63002, 16'd22668, 16'd39913, 16'd41191, 16'd2912, 16'd7088});
	test_expansion(128'hd0e541654585532abdb3541fbc024468, {16'd42314, 16'd37758, 16'd47359, 16'd33064, 16'd42274, 16'd7507, 16'd27587, 16'd49740, 16'd43068, 16'd59897, 16'd10790, 16'd58565, 16'd33311, 16'd41404, 16'd36411, 16'd51815, 16'd2187, 16'd63857, 16'd24912, 16'd61202, 16'd5814, 16'd3255, 16'd54089, 16'd27452, 16'd41601, 16'd62995});
	test_expansion(128'hcda3c0177518d65588fceb5dd593e4e3, {16'd2251, 16'd12128, 16'd59674, 16'd50701, 16'd59040, 16'd2063, 16'd55943, 16'd18127, 16'd46567, 16'd48778, 16'd13330, 16'd13043, 16'd38672, 16'd20840, 16'd29349, 16'd10094, 16'd10123, 16'd61284, 16'd30517, 16'd43216, 16'd43936, 16'd52297, 16'd32398, 16'd59405, 16'd55568, 16'd57387});
	test_expansion(128'hd7565986ffd0210c67fb9684c13ce05a, {16'd38707, 16'd20954, 16'd47629, 16'd18634, 16'd15379, 16'd4756, 16'd42103, 16'd4772, 16'd11877, 16'd39982, 16'd25853, 16'd27931, 16'd37889, 16'd20262, 16'd14669, 16'd43677, 16'd23604, 16'd52636, 16'd50997, 16'd33752, 16'd12267, 16'd52495, 16'd25670, 16'd35932, 16'd20604, 16'd638});
	test_expansion(128'hccffb5a6211a9727d30d65da1c68e1d9, {16'd5961, 16'd39356, 16'd12059, 16'd57832, 16'd58596, 16'd55504, 16'd13511, 16'd30850, 16'd1042, 16'd57045, 16'd50603, 16'd55407, 16'd31342, 16'd20197, 16'd21084, 16'd53854, 16'd13470, 16'd56867, 16'd22553, 16'd9723, 16'd3859, 16'd25546, 16'd58409, 16'd40852, 16'd58924, 16'd42272});
	test_expansion(128'h3578a8c47ee44fbdb94877ab090a070f, {16'd51557, 16'd29165, 16'd4086, 16'd24907, 16'd62028, 16'd37763, 16'd36737, 16'd48527, 16'd62640, 16'd37972, 16'd55937, 16'd1000, 16'd40365, 16'd19253, 16'd26503, 16'd42882, 16'd45426, 16'd42100, 16'd26292, 16'd41228, 16'd37183, 16'd8286, 16'd22178, 16'd59974, 16'd43958, 16'd34894});
	test_expansion(128'ha056cf96edcbd975f3e9654149652c56, {16'd29650, 16'd5220, 16'd45621, 16'd29847, 16'd13551, 16'd26788, 16'd10002, 16'd7429, 16'd29009, 16'd59389, 16'd24290, 16'd33827, 16'd1192, 16'd3653, 16'd25529, 16'd18028, 16'd12530, 16'd16982, 16'd36707, 16'd19692, 16'd35883, 16'd6932, 16'd54209, 16'd51960, 16'd16382, 16'd391});
	test_expansion(128'h671e61471ea270c8f3bd294825d376d2, {16'd16998, 16'd40466, 16'd15254, 16'd31640, 16'd60853, 16'd61337, 16'd31521, 16'd30022, 16'd11164, 16'd48933, 16'd50992, 16'd55951, 16'd34078, 16'd15127, 16'd30098, 16'd38801, 16'd6707, 16'd41874, 16'd32570, 16'd53068, 16'd28424, 16'd57056, 16'd87, 16'd42705, 16'd14059, 16'd42412});
	test_expansion(128'h2968312729f073d58a4936eecc61eb71, {16'd57121, 16'd2210, 16'd34014, 16'd54535, 16'd3566, 16'd18034, 16'd5487, 16'd6209, 16'd11318, 16'd18649, 16'd64942, 16'd12607, 16'd4608, 16'd26111, 16'd18623, 16'd64824, 16'd56622, 16'd24245, 16'd38553, 16'd22172, 16'd6977, 16'd40078, 16'd9400, 16'd14414, 16'd16276, 16'd31164});
	test_expansion(128'h465bef1bc9ed521294a14d8290b40951, {16'd11329, 16'd24270, 16'd14865, 16'd34121, 16'd21717, 16'd61576, 16'd31368, 16'd42215, 16'd46364, 16'd19955, 16'd44415, 16'd22456, 16'd953, 16'd6189, 16'd6752, 16'd28022, 16'd41634, 16'd63745, 16'd34426, 16'd60301, 16'd5136, 16'd40852, 16'd23884, 16'd63046, 16'd53720, 16'd14393});
	test_expansion(128'h46d41127c63224206da26f73ff189382, {16'd23300, 16'd24700, 16'd801, 16'd27800, 16'd34597, 16'd56286, 16'd4065, 16'd19857, 16'd39207, 16'd6850, 16'd50273, 16'd63254, 16'd23518, 16'd38461, 16'd61207, 16'd17837, 16'd3702, 16'd18965, 16'd36077, 16'd4856, 16'd1542, 16'd36376, 16'd1843, 16'd8411, 16'd7970, 16'd13566});
	test_expansion(128'h08b1f9d4a77b1cd2208c96f0e84219b8, {16'd31275, 16'd63102, 16'd6529, 16'd12112, 16'd35911, 16'd50150, 16'd43936, 16'd25529, 16'd59912, 16'd35042, 16'd19539, 16'd16342, 16'd40450, 16'd16577, 16'd26179, 16'd17500, 16'd34075, 16'd22607, 16'd63070, 16'd38789, 16'd29058, 16'd51295, 16'd44260, 16'd23353, 16'd52649, 16'd26906});
	test_expansion(128'h069c6e604e4f6521b572d5993737f457, {16'd14886, 16'd17753, 16'd45831, 16'd4534, 16'd57344, 16'd28886, 16'd28673, 16'd43305, 16'd63780, 16'd6836, 16'd3830, 16'd39369, 16'd47418, 16'd20474, 16'd36227, 16'd6170, 16'd62066, 16'd52308, 16'd17208, 16'd55517, 16'd13143, 16'd38701, 16'd53028, 16'd53986, 16'd22039, 16'd14620});
	test_expansion(128'h1ffffda8e5d1ea04c8fd8cd488f90034, {16'd20390, 16'd37982, 16'd44836, 16'd9997, 16'd57109, 16'd50332, 16'd22208, 16'd32710, 16'd55242, 16'd32576, 16'd2503, 16'd52227, 16'd47711, 16'd19928, 16'd49375, 16'd58907, 16'd25620, 16'd26454, 16'd30903, 16'd25697, 16'd37343, 16'd27146, 16'd44454, 16'd43347, 16'd16507, 16'd24912});
	test_expansion(128'h643ceb27fa2069c9858c1a850fe6262e, {16'd31364, 16'd29800, 16'd32055, 16'd9226, 16'd32103, 16'd10057, 16'd28651, 16'd60175, 16'd22974, 16'd1091, 16'd29178, 16'd5060, 16'd57176, 16'd50209, 16'd14599, 16'd39015, 16'd50262, 16'd28398, 16'd52490, 16'd13684, 16'd20137, 16'd46279, 16'd60616, 16'd54345, 16'd57351, 16'd19652});
	test_expansion(128'h9a50c6125fccd2d051a81e0aba22a9ef, {16'd42922, 16'd11076, 16'd31715, 16'd39429, 16'd33414, 16'd720, 16'd47252, 16'd4531, 16'd4838, 16'd53218, 16'd55971, 16'd25621, 16'd54169, 16'd596, 16'd3623, 16'd24976, 16'd2403, 16'd39979, 16'd41553, 16'd43912, 16'd55353, 16'd51471, 16'd63085, 16'd7503, 16'd23049, 16'd11054});
	test_expansion(128'hfdcb581b4a983742e089b9655f6f1daa, {16'd58120, 16'd20473, 16'd6383, 16'd52434, 16'd56435, 16'd30149, 16'd41049, 16'd14633, 16'd56378, 16'd48618, 16'd37164, 16'd58090, 16'd60565, 16'd25080, 16'd35233, 16'd8904, 16'd10563, 16'd40329, 16'd29997, 16'd41952, 16'd60960, 16'd122, 16'd57745, 16'd48721, 16'd43561, 16'd478});
	test_expansion(128'h5dd9914287f1cbc1b19924fc48db4838, {16'd42413, 16'd18535, 16'd41666, 16'd27676, 16'd40646, 16'd31480, 16'd33986, 16'd12118, 16'd11090, 16'd20732, 16'd48107, 16'd22126, 16'd35419, 16'd8026, 16'd58236, 16'd50888, 16'd58964, 16'd34045, 16'd3727, 16'd53452, 16'd13544, 16'd48068, 16'd23603, 16'd38595, 16'd53883, 16'd29119});
	test_expansion(128'h3f4801e4ee926af804367335e738ab03, {16'd56410, 16'd61162, 16'd61160, 16'd48115, 16'd4076, 16'd24477, 16'd29277, 16'd36363, 16'd56931, 16'd56510, 16'd1415, 16'd13861, 16'd26048, 16'd26929, 16'd59589, 16'd11664, 16'd26784, 16'd62163, 16'd1612, 16'd55436, 16'd58943, 16'd58040, 16'd25956, 16'd39527, 16'd54516, 16'd35781});
	test_expansion(128'h3faff8cf9863807d752033c0e4b29cbb, {16'd1699, 16'd51735, 16'd47969, 16'd3093, 16'd5131, 16'd59567, 16'd25803, 16'd3510, 16'd32296, 16'd51597, 16'd13590, 16'd50560, 16'd16773, 16'd17067, 16'd21376, 16'd50912, 16'd1361, 16'd22851, 16'd1509, 16'd2601, 16'd55143, 16'd31223, 16'd27548, 16'd45258, 16'd48041, 16'd11820});
	test_expansion(128'he90f691294588db85b4cccec828605ff, {16'd54879, 16'd24831, 16'd41596, 16'd64734, 16'd49881, 16'd13535, 16'd42380, 16'd24469, 16'd10955, 16'd53304, 16'd28383, 16'd50962, 16'd33416, 16'd38152, 16'd540, 16'd37166, 16'd19685, 16'd60195, 16'd27229, 16'd36304, 16'd62544, 16'd44790, 16'd16137, 16'd15750, 16'd64411, 16'd5530});
	test_expansion(128'h05b17054c0dd1af6a48a867a746f2f9c, {16'd55642, 16'd31344, 16'd52639, 16'd44875, 16'd26030, 16'd19919, 16'd2817, 16'd46256, 16'd47512, 16'd37717, 16'd43938, 16'd34581, 16'd60433, 16'd57222, 16'd43066, 16'd16470, 16'd44823, 16'd6978, 16'd11958, 16'd4945, 16'd28226, 16'd16561, 16'd18599, 16'd55423, 16'd48885, 16'd19563});
	test_expansion(128'h36bdab4c7ec61835242b916e789d01e2, {16'd28551, 16'd35579, 16'd56222, 16'd37832, 16'd46643, 16'd4498, 16'd57535, 16'd21498, 16'd23432, 16'd51581, 16'd37320, 16'd54203, 16'd63868, 16'd41272, 16'd48014, 16'd10677, 16'd7227, 16'd38470, 16'd12908, 16'd40496, 16'd17010, 16'd54656, 16'd64906, 16'd36917, 16'd31624, 16'd64987});
	test_expansion(128'h3926454de2f98fee7e33c279257dc5ad, {16'd6714, 16'd30353, 16'd19726, 16'd37236, 16'd9582, 16'd31566, 16'd2001, 16'd1894, 16'd38957, 16'd21993, 16'd53205, 16'd53854, 16'd44364, 16'd18085, 16'd8991, 16'd30690, 16'd22016, 16'd49718, 16'd11779, 16'd46862, 16'd26665, 16'd29876, 16'd58147, 16'd33222, 16'd52910, 16'd24616});
	test_expansion(128'h07cad447215a4003bc66b804df65812d, {16'd21420, 16'd10293, 16'd43296, 16'd50739, 16'd12867, 16'd14213, 16'd62833, 16'd26995, 16'd63494, 16'd16809, 16'd27880, 16'd41145, 16'd3276, 16'd5298, 16'd9710, 16'd11244, 16'd10726, 16'd28783, 16'd6023, 16'd35176, 16'd46042, 16'd60213, 16'd56300, 16'd58268, 16'd25497, 16'd15451});
	test_expansion(128'ha09b25bbd8b7203ce39e6b90692e607d, {16'd40397, 16'd55233, 16'd646, 16'd62894, 16'd28312, 16'd43692, 16'd26332, 16'd62439, 16'd10768, 16'd55483, 16'd5723, 16'd59847, 16'd48900, 16'd41023, 16'd39521, 16'd47776, 16'd63397, 16'd62431, 16'd48392, 16'd55932, 16'd5567, 16'd189, 16'd59504, 16'd389, 16'd52620, 16'd15407});
	test_expansion(128'hd927591f60af620d0f9ff9f232d3814c, {16'd4406, 16'd25734, 16'd63324, 16'd2218, 16'd32806, 16'd37044, 16'd8491, 16'd26133, 16'd27122, 16'd2239, 16'd40163, 16'd10323, 16'd62347, 16'd40670, 16'd57582, 16'd48965, 16'd25472, 16'd51439, 16'd37609, 16'd35855, 16'd49777, 16'd47232, 16'd16671, 16'd24214, 16'd7723, 16'd18425});
	test_expansion(128'h93eeab7e223f9b692c3d9d616ac9e007, {16'd32063, 16'd21967, 16'd27670, 16'd27831, 16'd46151, 16'd51112, 16'd55158, 16'd34720, 16'd27999, 16'd40925, 16'd49835, 16'd10003, 16'd37972, 16'd29657, 16'd61880, 16'd34628, 16'd39213, 16'd57596, 16'd6614, 16'd46139, 16'd30632, 16'd50708, 16'd62112, 16'd64040, 16'd34231, 16'd18121});
	test_expansion(128'h05aae9a2abd448f328fe7bedd6f3840f, {16'd24867, 16'd39563, 16'd45868, 16'd16649, 16'd37952, 16'd51442, 16'd63528, 16'd57187, 16'd28783, 16'd1171, 16'd24422, 16'd1649, 16'd35486, 16'd27875, 16'd29560, 16'd52974, 16'd20995, 16'd43993, 16'd45474, 16'd28283, 16'd10136, 16'd34571, 16'd30947, 16'd48157, 16'd63137, 16'd60461});
	test_expansion(128'h3044f632f194db68889c2280e0327587, {16'd53542, 16'd48871, 16'd31127, 16'd38243, 16'd11752, 16'd21405, 16'd40948, 16'd8430, 16'd32483, 16'd57252, 16'd42075, 16'd43388, 16'd34040, 16'd46735, 16'd56698, 16'd18687, 16'd54749, 16'd21774, 16'd16921, 16'd44695, 16'd53285, 16'd18437, 16'd64632, 16'd15367, 16'd61431, 16'd13895});
	test_expansion(128'hc6a1911128a288caed4dfeedd8bcdb41, {16'd2681, 16'd6276, 16'd60297, 16'd21111, 16'd52686, 16'd28776, 16'd39399, 16'd13047, 16'd65021, 16'd52540, 16'd24733, 16'd27000, 16'd35662, 16'd24054, 16'd3061, 16'd13977, 16'd10320, 16'd42731, 16'd33836, 16'd15599, 16'd18767, 16'd25083, 16'd40224, 16'd22959, 16'd56514, 16'd54733});
	test_expansion(128'hb57b5ca564806d861bd45ce589185f3b, {16'd515, 16'd11356, 16'd4195, 16'd56052, 16'd33559, 16'd13667, 16'd36370, 16'd14643, 16'd57491, 16'd58865, 16'd14721, 16'd10951, 16'd47037, 16'd28261, 16'd3255, 16'd64056, 16'd14182, 16'd11522, 16'd54553, 16'd40107, 16'd30645, 16'd22595, 16'd35209, 16'd10031, 16'd50483, 16'd3522});
	test_expansion(128'h795145d0d7cede339af0cde631b34b2e, {16'd61897, 16'd56109, 16'd62036, 16'd63772, 16'd50163, 16'd3687, 16'd61706, 16'd34812, 16'd40757, 16'd25161, 16'd6311, 16'd31101, 16'd30511, 16'd48841, 16'd61500, 16'd39735, 16'd54519, 16'd53075, 16'd32425, 16'd17750, 16'd20245, 16'd6797, 16'd4679, 16'd19374, 16'd5424, 16'd5844});
	test_expansion(128'h73577cd02f84a349785e1d4b07a8bf89, {16'd20006, 16'd24314, 16'd64018, 16'd47533, 16'd51360, 16'd25676, 16'd61860, 16'd15803, 16'd43806, 16'd31592, 16'd4814, 16'd18193, 16'd50785, 16'd14276, 16'd18828, 16'd35847, 16'd4258, 16'd10153, 16'd7317, 16'd63463, 16'd35069, 16'd21897, 16'd924, 16'd40401, 16'd12882, 16'd56328});
	test_expansion(128'h0c96a63205d505fd59a922747a2540a6, {16'd35473, 16'd34099, 16'd4744, 16'd9013, 16'd62641, 16'd5160, 16'd64189, 16'd38141, 16'd48758, 16'd42054, 16'd41554, 16'd38836, 16'd52585, 16'd15562, 16'd24927, 16'd8740, 16'd22141, 16'd5455, 16'd35529, 16'd47879, 16'd62511, 16'd38628, 16'd63610, 16'd1483, 16'd23318, 16'd26918});
	test_expansion(128'hf121cd4b377d078e9b4cce8b7ba13a89, {16'd35018, 16'd30957, 16'd40229, 16'd37094, 16'd36162, 16'd56445, 16'd15094, 16'd51033, 16'd55414, 16'd16651, 16'd936, 16'd36663, 16'd61320, 16'd30089, 16'd38961, 16'd5036, 16'd5128, 16'd28207, 16'd47729, 16'd4428, 16'd15622, 16'd63141, 16'd19788, 16'd63330, 16'd3869, 16'd40582});
	test_expansion(128'h0fda5532833fa36819fc6d609fb03661, {16'd17414, 16'd53009, 16'd45874, 16'd18375, 16'd62935, 16'd61027, 16'd640, 16'd27744, 16'd969, 16'd11677, 16'd57718, 16'd3468, 16'd3310, 16'd55187, 16'd37014, 16'd65255, 16'd36254, 16'd38120, 16'd1283, 16'd13879, 16'd57191, 16'd30821, 16'd8022, 16'd51869, 16'd8856, 16'd50455});
	test_expansion(128'hf7575217c5b8660ed46bfd8fff30f6af, {16'd40111, 16'd15382, 16'd33182, 16'd54714, 16'd50618, 16'd58834, 16'd27373, 16'd534, 16'd19818, 16'd29336, 16'd18567, 16'd19900, 16'd9264, 16'd28982, 16'd23595, 16'd9264, 16'd58576, 16'd57939, 16'd25927, 16'd14694, 16'd61580, 16'd9857, 16'd65513, 16'd38044, 16'd63548, 16'd47937});
	test_expansion(128'hefd5907b5ebbb103c034fd0a6e21889b, {16'd63265, 16'd38719, 16'd6898, 16'd17740, 16'd14034, 16'd38853, 16'd24564, 16'd29677, 16'd29826, 16'd61058, 16'd40933, 16'd31757, 16'd23947, 16'd8404, 16'd24550, 16'd43749, 16'd21836, 16'd7190, 16'd54834, 16'd30893, 16'd28213, 16'd57817, 16'd39405, 16'd58017, 16'd63614, 16'd32334});
	test_expansion(128'he6c5e09d9153424af44ba0bc28d4fd54, {16'd12, 16'd21797, 16'd51143, 16'd38907, 16'd29809, 16'd58010, 16'd6874, 16'd48557, 16'd39008, 16'd26303, 16'd36170, 16'd45453, 16'd45452, 16'd22499, 16'd23319, 16'd56307, 16'd41308, 16'd10762, 16'd43622, 16'd59396, 16'd11994, 16'd11, 16'd43012, 16'd34094, 16'd4609, 16'd40918});
	test_expansion(128'h455f27a09c82a995788b65b661f61e2b, {16'd63505, 16'd36459, 16'd36317, 16'd9835, 16'd51043, 16'd51525, 16'd39521, 16'd45247, 16'd13867, 16'd1523, 16'd60464, 16'd18518, 16'd32569, 16'd58047, 16'd24168, 16'd21290, 16'd37407, 16'd53127, 16'd50953, 16'd63208, 16'd29893, 16'd43767, 16'd22041, 16'd47867, 16'd45520, 16'd18517});
	test_expansion(128'h25c6479231ab4cba40e6a5cd2ef1fdce, {16'd50034, 16'd22553, 16'd24557, 16'd6873, 16'd54456, 16'd35144, 16'd28132, 16'd53903, 16'd65059, 16'd52102, 16'd23166, 16'd59909, 16'd57400, 16'd21113, 16'd52153, 16'd28554, 16'd51408, 16'd43750, 16'd57673, 16'd15444, 16'd59779, 16'd12055, 16'd51425, 16'd50878, 16'd48413, 16'd18215});
	test_expansion(128'hbe73bfd9194c77eedc2c9e4e5f91fcb0, {16'd36817, 16'd23707, 16'd23078, 16'd1448, 16'd23824, 16'd9973, 16'd17346, 16'd6448, 16'd8401, 16'd48076, 16'd63390, 16'd27638, 16'd13272, 16'd53822, 16'd33304, 16'd4818, 16'd22762, 16'd29283, 16'd18345, 16'd55932, 16'd56613, 16'd2952, 16'd24950, 16'd5857, 16'd40077, 16'd53772});
	test_expansion(128'h7f7c267a09f63d7c20e6803eafa9c39c, {16'd42683, 16'd16462, 16'd13586, 16'd33667, 16'd31504, 16'd6088, 16'd60884, 16'd41455, 16'd50802, 16'd12271, 16'd2750, 16'd7360, 16'd20665, 16'd32016, 16'd4508, 16'd19156, 16'd51641, 16'd60354, 16'd43909, 16'd10810, 16'd22646, 16'd63272, 16'd54687, 16'd2138, 16'd56617, 16'd30404});
	test_expansion(128'hd508e7c4784014a545075dec955ab8c9, {16'd57061, 16'd26090, 16'd20958, 16'd57075, 16'd7017, 16'd51986, 16'd51033, 16'd50549, 16'd33035, 16'd415, 16'd2338, 16'd28412, 16'd29252, 16'd50409, 16'd38005, 16'd590, 16'd55712, 16'd51795, 16'd59779, 16'd44623, 16'd46840, 16'd2204, 16'd13328, 16'd63128, 16'd30814, 16'd58586});
	test_expansion(128'he4032ca6ed839d64863e11369de7a465, {16'd31284, 16'd39048, 16'd17384, 16'd19279, 16'd30613, 16'd50129, 16'd35124, 16'd38420, 16'd56215, 16'd37642, 16'd36115, 16'd16862, 16'd43475, 16'd18036, 16'd64295, 16'd11828, 16'd45897, 16'd23213, 16'd30728, 16'd36269, 16'd61914, 16'd1672, 16'd24073, 16'd18125, 16'd13253, 16'd62889});
	test_expansion(128'h3c5e392f3f17752f5cf13f219a86e299, {16'd50320, 16'd37808, 16'd36240, 16'd33830, 16'd36239, 16'd2870, 16'd52790, 16'd24617, 16'd25935, 16'd11706, 16'd18216, 16'd37628, 16'd14174, 16'd11028, 16'd2613, 16'd64273, 16'd35497, 16'd33344, 16'd22455, 16'd26700, 16'd17105, 16'd23921, 16'd42937, 16'd49299, 16'd35048, 16'd6790});
	test_expansion(128'hf9d50ba86407005f9e2a3109ad3a7145, {16'd10479, 16'd34380, 16'd10247, 16'd4675, 16'd10357, 16'd23102, 16'd35168, 16'd24523, 16'd60107, 16'd41999, 16'd14852, 16'd1011, 16'd59111, 16'd44726, 16'd41062, 16'd14441, 16'd42875, 16'd17072, 16'd20490, 16'd1878, 16'd9904, 16'd3778, 16'd65145, 16'd347, 16'd10274, 16'd53796});
	test_expansion(128'hdb6b63195742a342ee6b5ea981160e71, {16'd48225, 16'd35956, 16'd46959, 16'd61896, 16'd44479, 16'd58135, 16'd41863, 16'd48210, 16'd11899, 16'd31087, 16'd62189, 16'd14861, 16'd38698, 16'd55703, 16'd27653, 16'd730, 16'd35471, 16'd620, 16'd20907, 16'd20109, 16'd40092, 16'd12746, 16'd10310, 16'd13786, 16'd26102, 16'd20199});
	test_expansion(128'h35e6d7a56e95fec8b6cadd15ba5ec375, {16'd47192, 16'd36921, 16'd33240, 16'd47551, 16'd40815, 16'd36182, 16'd27523, 16'd53399, 16'd40716, 16'd12793, 16'd22458, 16'd58922, 16'd56516, 16'd34960, 16'd59100, 16'd36631, 16'd44464, 16'd45823, 16'd23789, 16'd13954, 16'd62592, 16'd16759, 16'd15101, 16'd2065, 16'd12841, 16'd18344});
	test_expansion(128'h412086d1a7b182d07ce57db380b77834, {16'd28440, 16'd56824, 16'd27397, 16'd2664, 16'd38573, 16'd41375, 16'd13541, 16'd32254, 16'd55108, 16'd41144, 16'd25256, 16'd34961, 16'd43812, 16'd59690, 16'd29626, 16'd47475, 16'd35441, 16'd62683, 16'd16069, 16'd5932, 16'd24354, 16'd4788, 16'd3847, 16'd11405, 16'd12200, 16'd45591});
	test_expansion(128'hc60eabb88ea472046ea91ac5f0af292d, {16'd13986, 16'd25693, 16'd13626, 16'd36495, 16'd9689, 16'd43544, 16'd59831, 16'd21735, 16'd21070, 16'd64909, 16'd61202, 16'd7899, 16'd15772, 16'd16924, 16'd21845, 16'd15776, 16'd23417, 16'd64013, 16'd62263, 16'd60492, 16'd10756, 16'd23991, 16'd32972, 16'd6149, 16'd39266, 16'd5669});
	test_expansion(128'h6944dffbaba933e63457a528821e5b2d, {16'd43844, 16'd3458, 16'd39879, 16'd12339, 16'd55696, 16'd55368, 16'd24151, 16'd50341, 16'd43880, 16'd1452, 16'd30300, 16'd62104, 16'd7904, 16'd59643, 16'd44091, 16'd6369, 16'd23072, 16'd64299, 16'd31212, 16'd58332, 16'd15459, 16'd7380, 16'd62804, 16'd32198, 16'd60027, 16'd58530});
	test_expansion(128'hc888e92a2ac16c0e0c15abf31df9538b, {16'd37364, 16'd13946, 16'd32122, 16'd14818, 16'd57650, 16'd22298, 16'd9024, 16'd32132, 16'd38039, 16'd24612, 16'd36781, 16'd62188, 16'd51353, 16'd18700, 16'd51928, 16'd5456, 16'd9492, 16'd25752, 16'd22892, 16'd18451, 16'd52752, 16'd29230, 16'd62890, 16'd13764, 16'd26652, 16'd14535});
	test_expansion(128'h879f44de7e088e8f76007f76de9f752c, {16'd33117, 16'd58904, 16'd12552, 16'd2515, 16'd33073, 16'd13282, 16'd37487, 16'd51146, 16'd54888, 16'd48140, 16'd33262, 16'd30332, 16'd21505, 16'd35287, 16'd26146, 16'd56991, 16'd31753, 16'd38641, 16'd63737, 16'd34861, 16'd39179, 16'd14932, 16'd38892, 16'd16919, 16'd37308, 16'd24664});
	test_expansion(128'h3031b2d5796fafddb9abea822179bb6e, {16'd60261, 16'd42691, 16'd26700, 16'd26473, 16'd14706, 16'd62335, 16'd23978, 16'd56964, 16'd4202, 16'd46725, 16'd51579, 16'd1234, 16'd61892, 16'd5622, 16'd10137, 16'd19384, 16'd35825, 16'd60068, 16'd22393, 16'd37575, 16'd40285, 16'd42795, 16'd506, 16'd27095, 16'd49194, 16'd31236});
	test_expansion(128'h9334146c62469b77b54d100bd91de4e0, {16'd14516, 16'd20452, 16'd19739, 16'd16864, 16'd2367, 16'd35125, 16'd54224, 16'd42764, 16'd62432, 16'd46643, 16'd11850, 16'd4436, 16'd19994, 16'd49373, 16'd667, 16'd56084, 16'd61541, 16'd49494, 16'd12824, 16'd16874, 16'd32923, 16'd14338, 16'd36953, 16'd33998, 16'd36786, 16'd61540});
	test_expansion(128'h7aa16620b8c147de6b8797e7c0bf3169, {16'd20832, 16'd55478, 16'd52614, 16'd41496, 16'd47358, 16'd860, 16'd23514, 16'd6417, 16'd32319, 16'd12032, 16'd59130, 16'd29463, 16'd16019, 16'd37677, 16'd24267, 16'd11251, 16'd54481, 16'd9741, 16'd19211, 16'd9973, 16'd23772, 16'd62925, 16'd24393, 16'd24621, 16'd62351, 16'd48652});
	test_expansion(128'h02a7508194c319c0c793ac3b453e8c5e, {16'd4778, 16'd12061, 16'd33966, 16'd11544, 16'd41366, 16'd50938, 16'd21455, 16'd54340, 16'd11104, 16'd32032, 16'd6607, 16'd2402, 16'd5108, 16'd1373, 16'd37622, 16'd53618, 16'd13583, 16'd58789, 16'd21318, 16'd55248, 16'd37873, 16'd324, 16'd56209, 16'd59455, 16'd24993, 16'd42057});
	test_expansion(128'h5951de6f91fc5e14121d7a315c8149f8, {16'd28139, 16'd40988, 16'd8471, 16'd62405, 16'd34633, 16'd58250, 16'd13268, 16'd25218, 16'd5234, 16'd21600, 16'd24637, 16'd46490, 16'd24373, 16'd63156, 16'd15866, 16'd65197, 16'd64724, 16'd34290, 16'd50068, 16'd27774, 16'd62094, 16'd30557, 16'd7470, 16'd14464, 16'd29392, 16'd48091});
	test_expansion(128'h65b51779a8baa9049fd5403b253d773e, {16'd8012, 16'd8625, 16'd13896, 16'd40977, 16'd51064, 16'd19377, 16'd62636, 16'd53884, 16'd2773, 16'd65039, 16'd12162, 16'd15908, 16'd8026, 16'd5885, 16'd41763, 16'd25804, 16'd5776, 16'd32161, 16'd26771, 16'd2929, 16'd26258, 16'd8338, 16'd57100, 16'd63030, 16'd4374, 16'd2695});
	test_expansion(128'hcc4cbf6abc817aee57419de9d9439ffe, {16'd14914, 16'd37323, 16'd31670, 16'd63203, 16'd56547, 16'd57748, 16'd38888, 16'd10088, 16'd5410, 16'd35451, 16'd53927, 16'd31605, 16'd12823, 16'd26442, 16'd25923, 16'd15714, 16'd25478, 16'd58031, 16'd56376, 16'd40868, 16'd62295, 16'd42004, 16'd27686, 16'd48625, 16'd61596, 16'd41207});
	test_expansion(128'h035edd73ce1d582c92aae6106edc1a58, {16'd12181, 16'd9220, 16'd60577, 16'd20324, 16'd43834, 16'd49959, 16'd34842, 16'd55761, 16'd17186, 16'd14411, 16'd55355, 16'd50383, 16'd35326, 16'd24479, 16'd37087, 16'd44301, 16'd42904, 16'd12079, 16'd6994, 16'd18491, 16'd18255, 16'd42446, 16'd1306, 16'd50406, 16'd18222, 16'd36920});
	test_expansion(128'h360d89efb113d227ba7ae10375fcd046, {16'd13529, 16'd18415, 16'd55443, 16'd14359, 16'd42565, 16'd58529, 16'd60788, 16'd24061, 16'd6369, 16'd31501, 16'd15762, 16'd16072, 16'd1201, 16'd63514, 16'd16262, 16'd30808, 16'd15287, 16'd53033, 16'd22104, 16'd51218, 16'd14708, 16'd56194, 16'd24751, 16'd33985, 16'd19898, 16'd4231});
	test_expansion(128'h8e51b24c332a467283d0fcbdb8a588f8, {16'd56787, 16'd7436, 16'd432, 16'd37206, 16'd50005, 16'd43778, 16'd48120, 16'd47938, 16'd34709, 16'd46317, 16'd31827, 16'd53501, 16'd41718, 16'd35730, 16'd5972, 16'd59032, 16'd41240, 16'd62596, 16'd12428, 16'd39062, 16'd8497, 16'd37943, 16'd61183, 16'd53526, 16'd52765, 16'd52137});
	test_expansion(128'hd33f15e101f3176e6c1e685a102e987d, {16'd57183, 16'd63999, 16'd21056, 16'd6293, 16'd23911, 16'd50619, 16'd59063, 16'd65369, 16'd13869, 16'd23205, 16'd32770, 16'd15641, 16'd37453, 16'd33923, 16'd8546, 16'd25284, 16'd62233, 16'd41093, 16'd58091, 16'd37744, 16'd29748, 16'd24895, 16'd52775, 16'd61852, 16'd23079, 16'd60278});
	test_expansion(128'h8f6fece1508000a6ca9d1aa1195f65fe, {16'd48712, 16'd4927, 16'd61051, 16'd5815, 16'd5593, 16'd7527, 16'd48277, 16'd18735, 16'd7219, 16'd59037, 16'd51678, 16'd46556, 16'd43040, 16'd298, 16'd20263, 16'd23118, 16'd5879, 16'd37601, 16'd19367, 16'd10693, 16'd54494, 16'd59962, 16'd53701, 16'd19551, 16'd42857, 16'd46933});
	test_expansion(128'h80f6303c283232bc2bce3d19b616d8be, {16'd41815, 16'd4866, 16'd27405, 16'd63607, 16'd65534, 16'd1035, 16'd14499, 16'd47604, 16'd60276, 16'd45065, 16'd14728, 16'd29740, 16'd59630, 16'd47867, 16'd19699, 16'd34702, 16'd2209, 16'd28267, 16'd64352, 16'd32859, 16'd49136, 16'd16761, 16'd58826, 16'd34907, 16'd57172, 16'd5093});
	test_expansion(128'h0526566da75d834df314f999aac6a23b, {16'd1395, 16'd5895, 16'd49607, 16'd49838, 16'd27536, 16'd43923, 16'd25628, 16'd48482, 16'd47255, 16'd36320, 16'd1615, 16'd47963, 16'd26029, 16'd24929, 16'd46571, 16'd29138, 16'd63838, 16'd15198, 16'd28946, 16'd20462, 16'd8288, 16'd16436, 16'd14842, 16'd24436, 16'd11133, 16'd54591});
	test_expansion(128'hdfff3ee01e59106153d6084b2b29e0f4, {16'd32779, 16'd28570, 16'd43549, 16'd34787, 16'd63091, 16'd54801, 16'd48531, 16'd44566, 16'd34104, 16'd6245, 16'd26832, 16'd29737, 16'd9038, 16'd63410, 16'd53527, 16'd3357, 16'd56082, 16'd47969, 16'd51700, 16'd35795, 16'd52496, 16'd43018, 16'd51987, 16'd14530, 16'd6316, 16'd7491});
	test_expansion(128'h49b5a2017bb6d8a6a8ee2f762f743933, {16'd32507, 16'd43934, 16'd52708, 16'd27018, 16'd43046, 16'd30776, 16'd57965, 16'd28373, 16'd41186, 16'd37922, 16'd61920, 16'd29451, 16'd17273, 16'd64600, 16'd23947, 16'd3750, 16'd61319, 16'd23077, 16'd21743, 16'd37972, 16'd25387, 16'd36313, 16'd49876, 16'd47481, 16'd28653, 16'd54733});
	test_expansion(128'hc6530dce63fa047da6154fcb728d32e3, {16'd32444, 16'd55489, 16'd16848, 16'd54317, 16'd55560, 16'd29016, 16'd64504, 16'd42112, 16'd60608, 16'd14923, 16'd43187, 16'd57658, 16'd3605, 16'd54743, 16'd22920, 16'd32185, 16'd44949, 16'd13679, 16'd9034, 16'd43589, 16'd50163, 16'd44464, 16'd10865, 16'd8700, 16'd24890, 16'd5716});
	test_expansion(128'h43d9a29d0e824e04db30951de2ed7925, {16'd39230, 16'd22768, 16'd45483, 16'd47863, 16'd50799, 16'd53393, 16'd56716, 16'd41894, 16'd16557, 16'd54410, 16'd18582, 16'd25663, 16'd50020, 16'd26487, 16'd21428, 16'd19948, 16'd4145, 16'd32003, 16'd39997, 16'd25523, 16'd14711, 16'd43452, 16'd46435, 16'd47814, 16'd17445, 16'd11561});
	test_expansion(128'h48eaa8a3a7cedeef96576f2c2fa4adcf, {16'd4512, 16'd31108, 16'd6345, 16'd17000, 16'd36297, 16'd924, 16'd29295, 16'd49928, 16'd24093, 16'd41313, 16'd31588, 16'd31458, 16'd34275, 16'd12443, 16'd4207, 16'd8384, 16'd62854, 16'd39742, 16'd34585, 16'd19421, 16'd58697, 16'd3529, 16'd35701, 16'd2020, 16'd30101, 16'd3786});
	test_expansion(128'h7c7a52a58a4341d997a9a5081593dd53, {16'd16138, 16'd35612, 16'd33213, 16'd24067, 16'd63582, 16'd64504, 16'd31361, 16'd36493, 16'd3532, 16'd31243, 16'd58894, 16'd21240, 16'd4553, 16'd65219, 16'd42059, 16'd5785, 16'd61142, 16'd9139, 16'd32696, 16'd7377, 16'd10611, 16'd5277, 16'd2933, 16'd43578, 16'd36982, 16'd3642});
	test_expansion(128'ha520d59df5427d851e6e1f329906e958, {16'd54956, 16'd48551, 16'd37224, 16'd5043, 16'd14503, 16'd31065, 16'd37620, 16'd49122, 16'd50212, 16'd18256, 16'd28213, 16'd40392, 16'd43870, 16'd52852, 16'd20631, 16'd8781, 16'd41277, 16'd39950, 16'd56221, 16'd36758, 16'd27618, 16'd48471, 16'd61064, 16'd26061, 16'd9481, 16'd17760});
	test_expansion(128'hfd7e736f352d85eb1b1dcc29ecdb1f0d, {16'd51562, 16'd27913, 16'd26449, 16'd45894, 16'd41195, 16'd36803, 16'd15601, 16'd59093, 16'd60407, 16'd30044, 16'd24113, 16'd16499, 16'd45245, 16'd22436, 16'd53750, 16'd4497, 16'd48883, 16'd20093, 16'd54226, 16'd36813, 16'd63583, 16'd16780, 16'd58968, 16'd39446, 16'd36751, 16'd36231});
	test_expansion(128'hbc5c96ec8ce3f348f063ef75daed0ba3, {16'd17255, 16'd7832, 16'd26415, 16'd14717, 16'd47098, 16'd21822, 16'd42133, 16'd61508, 16'd23291, 16'd54560, 16'd19227, 16'd8984, 16'd6712, 16'd61138, 16'd41838, 16'd26435, 16'd38493, 16'd61561, 16'd19855, 16'd54324, 16'd7943, 16'd38336, 16'd47180, 16'd13831, 16'd25947, 16'd143});
	test_expansion(128'h05ddd34168c68e65a00d5090587715be, {16'd24408, 16'd16570, 16'd41266, 16'd32767, 16'd7141, 16'd45073, 16'd9816, 16'd17463, 16'd64642, 16'd1948, 16'd32420, 16'd14026, 16'd19853, 16'd12817, 16'd26141, 16'd36744, 16'd60826, 16'd63922, 16'd11054, 16'd20947, 16'd47116, 16'd34493, 16'd14832, 16'd41219, 16'd24077, 16'd61920});
	test_expansion(128'h12aca32cafa78a624b483a41cb4d09e1, {16'd35013, 16'd56675, 16'd50682, 16'd57034, 16'd8560, 16'd62824, 16'd42129, 16'd35945, 16'd48559, 16'd62837, 16'd13237, 16'd42407, 16'd53237, 16'd139, 16'd29864, 16'd39576, 16'd8917, 16'd29200, 16'd49199, 16'd8513, 16'd12131, 16'd15620, 16'd40172, 16'd41872, 16'd11397, 16'd18667});
	test_expansion(128'hf015ddfeec39fedaf17f7f17034caf90, {16'd49013, 16'd56445, 16'd41139, 16'd9038, 16'd47369, 16'd4539, 16'd2542, 16'd5817, 16'd37212, 16'd573, 16'd56777, 16'd48321, 16'd57984, 16'd1399, 16'd31780, 16'd60453, 16'd60244, 16'd47001, 16'd41507, 16'd10159, 16'd20434, 16'd21342, 16'd36244, 16'd26599, 16'd49575, 16'd47076});
	test_expansion(128'h15fa05c0548925199daeea57c4490a8d, {16'd60139, 16'd37725, 16'd4558, 16'd51657, 16'd23915, 16'd34279, 16'd31861, 16'd41713, 16'd50334, 16'd56854, 16'd49140, 16'd46556, 16'd13289, 16'd44383, 16'd60113, 16'd37587, 16'd64218, 16'd20786, 16'd20755, 16'd64495, 16'd13387, 16'd44212, 16'd37448, 16'd10517, 16'd48638, 16'd28335});
	test_expansion(128'h9268e4ae3867ddc2a305b8301712c481, {16'd62799, 16'd40427, 16'd35731, 16'd27378, 16'd27158, 16'd33165, 16'd51373, 16'd31534, 16'd6151, 16'd59337, 16'd39879, 16'd62080, 16'd4221, 16'd17610, 16'd51013, 16'd18808, 16'd63032, 16'd30892, 16'd25280, 16'd36754, 16'd25869, 16'd35047, 16'd28618, 16'd46561, 16'd62763, 16'd18694});
	test_expansion(128'h67cdf2dff1a3d20d6b07d2a535da6c11, {16'd47533, 16'd20401, 16'd22419, 16'd97, 16'd34461, 16'd20391, 16'd55952, 16'd48698, 16'd17564, 16'd62781, 16'd41681, 16'd38450, 16'd55756, 16'd8142, 16'd21375, 16'd11537, 16'd6081, 16'd12649, 16'd45493, 16'd11736, 16'd23869, 16'd27702, 16'd34548, 16'd60006, 16'd35175, 16'd8484});
	test_expansion(128'hbc0cfe388eea38d050af366fb89a2463, {16'd63242, 16'd21767, 16'd58412, 16'd53748, 16'd17450, 16'd63470, 16'd38874, 16'd62587, 16'd17283, 16'd36963, 16'd8485, 16'd47420, 16'd2614, 16'd55524, 16'd56696, 16'd59266, 16'd21154, 16'd53327, 16'd27573, 16'd29873, 16'd52376, 16'd7134, 16'd22586, 16'd30726, 16'd46542, 16'd39591});
	test_expansion(128'hbab5c07553b058840291c39a6d824a12, {16'd32476, 16'd60791, 16'd19537, 16'd11271, 16'd54501, 16'd35951, 16'd5158, 16'd57443, 16'd61719, 16'd25557, 16'd30274, 16'd3591, 16'd44927, 16'd4635, 16'd12821, 16'd53854, 16'd57711, 16'd51507, 16'd30413, 16'd38530, 16'd48007, 16'd46023, 16'd58885, 16'd38807, 16'd38029, 16'd9020});
	test_expansion(128'h3a42154698fc2db5dc710edacaa5fa79, {16'd9010, 16'd29812, 16'd52475, 16'd65248, 16'd58634, 16'd63299, 16'd22373, 16'd16326, 16'd35846, 16'd30187, 16'd61071, 16'd26532, 16'd55662, 16'd42630, 16'd38151, 16'd50927, 16'd5910, 16'd43214, 16'd47614, 16'd23172, 16'd3826, 16'd20639, 16'd20630, 16'd16055, 16'd18932, 16'd12306});
	test_expansion(128'h1690c2478ec5a3f4cf5f5dcfa3f1713e, {16'd58201, 16'd573, 16'd8837, 16'd7292, 16'd18177, 16'd39532, 16'd26530, 16'd58742, 16'd58020, 16'd20851, 16'd13132, 16'd37348, 16'd38009, 16'd12963, 16'd33913, 16'd43963, 16'd35475, 16'd42747, 16'd10101, 16'd46169, 16'd54059, 16'd23936, 16'd23777, 16'd25583, 16'd42366, 16'd28571});
	test_expansion(128'h7359ce5334413f89b087690c8aafe874, {16'd4928, 16'd11574, 16'd7480, 16'd11569, 16'd53573, 16'd56997, 16'd5788, 16'd31152, 16'd15680, 16'd40483, 16'd12935, 16'd61511, 16'd51858, 16'd35063, 16'd60031, 16'd42646, 16'd14669, 16'd39055, 16'd43582, 16'd43081, 16'd3537, 16'd55714, 16'd33669, 16'd6570, 16'd2860, 16'd36467});
	test_expansion(128'h24a4480131b73c05deb140466583ab3a, {16'd42728, 16'd45359, 16'd24506, 16'd44554, 16'd58744, 16'd15851, 16'd2165, 16'd14648, 16'd9925, 16'd33923, 16'd58292, 16'd23998, 16'd62464, 16'd42102, 16'd41441, 16'd21424, 16'd8240, 16'd57649, 16'd42612, 16'd46904, 16'd15566, 16'd33227, 16'd28613, 16'd12162, 16'd9119, 16'd60219});
	test_expansion(128'h7b6fda327236c0e2ea098e401396cdda, {16'd232, 16'd38232, 16'd38230, 16'd9759, 16'd11681, 16'd34441, 16'd15940, 16'd14041, 16'd17634, 16'd24701, 16'd27944, 16'd37772, 16'd914, 16'd39768, 16'd40662, 16'd48899, 16'd33419, 16'd18362, 16'd10705, 16'd9139, 16'd24691, 16'd28244, 16'd1031, 16'd34558, 16'd9504, 16'd5540});
	test_expansion(128'h009e8339c7dee695525cdb7a1e36ed4b, {16'd53502, 16'd50674, 16'd24637, 16'd32376, 16'd41571, 16'd53883, 16'd1218, 16'd18630, 16'd2413, 16'd25926, 16'd50155, 16'd34498, 16'd58161, 16'd4032, 16'd35822, 16'd25320, 16'd43383, 16'd26286, 16'd54567, 16'd35061, 16'd40175, 16'd1462, 16'd2944, 16'd39390, 16'd49156, 16'd35384});
	test_expansion(128'hdca8dcb0742c9b26436ac7470ee8eb01, {16'd29454, 16'd37795, 16'd2162, 16'd8843, 16'd3900, 16'd21903, 16'd10261, 16'd22816, 16'd33766, 16'd63241, 16'd52464, 16'd30804, 16'd57014, 16'd34526, 16'd17009, 16'd37080, 16'd641, 16'd47227, 16'd46757, 16'd30088, 16'd39029, 16'd36700, 16'd51683, 16'd62083, 16'd61170, 16'd58381});
	test_expansion(128'hcb8ec482ca3de53b2b69b946964e484c, {16'd36412, 16'd46162, 16'd32698, 16'd55977, 16'd59259, 16'd56606, 16'd56107, 16'd28202, 16'd36238, 16'd6789, 16'd39632, 16'd54424, 16'd20546, 16'd23138, 16'd54195, 16'd41435, 16'd11807, 16'd47201, 16'd51052, 16'd30067, 16'd30838, 16'd24163, 16'd13201, 16'd31450, 16'd9666, 16'd62579});
	test_expansion(128'hf939371deb55602a64b94f126f9c8d8a, {16'd11739, 16'd32821, 16'd36497, 16'd2279, 16'd33892, 16'd41846, 16'd47506, 16'd23564, 16'd63247, 16'd10078, 16'd60084, 16'd32553, 16'd38095, 16'd24831, 16'd46505, 16'd33060, 16'd21898, 16'd57408, 16'd50680, 16'd44102, 16'd23051, 16'd12710, 16'd21716, 16'd7658, 16'd16926, 16'd51579});
	test_expansion(128'hf8770b4e960516f166649b1abb7f09a3, {16'd29690, 16'd42975, 16'd6512, 16'd64332, 16'd32795, 16'd43006, 16'd57579, 16'd4940, 16'd56723, 16'd9658, 16'd29481, 16'd1176, 16'd4712, 16'd46273, 16'd22915, 16'd35442, 16'd16716, 16'd13542, 16'd54251, 16'd59265, 16'd25597, 16'd19312, 16'd18594, 16'd27247, 16'd61486, 16'd54475});
	test_expansion(128'h0762be53b1178a2cbbba12e6858970f2, {16'd5448, 16'd56388, 16'd40208, 16'd14393, 16'd10067, 16'd2332, 16'd43236, 16'd6133, 16'd27195, 16'd33683, 16'd50743, 16'd38725, 16'd31178, 16'd10061, 16'd52562, 16'd54594, 16'd7098, 16'd3818, 16'd3432, 16'd16766, 16'd49094, 16'd4698, 16'd52613, 16'd22174, 16'd18499, 16'd51046});
	test_expansion(128'h672a3ed7c53b3c28021bca18915a98e8, {16'd17579, 16'd33930, 16'd17564, 16'd21687, 16'd60894, 16'd44242, 16'd22359, 16'd30580, 16'd62922, 16'd46421, 16'd40601, 16'd18212, 16'd43062, 16'd45020, 16'd49765, 16'd13007, 16'd59607, 16'd63163, 16'd57457, 16'd1357, 16'd5720, 16'd30068, 16'd41052, 16'd9376, 16'd6632, 16'd56224});
	test_expansion(128'h9553d72559d3f5cfa8ac6bd12a428fd5, {16'd30312, 16'd30410, 16'd14117, 16'd29694, 16'd55303, 16'd19969, 16'd62415, 16'd44306, 16'd34002, 16'd7396, 16'd62985, 16'd43247, 16'd64468, 16'd3599, 16'd29333, 16'd43359, 16'd26545, 16'd1496, 16'd3581, 16'd38013, 16'd50109, 16'd15022, 16'd50121, 16'd10051, 16'd41463, 16'd63941});
	test_expansion(128'h7f64b890a007eec3c22472163f4f9970, {16'd29511, 16'd25264, 16'd28140, 16'd10083, 16'd37753, 16'd59180, 16'd54265, 16'd17541, 16'd48903, 16'd19633, 16'd35116, 16'd49436, 16'd63851, 16'd2842, 16'd12415, 16'd37096, 16'd33953, 16'd44449, 16'd43434, 16'd39231, 16'd20531, 16'd7874, 16'd8484, 16'd17109, 16'd6382, 16'd8550});
	test_expansion(128'h92b694724c88f9123f2d4a9aa5900e5e, {16'd3379, 16'd15399, 16'd6462, 16'd7105, 16'd42468, 16'd12066, 16'd11072, 16'd37991, 16'd34656, 16'd19541, 16'd15820, 16'd50138, 16'd39510, 16'd38358, 16'd35183, 16'd34985, 16'd53346, 16'd25882, 16'd62246, 16'd19576, 16'd42850, 16'd37975, 16'd45369, 16'd47066, 16'd3475, 16'd51809});
	test_expansion(128'h7e6de95fe61d83fbe8adea8d876e5d1c, {16'd29911, 16'd40040, 16'd8319, 16'd14470, 16'd970, 16'd20945, 16'd46708, 16'd56129, 16'd58301, 16'd3583, 16'd52717, 16'd47534, 16'd11084, 16'd43918, 16'd55141, 16'd60487, 16'd18718, 16'd24022, 16'd44857, 16'd32808, 16'd54427, 16'd56900, 16'd63883, 16'd50193, 16'd22096, 16'd5876});
	test_expansion(128'h09cb2f80cb6b9b89d2f532da97148063, {16'd41076, 16'd60804, 16'd53071, 16'd15742, 16'd24928, 16'd46493, 16'd63102, 16'd22801, 16'd6486, 16'd32546, 16'd15801, 16'd25193, 16'd30454, 16'd37824, 16'd23508, 16'd35820, 16'd9163, 16'd34011, 16'd34320, 16'd44652, 16'd46364, 16'd59407, 16'd40055, 16'd35734, 16'd39927, 16'd16670});
	test_expansion(128'h152c19809693b5fcbc9704238b65719c, {16'd47368, 16'd65424, 16'd18288, 16'd54937, 16'd33708, 16'd3262, 16'd35562, 16'd32197, 16'd27381, 16'd63609, 16'd54241, 16'd13362, 16'd53649, 16'd38722, 16'd52578, 16'd449, 16'd36530, 16'd12883, 16'd9900, 16'd43518, 16'd19214, 16'd64035, 16'd62339, 16'd35628, 16'd62219, 16'd55030});
	test_expansion(128'h44407243f73615beee35f90c6e8d2efb, {16'd60449, 16'd9058, 16'd1884, 16'd26889, 16'd7777, 16'd34717, 16'd65071, 16'd23990, 16'd45636, 16'd973, 16'd50486, 16'd33929, 16'd56778, 16'd53959, 16'd48469, 16'd22343, 16'd55929, 16'd31649, 16'd19047, 16'd38732, 16'd31531, 16'd6225, 16'd39323, 16'd27713, 16'd23538, 16'd12811});
	test_expansion(128'h61e956bfdf135bb4d218192ff4361cf1, {16'd13999, 16'd63409, 16'd12531, 16'd6484, 16'd49803, 16'd43066, 16'd12458, 16'd27931, 16'd61965, 16'd64256, 16'd48180, 16'd27184, 16'd36866, 16'd43259, 16'd65522, 16'd45088, 16'd21905, 16'd16212, 16'd27561, 16'd37239, 16'd30856, 16'd52967, 16'd48488, 16'd45569, 16'd8206, 16'd47354});
	test_expansion(128'h4a2f1cb87da12de60d01c0d4b01e29d9, {16'd58062, 16'd16931, 16'd2198, 16'd6985, 16'd39827, 16'd4462, 16'd10065, 16'd37526, 16'd1673, 16'd8978, 16'd5081, 16'd65524, 16'd412, 16'd38708, 16'd7637, 16'd55900, 16'd13557, 16'd52687, 16'd41270, 16'd28859, 16'd9029, 16'd53196, 16'd49805, 16'd8591, 16'd53590, 16'd5599});
	test_expansion(128'ha00a232edab3728e1f53a55cf3085e66, {16'd20158, 16'd8184, 16'd30633, 16'd36196, 16'd41398, 16'd16062, 16'd40894, 16'd3894, 16'd11871, 16'd38528, 16'd26085, 16'd57072, 16'd31130, 16'd37470, 16'd54017, 16'd42814, 16'd50888, 16'd58694, 16'd26100, 16'd35763, 16'd28300, 16'd59534, 16'd46963, 16'd3964, 16'd54896, 16'd51129});
	test_expansion(128'h80c68ff4af2d2777e3e30ba5f7a49e60, {16'd46457, 16'd64717, 16'd10390, 16'd50480, 16'd47915, 16'd14723, 16'd7277, 16'd57724, 16'd14849, 16'd8644, 16'd10266, 16'd16108, 16'd19125, 16'd25797, 16'd25284, 16'd61981, 16'd13920, 16'd40237, 16'd38269, 16'd1888, 16'd826, 16'd47117, 16'd15231, 16'd65123, 16'd52164, 16'd12703});
	test_expansion(128'hb6998ba3f40ff1dd666a6e21a03b027e, {16'd14763, 16'd60653, 16'd15613, 16'd1971, 16'd26608, 16'd9654, 16'd52368, 16'd26172, 16'd1352, 16'd65284, 16'd58297, 16'd56074, 16'd57574, 16'd8967, 16'd35009, 16'd35642, 16'd32150, 16'd61111, 16'd37790, 16'd62235, 16'd686, 16'd54555, 16'd27619, 16'd13165, 16'd1552, 16'd41979});
	test_expansion(128'h366d7f5fb0edca31ccaf82b75d9e35c8, {16'd49316, 16'd50036, 16'd42124, 16'd9122, 16'd3841, 16'd30203, 16'd42379, 16'd37118, 16'd49809, 16'd27684, 16'd14038, 16'd43308, 16'd60014, 16'd26573, 16'd33001, 16'd34990, 16'd60170, 16'd11793, 16'd37313, 16'd49361, 16'd7151, 16'd21577, 16'd50596, 16'd41039, 16'd51896, 16'd39547});
	test_expansion(128'hf4ffc857943111e64d0b8fe893e1b98b, {16'd51189, 16'd50156, 16'd23708, 16'd44482, 16'd49947, 16'd10856, 16'd766, 16'd37668, 16'd39262, 16'd53384, 16'd2134, 16'd60398, 16'd1414, 16'd19511, 16'd41581, 16'd30450, 16'd50898, 16'd34838, 16'd37525, 16'd34258, 16'd7126, 16'd29926, 16'd15279, 16'd47742, 16'd25459, 16'd51654});
	test_expansion(128'h2d49bc4e07fbc99b60ffcb42249dfdd4, {16'd36347, 16'd8662, 16'd3268, 16'd38740, 16'd58767, 16'd19351, 16'd12514, 16'd15598, 16'd4251, 16'd20784, 16'd14045, 16'd26485, 16'd2030, 16'd56895, 16'd36846, 16'd56729, 16'd58165, 16'd5679, 16'd37940, 16'd20902, 16'd33488, 16'd10078, 16'd29576, 16'd8281, 16'd58475, 16'd22331});
	test_expansion(128'h259d81403c842deaf68cd2fabd26e4ec, {16'd21741, 16'd15649, 16'd24994, 16'd43343, 16'd40987, 16'd16995, 16'd7624, 16'd12854, 16'd40906, 16'd39763, 16'd63577, 16'd45015, 16'd62351, 16'd30111, 16'd3627, 16'd61306, 16'd30521, 16'd24496, 16'd20056, 16'd54949, 16'd41071, 16'd54028, 16'd37186, 16'd35993, 16'd18376, 16'd8159});
	test_expansion(128'h906a163c741dc223302442b96e8b70dd, {16'd55590, 16'd14438, 16'd61113, 16'd48327, 16'd52983, 16'd12285, 16'd58272, 16'd21798, 16'd43744, 16'd26716, 16'd34725, 16'd9410, 16'd21265, 16'd1012, 16'd13046, 16'd65118, 16'd30353, 16'd56889, 16'd52756, 16'd18622, 16'd13949, 16'd21390, 16'd44881, 16'd53003, 16'd28333, 16'd24248});
	test_expansion(128'h35a081ef50c719eb467544fef8d12361, {16'd52575, 16'd63453, 16'd49763, 16'd27345, 16'd4975, 16'd61610, 16'd48956, 16'd30436, 16'd22170, 16'd42391, 16'd22545, 16'd56542, 16'd4401, 16'd35123, 16'd17124, 16'd12492, 16'd60404, 16'd32656, 16'd33277, 16'd24057, 16'd53308, 16'd33937, 16'd22943, 16'd11189, 16'd64361, 16'd18787});
	test_expansion(128'h3a0dcdb8f865be3ac025fc6680c64e33, {16'd16576, 16'd10861, 16'd50854, 16'd51019, 16'd5207, 16'd5671, 16'd9952, 16'd6562, 16'd50905, 16'd26867, 16'd65508, 16'd25978, 16'd44346, 16'd37245, 16'd28801, 16'd7922, 16'd125, 16'd4569, 16'd30897, 16'd38478, 16'd27594, 16'd35724, 16'd19037, 16'd41401, 16'd58565, 16'd2009});
	test_expansion(128'h68e1d900be3ba5ebbbad90cb202f174e, {16'd64778, 16'd11714, 16'd3176, 16'd54394, 16'd32500, 16'd51258, 16'd60765, 16'd58827, 16'd42672, 16'd7526, 16'd42916, 16'd23649, 16'd25776, 16'd23467, 16'd38847, 16'd2722, 16'd47806, 16'd53551, 16'd49545, 16'd47498, 16'd58619, 16'd20339, 16'd42356, 16'd25717, 16'd46251, 16'd10224});
	test_expansion(128'hc18baf4596d5f30bb431cbf755cc6b62, {16'd17158, 16'd27445, 16'd65068, 16'd28761, 16'd48880, 16'd9996, 16'd15582, 16'd42965, 16'd36175, 16'd56580, 16'd14409, 16'd20706, 16'd7724, 16'd18126, 16'd52230, 16'd20336, 16'd11363, 16'd12967, 16'd33143, 16'd9726, 16'd28298, 16'd853, 16'd47392, 16'd15770, 16'd42091, 16'd165});
	test_expansion(128'h2161ad6d5178aaa6aaf9bae4e214feb5, {16'd27171, 16'd58001, 16'd14315, 16'd15224, 16'd14435, 16'd49249, 16'd34668, 16'd32561, 16'd37643, 16'd27178, 16'd11079, 16'd10260, 16'd34647, 16'd61230, 16'd46210, 16'd24868, 16'd38306, 16'd55154, 16'd7387, 16'd3956, 16'd53085, 16'd6989, 16'd58513, 16'd65065, 16'd2102, 16'd2097});
	test_expansion(128'hc2a7033dc94770b7fd20e4032d2d886d, {16'd11522, 16'd52581, 16'd40540, 16'd59534, 16'd60788, 16'd37693, 16'd12791, 16'd65202, 16'd58247, 16'd29925, 16'd5177, 16'd62469, 16'd8459, 16'd31968, 16'd39028, 16'd35469, 16'd58850, 16'd38003, 16'd15890, 16'd63610, 16'd58118, 16'd3365, 16'd25847, 16'd6644, 16'd6059, 16'd58881});
	test_expansion(128'hb3eff25139c7fce2d116070b00854c09, {16'd54208, 16'd36168, 16'd23146, 16'd39510, 16'd53524, 16'd13502, 16'd49612, 16'd27819, 16'd51042, 16'd56922, 16'd18005, 16'd19109, 16'd55619, 16'd47815, 16'd18135, 16'd34080, 16'd14456, 16'd36464, 16'd39736, 16'd44096, 16'd57423, 16'd33477, 16'd40275, 16'd16254, 16'd7695, 16'd19947});
	test_expansion(128'h88a7b342ec7b48a44d3d573735214d9c, {16'd37264, 16'd36682, 16'd51990, 16'd29338, 16'd43954, 16'd28825, 16'd63910, 16'd49133, 16'd5112, 16'd22955, 16'd44914, 16'd5329, 16'd3885, 16'd63436, 16'd45547, 16'd48748, 16'd40391, 16'd23326, 16'd62140, 16'd16482, 16'd12523, 16'd8618, 16'd17926, 16'd56052, 16'd3899, 16'd3972});
	test_expansion(128'h9b07805655ca8ea5d9e1ba6bdbe9b3bf, {16'd5585, 16'd8040, 16'd31946, 16'd30186, 16'd174, 16'd58422, 16'd37481, 16'd64758, 16'd37461, 16'd8196, 16'd40812, 16'd2938, 16'd53731, 16'd48500, 16'd2511, 16'd2187, 16'd3270, 16'd22567, 16'd63297, 16'd44420, 16'd56882, 16'd16960, 16'd60441, 16'd33403, 16'd34981, 16'd44093});
	test_expansion(128'h98759bc71da539a92f586ffa710adbfa, {16'd46989, 16'd53879, 16'd59137, 16'd52129, 16'd33902, 16'd30739, 16'd26235, 16'd57303, 16'd3434, 16'd9876, 16'd60064, 16'd41360, 16'd56318, 16'd12638, 16'd43630, 16'd36107, 16'd62525, 16'd7167, 16'd49644, 16'd9577, 16'd29207, 16'd45170, 16'd1182, 16'd35570, 16'd38176, 16'd10346});
	test_expansion(128'hf7fe3284465f7404e4748c3c53d03f37, {16'd20405, 16'd41032, 16'd23637, 16'd57845, 16'd3212, 16'd6145, 16'd22368, 16'd8663, 16'd57786, 16'd33463, 16'd40582, 16'd7452, 16'd32157, 16'd20107, 16'd37048, 16'd3272, 16'd45492, 16'd23457, 16'd62365, 16'd31119, 16'd126, 16'd52905, 16'd7975, 16'd7337, 16'd42832, 16'd28127});
	test_expansion(128'hd1d2aeeacd32d6883854bf7d3a660eb6, {16'd42269, 16'd53679, 16'd64873, 16'd6988, 16'd50846, 16'd50203, 16'd46158, 16'd34566, 16'd29148, 16'd13383, 16'd22821, 16'd17125, 16'd25347, 16'd41422, 16'd43180, 16'd45970, 16'd29839, 16'd29853, 16'd59480, 16'd62414, 16'd14694, 16'd37634, 16'd9882, 16'd33411, 16'd54091, 16'd785});
	test_expansion(128'h687432c08f9eee7f89d39505909a8f6f, {16'd52369, 16'd56731, 16'd42746, 16'd5259, 16'd63481, 16'd45194, 16'd8228, 16'd9578, 16'd8075, 16'd35738, 16'd15111, 16'd1705, 16'd32515, 16'd20406, 16'd47171, 16'd2531, 16'd64230, 16'd28652, 16'd53506, 16'd14289, 16'd7286, 16'd43541, 16'd12958, 16'd14109, 16'd34387, 16'd6293});
	test_expansion(128'h629cbea305c1d7c8e0a9b49152a95341, {16'd34088, 16'd981, 16'd64934, 16'd49795, 16'd28106, 16'd31177, 16'd3178, 16'd59231, 16'd29964, 16'd47025, 16'd33858, 16'd12048, 16'd48918, 16'd43022, 16'd63940, 16'd31124, 16'd49259, 16'd6509, 16'd54924, 16'd60139, 16'd55095, 16'd12275, 16'd43457, 16'd1086, 16'd58421, 16'd25195});
	test_expansion(128'heb527856570ac02dfe2766d9fe26efc1, {16'd51449, 16'd85, 16'd15692, 16'd21531, 16'd55815, 16'd22479, 16'd9092, 16'd4565, 16'd46087, 16'd13554, 16'd8957, 16'd56009, 16'd32455, 16'd54722, 16'd36836, 16'd13256, 16'd25498, 16'd58799, 16'd60494, 16'd8434, 16'd53972, 16'd6528, 16'd25032, 16'd14896, 16'd31383, 16'd23990});
	test_expansion(128'h79d8182dd40eeb329758a7b3c4d23216, {16'd50592, 16'd26302, 16'd7724, 16'd15806, 16'd56067, 16'd11305, 16'd292, 16'd24570, 16'd944, 16'd34073, 16'd10083, 16'd35090, 16'd34975, 16'd54834, 16'd56598, 16'd41092, 16'd48209, 16'd7642, 16'd21042, 16'd50579, 16'd55460, 16'd20303, 16'd60056, 16'd3257, 16'd55134, 16'd42882});
	test_expansion(128'ha36d02c170d54946c30ea4dc8c2e07b2, {16'd19921, 16'd35495, 16'd21884, 16'd64161, 16'd19561, 16'd64588, 16'd16506, 16'd13155, 16'd64621, 16'd48664, 16'd27674, 16'd10128, 16'd19186, 16'd38332, 16'd34610, 16'd33441, 16'd60435, 16'd22992, 16'd19815, 16'd22155, 16'd4425, 16'd14502, 16'd12844, 16'd33631, 16'd10585, 16'd42727});
	test_expansion(128'hff5aa76ef9a37c7bede3bb66da8131e6, {16'd44270, 16'd59215, 16'd54562, 16'd37011, 16'd50882, 16'd17234, 16'd17107, 16'd53494, 16'd41174, 16'd32564, 16'd25264, 16'd51654, 16'd30116, 16'd44276, 16'd19966, 16'd60507, 16'd14862, 16'd32508, 16'd57185, 16'd37051, 16'd27479, 16'd36523, 16'd57446, 16'd36756, 16'd62368, 16'd3486});
	test_expansion(128'h2172ccad7ae3f5847d7fbfdc02c6d771, {16'd8331, 16'd1202, 16'd55187, 16'd34307, 16'd41389, 16'd46980, 16'd52722, 16'd20941, 16'd22100, 16'd52014, 16'd47245, 16'd22986, 16'd39914, 16'd39357, 16'd28430, 16'd12690, 16'd37843, 16'd52253, 16'd36428, 16'd7063, 16'd10528, 16'd42581, 16'd16477, 16'd47384, 16'd44055, 16'd55157});
	test_expansion(128'hd8d98251e944c4539a68e2aae60f2f30, {16'd1053, 16'd5182, 16'd33996, 16'd49209, 16'd33677, 16'd37708, 16'd48870, 16'd11994, 16'd39915, 16'd2905, 16'd15974, 16'd12148, 16'd51543, 16'd39200, 16'd7301, 16'd31406, 16'd30086, 16'd12820, 16'd58949, 16'd169, 16'd64142, 16'd62036, 16'd3434, 16'd16600, 16'd53837, 16'd63126});
	test_expansion(128'hdab2007550a1af0ee80d022eededc1a7, {16'd3779, 16'd52129, 16'd8424, 16'd39967, 16'd32349, 16'd56965, 16'd65381, 16'd648, 16'd27913, 16'd47273, 16'd20441, 16'd25179, 16'd60733, 16'd14911, 16'd41748, 16'd59197, 16'd40541, 16'd29937, 16'd18407, 16'd25392, 16'd26028, 16'd28811, 16'd37530, 16'd53912, 16'd15673, 16'd57641});
	test_expansion(128'h0cbaf82e230f3c30997470fba11a9d57, {16'd17619, 16'd12645, 16'd2843, 16'd64438, 16'd59834, 16'd58008, 16'd56658, 16'd33738, 16'd1664, 16'd47448, 16'd65181, 16'd46456, 16'd34544, 16'd46798, 16'd36877, 16'd19483, 16'd38439, 16'd12637, 16'd23154, 16'd45710, 16'd27441, 16'd65036, 16'd12575, 16'd4402, 16'd9910, 16'd34002});
	test_expansion(128'ha0642fe2b0a725e4f0b71e81d4857bdc, {16'd45662, 16'd32873, 16'd50070, 16'd1955, 16'd36271, 16'd35198, 16'd37587, 16'd21381, 16'd14720, 16'd8711, 16'd30736, 16'd11994, 16'd28325, 16'd36769, 16'd59165, 16'd22548, 16'd38002, 16'd12917, 16'd12947, 16'd51332, 16'd59084, 16'd56162, 16'd64452, 16'd61555, 16'd19397, 16'd46722});
	test_expansion(128'hde5e10048fe6b6d0b2c6c55c7048989c, {16'd11733, 16'd44410, 16'd28647, 16'd57901, 16'd35362, 16'd13488, 16'd7626, 16'd54903, 16'd55153, 16'd31754, 16'd4713, 16'd59044, 16'd36528, 16'd42238, 16'd52376, 16'd57657, 16'd32117, 16'd18335, 16'd48776, 16'd45550, 16'd17603, 16'd7630, 16'd39224, 16'd47915, 16'd7886, 16'd60974});
	test_expansion(128'hbc7775f719c0b653c2ff20dbb01db494, {16'd65007, 16'd64950, 16'd29576, 16'd34672, 16'd23232, 16'd4886, 16'd62886, 16'd53758, 16'd35855, 16'd64862, 16'd63141, 16'd38679, 16'd54048, 16'd19473, 16'd49153, 16'd65154, 16'd33822, 16'd16820, 16'd65389, 16'd22107, 16'd12406, 16'd50295, 16'd43643, 16'd59474, 16'd20267, 16'd43298});
	test_expansion(128'h96230c68fcada2621a569c54c17c3674, {16'd43562, 16'd31567, 16'd64900, 16'd30931, 16'd60999, 16'd63652, 16'd24118, 16'd26864, 16'd34070, 16'd34794, 16'd52020, 16'd42215, 16'd34587, 16'd43299, 16'd16527, 16'd36123, 16'd27300, 16'd63048, 16'd61644, 16'd4047, 16'd2198, 16'd16130, 16'd24135, 16'd30103, 16'd6699, 16'd21011});
	test_expansion(128'hda174610e3dbbe8d3051285d140cbaab, {16'd22485, 16'd16164, 16'd24837, 16'd4593, 16'd52667, 16'd12724, 16'd39825, 16'd52562, 16'd51899, 16'd2162, 16'd5605, 16'd56296, 16'd49177, 16'd18480, 16'd23092, 16'd26908, 16'd65353, 16'd10948, 16'd39189, 16'd11384, 16'd37582, 16'd41852, 16'd32798, 16'd33404, 16'd8265, 16'd49430});
	test_expansion(128'h9a62cdd83728aa48dac9a6810c1b24da, {16'd60526, 16'd22079, 16'd11693, 16'd49060, 16'd41525, 16'd20977, 16'd47395, 16'd24171, 16'd19542, 16'd10395, 16'd39355, 16'd51556, 16'd18690, 16'd54392, 16'd52759, 16'd7858, 16'd6681, 16'd33012, 16'd29481, 16'd25778, 16'd41744, 16'd57425, 16'd60714, 16'd57744, 16'd20204, 16'd61217});
	test_expansion(128'hf69e39ae662d30abf9cf3fb9ebd5c831, {16'd12728, 16'd63814, 16'd98, 16'd34596, 16'd32364, 16'd52013, 16'd50945, 16'd47090, 16'd42193, 16'd2957, 16'd36449, 16'd25308, 16'd20089, 16'd35670, 16'd15104, 16'd14124, 16'd59267, 16'd18679, 16'd16033, 16'd14676, 16'd6896, 16'd42041, 16'd59093, 16'd49388, 16'd22145, 16'd43362});
	test_expansion(128'h5837e2e49a68b39e1b56ec3701b5b0f5, {16'd36568, 16'd55594, 16'd47113, 16'd57994, 16'd12476, 16'd17901, 16'd24105, 16'd30634, 16'd22601, 16'd54964, 16'd3057, 16'd54987, 16'd15348, 16'd63050, 16'd12221, 16'd28500, 16'd12785, 16'd62681, 16'd39482, 16'd25041, 16'd37492, 16'd35648, 16'd41630, 16'd740, 16'd33156, 16'd27477});
	test_expansion(128'ha831dca9b2697112082d6ab90ff7f20a, {16'd19676, 16'd57877, 16'd2203, 16'd1128, 16'd13952, 16'd12916, 16'd3579, 16'd4330, 16'd9482, 16'd51728, 16'd19309, 16'd22189, 16'd57021, 16'd36654, 16'd37821, 16'd61880, 16'd58588, 16'd7963, 16'd65503, 16'd8651, 16'd55304, 16'd44792, 16'd33152, 16'd29103, 16'd47825, 16'd43999});
	test_expansion(128'hcf10dd88ccdfe29e3fc32105b235408b, {16'd15419, 16'd1727, 16'd56438, 16'd64373, 16'd53042, 16'd18078, 16'd8996, 16'd48249, 16'd39355, 16'd56179, 16'd4195, 16'd15178, 16'd4371, 16'd21703, 16'd12555, 16'd18435, 16'd56004, 16'd46664, 16'd13899, 16'd11940, 16'd37728, 16'd46848, 16'd15370, 16'd21661, 16'd39307, 16'd12493});
	test_expansion(128'hb6ed425f3d49ab8eb40403b28344a240, {16'd19020, 16'd36933, 16'd18506, 16'd33703, 16'd47641, 16'd44568, 16'd29786, 16'd15955, 16'd27456, 16'd53857, 16'd49558, 16'd47648, 16'd62359, 16'd27653, 16'd55460, 16'd23467, 16'd9264, 16'd13825, 16'd55759, 16'd8186, 16'd3201, 16'd16366, 16'd26214, 16'd40903, 16'd27014, 16'd58303});
	test_expansion(128'h36e8a00320c74e253608d7a66986cd82, {16'd35976, 16'd19771, 16'd8286, 16'd28399, 16'd8841, 16'd44479, 16'd26109, 16'd24808, 16'd10443, 16'd33762, 16'd14967, 16'd59048, 16'd38032, 16'd61107, 16'd50976, 16'd51285, 16'd51462, 16'd8713, 16'd59190, 16'd18183, 16'd793, 16'd24160, 16'd28850, 16'd61081, 16'd11532, 16'd60847});
	test_expansion(128'h9a2f4184f9c4ee51d0aebddcbd8a6f8a, {16'd18641, 16'd52362, 16'd14996, 16'd7016, 16'd23564, 16'd6118, 16'd53660, 16'd1746, 16'd678, 16'd1368, 16'd31174, 16'd33241, 16'd37618, 16'd59091, 16'd15467, 16'd48584, 16'd17002, 16'd28087, 16'd29266, 16'd51568, 16'd39520, 16'd28632, 16'd38034, 16'd57592, 16'd22411, 16'd57704});
	test_expansion(128'hdee2a4423213c23424bf0e7c76193e03, {16'd41514, 16'd6776, 16'd54918, 16'd11698, 16'd41697, 16'd8555, 16'd6579, 16'd53391, 16'd16368, 16'd14936, 16'd51549, 16'd51595, 16'd42540, 16'd2887, 16'd43372, 16'd29366, 16'd39968, 16'd25734, 16'd14462, 16'd3841, 16'd18004, 16'd62024, 16'd616, 16'd50750, 16'd36611, 16'd49844});
	test_expansion(128'h837ed6a3a8db80712731b8c5f577130b, {16'd5017, 16'd7594, 16'd9508, 16'd39346, 16'd63142, 16'd50626, 16'd35527, 16'd4669, 16'd35604, 16'd20240, 16'd61980, 16'd4804, 16'd17902, 16'd35552, 16'd34395, 16'd55220, 16'd40191, 16'd43, 16'd35349, 16'd15295, 16'd32437, 16'd19783, 16'd25973, 16'd20089, 16'd58831, 16'd34281});
	test_expansion(128'h644599e5bd529feefeebc948877d0602, {16'd38516, 16'd26247, 16'd45172, 16'd52332, 16'd62117, 16'd27248, 16'd763, 16'd21389, 16'd21271, 16'd49507, 16'd15418, 16'd19073, 16'd33348, 16'd21931, 16'd51198, 16'd36780, 16'd2652, 16'd41123, 16'd36441, 16'd52203, 16'd59526, 16'd34727, 16'd18199, 16'd28982, 16'd27698, 16'd8180});
	test_expansion(128'hc46d88e02a0f0712321e514677fb0542, {16'd14904, 16'd12904, 16'd20291, 16'd16308, 16'd6988, 16'd17487, 16'd40732, 16'd10847, 16'd9241, 16'd24237, 16'd33664, 16'd58169, 16'd59163, 16'd48797, 16'd64145, 16'd49814, 16'd36293, 16'd43559, 16'd24179, 16'd53543, 16'd10764, 16'd55542, 16'd47482, 16'd13556, 16'd2943, 16'd18238});
	test_expansion(128'h01760f63fcc2cd292b88b0a685579a33, {16'd2085, 16'd49916, 16'd62587, 16'd48226, 16'd2901, 16'd17464, 16'd7190, 16'd2739, 16'd58555, 16'd26210, 16'd40642, 16'd51308, 16'd32500, 16'd51153, 16'd36874, 16'd41146, 16'd30583, 16'd51898, 16'd11885, 16'd6268, 16'd48497, 16'd31728, 16'd43030, 16'd49359, 16'd6735, 16'd46590});
	test_expansion(128'h13fc90c83f180eaf42e7cdd1c2f81264, {16'd43702, 16'd35053, 16'd44204, 16'd9287, 16'd3227, 16'd58460, 16'd59854, 16'd64681, 16'd26071, 16'd41880, 16'd63605, 16'd40767, 16'd529, 16'd1950, 16'd18087, 16'd57316, 16'd17507, 16'd38144, 16'd64599, 16'd17329, 16'd51343, 16'd64793, 16'd50544, 16'd59190, 16'd28655, 16'd1157});
	test_expansion(128'h96937dfa6a0b961b5ceaed2326070fd2, {16'd49584, 16'd56189, 16'd53794, 16'd27934, 16'd37803, 16'd56233, 16'd58758, 16'd11516, 16'd59058, 16'd17757, 16'd44739, 16'd1084, 16'd41752, 16'd22297, 16'd33914, 16'd15891, 16'd2412, 16'd57411, 16'd23788, 16'd29095, 16'd56381, 16'd468, 16'd41581, 16'd30239, 16'd54628, 16'd63244});
	test_expansion(128'h5b9857f6059893d9ec9e3d8f39e142c9, {16'd55593, 16'd32193, 16'd40577, 16'd63853, 16'd6311, 16'd18149, 16'd50156, 16'd8678, 16'd1773, 16'd38139, 16'd36223, 16'd32325, 16'd16747, 16'd34741, 16'd21977, 16'd50805, 16'd33749, 16'd12484, 16'd2762, 16'd48166, 16'd43360, 16'd28320, 16'd9523, 16'd23718, 16'd5014, 16'd47892});
	test_expansion(128'h2ca77a06aeb0a21cb69011c83a160bf3, {16'd26641, 16'd47377, 16'd3178, 16'd14182, 16'd28061, 16'd28223, 16'd37464, 16'd56450, 16'd6481, 16'd43207, 16'd62446, 16'd61335, 16'd38582, 16'd43469, 16'd25363, 16'd19396, 16'd56969, 16'd39446, 16'd27003, 16'd30637, 16'd60501, 16'd7122, 16'd2302, 16'd42784, 16'd8114, 16'd39552});
	test_expansion(128'hbb3c55dac764b0200cbc162098bf3dc6, {16'd30560, 16'd17309, 16'd23220, 16'd27107, 16'd62977, 16'd50825, 16'd3262, 16'd63450, 16'd5247, 16'd57374, 16'd62815, 16'd47298, 16'd27721, 16'd8855, 16'd21257, 16'd37956, 16'd46150, 16'd34691, 16'd2276, 16'd65235, 16'd3610, 16'd31525, 16'd21420, 16'd4062, 16'd56225, 16'd22360});
	test_expansion(128'hc04208c478a1a9dec6b50c9cd8f675c9, {16'd57526, 16'd64181, 16'd17271, 16'd25534, 16'd21364, 16'd29015, 16'd3986, 16'd62010, 16'd29596, 16'd20394, 16'd18059, 16'd32457, 16'd9631, 16'd9401, 16'd3036, 16'd14516, 16'd29, 16'd36317, 16'd12968, 16'd57671, 16'd2504, 16'd2549, 16'd63257, 16'd31119, 16'd15734, 16'd35184});
	test_expansion(128'h789ef5f77697653fbc02193a245b359a, {16'd25395, 16'd51495, 16'd13870, 16'd9388, 16'd62069, 16'd21882, 16'd33731, 16'd33970, 16'd37716, 16'd53395, 16'd835, 16'd59766, 16'd11735, 16'd17213, 16'd57657, 16'd61637, 16'd7561, 16'd21950, 16'd55366, 16'd61185, 16'd11043, 16'd21427, 16'd64352, 16'd5122, 16'd20142, 16'd34531});
	test_expansion(128'hb2eb9cf81484dfbde9ffda8400a8fa2f, {16'd53164, 16'd18365, 16'd43581, 16'd39565, 16'd34744, 16'd63750, 16'd28089, 16'd14080, 16'd17687, 16'd48504, 16'd3278, 16'd62805, 16'd56691, 16'd13555, 16'd55617, 16'd63785, 16'd53024, 16'd55630, 16'd43463, 16'd30005, 16'd9047, 16'd25261, 16'd41474, 16'd21178, 16'd38757, 16'd64674});
	test_expansion(128'hf0e55e9834502417234dffc5683624e2, {16'd20312, 16'd46157, 16'd19336, 16'd42676, 16'd42922, 16'd145, 16'd56653, 16'd16439, 16'd65074, 16'd57474, 16'd54847, 16'd3036, 16'd5352, 16'd47649, 16'd15022, 16'd37680, 16'd60951, 16'd23698, 16'd63906, 16'd52257, 16'd62458, 16'd41162, 16'd29772, 16'd45070, 16'd25153, 16'd52578});
	test_expansion(128'h772ee68d1f162478028b3271b9d15219, {16'd37445, 16'd44843, 16'd6263, 16'd13027, 16'd44031, 16'd63717, 16'd41440, 16'd55204, 16'd11285, 16'd3729, 16'd87, 16'd8446, 16'd10750, 16'd35179, 16'd62833, 16'd31811, 16'd10385, 16'd39652, 16'd22909, 16'd55669, 16'd16333, 16'd24703, 16'd43444, 16'd15006, 16'd11590, 16'd43430});
	test_expansion(128'hb6a15594f78663772782da16f422ee1f, {16'd52034, 16'd52100, 16'd12945, 16'd42085, 16'd62566, 16'd50948, 16'd36152, 16'd41022, 16'd14316, 16'd48338, 16'd12277, 16'd11605, 16'd34705, 16'd65534, 16'd60957, 16'd56987, 16'd40718, 16'd51580, 16'd19577, 16'd19637, 16'd17381, 16'd55675, 16'd6890, 16'd39091, 16'd51526, 16'd63760});
	test_expansion(128'h601ee781c53572579df24696c6addc1d, {16'd3636, 16'd51865, 16'd38029, 16'd1247, 16'd19670, 16'd11375, 16'd20351, 16'd61915, 16'd14159, 16'd13795, 16'd33666, 16'd37221, 16'd41180, 16'd39705, 16'd14883, 16'd62809, 16'd62429, 16'd1547, 16'd57, 16'd61882, 16'd45074, 16'd54669, 16'd25351, 16'd54968, 16'd3200, 16'd51403});
	test_expansion(128'ha6d3bb5101de34b5ddc8887a6dc846c9, {16'd17426, 16'd39166, 16'd11729, 16'd5184, 16'd23620, 16'd15804, 16'd41076, 16'd35204, 16'd32852, 16'd19357, 16'd60460, 16'd28404, 16'd35011, 16'd58609, 16'd29587, 16'd18356, 16'd35858, 16'd10597, 16'd45779, 16'd33814, 16'd26409, 16'd59000, 16'd61811, 16'd8424, 16'd29789, 16'd50895});
	test_expansion(128'hc21e781c2268166d11cb93d8ac710144, {16'd39311, 16'd43801, 16'd3503, 16'd23206, 16'd5486, 16'd36480, 16'd58039, 16'd11145, 16'd40755, 16'd40493, 16'd64564, 16'd30989, 16'd54810, 16'd40181, 16'd32580, 16'd15422, 16'd4696, 16'd6229, 16'd12784, 16'd35021, 16'd53116, 16'd36723, 16'd23941, 16'd25226, 16'd17380, 16'd523});
	test_expansion(128'h92ed17e7b19953196cb9a3b62f5c220b, {16'd16599, 16'd916, 16'd24656, 16'd61701, 16'd36864, 16'd43169, 16'd21469, 16'd53126, 16'd59161, 16'd12891, 16'd3942, 16'd1156, 16'd39372, 16'd12140, 16'd20129, 16'd9285, 16'd1170, 16'd34885, 16'd3883, 16'd6894, 16'd2456, 16'd12734, 16'd22815, 16'd5410, 16'd6335, 16'd52710});
	test_expansion(128'h34d8e86f64ebe54e4566fdb3a7355060, {16'd54455, 16'd14703, 16'd57201, 16'd45411, 16'd8085, 16'd11203, 16'd5850, 16'd12434, 16'd24885, 16'd28546, 16'd14800, 16'd9468, 16'd48038, 16'd41044, 16'd62486, 16'd56754, 16'd708, 16'd15615, 16'd33052, 16'd22609, 16'd31961, 16'd45814, 16'd19793, 16'd35116, 16'd24704, 16'd43257});
	test_expansion(128'hb41eb5746ec0fe370002209337741ba9, {16'd14050, 16'd36239, 16'd6466, 16'd29547, 16'd43752, 16'd45267, 16'd34364, 16'd55960, 16'd56976, 16'd10106, 16'd58093, 16'd52771, 16'd38604, 16'd10976, 16'd46227, 16'd53849, 16'd23669, 16'd27440, 16'd45418, 16'd53727, 16'd25668, 16'd24373, 16'd7892, 16'd30388, 16'd62988, 16'd64329});
	test_expansion(128'h89f02ff4bf8bc6136c86eb66b46768a0, {16'd58239, 16'd26226, 16'd35695, 16'd2266, 16'd12645, 16'd41390, 16'd54009, 16'd32350, 16'd37021, 16'd39285, 16'd30384, 16'd62801, 16'd57449, 16'd30691, 16'd18206, 16'd9361, 16'd31930, 16'd62043, 16'd61460, 16'd14784, 16'd47771, 16'd32469, 16'd49426, 16'd18472, 16'd13848, 16'd6572});
	test_expansion(128'h6afef431460a7a2b31e74bc08f95788d, {16'd16786, 16'd43800, 16'd32696, 16'd43371, 16'd25356, 16'd53518, 16'd58399, 16'd16381, 16'd43337, 16'd2756, 16'd60315, 16'd62547, 16'd9827, 16'd16365, 16'd51, 16'd50723, 16'd57926, 16'd17537, 16'd10031, 16'd56694, 16'd24891, 16'd51255, 16'd43262, 16'd20463, 16'd54364, 16'd7371});
	test_expansion(128'h41fecf7fb6ff2be16de41d2f6e9f5d06, {16'd52059, 16'd63381, 16'd4906, 16'd36661, 16'd38077, 16'd18913, 16'd49493, 16'd20743, 16'd62740, 16'd3082, 16'd30488, 16'd7598, 16'd14560, 16'd10802, 16'd16267, 16'd49526, 16'd21803, 16'd12590, 16'd21127, 16'd49871, 16'd25328, 16'd43381, 16'd49150, 16'd35485, 16'd57866, 16'd18016});
	test_expansion(128'h94b019f8994634eed639d04301e9d7b4, {16'd38476, 16'd43031, 16'd27277, 16'd48277, 16'd31388, 16'd6621, 16'd64667, 16'd44584, 16'd24565, 16'd25815, 16'd46162, 16'd25390, 16'd21822, 16'd21240, 16'd2091, 16'd45624, 16'd2803, 16'd18627, 16'd10087, 16'd58889, 16'd64462, 16'd60509, 16'd5892, 16'd29990, 16'd29421, 16'd36788});
	test_expansion(128'ha6830bb2c51b95e65d7836351d536e3d, {16'd48943, 16'd58790, 16'd7257, 16'd54570, 16'd2401, 16'd20230, 16'd12747, 16'd58865, 16'd10217, 16'd38611, 16'd64245, 16'd63647, 16'd34060, 16'd11321, 16'd6659, 16'd6807, 16'd61054, 16'd49600, 16'd14481, 16'd1242, 16'd31116, 16'd35843, 16'd11404, 16'd4318, 16'd23716, 16'd23111});
	test_expansion(128'h8d02efd15073482cc1f3b39949050b6e, {16'd31189, 16'd44797, 16'd53111, 16'd14114, 16'd45677, 16'd19079, 16'd64899, 16'd14289, 16'd52221, 16'd44135, 16'd60077, 16'd33629, 16'd14013, 16'd14767, 16'd24317, 16'd45944, 16'd16776, 16'd43085, 16'd437, 16'd30818, 16'd14662, 16'd43020, 16'd24622, 16'd49947, 16'd41759, 16'd36992});
	test_expansion(128'h0590cab4a4dd6cc4a4bbfc0b3e613f54, {16'd12617, 16'd7758, 16'd18745, 16'd50989, 16'd14833, 16'd39917, 16'd56459, 16'd36203, 16'd4136, 16'd18067, 16'd32348, 16'd43504, 16'd10944, 16'd36436, 16'd62041, 16'd16801, 16'd9570, 16'd15264, 16'd19470, 16'd23002, 16'd5419, 16'd3707, 16'd17974, 16'd58172, 16'd60909, 16'd10982});
	test_expansion(128'ha4ceca35f4779a7e88c3a9abca283f48, {16'd56568, 16'd47380, 16'd57027, 16'd59760, 16'd36396, 16'd15575, 16'd22618, 16'd49095, 16'd46038, 16'd15856, 16'd46620, 16'd38524, 16'd31104, 16'd61153, 16'd28291, 16'd33112, 16'd57434, 16'd63568, 16'd50203, 16'd50472, 16'd36262, 16'd5385, 16'd53425, 16'd33656, 16'd49828, 16'd38040});
	test_expansion(128'h50e9e7651692d93c9131ac5cb9c03827, {16'd33125, 16'd43011, 16'd39080, 16'd49184, 16'd62452, 16'd45923, 16'd44958, 16'd45679, 16'd837, 16'd21057, 16'd58964, 16'd55092, 16'd15070, 16'd40896, 16'd5433, 16'd27371, 16'd23771, 16'd21393, 16'd42833, 16'd65159, 16'd28900, 16'd6166, 16'd50992, 16'd56675, 16'd30724, 16'd49230});
	test_expansion(128'hc700ac470da4334673268ac9432c4570, {16'd34355, 16'd48123, 16'd51771, 16'd61757, 16'd8127, 16'd5293, 16'd59129, 16'd41747, 16'd24297, 16'd37907, 16'd18199, 16'd53301, 16'd57132, 16'd19916, 16'd6570, 16'd17971, 16'd30104, 16'd61952, 16'd43382, 16'd15394, 16'd50292, 16'd42117, 16'd6145, 16'd8970, 16'd12300, 16'd17673});
	test_expansion(128'h2b5b339613d73df0d678e3cce2c44065, {16'd508, 16'd53489, 16'd25404, 16'd27107, 16'd3357, 16'd57680, 16'd48607, 16'd29806, 16'd2865, 16'd26313, 16'd55093, 16'd32194, 16'd43162, 16'd46822, 16'd53589, 16'd19755, 16'd61382, 16'd44101, 16'd27700, 16'd54117, 16'd43857, 16'd3374, 16'd43338, 16'd5800, 16'd7682, 16'd8011});
	test_expansion(128'h6bd9088524a5feadad233178ca68aa17, {16'd17320, 16'd59349, 16'd9684, 16'd22041, 16'd10149, 16'd17131, 16'd2388, 16'd32183, 16'd20241, 16'd2038, 16'd50140, 16'd1908, 16'd48021, 16'd18699, 16'd52792, 16'd53224, 16'd57487, 16'd56143, 16'd22984, 16'd32607, 16'd19786, 16'd48602, 16'd11601, 16'd56718, 16'd1679, 16'd22369});
	test_expansion(128'h76adeed4e3f31d67b9aff1fea23bea0d, {16'd54392, 16'd56946, 16'd5646, 16'd16130, 16'd34285, 16'd61965, 16'd15205, 16'd34308, 16'd58498, 16'd61166, 16'd58363, 16'd54766, 16'd9624, 16'd59292, 16'd15118, 16'd33217, 16'd18533, 16'd54767, 16'd19896, 16'd43625, 16'd46872, 16'd39768, 16'd49655, 16'd60157, 16'd24259, 16'd12518});
	test_expansion(128'h18b1f97a567290b00a77842b466306ea, {16'd53943, 16'd11987, 16'd21947, 16'd56856, 16'd703, 16'd37425, 16'd52724, 16'd41816, 16'd36248, 16'd14225, 16'd27802, 16'd28331, 16'd63593, 16'd21527, 16'd39624, 16'd6484, 16'd17246, 16'd48165, 16'd11808, 16'd34181, 16'd49365, 16'd12602, 16'd37727, 16'd27865, 16'd13566, 16'd60332});
	test_expansion(128'h91d369c0cf4a1fbb153ca5e0e8220416, {16'd49467, 16'd1301, 16'd37318, 16'd21926, 16'd5351, 16'd21123, 16'd36953, 16'd24108, 16'd56968, 16'd57657, 16'd3311, 16'd54556, 16'd17717, 16'd64431, 16'd28636, 16'd448, 16'd20379, 16'd38792, 16'd21070, 16'd61435, 16'd36186, 16'd8601, 16'd62321, 16'd54971, 16'd3741, 16'd4944});
	test_expansion(128'h41dc45c8aebff393dbe164eb00b6df28, {16'd59674, 16'd1681, 16'd15213, 16'd33801, 16'd17905, 16'd6259, 16'd6250, 16'd56886, 16'd44649, 16'd63735, 16'd4260, 16'd59706, 16'd34572, 16'd11720, 16'd53162, 16'd21602, 16'd21519, 16'd45023, 16'd60609, 16'd39957, 16'd56632, 16'd54541, 16'd45999, 16'd27404, 16'd41767, 16'd60731});
	test_expansion(128'hc7a476c4480ca19185391178065df428, {16'd60468, 16'd35014, 16'd24750, 16'd1725, 16'd9167, 16'd9306, 16'd4640, 16'd9828, 16'd3575, 16'd11203, 16'd42388, 16'd62773, 16'd61733, 16'd27559, 16'd27874, 16'd15296, 16'd46372, 16'd60444, 16'd38960, 16'd50441, 16'd15008, 16'd64117, 16'd7277, 16'd64014, 16'd36417, 16'd7338});
	test_expansion(128'hcfe602f0a4e32ea8008c1009816e1d68, {16'd9522, 16'd20992, 16'd60695, 16'd1555, 16'd40293, 16'd48122, 16'd47627, 16'd1228, 16'd25926, 16'd61904, 16'd55292, 16'd60152, 16'd21520, 16'd42908, 16'd29642, 16'd64246, 16'd10573, 16'd17663, 16'd17383, 16'd58431, 16'd60366, 16'd44580, 16'd35669, 16'd38912, 16'd29387, 16'd21867});
	test_expansion(128'h465ea18533861d9b7689146b08cf59fb, {16'd14136, 16'd65524, 16'd23940, 16'd47870, 16'd33696, 16'd21935, 16'd65426, 16'd62662, 16'd31987, 16'd8749, 16'd41823, 16'd61398, 16'd65021, 16'd9738, 16'd7821, 16'd62480, 16'd47111, 16'd42333, 16'd19354, 16'd48525, 16'd39839, 16'd17297, 16'd38449, 16'd13259, 16'd11692, 16'd61462});
	test_expansion(128'hed11afe2f52e0c7a20c7757cb3c09db2, {16'd63490, 16'd56360, 16'd22436, 16'd11841, 16'd45857, 16'd31220, 16'd64768, 16'd9156, 16'd41038, 16'd44034, 16'd29809, 16'd40719, 16'd22698, 16'd952, 16'd64093, 16'd9287, 16'd14751, 16'd54231, 16'd37544, 16'd57763, 16'd40327, 16'd52641, 16'd28314, 16'd27823, 16'd49542, 16'd21687});
	test_expansion(128'he798ced78f03882e815ea3cf1fc061b2, {16'd33829, 16'd27160, 16'd24747, 16'd32296, 16'd18206, 16'd14003, 16'd32647, 16'd24727, 16'd35920, 16'd34294, 16'd4597, 16'd42905, 16'd58737, 16'd52570, 16'd22953, 16'd32549, 16'd22135, 16'd35968, 16'd52888, 16'd16614, 16'd20541, 16'd58527, 16'd40784, 16'd26962, 16'd62310, 16'd17224});
	test_expansion(128'h796b0d9a3d060c04dd45733f72c09b7f, {16'd27046, 16'd59332, 16'd33144, 16'd23371, 16'd40096, 16'd38303, 16'd47187, 16'd25200, 16'd45487, 16'd9900, 16'd30202, 16'd3853, 16'd13983, 16'd64044, 16'd17554, 16'd58240, 16'd45659, 16'd54348, 16'd34742, 16'd22686, 16'd7471, 16'd37785, 16'd22181, 16'd6849, 16'd34812, 16'd50303});
	test_expansion(128'h498254052d585c2b89da9a238e92b381, {16'd42321, 16'd54023, 16'd1469, 16'd54210, 16'd29128, 16'd61347, 16'd13152, 16'd51926, 16'd39027, 16'd64795, 16'd23504, 16'd11283, 16'd51015, 16'd17730, 16'd34144, 16'd33630, 16'd35199, 16'd51887, 16'd43352, 16'd41828, 16'd8032, 16'd58033, 16'd14297, 16'd6420, 16'd56571, 16'd4719});
	test_expansion(128'hada6583efafa5afbbbfd1b8bbb18fb41, {16'd51438, 16'd4840, 16'd62985, 16'd11774, 16'd9788, 16'd2875, 16'd18492, 16'd51514, 16'd51734, 16'd50449, 16'd29859, 16'd22091, 16'd20907, 16'd57999, 16'd53160, 16'd47450, 16'd22009, 16'd6520, 16'd27717, 16'd17138, 16'd57255, 16'd57884, 16'd22336, 16'd23515, 16'd29496, 16'd28396});
	test_expansion(128'hc03a60954e7b0edbdf2f07ca3a45fc57, {16'd26156, 16'd23137, 16'd29375, 16'd34162, 16'd45663, 16'd24622, 16'd55744, 16'd14823, 16'd4309, 16'd56349, 16'd17503, 16'd10447, 16'd54807, 16'd62093, 16'd4394, 16'd23584, 16'd60288, 16'd5796, 16'd51453, 16'd61658, 16'd54738, 16'd30944, 16'd58801, 16'd56829, 16'd57158, 16'd59591});
	test_expansion(128'hd6347d67ed8a3541bb9b5761a318be6c, {16'd54197, 16'd51309, 16'd37686, 16'd30227, 16'd830, 16'd11492, 16'd12699, 16'd6185, 16'd64858, 16'd50926, 16'd8752, 16'd62121, 16'd38478, 16'd16527, 16'd6018, 16'd46565, 16'd55412, 16'd38028, 16'd7202, 16'd12040, 16'd28515, 16'd246, 16'd21375, 16'd7251, 16'd48378, 16'd64048});
	test_expansion(128'h2998227b04e365e03b687f3cf8bd38f3, {16'd62339, 16'd5967, 16'd32470, 16'd36464, 16'd51185, 16'd34020, 16'd49118, 16'd46644, 16'd8298, 16'd49225, 16'd55840, 16'd33925, 16'd24882, 16'd50112, 16'd35699, 16'd33904, 16'd53491, 16'd17153, 16'd3323, 16'd51722, 16'd59184, 16'd8008, 16'd27498, 16'd38649, 16'd64522, 16'd37861});
	test_expansion(128'h6577fb646ee07d640bec4d22401d9c2c, {16'd39534, 16'd9438, 16'd30569, 16'd60606, 16'd53690, 16'd39646, 16'd44106, 16'd41444, 16'd52182, 16'd31508, 16'd18657, 16'd34515, 16'd18202, 16'd10586, 16'd15925, 16'd15023, 16'd21556, 16'd39176, 16'd62413, 16'd38767, 16'd12878, 16'd14447, 16'd22182, 16'd61115, 16'd28268, 16'd47473});
	test_expansion(128'hfa67e76176d47fc1599c1cca51df9bd1, {16'd11039, 16'd6829, 16'd50483, 16'd36795, 16'd17175, 16'd30069, 16'd22692, 16'd39797, 16'd16219, 16'd22591, 16'd19976, 16'd4096, 16'd8303, 16'd1675, 16'd12259, 16'd47309, 16'd17995, 16'd3941, 16'd42354, 16'd27802, 16'd60176, 16'd43713, 16'd65460, 16'd4624, 16'd25729, 16'd13958});
	test_expansion(128'h86ebdf3aba0fde209778ea3b537a1437, {16'd44327, 16'd20261, 16'd19347, 16'd2634, 16'd22142, 16'd30092, 16'd60385, 16'd32442, 16'd6690, 16'd16283, 16'd58125, 16'd5770, 16'd39001, 16'd51275, 16'd34053, 16'd49810, 16'd1361, 16'd61657, 16'd36796, 16'd5362, 16'd10797, 16'd8481, 16'd47871, 16'd8016, 16'd30565, 16'd43948});
	test_expansion(128'hd565dde95f1c2ec605a72433512094b6, {16'd46033, 16'd53725, 16'd13711, 16'd18442, 16'd34009, 16'd64524, 16'd45154, 16'd29026, 16'd57776, 16'd25048, 16'd43153, 16'd48592, 16'd37012, 16'd28305, 16'd24821, 16'd16511, 16'd18260, 16'd41039, 16'd7537, 16'd6126, 16'd6660, 16'd63111, 16'd21001, 16'd57834, 16'd20047, 16'd49316});
	test_expansion(128'h29257c2987e9803a1a69e82b251c993f, {16'd43418, 16'd55460, 16'd19136, 16'd27544, 16'd29000, 16'd5819, 16'd1369, 16'd42788, 16'd58791, 16'd3578, 16'd32014, 16'd35100, 16'd60659, 16'd44838, 16'd31864, 16'd23826, 16'd65486, 16'd22887, 16'd48773, 16'd41066, 16'd23359, 16'd56497, 16'd19844, 16'd20887, 16'd54508, 16'd42271});
	test_expansion(128'h4288b4bab1ca0a732177dff7d863f631, {16'd54758, 16'd28140, 16'd16992, 16'd64502, 16'd61416, 16'd46361, 16'd33727, 16'd57071, 16'd61888, 16'd1917, 16'd12110, 16'd16091, 16'd23020, 16'd31472, 16'd44373, 16'd2494, 16'd23108, 16'd46989, 16'd18049, 16'd19878, 16'd58661, 16'd40432, 16'd26464, 16'd43476, 16'd21751, 16'd49229});
	test_expansion(128'h08600e34db62f07c1e8863f1ebab8eb2, {16'd55773, 16'd29362, 16'd54745, 16'd13191, 16'd17267, 16'd36782, 16'd15892, 16'd62287, 16'd53542, 16'd36670, 16'd65350, 16'd20589, 16'd23983, 16'd47159, 16'd52374, 16'd37284, 16'd55457, 16'd13245, 16'd57488, 16'd2853, 16'd10650, 16'd55976, 16'd42608, 16'd59203, 16'd55034, 16'd9211});
	test_expansion(128'he9a558c66e82490efbf0bb0b49586e71, {16'd11510, 16'd9304, 16'd30258, 16'd28711, 16'd64302, 16'd51087, 16'd27771, 16'd7968, 16'd7001, 16'd58394, 16'd51623, 16'd13161, 16'd15453, 16'd56955, 16'd59230, 16'd56397, 16'd53454, 16'd3414, 16'd61211, 16'd48812, 16'd26539, 16'd27362, 16'd16418, 16'd3398, 16'd54762, 16'd42615});
	test_expansion(128'h11bef61495110d33e4620c2d0cb73a57, {16'd70, 16'd21027, 16'd18721, 16'd45346, 16'd48783, 16'd65062, 16'd45931, 16'd58269, 16'd15492, 16'd9591, 16'd46716, 16'd18409, 16'd25533, 16'd38224, 16'd64309, 16'd9451, 16'd50477, 16'd9317, 16'd55119, 16'd42411, 16'd50080, 16'd38187, 16'd15724, 16'd48649, 16'd26692, 16'd39155});
	test_expansion(128'h3bcc7d021cb18c19947919ff235366f0, {16'd63840, 16'd36640, 16'd56206, 16'd17520, 16'd41968, 16'd35389, 16'd4749, 16'd2042, 16'd55411, 16'd56606, 16'd12895, 16'd23696, 16'd6007, 16'd7939, 16'd35505, 16'd14961, 16'd43748, 16'd23116, 16'd8549, 16'd51219, 16'd18453, 16'd25912, 16'd60456, 16'd8662, 16'd36811, 16'd46666});
	test_expansion(128'h68204305bdeaf8e294b6a4f7d35b238a, {16'd46207, 16'd4565, 16'd38629, 16'd37998, 16'd1221, 16'd545, 16'd30322, 16'd25729, 16'd19804, 16'd1265, 16'd27799, 16'd37743, 16'd41364, 16'd47123, 16'd6951, 16'd19979, 16'd24726, 16'd28760, 16'd24849, 16'd37750, 16'd7122, 16'd57624, 16'd57178, 16'd20520, 16'd28406, 16'd45084});
	test_expansion(128'h8a7d93226550514ac779615fcfb7d81c, {16'd22614, 16'd61874, 16'd29542, 16'd62315, 16'd57147, 16'd199, 16'd54667, 16'd36910, 16'd23813, 16'd2482, 16'd4902, 16'd39013, 16'd62340, 16'd39584, 16'd29091, 16'd64531, 16'd32840, 16'd55311, 16'd33214, 16'd12014, 16'd59451, 16'd9547, 16'd48916, 16'd42475, 16'd44280, 16'd38277});
	test_expansion(128'h49214bd930eb3b404fc4a03c578dd6f3, {16'd17213, 16'd63722, 16'd28664, 16'd22616, 16'd38897, 16'd46531, 16'd36127, 16'd36327, 16'd34273, 16'd17940, 16'd34548, 16'd54614, 16'd47516, 16'd46855, 16'd47197, 16'd26717, 16'd22533, 16'd2986, 16'd13325, 16'd40418, 16'd52571, 16'd17158, 16'd51268, 16'd10934, 16'd44935, 16'd34204});
	test_expansion(128'h1be5e6b8a344961f5b8e1ded785d42ff, {16'd6245, 16'd34361, 16'd9896, 16'd17589, 16'd24386, 16'd1018, 16'd27866, 16'd50506, 16'd6015, 16'd50233, 16'd51995, 16'd11795, 16'd37130, 16'd38226, 16'd57686, 16'd2802, 16'd43219, 16'd750, 16'd57482, 16'd3996, 16'd47787, 16'd43573, 16'd8705, 16'd1519, 16'd53307, 16'd22367});
	test_expansion(128'hc3b3999904dc5fa98f03ceacfd6a2324, {16'd19310, 16'd65240, 16'd64328, 16'd46782, 16'd50256, 16'd32419, 16'd42817, 16'd43548, 16'd27534, 16'd49260, 16'd11471, 16'd36795, 16'd19, 16'd10596, 16'd30453, 16'd38426, 16'd59269, 16'd13015, 16'd21513, 16'd30245, 16'd34739, 16'd8938, 16'd12364, 16'd4005, 16'd15406, 16'd1514});
	test_expansion(128'h1775f2c6f0ee0f524cbeef3305509028, {16'd12274, 16'd48651, 16'd12278, 16'd48493, 16'd58901, 16'd47350, 16'd6967, 16'd26887, 16'd889, 16'd6502, 16'd10633, 16'd15951, 16'd63717, 16'd39351, 16'd47121, 16'd12055, 16'd30336, 16'd31568, 16'd26526, 16'd45981, 16'd1614, 16'd54819, 16'd56699, 16'd43401, 16'd5309, 16'd8868});
	test_expansion(128'h0ec6208be8e4ceab0c74b74db304332f, {16'd18887, 16'd13340, 16'd12230, 16'd21142, 16'd21852, 16'd58086, 16'd52241, 16'd55795, 16'd33881, 16'd3334, 16'd45676, 16'd21222, 16'd55733, 16'd13596, 16'd56595, 16'd39868, 16'd5298, 16'd37146, 16'd17997, 16'd11913, 16'd43817, 16'd2844, 16'd34095, 16'd17439, 16'd26857, 16'd49003});
	test_expansion(128'hbaf8cad7daecdc9285946607485dc314, {16'd16937, 16'd21861, 16'd4823, 16'd26521, 16'd57397, 16'd30276, 16'd46816, 16'd39018, 16'd12798, 16'd45274, 16'd53009, 16'd20147, 16'd34888, 16'd64301, 16'd43210, 16'd42349, 16'd41895, 16'd48250, 16'd12500, 16'd26341, 16'd39144, 16'd64816, 16'd33453, 16'd29957, 16'd43696, 16'd53517});
	test_expansion(128'hb209e881852369fd386c106f28ce9cba, {16'd18455, 16'd4736, 16'd2228, 16'd49779, 16'd10347, 16'd33569, 16'd39085, 16'd16477, 16'd11011, 16'd49902, 16'd61434, 16'd3575, 16'd20452, 16'd21752, 16'd33655, 16'd34627, 16'd27059, 16'd49387, 16'd32878, 16'd35326, 16'd27449, 16'd10516, 16'd61509, 16'd61977, 16'd9604, 16'd36009});
	test_expansion(128'h27d259b47e9368c40dff9f609d0123d9, {16'd59557, 16'd38724, 16'd40816, 16'd38252, 16'd2707, 16'd46023, 16'd3682, 16'd2698, 16'd42218, 16'd28725, 16'd16659, 16'd21821, 16'd10194, 16'd42002, 16'd61364, 16'd30150, 16'd15556, 16'd43308, 16'd16196, 16'd32396, 16'd47104, 16'd22477, 16'd31882, 16'd19078, 16'd22676, 16'd47327});
	test_expansion(128'h43f8c24171c6f12a84f7ad9d23b94f52, {16'd559, 16'd49465, 16'd27952, 16'd60523, 16'd37426, 16'd63299, 16'd62498, 16'd222, 16'd50418, 16'd25448, 16'd60933, 16'd24743, 16'd33999, 16'd21311, 16'd63593, 16'd54691, 16'd11733, 16'd6048, 16'd55457, 16'd57360, 16'd13434, 16'd35277, 16'd29772, 16'd6526, 16'd7317, 16'd46695});
	test_expansion(128'hcba8605b6912d0d3fbcc8489fe0848c6, {16'd63837, 16'd22144, 16'd30865, 16'd30813, 16'd64989, 16'd33872, 16'd48603, 16'd36184, 16'd44492, 16'd30952, 16'd47891, 16'd51984, 16'd34819, 16'd26780, 16'd11799, 16'd5937, 16'd32078, 16'd5058, 16'd65510, 16'd1885, 16'd6226, 16'd1187, 16'd55721, 16'd33677, 16'd39777, 16'd17746});
	test_expansion(128'h18339d2329c323c4af3075762d5a8ab3, {16'd63299, 16'd9623, 16'd17260, 16'd40313, 16'd1693, 16'd22595, 16'd48177, 16'd46348, 16'd12539, 16'd55879, 16'd20515, 16'd15094, 16'd53210, 16'd10819, 16'd21994, 16'd10053, 16'd43918, 16'd47948, 16'd25826, 16'd48513, 16'd61489, 16'd65080, 16'd12511, 16'd46241, 16'd39457, 16'd59102});
	test_expansion(128'h843691e4ff4a3106400bbb73918079ab, {16'd25793, 16'd17660, 16'd14711, 16'd41577, 16'd40047, 16'd16997, 16'd32465, 16'd33828, 16'd34695, 16'd44513, 16'd7157, 16'd55709, 16'd29403, 16'd20116, 16'd414, 16'd6956, 16'd7710, 16'd54942, 16'd64643, 16'd12731, 16'd11653, 16'd64553, 16'd43659, 16'd48241, 16'd64308, 16'd63110});
	test_expansion(128'h442d7d8f968d520b21dca94d434fe5b1, {16'd1256, 16'd35214, 16'd19657, 16'd35660, 16'd37297, 16'd51772, 16'd43294, 16'd2232, 16'd62957, 16'd4868, 16'd34065, 16'd64367, 16'd44939, 16'd42470, 16'd28490, 16'd196, 16'd18371, 16'd24671, 16'd22342, 16'd2186, 16'd39211, 16'd5996, 16'd36044, 16'd6740, 16'd16031, 16'd43018});
	test_expansion(128'h5bf38c0e1dc2069aaf194cc963155e9a, {16'd1694, 16'd35906, 16'd7152, 16'd51338, 16'd39646, 16'd52568, 16'd29214, 16'd16026, 16'd56486, 16'd36881, 16'd42430, 16'd8697, 16'd50159, 16'd5667, 16'd57457, 16'd59107, 16'd63066, 16'd64603, 16'd35661, 16'd38396, 16'd48747, 16'd4849, 16'd20682, 16'd63047, 16'd31153, 16'd31233});
	test_expansion(128'h2689fe5dc0e775e13a04c34bc5d720e6, {16'd38790, 16'd49084, 16'd8938, 16'd3572, 16'd40948, 16'd54341, 16'd27090, 16'd49778, 16'd45750, 16'd39949, 16'd13261, 16'd20118, 16'd40497, 16'd53042, 16'd6653, 16'd35239, 16'd34889, 16'd12837, 16'd4857, 16'd33737, 16'd15876, 16'd8867, 16'd39479, 16'd47899, 16'd52474, 16'd22588});
	test_expansion(128'h5b1c92f2e2a1f4ce332f901ea8fe1dbe, {16'd56426, 16'd36663, 16'd27674, 16'd5701, 16'd24602, 16'd52996, 16'd27293, 16'd36953, 16'd14168, 16'd9463, 16'd14737, 16'd6422, 16'd36161, 16'd62988, 16'd31984, 16'd32937, 16'd29668, 16'd6100, 16'd35730, 16'd40401, 16'd11884, 16'd30255, 16'd33116, 16'd11894, 16'd13367, 16'd9370});
	test_expansion(128'h818796cd758663bb92ddc1aac018bdcf, {16'd1570, 16'd7641, 16'd58311, 16'd20386, 16'd40321, 16'd43521, 16'd57715, 16'd40941, 16'd10580, 16'd5181, 16'd23477, 16'd30799, 16'd36400, 16'd5185, 16'd18671, 16'd15694, 16'd48926, 16'd28552, 16'd14677, 16'd40766, 16'd35448, 16'd18814, 16'd27872, 16'd50564, 16'd60395, 16'd8085});
	test_expansion(128'h65d2544720595643a924ad71edb2f1a2, {16'd63502, 16'd41534, 16'd23404, 16'd37334, 16'd54845, 16'd41237, 16'd20693, 16'd15657, 16'd61564, 16'd48023, 16'd48096, 16'd19170, 16'd57077, 16'd24461, 16'd17838, 16'd41561, 16'd48296, 16'd55952, 16'd33745, 16'd36680, 16'd28992, 16'd10398, 16'd36066, 16'd57820, 16'd40364, 16'd39062});
	test_expansion(128'h1d63bc3624034970043f6de7f2e4b951, {16'd44772, 16'd15344, 16'd50846, 16'd22115, 16'd22624, 16'd32482, 16'd4374, 16'd25427, 16'd8947, 16'd23796, 16'd38290, 16'd31111, 16'd62613, 16'd5822, 16'd33855, 16'd20093, 16'd23866, 16'd20672, 16'd59764, 16'd64064, 16'd22114, 16'd26902, 16'd19459, 16'd49879, 16'd59841, 16'd51579});
	test_expansion(128'h42851ce209df969dacbc27078350dea7, {16'd16462, 16'd51684, 16'd41060, 16'd25223, 16'd2098, 16'd34097, 16'd15652, 16'd54768, 16'd33852, 16'd52171, 16'd1520, 16'd46216, 16'd35263, 16'd33323, 16'd44869, 16'd18240, 16'd44710, 16'd9323, 16'd30658, 16'd33877, 16'd44756, 16'd63449, 16'd60652, 16'd24121, 16'd60258, 16'd48321});
	test_expansion(128'hea766acdf6b6cc32baa461d31ef082ec, {16'd64116, 16'd35675, 16'd52631, 16'd49520, 16'd28797, 16'd59234, 16'd40718, 16'd9825, 16'd20052, 16'd51101, 16'd5616, 16'd63652, 16'd59668, 16'd13468, 16'd14764, 16'd10147, 16'd31047, 16'd20741, 16'd14854, 16'd6256, 16'd14517, 16'd6462, 16'd12638, 16'd58923, 16'd15382, 16'd43608});
	test_expansion(128'h9074f32d9a1848c5c9abf6e7a3577169, {16'd10438, 16'd56998, 16'd53051, 16'd20838, 16'd65309, 16'd56754, 16'd63269, 16'd52282, 16'd620, 16'd23623, 16'd19261, 16'd1485, 16'd22994, 16'd9148, 16'd13293, 16'd26522, 16'd9805, 16'd41768, 16'd59108, 16'd33247, 16'd64022, 16'd34838, 16'd23628, 16'd16040, 16'd61284, 16'd22429});
	test_expansion(128'h77527fc96f207cb19b79b6c777ab68d1, {16'd58040, 16'd42751, 16'd3798, 16'd41929, 16'd41622, 16'd57902, 16'd58849, 16'd34082, 16'd16371, 16'd36399, 16'd54481, 16'd11363, 16'd4353, 16'd18822, 16'd2599, 16'd31075, 16'd48814, 16'd20154, 16'd34417, 16'd30814, 16'd64546, 16'd18368, 16'd56344, 16'd38123, 16'd49456, 16'd28716});
	test_expansion(128'hd07bda67611c1f6b250a3981248b533b, {16'd32258, 16'd31665, 16'd26108, 16'd48915, 16'd31495, 16'd8202, 16'd8933, 16'd51233, 16'd29165, 16'd15372, 16'd61890, 16'd48611, 16'd28042, 16'd57051, 16'd47854, 16'd61873, 16'd16853, 16'd6923, 16'd26238, 16'd23384, 16'd15368, 16'd40252, 16'd6273, 16'd49604, 16'd12476, 16'd43362});
	test_expansion(128'h51777a3f27d42c1f56ad9e17ad434e53, {16'd40361, 16'd25459, 16'd17088, 16'd48270, 16'd8479, 16'd50404, 16'd35505, 16'd50839, 16'd8631, 16'd7663, 16'd21148, 16'd17341, 16'd65419, 16'd54596, 16'd56858, 16'd1393, 16'd9824, 16'd9771, 16'd21124, 16'd52850, 16'd248, 16'd34281, 16'd52123, 16'd30902, 16'd20499, 16'd9680});
	test_expansion(128'h42948557b1b8dde3c7036947c6854c73, {16'd18564, 16'd63216, 16'd14450, 16'd7576, 16'd13818, 16'd35679, 16'd14429, 16'd3931, 16'd55453, 16'd26420, 16'd47963, 16'd14192, 16'd18718, 16'd16214, 16'd31515, 16'd14561, 16'd54263, 16'd53886, 16'd21243, 16'd37945, 16'd54386, 16'd17794, 16'd38047, 16'd156, 16'd40186, 16'd61531});
	test_expansion(128'hfaa449b80cb266b28709b6ddacafaa73, {16'd57984, 16'd50889, 16'd65449, 16'd42113, 16'd58823, 16'd26256, 16'd30599, 16'd48435, 16'd57311, 16'd8001, 16'd6815, 16'd53092, 16'd53026, 16'd27268, 16'd677, 16'd54693, 16'd41069, 16'd24702, 16'd8827, 16'd21921, 16'd29200, 16'd12335, 16'd16954, 16'd30069, 16'd42183, 16'd15805});
	test_expansion(128'h1c3fa4c338b4677333c8c782b0fe244c, {16'd39534, 16'd1409, 16'd6245, 16'd32202, 16'd2631, 16'd5469, 16'd6995, 16'd64803, 16'd56484, 16'd52189, 16'd48711, 16'd10069, 16'd33130, 16'd61420, 16'd22337, 16'd10341, 16'd64334, 16'd58500, 16'd49020, 16'd931, 16'd63067, 16'd5990, 16'd22929, 16'd30707, 16'd50009, 16'd3821});
	test_expansion(128'h089b0cb3ef6ab1482e860a10c692016e, {16'd35246, 16'd62470, 16'd37703, 16'd29943, 16'd39036, 16'd64706, 16'd65499, 16'd55449, 16'd6862, 16'd16007, 16'd44740, 16'd6915, 16'd65505, 16'd51520, 16'd38400, 16'd36011, 16'd54902, 16'd34142, 16'd47637, 16'd36588, 16'd40073, 16'd42166, 16'd19020, 16'd22397, 16'd42861, 16'd5690});
	test_expansion(128'he48f83b8b7a8ca426e5b616e5681c9e8, {16'd29797, 16'd47427, 16'd16416, 16'd1556, 16'd7335, 16'd46651, 16'd56316, 16'd41535, 16'd11461, 16'd26428, 16'd16031, 16'd30789, 16'd10784, 16'd2741, 16'd16060, 16'd39441, 16'd23072, 16'd61597, 16'd19089, 16'd20195, 16'd59312, 16'd52307, 16'd27960, 16'd27827, 16'd7245, 16'd675});
	test_expansion(128'hc1f65e671027aa81f444c35dbb5fa2b6, {16'd56661, 16'd48444, 16'd35888, 16'd19620, 16'd51229, 16'd27035, 16'd543, 16'd45678, 16'd10761, 16'd38744, 16'd4096, 16'd37614, 16'd40466, 16'd21745, 16'd5828, 16'd16771, 16'd63656, 16'd60686, 16'd15483, 16'd21339, 16'd51162, 16'd12924, 16'd21487, 16'd41028, 16'd3094, 16'd3169});
	test_expansion(128'h7c3bc680beab9a31f51c6b5bb66307f8, {16'd7471, 16'd65442, 16'd52556, 16'd40570, 16'd35368, 16'd48813, 16'd41088, 16'd13214, 16'd345, 16'd4708, 16'd11058, 16'd44198, 16'd30070, 16'd235, 16'd33453, 16'd63341, 16'd2978, 16'd4307, 16'd63143, 16'd7790, 16'd1336, 16'd17272, 16'd48337, 16'd14858, 16'd65041, 16'd6850});
	test_expansion(128'h865380613855eb16b351e8f4368ae05e, {16'd32116, 16'd31267, 16'd52632, 16'd37030, 16'd19345, 16'd42503, 16'd34387, 16'd2544, 16'd53677, 16'd41632, 16'd19134, 16'd46276, 16'd54641, 16'd45129, 16'd6315, 16'd44489, 16'd42305, 16'd34729, 16'd29218, 16'd31322, 16'd44077, 16'd1029, 16'd53348, 16'd35559, 16'd26947, 16'd54424});
	test_expansion(128'h31e6d98e6682d75709671836a5afe0cf, {16'd35249, 16'd6133, 16'd9947, 16'd14802, 16'd53386, 16'd1562, 16'd26151, 16'd46731, 16'd14755, 16'd27214, 16'd9177, 16'd12957, 16'd62733, 16'd7593, 16'd10818, 16'd5096, 16'd54931, 16'd18914, 16'd14939, 16'd10847, 16'd40373, 16'd28393, 16'd19423, 16'd3850, 16'd47914, 16'd55363});
	test_expansion(128'h5be5acb9ac60961c9725062b0aa80235, {16'd4672, 16'd9137, 16'd63282, 16'd31817, 16'd33243, 16'd58381, 16'd30304, 16'd32780, 16'd63957, 16'd61017, 16'd1890, 16'd54508, 16'd52270, 16'd43852, 16'd45797, 16'd43380, 16'd33372, 16'd35747, 16'd9826, 16'd40598, 16'd42989, 16'd39202, 16'd35025, 16'd47122, 16'd63837, 16'd49324});
	test_expansion(128'h22212b9b3bfb5844615ce29b6687820c, {16'd34534, 16'd32324, 16'd12933, 16'd25004, 16'd4981, 16'd50647, 16'd57600, 16'd29517, 16'd19885, 16'd62250, 16'd17896, 16'd30905, 16'd10441, 16'd60121, 16'd1857, 16'd52962, 16'd63116, 16'd33328, 16'd45933, 16'd12270, 16'd64385, 16'd13658, 16'd12191, 16'd46752, 16'd41238, 16'd6718});
	test_expansion(128'h181364d2696c30532c725c9aa8534651, {16'd52873, 16'd1067, 16'd54264, 16'd620, 16'd30981, 16'd27301, 16'd14527, 16'd64053, 16'd38088, 16'd10563, 16'd26757, 16'd27171, 16'd58679, 16'd62285, 16'd35441, 16'd30913, 16'd43450, 16'd24043, 16'd53689, 16'd19461, 16'd62163, 16'd23806, 16'd25554, 16'd49352, 16'd52677, 16'd30763});
	test_expansion(128'hb6c9ae949ade5d3e5076d1575adf23cc, {16'd41865, 16'd36925, 16'd6857, 16'd15875, 16'd37221, 16'd25765, 16'd25817, 16'd45750, 16'd24975, 16'd46804, 16'd44549, 16'd7904, 16'd1652, 16'd62564, 16'd21552, 16'd57550, 16'd4410, 16'd6344, 16'd56476, 16'd16771, 16'd46628, 16'd36526, 16'd5749, 16'd59453, 16'd54203, 16'd41699});
	test_expansion(128'ha4085c5ba6137b0c555d6973d95edc0e, {16'd3147, 16'd663, 16'd27380, 16'd7866, 16'd38358, 16'd4507, 16'd41122, 16'd13014, 16'd17811, 16'd51847, 16'd41835, 16'd40730, 16'd16429, 16'd30011, 16'd29188, 16'd54026, 16'd13179, 16'd44359, 16'd8842, 16'd30987, 16'd61481, 16'd3138, 16'd47746, 16'd38533, 16'd19771, 16'd61744});
	test_expansion(128'h2045e893f2d84a878081ba66b1096e30, {16'd54854, 16'd19822, 16'd28290, 16'd28630, 16'd30662, 16'd12255, 16'd19133, 16'd58913, 16'd28197, 16'd13713, 16'd13433, 16'd48473, 16'd31067, 16'd22208, 16'd59702, 16'd60944, 16'd10390, 16'd20816, 16'd28865, 16'd12629, 16'd61908, 16'd30380, 16'd52961, 16'd31125, 16'd47056, 16'd7678});
	test_expansion(128'h666a8ebdad6e9a6770537397b56d921f, {16'd9649, 16'd3087, 16'd62797, 16'd31546, 16'd51313, 16'd11356, 16'd18238, 16'd61813, 16'd7164, 16'd26147, 16'd60745, 16'd19470, 16'd43785, 16'd52810, 16'd32830, 16'd55487, 16'd21737, 16'd40074, 16'd61831, 16'd63783, 16'd19460, 16'd46279, 16'd16435, 16'd39049, 16'd9969, 16'd27622});
	test_expansion(128'h9f27a7ba328a644bc21211d7b46eb6bc, {16'd17896, 16'd12376, 16'd10349, 16'd52109, 16'd12248, 16'd8540, 16'd33615, 16'd2801, 16'd4212, 16'd18285, 16'd13094, 16'd51271, 16'd39360, 16'd11561, 16'd53991, 16'd61402, 16'd42933, 16'd37054, 16'd46321, 16'd19462, 16'd32129, 16'd50763, 16'd36003, 16'd46340, 16'd44278, 16'd7613});
	test_expansion(128'h3cf9ca07069e076288894bf6d9156be4, {16'd7765, 16'd58754, 16'd56428, 16'd11722, 16'd48442, 16'd55819, 16'd20151, 16'd52466, 16'd3380, 16'd32565, 16'd32683, 16'd1979, 16'd61293, 16'd20078, 16'd3903, 16'd33319, 16'd21675, 16'd31023, 16'd14585, 16'd50635, 16'd2542, 16'd25304, 16'd17145, 16'd32778, 16'd20537, 16'd29880});
	test_expansion(128'h31f676e93a292cf5b1500b159fed5316, {16'd7832, 16'd31006, 16'd38011, 16'd13383, 16'd55368, 16'd31376, 16'd4374, 16'd62064, 16'd43526, 16'd61496, 16'd38475, 16'd64091, 16'd54625, 16'd43912, 16'd1300, 16'd32941, 16'd13020, 16'd29391, 16'd51261, 16'd58581, 16'd46842, 16'd23861, 16'd40764, 16'd46883, 16'd61784, 16'd27489});
	test_expansion(128'h564b828f6db3fe8b34fb7a55aeb38116, {16'd16431, 16'd15081, 16'd27721, 16'd48222, 16'd23770, 16'd10315, 16'd36155, 16'd33254, 16'd43671, 16'd16422, 16'd37305, 16'd54129, 16'd49571, 16'd61864, 16'd18949, 16'd46211, 16'd46212, 16'd5506, 16'd54563, 16'd49759, 16'd33741, 16'd27160, 16'd25053, 16'd16669, 16'd62025, 16'd60533});
	test_expansion(128'hbb82123dba88359df836913b78951f36, {16'd44144, 16'd8737, 16'd32668, 16'd32146, 16'd40156, 16'd14438, 16'd14584, 16'd1091, 16'd24860, 16'd8572, 16'd23397, 16'd5115, 16'd42242, 16'd14675, 16'd61841, 16'd45005, 16'd10663, 16'd49776, 16'd20137, 16'd17344, 16'd10177, 16'd33987, 16'd49217, 16'd10630, 16'd12561, 16'd17937});
	test_expansion(128'ha8a19b73126ead6cfa0940f669b74636, {16'd13034, 16'd48035, 16'd16484, 16'd22313, 16'd60262, 16'd12193, 16'd34759, 16'd60222, 16'd23400, 16'd19261, 16'd3584, 16'd24164, 16'd31229, 16'd28965, 16'd46923, 16'd56670, 16'd35136, 16'd61263, 16'd53995, 16'd61537, 16'd11537, 16'd16990, 16'd25716, 16'd40139, 16'd55695, 16'd6569});
	test_expansion(128'h92cb48d0ade9c8d5159df3825a5dcd28, {16'd46396, 16'd504, 16'd50853, 16'd44337, 16'd43644, 16'd29632, 16'd39014, 16'd43078, 16'd6379, 16'd58998, 16'd39021, 16'd53506, 16'd18246, 16'd657, 16'd25908, 16'd2559, 16'd42381, 16'd38628, 16'd10879, 16'd23070, 16'd5842, 16'd5643, 16'd32633, 16'd1284, 16'd1807, 16'd49085});
	test_expansion(128'hef9359c5f64045ebbef54550621176a5, {16'd27158, 16'd42875, 16'd39774, 16'd61013, 16'd43002, 16'd47371, 16'd16215, 16'd33970, 16'd63938, 16'd55780, 16'd44767, 16'd50308, 16'd4175, 16'd28755, 16'd17930, 16'd34725, 16'd56034, 16'd29246, 16'd35274, 16'd11798, 16'd9653, 16'd65288, 16'd10380, 16'd10718, 16'd19813, 16'd50213});
	test_expansion(128'h315783f9db121f3ce54fd7b6c64a2331, {16'd38119, 16'd34665, 16'd25175, 16'd22539, 16'd35631, 16'd18472, 16'd30319, 16'd29119, 16'd2097, 16'd6054, 16'd31021, 16'd24448, 16'd27251, 16'd53997, 16'd54693, 16'd33401, 16'd6588, 16'd36983, 16'd20189, 16'd8233, 16'd54722, 16'd15340, 16'd63017, 16'd60257, 16'd41999, 16'd22156});
	test_expansion(128'h40c74c2bbe34789638bd7daa7de56d2b, {16'd3443, 16'd14669, 16'd13696, 16'd63900, 16'd48387, 16'd18465, 16'd41827, 16'd35353, 16'd25754, 16'd31448, 16'd61083, 16'd40352, 16'd13494, 16'd47350, 16'd27576, 16'd58819, 16'd57620, 16'd46784, 16'd8754, 16'd36891, 16'd22980, 16'd1756, 16'd17264, 16'd22974, 16'd34586, 16'd51949});
	test_expansion(128'hd0c6c17d9b66f5a884418719255a1134, {16'd35433, 16'd58635, 16'd2855, 16'd41342, 16'd26533, 16'd35844, 16'd4324, 16'd47275, 16'd32200, 16'd31906, 16'd32092, 16'd31731, 16'd33300, 16'd38776, 16'd29588, 16'd23861, 16'd33147, 16'd34843, 16'd26995, 16'd7799, 16'd31216, 16'd35468, 16'd18404, 16'd17746, 16'd40580, 16'd62206});
	test_expansion(128'he39e6dd98bd8a5f9f9bb5717c82ae167, {16'd33557, 16'd22921, 16'd23814, 16'd11104, 16'd46612, 16'd44210, 16'd9261, 16'd23374, 16'd49507, 16'd11028, 16'd43842, 16'd2924, 16'd44219, 16'd65004, 16'd60024, 16'd58636, 16'd37969, 16'd20247, 16'd46801, 16'd60148, 16'd49580, 16'd11728, 16'd16281, 16'd52373, 16'd58551, 16'd53431});
	test_expansion(128'h75f19337fc916ea5fe935922bc8473ba, {16'd1428, 16'd35169, 16'd63519, 16'd47117, 16'd46235, 16'd22683, 16'd43665, 16'd5507, 16'd12563, 16'd18491, 16'd41080, 16'd63858, 16'd17138, 16'd57161, 16'd27271, 16'd12839, 16'd63599, 16'd36851, 16'd55241, 16'd15261, 16'd13079, 16'd65302, 16'd47243, 16'd52807, 16'd56178, 16'd9377});
	test_expansion(128'hf6add0071f0208acc392eca4c590a0d7, {16'd16065, 16'd53001, 16'd58898, 16'd20596, 16'd41381, 16'd13566, 16'd39063, 16'd22082, 16'd55931, 16'd1021, 16'd13589, 16'd8736, 16'd27190, 16'd29653, 16'd49231, 16'd21237, 16'd48052, 16'd47962, 16'd37391, 16'd55002, 16'd46190, 16'd337, 16'd44146, 16'd37754, 16'd17345, 16'd56552});
	test_expansion(128'h361f8d1a495a8ac31b65057a29bd1e9c, {16'd17983, 16'd8647, 16'd10659, 16'd64205, 16'd64251, 16'd55131, 16'd26967, 16'd45310, 16'd3722, 16'd58858, 16'd45769, 16'd14443, 16'd63811, 16'd46594, 16'd48945, 16'd4025, 16'd61306, 16'd45887, 16'd54178, 16'd11698, 16'd61260, 16'd391, 16'd36396, 16'd43350, 16'd14388, 16'd62590});
	test_expansion(128'h708f0baeaef874aeeb8f6756becd7f79, {16'd696, 16'd39804, 16'd56337, 16'd38045, 16'd64737, 16'd14702, 16'd888, 16'd36607, 16'd40732, 16'd4367, 16'd29047, 16'd47285, 16'd53125, 16'd42814, 16'd47002, 16'd14429, 16'd14518, 16'd56288, 16'd3611, 16'd60519, 16'd23898, 16'd5117, 16'd64799, 16'd61544, 16'd40545, 16'd48740});
	test_expansion(128'ha1f279901c2f8e8572d5cf9d9b18a415, {16'd17192, 16'd18224, 16'd9857, 16'd61666, 16'd49301, 16'd29987, 16'd47498, 16'd19032, 16'd7245, 16'd2499, 16'd47176, 16'd54007, 16'd40218, 16'd47225, 16'd35721, 16'd9585, 16'd30852, 16'd29855, 16'd32429, 16'd40070, 16'd38060, 16'd19778, 16'd59854, 16'd24837, 16'd4726, 16'd30615});
	test_expansion(128'h3660608ff3136240a95db857c18e999b, {16'd39616, 16'd24625, 16'd31409, 16'd57781, 16'd51529, 16'd60821, 16'd14544, 16'd36023, 16'd59574, 16'd38912, 16'd16795, 16'd57287, 16'd28917, 16'd32919, 16'd53071, 16'd47522, 16'd18885, 16'd58068, 16'd39613, 16'd79, 16'd12989, 16'd43108, 16'd5236, 16'd62446, 16'd61033, 16'd21031});
	test_expansion(128'hc39e73cceae4e7a83ef59679ba9b56b7, {16'd7595, 16'd30443, 16'd62510, 16'd33858, 16'd5486, 16'd3042, 16'd8188, 16'd27234, 16'd64750, 16'd32701, 16'd35074, 16'd20618, 16'd34647, 16'd56197, 16'd14552, 16'd21290, 16'd12867, 16'd12475, 16'd57867, 16'd23949, 16'd27390, 16'd43539, 16'd47755, 16'd62116, 16'd54553, 16'd23822});
	test_expansion(128'h2394c8b89a14ccb656789275f7a0e715, {16'd61866, 16'd12397, 16'd29132, 16'd60079, 16'd12750, 16'd57408, 16'd21762, 16'd36196, 16'd8878, 16'd29550, 16'd34351, 16'd56344, 16'd51103, 16'd4054, 16'd13867, 16'd22945, 16'd48922, 16'd49434, 16'd37997, 16'd61964, 16'd24392, 16'd34357, 16'd44804, 16'd15948, 16'd61054, 16'd8777});
	test_expansion(128'h8d2c7b2d8d1a06a4612503e269e4036a, {16'd22913, 16'd59416, 16'd43540, 16'd61614, 16'd1176, 16'd54251, 16'd15476, 16'd43257, 16'd27586, 16'd18470, 16'd64404, 16'd23345, 16'd20324, 16'd2729, 16'd6968, 16'd48101, 16'd5265, 16'd19953, 16'd62195, 16'd184, 16'd16787, 16'd38063, 16'd46817, 16'd25709, 16'd55820, 16'd63065});
	test_expansion(128'hb7244477f882204fa3b0a6ab6ef3fda3, {16'd53553, 16'd8481, 16'd2139, 16'd41545, 16'd10351, 16'd5361, 16'd54273, 16'd19536, 16'd1869, 16'd4682, 16'd5471, 16'd58048, 16'd12565, 16'd9539, 16'd27139, 16'd7570, 16'd11189, 16'd24336, 16'd38307, 16'd55711, 16'd35273, 16'd54645, 16'd59944, 16'd52650, 16'd37042, 16'd49866});
	test_expansion(128'hba8c8b7ceec34d58eb84204fa95578c7, {16'd17644, 16'd10851, 16'd23443, 16'd39829, 16'd57917, 16'd41072, 16'd45867, 16'd59027, 16'd64305, 16'd43146, 16'd42350, 16'd12309, 16'd21416, 16'd17209, 16'd36696, 16'd3483, 16'd33703, 16'd64224, 16'd38667, 16'd4162, 16'd8081, 16'd47889, 16'd64451, 16'd33998, 16'd57381, 16'd4246});
	test_expansion(128'h0e902858e6ef95bda30588ba68d42e03, {16'd8601, 16'd57390, 16'd30477, 16'd59781, 16'd40155, 16'd61968, 16'd38487, 16'd40696, 16'd40661, 16'd7746, 16'd26087, 16'd24511, 16'd51882, 16'd27360, 16'd63533, 16'd44681, 16'd55275, 16'd55140, 16'd13296, 16'd63046, 16'd52637, 16'd24850, 16'd7927, 16'd41428, 16'd38707, 16'd55584});
	test_expansion(128'hebff2fbcee9f0e005c8ca5aa0ae9b0db, {16'd60586, 16'd47913, 16'd63122, 16'd3740, 16'd9842, 16'd30226, 16'd28182, 16'd20738, 16'd23501, 16'd7850, 16'd55031, 16'd29752, 16'd56121, 16'd59415, 16'd28351, 16'd55330, 16'd61083, 16'd60270, 16'd4188, 16'd272, 16'd43507, 16'd3578, 16'd43301, 16'd21505, 16'd6081, 16'd62026});
	test_expansion(128'hf9993070ecb98b558761718c31c99c34, {16'd10895, 16'd65406, 16'd48816, 16'd56674, 16'd50741, 16'd13263, 16'd20743, 16'd4924, 16'd627, 16'd42696, 16'd9314, 16'd1199, 16'd60717, 16'd19268, 16'd60643, 16'd14025, 16'd702, 16'd55592, 16'd29901, 16'd10082, 16'd25560, 16'd52602, 16'd28117, 16'd30558, 16'd64318, 16'd46124});
	test_expansion(128'h5deacbd5bc3dca9ca9f6d86fff08341c, {16'd51077, 16'd44838, 16'd25451, 16'd39120, 16'd30490, 16'd50188, 16'd27286, 16'd47951, 16'd11809, 16'd28859, 16'd36470, 16'd41685, 16'd54673, 16'd55376, 16'd36844, 16'd62964, 16'd39823, 16'd38539, 16'd45229, 16'd10143, 16'd14889, 16'd51753, 16'd53741, 16'd1141, 16'd1450, 16'd8743});
	test_expansion(128'h7f5bf86eb5fa1bbd15f10c3c9d9b0301, {16'd47964, 16'd35685, 16'd57474, 16'd18433, 16'd22488, 16'd64877, 16'd10165, 16'd24965, 16'd62643, 16'd21441, 16'd27184, 16'd40615, 16'd8736, 16'd18080, 16'd52780, 16'd48726, 16'd40499, 16'd7416, 16'd48347, 16'd53688, 16'd23696, 16'd19730, 16'd47530, 16'd26572, 16'd20184, 16'd13572});
	test_expansion(128'h8606c6059f4d3b4baa4c4ec2e2eb92ca, {16'd26273, 16'd44245, 16'd12860, 16'd3981, 16'd1141, 16'd28537, 16'd56440, 16'd50508, 16'd58827, 16'd45961, 16'd56861, 16'd26955, 16'd30639, 16'd12849, 16'd4345, 16'd39446, 16'd64672, 16'd18160, 16'd21347, 16'd33548, 16'd57899, 16'd52401, 16'd33336, 16'd53329, 16'd57354, 16'd50003});
	test_expansion(128'h451d6247b15b3f7f7e094b5a22c158b1, {16'd30140, 16'd9996, 16'd12639, 16'd63976, 16'd35730, 16'd23753, 16'd4533, 16'd42260, 16'd6175, 16'd46113, 16'd50537, 16'd4942, 16'd42363, 16'd54447, 16'd11754, 16'd26444, 16'd53661, 16'd48685, 16'd17812, 16'd29293, 16'd44709, 16'd43132, 16'd11159, 16'd36747, 16'd25610, 16'd50879});
	test_expansion(128'h3b5916ca68d482002698cda5f4472d9e, {16'd15523, 16'd32332, 16'd33035, 16'd20375, 16'd33088, 16'd34880, 16'd23369, 16'd51876, 16'd60815, 16'd22491, 16'd18752, 16'd33426, 16'd16907, 16'd3592, 16'd18734, 16'd1382, 16'd10052, 16'd24742, 16'd42715, 16'd58981, 16'd16692, 16'd34518, 16'd55243, 16'd21310, 16'd42370, 16'd52754});
	test_expansion(128'hc8c967758a9bae14bc1c2cfd06a629c5, {16'd57683, 16'd44541, 16'd31303, 16'd15686, 16'd51382, 16'd7841, 16'd54338, 16'd39277, 16'd49138, 16'd28988, 16'd35995, 16'd49986, 16'd59531, 16'd2972, 16'd32401, 16'd56923, 16'd40827, 16'd30144, 16'd14072, 16'd64873, 16'd35738, 16'd17872, 16'd25669, 16'd4539, 16'd45563, 16'd45277});
	test_expansion(128'hb205628ed5308b690e0e9099dd0aba1f, {16'd33732, 16'd38179, 16'd49839, 16'd61828, 16'd41755, 16'd14655, 16'd38947, 16'd63577, 16'd4552, 16'd34951, 16'd51214, 16'd28300, 16'd45998, 16'd56332, 16'd4175, 16'd48442, 16'd28561, 16'd47478, 16'd65114, 16'd22028, 16'd57727, 16'd64953, 16'd47083, 16'd26954, 16'd19779, 16'd33538});
	test_expansion(128'hac0667099d5ad87312b380bf3ff56f55, {16'd46385, 16'd36105, 16'd12571, 16'd42461, 16'd17566, 16'd1715, 16'd835, 16'd55260, 16'd45554, 16'd19231, 16'd19709, 16'd41732, 16'd56397, 16'd19732, 16'd31272, 16'd56979, 16'd1757, 16'd7953, 16'd53707, 16'd57010, 16'd46394, 16'd18355, 16'd52713, 16'd20019, 16'd36670, 16'd2831});
	test_expansion(128'hc18888686974526cdc5c2fb4136e2580, {16'd44137, 16'd22452, 16'd39100, 16'd40748, 16'd30752, 16'd19231, 16'd1765, 16'd64315, 16'd30076, 16'd21219, 16'd16646, 16'd31437, 16'd33294, 16'd13735, 16'd41127, 16'd60411, 16'd46219, 16'd32135, 16'd18868, 16'd37431, 16'd12198, 16'd17766, 16'd15433, 16'd17157, 16'd42783, 16'd11582});
	test_expansion(128'h98401371d6235cd6db8978d00069a970, {16'd13570, 16'd14047, 16'd1428, 16'd35711, 16'd30306, 16'd62026, 16'd21298, 16'd30037, 16'd4998, 16'd39340, 16'd16215, 16'd3927, 16'd42957, 16'd42553, 16'd38926, 16'd8001, 16'd42935, 16'd36158, 16'd17114, 16'd13627, 16'd16846, 16'd30628, 16'd39196, 16'd23535, 16'd56337, 16'd38397});
	test_expansion(128'hdd8a119c2c01481c7d4d4ccc912668db, {16'd43756, 16'd23610, 16'd49155, 16'd36851, 16'd57933, 16'd46693, 16'd20431, 16'd16607, 16'd18927, 16'd30530, 16'd36661, 16'd37264, 16'd1512, 16'd64814, 16'd61687, 16'd8965, 16'd29721, 16'd54694, 16'd35464, 16'd23827, 16'd3367, 16'd33987, 16'd59889, 16'd50879, 16'd13005, 16'd46058});
	test_expansion(128'h9e71f82bc6b5ff8e3ea2d94adb427713, {16'd39820, 16'd5598, 16'd21054, 16'd42910, 16'd45251, 16'd19568, 16'd45255, 16'd36705, 16'd36847, 16'd25570, 16'd8796, 16'd20155, 16'd36577, 16'd55937, 16'd8105, 16'd51319, 16'd23967, 16'd59958, 16'd36159, 16'd57355, 16'd27206, 16'd64862, 16'd14906, 16'd25265, 16'd22448, 16'd49884});
	test_expansion(128'hfbe003883cf765e1f27767b027e6d1ec, {16'd59269, 16'd17361, 16'd20556, 16'd52618, 16'd52587, 16'd27107, 16'd18511, 16'd48023, 16'd4502, 16'd64088, 16'd57777, 16'd63905, 16'd51607, 16'd52559, 16'd33226, 16'd9052, 16'd57892, 16'd63921, 16'd660, 16'd25223, 16'd61450, 16'd24731, 16'd18762, 16'd31877, 16'd50809, 16'd19145});
	test_expansion(128'h99936718fba656bd3c3e0285a5d9bbe1, {16'd29579, 16'd15669, 16'd41414, 16'd51623, 16'd54932, 16'd15352, 16'd44390, 16'd56345, 16'd38013, 16'd62660, 16'd24858, 16'd44754, 16'd35207, 16'd43518, 16'd39861, 16'd58054, 16'd12355, 16'd8375, 16'd64880, 16'd30718, 16'd10036, 16'd64935, 16'd48286, 16'd61911, 16'd14550, 16'd6561});
	test_expansion(128'h0b64ad03cce39099a08bedbfeb174fa3, {16'd24065, 16'd7241, 16'd34165, 16'd9170, 16'd4246, 16'd63862, 16'd41955, 16'd15554, 16'd2200, 16'd39341, 16'd37324, 16'd53669, 16'd14305, 16'd39169, 16'd5221, 16'd16001, 16'd61982, 16'd49255, 16'd26152, 16'd27692, 16'd41053, 16'd41488, 16'd54415, 16'd14447, 16'd47509, 16'd21382});
	test_expansion(128'he1e2e6baddd8393cba28208c3642be24, {16'd24730, 16'd35337, 16'd62844, 16'd17112, 16'd31273, 16'd25253, 16'd32700, 16'd12192, 16'd23998, 16'd23509, 16'd24634, 16'd9298, 16'd65157, 16'd14518, 16'd31954, 16'd56590, 16'd57574, 16'd46290, 16'd12208, 16'd23047, 16'd61818, 16'd63096, 16'd17074, 16'd30813, 16'd48209, 16'd48590});
	test_expansion(128'h0af1fa7d8dc49fd3aa38329c24bd479b, {16'd44229, 16'd37924, 16'd28016, 16'd35848, 16'd64689, 16'd31921, 16'd51543, 16'd59175, 16'd17536, 16'd31809, 16'd25146, 16'd15281, 16'd19170, 16'd58578, 16'd43808, 16'd60267, 16'd40585, 16'd64600, 16'd59101, 16'd5921, 16'd63126, 16'd47637, 16'd30889, 16'd20288, 16'd44326, 16'd49592});
	test_expansion(128'hc1a4a5a4b4f9c2745716b6096d27a369, {16'd49275, 16'd9084, 16'd7218, 16'd4818, 16'd54356, 16'd4176, 16'd43530, 16'd26239, 16'd8012, 16'd28531, 16'd56736, 16'd49074, 16'd17939, 16'd57586, 16'd15053, 16'd26689, 16'd33358, 16'd22172, 16'd15917, 16'd60808, 16'd54337, 16'd29925, 16'd35464, 16'd53262, 16'd58453, 16'd13086});
	test_expansion(128'hd6ede31747278b6af5dc92fc0c97b577, {16'd29786, 16'd17215, 16'd27352, 16'd983, 16'd44488, 16'd36432, 16'd35216, 16'd3001, 16'd27183, 16'd47880, 16'd52878, 16'd26735, 16'd17472, 16'd23255, 16'd55591, 16'd23375, 16'd36706, 16'd49302, 16'd61623, 16'd4798, 16'd39193, 16'd8392, 16'd11695, 16'd33688, 16'd16374, 16'd58046});
	test_expansion(128'h5d8db4a6ffa440d3416e97a21b8e5b36, {16'd45938, 16'd12867, 16'd53272, 16'd61672, 16'd22984, 16'd6348, 16'd59154, 16'd23857, 16'd59216, 16'd26622, 16'd32564, 16'd28339, 16'd7904, 16'd17870, 16'd53412, 16'd9449, 16'd43719, 16'd15013, 16'd63019, 16'd19993, 16'd50830, 16'd49309, 16'd48870, 16'd64190, 16'd41630, 16'd59576});
	test_expansion(128'h9cfcd6e9e5fab2a175fce36053060c8e, {16'd42260, 16'd49468, 16'd45433, 16'd18521, 16'd26199, 16'd44430, 16'd10851, 16'd20787, 16'd47991, 16'd31297, 16'd30218, 16'd9050, 16'd65174, 16'd13716, 16'd12973, 16'd57030, 16'd38685, 16'd53251, 16'd20100, 16'd11334, 16'd40400, 16'd58551, 16'd57011, 16'd58010, 16'd26878, 16'd50329});
	test_expansion(128'h6cb03346901730f6257b02fe58a4e149, {16'd6605, 16'd32340, 16'd41553, 16'd42571, 16'd37865, 16'd37217, 16'd3543, 16'd12522, 16'd63498, 16'd47463, 16'd12361, 16'd62934, 16'd26316, 16'd40874, 16'd53225, 16'd18802, 16'd64756, 16'd48224, 16'd7040, 16'd57319, 16'd54412, 16'd63203, 16'd48199, 16'd46829, 16'd8856, 16'd436});
	test_expansion(128'h12667f7eec1c9a9b7e637041b88723a2, {16'd58417, 16'd56281, 16'd14976, 16'd10044, 16'd45056, 16'd64710, 16'd43009, 16'd48221, 16'd21433, 16'd46270, 16'd12202, 16'd48979, 16'd1483, 16'd20840, 16'd3716, 16'd7446, 16'd19856, 16'd22553, 16'd12055, 16'd10797, 16'd64054, 16'd54337, 16'd42031, 16'd17471, 16'd11990, 16'd17769});
	test_expansion(128'ha3e8c58dbf7af2a970518dc848cf25d5, {16'd54343, 16'd8865, 16'd60073, 16'd65303, 16'd38336, 16'd4575, 16'd59911, 16'd48574, 16'd38106, 16'd62146, 16'd48289, 16'd7789, 16'd41133, 16'd23158, 16'd57527, 16'd40077, 16'd57316, 16'd30496, 16'd8136, 16'd54718, 16'd4519, 16'd23665, 16'd26088, 16'd43462, 16'd39430, 16'd51549});
	test_expansion(128'hf3e9a1e68ab5a93e8d5b616bfe541877, {16'd59595, 16'd59043, 16'd31472, 16'd2597, 16'd59545, 16'd36362, 16'd30169, 16'd63912, 16'd52188, 16'd3593, 16'd54562, 16'd63352, 16'd181, 16'd64773, 16'd50944, 16'd11763, 16'd58291, 16'd64518, 16'd49973, 16'd36753, 16'd35300, 16'd41701, 16'd64718, 16'd7449, 16'd19013, 16'd31918});
	test_expansion(128'h732f8d1fcc187290630032bd8d7a8277, {16'd7255, 16'd52053, 16'd31277, 16'd4745, 16'd7578, 16'd43018, 16'd38040, 16'd48532, 16'd19874, 16'd35373, 16'd16227, 16'd21494, 16'd19497, 16'd54468, 16'd27253, 16'd61493, 16'd57491, 16'd6742, 16'd39656, 16'd19903, 16'd36826, 16'd63379, 16'd38549, 16'd48877, 16'd748, 16'd31219});
	test_expansion(128'he0b8e2a4e65970332632a80109393629, {16'd56735, 16'd48963, 16'd14215, 16'd35095, 16'd42292, 16'd61777, 16'd35565, 16'd64717, 16'd23548, 16'd22013, 16'd29423, 16'd42176, 16'd13945, 16'd23538, 16'd22513, 16'd50294, 16'd3401, 16'd30334, 16'd61502, 16'd19698, 16'd5817, 16'd3034, 16'd2915, 16'd53741, 16'd64091, 16'd3337});
	test_expansion(128'h600145cc512bf2b981a7c43c52ddffdd, {16'd26959, 16'd5029, 16'd3303, 16'd1474, 16'd20364, 16'd40711, 16'd38553, 16'd63183, 16'd44453, 16'd65122, 16'd33930, 16'd65421, 16'd42495, 16'd40007, 16'd52995, 16'd23091, 16'd32228, 16'd39897, 16'd52015, 16'd34503, 16'd25823, 16'd46042, 16'd16156, 16'd12883, 16'd64007, 16'd39525});
	test_expansion(128'h74c60f32c1f37d2e29afa70850a10dae, {16'd25239, 16'd13315, 16'd37823, 16'd51670, 16'd57429, 16'd55859, 16'd5851, 16'd55792, 16'd15807, 16'd15654, 16'd49455, 16'd63649, 16'd18416, 16'd30107, 16'd37259, 16'd34261, 16'd18835, 16'd21717, 16'd12568, 16'd15524, 16'd39820, 16'd4154, 16'd36262, 16'd2423, 16'd29259, 16'd17075});
	test_expansion(128'had5414c47d5d32915142ef982fb50590, {16'd25461, 16'd6182, 16'd49698, 16'd31170, 16'd60970, 16'd23996, 16'd24355, 16'd45553, 16'd44354, 16'd63741, 16'd32066, 16'd19967, 16'd4425, 16'd19811, 16'd48681, 16'd13178, 16'd43803, 16'd9531, 16'd52344, 16'd52981, 16'd18381, 16'd31566, 16'd37370, 16'd37491, 16'd64721, 16'd52403});
	test_expansion(128'h8a78019aa8d3988a34e00bc421209fd7, {16'd39740, 16'd15003, 16'd54911, 16'd24765, 16'd18607, 16'd5232, 16'd62000, 16'd9852, 16'd32290, 16'd53799, 16'd1575, 16'd637, 16'd55757, 16'd38079, 16'd10286, 16'd59984, 16'd37253, 16'd19228, 16'd1321, 16'd4091, 16'd52449, 16'd54089, 16'd6350, 16'd63235, 16'd26979, 16'd56411});
	test_expansion(128'h405887a8a8a81d261c8312121e2cf032, {16'd48810, 16'd22356, 16'd49227, 16'd11425, 16'd15962, 16'd17163, 16'd51481, 16'd42644, 16'd44924, 16'd43877, 16'd35271, 16'd6523, 16'd26691, 16'd14282, 16'd17067, 16'd54214, 16'd50845, 16'd20063, 16'd60938, 16'd33350, 16'd15785, 16'd26560, 16'd47186, 16'd7046, 16'd49351, 16'd18802});
	test_expansion(128'h8a5bbea82b9fb077515c99ae6b75484e, {16'd50812, 16'd36990, 16'd36165, 16'd45594, 16'd26043, 16'd11086, 16'd63433, 16'd10550, 16'd54870, 16'd9516, 16'd55652, 16'd9077, 16'd42549, 16'd133, 16'd44346, 16'd30233, 16'd36349, 16'd51869, 16'd18307, 16'd62863, 16'd3288, 16'd58786, 16'd36768, 16'd33892, 16'd63928, 16'd28686});
	test_expansion(128'h8997b94130866e3c9fdee1644d6780df, {16'd30769, 16'd3447, 16'd40797, 16'd29106, 16'd26642, 16'd32139, 16'd57778, 16'd48336, 16'd19710, 16'd5911, 16'd49149, 16'd52677, 16'd1442, 16'd16941, 16'd45249, 16'd62277, 16'd36787, 16'd1320, 16'd33941, 16'd28694, 16'd10644, 16'd55941, 16'd27797, 16'd31775, 16'd43937, 16'd44018});
	test_expansion(128'hdb43506a53d5663118700638ce4e6c50, {16'd60057, 16'd12552, 16'd48693, 16'd18117, 16'd52256, 16'd20619, 16'd10153, 16'd4140, 16'd28877, 16'd39917, 16'd7707, 16'd40434, 16'd42460, 16'd6716, 16'd22639, 16'd41367, 16'd18809, 16'd45653, 16'd59488, 16'd37325, 16'd27929, 16'd23767, 16'd38284, 16'd573, 16'd52143, 16'd14641});
	test_expansion(128'h028b8063c31564e805052d031cd67af6, {16'd1290, 16'd32842, 16'd52965, 16'd45448, 16'd9731, 16'd22953, 16'd12293, 16'd12392, 16'd21962, 16'd59728, 16'd9055, 16'd18578, 16'd46533, 16'd33277, 16'd44100, 16'd44874, 16'd28478, 16'd7074, 16'd31703, 16'd32782, 16'd63947, 16'd59792, 16'd41857, 16'd4578, 16'd35506, 16'd37116});
	test_expansion(128'hb9838efdd411ac50d79390dd4164a334, {16'd10627, 16'd20958, 16'd41671, 16'd4609, 16'd64548, 16'd4014, 16'd6269, 16'd38221, 16'd12588, 16'd17647, 16'd36207, 16'd28433, 16'd46021, 16'd29221, 16'd38483, 16'd29435, 16'd60550, 16'd7514, 16'd43563, 16'd49904, 16'd25846, 16'd61255, 16'd14671, 16'd50597, 16'd8011, 16'd31225});
	test_expansion(128'h0dea5994c105d694010229c0ac72458a, {16'd28532, 16'd44906, 16'd4249, 16'd43484, 16'd6973, 16'd22985, 16'd47194, 16'd3160, 16'd14167, 16'd55525, 16'd59771, 16'd39526, 16'd56713, 16'd43270, 16'd25886, 16'd8367, 16'd8285, 16'd49404, 16'd46479, 16'd42330, 16'd56462, 16'd55489, 16'd11648, 16'd24744, 16'd59612, 16'd50474});
	test_expansion(128'h37d6a696c80442f02421ef96894a0324, {16'd42393, 16'd33600, 16'd46299, 16'd15673, 16'd11672, 16'd64870, 16'd55094, 16'd60263, 16'd38893, 16'd4386, 16'd30598, 16'd965, 16'd45702, 16'd64222, 16'd64851, 16'd46563, 16'd36858, 16'd16520, 16'd46952, 16'd167, 16'd58694, 16'd32124, 16'd55951, 16'd47353, 16'd11599, 16'd26611});
	test_expansion(128'h4844cc4e313eec1f68eae0330ab9134a, {16'd60162, 16'd47448, 16'd10764, 16'd37216, 16'd47126, 16'd30608, 16'd43580, 16'd35422, 16'd19104, 16'd27552, 16'd56589, 16'd8736, 16'd12586, 16'd37265, 16'd5738, 16'd34328, 16'd61390, 16'd47758, 16'd63777, 16'd39931, 16'd26875, 16'd23100, 16'd42205, 16'd26383, 16'd35248, 16'd63688});
	test_expansion(128'hd4d9a46d992466e03a9b6e1fd7f0d293, {16'd25276, 16'd56987, 16'd6967, 16'd52039, 16'd5904, 16'd27191, 16'd47670, 16'd30217, 16'd34305, 16'd15573, 16'd62474, 16'd38231, 16'd8888, 16'd62754, 16'd20745, 16'd3625, 16'd21767, 16'd31043, 16'd39344, 16'd2468, 16'd5262, 16'd42044, 16'd26225, 16'd21167, 16'd11329, 16'd27272});
	test_expansion(128'h05bd2291fbe9a5e9023333aaa907120c, {16'd20343, 16'd63261, 16'd27591, 16'd26540, 16'd8166, 16'd18331, 16'd17791, 16'd62963, 16'd47289, 16'd52001, 16'd29852, 16'd50857, 16'd19592, 16'd60183, 16'd59562, 16'd60396, 16'd16506, 16'd19558, 16'd5072, 16'd53804, 16'd9354, 16'd60243, 16'd40807, 16'd33291, 16'd7580, 16'd47050});
	test_expansion(128'h6aa4d5b0b199a5d57e581cff3bb1f813, {16'd30500, 16'd58283, 16'd4471, 16'd39674, 16'd12428, 16'd59465, 16'd40304, 16'd18506, 16'd5211, 16'd59067, 16'd18742, 16'd59579, 16'd17377, 16'd53061, 16'd12554, 16'd5259, 16'd56661, 16'd17168, 16'd24624, 16'd17281, 16'd2550, 16'd62838, 16'd60735, 16'd45707, 16'd11637, 16'd49882});
	test_expansion(128'hcee0650a74720dd4d6858a9abc82dead, {16'd60242, 16'd6997, 16'd36226, 16'd35868, 16'd48752, 16'd52878, 16'd60910, 16'd64655, 16'd18366, 16'd56722, 16'd57769, 16'd42081, 16'd30915, 16'd51504, 16'd26912, 16'd38320, 16'd62051, 16'd57784, 16'd21141, 16'd21776, 16'd21870, 16'd17486, 16'd6828, 16'd45260, 16'd39015, 16'd15986});
	test_expansion(128'ha1072d76f9b63cf5caff78091739dbb2, {16'd373, 16'd22289, 16'd17534, 16'd42091, 16'd40893, 16'd51361, 16'd3231, 16'd50389, 16'd10082, 16'd3889, 16'd11191, 16'd44127, 16'd19115, 16'd31283, 16'd9399, 16'd7660, 16'd53346, 16'd22386, 16'd5561, 16'd38833, 16'd47210, 16'd13252, 16'd42594, 16'd10911, 16'd14575, 16'd64292});
	test_expansion(128'he4fcd63e76f42ad923ef0bfae2e3434b, {16'd18580, 16'd27169, 16'd62473, 16'd34944, 16'd55794, 16'd19021, 16'd6735, 16'd5344, 16'd41353, 16'd48082, 16'd41737, 16'd27633, 16'd28175, 16'd18887, 16'd4478, 16'd43670, 16'd46697, 16'd44818, 16'd56602, 16'd42228, 16'd3692, 16'd3021, 16'd50927, 16'd11753, 16'd23633, 16'd62750});
	test_expansion(128'hf8616c1d0650a18b9ae2f780a643face, {16'd28341, 16'd46791, 16'd64823, 16'd47999, 16'd5593, 16'd65052, 16'd27123, 16'd7430, 16'd27080, 16'd2754, 16'd19027, 16'd61768, 16'd38679, 16'd46924, 16'd56561, 16'd13339, 16'd20891, 16'd48488, 16'd16177, 16'd47297, 16'd31902, 16'd46684, 16'd17073, 16'd25152, 16'd37656, 16'd3426});
	test_expansion(128'h227ca16be7a3e1715913a271475d5b00, {16'd6015, 16'd32180, 16'd46242, 16'd1642, 16'd14118, 16'd1463, 16'd56929, 16'd13984, 16'd25668, 16'd43577, 16'd25484, 16'd28324, 16'd28930, 16'd28337, 16'd23033, 16'd64386, 16'd58289, 16'd25678, 16'd55946, 16'd34554, 16'd30613, 16'd57332, 16'd18154, 16'd24183, 16'd41756, 16'd59915});
	test_expansion(128'h063c48b761f0f33412257f4426e70354, {16'd26000, 16'd23010, 16'd16172, 16'd19114, 16'd53189, 16'd2739, 16'd19948, 16'd31997, 16'd19603, 16'd5526, 16'd25896, 16'd1923, 16'd1586, 16'd36499, 16'd20902, 16'd36845, 16'd38929, 16'd5195, 16'd7313, 16'd2663, 16'd11268, 16'd31568, 16'd50868, 16'd36343, 16'd10757, 16'd31614});
	test_expansion(128'h1770ad104ee8f097aaab8692a210b993, {16'd2900, 16'd9426, 16'd53461, 16'd32583, 16'd36674, 16'd62365, 16'd41087, 16'd3961, 16'd9522, 16'd10168, 16'd60472, 16'd13714, 16'd26453, 16'd39278, 16'd50648, 16'd40192, 16'd2189, 16'd56995, 16'd423, 16'd35366, 16'd37755, 16'd22339, 16'd53255, 16'd51042, 16'd56820, 16'd32693});
	test_expansion(128'hd7822e8982e9400f8fdd72e5ff150e2c, {16'd64430, 16'd19002, 16'd54803, 16'd38390, 16'd18511, 16'd34215, 16'd19737, 16'd55022, 16'd16515, 16'd11393, 16'd3539, 16'd28190, 16'd12927, 16'd30754, 16'd35584, 16'd12757, 16'd62509, 16'd53223, 16'd18606, 16'd44564, 16'd58052, 16'd39507, 16'd10659, 16'd51504, 16'd36250, 16'd32954});
	test_expansion(128'hb3897ad5e649a743a725dc771ba0b8fb, {16'd58304, 16'd40863, 16'd4956, 16'd7624, 16'd7609, 16'd38167, 16'd14793, 16'd7283, 16'd16069, 16'd50715, 16'd62793, 16'd47427, 16'd63086, 16'd21469, 16'd44993, 16'd23059, 16'd45588, 16'd32581, 16'd10511, 16'd10882, 16'd11315, 16'd28059, 16'd13366, 16'd3917, 16'd52442, 16'd46707});
	test_expansion(128'h4c7c29788a22c1a304f1e509292dbd0c, {16'd7180, 16'd55844, 16'd55331, 16'd34726, 16'd42970, 16'd1336, 16'd42493, 16'd23254, 16'd14946, 16'd3688, 16'd38356, 16'd1332, 16'd52915, 16'd27698, 16'd23617, 16'd16119, 16'd41771, 16'd48644, 16'd59636, 16'd37145, 16'd7932, 16'd25460, 16'd47771, 16'd23899, 16'd61393, 16'd1070});
	test_expansion(128'hfd5dd7628e1a0fed5c8a6614f955dd2b, {16'd31778, 16'd23167, 16'd26125, 16'd43750, 16'd148, 16'd9446, 16'd62069, 16'd62841, 16'd29753, 16'd12123, 16'd38235, 16'd29769, 16'd8749, 16'd56134, 16'd15362, 16'd2000, 16'd45134, 16'd47572, 16'd7407, 16'd5005, 16'd38889, 16'd10161, 16'd58375, 16'd5718, 16'd4646, 16'd49258});
	test_expansion(128'hed1c65e01e100d96a37a27b089588ce9, {16'd44171, 16'd46210, 16'd30503, 16'd30366, 16'd56657, 16'd48953, 16'd41018, 16'd8199, 16'd7281, 16'd44248, 16'd15704, 16'd55404, 16'd17791, 16'd65479, 16'd43849, 16'd60878, 16'd6531, 16'd49568, 16'd8530, 16'd37012, 16'd63335, 16'd17159, 16'd26669, 16'd8509, 16'd55548, 16'd19822});
	test_expansion(128'hd523e71a34cc0f10fa4d2bcd1faeaa3f, {16'd28467, 16'd1451, 16'd33614, 16'd40047, 16'd40159, 16'd49643, 16'd29025, 16'd46498, 16'd53658, 16'd44496, 16'd20161, 16'd770, 16'd8643, 16'd10153, 16'd38920, 16'd8101, 16'd37115, 16'd1930, 16'd31769, 16'd5941, 16'd35964, 16'd56470, 16'd48939, 16'd53540, 16'd60162, 16'd22929});
	test_expansion(128'hb519fe770f15afea3763cd0fa6ad8c24, {16'd56251, 16'd56146, 16'd29402, 16'd33340, 16'd43788, 16'd15781, 16'd19254, 16'd60941, 16'd15488, 16'd23302, 16'd23946, 16'd24608, 16'd7419, 16'd5630, 16'd50970, 16'd28713, 16'd9549, 16'd55588, 16'd2049, 16'd2752, 16'd19983, 16'd59313, 16'd50355, 16'd58812, 16'd43397, 16'd10499});
	test_expansion(128'h3239331d0e9aa55fad25b1694d90a902, {16'd43862, 16'd64845, 16'd11893, 16'd53486, 16'd32539, 16'd6091, 16'd41531, 16'd47339, 16'd33379, 16'd43329, 16'd52360, 16'd29918, 16'd46880, 16'd54288, 16'd56273, 16'd7382, 16'd29649, 16'd3898, 16'd9786, 16'd1365, 16'd50077, 16'd33311, 16'd27752, 16'd45, 16'd47297, 16'd58602});
	test_expansion(128'h7a17251e484fc14ef329ee7128292378, {16'd18101, 16'd44967, 16'd43153, 16'd3549, 16'd45691, 16'd49182, 16'd51259, 16'd7594, 16'd52800, 16'd21628, 16'd54367, 16'd62743, 16'd51319, 16'd59336, 16'd22995, 16'd32331, 16'd61065, 16'd8199, 16'd51773, 16'd65427, 16'd3274, 16'd7871, 16'd49149, 16'd56245, 16'd12697, 16'd52341});
	test_expansion(128'h399dc6c646bcd90950b4efa2ede807d9, {16'd5058, 16'd5735, 16'd17990, 16'd1389, 16'd43814, 16'd56208, 16'd25376, 16'd17832, 16'd35152, 16'd38523, 16'd1046, 16'd19181, 16'd23906, 16'd62473, 16'd56412, 16'd63258, 16'd52103, 16'd5539, 16'd25848, 16'd32217, 16'd28457, 16'd28633, 16'd28323, 16'd11706, 16'd14627, 16'd50523});
	test_expansion(128'h20caf4f186b0d548a606649533bc0b24, {16'd63686, 16'd50018, 16'd33463, 16'd64215, 16'd38646, 16'd60991, 16'd59703, 16'd64521, 16'd10791, 16'd52976, 16'd44785, 16'd60323, 16'd48586, 16'd90, 16'd34528, 16'd27531, 16'd58910, 16'd15502, 16'd39828, 16'd34316, 16'd58490, 16'd42336, 16'd57687, 16'd48533, 16'd9629, 16'd63829});
	test_expansion(128'hb4ffaf0596f140cde04d309b5cbfa0a9, {16'd60299, 16'd19836, 16'd51829, 16'd16813, 16'd53105, 16'd24223, 16'd41321, 16'd42264, 16'd39641, 16'd62484, 16'd9405, 16'd18315, 16'd53693, 16'd50092, 16'd14180, 16'd8891, 16'd17899, 16'd47733, 16'd36557, 16'd33684, 16'd2512, 16'd13173, 16'd42935, 16'd233, 16'd48184, 16'd51442});
	test_expansion(128'hc127830d731a7f4fa2caae66e1bf052c, {16'd13559, 16'd51403, 16'd35771, 16'd49311, 16'd10529, 16'd1029, 16'd48132, 16'd53548, 16'd28067, 16'd2807, 16'd64233, 16'd18775, 16'd10061, 16'd18567, 16'd43702, 16'd27940, 16'd40577, 16'd48709, 16'd42883, 16'd63727, 16'd54900, 16'd30364, 16'd22598, 16'd11009, 16'd42145, 16'd48261});
	test_expansion(128'h087542d59b78a9f7411c481f83c58d8d, {16'd54522, 16'd48902, 16'd58147, 16'd32835, 16'd29533, 16'd19804, 16'd668, 16'd60517, 16'd51593, 16'd21139, 16'd30426, 16'd24865, 16'd30548, 16'd47414, 16'd22084, 16'd25548, 16'd62038, 16'd51449, 16'd30004, 16'd59102, 16'd13292, 16'd45010, 16'd9924, 16'd2125, 16'd18145, 16'd7260});
	test_expansion(128'h77540f7311750ab55a36a572a9480484, {16'd59639, 16'd32576, 16'd21449, 16'd45089, 16'd35776, 16'd12302, 16'd53867, 16'd13235, 16'd8937, 16'd56828, 16'd26998, 16'd13581, 16'd2674, 16'd13984, 16'd34609, 16'd49519, 16'd60453, 16'd3505, 16'd17902, 16'd60490, 16'd12591, 16'd9475, 16'd5872, 16'd17099, 16'd47552, 16'd33326});
	test_expansion(128'h696f77e92720c2a686e5afd52732830c, {16'd15251, 16'd5934, 16'd35660, 16'd31531, 16'd3943, 16'd40904, 16'd9281, 16'd46390, 16'd52130, 16'd10951, 16'd11418, 16'd43073, 16'd42971, 16'd42716, 16'd64688, 16'd17451, 16'd4620, 16'd16808, 16'd3075, 16'd51301, 16'd32345, 16'd16832, 16'd4202, 16'd3481, 16'd48829, 16'd52950});
	test_expansion(128'h22a31c76f3a7295571e4627754f165a6, {16'd47294, 16'd36210, 16'd51083, 16'd50355, 16'd32786, 16'd10815, 16'd20647, 16'd56726, 16'd7450, 16'd62233, 16'd27934, 16'd54903, 16'd49373, 16'd42129, 16'd21229, 16'd65226, 16'd3294, 16'd19097, 16'd13047, 16'd56442, 16'd18216, 16'd17174, 16'd20112, 16'd43127, 16'd50971, 16'd40308});
	test_expansion(128'h995ac91cbccad31d0bbed38474213f3c, {16'd38810, 16'd48442, 16'd28243, 16'd13316, 16'd50099, 16'd52878, 16'd7133, 16'd51655, 16'd47941, 16'd48313, 16'd40563, 16'd15863, 16'd64152, 16'd60927, 16'd42786, 16'd14590, 16'd18505, 16'd55380, 16'd6428, 16'd61446, 16'd47330, 16'd53344, 16'd60135, 16'd45704, 16'd52417, 16'd42328});
	test_expansion(128'ha3c7284cf0f68bede3c53c3d09a41a5a, {16'd43225, 16'd47871, 16'd4821, 16'd57852, 16'd18712, 16'd16921, 16'd56551, 16'd48144, 16'd13550, 16'd54635, 16'd49436, 16'd29116, 16'd38341, 16'd8315, 16'd17715, 16'd48774, 16'd112, 16'd29079, 16'd16500, 16'd5526, 16'd34882, 16'd30195, 16'd33497, 16'd60149, 16'd42841, 16'd61025});
	test_expansion(128'h19a00ee77b8b81ff0c5835a82bf5e5d9, {16'd10075, 16'd45496, 16'd19727, 16'd65501, 16'd6192, 16'd58853, 16'd10326, 16'd60025, 16'd49067, 16'd39221, 16'd35170, 16'd11009, 16'd15458, 16'd52811, 16'd43539, 16'd22483, 16'd40884, 16'd3522, 16'd59696, 16'd9276, 16'd20423, 16'd3241, 16'd14601, 16'd58928, 16'd533, 16'd61306});
	test_expansion(128'h4bbacd9b4f4b9d9f85f4d6ecdcf327d3, {16'd47261, 16'd3553, 16'd28854, 16'd12195, 16'd13576, 16'd24947, 16'd9569, 16'd34264, 16'd2577, 16'd35445, 16'd51709, 16'd50461, 16'd33590, 16'd25888, 16'd13557, 16'd46635, 16'd9688, 16'd45663, 16'd22558, 16'd34593, 16'd33086, 16'd32459, 16'd4215, 16'd46962, 16'd63246, 16'd61374});
	test_expansion(128'h1c2aa40f554f2f803560c700e7faa056, {16'd29068, 16'd30874, 16'd32649, 16'd979, 16'd56099, 16'd63841, 16'd40685, 16'd15269, 16'd48387, 16'd12547, 16'd23429, 16'd50290, 16'd57482, 16'd56158, 16'd28929, 16'd22543, 16'd56578, 16'd40161, 16'd7493, 16'd23374, 16'd52151, 16'd37916, 16'd46857, 16'd42115, 16'd10854, 16'd43985});
	test_expansion(128'he01eb91dd478762f22960cc0b70eef44, {16'd34961, 16'd34984, 16'd13021, 16'd1721, 16'd1209, 16'd56325, 16'd21383, 16'd65114, 16'd36974, 16'd1672, 16'd59002, 16'd40245, 16'd42220, 16'd10519, 16'd42190, 16'd3388, 16'd54007, 16'd38814, 16'd64162, 16'd27282, 16'd36612, 16'd23664, 16'd7087, 16'd2822, 16'd47530, 16'd33492});
	test_expansion(128'h6f4295c4cbe98ff46b992e37c59f1dc5, {16'd56016, 16'd63586, 16'd43862, 16'd6821, 16'd37517, 16'd41602, 16'd951, 16'd15334, 16'd4079, 16'd42522, 16'd41702, 16'd3835, 16'd26526, 16'd62082, 16'd53574, 16'd36590, 16'd4422, 16'd58652, 16'd42749, 16'd10387, 16'd59541, 16'd33385, 16'd7380, 16'd42616, 16'd16345, 16'd18369});
	test_expansion(128'hf21457749559a7b9c380fe3743fa838d, {16'd20831, 16'd24609, 16'd31980, 16'd20019, 16'd31441, 16'd7049, 16'd43301, 16'd54776, 16'd57453, 16'd33802, 16'd58046, 16'd3243, 16'd11192, 16'd41803, 16'd21337, 16'd22179, 16'd63258, 16'd43096, 16'd31122, 16'd18017, 16'd48551, 16'd51096, 16'd7103, 16'd54932, 16'd2590, 16'd47642});
	test_expansion(128'hffa78825290d3216ecdfe306c5ed1465, {16'd17514, 16'd4339, 16'd38461, 16'd905, 16'd46090, 16'd48579, 16'd60487, 16'd41534, 16'd43106, 16'd31863, 16'd49231, 16'd6512, 16'd1117, 16'd6852, 16'd13507, 16'd17690, 16'd32401, 16'd60198, 16'd54267, 16'd373, 16'd32493, 16'd14521, 16'd63277, 16'd50067, 16'd46517, 16'd2510});
	test_expansion(128'h1800aaa23517968b916933adc7438858, {16'd44338, 16'd9119, 16'd64880, 16'd42334, 16'd45907, 16'd43032, 16'd59296, 16'd5181, 16'd43037, 16'd17497, 16'd15896, 16'd1453, 16'd1150, 16'd46530, 16'd20722, 16'd19592, 16'd31273, 16'd595, 16'd3038, 16'd42626, 16'd26266, 16'd33433, 16'd28792, 16'd7849, 16'd24790, 16'd21012});
	test_expansion(128'h6c865f6c21b887102e8df04cc2381977, {16'd7543, 16'd37305, 16'd36767, 16'd51187, 16'd12936, 16'd30763, 16'd46589, 16'd24758, 16'd32444, 16'd55673, 16'd23462, 16'd61329, 16'd42759, 16'd64490, 16'd20782, 16'd60142, 16'd842, 16'd13370, 16'd22655, 16'd53255, 16'd19910, 16'd29338, 16'd34227, 16'd52850, 16'd35063, 16'd54405});
	test_expansion(128'h6edaf7ef4a00eeb66afcbe3d49ba081d, {16'd55127, 16'd35572, 16'd52829, 16'd12043, 16'd18430, 16'd33110, 16'd27239, 16'd62005, 16'd21601, 16'd60315, 16'd5413, 16'd51751, 16'd62716, 16'd11928, 16'd60082, 16'd44703, 16'd39978, 16'd52544, 16'd46277, 16'd59914, 16'd63322, 16'd21576, 16'd63390, 16'd64726, 16'd14531, 16'd6634});
	test_expansion(128'h5c2efdbf1f2e8179be4f393492dbe9fb, {16'd4340, 16'd2040, 16'd54244, 16'd31618, 16'd12984, 16'd50575, 16'd53010, 16'd40980, 16'd45210, 16'd9040, 16'd52255, 16'd54879, 16'd45575, 16'd41935, 16'd42950, 16'd57365, 16'd54588, 16'd45247, 16'd43700, 16'd51520, 16'd41568, 16'd1400, 16'd36094, 16'd22612, 16'd22853, 16'd19087});
	test_expansion(128'h4d8fe4758f0711142ffffa66f8affff6, {16'd50503, 16'd26683, 16'd42767, 16'd3347, 16'd48969, 16'd38343, 16'd65409, 16'd43095, 16'd4914, 16'd11632, 16'd36962, 16'd26804, 16'd37343, 16'd55310, 16'd23588, 16'd41049, 16'd50756, 16'd12975, 16'd34987, 16'd6475, 16'd52905, 16'd59212, 16'd49629, 16'd51544, 16'd30336, 16'd12617});
	test_expansion(128'heaf5d759a7e7879fa376913ddda3fde4, {16'd13768, 16'd14770, 16'd7724, 16'd56640, 16'd42900, 16'd62577, 16'd44039, 16'd57355, 16'd65229, 16'd6440, 16'd54753, 16'd19405, 16'd29248, 16'd45870, 16'd15927, 16'd39192, 16'd63129, 16'd31584, 16'd38574, 16'd53654, 16'd38588, 16'd43252, 16'd16717, 16'd17550, 16'd14203, 16'd38287});
	test_expansion(128'h370309f7de13b5342d6dab3abff1eb43, {16'd62797, 16'd6728, 16'd32996, 16'd37063, 16'd17784, 16'd6759, 16'd33892, 16'd46776, 16'd5245, 16'd2464, 16'd42447, 16'd16199, 16'd57004, 16'd3595, 16'd13935, 16'd26552, 16'd59603, 16'd20037, 16'd44048, 16'd27520, 16'd59448, 16'd51495, 16'd46934, 16'd31238, 16'd58567, 16'd5362});
	test_expansion(128'h76cc30bd3d67aab220be3c6356bec12b, {16'd55548, 16'd21842, 16'd25564, 16'd50742, 16'd15604, 16'd62051, 16'd24597, 16'd8800, 16'd11326, 16'd3519, 16'd55703, 16'd49527, 16'd21998, 16'd26590, 16'd23243, 16'd5743, 16'd5572, 16'd4477, 16'd36451, 16'd22338, 16'd27229, 16'd52261, 16'd59220, 16'd22671, 16'd21356, 16'd12928});
	test_expansion(128'he45da416531dff22cd238c9cc55fcd11, {16'd51293, 16'd32662, 16'd53454, 16'd3855, 16'd2931, 16'd10768, 16'd49773, 16'd46039, 16'd21721, 16'd63480, 16'd53483, 16'd9270, 16'd50966, 16'd1056, 16'd30332, 16'd3259, 16'd19234, 16'd22684, 16'd43803, 16'd58798, 16'd27323, 16'd8162, 16'd55978, 16'd51421, 16'd4322, 16'd46890});
	test_expansion(128'hbfaed1e037fcd1fad2331a88da78b40c, {16'd39978, 16'd25149, 16'd20997, 16'd14422, 16'd39220, 16'd63519, 16'd19122, 16'd20731, 16'd39988, 16'd38262, 16'd47846, 16'd5577, 16'd16751, 16'd37322, 16'd40854, 16'd27987, 16'd51195, 16'd38977, 16'd30494, 16'd7379, 16'd5983, 16'd23342, 16'd1510, 16'd56342, 16'd32954, 16'd40950});
	test_expansion(128'h051bfe603f9f43488c5be3099ca96131, {16'd33094, 16'd46297, 16'd13810, 16'd41405, 16'd31389, 16'd4518, 16'd4748, 16'd49718, 16'd9319, 16'd4853, 16'd40582, 16'd176, 16'd62302, 16'd59267, 16'd15624, 16'd51088, 16'd14479, 16'd17242, 16'd42785, 16'd48475, 16'd46074, 16'd57602, 16'd10137, 16'd5488, 16'd3271, 16'd17966});
	test_expansion(128'hadf899a3096c357d3deda4b07323dce1, {16'd11816, 16'd18144, 16'd33711, 16'd58953, 16'd18075, 16'd24898, 16'd45397, 16'd62115, 16'd64570, 16'd31646, 16'd46936, 16'd12062, 16'd53053, 16'd62616, 16'd9155, 16'd17491, 16'd2050, 16'd49149, 16'd54715, 16'd14806, 16'd29774, 16'd12283, 16'd33694, 16'd25754, 16'd49694, 16'd12313});
	test_expansion(128'h6ba60e4b126af79da5855db6c3538359, {16'd62808, 16'd5760, 16'd30866, 16'd23225, 16'd50498, 16'd56141, 16'd3924, 16'd35105, 16'd53842, 16'd47911, 16'd25252, 16'd33991, 16'd23256, 16'd7701, 16'd11944, 16'd6979, 16'd43441, 16'd24674, 16'd13228, 16'd20313, 16'd59223, 16'd49656, 16'd32080, 16'd63564, 16'd61405, 16'd29172});
	test_expansion(128'he51128620e72b74468b730c9c7fe7475, {16'd47903, 16'd26188, 16'd45886, 16'd41076, 16'd21877, 16'd45160, 16'd55000, 16'd3591, 16'd7177, 16'd18762, 16'd59414, 16'd61728, 16'd21241, 16'd52566, 16'd3061, 16'd644, 16'd47720, 16'd27163, 16'd53632, 16'd16143, 16'd54882, 16'd29940, 16'd8532, 16'd44445, 16'd2318, 16'd33244});
	test_expansion(128'hc842c8250b4ea989d4927a97f2ae6951, {16'd58050, 16'd15622, 16'd64946, 16'd41911, 16'd12595, 16'd16202, 16'd60365, 16'd9244, 16'd14643, 16'd26199, 16'd10869, 16'd51049, 16'd20896, 16'd35907, 16'd26187, 16'd25574, 16'd16639, 16'd39632, 16'd8998, 16'd22589, 16'd17297, 16'd40110, 16'd30338, 16'd53632, 16'd64590, 16'd36694});
	test_expansion(128'h0ecfb6a5cfb30a0ed7a3d32de6c68bcf, {16'd49680, 16'd50580, 16'd34644, 16'd64346, 16'd60259, 16'd43113, 16'd17519, 16'd19520, 16'd33789, 16'd15881, 16'd33919, 16'd14817, 16'd49055, 16'd25242, 16'd22708, 16'd31050, 16'd55957, 16'd25267, 16'd37628, 16'd63952, 16'd53441, 16'd27298, 16'd53, 16'd46732, 16'd34529, 16'd43428});
	test_expansion(128'h7c1fc5a5933f9ea74415dfe2829ab603, {16'd53995, 16'd9971, 16'd63939, 16'd12106, 16'd21453, 16'd13251, 16'd50426, 16'd47233, 16'd57, 16'd31745, 16'd27557, 16'd59834, 16'd8393, 16'd52454, 16'd55030, 16'd12963, 16'd20590, 16'd58498, 16'd43769, 16'd63800, 16'd24248, 16'd33934, 16'd19147, 16'd20907, 16'd29684, 16'd20461});
	test_expansion(128'h0084dfcdaed10a3e8aa59ecf94d42e55, {16'd10718, 16'd11491, 16'd50587, 16'd54161, 16'd34632, 16'd19117, 16'd14813, 16'd40662, 16'd5477, 16'd13943, 16'd16942, 16'd57779, 16'd33946, 16'd2937, 16'd34453, 16'd48612, 16'd4453, 16'd18436, 16'd38037, 16'd23941, 16'd6277, 16'd27303, 16'd39751, 16'd51994, 16'd61237, 16'd5675});
	test_expansion(128'h3ec950f025386544bdf234f071817275, {16'd61335, 16'd63038, 16'd2647, 16'd54204, 16'd16721, 16'd6662, 16'd23185, 16'd63985, 16'd56996, 16'd65236, 16'd9535, 16'd12938, 16'd6163, 16'd16958, 16'd59715, 16'd20285, 16'd41030, 16'd32709, 16'd23869, 16'd21449, 16'd4412, 16'd57930, 16'd13033, 16'd19369, 16'd60404, 16'd502});
	test_expansion(128'h5711805ca80ab58b1810f5f5aba2d665, {16'd4823, 16'd25100, 16'd54165, 16'd21605, 16'd29006, 16'd63269, 16'd54947, 16'd16657, 16'd38325, 16'd47131, 16'd22669, 16'd56234, 16'd36322, 16'd33531, 16'd59237, 16'd52270, 16'd44077, 16'd64362, 16'd27557, 16'd6029, 16'd58117, 16'd56074, 16'd46022, 16'd31423, 16'd10824, 16'd5981});
	test_expansion(128'hf085e95b21ae831cac06400d12739a09, {16'd45965, 16'd2679, 16'd60282, 16'd55536, 16'd4831, 16'd30110, 16'd59860, 16'd4273, 16'd890, 16'd25046, 16'd20836, 16'd65233, 16'd1986, 16'd56844, 16'd33875, 16'd53817, 16'd20522, 16'd43070, 16'd50542, 16'd32239, 16'd8512, 16'd54746, 16'd16792, 16'd28865, 16'd4522, 16'd6025});
	test_expansion(128'hfeb6e612be6654bba32d5f37520b7465, {16'd56707, 16'd38223, 16'd54045, 16'd33840, 16'd20875, 16'd21605, 16'd43113, 16'd2961, 16'd7344, 16'd33872, 16'd52353, 16'd30811, 16'd13825, 16'd34823, 16'd35554, 16'd42685, 16'd45258, 16'd61081, 16'd18122, 16'd59907, 16'd50808, 16'd5761, 16'd19822, 16'd7096, 16'd8245, 16'd24156});
	test_expansion(128'ha6279bcb7fddce3e54c8a2a323f04596, {16'd11070, 16'd11776, 16'd31079, 16'd45891, 16'd13294, 16'd56192, 16'd22860, 16'd7942, 16'd45443, 16'd41947, 16'd55986, 16'd61014, 16'd49212, 16'd63198, 16'd59304, 16'd58336, 16'd28981, 16'd59520, 16'd20326, 16'd48635, 16'd25974, 16'd6226, 16'd22997, 16'd36028, 16'd60320, 16'd7643});
	test_expansion(128'he25e22f16c61834c2fb660ddecccb77a, {16'd34587, 16'd55081, 16'd9317, 16'd53469, 16'd25858, 16'd6988, 16'd54490, 16'd36213, 16'd49339, 16'd11558, 16'd47775, 16'd13293, 16'd62123, 16'd46216, 16'd11081, 16'd60883, 16'd38700, 16'd12252, 16'd2403, 16'd63077, 16'd2200, 16'd54270, 16'd408, 16'd29182, 16'd10483, 16'd2945});
	test_expansion(128'h40ae91e0530942f43e764205c61441d6, {16'd10193, 16'd11664, 16'd36852, 16'd33894, 16'd21037, 16'd64932, 16'd1225, 16'd33432, 16'd7470, 16'd42646, 16'd38111, 16'd27521, 16'd16977, 16'd39878, 16'd56761, 16'd62201, 16'd55241, 16'd33870, 16'd58566, 16'd3636, 16'd23064, 16'd7977, 16'd57970, 16'd27687, 16'd1705, 16'd18779});
	test_expansion(128'haf7a41fc0f543e02bb616f612f14a2f3, {16'd58925, 16'd12124, 16'd23217, 16'd14528, 16'd12894, 16'd37719, 16'd41351, 16'd46845, 16'd37581, 16'd60434, 16'd15546, 16'd56253, 16'd41244, 16'd17568, 16'd32757, 16'd10462, 16'd13133, 16'd24265, 16'd26820, 16'd1679, 16'd29319, 16'd11783, 16'd2733, 16'd23113, 16'd53455, 16'd4209});
	test_expansion(128'hc52fe90ac9dd0f14f48b9cc406d45571, {16'd51348, 16'd27209, 16'd11342, 16'd27893, 16'd47285, 16'd54481, 16'd37996, 16'd14933, 16'd64449, 16'd14341, 16'd41848, 16'd13052, 16'd5821, 16'd39633, 16'd51294, 16'd30174, 16'd25026, 16'd16970, 16'd36833, 16'd38438, 16'd48586, 16'd38562, 16'd46238, 16'd50018, 16'd7815, 16'd36300});
	test_expansion(128'h16d8396ad95b8c2aee91206ba41d9ecd, {16'd10431, 16'd11183, 16'd21853, 16'd43788, 16'd53125, 16'd58963, 16'd7565, 16'd40189, 16'd1251, 16'd7971, 16'd11184, 16'd45525, 16'd25628, 16'd15584, 16'd568, 16'd29055, 16'd55699, 16'd11728, 16'd55181, 16'd224, 16'd674, 16'd27985, 16'd24242, 16'd28374, 16'd11698, 16'd49368});
	test_expansion(128'h7f6bfd9ada82021319ea2b03920a9237, {16'd11982, 16'd55395, 16'd33103, 16'd14572, 16'd16802, 16'd50563, 16'd25696, 16'd9845, 16'd26636, 16'd19824, 16'd23768, 16'd61827, 16'd64796, 16'd48647, 16'd17954, 16'd18519, 16'd32353, 16'd42651, 16'd49080, 16'd35303, 16'd1159, 16'd55251, 16'd22745, 16'd7132, 16'd48903, 16'd12875});
	test_expansion(128'hb758b30151e27ed22e1cc48133703e8a, {16'd25575, 16'd47629, 16'd3857, 16'd57783, 16'd34280, 16'd33537, 16'd52812, 16'd364, 16'd21106, 16'd3716, 16'd44157, 16'd62384, 16'd33457, 16'd54327, 16'd14455, 16'd41276, 16'd2166, 16'd11288, 16'd53483, 16'd21848, 16'd9170, 16'd16183, 16'd31659, 16'd60653, 16'd20799, 16'd23141});
	test_expansion(128'ha53c1713c2dbfeac62bec3052049fca3, {16'd33976, 16'd54749, 16'd30038, 16'd46041, 16'd42034, 16'd61270, 16'd5041, 16'd38972, 16'd28275, 16'd27791, 16'd37443, 16'd9379, 16'd20021, 16'd32068, 16'd64211, 16'd60516, 16'd7117, 16'd21328, 16'd11499, 16'd39028, 16'd3256, 16'd12831, 16'd59166, 16'd14964, 16'd4149, 16'd5986});
	test_expansion(128'hf4de2e42ff15e1f62e64f71e88848f29, {16'd26250, 16'd33993, 16'd6233, 16'd48054, 16'd18679, 16'd55415, 16'd57976, 16'd17196, 16'd9939, 16'd33503, 16'd47678, 16'd13058, 16'd5270, 16'd62758, 16'd17369, 16'd63415, 16'd59287, 16'd36335, 16'd48270, 16'd30542, 16'd3227, 16'd35674, 16'd61547, 16'd8966, 16'd22108, 16'd47754});
	test_expansion(128'hc7a63344751291953868057e6dd879ba, {16'd6234, 16'd4232, 16'd42287, 16'd18213, 16'd38718, 16'd42372, 16'd35886, 16'd36805, 16'd4755, 16'd16459, 16'd40132, 16'd15696, 16'd9917, 16'd28610, 16'd42553, 16'd17629, 16'd60067, 16'd33248, 16'd19320, 16'd35286, 16'd53143, 16'd6572, 16'd1126, 16'd40881, 16'd64756, 16'd31535});
	test_expansion(128'h0678a9feda071e48d8f554059396d5f8, {16'd12712, 16'd51966, 16'd11291, 16'd43866, 16'd46030, 16'd34145, 16'd34179, 16'd64545, 16'd48027, 16'd24776, 16'd1551, 16'd30044, 16'd46395, 16'd40736, 16'd2668, 16'd45760, 16'd55030, 16'd45211, 16'd63190, 16'd22661, 16'd60510, 16'd48847, 16'd57891, 16'd43743, 16'd12079, 16'd62588});
	test_expansion(128'h32f4ca130492c64aa9e4dc93cfd2d139, {16'd13978, 16'd14341, 16'd26452, 16'd15887, 16'd28785, 16'd2103, 16'd59267, 16'd34180, 16'd976, 16'd30120, 16'd13094, 16'd57284, 16'd64561, 16'd54509, 16'd37730, 16'd42414, 16'd38479, 16'd29998, 16'd24305, 16'd45573, 16'd23476, 16'd3163, 16'd29135, 16'd47072, 16'd46360, 16'd23015});
	test_expansion(128'h778993239202e3bcd4928b5a17ff5ba9, {16'd58031, 16'd16922, 16'd9841, 16'd25096, 16'd59915, 16'd29640, 16'd37710, 16'd2450, 16'd25202, 16'd7371, 16'd13059, 16'd25160, 16'd64505, 16'd44767, 16'd15636, 16'd17079, 16'd42659, 16'd39380, 16'd46230, 16'd63391, 16'd21581, 16'd24605, 16'd4158, 16'd33769, 16'd14949, 16'd61764});
	test_expansion(128'hd121ae484792202f6a5184b35cb1cb53, {16'd34757, 16'd39476, 16'd44850, 16'd11994, 16'd13321, 16'd36273, 16'd30394, 16'd48032, 16'd46284, 16'd42251, 16'd35243, 16'd23725, 16'd61609, 16'd22932, 16'd38093, 16'd3774, 16'd54563, 16'd41512, 16'd35522, 16'd30089, 16'd9427, 16'd56595, 16'd10033, 16'd4673, 16'd681, 16'd25270});
	test_expansion(128'hb2766d4391f15a6064796f0dbff20e87, {16'd1172, 16'd60994, 16'd48806, 16'd45853, 16'd16166, 16'd7494, 16'd45474, 16'd2933, 16'd25444, 16'd21682, 16'd64739, 16'd65206, 16'd26308, 16'd46246, 16'd24272, 16'd18508, 16'd40792, 16'd31085, 16'd26911, 16'd45625, 16'd52370, 16'd50358, 16'd36252, 16'd33842, 16'd19063, 16'd55901});
	test_expansion(128'hd5fd52fb667c439c5e8a420eeafd6ff0, {16'd54719, 16'd45413, 16'd26978, 16'd25276, 16'd63337, 16'd9928, 16'd28922, 16'd24050, 16'd30469, 16'd54532, 16'd333, 16'd44278, 16'd17223, 16'd955, 16'd54688, 16'd43851, 16'd61445, 16'd41332, 16'd55092, 16'd17012, 16'd7356, 16'd35218, 16'd23701, 16'd57330, 16'd25806, 16'd10460});
	test_expansion(128'h7231a52c77d1e080cd7311c267cf21c6, {16'd6494, 16'd50547, 16'd21025, 16'd59651, 16'd56311, 16'd1141, 16'd24160, 16'd26084, 16'd31780, 16'd65047, 16'd16336, 16'd44352, 16'd27997, 16'd47762, 16'd4464, 16'd25682, 16'd319, 16'd12973, 16'd56160, 16'd14990, 16'd38379, 16'd25267, 16'd10269, 16'd21753, 16'd23322, 16'd49473});
	test_expansion(128'h782c2468316a5a7942a3c0faf34faedb, {16'd54051, 16'd30156, 16'd19880, 16'd2553, 16'd29896, 16'd37140, 16'd44675, 16'd53401, 16'd23400, 16'd28198, 16'd59025, 16'd34609, 16'd21139, 16'd40378, 16'd39795, 16'd13146, 16'd5575, 16'd36476, 16'd9372, 16'd24246, 16'd10740, 16'd4143, 16'd38559, 16'd16614, 16'd62015, 16'd54365});
	test_expansion(128'he73dc620b7c3532fc2c074e4195f77a0, {16'd25625, 16'd63077, 16'd56363, 16'd48263, 16'd48202, 16'd43262, 16'd58211, 16'd28047, 16'd56937, 16'd32096, 16'd12528, 16'd34276, 16'd60277, 16'd14265, 16'd19007, 16'd33, 16'd56340, 16'd62744, 16'd51639, 16'd3841, 16'd122, 16'd4320, 16'd15817, 16'd3469, 16'd47430, 16'd27561});
	test_expansion(128'h1a3c5819c9f249bf277f348e07075022, {16'd49267, 16'd4718, 16'd63366, 16'd35475, 16'd46793, 16'd25262, 16'd37384, 16'd55868, 16'd35290, 16'd8847, 16'd10060, 16'd60011, 16'd41635, 16'd45086, 16'd20296, 16'd59424, 16'd7817, 16'd31246, 16'd47882, 16'd47943, 16'd60631, 16'd17147, 16'd24186, 16'd13456, 16'd47808, 16'd41153});
	test_expansion(128'h80ce0c88651c2405f07d5309ffd47c89, {16'd15125, 16'd44936, 16'd26312, 16'd29946, 16'd20077, 16'd39554, 16'd57897, 16'd45974, 16'd19831, 16'd46430, 16'd38614, 16'd30823, 16'd18221, 16'd36916, 16'd51937, 16'd59090, 16'd53160, 16'd36455, 16'd2693, 16'd7288, 16'd47252, 16'd46543, 16'd60104, 16'd16890, 16'd54905, 16'd61582});
	test_expansion(128'ha27981d7a26dfbad6c03a7b138a78721, {16'd37663, 16'd401, 16'd16384, 16'd33057, 16'd17766, 16'd19985, 16'd63810, 16'd58825, 16'd10975, 16'd65398, 16'd2810, 16'd38765, 16'd15060, 16'd14736, 16'd21536, 16'd41222, 16'd1142, 16'd1917, 16'd21433, 16'd33292, 16'd45898, 16'd45379, 16'd4544, 16'd61484, 16'd23458, 16'd37540});
	test_expansion(128'h956b451887379b262298d7ade762a901, {16'd18144, 16'd46181, 16'd62945, 16'd11647, 16'd27404, 16'd49665, 16'd48869, 16'd61994, 16'd3060, 16'd52258, 16'd23132, 16'd20185, 16'd56587, 16'd56306, 16'd61130, 16'd2165, 16'd47730, 16'd60584, 16'd50870, 16'd28892, 16'd55660, 16'd6101, 16'd51812, 16'd31407, 16'd52720, 16'd17416});
	test_expansion(128'h5f47ffa088f5fec15189224cc0f1eb59, {16'd18746, 16'd47300, 16'd10097, 16'd50989, 16'd26448, 16'd5067, 16'd43764, 16'd55996, 16'd64961, 16'd62364, 16'd61638, 16'd1486, 16'd37114, 16'd43938, 16'd17940, 16'd46220, 16'd54749, 16'd12844, 16'd32270, 16'd53647, 16'd30328, 16'd40890, 16'd32183, 16'd25530, 16'd11515, 16'd13751});
	test_expansion(128'h947804494d58f1159399dae4e2ca444c, {16'd60810, 16'd32783, 16'd28317, 16'd47178, 16'd24300, 16'd14692, 16'd49008, 16'd39993, 16'd37193, 16'd38842, 16'd20988, 16'd52003, 16'd58059, 16'd59127, 16'd15546, 16'd35287, 16'd30314, 16'd29638, 16'd62497, 16'd26513, 16'd51628, 16'd39008, 16'd16755, 16'd24192, 16'd47122, 16'd53530});
	test_expansion(128'hf9aa9203564babbd1aee1ec85e927b3e, {16'd40318, 16'd34589, 16'd1173, 16'd19950, 16'd20339, 16'd54769, 16'd52954, 16'd7097, 16'd30457, 16'd21553, 16'd28795, 16'd18064, 16'd24124, 16'd46508, 16'd44621, 16'd973, 16'd33145, 16'd994, 16'd60902, 16'd61895, 16'd21364, 16'd35419, 16'd27963, 16'd28674, 16'd42546, 16'd7737});
	test_expansion(128'heea343f38fbfa32d5f6039d8c9ec929e, {16'd21271, 16'd42719, 16'd14444, 16'd45544, 16'd43930, 16'd62753, 16'd64167, 16'd28419, 16'd50654, 16'd52167, 16'd64035, 16'd56662, 16'd7543, 16'd44919, 16'd55335, 16'd40268, 16'd1961, 16'd50800, 16'd4276, 16'd5941, 16'd50057, 16'd33210, 16'd21908, 16'd37935, 16'd64525, 16'd24385});
	test_expansion(128'h41a882cb8f1f697b43679d3b81b58341, {16'd31456, 16'd59570, 16'd27708, 16'd51264, 16'd23673, 16'd60952, 16'd45840, 16'd33779, 16'd19342, 16'd39611, 16'd15771, 16'd1035, 16'd5720, 16'd16183, 16'd43845, 16'd12891, 16'd55848, 16'd9645, 16'd6688, 16'd40576, 16'd28405, 16'd25877, 16'd17860, 16'd16581, 16'd27554, 16'd3408});
	test_expansion(128'h001d4b8f8af3bf3e1a881d854f3b45c2, {16'd52077, 16'd26136, 16'd50354, 16'd56243, 16'd35660, 16'd28641, 16'd35335, 16'd52557, 16'd42730, 16'd20152, 16'd12229, 16'd54907, 16'd43347, 16'd39240, 16'd62024, 16'd29241, 16'd17216, 16'd35291, 16'd29397, 16'd3706, 16'd33191, 16'd44248, 16'd51107, 16'd22103, 16'd37770, 16'd14208});
	test_expansion(128'h7b2d97b91427df13a793c1fea1c57180, {16'd34015, 16'd6506, 16'd34237, 16'd41289, 16'd11806, 16'd18253, 16'd49220, 16'd65028, 16'd8421, 16'd24424, 16'd65037, 16'd2897, 16'd48949, 16'd222, 16'd29872, 16'd42372, 16'd10402, 16'd62834, 16'd28631, 16'd41183, 16'd31850, 16'd25416, 16'd6065, 16'd24112, 16'd51890, 16'd8495});
	test_expansion(128'h111d9df63fdfbc47e9d232900ec6c056, {16'd63389, 16'd37947, 16'd9725, 16'd56351, 16'd23664, 16'd3095, 16'd35149, 16'd35908, 16'd31265, 16'd34119, 16'd56811, 16'd34437, 16'd25467, 16'd45979, 16'd61022, 16'd34283, 16'd41418, 16'd14489, 16'd13498, 16'd22215, 16'd59458, 16'd32281, 16'd15934, 16'd19458, 16'd31584, 16'd28846});
	test_expansion(128'hd97e118390d060e934e4c70a90303e0a, {16'd5495, 16'd64784, 16'd35764, 16'd42962, 16'd56470, 16'd43876, 16'd21909, 16'd53440, 16'd25369, 16'd24608, 16'd39861, 16'd17116, 16'd63609, 16'd14443, 16'd57680, 16'd46054, 16'd51994, 16'd24145, 16'd20596, 16'd13471, 16'd24992, 16'd4263, 16'd42995, 16'd3815, 16'd39669, 16'd47769});
	test_expansion(128'hef439a12d4564b67d7b4b0a5f8605559, {16'd34790, 16'd26569, 16'd52, 16'd62240, 16'd8175, 16'd19605, 16'd37901, 16'd64218, 16'd5406, 16'd2857, 16'd2341, 16'd51551, 16'd56558, 16'd57115, 16'd23594, 16'd52064, 16'd9660, 16'd37201, 16'd47979, 16'd59156, 16'd37283, 16'd7599, 16'd29732, 16'd39131, 16'd8120, 16'd12003});
	test_expansion(128'hd1eb5ed7c0b5f7e0e2f0eaa9a5663e05, {16'd56104, 16'd2705, 16'd62168, 16'd62989, 16'd11684, 16'd33864, 16'd7782, 16'd21434, 16'd59851, 16'd17094, 16'd5993, 16'd54046, 16'd45147, 16'd33878, 16'd57608, 16'd36878, 16'd64079, 16'd51203, 16'd45500, 16'd60175, 16'd34160, 16'd27132, 16'd54447, 16'd5879, 16'd8456, 16'd22726});
	test_expansion(128'h55d1d726f0b3408233572897294e2a42, {16'd56236, 16'd31530, 16'd33686, 16'd47978, 16'd50569, 16'd41999, 16'd24403, 16'd40247, 16'd31348, 16'd15399, 16'd50675, 16'd54506, 16'd54776, 16'd21698, 16'd49883, 16'd31956, 16'd6349, 16'd22699, 16'd16549, 16'd23478, 16'd48220, 16'd7029, 16'd12659, 16'd64351, 16'd52007, 16'd54650});
	test_expansion(128'h968dc150feea8ff76de1606c7200072d, {16'd3185, 16'd50082, 16'd32841, 16'd51687, 16'd24432, 16'd30614, 16'd1640, 16'd3143, 16'd35322, 16'd54138, 16'd2685, 16'd56975, 16'd8192, 16'd31067, 16'd8147, 16'd51679, 16'd7222, 16'd31071, 16'd52677, 16'd14908, 16'd21004, 16'd56433, 16'd34408, 16'd61607, 16'd47816, 16'd52964});
	test_expansion(128'h5bc394596545dbd064652cf2f7635d5e, {16'd3374, 16'd60057, 16'd27342, 16'd49982, 16'd319, 16'd52061, 16'd3349, 16'd61693, 16'd4814, 16'd25177, 16'd19204, 16'd38795, 16'd32428, 16'd1401, 16'd39246, 16'd29898, 16'd40892, 16'd61882, 16'd63848, 16'd10833, 16'd9171, 16'd45776, 16'd28490, 16'd13968, 16'd1406, 16'd27655});
	test_expansion(128'hc31ec17837ffe85783506bbbce31e17b, {16'd23765, 16'd12242, 16'd7313, 16'd39992, 16'd31638, 16'd34797, 16'd2229, 16'd56039, 16'd36004, 16'd25123, 16'd35616, 16'd47396, 16'd21627, 16'd26863, 16'd23005, 16'd45126, 16'd20641, 16'd62202, 16'd46780, 16'd51799, 16'd30417, 16'd54078, 16'd55060, 16'd9684, 16'd6032, 16'd62940});
	test_expansion(128'h6c2254c3988c720e962ba815c8ac1cbf, {16'd54337, 16'd39878, 16'd1937, 16'd15085, 16'd2010, 16'd19087, 16'd58684, 16'd59418, 16'd50241, 16'd64007, 16'd14181, 16'd6719, 16'd13677, 16'd65501, 16'd51862, 16'd58105, 16'd36892, 16'd54839, 16'd39716, 16'd6838, 16'd63134, 16'd16726, 16'd45617, 16'd12712, 16'd21229, 16'd16993});
	test_expansion(128'h0e66341950d63f14083bc53e9b3a2cc6, {16'd269, 16'd54468, 16'd31582, 16'd22252, 16'd14806, 16'd50045, 16'd64911, 16'd65422, 16'd18985, 16'd21463, 16'd8529, 16'd3594, 16'd7560, 16'd26267, 16'd30706, 16'd42466, 16'd29618, 16'd58437, 16'd15199, 16'd19840, 16'd27053, 16'd49045, 16'd470, 16'd62016, 16'd26342, 16'd1027});
	test_expansion(128'h50fcfc268983211a2c2e9a1976da847a, {16'd41593, 16'd11676, 16'd37712, 16'd20288, 16'd28801, 16'd5639, 16'd34880, 16'd64083, 16'd48749, 16'd2715, 16'd22636, 16'd52871, 16'd5595, 16'd5848, 16'd25623, 16'd57867, 16'd23818, 16'd52934, 16'd12171, 16'd21461, 16'd44526, 16'd9606, 16'd32267, 16'd39253, 16'd31332, 16'd10664});
	test_expansion(128'hbea1d16415d803a7439d325d7e713487, {16'd42526, 16'd2976, 16'd3430, 16'd16260, 16'd19403, 16'd56710, 16'd52023, 16'd716, 16'd22993, 16'd19583, 16'd60009, 16'd58799, 16'd19126, 16'd41779, 16'd52368, 16'd962, 16'd62006, 16'd12343, 16'd52756, 16'd54623, 16'd45833, 16'd44157, 16'd19901, 16'd60598, 16'd63894, 16'd117});
	test_expansion(128'h920dada8943f014085cdd64752d27db8, {16'd49640, 16'd24376, 16'd30814, 16'd10972, 16'd55866, 16'd28827, 16'd31202, 16'd44393, 16'd49940, 16'd38593, 16'd4464, 16'd9342, 16'd36421, 16'd981, 16'd57833, 16'd24158, 16'd3094, 16'd22292, 16'd54199, 16'd19053, 16'd59819, 16'd19599, 16'd26593, 16'd53390, 16'd22571, 16'd17361});
	test_expansion(128'h028bbcf18d659a138b70cfb028cb09e1, {16'd9574, 16'd43621, 16'd21860, 16'd61202, 16'd43572, 16'd52822, 16'd51578, 16'd946, 16'd51432, 16'd44989, 16'd11795, 16'd53336, 16'd36023, 16'd9025, 16'd3629, 16'd52792, 16'd17510, 16'd32814, 16'd35432, 16'd28280, 16'd40040, 16'd20400, 16'd20407, 16'd31147, 16'd18089, 16'd15756});
	test_expansion(128'hf724253cac72bdf13fb11ae1c78d7cde, {16'd16434, 16'd56545, 16'd61686, 16'd56893, 16'd7739, 16'd44639, 16'd46992, 16'd22893, 16'd63445, 16'd15389, 16'd23773, 16'd14531, 16'd30084, 16'd47393, 16'd42513, 16'd44824, 16'd60609, 16'd61913, 16'd57320, 16'd521, 16'd45233, 16'd23341, 16'd4719, 16'd13507, 16'd5926, 16'd43120});
	test_expansion(128'hd5ce037f237216ff373bfa2886dcf73b, {16'd20356, 16'd8562, 16'd29202, 16'd15467, 16'd19020, 16'd18125, 16'd7687, 16'd31221, 16'd20250, 16'd60224, 16'd59645, 16'd52134, 16'd18552, 16'd49472, 16'd42629, 16'd64026, 16'd49168, 16'd5912, 16'd4768, 16'd43980, 16'd4056, 16'd46986, 16'd47313, 16'd9436, 16'd42293, 16'd20201});
	test_expansion(128'ha76670bdf40d4ce27f8514c519b91d8c, {16'd37561, 16'd14606, 16'd15073, 16'd34511, 16'd28773, 16'd40349, 16'd10624, 16'd55386, 16'd9889, 16'd11638, 16'd32149, 16'd22410, 16'd26049, 16'd30605, 16'd42142, 16'd21711, 16'd336, 16'd21741, 16'd22568, 16'd33581, 16'd42316, 16'd5292, 16'd38615, 16'd11107, 16'd11991, 16'd49772});
	test_expansion(128'h069cdef6e92020fc1b6a0b09bdbf2d77, {16'd43555, 16'd47392, 16'd10217, 16'd24464, 16'd36071, 16'd14509, 16'd43485, 16'd36523, 16'd47677, 16'd39156, 16'd45100, 16'd11882, 16'd64742, 16'd51028, 16'd2781, 16'd57239, 16'd23541, 16'd17365, 16'd55099, 16'd6633, 16'd37304, 16'd9740, 16'd36757, 16'd14652, 16'd16688, 16'd5664});
	test_expansion(128'h5f8a62c3623545565714870b75559b41, {16'd40883, 16'd51721, 16'd58994, 16'd32548, 16'd8218, 16'd18015, 16'd4504, 16'd58899, 16'd53919, 16'd15191, 16'd29008, 16'd11641, 16'd13863, 16'd41138, 16'd35138, 16'd28343, 16'd35319, 16'd22024, 16'd39244, 16'd5209, 16'd63323, 16'd12820, 16'd15944, 16'd16012, 16'd29879, 16'd55313});
	test_expansion(128'h859fc247d97ad5bbf8b23321b536f96c, {16'd51611, 16'd24418, 16'd47567, 16'd40213, 16'd59012, 16'd8558, 16'd48508, 16'd26108, 16'd36099, 16'd31772, 16'd32187, 16'd24344, 16'd43727, 16'd7237, 16'd45493, 16'd11235, 16'd43493, 16'd27590, 16'd32435, 16'd3888, 16'd21967, 16'd61108, 16'd17179, 16'd33804, 16'd55730, 16'd31142});
	test_expansion(128'hc7dfb5e81647e3bde893fe90e97615aa, {16'd53929, 16'd24559, 16'd15318, 16'd30027, 16'd55697, 16'd44308, 16'd50328, 16'd2651, 16'd7805, 16'd1514, 16'd53328, 16'd4068, 16'd57943, 16'd54787, 16'd57360, 16'd37341, 16'd57062, 16'd36677, 16'd47633, 16'd43800, 16'd3789, 16'd21453, 16'd6441, 16'd45394, 16'd4029, 16'd52754});
	test_expansion(128'h6729b62046aa8b0b7fa7f3addabaf6f6, {16'd39282, 16'd5979, 16'd4100, 16'd62049, 16'd17395, 16'd14574, 16'd38081, 16'd15529, 16'd10222, 16'd60197, 16'd38395, 16'd8066, 16'd34890, 16'd56911, 16'd42322, 16'd20190, 16'd20176, 16'd17895, 16'd1252, 16'd50307, 16'd57299, 16'd270, 16'd16743, 16'd22469, 16'd34315, 16'd51546});
	test_expansion(128'h888628cd27ca02e0e265af81ac4d1a30, {16'd56515, 16'd8305, 16'd18187, 16'd12142, 16'd64524, 16'd39586, 16'd42458, 16'd37570, 16'd5359, 16'd29178, 16'd58920, 16'd36923, 16'd58644, 16'd45433, 16'd4884, 16'd58647, 16'd47944, 16'd13900, 16'd37402, 16'd61489, 16'd17319, 16'd46048, 16'd34478, 16'd53810, 16'd42125, 16'd6610});
	test_expansion(128'h56a3756aea3f3c68aa2893fd126d9b6a, {16'd24156, 16'd14124, 16'd56969, 16'd40852, 16'd12544, 16'd41399, 16'd23214, 16'd45049, 16'd56271, 16'd53685, 16'd17248, 16'd8735, 16'd64154, 16'd53542, 16'd26877, 16'd64456, 16'd59296, 16'd61585, 16'd34267, 16'd17339, 16'd58055, 16'd33957, 16'd53568, 16'd29199, 16'd6952, 16'd43041});
	test_expansion(128'hfddf6699cd27e53dbcbc89512c3b0f60, {16'd26786, 16'd33961, 16'd12645, 16'd1030, 16'd974, 16'd38265, 16'd29686, 16'd29070, 16'd3603, 16'd53008, 16'd53936, 16'd35376, 16'd34771, 16'd11527, 16'd62755, 16'd26666, 16'd64405, 16'd47527, 16'd22928, 16'd37602, 16'd57405, 16'd8610, 16'd5107, 16'd41844, 16'd62145, 16'd65343});
	test_expansion(128'hb0a045dd420ce5454e8ebb0584c88377, {16'd57766, 16'd54174, 16'd57535, 16'd60694, 16'd44415, 16'd27381, 16'd10534, 16'd37488, 16'd25489, 16'd16429, 16'd48159, 16'd7759, 16'd64910, 16'd12230, 16'd45875, 16'd30512, 16'd423, 16'd7703, 16'd42471, 16'd15684, 16'd8248, 16'd15330, 16'd64250, 16'd51114, 16'd49509, 16'd50276});
	test_expansion(128'h496a1d1df53a0a08f3c9f7a89e92c65e, {16'd3433, 16'd12368, 16'd44352, 16'd22602, 16'd8195, 16'd19326, 16'd45500, 16'd9447, 16'd41850, 16'd7734, 16'd27914, 16'd43090, 16'd51708, 16'd14571, 16'd2362, 16'd24328, 16'd45795, 16'd43982, 16'd12054, 16'd20437, 16'd45646, 16'd39998, 16'd19811, 16'd3924, 16'd58272, 16'd721});
	test_expansion(128'h16fb8d14d894d349632b79cda65aad9e, {16'd54432, 16'd65430, 16'd16614, 16'd40517, 16'd44572, 16'd48975, 16'd12228, 16'd29587, 16'd59559, 16'd39699, 16'd1582, 16'd7896, 16'd45056, 16'd59708, 16'd1925, 16'd2289, 16'd29688, 16'd26219, 16'd3310, 16'd11456, 16'd31251, 16'd1358, 16'd10894, 16'd23644, 16'd58666, 16'd26522});
	test_expansion(128'h206b7742a719d6a4f12b9e46547d6d11, {16'd1076, 16'd55693, 16'd34221, 16'd19004, 16'd60592, 16'd8962, 16'd56835, 16'd25299, 16'd42614, 16'd57281, 16'd31610, 16'd34086, 16'd14524, 16'd60268, 16'd41009, 16'd35128, 16'd39447, 16'd23632, 16'd43517, 16'd35745, 16'd22628, 16'd21124, 16'd5190, 16'd4450, 16'd52700, 16'd35480});
	test_expansion(128'hb21a6979ae7310b26e4fdb01c9834449, {16'd18663, 16'd41653, 16'd837, 16'd58858, 16'd12075, 16'd5493, 16'd60533, 16'd61711, 16'd11403, 16'd43991, 16'd35351, 16'd57661, 16'd60650, 16'd182, 16'd30979, 16'd33679, 16'd22395, 16'd6646, 16'd6955, 16'd38302, 16'd2778, 16'd64720, 16'd41125, 16'd29873, 16'd17481, 16'd26770});
	test_expansion(128'h044be056abfdc64dcea17c19392feb8b, {16'd61739, 16'd53145, 16'd23412, 16'd34258, 16'd48324, 16'd18435, 16'd36506, 16'd46835, 16'd20240, 16'd58077, 16'd18606, 16'd42880, 16'd45197, 16'd16441, 16'd50742, 16'd21520, 16'd9187, 16'd49656, 16'd13563, 16'd40687, 16'd34741, 16'd57796, 16'd25185, 16'd12116, 16'd32102, 16'd54397});
	test_expansion(128'hd55b727abe056295b81a806690cda98e, {16'd8611, 16'd61544, 16'd14562, 16'd32899, 16'd22128, 16'd47352, 16'd52279, 16'd3792, 16'd43360, 16'd54679, 16'd46449, 16'd34535, 16'd42704, 16'd33056, 16'd65052, 16'd55678, 16'd52838, 16'd59, 16'd23168, 16'd62097, 16'd43137, 16'd54426, 16'd30164, 16'd59618, 16'd20074, 16'd8444});
	test_expansion(128'hb01dcaf7a9439ce5bb01186be1db2188, {16'd4909, 16'd37680, 16'd752, 16'd41084, 16'd12391, 16'd57337, 16'd10425, 16'd60286, 16'd14259, 16'd19455, 16'd54196, 16'd10766, 16'd50144, 16'd18681, 16'd31854, 16'd27680, 16'd47235, 16'd11291, 16'd2015, 16'd54418, 16'd52326, 16'd40761, 16'd2452, 16'd32049, 16'd41999, 16'd37773});
	test_expansion(128'h47f48640cf1156f7f7f53f374183398b, {16'd16709, 16'd20298, 16'd49776, 16'd52714, 16'd65229, 16'd8466, 16'd54716, 16'd56038, 16'd30718, 16'd28564, 16'd35301, 16'd36489, 16'd62407, 16'd40500, 16'd4881, 16'd16280, 16'd25571, 16'd54590, 16'd40400, 16'd40298, 16'd37448, 16'd23145, 16'd53987, 16'd20170, 16'd59924, 16'd4797});
	test_expansion(128'hca02030689e3693caf7ad5d6695aadd9, {16'd56702, 16'd50805, 16'd40545, 16'd4403, 16'd48442, 16'd27834, 16'd41250, 16'd4185, 16'd46320, 16'd57428, 16'd45077, 16'd15854, 16'd28251, 16'd64578, 16'd35203, 16'd64243, 16'd23169, 16'd50373, 16'd8736, 16'd6053, 16'd46815, 16'd48807, 16'd6868, 16'd41178, 16'd44595, 16'd63342});
	test_expansion(128'h611d491181624ffd044e6ca95558fb21, {16'd21268, 16'd51149, 16'd29289, 16'd15080, 16'd64802, 16'd32097, 16'd16283, 16'd21542, 16'd27150, 16'd15765, 16'd27541, 16'd7051, 16'd26089, 16'd41485, 16'd59042, 16'd29962, 16'd37355, 16'd65286, 16'd9550, 16'd14633, 16'd7901, 16'd29289, 16'd51280, 16'd44564, 16'd16793, 16'd24127});
	test_expansion(128'hb99e18ae4b5a80624a41951028c67013, {16'd2664, 16'd45148, 16'd58002, 16'd23362, 16'd55892, 16'd54377, 16'd19378, 16'd50891, 16'd46276, 16'd32507, 16'd101, 16'd48437, 16'd65264, 16'd19157, 16'd52898, 16'd20513, 16'd48107, 16'd14436, 16'd47432, 16'd65277, 16'd38751, 16'd28460, 16'd46909, 16'd2298, 16'd3278, 16'd33769});
	test_expansion(128'h7d2e16ab43a52589b46a67199ba55841, {16'd36967, 16'd16371, 16'd27209, 16'd53723, 16'd13401, 16'd53798, 16'd2416, 16'd9542, 16'd13663, 16'd5859, 16'd39508, 16'd48627, 16'd39595, 16'd15829, 16'd22220, 16'd58, 16'd35724, 16'd50489, 16'd27992, 16'd45227, 16'd21694, 16'd25210, 16'd51473, 16'd63936, 16'd31942, 16'd54202});
	test_expansion(128'h0eb6adaff29934c6f427f101f915a854, {16'd239, 16'd16571, 16'd51008, 16'd25809, 16'd22608, 16'd40031, 16'd443, 16'd47230, 16'd44329, 16'd25620, 16'd46728, 16'd47376, 16'd32876, 16'd37634, 16'd58034, 16'd38007, 16'd45362, 16'd64404, 16'd1350, 16'd17780, 16'd11424, 16'd5035, 16'd6942, 16'd62914, 16'd44538, 16'd52916});
	test_expansion(128'h4f6fd2d4915456f8f7a7a503dc799557, {16'd2285, 16'd20368, 16'd42038, 16'd4332, 16'd4624, 16'd29201, 16'd58478, 16'd27847, 16'd37084, 16'd58297, 16'd31718, 16'd59297, 16'd13810, 16'd3492, 16'd59731, 16'd62484, 16'd22815, 16'd58125, 16'd36377, 16'd23476, 16'd37057, 16'd52669, 16'd13742, 16'd36578, 16'd61113, 16'd41963});
	test_expansion(128'h7f701734c3ce2bc541b63bd75aed5ec5, {16'd57524, 16'd16468, 16'd50452, 16'd50120, 16'd36932, 16'd31493, 16'd26477, 16'd39501, 16'd2600, 16'd5398, 16'd45919, 16'd8323, 16'd30315, 16'd23079, 16'd29921, 16'd33608, 16'd10152, 16'd32795, 16'd64468, 16'd7121, 16'd45454, 16'd54599, 16'd26495, 16'd33953, 16'd61177, 16'd47817});
	test_expansion(128'hfcd3760b0f4be68547507fa1b68519c1, {16'd8902, 16'd59172, 16'd61152, 16'd58188, 16'd23764, 16'd39646, 16'd20778, 16'd13533, 16'd13630, 16'd35835, 16'd60445, 16'd7772, 16'd12168, 16'd12654, 16'd61579, 16'd64297, 16'd55776, 16'd8456, 16'd30852, 16'd5237, 16'd33242, 16'd12981, 16'd45680, 16'd43410, 16'd7136, 16'd37410});
	test_expansion(128'h818bb2a872920aea9760713da553b948, {16'd59275, 16'd23223, 16'd28683, 16'd34773, 16'd57371, 16'd33500, 16'd61845, 16'd40093, 16'd36254, 16'd27369, 16'd11438, 16'd44585, 16'd42627, 16'd27863, 16'd17722, 16'd44861, 16'd40949, 16'd33133, 16'd48067, 16'd9076, 16'd39126, 16'd33269, 16'd47681, 16'd389, 16'd40176, 16'd14132});
	test_expansion(128'h900092a924c1205b400b75e96c0821f0, {16'd55222, 16'd15837, 16'd37463, 16'd12444, 16'd54894, 16'd19695, 16'd17078, 16'd47422, 16'd37333, 16'd34709, 16'd9157, 16'd34250, 16'd49836, 16'd15792, 16'd49518, 16'd31595, 16'd48130, 16'd18144, 16'd21798, 16'd57731, 16'd62246, 16'd54935, 16'd60410, 16'd28511, 16'd25667, 16'd28301});
	test_expansion(128'h46b58035c6a4f882acfe9516b19eef41, {16'd6484, 16'd17436, 16'd8067, 16'd40103, 16'd23031, 16'd6023, 16'd30891, 16'd59100, 16'd5430, 16'd32235, 16'd4273, 16'd39586, 16'd56638, 16'd43251, 16'd20711, 16'd42372, 16'd57168, 16'd35563, 16'd16734, 16'd59380, 16'd63490, 16'd22106, 16'd23079, 16'd50992, 16'd22670, 16'd1526});
	test_expansion(128'h5cca3046ffb8e9e68ab768df4e238ffa, {16'd42683, 16'd45970, 16'd40464, 16'd14706, 16'd45098, 16'd12204, 16'd49124, 16'd4679, 16'd350, 16'd56115, 16'd33054, 16'd50359, 16'd59739, 16'd41375, 16'd24811, 16'd38549, 16'd44720, 16'd38406, 16'd50066, 16'd28213, 16'd4540, 16'd19488, 16'd3162, 16'd39888, 16'd36355, 16'd9239});
	test_expansion(128'hd63ae7f721f7b7f8fd72a7d234821031, {16'd45948, 16'd56261, 16'd32560, 16'd757, 16'd28641, 16'd60785, 16'd5997, 16'd7712, 16'd53710, 16'd41561, 16'd20680, 16'd44718, 16'd10305, 16'd50892, 16'd22708, 16'd63255, 16'd35838, 16'd59841, 16'd117, 16'd11049, 16'd64235, 16'd49475, 16'd48647, 16'd54511, 16'd5038, 16'd46801});
	test_expansion(128'h0bf4b05f10fbd285f80efe6b0ac57a7e, {16'd11708, 16'd20922, 16'd58687, 16'd36722, 16'd5832, 16'd58495, 16'd56794, 16'd54250, 16'd5247, 16'd42573, 16'd44603, 16'd8995, 16'd57633, 16'd16523, 16'd42526, 16'd43248, 16'd59613, 16'd41293, 16'd56618, 16'd49135, 16'd46961, 16'd56552, 16'd13450, 16'd50161, 16'd22185, 16'd43731});
	test_expansion(128'h0ef0d0935f20a4b91f66f016f65b9928, {16'd18103, 16'd17061, 16'd41932, 16'd30052, 16'd37616, 16'd45000, 16'd45763, 16'd20734, 16'd2226, 16'd2823, 16'd51994, 16'd36936, 16'd6784, 16'd51808, 16'd10839, 16'd64478, 16'd2595, 16'd41474, 16'd7854, 16'd26304, 16'd55581, 16'd57297, 16'd48095, 16'd7376, 16'd20455, 16'd44219});
	test_expansion(128'h5a1ac059334b1bdfebe8ef7fe3da8be9, {16'd9125, 16'd59639, 16'd48624, 16'd51357, 16'd40895, 16'd8612, 16'd58106, 16'd26105, 16'd30229, 16'd13153, 16'd30050, 16'd6082, 16'd46075, 16'd6064, 16'd36168, 16'd36267, 16'd63968, 16'd64889, 16'd32475, 16'd26804, 16'd40498, 16'd34104, 16'd18498, 16'd54697, 16'd63318, 16'd3092});
	test_expansion(128'h16711974cfdf9aae26c27c1e12fcb7e6, {16'd9023, 16'd41249, 16'd64198, 16'd47227, 16'd20002, 16'd23567, 16'd16794, 16'd51635, 16'd37991, 16'd53086, 16'd17637, 16'd46843, 16'd14577, 16'd13245, 16'd62778, 16'd4841, 16'd54282, 16'd36293, 16'd7836, 16'd59107, 16'd28621, 16'd42564, 16'd5995, 16'd21682, 16'd40683, 16'd14134});
	test_expansion(128'h969b0dcb9ec37c253fa19a9e8a4203a8, {16'd13505, 16'd14904, 16'd41169, 16'd34510, 16'd10952, 16'd36745, 16'd2148, 16'd39428, 16'd20976, 16'd21415, 16'd29935, 16'd62586, 16'd49341, 16'd56368, 16'd14437, 16'd7486, 16'd34155, 16'd49426, 16'd23414, 16'd5301, 16'd968, 16'd14715, 16'd2722, 16'd37607, 16'd32192, 16'd10433});
	test_expansion(128'h2ca934ed6eb597391ffe5b821868b4da, {16'd40199, 16'd30011, 16'd37232, 16'd19467, 16'd21162, 16'd31166, 16'd47134, 16'd472, 16'd47957, 16'd61743, 16'd2029, 16'd62127, 16'd58951, 16'd5226, 16'd1787, 16'd47980, 16'd37027, 16'd23237, 16'd55374, 16'd43821, 16'd41263, 16'd11413, 16'd23075, 16'd40385, 16'd279, 16'd43995});
	test_expansion(128'hb79cff28f648a18cdf1cac975cd94b8b, {16'd29501, 16'd47903, 16'd53085, 16'd11648, 16'd30542, 16'd16421, 16'd34068, 16'd11267, 16'd48451, 16'd52321, 16'd14088, 16'd61980, 16'd58251, 16'd63369, 16'd59635, 16'd22508, 16'd27568, 16'd63906, 16'd6335, 16'd29212, 16'd56360, 16'd50646, 16'd54167, 16'd63005, 16'd18207, 16'd21007});
	test_expansion(128'h230f89f7f12dce26d9811b57fd4e3c36, {16'd25097, 16'd6993, 16'd49494, 16'd53379, 16'd14633, 16'd34267, 16'd55708, 16'd45359, 16'd45736, 16'd34121, 16'd62028, 16'd24396, 16'd46137, 16'd45387, 16'd37570, 16'd2158, 16'd10275, 16'd42608, 16'd53391, 16'd52004, 16'd51909, 16'd58471, 16'd41492, 16'd49839, 16'd10838, 16'd14635});
	test_expansion(128'h26ad9e5da416516fa6bddeeada31bdd9, {16'd29540, 16'd30794, 16'd2321, 16'd1566, 16'd3194, 16'd26732, 16'd25488, 16'd33880, 16'd35874, 16'd7694, 16'd12736, 16'd51403, 16'd22384, 16'd63221, 16'd61225, 16'd34386, 16'd59566, 16'd9629, 16'd35910, 16'd23449, 16'd24019, 16'd20131, 16'd5523, 16'd61504, 16'd14615, 16'd8167});
	test_expansion(128'h1c08d9e2240498cce3b2221ded7d4c52, {16'd17315, 16'd24125, 16'd19351, 16'd2757, 16'd19000, 16'd43104, 16'd32861, 16'd62610, 16'd36522, 16'd30495, 16'd63190, 16'd9948, 16'd24242, 16'd51990, 16'd31986, 16'd13288, 16'd19368, 16'd63286, 16'd43224, 16'd48266, 16'd16862, 16'd30387, 16'd23496, 16'd10429, 16'd44058, 16'd12081});
	test_expansion(128'h353fc4f93ea24c1d497ae715d2339b35, {16'd46824, 16'd5454, 16'd23600, 16'd21655, 16'd17752, 16'd49124, 16'd55309, 16'd45533, 16'd38844, 16'd61440, 16'd51959, 16'd53126, 16'd54971, 16'd64033, 16'd8031, 16'd8509, 16'd1069, 16'd61319, 16'd57876, 16'd52586, 16'd29577, 16'd45474, 16'd6155, 16'd6309, 16'd81, 16'd16484});
	test_expansion(128'hb086698c39df2ab4d7791cbc18d8c1d3, {16'd3747, 16'd43316, 16'd1445, 16'd65456, 16'd31560, 16'd47306, 16'd59856, 16'd25638, 16'd16811, 16'd45132, 16'd23579, 16'd36297, 16'd11123, 16'd16401, 16'd60221, 16'd16757, 16'd26458, 16'd35431, 16'd52491, 16'd54992, 16'd58586, 16'd18849, 16'd34739, 16'd55811, 16'd10840, 16'd13360});
	test_expansion(128'h1883620ef789dbc409dc57391162a97d, {16'd43003, 16'd4792, 16'd63601, 16'd23607, 16'd20441, 16'd15275, 16'd11514, 16'd26552, 16'd54147, 16'd51932, 16'd44133, 16'd47048, 16'd32136, 16'd55084, 16'd34450, 16'd52812, 16'd3949, 16'd5709, 16'd13718, 16'd47712, 16'd19084, 16'd65434, 16'd41483, 16'd38429, 16'd32378, 16'd45682});
	test_expansion(128'h2fa81c494d03a35b84ac95bd6c58ef29, {16'd55677, 16'd40841, 16'd27559, 16'd18437, 16'd63591, 16'd60383, 16'd35797, 16'd35184, 16'd25237, 16'd55200, 16'd30597, 16'd17879, 16'd22392, 16'd9235, 16'd65444, 16'd62734, 16'd58501, 16'd52474, 16'd48984, 16'd17446, 16'd30334, 16'd35442, 16'd54422, 16'd14464, 16'd62326, 16'd27077});
	test_expansion(128'h00fec83eeab53f950d4cf9b221094930, {16'd53847, 16'd12059, 16'd36779, 16'd35022, 16'd9738, 16'd62231, 16'd25813, 16'd58849, 16'd16572, 16'd11367, 16'd44178, 16'd27101, 16'd27437, 16'd9552, 16'd17669, 16'd18357, 16'd18137, 16'd34329, 16'd59208, 16'd29724, 16'd1943, 16'd28858, 16'd11902, 16'd33847, 16'd65176, 16'd54860});
	test_expansion(128'h9448b7d040640b7e0cf19734680b6239, {16'd32173, 16'd49346, 16'd9240, 16'd43536, 16'd5659, 16'd21528, 16'd12363, 16'd47399, 16'd42165, 16'd1226, 16'd57721, 16'd62248, 16'd56221, 16'd18459, 16'd52954, 16'd60205, 16'd49245, 16'd16855, 16'd36763, 16'd3311, 16'd26926, 16'd62347, 16'd50258, 16'd35447, 16'd50686, 16'd48293});
	test_expansion(128'hc4bb51fe833fa56d825f6257b20d8f42, {16'd19899, 16'd29363, 16'd15911, 16'd22925, 16'd8239, 16'd19309, 16'd45670, 16'd37347, 16'd39465, 16'd49454, 16'd46409, 16'd8416, 16'd9420, 16'd7506, 16'd4641, 16'd29082, 16'd64313, 16'd29029, 16'd4004, 16'd2695, 16'd19288, 16'd29526, 16'd34602, 16'd8760, 16'd12054, 16'd34957});
	test_expansion(128'he2d23e5df8f2ebe6315360c96cbb9a89, {16'd53827, 16'd12370, 16'd25741, 16'd28922, 16'd10300, 16'd25957, 16'd59139, 16'd7371, 16'd5302, 16'd40427, 16'd12800, 16'd51952, 16'd26000, 16'd7823, 16'd58616, 16'd58465, 16'd21322, 16'd10962, 16'd65093, 16'd19499, 16'd64807, 16'd9193, 16'd16664, 16'd6525, 16'd51193, 16'd16953});
	test_expansion(128'h89fa8daf6ea0ed9cc4e93d56fee90839, {16'd52812, 16'd42053, 16'd36948, 16'd34210, 16'd5253, 16'd52628, 16'd56363, 16'd18879, 16'd25743, 16'd4084, 16'd27412, 16'd41995, 16'd53074, 16'd44477, 16'd26356, 16'd19118, 16'd18921, 16'd13595, 16'd24630, 16'd45281, 16'd3850, 16'd55820, 16'd62088, 16'd32296, 16'd31953, 16'd38969});
	test_expansion(128'h55fed30161716a9531a19dbd4364c79e, {16'd56076, 16'd24596, 16'd55784, 16'd9446, 16'd26082, 16'd59967, 16'd22512, 16'd27950, 16'd39307, 16'd42628, 16'd30781, 16'd29288, 16'd51439, 16'd38052, 16'd54059, 16'd36123, 16'd34892, 16'd57217, 16'd24708, 16'd57831, 16'd35257, 16'd17970, 16'd53995, 16'd59790, 16'd62192, 16'd5203});
	test_expansion(128'h1833d3aa1e592473c54816dcd7d1e208, {16'd1396, 16'd4355, 16'd39056, 16'd30540, 16'd55103, 16'd1392, 16'd63950, 16'd5735, 16'd25759, 16'd62563, 16'd24519, 16'd59810, 16'd41511, 16'd15629, 16'd65321, 16'd61676, 16'd53834, 16'd62793, 16'd6472, 16'd32808, 16'd40894, 16'd23749, 16'd28150, 16'd10664, 16'd46198, 16'd7529});
	test_expansion(128'h221a4248935e5936164e3272193141c4, {16'd16723, 16'd41763, 16'd14920, 16'd60506, 16'd25450, 16'd24937, 16'd51785, 16'd52235, 16'd1618, 16'd19936, 16'd35576, 16'd17045, 16'd45415, 16'd1020, 16'd4073, 16'd48984, 16'd4111, 16'd28130, 16'd10925, 16'd21377, 16'd15212, 16'd12520, 16'd52239, 16'd33676, 16'd54553, 16'd28659});
	test_expansion(128'h0a25693da63065362f33687a90b5c603, {16'd4811, 16'd64825, 16'd29726, 16'd55152, 16'd55302, 16'd19442, 16'd25204, 16'd15861, 16'd3634, 16'd63341, 16'd16250, 16'd41105, 16'd37883, 16'd55970, 16'd61692, 16'd35850, 16'd32977, 16'd51430, 16'd53589, 16'd54330, 16'd5226, 16'd16343, 16'd18962, 16'd11507, 16'd6258, 16'd20209});
	test_expansion(128'h8181e50248e90da60c70425067ed00f3, {16'd32029, 16'd41022, 16'd51760, 16'd63326, 16'd21297, 16'd39400, 16'd64948, 16'd32190, 16'd28974, 16'd44007, 16'd45814, 16'd55920, 16'd1180, 16'd32135, 16'd45726, 16'd54539, 16'd32236, 16'd3614, 16'd22603, 16'd14230, 16'd31009, 16'd10101, 16'd38433, 16'd63215, 16'd54655, 16'd64070});
	test_expansion(128'h5894956ab63c51e99f4f5f92424bff17, {16'd12400, 16'd43143, 16'd41038, 16'd64605, 16'd8572, 16'd2159, 16'd19656, 16'd41391, 16'd31356, 16'd59302, 16'd3934, 16'd16755, 16'd51529, 16'd2796, 16'd12153, 16'd11969, 16'd31163, 16'd47036, 16'd3340, 16'd18078, 16'd60760, 16'd21187, 16'd32986, 16'd40568, 16'd3577, 16'd59326});
	test_expansion(128'hd402b68a063e3f47df94a0d980790a23, {16'd38488, 16'd32189, 16'd18932, 16'd4862, 16'd48143, 16'd47673, 16'd3301, 16'd25915, 16'd33216, 16'd45212, 16'd36548, 16'd23832, 16'd43698, 16'd57395, 16'd13091, 16'd627, 16'd22773, 16'd6322, 16'd55394, 16'd8574, 16'd20892, 16'd26942, 16'd22477, 16'd3553, 16'd33092, 16'd7248});
	test_expansion(128'h4daf1f18581afeeac1aa3ea533ee879e, {16'd22444, 16'd62675, 16'd42319, 16'd4726, 16'd22745, 16'd22915, 16'd63927, 16'd30462, 16'd49595, 16'd47585, 16'd59711, 16'd11569, 16'd11521, 16'd17779, 16'd65045, 16'd60514, 16'd54916, 16'd39074, 16'd7064, 16'd35232, 16'd1650, 16'd2605, 16'd48310, 16'd58937, 16'd20358, 16'd19079});
	test_expansion(128'h2bfed9d12bf9555a8c694e444aac6ada, {16'd26266, 16'd58548, 16'd22071, 16'd50536, 16'd20775, 16'd26444, 16'd40486, 16'd3464, 16'd64228, 16'd13465, 16'd8509, 16'd42179, 16'd821, 16'd19809, 16'd27959, 16'd14509, 16'd53550, 16'd59273, 16'd65437, 16'd46282, 16'd54523, 16'd37237, 16'd53094, 16'd41655, 16'd10558, 16'd42101});
	test_expansion(128'h82b1638b24fda77da7b6449d4931bd9e, {16'd9391, 16'd46849, 16'd29164, 16'd37600, 16'd22494, 16'd9520, 16'd19711, 16'd50087, 16'd55782, 16'd19225, 16'd31158, 16'd42857, 16'd48803, 16'd38922, 16'd24239, 16'd3636, 16'd39119, 16'd42523, 16'd40378, 16'd31108, 16'd18233, 16'd52070, 16'd35831, 16'd45686, 16'd18975, 16'd33628});
	test_expansion(128'hd056c3104b0563bf87e66654ba65d87d, {16'd27543, 16'd51456, 16'd37002, 16'd58172, 16'd10425, 16'd26008, 16'd35317, 16'd41935, 16'd5676, 16'd42921, 16'd33678, 16'd65231, 16'd43722, 16'd64433, 16'd12698, 16'd37322, 16'd1444, 16'd57033, 16'd17333, 16'd251, 16'd34086, 16'd63588, 16'd35439, 16'd57795, 16'd28732, 16'd53285});
	test_expansion(128'hf3c20f54d975f57e56857bbc58d41d86, {16'd34848, 16'd14608, 16'd64762, 16'd27270, 16'd32167, 16'd43514, 16'd47497, 16'd47568, 16'd18196, 16'd33455, 16'd898, 16'd41143, 16'd53533, 16'd46529, 16'd17072, 16'd64193, 16'd25147, 16'd18153, 16'd40729, 16'd15773, 16'd30600, 16'd3843, 16'd17160, 16'd59601, 16'd1369, 16'd18103});
	test_expansion(128'hdfb8c5052dfccb65a06e49d6a54ef9cc, {16'd20916, 16'd54721, 16'd13043, 16'd38986, 16'd56272, 16'd7921, 16'd62531, 16'd4767, 16'd63965, 16'd53276, 16'd36958, 16'd54093, 16'd4777, 16'd18537, 16'd4719, 16'd19128, 16'd18025, 16'd63969, 16'd43154, 16'd45181, 16'd45782, 16'd61732, 16'd15947, 16'd8334, 16'd16252, 16'd39931});
	test_expansion(128'h23a08bebb1172f4e4e8762c68123293a, {16'd41639, 16'd39978, 16'd42923, 16'd14939, 16'd23505, 16'd20695, 16'd53411, 16'd59682, 16'd22533, 16'd47317, 16'd22570, 16'd55504, 16'd47782, 16'd33589, 16'd53225, 16'd41006, 16'd43200, 16'd8622, 16'd13725, 16'd18692, 16'd46745, 16'd12583, 16'd24090, 16'd46448, 16'd29791, 16'd5737});
	test_expansion(128'h71ffd54194d708f399392b33f21517c5, {16'd27564, 16'd27975, 16'd60779, 16'd18604, 16'd11747, 16'd19267, 16'd23204, 16'd42904, 16'd4171, 16'd7329, 16'd62258, 16'd14857, 16'd20959, 16'd38652, 16'd28959, 16'd64606, 16'd32421, 16'd16330, 16'd34806, 16'd14447, 16'd4920, 16'd34517, 16'd59882, 16'd33415, 16'd5471, 16'd48383});
	test_expansion(128'h1daa833c2998601b965e8fbc2b309f9a, {16'd3926, 16'd59076, 16'd15632, 16'd14666, 16'd46798, 16'd3694, 16'd6035, 16'd40677, 16'd63738, 16'd23229, 16'd40678, 16'd26433, 16'd15350, 16'd1857, 16'd36023, 16'd25101, 16'd63584, 16'd41412, 16'd216, 16'd18552, 16'd21949, 16'd39343, 16'd11212, 16'd14049, 16'd57477, 16'd52915});
	test_expansion(128'had351855334e8023ad25b2c35031d6b4, {16'd13489, 16'd50842, 16'd45671, 16'd9133, 16'd32388, 16'd28330, 16'd24690, 16'd7756, 16'd25720, 16'd2260, 16'd15937, 16'd61594, 16'd45389, 16'd54124, 16'd24646, 16'd18985, 16'd49097, 16'd58431, 16'd60874, 16'd7340, 16'd36253, 16'd23114, 16'd29317, 16'd60050, 16'd59592, 16'd7197});
	test_expansion(128'h14341e3b2353246b3be4a22f7c19a269, {16'd42488, 16'd26260, 16'd29083, 16'd45528, 16'd45856, 16'd2605, 16'd63329, 16'd38235, 16'd10605, 16'd57227, 16'd55399, 16'd25072, 16'd42897, 16'd39397, 16'd17763, 16'd32808, 16'd13286, 16'd9798, 16'd61231, 16'd53369, 16'd19432, 16'd49148, 16'd32146, 16'd35807, 16'd13561, 16'd239});
	test_expansion(128'h114d7bb570e7b8041b1a9379b58a77a2, {16'd28080, 16'd51897, 16'd15866, 16'd23750, 16'd64362, 16'd53942, 16'd18305, 16'd9095, 16'd43765, 16'd29638, 16'd39016, 16'd27275, 16'd29480, 16'd5963, 16'd63968, 16'd8171, 16'd61622, 16'd50675, 16'd2363, 16'd60290, 16'd55945, 16'd26923, 16'd37145, 16'd6419, 16'd61625, 16'd22761});
	test_expansion(128'h4a8dbf00269161bc5a21bcde8061de99, {16'd26219, 16'd20994, 16'd39076, 16'd5644, 16'd44176, 16'd24476, 16'd497, 16'd32094, 16'd20110, 16'd32193, 16'd44860, 16'd20844, 16'd28085, 16'd29871, 16'd22949, 16'd39002, 16'd64385, 16'd55330, 16'd49339, 16'd51985, 16'd64456, 16'd46532, 16'd18126, 16'd41570, 16'd24427, 16'd20492});
	test_expansion(128'h13e40df7f5d538884f0905203ffed980, {16'd31393, 16'd25102, 16'd4377, 16'd4067, 16'd40132, 16'd58756, 16'd46927, 16'd43982, 16'd60624, 16'd54247, 16'd18679, 16'd41142, 16'd884, 16'd45036, 16'd43032, 16'd13860, 16'd41082, 16'd29568, 16'd37544, 16'd13996, 16'd30611, 16'd6541, 16'd20702, 16'd11845, 16'd14180, 16'd54988});
	test_expansion(128'h1a716bd6dc298836673ff5e0939db08c, {16'd32519, 16'd48177, 16'd12451, 16'd1779, 16'd1356, 16'd51557, 16'd38124, 16'd40066, 16'd61317, 16'd30991, 16'd4526, 16'd6145, 16'd39182, 16'd41714, 16'd25509, 16'd13141, 16'd50042, 16'd874, 16'd7990, 16'd60591, 16'd25278, 16'd14849, 16'd40737, 16'd63795, 16'd41685, 16'd48592});
	test_expansion(128'h8b283616c7c8184b84ec70b1a409eef6, {16'd56167, 16'd19482, 16'd14878, 16'd42359, 16'd37589, 16'd54538, 16'd50536, 16'd61774, 16'd59167, 16'd10582, 16'd14180, 16'd8065, 16'd59353, 16'd62465, 16'd12268, 16'd57546, 16'd1341, 16'd42584, 16'd55525, 16'd2682, 16'd43012, 16'd27916, 16'd54914, 16'd11471, 16'd17682, 16'd4451});
	test_expansion(128'h1230803adc736b01ff7f3ef57638f533, {16'd23694, 16'd3933, 16'd50747, 16'd16471, 16'd20620, 16'd42688, 16'd58307, 16'd59096, 16'd39198, 16'd37501, 16'd28210, 16'd16415, 16'd59911, 16'd42854, 16'd41113, 16'd47811, 16'd52861, 16'd63946, 16'd17295, 16'd64750, 16'd29125, 16'd4835, 16'd18950, 16'd47300, 16'd12009, 16'd35314});
	test_expansion(128'hee7f6ed39397e499e22033d935778b85, {16'd20835, 16'd20542, 16'd29863, 16'd39192, 16'd64393, 16'd26299, 16'd24260, 16'd1779, 16'd28505, 16'd36446, 16'd18300, 16'd47094, 16'd5609, 16'd20489, 16'd23282, 16'd15441, 16'd60045, 16'd14125, 16'd28630, 16'd34966, 16'd4477, 16'd23917, 16'd54644, 16'd52653, 16'd7172, 16'd37854});
	test_expansion(128'h3a8ad3f7b0563bde66f77fbdfb23cd49, {16'd57875, 16'd13075, 16'd35024, 16'd12186, 16'd29252, 16'd57766, 16'd25815, 16'd48275, 16'd40511, 16'd581, 16'd54120, 16'd37248, 16'd40471, 16'd41763, 16'd2699, 16'd49650, 16'd10227, 16'd41358, 16'd22924, 16'd30137, 16'd21190, 16'd54325, 16'd50652, 16'd40165, 16'd28487, 16'd22347});
	test_expansion(128'hda592a8a4e16e3026190f8c73e17003f, {16'd54050, 16'd9018, 16'd3594, 16'd14735, 16'd55172, 16'd21116, 16'd10468, 16'd38870, 16'd62522, 16'd54706, 16'd47358, 16'd26711, 16'd3385, 16'd56998, 16'd64908, 16'd614, 16'd56646, 16'd26664, 16'd28434, 16'd29491, 16'd536, 16'd50253, 16'd40595, 16'd51518, 16'd804, 16'd21511});
	test_expansion(128'hfef01712c2943e9a7f40a691c597d40d, {16'd49984, 16'd21865, 16'd54529, 16'd64143, 16'd8250, 16'd19847, 16'd62393, 16'd15024, 16'd14874, 16'd31690, 16'd59626, 16'd15222, 16'd32760, 16'd48982, 16'd17541, 16'd46345, 16'd1185, 16'd55992, 16'd53224, 16'd53389, 16'd2709, 16'd31041, 16'd11866, 16'd54628, 16'd14486, 16'd59090});
	test_expansion(128'he19bbe389c37bc7ec5c4ae82d8eca24f, {16'd41622, 16'd3726, 16'd22373, 16'd56656, 16'd44541, 16'd34824, 16'd65420, 16'd1652, 16'd26577, 16'd45819, 16'd36071, 16'd35798, 16'd50145, 16'd15963, 16'd35128, 16'd32117, 16'd4160, 16'd18338, 16'd48058, 16'd29545, 16'd36067, 16'd44484, 16'd60862, 16'd35092, 16'd60923, 16'd41684});
	test_expansion(128'h5176a769fbf87e0e22f60f64037bf788, {16'd46902, 16'd23601, 16'd27452, 16'd43697, 16'd7338, 16'd33508, 16'd19071, 16'd30852, 16'd18047, 16'd58098, 16'd58963, 16'd46965, 16'd27603, 16'd4581, 16'd4930, 16'd9179, 16'd40752, 16'd63194, 16'd64593, 16'd3539, 16'd34458, 16'd57231, 16'd26736, 16'd5526, 16'd40306, 16'd52947});
	test_expansion(128'hfb5e1d2e796e491c26430c9faffd0522, {16'd30698, 16'd33976, 16'd38936, 16'd17054, 16'd33730, 16'd42450, 16'd50195, 16'd58502, 16'd51855, 16'd55005, 16'd40042, 16'd53094, 16'd6077, 16'd31911, 16'd59041, 16'd29936, 16'd63577, 16'd55754, 16'd23160, 16'd18468, 16'd38007, 16'd60748, 16'd64480, 16'd51385, 16'd9148, 16'd17314});
	test_expansion(128'h8ad85d049fe5d020a8f2ce5a769b7eb5, {16'd47049, 16'd38378, 16'd52621, 16'd55530, 16'd57833, 16'd47210, 16'd46052, 16'd57749, 16'd55094, 16'd17777, 16'd6822, 16'd7300, 16'd43336, 16'd4192, 16'd37263, 16'd18739, 16'd5632, 16'd28240, 16'd28208, 16'd57259, 16'd52570, 16'd49915, 16'd17219, 16'd54802, 16'd12557, 16'd52331});
	test_expansion(128'h9f779294a24996f664fe71a1f574dd5d, {16'd8835, 16'd22966, 16'd19961, 16'd57563, 16'd44705, 16'd30600, 16'd35562, 16'd3165, 16'd65346, 16'd51691, 16'd65437, 16'd60234, 16'd44807, 16'd24697, 16'd24189, 16'd51500, 16'd29597, 16'd6286, 16'd50189, 16'd38273, 16'd11302, 16'd41361, 16'd52673, 16'd64092, 16'd39671, 16'd18555});
	test_expansion(128'hf00211bfd6d8a87e3476b621abc92202, {16'd59009, 16'd15667, 16'd62848, 16'd17247, 16'd11528, 16'd8373, 16'd36672, 16'd54074, 16'd12731, 16'd49293, 16'd3257, 16'd30173, 16'd60870, 16'd35019, 16'd6005, 16'd30076, 16'd34216, 16'd51457, 16'd52711, 16'd56615, 16'd22196, 16'd59471, 16'd46354, 16'd25927, 16'd21031, 16'd25141});
	test_expansion(128'h00b9ef7c50502e521ea74356e228d0d6, {16'd14846, 16'd37241, 16'd27317, 16'd17123, 16'd10773, 16'd25301, 16'd47761, 16'd53414, 16'd9552, 16'd41382, 16'd48533, 16'd28878, 16'd42572, 16'd52029, 16'd23042, 16'd47325, 16'd61844, 16'd35788, 16'd52570, 16'd45415, 16'd28211, 16'd30394, 16'd47902, 16'd16080, 16'd62458, 16'd40450});
	test_expansion(128'hf9f22ac5ae9fd06d702d9d83a6f59d9f, {16'd63199, 16'd56149, 16'd49641, 16'd6214, 16'd50252, 16'd46066, 16'd11212, 16'd42387, 16'd887, 16'd22872, 16'd26423, 16'd59953, 16'd29484, 16'd37978, 16'd18705, 16'd18119, 16'd56629, 16'd32473, 16'd57000, 16'd16877, 16'd57812, 16'd55357, 16'd30139, 16'd18220, 16'd11471, 16'd41067});
	test_expansion(128'hf6367a6ed3c031ad36ffae93f686a61f, {16'd12200, 16'd55511, 16'd38634, 16'd48990, 16'd45815, 16'd10057, 16'd33800, 16'd24611, 16'd32167, 16'd25407, 16'd61932, 16'd39432, 16'd62331, 16'd62933, 16'd38547, 16'd33658, 16'd6685, 16'd23592, 16'd25510, 16'd22756, 16'd47615, 16'd37866, 16'd35412, 16'd27450, 16'd56768, 16'd27496});
	test_expansion(128'hf71d3b9c00b0c00391fddd056269b1dd, {16'd20648, 16'd6876, 16'd55118, 16'd61537, 16'd64904, 16'd11311, 16'd63491, 16'd17418, 16'd48121, 16'd26355, 16'd25044, 16'd15249, 16'd61178, 16'd53796, 16'd62867, 16'd58520, 16'd10906, 16'd27464, 16'd62139, 16'd58501, 16'd35321, 16'd33243, 16'd58594, 16'd40310, 16'd48300, 16'd27712});
	test_expansion(128'hb3eeb64270847e9527458dd7a2e2180e, {16'd54342, 16'd41107, 16'd30763, 16'd42820, 16'd55547, 16'd10615, 16'd37374, 16'd37114, 16'd61305, 16'd42370, 16'd57628, 16'd29300, 16'd36340, 16'd15053, 16'd64242, 16'd51594, 16'd56411, 16'd63019, 16'd26178, 16'd45279, 16'd42917, 16'd3635, 16'd43792, 16'd40638, 16'd55390, 16'd16642});
	test_expansion(128'h9fa990d88664a3570e9f05e8bd740652, {16'd57615, 16'd55317, 16'd46492, 16'd37153, 16'd22721, 16'd54786, 16'd52905, 16'd57542, 16'd8838, 16'd28231, 16'd48442, 16'd36931, 16'd24547, 16'd36695, 16'd21673, 16'd33135, 16'd22442, 16'd28814, 16'd34321, 16'd23729, 16'd8605, 16'd19981, 16'd44845, 16'd13416, 16'd16456, 16'd52580});
	test_expansion(128'h357f1429a5b223581380fe5015267dd7, {16'd60522, 16'd39229, 16'd59603, 16'd46015, 16'd57131, 16'd51992, 16'd59510, 16'd13527, 16'd55226, 16'd11402, 16'd8611, 16'd29018, 16'd17497, 16'd37005, 16'd10828, 16'd49185, 16'd29136, 16'd4580, 16'd53699, 16'd21844, 16'd54701, 16'd53280, 16'd10020, 16'd13012, 16'd35941, 16'd55877});
	test_expansion(128'h87aa23d8f614d8a99b40652909baf3f1, {16'd42573, 16'd27985, 16'd37916, 16'd26083, 16'd13980, 16'd38481, 16'd17557, 16'd11673, 16'd16317, 16'd36716, 16'd8337, 16'd46779, 16'd3553, 16'd64998, 16'd63372, 16'd61887, 16'd40086, 16'd25353, 16'd42588, 16'd40344, 16'd8332, 16'd21202, 16'd29975, 16'd46023, 16'd916, 16'd38213});
	test_expansion(128'hf9a821a7764285aa35d19cadf47d4a02, {16'd38768, 16'd25176, 16'd47837, 16'd15735, 16'd40481, 16'd60137, 16'd11229, 16'd44633, 16'd3696, 16'd3247, 16'd10769, 16'd50308, 16'd43963, 16'd14444, 16'd295, 16'd28135, 16'd7803, 16'd59594, 16'd16794, 16'd27490, 16'd8331, 16'd48740, 16'd17094, 16'd46826, 16'd5788, 16'd2403});
	test_expansion(128'hcd015781f3937bf7ab54ae44addf9b00, {16'd48933, 16'd58769, 16'd21852, 16'd19369, 16'd24785, 16'd48070, 16'd5428, 16'd10426, 16'd50557, 16'd36003, 16'd34418, 16'd23831, 16'd12309, 16'd49588, 16'd31298, 16'd63514, 16'd30750, 16'd11860, 16'd12760, 16'd33982, 16'd44475, 16'd48692, 16'd64388, 16'd12315, 16'd10083, 16'd47542});
	test_expansion(128'hd6285a42cd022371e48df3ea06ad6499, {16'd54111, 16'd20632, 16'd40487, 16'd40502, 16'd19751, 16'd58704, 16'd58040, 16'd9246, 16'd18674, 16'd2983, 16'd27047, 16'd516, 16'd65425, 16'd24728, 16'd45305, 16'd10570, 16'd47547, 16'd52514, 16'd23538, 16'd52524, 16'd65330, 16'd61429, 16'd225, 16'd62196, 16'd45063, 16'd31381});
	test_expansion(128'h9e174bd838eb22a19fc39e91e62337a8, {16'd20107, 16'd10559, 16'd55120, 16'd12965, 16'd26826, 16'd42346, 16'd64221, 16'd24254, 16'd25434, 16'd43624, 16'd2366, 16'd18860, 16'd15201, 16'd28787, 16'd244, 16'd62924, 16'd10540, 16'd23868, 16'd27980, 16'd15329, 16'd48842, 16'd23191, 16'd11993, 16'd38357, 16'd52971, 16'd61560});
	test_expansion(128'h97b6845371bd379ba9f955a78b9c8d68, {16'd37017, 16'd63498, 16'd48723, 16'd19435, 16'd60929, 16'd50974, 16'd16480, 16'd46960, 16'd42285, 16'd30514, 16'd55988, 16'd46671, 16'd20318, 16'd10207, 16'd32612, 16'd31149, 16'd56993, 16'd63726, 16'd36329, 16'd46614, 16'd22390, 16'd16799, 16'd22564, 16'd34437, 16'd44154, 16'd57562});
	test_expansion(128'hbafb08641ca98253a8fdeb711f7a685a, {16'd29923, 16'd29184, 16'd10230, 16'd50462, 16'd45799, 16'd6284, 16'd32439, 16'd50594, 16'd18985, 16'd23056, 16'd48973, 16'd22820, 16'd59120, 16'd23715, 16'd45991, 16'd37497, 16'd51302, 16'd39298, 16'd55866, 16'd9590, 16'd32709, 16'd45045, 16'd19677, 16'd58736, 16'd37335, 16'd22090});
	test_expansion(128'h4fe156f40811c1e73b98f9a03d521dbc, {16'd32741, 16'd35653, 16'd42454, 16'd61990, 16'd1690, 16'd33644, 16'd28528, 16'd52247, 16'd18468, 16'd48580, 16'd54702, 16'd3697, 16'd65202, 16'd55429, 16'd58682, 16'd49671, 16'd52109, 16'd24160, 16'd52266, 16'd63070, 16'd26667, 16'd34947, 16'd33330, 16'd29378, 16'd44675, 16'd38371});
	test_expansion(128'h445566e2cfef135df7d6cef463774bbc, {16'd23317, 16'd36294, 16'd44976, 16'd9241, 16'd2672, 16'd11358, 16'd29458, 16'd32973, 16'd27297, 16'd5422, 16'd22843, 16'd46078, 16'd44853, 16'd8551, 16'd37923, 16'd57103, 16'd38010, 16'd20301, 16'd41299, 16'd34890, 16'd68, 16'd6326, 16'd29607, 16'd44800, 16'd49885, 16'd9891});
	test_expansion(128'h83439480b38ef542a7267c84cd429b35, {16'd49364, 16'd43477, 16'd3072, 16'd1127, 16'd47032, 16'd33892, 16'd59011, 16'd58693, 16'd42371, 16'd5998, 16'd8910, 16'd56976, 16'd53713, 16'd36345, 16'd42929, 16'd38424, 16'd4386, 16'd14713, 16'd10596, 16'd40388, 16'd63762, 16'd35601, 16'd62004, 16'd51968, 16'd23657, 16'd25974});
	test_expansion(128'h7d24ac2726b7677bccb78e1022a5d988, {16'd18779, 16'd56905, 16'd15247, 16'd49381, 16'd20700, 16'd4372, 16'd58389, 16'd63328, 16'd51689, 16'd42899, 16'd14743, 16'd33340, 16'd48942, 16'd53575, 16'd60569, 16'd59272, 16'd53094, 16'd51296, 16'd4974, 16'd31770, 16'd10032, 16'd7932, 16'd8222, 16'd23077, 16'd52548, 16'd18198});
	test_expansion(128'he22e0f6579e0ce52018dcb1d78f100f5, {16'd56233, 16'd35154, 16'd35198, 16'd49661, 16'd35707, 16'd57782, 16'd25069, 16'd40793, 16'd16028, 16'd57355, 16'd39715, 16'd15272, 16'd44826, 16'd45625, 16'd15460, 16'd759, 16'd4634, 16'd9826, 16'd12054, 16'd20415, 16'd51597, 16'd19483, 16'd17254, 16'd30822, 16'd26257, 16'd43806});
	test_expansion(128'h8259bc52e7cb252913f2c3196566c206, {16'd15504, 16'd45132, 16'd14795, 16'd18434, 16'd18130, 16'd23604, 16'd63164, 16'd17818, 16'd58031, 16'd3454, 16'd11844, 16'd19358, 16'd52029, 16'd48639, 16'd38201, 16'd39361, 16'd5470, 16'd52711, 16'd44473, 16'd34189, 16'd58038, 16'd41830, 16'd48370, 16'd57554, 16'd2103, 16'd37324});
	test_expansion(128'hf5b9231407a5c1978d74dd35b2acdc87, {16'd11683, 16'd53785, 16'd51412, 16'd27856, 16'd31312, 16'd3692, 16'd55578, 16'd31015, 16'd55622, 16'd58983, 16'd31734, 16'd47614, 16'd59190, 16'd9752, 16'd24384, 16'd31297, 16'd13118, 16'd57138, 16'd15909, 16'd51796, 16'd24375, 16'd35441, 16'd43504, 16'd42689, 16'd1138, 16'd24502});
	test_expansion(128'hb02a146669092a577d276d1412e05e96, {16'd18173, 16'd4657, 16'd34326, 16'd49117, 16'd55778, 16'd39686, 16'd25282, 16'd25430, 16'd22398, 16'd7684, 16'd13505, 16'd13155, 16'd53200, 16'd62221, 16'd5535, 16'd26459, 16'd44744, 16'd51338, 16'd47274, 16'd54108, 16'd27258, 16'd28713, 16'd18639, 16'd52646, 16'd25018, 16'd1879});
	test_expansion(128'h6a1211edfd87408cf7f567096bfe62a2, {16'd42796, 16'd54893, 16'd12625, 16'd59276, 16'd57812, 16'd58172, 16'd58441, 16'd10510, 16'd43203, 16'd12417, 16'd7625, 16'd28076, 16'd2696, 16'd53761, 16'd37833, 16'd17316, 16'd12167, 16'd60408, 16'd83, 16'd9334, 16'd56586, 16'd53038, 16'd12108, 16'd58896, 16'd29833, 16'd30430});
	test_expansion(128'h047fe01235e12fd3b9f769f81c46d945, {16'd10075, 16'd8971, 16'd21768, 16'd36174, 16'd2214, 16'd2866, 16'd40709, 16'd47504, 16'd14202, 16'd23587, 16'd46464, 16'd16366, 16'd45193, 16'd46022, 16'd9373, 16'd48358, 16'd23048, 16'd1151, 16'd6488, 16'd56348, 16'd62840, 16'd27142, 16'd50148, 16'd30648, 16'd55444, 16'd35052});
	test_expansion(128'h4e734141a05c0e3e5f66b51467a4c87a, {16'd42055, 16'd30036, 16'd17817, 16'd60191, 16'd25284, 16'd52455, 16'd48285, 16'd27259, 16'd64475, 16'd30841, 16'd53933, 16'd27879, 16'd51997, 16'd56794, 16'd3473, 16'd39361, 16'd24294, 16'd30592, 16'd58126, 16'd55103, 16'd2658, 16'd37881, 16'd46549, 16'd39853, 16'd24027, 16'd11044});
	test_expansion(128'hb76fc69c937cfe752ba2d272c3253ccc, {16'd2532, 16'd9548, 16'd62475, 16'd2854, 16'd41488, 16'd20007, 16'd21560, 16'd5431, 16'd22186, 16'd52159, 16'd25549, 16'd64082, 16'd52499, 16'd17406, 16'd44525, 16'd21139, 16'd65254, 16'd46803, 16'd37142, 16'd25211, 16'd61926, 16'd19621, 16'd52631, 16'd29533, 16'd34686, 16'd18042});
	test_expansion(128'hd7219e1bcd444aa85cf26cdeb06db1ee, {16'd12133, 16'd38007, 16'd61774, 16'd61801, 16'd54280, 16'd45371, 16'd34253, 16'd14783, 16'd14148, 16'd29223, 16'd12551, 16'd57144, 16'd22950, 16'd2194, 16'd52961, 16'd15557, 16'd41179, 16'd26165, 16'd22939, 16'd492, 16'd52326, 16'd3219, 16'd40768, 16'd11645, 16'd22348, 16'd30820});
	test_expansion(128'h6f2877f096f9160f6e56034ae21a04bf, {16'd16126, 16'd25434, 16'd29510, 16'd55088, 16'd51336, 16'd30525, 16'd56962, 16'd11255, 16'd58324, 16'd56651, 16'd21073, 16'd12152, 16'd22244, 16'd8311, 16'd4435, 16'd47162, 16'd38898, 16'd131, 16'd63332, 16'd23421, 16'd34460, 16'd6346, 16'd29657, 16'd26116, 16'd20988, 16'd20573});
	test_expansion(128'h4c7d87a337c1898e72c995898fb61ac3, {16'd42980, 16'd56227, 16'd51020, 16'd60779, 16'd6955, 16'd51368, 16'd23939, 16'd40087, 16'd60750, 16'd9268, 16'd34095, 16'd26669, 16'd18779, 16'd37640, 16'd8178, 16'd47514, 16'd11739, 16'd56196, 16'd49363, 16'd35038, 16'd63116, 16'd43463, 16'd20940, 16'd55889, 16'd2674, 16'd36540});
	test_expansion(128'h25d33c3fb4f1236b40dd1974148411ac, {16'd53312, 16'd46803, 16'd21901, 16'd48552, 16'd52652, 16'd64544, 16'd52297, 16'd43152, 16'd44157, 16'd9908, 16'd46077, 16'd3834, 16'd47140, 16'd45816, 16'd10115, 16'd12574, 16'd61485, 16'd32577, 16'd758, 16'd42022, 16'd9922, 16'd55565, 16'd37830, 16'd17741, 16'd27113, 16'd31391});
	test_expansion(128'h1a8728805bedaba2033815a7af4c0068, {16'd34020, 16'd29934, 16'd21367, 16'd33810, 16'd32671, 16'd20997, 16'd20031, 16'd27994, 16'd11924, 16'd31020, 16'd61656, 16'd21719, 16'd15104, 16'd30822, 16'd32762, 16'd7106, 16'd50479, 16'd28447, 16'd20273, 16'd4335, 16'd31920, 16'd36843, 16'd5632, 16'd22949, 16'd57698, 16'd57594});
	test_expansion(128'h30d38567e59b46de853f2b64efad0391, {16'd11454, 16'd63347, 16'd11640, 16'd2605, 16'd24323, 16'd8218, 16'd3511, 16'd49214, 16'd19811, 16'd43076, 16'd54528, 16'd58088, 16'd35881, 16'd41675, 16'd63696, 16'd27644, 16'd49301, 16'd41582, 16'd55561, 16'd46147, 16'd37867, 16'd1315, 16'd53390, 16'd47569, 16'd43079, 16'd18270});
	test_expansion(128'hd124b438842466487963f6b5e12dd3ef, {16'd2450, 16'd65166, 16'd1989, 16'd32861, 16'd53094, 16'd14911, 16'd36840, 16'd32968, 16'd6360, 16'd14051, 16'd30431, 16'd33368, 16'd862, 16'd15787, 16'd18931, 16'd49298, 16'd16656, 16'd25244, 16'd10076, 16'd44945, 16'd10701, 16'd25250, 16'd58887, 16'd17978, 16'd14750, 16'd8211});
	test_expansion(128'hb5458de398dbc3233205e57a5bc5ecad, {16'd40568, 16'd8703, 16'd34488, 16'd2782, 16'd48540, 16'd41482, 16'd28278, 16'd14520, 16'd56732, 16'd51560, 16'd58843, 16'd4434, 16'd7113, 16'd37067, 16'd19717, 16'd30935, 16'd17481, 16'd59480, 16'd24869, 16'd25856, 16'd28695, 16'd1063, 16'd18933, 16'd60069, 16'd21393, 16'd34084});
	test_expansion(128'hd0cd61acaa04480f9404b809c310dec9, {16'd3129, 16'd25943, 16'd24539, 16'd30882, 16'd42820, 16'd10964, 16'd33965, 16'd40145, 16'd58850, 16'd22789, 16'd50847, 16'd43436, 16'd42980, 16'd35556, 16'd34416, 16'd17825, 16'd26698, 16'd15333, 16'd6843, 16'd3190, 16'd24258, 16'd41358, 16'd53105, 16'd40069, 16'd51278, 16'd61645});
	test_expansion(128'h251e27b83868e4d022c84c7a242efa3c, {16'd54183, 16'd33742, 16'd33802, 16'd13070, 16'd267, 16'd60102, 16'd62085, 16'd46820, 16'd26221, 16'd16531, 16'd46617, 16'd44299, 16'd61269, 16'd49153, 16'd3926, 16'd49549, 16'd25993, 16'd18162, 16'd13848, 16'd49190, 16'd8454, 16'd17551, 16'd14582, 16'd22408, 16'd61871, 16'd8388});
	test_expansion(128'h9920bf46afe64d2a5c41a7208de71139, {16'd44163, 16'd42513, 16'd51394, 16'd64069, 16'd5411, 16'd1643, 16'd40817, 16'd64192, 16'd39413, 16'd57384, 16'd33713, 16'd57974, 16'd46116, 16'd31151, 16'd55772, 16'd37801, 16'd37961, 16'd31719, 16'd32567, 16'd34867, 16'd36142, 16'd6412, 16'd34939, 16'd63439, 16'd41684, 16'd16901});
	test_expansion(128'h3c58963de36d318dc9f320bcf8f32bee, {16'd27193, 16'd54084, 16'd56905, 16'd6791, 16'd4451, 16'd59298, 16'd20197, 16'd64802, 16'd10272, 16'd18226, 16'd24128, 16'd37749, 16'd64797, 16'd2300, 16'd34450, 16'd59983, 16'd28029, 16'd50679, 16'd35479, 16'd57067, 16'd46077, 16'd39506, 16'd41383, 16'd31526, 16'd16018, 16'd5279});
	test_expansion(128'h29380993d3f281d89d3ba3ce09b1bd76, {16'd10165, 16'd12699, 16'd42592, 16'd40007, 16'd51761, 16'd45884, 16'd13250, 16'd35068, 16'd2447, 16'd41871, 16'd61868, 16'd1859, 16'd56472, 16'd8667, 16'd27551, 16'd61380, 16'd6736, 16'd46826, 16'd37803, 16'd46696, 16'd50596, 16'd420, 16'd1530, 16'd11830, 16'd33081, 16'd62884});
	test_expansion(128'hac30758685d69a3d4b03a12d78cf796f, {16'd57689, 16'd55266, 16'd51487, 16'd54979, 16'd39488, 16'd31952, 16'd45288, 16'd63772, 16'd56708, 16'd10345, 16'd846, 16'd31792, 16'd46031, 16'd44990, 16'd5599, 16'd60785, 16'd46665, 16'd64743, 16'd35532, 16'd19824, 16'd53523, 16'd14407, 16'd14372, 16'd38520, 16'd27003, 16'd11650});
	test_expansion(128'h60439a7e5e924d5d251bdb14a72ec9b9, {16'd1705, 16'd7549, 16'd56981, 16'd51958, 16'd2686, 16'd3217, 16'd49354, 16'd30739, 16'd63596, 16'd51069, 16'd22067, 16'd58881, 16'd7882, 16'd48494, 16'd60632, 16'd63897, 16'd25984, 16'd52789, 16'd62278, 16'd20094, 16'd19325, 16'd44004, 16'd13419, 16'd43953, 16'd32070, 16'd1035});
	test_expansion(128'hd78bb3745ecd06fa877ba484c07ffa72, {16'd31047, 16'd11440, 16'd19264, 16'd15719, 16'd37340, 16'd43329, 16'd35202, 16'd57659, 16'd7104, 16'd37167, 16'd1000, 16'd62397, 16'd30345, 16'd25013, 16'd26280, 16'd2683, 16'd56077, 16'd62301, 16'd54381, 16'd28746, 16'd16133, 16'd61469, 16'd60017, 16'd36878, 16'd44488, 16'd36168});
	test_expansion(128'h188527acb3aa5dff1f35526ed42ed211, {16'd47895, 16'd56158, 16'd41867, 16'd49556, 16'd33556, 16'd4463, 16'd42042, 16'd41589, 16'd59040, 16'd60909, 16'd8701, 16'd39760, 16'd28717, 16'd18978, 16'd1533, 16'd55039, 16'd20290, 16'd12114, 16'd42409, 16'd65455, 16'd11194, 16'd23370, 16'd14297, 16'd33582, 16'd63064, 16'd18834});
	test_expansion(128'h4a7409c3922039d70c19ee04f6db5f92, {16'd35833, 16'd12650, 16'd49636, 16'd46970, 16'd55292, 16'd39242, 16'd29988, 16'd17683, 16'd1135, 16'd969, 16'd25616, 16'd22843, 16'd44802, 16'd57302, 16'd53228, 16'd32501, 16'd45226, 16'd48956, 16'd1599, 16'd28330, 16'd3847, 16'd23098, 16'd4385, 16'd12960, 16'd12012, 16'd20899});
	test_expansion(128'h5f2b9b78f23b397424157a78b66776d2, {16'd22004, 16'd3326, 16'd19486, 16'd22478, 16'd11982, 16'd47124, 16'd32040, 16'd21773, 16'd36703, 16'd16866, 16'd31413, 16'd55598, 16'd57709, 16'd46851, 16'd37996, 16'd24661, 16'd65457, 16'd5517, 16'd30420, 16'd13210, 16'd11423, 16'd28833, 16'd33522, 16'd53906, 16'd38515, 16'd31187});
	test_expansion(128'hd4c9b51fb6dea3d04ae4311740e70919, {16'd24564, 16'd50903, 16'd60062, 16'd4400, 16'd48607, 16'd6468, 16'd45397, 16'd21232, 16'd4375, 16'd4194, 16'd4190, 16'd18472, 16'd28412, 16'd17381, 16'd25924, 16'd58783, 16'd32795, 16'd33151, 16'd65452, 16'd33054, 16'd26976, 16'd26981, 16'd63056, 16'd6775, 16'd55067, 16'd28712});
	test_expansion(128'h8c09e3e5ea4a043743337068c3b6c99a, {16'd30705, 16'd13697, 16'd27913, 16'd63986, 16'd57909, 16'd42993, 16'd43488, 16'd59870, 16'd26549, 16'd31236, 16'd49589, 16'd26701, 16'd7873, 16'd20135, 16'd57318, 16'd59462, 16'd50857, 16'd17804, 16'd24561, 16'd64446, 16'd24521, 16'd32074, 16'd50394, 16'd26152, 16'd41752, 16'd14689});
	test_expansion(128'h886b38b5bcbbc08d42071e2e5a89652f, {16'd28574, 16'd16730, 16'd44452, 16'd40080, 16'd61430, 16'd6862, 16'd5190, 16'd23084, 16'd31519, 16'd9582, 16'd58151, 16'd284, 16'd12734, 16'd10704, 16'd2297, 16'd52540, 16'd12403, 16'd32116, 16'd17130, 16'd43832, 16'd39939, 16'd63293, 16'd14201, 16'd3441, 16'd30774, 16'd52372});
	test_expansion(128'h1c8a4714e90acbd714dc96014635c07b, {16'd2582, 16'd17915, 16'd25952, 16'd18466, 16'd54529, 16'd4466, 16'd43528, 16'd17130, 16'd45590, 16'd29552, 16'd8493, 16'd2926, 16'd19241, 16'd59798, 16'd15046, 16'd12271, 16'd24190, 16'd45041, 16'd37699, 16'd63516, 16'd26929, 16'd17062, 16'd2455, 16'd36080, 16'd51516, 16'd19462});
	test_expansion(128'hd44a69694726e5e1fba2bb910a82510a, {16'd49541, 16'd29941, 16'd6428, 16'd34835, 16'd59213, 16'd46219, 16'd32009, 16'd55209, 16'd23258, 16'd31065, 16'd22541, 16'd56034, 16'd6020, 16'd34571, 16'd11046, 16'd11232, 16'd1341, 16'd46403, 16'd7168, 16'd15831, 16'd62356, 16'd30789, 16'd11914, 16'd9986, 16'd33870, 16'd653});
	test_expansion(128'h46b980f6cde587710c594e997b41997c, {16'd24487, 16'd31659, 16'd37390, 16'd42796, 16'd38290, 16'd28534, 16'd50775, 16'd9031, 16'd64497, 16'd57493, 16'd11238, 16'd31280, 16'd38911, 16'd15744, 16'd8969, 16'd43107, 16'd40185, 16'd27004, 16'd24886, 16'd31982, 16'd49342, 16'd7089, 16'd37605, 16'd49332, 16'd17368, 16'd56341});
	test_expansion(128'h599652a5a191fae64fa41333e99237b0, {16'd17170, 16'd43604, 16'd15593, 16'd56198, 16'd3566, 16'd20896, 16'd11939, 16'd23629, 16'd26166, 16'd17273, 16'd7536, 16'd14590, 16'd63861, 16'd57969, 16'd14863, 16'd53676, 16'd51908, 16'd60019, 16'd43882, 16'd52829, 16'd52234, 16'd3928, 16'd38073, 16'd40406, 16'd18340, 16'd60112});
	test_expansion(128'h39b92cf301c2108bf5073d61d9cc7c40, {16'd12292, 16'd52036, 16'd13428, 16'd37914, 16'd64774, 16'd50152, 16'd48075, 16'd14807, 16'd35850, 16'd1047, 16'd21693, 16'd30336, 16'd57446, 16'd4496, 16'd4973, 16'd22276, 16'd55888, 16'd23610, 16'd17701, 16'd49459, 16'd30873, 16'd38124, 16'd751, 16'd642, 16'd63771, 16'd46399});
	test_expansion(128'h8a90f3c3a7e860b47a02ab47cc4f81f1, {16'd2215, 16'd49190, 16'd58301, 16'd43502, 16'd57088, 16'd14211, 16'd24825, 16'd54245, 16'd28708, 16'd40997, 16'd8486, 16'd52100, 16'd46812, 16'd29576, 16'd6267, 16'd58731, 16'd44964, 16'd18457, 16'd38825, 16'd7787, 16'd13989, 16'd29221, 16'd40238, 16'd20011, 16'd20924, 16'd30929});
	test_expansion(128'hdcee5ee6bd6f7cd2ca77f8f5eaf6db5b, {16'd2209, 16'd54717, 16'd4669, 16'd34131, 16'd58050, 16'd61412, 16'd11251, 16'd60237, 16'd21020, 16'd1797, 16'd57480, 16'd2064, 16'd15440, 16'd19472, 16'd46558, 16'd58650, 16'd1977, 16'd15959, 16'd37070, 16'd24666, 16'd39116, 16'd42834, 16'd65511, 16'd48351, 16'd37281, 16'd19906});
	test_expansion(128'hb99b7ec907de5e98baf8ffb895f0c183, {16'd39623, 16'd6732, 16'd13280, 16'd29485, 16'd14588, 16'd14890, 16'd47747, 16'd57219, 16'd13998, 16'd25949, 16'd14420, 16'd5155, 16'd20211, 16'd17184, 16'd11286, 16'd15473, 16'd63484, 16'd51118, 16'd61293, 16'd47327, 16'd29052, 16'd4850, 16'd25460, 16'd23676, 16'd4648, 16'd54179});
	test_expansion(128'ha122246a70cd48632d4edc7a9f95be41, {16'd59843, 16'd58592, 16'd47217, 16'd19244, 16'd36350, 16'd5777, 16'd15247, 16'd55764, 16'd9743, 16'd57542, 16'd43633, 16'd5159, 16'd30053, 16'd43499, 16'd29650, 16'd51332, 16'd23342, 16'd29621, 16'd19351, 16'd21253, 16'd23115, 16'd14317, 16'd10381, 16'd46111, 16'd29486, 16'd63344});
	test_expansion(128'hcd86d0d67c804034cb767a0543e4757c, {16'd5300, 16'd60523, 16'd18658, 16'd58770, 16'd29991, 16'd27586, 16'd5180, 16'd47587, 16'd6507, 16'd39336, 16'd11423, 16'd12293, 16'd35849, 16'd30884, 16'd36083, 16'd15749, 16'd20685, 16'd62350, 16'd62251, 16'd23807, 16'd17541, 16'd60382, 16'd13594, 16'd42565, 16'd20130, 16'd49126});
	test_expansion(128'h7f4e14248bb8bc49518c25a64737e6cc, {16'd209, 16'd49026, 16'd47011, 16'd34886, 16'd60460, 16'd5564, 16'd51167, 16'd12456, 16'd5336, 16'd4099, 16'd55271, 16'd810, 16'd42258, 16'd21094, 16'd21010, 16'd20277, 16'd4947, 16'd9150, 16'd38587, 16'd50567, 16'd46776, 16'd46429, 16'd21923, 16'd40570, 16'd5001, 16'd41175});
	test_expansion(128'h844759904462ab66c57f387cdd2d1b9e, {16'd43203, 16'd53617, 16'd45454, 16'd15193, 16'd5858, 16'd8324, 16'd308, 16'd61734, 16'd65392, 16'd44205, 16'd47256, 16'd43944, 16'd60142, 16'd53113, 16'd46088, 16'd16214, 16'd31978, 16'd49998, 16'd32714, 16'd60823, 16'd57546, 16'd53776, 16'd63297, 16'd6936, 16'd56349, 16'd28782});
	test_expansion(128'h9304cc95952dc2e25fb36f8819f6511e, {16'd54864, 16'd8114, 16'd1026, 16'd22094, 16'd28941, 16'd6890, 16'd29355, 16'd41326, 16'd20337, 16'd62843, 16'd5447, 16'd59758, 16'd43804, 16'd28207, 16'd10806, 16'd21197, 16'd3139, 16'd14118, 16'd23309, 16'd21372, 16'd56667, 16'd56615, 16'd48427, 16'd64813, 16'd35141, 16'd46230});
	test_expansion(128'h1bc6e3b747ddda31d59d9432a687a32c, {16'd65378, 16'd19030, 16'd45867, 16'd30319, 16'd3750, 16'd39876, 16'd50252, 16'd12691, 16'd64129, 16'd16754, 16'd15260, 16'd4064, 16'd32645, 16'd25802, 16'd34385, 16'd52806, 16'd18535, 16'd30293, 16'd8476, 16'd21736, 16'd11371, 16'd45189, 16'd49890, 16'd27817, 16'd44010, 16'd64272});
	test_expansion(128'hcb7a8f860c41d83e2e8df49a523e0429, {16'd19484, 16'd31696, 16'd14643, 16'd62136, 16'd36820, 16'd13195, 16'd33171, 16'd19090, 16'd16660, 16'd19599, 16'd27510, 16'd26172, 16'd54, 16'd27480, 16'd12760, 16'd24659, 16'd50348, 16'd41589, 16'd52648, 16'd34351, 16'd21028, 16'd18424, 16'd28541, 16'd4109, 16'd41695, 16'd19150});
	test_expansion(128'hf73071d6e5f8381542f55845151a3bf0, {16'd25732, 16'd51800, 16'd54047, 16'd36171, 16'd34775, 16'd16911, 16'd64114, 16'd2301, 16'd20550, 16'd64640, 16'd13349, 16'd3424, 16'd26349, 16'd58269, 16'd14721, 16'd35606, 16'd60296, 16'd32156, 16'd37508, 16'd47305, 16'd48591, 16'd60478, 16'd58452, 16'd23777, 16'd7459, 16'd30435});
	test_expansion(128'h3e8b896d6fe8a1bc9b91963214810631, {16'd5805, 16'd4375, 16'd9853, 16'd12848, 16'd24005, 16'd5045, 16'd49729, 16'd52147, 16'd5251, 16'd45764, 16'd4353, 16'd7810, 16'd42246, 16'd50965, 16'd63910, 16'd58734, 16'd37785, 16'd18628, 16'd48049, 16'd40540, 16'd53761, 16'd19037, 16'd55250, 16'd30442, 16'd5724, 16'd18006});
	test_expansion(128'hf7d7d0e7f5073b41251302559954dba5, {16'd40578, 16'd42515, 16'd43270, 16'd18936, 16'd48645, 16'd24549, 16'd31694, 16'd16156, 16'd5518, 16'd49827, 16'd47318, 16'd60474, 16'd2503, 16'd14148, 16'd42168, 16'd17449, 16'd65459, 16'd12103, 16'd64907, 16'd5593, 16'd55317, 16'd13616, 16'd18176, 16'd43211, 16'd6689, 16'd460});
	test_expansion(128'h152de9fe1f3e0a16269180b9e8d403ac, {16'd959, 16'd52010, 16'd20473, 16'd37434, 16'd22290, 16'd35104, 16'd13957, 16'd12111, 16'd49125, 16'd2259, 16'd26009, 16'd25036, 16'd63185, 16'd43573, 16'd4248, 16'd63187, 16'd52230, 16'd7428, 16'd46157, 16'd13005, 16'd49951, 16'd14350, 16'd60455, 16'd6594, 16'd13615, 16'd10677});
	test_expansion(128'h76454fa56208123971550cf59d3c0e19, {16'd44871, 16'd40840, 16'd35461, 16'd48676, 16'd7652, 16'd2356, 16'd15054, 16'd54190, 16'd19048, 16'd17034, 16'd61203, 16'd10009, 16'd5731, 16'd5770, 16'd21149, 16'd6686, 16'd18815, 16'd60713, 16'd11530, 16'd45398, 16'd49431, 16'd22055, 16'd17325, 16'd64415, 16'd33730, 16'd59214});
	test_expansion(128'h8acba7ccc88a13c3f08042377501707f, {16'd4874, 16'd29180, 16'd26320, 16'd26737, 16'd39416, 16'd2743, 16'd29369, 16'd5249, 16'd6507, 16'd15345, 16'd16835, 16'd59442, 16'd48368, 16'd43286, 16'd62384, 16'd55841, 16'd64660, 16'd6013, 16'd59342, 16'd64500, 16'd23444, 16'd12121, 16'd9110, 16'd51216, 16'd17392, 16'd38577});
	test_expansion(128'h7267000be85d0b206d05f9050c73c449, {16'd23812, 16'd21662, 16'd9114, 16'd1700, 16'd25443, 16'd59438, 16'd25021, 16'd12318, 16'd7029, 16'd30534, 16'd51911, 16'd65004, 16'd31319, 16'd923, 16'd18860, 16'd2464, 16'd31908, 16'd13783, 16'd792, 16'd43026, 16'd59835, 16'd32286, 16'd26124, 16'd26662, 16'd32515, 16'd61741});
	test_expansion(128'h78a7747ed87efbf1a8fa5f07047efe27, {16'd58474, 16'd57134, 16'd3699, 16'd23214, 16'd55110, 16'd7629, 16'd16070, 16'd15435, 16'd39486, 16'd6807, 16'd55808, 16'd12026, 16'd24857, 16'd36059, 16'd12253, 16'd33928, 16'd6435, 16'd35692, 16'd38115, 16'd59118, 16'd12951, 16'd45228, 16'd37542, 16'd48061, 16'd46067, 16'd8198});
	test_expansion(128'h77a8c2133790059187911ac139abb7ec, {16'd18818, 16'd28472, 16'd14899, 16'd19332, 16'd39465, 16'd8975, 16'd7714, 16'd20420, 16'd35339, 16'd52684, 16'd57335, 16'd47219, 16'd56665, 16'd16956, 16'd44879, 16'd20388, 16'd30072, 16'd26708, 16'd28510, 16'd45037, 16'd24982, 16'd5739, 16'd17517, 16'd36570, 16'd51252, 16'd19688});
	test_expansion(128'h0eb15583ae94d5be894abf5387855530, {16'd24477, 16'd64572, 16'd13187, 16'd56127, 16'd28698, 16'd44626, 16'd43604, 16'd51494, 16'd51301, 16'd34706, 16'd284, 16'd41731, 16'd11375, 16'd63971, 16'd58444, 16'd17729, 16'd63427, 16'd47923, 16'd25978, 16'd5246, 16'd42276, 16'd20664, 16'd50003, 16'd32537, 16'd39771, 16'd34573});
	test_expansion(128'h348edb327f96214dba09f30046245bc8, {16'd34597, 16'd57200, 16'd46013, 16'd1754, 16'd13182, 16'd7604, 16'd12813, 16'd42158, 16'd38934, 16'd44988, 16'd62560, 16'd39120, 16'd1749, 16'd48689, 16'd55639, 16'd57768, 16'd16866, 16'd38810, 16'd29284, 16'd41650, 16'd62005, 16'd30882, 16'd46585, 16'd33539, 16'd45714, 16'd10887});
	test_expansion(128'h08722a39e40415ea485278c0ad01757b, {16'd45847, 16'd63524, 16'd8419, 16'd59445, 16'd36358, 16'd33359, 16'd46441, 16'd14276, 16'd31756, 16'd13302, 16'd50085, 16'd15587, 16'd52661, 16'd41114, 16'd19674, 16'd46073, 16'd39723, 16'd7109, 16'd11477, 16'd20222, 16'd45431, 16'd55968, 16'd58966, 16'd42234, 16'd28881, 16'd47130});
	test_expansion(128'h2463256b8465738ea43e61626c3a72b3, {16'd61566, 16'd74, 16'd50591, 16'd59162, 16'd29234, 16'd49471, 16'd25738, 16'd16221, 16'd33573, 16'd38440, 16'd63468, 16'd35613, 16'd1015, 16'd10321, 16'd20335, 16'd56334, 16'd4828, 16'd22078, 16'd53308, 16'd53704, 16'd30250, 16'd36769, 16'd17804, 16'd56502, 16'd62909, 16'd40192});
	test_expansion(128'h2d34d97f6cbec6a5bfefc57978b05d7a, {16'd31338, 16'd40176, 16'd4135, 16'd53054, 16'd1335, 16'd44945, 16'd8448, 16'd5161, 16'd55167, 16'd36356, 16'd22921, 16'd3592, 16'd17239, 16'd56969, 16'd29250, 16'd14349, 16'd9043, 16'd4210, 16'd61883, 16'd15135, 16'd17381, 16'd21314, 16'd15295, 16'd64044, 16'd34191, 16'd13357});
	test_expansion(128'h191411783e1b31088f9090bec3781a80, {16'd39753, 16'd31130, 16'd4595, 16'd50877, 16'd57040, 16'd52869, 16'd18250, 16'd9037, 16'd14991, 16'd33924, 16'd42268, 16'd38308, 16'd55222, 16'd28163, 16'd19698, 16'd61964, 16'd945, 16'd61776, 16'd4744, 16'd44324, 16'd39328, 16'd4948, 16'd13020, 16'd61894, 16'd11921, 16'd60936});
	test_expansion(128'h8d1f6eab5cb8b17b3272f6bc156802a0, {16'd7657, 16'd21922, 16'd17542, 16'd26037, 16'd14992, 16'd11266, 16'd54391, 16'd46093, 16'd47239, 16'd12665, 16'd56010, 16'd3904, 16'd62030, 16'd46865, 16'd4160, 16'd45075, 16'd26691, 16'd32879, 16'd6583, 16'd15621, 16'd37459, 16'd28747, 16'd61412, 16'd9973, 16'd21814, 16'd4838});
	test_expansion(128'h41c886bf67293f373b15b3131660a071, {16'd65196, 16'd7665, 16'd13488, 16'd49981, 16'd36778, 16'd54192, 16'd7737, 16'd51918, 16'd56668, 16'd11845, 16'd16967, 16'd50297, 16'd1312, 16'd14152, 16'd1101, 16'd14707, 16'd6619, 16'd18326, 16'd14981, 16'd51707, 16'd32020, 16'd25271, 16'd44063, 16'd28244, 16'd15403, 16'd24180});
	test_expansion(128'hcf7706956895a23f43035cd928b185ee, {16'd18712, 16'd33220, 16'd57859, 16'd9198, 16'd63059, 16'd23260, 16'd1282, 16'd20247, 16'd2436, 16'd63129, 16'd59238, 16'd33427, 16'd35330, 16'd22253, 16'd17170, 16'd7015, 16'd16349, 16'd6353, 16'd57466, 16'd10857, 16'd31898, 16'd2713, 16'd2081, 16'd914, 16'd29364, 16'd18712});
	test_expansion(128'h6cdf5dac9d533c9f5451f447bfd9e295, {16'd13015, 16'd54351, 16'd63397, 16'd5970, 16'd828, 16'd43904, 16'd4803, 16'd61476, 16'd29127, 16'd7239, 16'd23583, 16'd15710, 16'd2773, 16'd45456, 16'd18960, 16'd22654, 16'd42787, 16'd14669, 16'd47124, 16'd15335, 16'd47592, 16'd64677, 16'd42053, 16'd45982, 16'd44988, 16'd3232});
	test_expansion(128'h83a6a9904b011c9fd3603222e7b191c0, {16'd44987, 16'd54825, 16'd37297, 16'd48557, 16'd30484, 16'd6237, 16'd61122, 16'd27797, 16'd59861, 16'd63711, 16'd50980, 16'd56623, 16'd37283, 16'd21092, 16'd62571, 16'd64951, 16'd50165, 16'd53057, 16'd1559, 16'd1183, 16'd41386, 16'd16240, 16'd14695, 16'd26915, 16'd47428, 16'd58494});
	test_expansion(128'h4fb34069b904596d03b36d4f9e2c757f, {16'd10465, 16'd44131, 16'd50081, 16'd46763, 16'd22605, 16'd60386, 16'd59947, 16'd43070, 16'd14260, 16'd39594, 16'd32017, 16'd17140, 16'd51761, 16'd35575, 16'd26808, 16'd65023, 16'd41772, 16'd33709, 16'd24479, 16'd49978, 16'd53629, 16'd6665, 16'd51300, 16'd4350, 16'd344, 16'd1828});
	test_expansion(128'hb8b20726eb4511bf94f341cb52bb2eef, {16'd30411, 16'd9842, 16'd17106, 16'd60168, 16'd41429, 16'd64263, 16'd5496, 16'd25680, 16'd42999, 16'd30467, 16'd58694, 16'd60199, 16'd33119, 16'd26139, 16'd39207, 16'd54430, 16'd59122, 16'd37012, 16'd20137, 16'd63163, 16'd34918, 16'd63321, 16'd15732, 16'd38969, 16'd32069, 16'd34917});
	test_expansion(128'h4639c714a823621fc3ec468f8cd1824a, {16'd19109, 16'd9087, 16'd12993, 16'd28821, 16'd2177, 16'd28921, 16'd39963, 16'd16528, 16'd12309, 16'd21840, 16'd53395, 16'd16110, 16'd15775, 16'd31195, 16'd34392, 16'd16035, 16'd28672, 16'd58626, 16'd29231, 16'd775, 16'd33147, 16'd32655, 16'd10375, 16'd25950, 16'd53923, 16'd7869});
	test_expansion(128'h9f4470bec60ee679d5e3f23216276b3d, {16'd29221, 16'd65522, 16'd54515, 16'd6292, 16'd32071, 16'd43186, 16'd18761, 16'd5902, 16'd55364, 16'd41451, 16'd53983, 16'd5009, 16'd1252, 16'd2326, 16'd10593, 16'd27226, 16'd52160, 16'd24901, 16'd54428, 16'd10528, 16'd52775, 16'd15158, 16'd36780, 16'd16689, 16'd59437, 16'd21133});
	test_expansion(128'h4838a97d2dea626e76b9fd188cddec15, {16'd34106, 16'd30800, 16'd51094, 16'd46738, 16'd64129, 16'd51293, 16'd27958, 16'd12200, 16'd4494, 16'd56456, 16'd62495, 16'd55599, 16'd16400, 16'd40288, 16'd2794, 16'd26699, 16'd22571, 16'd39357, 16'd23303, 16'd40226, 16'd35990, 16'd18497, 16'd13644, 16'd11458, 16'd18202, 16'd44006});
	test_expansion(128'he122eb2f3de44d6461149fd81e915e48, {16'd6743, 16'd13261, 16'd4017, 16'd4968, 16'd64377, 16'd54815, 16'd55321, 16'd5474, 16'd24646, 16'd47379, 16'd11912, 16'd39201, 16'd6176, 16'd44208, 16'd27534, 16'd48278, 16'd35835, 16'd6607, 16'd6184, 16'd49115, 16'd59202, 16'd58258, 16'd62618, 16'd29989, 16'd37, 16'd43643});
	test_expansion(128'hf8257c36af7044b9c9ff09a3f3c1e3ca, {16'd42360, 16'd61129, 16'd64221, 16'd47317, 16'd58267, 16'd10023, 16'd29298, 16'd8354, 16'd12835, 16'd54440, 16'd52267, 16'd50862, 16'd59143, 16'd1613, 16'd39452, 16'd54590, 16'd65240, 16'd55667, 16'd15795, 16'd61428, 16'd65330, 16'd8379, 16'd38717, 16'd4953, 16'd10163, 16'd46557});
	test_expansion(128'ha9d44d8a642789f56bc5dea7575768a6, {16'd9942, 16'd26359, 16'd31721, 16'd52141, 16'd11431, 16'd16481, 16'd55912, 16'd60570, 16'd10885, 16'd15661, 16'd56848, 16'd18267, 16'd65106, 16'd11544, 16'd47288, 16'd48615, 16'd1207, 16'd63613, 16'd29337, 16'd30305, 16'd52309, 16'd40658, 16'd48070, 16'd14585, 16'd24726, 16'd51872});
	test_expansion(128'hfde83215e3c65963017c36270b22bb49, {16'd46545, 16'd13410, 16'd10458, 16'd35399, 16'd10860, 16'd35883, 16'd11316, 16'd11700, 16'd55060, 16'd228, 16'd59768, 16'd28844, 16'd40149, 16'd49227, 16'd6791, 16'd50970, 16'd35857, 16'd2804, 16'd52698, 16'd49524, 16'd29033, 16'd24040, 16'd46348, 16'd26686, 16'd13454, 16'd62110});
	test_expansion(128'h84d626371c4dbd514775adcfd89b48e2, {16'd60458, 16'd43381, 16'd51778, 16'd59224, 16'd21937, 16'd51805, 16'd15422, 16'd33593, 16'd16320, 16'd64763, 16'd1959, 16'd11524, 16'd55381, 16'd64649, 16'd26453, 16'd6991, 16'd41442, 16'd41109, 16'd60317, 16'd45392, 16'd24563, 16'd35111, 16'd51322, 16'd65134, 16'd43513, 16'd24679});
	test_expansion(128'h7f616dba1e043b0cd3f61ddc0e4a1493, {16'd48925, 16'd38300, 16'd21849, 16'd1081, 16'd21584, 16'd2877, 16'd42425, 16'd1422, 16'd28738, 16'd63223, 16'd56968, 16'd32569, 16'd29255, 16'd63423, 16'd32699, 16'd16233, 16'd2511, 16'd21903, 16'd60889, 16'd40153, 16'd64128, 16'd61937, 16'd55776, 16'd57606, 16'd17114, 16'd57228});
	test_expansion(128'h5a4072b9cd218763e176714b51a48067, {16'd20901, 16'd7736, 16'd37457, 16'd15730, 16'd39581, 16'd35137, 16'd18988, 16'd4776, 16'd51186, 16'd50834, 16'd17792, 16'd5763, 16'd8457, 16'd51831, 16'd10033, 16'd41704, 16'd34841, 16'd39321, 16'd57818, 16'd18450, 16'd10812, 16'd10507, 16'd40025, 16'd56529, 16'd46902, 16'd43168});
	test_expansion(128'hc6ab672ef94475cf2f6e4013eb8b9a20, {16'd40548, 16'd16099, 16'd21503, 16'd28292, 16'd12924, 16'd18702, 16'd56157, 16'd4765, 16'd27668, 16'd9744, 16'd56946, 16'd14107, 16'd60230, 16'd51807, 16'd28046, 16'd61848, 16'd15844, 16'd6345, 16'd5410, 16'd11721, 16'd8748, 16'd25125, 16'd57223, 16'd48108, 16'd59827, 16'd1831});
	test_expansion(128'h34196e4d5f2819124e48f16603319acc, {16'd11416, 16'd28588, 16'd12453, 16'd40740, 16'd16937, 16'd60041, 16'd31254, 16'd41099, 16'd39512, 16'd38949, 16'd519, 16'd30741, 16'd40210, 16'd14376, 16'd19066, 16'd21320, 16'd17487, 16'd18540, 16'd20238, 16'd57613, 16'd35425, 16'd13127, 16'd52241, 16'd33587, 16'd2192, 16'd16451});
	test_expansion(128'h165d02e6a8d51a0f7b58a5ec09aa47ce, {16'd58273, 16'd57773, 16'd25081, 16'd54080, 16'd23533, 16'd58484, 16'd31190, 16'd24792, 16'd40638, 16'd26124, 16'd25271, 16'd43188, 16'd61116, 16'd34713, 16'd41444, 16'd17285, 16'd25776, 16'd56812, 16'd8707, 16'd55759, 16'd57566, 16'd6104, 16'd46955, 16'd32761, 16'd64203, 16'd57966});
	test_expansion(128'h67cc77a6464e4bd6bd5fcb6538a46236, {16'd27011, 16'd63814, 16'd63697, 16'd1061, 16'd65198, 16'd43438, 16'd12551, 16'd47913, 16'd35730, 16'd60917, 16'd40611, 16'd47206, 16'd8447, 16'd61660, 16'd23003, 16'd2243, 16'd33064, 16'd38851, 16'd2871, 16'd40810, 16'd58792, 16'd15452, 16'd42193, 16'd50454, 16'd38920, 16'd40220});
	test_expansion(128'habe6e419ca5860e9b7f473b93b45d57b, {16'd26238, 16'd30518, 16'd18054, 16'd60509, 16'd25330, 16'd51524, 16'd16683, 16'd9671, 16'd12433, 16'd41125, 16'd51450, 16'd10509, 16'd18048, 16'd62370, 16'd14367, 16'd63412, 16'd54302, 16'd19557, 16'd53284, 16'd52436, 16'd6260, 16'd34806, 16'd60309, 16'd45193, 16'd21256, 16'd23078});
	test_expansion(128'h645894727dceddfe54c6cdec592e0d83, {16'd25580, 16'd31458, 16'd56984, 16'd42003, 16'd64515, 16'd35471, 16'd23804, 16'd25787, 16'd24611, 16'd53644, 16'd6548, 16'd27257, 16'd39132, 16'd10894, 16'd31742, 16'd22996, 16'd44876, 16'd13168, 16'd22871, 16'd2146, 16'd38351, 16'd49974, 16'd38789, 16'd4941, 16'd6947, 16'd10015});
	test_expansion(128'hd5256d96c32c78cb50739b5866c0e6e3, {16'd28248, 16'd55633, 16'd33879, 16'd5432, 16'd63788, 16'd45975, 16'd33173, 16'd60450, 16'd8520, 16'd33820, 16'd62686, 16'd15303, 16'd20629, 16'd27787, 16'd49379, 16'd58703, 16'd33264, 16'd32426, 16'd59771, 16'd9707, 16'd30953, 16'd1125, 16'd49084, 16'd37030, 16'd37194, 16'd56081});
	test_expansion(128'h99edcf83918d630bbfb3a471c8dc1041, {16'd17809, 16'd46055, 16'd12861, 16'd55729, 16'd26353, 16'd60300, 16'd22511, 16'd9909, 16'd31363, 16'd42113, 16'd40255, 16'd2565, 16'd49490, 16'd19464, 16'd54433, 16'd28162, 16'd36153, 16'd54585, 16'd15653, 16'd57658, 16'd64020, 16'd197, 16'd397, 16'd59866, 16'd36169, 16'd61073});
	test_expansion(128'hb39e734c766451c304da6fdee7e9ad37, {16'd11640, 16'd21222, 16'd32692, 16'd8718, 16'd36482, 16'd16684, 16'd23954, 16'd19862, 16'd62915, 16'd36976, 16'd40514, 16'd61968, 16'd19935, 16'd21119, 16'd5905, 16'd43541, 16'd63879, 16'd62841, 16'd31791, 16'd12689, 16'd52568, 16'd27836, 16'd61250, 16'd16329, 16'd35397, 16'd4069});
	test_expansion(128'h42313a1d3fbb86b62720bb1b65da57c8, {16'd16611, 16'd49563, 16'd54444, 16'd24994, 16'd55383, 16'd62804, 16'd49337, 16'd62851, 16'd54713, 16'd38709, 16'd18639, 16'd4701, 16'd39527, 16'd18432, 16'd17017, 16'd19554, 16'd5564, 16'd26038, 16'd10790, 16'd43991, 16'd30056, 16'd47313, 16'd18073, 16'd13869, 16'd35943, 16'd61793});
	test_expansion(128'he6b818f0d0d7dcd874d3941bc723c33f, {16'd59877, 16'd45448, 16'd44110, 16'd16145, 16'd13124, 16'd61239, 16'd57887, 16'd55741, 16'd12253, 16'd62647, 16'd49107, 16'd57241, 16'd34225, 16'd55493, 16'd10775, 16'd59369, 16'd5456, 16'd44780, 16'd60476, 16'd51852, 16'd1182, 16'd6066, 16'd52199, 16'd4471, 16'd12843, 16'd4694});
	test_expansion(128'ha6758822a63358c8cf1526a96a03a2a6, {16'd19985, 16'd51357, 16'd54136, 16'd2091, 16'd9317, 16'd54451, 16'd58638, 16'd40052, 16'd24337, 16'd32359, 16'd13257, 16'd32268, 16'd12630, 16'd3177, 16'd61724, 16'd23710, 16'd17181, 16'd47651, 16'd29491, 16'd45527, 16'd3988, 16'd14191, 16'd34701, 16'd52755, 16'd51266, 16'd59500});
	test_expansion(128'h239031f56114a43bf2fcfa74a533f4c6, {16'd59375, 16'd29743, 16'd5972, 16'd6280, 16'd60940, 16'd36576, 16'd6986, 16'd23250, 16'd22905, 16'd33204, 16'd19337, 16'd39167, 16'd65373, 16'd918, 16'd14802, 16'd43844, 16'd8549, 16'd35081, 16'd29702, 16'd61721, 16'd6929, 16'd53887, 16'd34324, 16'd54004, 16'd48474, 16'd56996});
	test_expansion(128'h9ef08439cc7e86db2b4fd5a0046c2ba4, {16'd22699, 16'd54434, 16'd33301, 16'd43578, 16'd27561, 16'd30429, 16'd50451, 16'd21121, 16'd42646, 16'd8039, 16'd64539, 16'd13135, 16'd3606, 16'd55373, 16'd58365, 16'd50376, 16'd40375, 16'd7094, 16'd34380, 16'd43277, 16'd45079, 16'd56982, 16'd61209, 16'd59131, 16'd49487, 16'd41644});
	test_expansion(128'h940cd6cc391681f5598948b6fee7d38b, {16'd27664, 16'd64421, 16'd26653, 16'd53050, 16'd42750, 16'd45057, 16'd40095, 16'd49064, 16'd18928, 16'd54957, 16'd46261, 16'd27001, 16'd52514, 16'd23243, 16'd64013, 16'd3523, 16'd27804, 16'd65174, 16'd18973, 16'd13100, 16'd44849, 16'd21232, 16'd42942, 16'd64078, 16'd41271, 16'd10749});
	test_expansion(128'hfb3de39eac5845b08231e3c1c79069cb, {16'd62104, 16'd40951, 16'd28497, 16'd49518, 16'd13262, 16'd54301, 16'd17065, 16'd8347, 16'd39650, 16'd18313, 16'd18593, 16'd34780, 16'd31660, 16'd41201, 16'd2045, 16'd35979, 16'd24061, 16'd51861, 16'd35918, 16'd37247, 16'd44957, 16'd57349, 16'd38724, 16'd8948, 16'd49132, 16'd44180});
	test_expansion(128'hee9cfeb62df4db740963bd5c90bfedf8, {16'd30530, 16'd29596, 16'd26788, 16'd58300, 16'd17973, 16'd33727, 16'd17312, 16'd19763, 16'd31356, 16'd39723, 16'd39139, 16'd12697, 16'd4891, 16'd32170, 16'd14581, 16'd21755, 16'd51588, 16'd7849, 16'd10770, 16'd13820, 16'd41190, 16'd32834, 16'd60270, 16'd49017, 16'd49559, 16'd3400});
	test_expansion(128'h02d0979609dc7240d43d8244d755f10d, {16'd57342, 16'd36220, 16'd36446, 16'd63572, 16'd23724, 16'd22615, 16'd27350, 16'd35078, 16'd40593, 16'd59780, 16'd64610, 16'd10135, 16'd8304, 16'd59632, 16'd37304, 16'd32589, 16'd47356, 16'd11673, 16'd65189, 16'd35770, 16'd13264, 16'd2521, 16'd42679, 16'd14242, 16'd58325, 16'd30103});
	test_expansion(128'he05595168f331545254f79c47080c80d, {16'd47907, 16'd58990, 16'd17537, 16'd38147, 16'd23166, 16'd24523, 16'd30928, 16'd39982, 16'd30444, 16'd58318, 16'd43168, 16'd51612, 16'd37480, 16'd30584, 16'd41117, 16'd22728, 16'd24743, 16'd63734, 16'd11948, 16'd15503, 16'd64889, 16'd49738, 16'd13970, 16'd439, 16'd43466, 16'd38978});
	test_expansion(128'hbf2c4692e5f178420070c46ec9443810, {16'd56036, 16'd46710, 16'd39056, 16'd62375, 16'd3197, 16'd50839, 16'd34448, 16'd56962, 16'd34847, 16'd15437, 16'd35932, 16'd61968, 16'd16127, 16'd42335, 16'd16791, 16'd49444, 16'd62394, 16'd10423, 16'd42161, 16'd6671, 16'd21277, 16'd6427, 16'd37401, 16'd14604, 16'd14566, 16'd29119});
	test_expansion(128'h7b34a665c3796c8d16dd280d6a9083cb, {16'd57052, 16'd26734, 16'd3217, 16'd43531, 16'd30149, 16'd46789, 16'd36190, 16'd2730, 16'd49367, 16'd54280, 16'd35983, 16'd15766, 16'd62839, 16'd41865, 16'd60728, 16'd34667, 16'd2921, 16'd37013, 16'd35736, 16'd45554, 16'd35781, 16'd8681, 16'd39946, 16'd13137, 16'd48955, 16'd27939});
	test_expansion(128'h1e0a50e5cd24bfcd9f3631587f20b8e2, {16'd27599, 16'd26503, 16'd30822, 16'd5255, 16'd25242, 16'd54903, 16'd15552, 16'd6176, 16'd41951, 16'd15936, 16'd41587, 16'd52223, 16'd57284, 16'd49783, 16'd19553, 16'd9909, 16'd15205, 16'd37346, 16'd63294, 16'd48727, 16'd5840, 16'd25163, 16'd44037, 16'd65479, 16'd26720, 16'd4737});
	test_expansion(128'h0a6dc1d7549dc4aff340b42831fb6b13, {16'd7825, 16'd60799, 16'd3753, 16'd52756, 16'd34453, 16'd35274, 16'd22349, 16'd42657, 16'd57863, 16'd64136, 16'd39384, 16'd12023, 16'd18100, 16'd6748, 16'd25359, 16'd63984, 16'd41675, 16'd32760, 16'd11995, 16'd51862, 16'd47564, 16'd51229, 16'd3931, 16'd63624, 16'd3808, 16'd62392});
	test_expansion(128'h2d348a0ca8aa25e30a86e39ba619331a, {16'd12752, 16'd36120, 16'd36071, 16'd31617, 16'd47838, 16'd30221, 16'd22297, 16'd49110, 16'd36277, 16'd22854, 16'd29456, 16'd64284, 16'd7454, 16'd17194, 16'd41681, 16'd2075, 16'd14077, 16'd43581, 16'd8763, 16'd38953, 16'd43457, 16'd52015, 16'd27791, 16'd41954, 16'd18884, 16'd154});
	test_expansion(128'h488dcde8ef8754a1f6d1449b8f6dfcbf, {16'd47830, 16'd18697, 16'd19209, 16'd20267, 16'd15597, 16'd1568, 16'd37535, 16'd58427, 16'd41411, 16'd30706, 16'd30445, 16'd5462, 16'd16137, 16'd22956, 16'd33558, 16'd46728, 16'd7718, 16'd18389, 16'd9435, 16'd5829, 16'd64268, 16'd19118, 16'd52513, 16'd438, 16'd48665, 16'd62934});
	test_expansion(128'h91ea79fa8a825d52b8426b247dc6efc9, {16'd1728, 16'd2297, 16'd35644, 16'd14850, 16'd26056, 16'd17453, 16'd46717, 16'd50381, 16'd26539, 16'd45784, 16'd21599, 16'd12796, 16'd13387, 16'd55193, 16'd52759, 16'd59989, 16'd43173, 16'd60614, 16'd24251, 16'd33891, 16'd61976, 16'd58792, 16'd34942, 16'd21452, 16'd7569, 16'd49726});
	test_expansion(128'h296250d0fbf717f66046e14f11e6c500, {16'd27374, 16'd917, 16'd59678, 16'd21011, 16'd14993, 16'd25279, 16'd42319, 16'd4636, 16'd45412, 16'd13796, 16'd21859, 16'd55955, 16'd1195, 16'd54289, 16'd15527, 16'd27134, 16'd25531, 16'd62051, 16'd10380, 16'd31853, 16'd10413, 16'd37083, 16'd38955, 16'd27962, 16'd65168, 16'd25166});
	test_expansion(128'h0e28ab3f9bfe89c0e622684c0c86bbc4, {16'd27100, 16'd56066, 16'd9943, 16'd32756, 16'd47816, 16'd7968, 16'd51988, 16'd46233, 16'd4313, 16'd53260, 16'd12466, 16'd45859, 16'd45570, 16'd7202, 16'd3275, 16'd4286, 16'd43557, 16'd26435, 16'd27324, 16'd29368, 16'd22069, 16'd8332, 16'd8100, 16'd22654, 16'd51364, 16'd47852});
	test_expansion(128'h4cad50f17e22c25a54e6fe99b67ae631, {16'd18004, 16'd20273, 16'd15103, 16'd35876, 16'd16984, 16'd27751, 16'd46709, 16'd39795, 16'd12172, 16'd64480, 16'd31152, 16'd3294, 16'd6126, 16'd51326, 16'd10466, 16'd65448, 16'd27933, 16'd17225, 16'd36383, 16'd11081, 16'd6444, 16'd11593, 16'd46877, 16'd46659, 16'd53366, 16'd13413});
	test_expansion(128'h8d428120a42e5a851254aaad91075dcd, {16'd8131, 16'd61200, 16'd64904, 16'd22559, 16'd15208, 16'd36925, 16'd38571, 16'd9745, 16'd6945, 16'd33832, 16'd52756, 16'd49953, 16'd38222, 16'd16872, 16'd43650, 16'd376, 16'd8742, 16'd29530, 16'd43373, 16'd33851, 16'd27435, 16'd31259, 16'd32746, 16'd57802, 16'd39351, 16'd55397});
	test_expansion(128'hbba5991470235d0a01a92af4993491cb, {16'd45389, 16'd19344, 16'd61566, 16'd55741, 16'd11128, 16'd31037, 16'd39734, 16'd56433, 16'd55029, 16'd9913, 16'd47971, 16'd65317, 16'd11382, 16'd34602, 16'd58508, 16'd54737, 16'd50754, 16'd18515, 16'd37358, 16'd42525, 16'd7803, 16'd60720, 16'd54705, 16'd4538, 16'd64920, 16'd24210});
	test_expansion(128'h12c1c21599cd4cb3b0d16c356728264f, {16'd50016, 16'd5092, 16'd10259, 16'd27471, 16'd58079, 16'd27075, 16'd36176, 16'd25561, 16'd49431, 16'd8007, 16'd21722, 16'd52464, 16'd11750, 16'd32538, 16'd42694, 16'd54324, 16'd2771, 16'd24606, 16'd58101, 16'd12738, 16'd1674, 16'd3597, 16'd61014, 16'd35112, 16'd45546, 16'd9907});
	test_expansion(128'hf3a038ac1599e17ddc0a83164a68d749, {16'd39628, 16'd32950, 16'd33673, 16'd16597, 16'd49213, 16'd11877, 16'd9625, 16'd50716, 16'd9669, 16'd45779, 16'd32558, 16'd40169, 16'd14892, 16'd6851, 16'd20551, 16'd29247, 16'd43487, 16'd55747, 16'd42316, 16'd23533, 16'd6817, 16'd32513, 16'd28905, 16'd35603, 16'd23583, 16'd61667});
	test_expansion(128'h993924a92dcb160f073f56a5238801d4, {16'd52247, 16'd26957, 16'd46523, 16'd39301, 16'd51761, 16'd46759, 16'd50981, 16'd38582, 16'd14517, 16'd31520, 16'd19175, 16'd13389, 16'd28948, 16'd8728, 16'd38235, 16'd12860, 16'd13725, 16'd55448, 16'd28934, 16'd27626, 16'd48849, 16'd53609, 16'd27509, 16'd30763, 16'd61941, 16'd505});
	test_expansion(128'h140b1c27c09e7992012b06fc92960da8, {16'd24847, 16'd7870, 16'd35793, 16'd37949, 16'd22094, 16'd181, 16'd26129, 16'd61103, 16'd31969, 16'd61181, 16'd20363, 16'd56473, 16'd9449, 16'd26419, 16'd64636, 16'd15278, 16'd55485, 16'd64246, 16'd45955, 16'd19205, 16'd13643, 16'd53310, 16'd47157, 16'd38331, 16'd30980, 16'd33689});
	test_expansion(128'hd3c8db69c71c9145a6a42cec69dda943, {16'd46230, 16'd42039, 16'd56172, 16'd11412, 16'd41703, 16'd54734, 16'd57181, 16'd633, 16'd50021, 16'd26507, 16'd33375, 16'd44423, 16'd18395, 16'd419, 16'd7964, 16'd31165, 16'd6631, 16'd24037, 16'd31204, 16'd58613, 16'd21367, 16'd15672, 16'd41965, 16'd49921, 16'd16689, 16'd59919});
	test_expansion(128'hd85044793ddd08b1b12dcba51a4050d1, {16'd32760, 16'd19072, 16'd55593, 16'd14323, 16'd42197, 16'd1857, 16'd5588, 16'd29257, 16'd35253, 16'd21265, 16'd50790, 16'd22829, 16'd17207, 16'd11731, 16'd38078, 16'd51857, 16'd29355, 16'd6037, 16'd39812, 16'd41502, 16'd60695, 16'd60161, 16'd28045, 16'd21400, 16'd20907, 16'd62261});
	test_expansion(128'h2f54f117aa3241be5fd0a47956ceabac, {16'd25391, 16'd1066, 16'd58547, 16'd64057, 16'd17354, 16'd40235, 16'd39812, 16'd45616, 16'd198, 16'd23261, 16'd38203, 16'd57482, 16'd56303, 16'd476, 16'd62018, 16'd62442, 16'd28534, 16'd7895, 16'd26896, 16'd60987, 16'd53069, 16'd10834, 16'd55749, 16'd2241, 16'd18738, 16'd49797});
	test_expansion(128'h14cfa768ecebdb80efc0540a527adcf8, {16'd21139, 16'd29383, 16'd45455, 16'd673, 16'd45817, 16'd29381, 16'd18736, 16'd54434, 16'd31534, 16'd51023, 16'd9586, 16'd13666, 16'd54999, 16'd58780, 16'd33028, 16'd10523, 16'd56717, 16'd21168, 16'd50476, 16'd1683, 16'd59604, 16'd64581, 16'd21745, 16'd29984, 16'd2485, 16'd6084});
	test_expansion(128'h096e2449f4a9488e369f5d99967c497e, {16'd63516, 16'd56532, 16'd17594, 16'd47998, 16'd60438, 16'd18498, 16'd27030, 16'd42072, 16'd19186, 16'd60648, 16'd42390, 16'd6343, 16'd64134, 16'd49526, 16'd25991, 16'd16228, 16'd4185, 16'd44183, 16'd37296, 16'd5329, 16'd60210, 16'd24029, 16'd49864, 16'd22962, 16'd22909, 16'd44455});
	test_expansion(128'h56ff1f1eac3213ea000d63431db1aec3, {16'd16385, 16'd12395, 16'd55259, 16'd38128, 16'd26913, 16'd36065, 16'd11072, 16'd17930, 16'd34957, 16'd25198, 16'd65458, 16'd35655, 16'd33140, 16'd17483, 16'd38996, 16'd18643, 16'd59515, 16'd47077, 16'd13185, 16'd42584, 16'd27297, 16'd15043, 16'd43847, 16'd30016, 16'd4158, 16'd34477});
	test_expansion(128'hba7758cf81a1bab44ed605de4d008b36, {16'd38577, 16'd61196, 16'd58332, 16'd46280, 16'd6159, 16'd48418, 16'd54966, 16'd40611, 16'd22605, 16'd17484, 16'd3136, 16'd55603, 16'd55594, 16'd53849, 16'd5049, 16'd53601, 16'd12756, 16'd4935, 16'd21323, 16'd38529, 16'd48946, 16'd27880, 16'd19283, 16'd12166, 16'd59041, 16'd35865});
	test_expansion(128'hfce4d88daf3e03e052b1ccc9ea9f208c, {16'd36423, 16'd8346, 16'd23220, 16'd56063, 16'd58070, 16'd40493, 16'd16140, 16'd48097, 16'd9467, 16'd22529, 16'd32240, 16'd54651, 16'd45379, 16'd49087, 16'd43035, 16'd25469, 16'd26196, 16'd61346, 16'd8241, 16'd52785, 16'd43294, 16'd35850, 16'd12481, 16'd20531, 16'd17757, 16'd31557});
	test_expansion(128'hc1b763e0b85448be96fb83065907697e, {16'd10074, 16'd29101, 16'd32468, 16'd53254, 16'd1203, 16'd60567, 16'd44493, 16'd50406, 16'd29353, 16'd16031, 16'd38029, 16'd9224, 16'd15614, 16'd35851, 16'd58937, 16'd16902, 16'd34828, 16'd2386, 16'd15818, 16'd57006, 16'd28869, 16'd17008, 16'd61028, 16'd17116, 16'd14381, 16'd326});
	test_expansion(128'h7f75bc51cbde054c8c96f09e9c38f941, {16'd64684, 16'd28541, 16'd30128, 16'd55356, 16'd31612, 16'd41013, 16'd51032, 16'd6173, 16'd55965, 16'd24263, 16'd20388, 16'd30619, 16'd8608, 16'd25298, 16'd36066, 16'd63828, 16'd28045, 16'd62503, 16'd14077, 16'd19045, 16'd35354, 16'd35811, 16'd43564, 16'd24898, 16'd61679, 16'd62450});
	test_expansion(128'h21cdcdd2ee45560eb0f1af80c44336fe, {16'd58494, 16'd10635, 16'd5417, 16'd4099, 16'd35644, 16'd27067, 16'd6830, 16'd4452, 16'd13156, 16'd57876, 16'd34249, 16'd60572, 16'd24328, 16'd64008, 16'd54220, 16'd36109, 16'd44271, 16'd50895, 16'd23652, 16'd26119, 16'd31393, 16'd3274, 16'd4805, 16'd29688, 16'd12051, 16'd36702});
	test_expansion(128'hc56692755c2523ae47ee35ad0707a4d7, {16'd13165, 16'd55348, 16'd51600, 16'd39715, 16'd15476, 16'd53944, 16'd816, 16'd41663, 16'd23294, 16'd29244, 16'd30043, 16'd5659, 16'd11332, 16'd51334, 16'd39986, 16'd28298, 16'd48082, 16'd40907, 16'd14153, 16'd53144, 16'd40547, 16'd61809, 16'd21237, 16'd10020, 16'd55352, 16'd5819});
	test_expansion(128'h4eaaea1b08009db89a4cac95e1a3a264, {16'd49022, 16'd12826, 16'd62340, 16'd8199, 16'd55663, 16'd33914, 16'd42616, 16'd53254, 16'd51324, 16'd42041, 16'd40154, 16'd9737, 16'd2413, 16'd60243, 16'd39498, 16'd5251, 16'd13053, 16'd7962, 16'd39326, 16'd58063, 16'd18120, 16'd51101, 16'd35883, 16'd24308, 16'd29157, 16'd53875});
	test_expansion(128'hb884d164b03b1b06d3dc1df6caba6b6f, {16'd50179, 16'd54132, 16'd21875, 16'd55430, 16'd49614, 16'd35170, 16'd33298, 16'd54500, 16'd43679, 16'd37600, 16'd57031, 16'd23633, 16'd47019, 16'd5487, 16'd41678, 16'd4071, 16'd59480, 16'd58039, 16'd3069, 16'd39759, 16'd5816, 16'd65496, 16'd20989, 16'd53502, 16'd44175, 16'd4844});
	test_expansion(128'hf81fac03191f137316fff75186a3ff4e, {16'd22586, 16'd33466, 16'd47249, 16'd23444, 16'd14016, 16'd19441, 16'd24227, 16'd36844, 16'd53628, 16'd25897, 16'd43448, 16'd47974, 16'd20879, 16'd19418, 16'd36807, 16'd8819, 16'd58986, 16'd16113, 16'd61594, 16'd11829, 16'd39456, 16'd63514, 16'd51644, 16'd63500, 16'd63956, 16'd18431});
	test_expansion(128'hfba9467ce53305ac64d2205f49ead0bd, {16'd40424, 16'd34091, 16'd7115, 16'd55667, 16'd59625, 16'd34659, 16'd27583, 16'd60149, 16'd63827, 16'd30611, 16'd18638, 16'd56635, 16'd39291, 16'd14683, 16'd28769, 16'd52053, 16'd22226, 16'd3452, 16'd40429, 16'd35496, 16'd65472, 16'd27865, 16'd58091, 16'd18577, 16'd38655, 16'd13286});
	test_expansion(128'ha8b35a78d376fd6bd35142936b5834a2, {16'd41179, 16'd55034, 16'd64015, 16'd2669, 16'd57671, 16'd59264, 16'd43279, 16'd25464, 16'd6148, 16'd36016, 16'd49938, 16'd46564, 16'd2393, 16'd37543, 16'd45462, 16'd50951, 16'd29413, 16'd56064, 16'd52835, 16'd33464, 16'd8020, 16'd64022, 16'd33725, 16'd57987, 16'd24563, 16'd21180});
	test_expansion(128'hb1a65bdf3d406f489382c87586fb30ed, {16'd3539, 16'd9097, 16'd51160, 16'd29103, 16'd42402, 16'd60512, 16'd54680, 16'd36737, 16'd47162, 16'd32048, 16'd14591, 16'd20352, 16'd21579, 16'd65225, 16'd20422, 16'd63530, 16'd51873, 16'd18697, 16'd37339, 16'd17847, 16'd24003, 16'd51547, 16'd50730, 16'd60078, 16'd19253, 16'd52279});
	test_expansion(128'h5bebd45193fa75131b96b7e82f0b5a22, {16'd46646, 16'd47330, 16'd63598, 16'd29319, 16'd57596, 16'd52831, 16'd16421, 16'd1296, 16'd14367, 16'd12601, 16'd42008, 16'd16426, 16'd7292, 16'd7888, 16'd17732, 16'd54385, 16'd28200, 16'd35943, 16'd35912, 16'd40596, 16'd47941, 16'd13934, 16'd35245, 16'd53532, 16'd53612, 16'd10941});
	test_expansion(128'ha91d2cfa81a3d8e175a4d570485bd36c, {16'd37710, 16'd48373, 16'd62004, 16'd33082, 16'd10687, 16'd61166, 16'd5300, 16'd34194, 16'd64926, 16'd62981, 16'd22492, 16'd42039, 16'd37934, 16'd33563, 16'd38152, 16'd22942, 16'd21948, 16'd50198, 16'd242, 16'd14809, 16'd28426, 16'd33940, 16'd38494, 16'd43182, 16'd37503, 16'd13772});
	test_expansion(128'he710c4a0b77dc7e57c6306f1cf82e42a, {16'd5680, 16'd2924, 16'd50010, 16'd47539, 16'd20082, 16'd11426, 16'd55560, 16'd13987, 16'd458, 16'd46345, 16'd21161, 16'd14299, 16'd33117, 16'd33574, 16'd48986, 16'd6435, 16'd25287, 16'd2654, 16'd35817, 16'd21178, 16'd62211, 16'd33276, 16'd61974, 16'd38767, 16'd55351, 16'd14179});
	test_expansion(128'h65cc9f2e6a998a230c1d4fc92043840c, {16'd20692, 16'd63981, 16'd29305, 16'd2700, 16'd4309, 16'd30053, 16'd20077, 16'd60040, 16'd58652, 16'd32242, 16'd10644, 16'd55161, 16'd16420, 16'd41939, 16'd18983, 16'd15618, 16'd27746, 16'd54573, 16'd40725, 16'd15208, 16'd61931, 16'd39803, 16'd14669, 16'd64847, 16'd10067, 16'd1933});
	test_expansion(128'h6790ac19a23c2c7adad678aa996f32c2, {16'd40774, 16'd50665, 16'd52548, 16'd51854, 16'd18767, 16'd42374, 16'd32816, 16'd62607, 16'd1382, 16'd42272, 16'd53305, 16'd3557, 16'd9028, 16'd11749, 16'd64886, 16'd21883, 16'd20710, 16'd2566, 16'd29536, 16'd60211, 16'd50414, 16'd27937, 16'd30201, 16'd26443, 16'd24857, 16'd32037});
	test_expansion(128'he57626639105126769e0174a0d784f3e, {16'd12904, 16'd36147, 16'd4662, 16'd63553, 16'd22296, 16'd37221, 16'd42439, 16'd412, 16'd5533, 16'd48713, 16'd11489, 16'd7769, 16'd26901, 16'd18362, 16'd28211, 16'd23427, 16'd26822, 16'd47835, 16'd19660, 16'd39920, 16'd63257, 16'd42595, 16'd14177, 16'd64298, 16'd18646, 16'd22098});
	test_expansion(128'hedccc9fd52b190894f97f1df61c1b177, {16'd37730, 16'd5710, 16'd14394, 16'd38744, 16'd56810, 16'd11040, 16'd5065, 16'd18230, 16'd36046, 16'd56167, 16'd62831, 16'd54690, 16'd16723, 16'd44757, 16'd47285, 16'd47655, 16'd8298, 16'd44025, 16'd9155, 16'd60218, 16'd17008, 16'd47229, 16'd4609, 16'd21117, 16'd49039, 16'd20159});
	test_expansion(128'h00287c94c95b746df11e05b64df87dae, {16'd22630, 16'd52947, 16'd17052, 16'd15132, 16'd20392, 16'd36815, 16'd14279, 16'd31455, 16'd52805, 16'd13678, 16'd31313, 16'd18543, 16'd11399, 16'd56663, 16'd19424, 16'd43196, 16'd40743, 16'd64416, 16'd9493, 16'd64727, 16'd60679, 16'd384, 16'd3788, 16'd25122, 16'd6162, 16'd30175});
	test_expansion(128'hb89a78a40472dfb48301ea5236831373, {16'd47276, 16'd12707, 16'd8691, 16'd25382, 16'd65214, 16'd49206, 16'd55369, 16'd27428, 16'd35289, 16'd60529, 16'd64233, 16'd51764, 16'd32228, 16'd47733, 16'd53842, 16'd24950, 16'd56941, 16'd57610, 16'd266, 16'd61482, 16'd27689, 16'd19970, 16'd10502, 16'd54362, 16'd55913, 16'd26629});
	test_expansion(128'h3f60e26f0d78f3065cfbe352105795c0, {16'd2049, 16'd46026, 16'd25562, 16'd32993, 16'd52589, 16'd48357, 16'd23100, 16'd23061, 16'd3717, 16'd28388, 16'd24726, 16'd17481, 16'd43273, 16'd55496, 16'd45147, 16'd6006, 16'd28885, 16'd10157, 16'd58227, 16'd11477, 16'd48927, 16'd15443, 16'd20471, 16'd46315, 16'd2136, 16'd3152});
	test_expansion(128'hc33cab8a43c1c310a364f626876ff911, {16'd24097, 16'd2138, 16'd57753, 16'd17568, 16'd10108, 16'd59685, 16'd60758, 16'd16233, 16'd55554, 16'd18112, 16'd45739, 16'd37529, 16'd19395, 16'd61231, 16'd22780, 16'd8448, 16'd27915, 16'd35982, 16'd44083, 16'd60222, 16'd57265, 16'd26731, 16'd26465, 16'd35156, 16'd61821, 16'd43721});
	test_expansion(128'hbde0c081a3f51b149dc5b162198653e9, {16'd9826, 16'd35586, 16'd1147, 16'd64577, 16'd56322, 16'd35941, 16'd56078, 16'd26317, 16'd39125, 16'd57163, 16'd45571, 16'd24078, 16'd26074, 16'd36351, 16'd20799, 16'd14031, 16'd32707, 16'd59938, 16'd62620, 16'd23493, 16'd60371, 16'd53576, 16'd46318, 16'd8205, 16'd17125, 16'd21048});
	test_expansion(128'hfa4071268afc138345048da2ed1c893d, {16'd13314, 16'd49255, 16'd4451, 16'd13658, 16'd27903, 16'd57760, 16'd46548, 16'd23489, 16'd12556, 16'd34837, 16'd63220, 16'd50845, 16'd51680, 16'd38106, 16'd35244, 16'd47704, 16'd27094, 16'd38237, 16'd8720, 16'd14042, 16'd37547, 16'd18715, 16'd64014, 16'd26648, 16'd20694, 16'd56559});
	test_expansion(128'hdb61dde88de72eda498d7471e6809d1f, {16'd36005, 16'd59252, 16'd23128, 16'd54294, 16'd46049, 16'd3744, 16'd65325, 16'd37260, 16'd58485, 16'd41166, 16'd50170, 16'd64994, 16'd57577, 16'd18638, 16'd54414, 16'd64728, 16'd25564, 16'd29432, 16'd34726, 16'd37710, 16'd43805, 16'd4723, 16'd39927, 16'd12830, 16'd25925, 16'd7938});
	test_expansion(128'hf4e41e9f8ebb706f82a88d78689d04d5, {16'd557, 16'd37039, 16'd23240, 16'd3529, 16'd10629, 16'd54775, 16'd47083, 16'd28503, 16'd31213, 16'd3964, 16'd29456, 16'd32401, 16'd44867, 16'd2190, 16'd61203, 16'd30679, 16'd59464, 16'd8948, 16'd13765, 16'd15703, 16'd16117, 16'd37719, 16'd28846, 16'd48470, 16'd37011, 16'd38269});
	test_expansion(128'h4d55a65c3bc586e2d4fe5fa73711181d, {16'd16089, 16'd22945, 16'd38469, 16'd61071, 16'd16111, 16'd46653, 16'd62021, 16'd42394, 16'd23539, 16'd50333, 16'd12651, 16'd29525, 16'd17954, 16'd43819, 16'd7266, 16'd44611, 16'd61915, 16'd26897, 16'd41423, 16'd21615, 16'd45342, 16'd64105, 16'd45069, 16'd3954, 16'd6291, 16'd41441});
	test_expansion(128'h48e52a0e1ae0c5f33e25692536200393, {16'd46962, 16'd51406, 16'd62402, 16'd38787, 16'd52326, 16'd29427, 16'd47285, 16'd1616, 16'd30382, 16'd12416, 16'd44320, 16'd59209, 16'd30540, 16'd12145, 16'd19012, 16'd34494, 16'd34166, 16'd27708, 16'd48623, 16'd24931, 16'd9157, 16'd58041, 16'd15163, 16'd57172, 16'd46917, 16'd23631});
	test_expansion(128'h3bf1fac81b2f9a6d85ac52bbf72263fd, {16'd10787, 16'd10539, 16'd32694, 16'd17552, 16'd20430, 16'd13908, 16'd18265, 16'd40298, 16'd49264, 16'd26664, 16'd49522, 16'd5430, 16'd23488, 16'd24849, 16'd53868, 16'd24665, 16'd56824, 16'd59970, 16'd20995, 16'd44390, 16'd37665, 16'd53738, 16'd24321, 16'd6694, 16'd16253, 16'd28398});
	test_expansion(128'h1b5a18dc47cd67c379d03d278c83c381, {16'd42569, 16'd46150, 16'd40248, 16'd35066, 16'd60743, 16'd23210, 16'd8338, 16'd44369, 16'd48057, 16'd4811, 16'd37215, 16'd64931, 16'd12164, 16'd57819, 16'd43978, 16'd57901, 16'd42399, 16'd51079, 16'd23830, 16'd29975, 16'd47325, 16'd6281, 16'd13677, 16'd27321, 16'd61753, 16'd39032});
	test_expansion(128'hd02d438fbd866bfd5d8f8e3267a1eb2f, {16'd30326, 16'd43811, 16'd8335, 16'd58098, 16'd33852, 16'd55518, 16'd3013, 16'd11638, 16'd53044, 16'd52345, 16'd18380, 16'd55849, 16'd2361, 16'd29897, 16'd21205, 16'd59908, 16'd30479, 16'd11030, 16'd32774, 16'd37634, 16'd39446, 16'd41928, 16'd54807, 16'd37823, 16'd52974, 16'd62094});
	test_expansion(128'hb73f0a96ce9fdbe88169bb0736194c98, {16'd25739, 16'd12507, 16'd13231, 16'd20060, 16'd13244, 16'd16254, 16'd50323, 16'd14440, 16'd57358, 16'd18452, 16'd59181, 16'd25489, 16'd60561, 16'd41906, 16'd11320, 16'd39972, 16'd34928, 16'd18054, 16'd26478, 16'd11142, 16'd32314, 16'd44366, 16'd58491, 16'd30345, 16'd1323, 16'd979});
	test_expansion(128'h4c713d2b3df540317262141d47ce24b1, {16'd64110, 16'd4129, 16'd57030, 16'd59364, 16'd57883, 16'd49336, 16'd48200, 16'd10515, 16'd11447, 16'd11558, 16'd28206, 16'd36029, 16'd35928, 16'd55648, 16'd51351, 16'd23950, 16'd12656, 16'd20644, 16'd14258, 16'd23464, 16'd30411, 16'd32534, 16'd51065, 16'd50009, 16'd15238, 16'd43729});
	test_expansion(128'h726e2d6e8c0c800e84c15123ac590c99, {16'd8504, 16'd46217, 16'd50276, 16'd23524, 16'd9173, 16'd12126, 16'd57392, 16'd19132, 16'd55183, 16'd14998, 16'd44177, 16'd53184, 16'd21871, 16'd44212, 16'd50675, 16'd27010, 16'd54801, 16'd39493, 16'd30988, 16'd3933, 16'd50833, 16'd43369, 16'd55734, 16'd29868, 16'd40978, 16'd6341});
	test_expansion(128'h446f2cd22850c496cc30bac54e92e8ed, {16'd59302, 16'd23211, 16'd42667, 16'd30522, 16'd37766, 16'd8977, 16'd35633, 16'd47838, 16'd48826, 16'd16989, 16'd56970, 16'd1292, 16'd11151, 16'd14855, 16'd29559, 16'd62810, 16'd1727, 16'd16201, 16'd39268, 16'd48300, 16'd38233, 16'd53500, 16'd56685, 16'd52615, 16'd20188, 16'd52325});
	test_expansion(128'h784619d74e3585bc06cadf672a5c23ff, {16'd64101, 16'd36618, 16'd1955, 16'd18022, 16'd19222, 16'd31378, 16'd36429, 16'd8089, 16'd31858, 16'd40818, 16'd6322, 16'd5286, 16'd15706, 16'd61734, 16'd2646, 16'd56161, 16'd20122, 16'd34623, 16'd471, 16'd45410, 16'd7851, 16'd8956, 16'd18384, 16'd1084, 16'd40973, 16'd57973});
	test_expansion(128'h38f3c7457a19751538f636aadcec8239, {16'd58735, 16'd27249, 16'd17564, 16'd35419, 16'd35821, 16'd19743, 16'd37432, 16'd51453, 16'd32567, 16'd38972, 16'd19011, 16'd32004, 16'd50900, 16'd53484, 16'd32610, 16'd16600, 16'd30343, 16'd35827, 16'd4753, 16'd34419, 16'd42742, 16'd43682, 16'd4839, 16'd30291, 16'd26310, 16'd41823});
	test_expansion(128'he8f25cc6584f4af1acd56c9e049a94a5, {16'd6415, 16'd60019, 16'd37986, 16'd37658, 16'd12851, 16'd7696, 16'd6441, 16'd35269, 16'd44410, 16'd43202, 16'd16732, 16'd23017, 16'd8703, 16'd24718, 16'd31709, 16'd7112, 16'd4435, 16'd13503, 16'd59304, 16'd27594, 16'd36711, 16'd62506, 16'd28208, 16'd46391, 16'd20755, 16'd21801});
	test_expansion(128'h9ccbf5ad7affe28ef459fac13c450542, {16'd56652, 16'd53471, 16'd42028, 16'd52186, 16'd6509, 16'd31412, 16'd22731, 16'd34986, 16'd16851, 16'd805, 16'd41705, 16'd30528, 16'd11387, 16'd14241, 16'd30147, 16'd41473, 16'd27208, 16'd20288, 16'd32008, 16'd12660, 16'd38865, 16'd60486, 16'd22111, 16'd65129, 16'd39457, 16'd55617});
	test_expansion(128'h43716495ac7b24b0f90470c8859d1454, {16'd40305, 16'd61538, 16'd61181, 16'd28048, 16'd59865, 16'd5290, 16'd12976, 16'd14418, 16'd19575, 16'd7112, 16'd14307, 16'd20451, 16'd23850, 16'd64070, 16'd36314, 16'd6715, 16'd12429, 16'd45425, 16'd36452, 16'd47999, 16'd34803, 16'd7944, 16'd19211, 16'd18971, 16'd28321, 16'd36699});
	test_expansion(128'h94a517d3e8299140c8bb3ee1bd2aa5fd, {16'd4242, 16'd54205, 16'd64646, 16'd45568, 16'd34359, 16'd30325, 16'd35296, 16'd61492, 16'd65335, 16'd34706, 16'd10248, 16'd6746, 16'd19180, 16'd31004, 16'd12091, 16'd15939, 16'd27215, 16'd61238, 16'd49738, 16'd36657, 16'd60346, 16'd56347, 16'd1675, 16'd3804, 16'd36416, 16'd52251});
	test_expansion(128'hb358df9855306d078e2fa5b8d3a539f2, {16'd37641, 16'd36154, 16'd37861, 16'd18440, 16'd778, 16'd64791, 16'd37491, 16'd34646, 16'd38567, 16'd42760, 16'd30925, 16'd9808, 16'd47949, 16'd59380, 16'd38499, 16'd60307, 16'd4499, 16'd31568, 16'd35278, 16'd8772, 16'd11845, 16'd13744, 16'd37609, 16'd60829, 16'd11542, 16'd55250});
	test_expansion(128'h6d4454b82b83ea122b1ddecfd7e35a8f, {16'd31701, 16'd12045, 16'd29613, 16'd28506, 16'd34513, 16'd52291, 16'd34265, 16'd32459, 16'd38081, 16'd37332, 16'd35763, 16'd27260, 16'd11678, 16'd29362, 16'd38657, 16'd9748, 16'd15199, 16'd11143, 16'd45841, 16'd10000, 16'd46094, 16'd13481, 16'd62541, 16'd32185, 16'd33106, 16'd39855});
	test_expansion(128'h91dc9c32456cd5350e260429e201c63f, {16'd58407, 16'd56818, 16'd63128, 16'd16653, 16'd17973, 16'd33980, 16'd62442, 16'd46907, 16'd2088, 16'd24905, 16'd60373, 16'd59994, 16'd43965, 16'd34180, 16'd52616, 16'd2880, 16'd8624, 16'd39834, 16'd15386, 16'd11043, 16'd3537, 16'd9309, 16'd116, 16'd4780, 16'd41364, 16'd31414});
	test_expansion(128'h68053b38c28d44263366092395478c31, {16'd25316, 16'd65141, 16'd30499, 16'd17653, 16'd31960, 16'd418, 16'd39017, 16'd20958, 16'd5777, 16'd36989, 16'd11126, 16'd55184, 16'd36435, 16'd38040, 16'd17043, 16'd14906, 16'd27967, 16'd57997, 16'd8353, 16'd52882, 16'd29868, 16'd42136, 16'd42394, 16'd62453, 16'd27982, 16'd53028});
	test_expansion(128'h88334b77581a30550c53b606a8250330, {16'd2137, 16'd40872, 16'd52354, 16'd45400, 16'd30912, 16'd10880, 16'd33245, 16'd14287, 16'd46581, 16'd56997, 16'd59105, 16'd23825, 16'd39610, 16'd25638, 16'd26175, 16'd12431, 16'd49166, 16'd46631, 16'd61734, 16'd31362, 16'd51387, 16'd29458, 16'd57520, 16'd8050, 16'd3706, 16'd16633});
	test_expansion(128'h963080f81e1f20df7f36712ba26cd3bb, {16'd9334, 16'd1781, 16'd34403, 16'd56460, 16'd17834, 16'd46258, 16'd36599, 16'd4730, 16'd5023, 16'd64964, 16'd7795, 16'd23541, 16'd27565, 16'd42400, 16'd33348, 16'd33453, 16'd14878, 16'd32544, 16'd39924, 16'd58662, 16'd35238, 16'd53969, 16'd35859, 16'd49471, 16'd9220, 16'd51294});
	test_expansion(128'he4a318910aa4ec3ceaa02d010a49d104, {16'd47438, 16'd33081, 16'd22215, 16'd17683, 16'd56001, 16'd24383, 16'd20576, 16'd57819, 16'd22410, 16'd39993, 16'd11703, 16'd35750, 16'd6266, 16'd28193, 16'd34878, 16'd35049, 16'd31155, 16'd127, 16'd53705, 16'd42670, 16'd51344, 16'd39685, 16'd236, 16'd30952, 16'd12780, 16'd48623});
	test_expansion(128'h5245f28936957f1ee6a9c185652f55bc, {16'd8844, 16'd25187, 16'd40873, 16'd56941, 16'd26289, 16'd60030, 16'd42579, 16'd58804, 16'd21963, 16'd59603, 16'd58593, 16'd57459, 16'd20864, 16'd53023, 16'd24608, 16'd29866, 16'd58606, 16'd60987, 16'd28802, 16'd40469, 16'd36956, 16'd28582, 16'd7795, 16'd44196, 16'd49896, 16'd43927});
	test_expansion(128'hdebc2fbf927a827470f8c6533f1f435f, {16'd65140, 16'd43299, 16'd42562, 16'd57308, 16'd33266, 16'd47339, 16'd53530, 16'd44935, 16'd58170, 16'd48382, 16'd20338, 16'd47257, 16'd39766, 16'd62557, 16'd731, 16'd25676, 16'd249, 16'd33829, 16'd9943, 16'd14549, 16'd49359, 16'd6479, 16'd53365, 16'd3506, 16'd25060, 16'd47202});
	test_expansion(128'h1488c1d44a01bf4249db3a260d69cab4, {16'd43594, 16'd62364, 16'd56240, 16'd58949, 16'd62104, 16'd15345, 16'd60830, 16'd7539, 16'd37074, 16'd53343, 16'd62722, 16'd51699, 16'd50221, 16'd33803, 16'd56303, 16'd36173, 16'd54538, 16'd16467, 16'd28884, 16'd53461, 16'd35438, 16'd12606, 16'd872, 16'd9784, 16'd53221, 16'd20015});
	test_expansion(128'hfe3a7149227c0242bcefc892ee3d810c, {16'd39900, 16'd32317, 16'd9565, 16'd63793, 16'd35706, 16'd32668, 16'd16108, 16'd21211, 16'd52967, 16'd46893, 16'd48214, 16'd3309, 16'd28064, 16'd31034, 16'd43569, 16'd62239, 16'd48837, 16'd48751, 16'd15090, 16'd62549, 16'd55903, 16'd54278, 16'd40818, 16'd60344, 16'd1419, 16'd28136});
	test_expansion(128'h73a72d72cf39ac992016dbef69278bcd, {16'd29988, 16'd21483, 16'd8540, 16'd26515, 16'd40047, 16'd43328, 16'd55067, 16'd34213, 16'd14804, 16'd38821, 16'd53614, 16'd52527, 16'd11727, 16'd59509, 16'd62178, 16'd7884, 16'd41035, 16'd40997, 16'd27813, 16'd56725, 16'd30062, 16'd63900, 16'd43211, 16'd56053, 16'd36938, 16'd44433});
	test_expansion(128'hbc5f071d44c1caf7641550e5af4be482, {16'd58448, 16'd46732, 16'd21486, 16'd45828, 16'd5102, 16'd35448, 16'd56997, 16'd50056, 16'd3061, 16'd43908, 16'd16700, 16'd64906, 16'd12419, 16'd55291, 16'd55908, 16'd48082, 16'd13949, 16'd25201, 16'd38979, 16'd930, 16'd11319, 16'd32434, 16'd26317, 16'd23365, 16'd47108, 16'd11175});
	test_expansion(128'h828c729a78221a9ffb67c008f457ae77, {16'd52522, 16'd53405, 16'd58306, 16'd3568, 16'd51284, 16'd58707, 16'd1505, 16'd2863, 16'd60022, 16'd46790, 16'd12862, 16'd51595, 16'd48312, 16'd42945, 16'd54998, 16'd4548, 16'd12705, 16'd39968, 16'd54885, 16'd4354, 16'd6083, 16'd62710, 16'd60245, 16'd32829, 16'd48330, 16'd45171});
	test_expansion(128'h37b243bbb60a2a79044c02390add8bff, {16'd31065, 16'd47539, 16'd61392, 16'd1362, 16'd6717, 16'd5728, 16'd2347, 16'd51602, 16'd54935, 16'd17731, 16'd26621, 16'd39958, 16'd35898, 16'd24266, 16'd10425, 16'd3722, 16'd62908, 16'd4207, 16'd126, 16'd53854, 16'd17301, 16'd54615, 16'd57878, 16'd50536, 16'd13795, 16'd27167});
	test_expansion(128'h56d9cd2847ba2bf53446afba5555cfce, {16'd47351, 16'd11704, 16'd10303, 16'd18165, 16'd50230, 16'd35661, 16'd23977, 16'd17196, 16'd50202, 16'd52821, 16'd49192, 16'd9477, 16'd21960, 16'd64957, 16'd18925, 16'd8120, 16'd31081, 16'd57420, 16'd42380, 16'd32803, 16'd14791, 16'd13576, 16'd35653, 16'd26652, 16'd14008, 16'd40302});
	test_expansion(128'hda7a0d22e73d86726c949c8a5cb98764, {16'd56203, 16'd14549, 16'd29924, 16'd61377, 16'd6625, 16'd9055, 16'd55788, 16'd10408, 16'd38045, 16'd40933, 16'd5607, 16'd23565, 16'd48734, 16'd57512, 16'd56497, 16'd6312, 16'd13585, 16'd19709, 16'd34389, 16'd59546, 16'd57840, 16'd16284, 16'd1995, 16'd55790, 16'd21433, 16'd19139});
	test_expansion(128'hbe00389fdce00a389a0671fb7e4dbd36, {16'd50117, 16'd22049, 16'd5275, 16'd17185, 16'd44627, 16'd10734, 16'd29134, 16'd21311, 16'd14681, 16'd6650, 16'd11968, 16'd13705, 16'd10021, 16'd44535, 16'd57954, 16'd54578, 16'd40851, 16'd54235, 16'd49012, 16'd18884, 16'd34602, 16'd9476, 16'd30254, 16'd41513, 16'd14301, 16'd60693});
	test_expansion(128'hb32a61acdf6ba494f240c1745752c626, {16'd1575, 16'd7363, 16'd30401, 16'd38641, 16'd63794, 16'd55438, 16'd28788, 16'd34429, 16'd51849, 16'd11808, 16'd15889, 16'd35947, 16'd6957, 16'd28074, 16'd27105, 16'd65249, 16'd48723, 16'd1367, 16'd28937, 16'd16658, 16'd12945, 16'd51162, 16'd54123, 16'd9873, 16'd28903, 16'd10110});
	test_expansion(128'h418f1e64bf1b34522003945dd1058acc, {16'd23527, 16'd60578, 16'd534, 16'd62359, 16'd58277, 16'd50550, 16'd23473, 16'd22104, 16'd65227, 16'd7221, 16'd65366, 16'd1669, 16'd28507, 16'd36924, 16'd42936, 16'd7618, 16'd35150, 16'd59587, 16'd1708, 16'd39843, 16'd21404, 16'd60485, 16'd1272, 16'd62295, 16'd40706, 16'd42826});
	test_expansion(128'h6226df64e9d36824bbaa634ac6ba54f4, {16'd5663, 16'd41202, 16'd60061, 16'd5570, 16'd59539, 16'd44768, 16'd23586, 16'd20000, 16'd31115, 16'd39959, 16'd8414, 16'd17362, 16'd60986, 16'd35705, 16'd24033, 16'd19594, 16'd3051, 16'd277, 16'd6652, 16'd32993, 16'd4019, 16'd5633, 16'd62464, 16'd27153, 16'd3804, 16'd26030});
	test_expansion(128'hdeeb462ec8fc7b44e8d3afec11a30c62, {16'd21860, 16'd27897, 16'd53771, 16'd57919, 16'd55922, 16'd17714, 16'd64792, 16'd2511, 16'd52724, 16'd33272, 16'd23785, 16'd33764, 16'd34884, 16'd27052, 16'd48856, 16'd47250, 16'd61976, 16'd58963, 16'd48661, 16'd20509, 16'd13346, 16'd56329, 16'd50508, 16'd15297, 16'd56861, 16'd361});
	test_expansion(128'hb7aff68155a6ad53f1977590354c17a8, {16'd11367, 16'd5194, 16'd45475, 16'd11621, 16'd21814, 16'd30257, 16'd65392, 16'd11423, 16'd57528, 16'd3641, 16'd20237, 16'd25074, 16'd35352, 16'd30090, 16'd43738, 16'd54562, 16'd62170, 16'd48061, 16'd9229, 16'd64239, 16'd47870, 16'd56483, 16'd26118, 16'd56918, 16'd13872, 16'd31768});
	test_expansion(128'hc6e542b7d77bbc246376635aefd60be3, {16'd36239, 16'd871, 16'd10387, 16'd33077, 16'd54313, 16'd60691, 16'd25917, 16'd7189, 16'd19002, 16'd19725, 16'd64416, 16'd23756, 16'd9954, 16'd12921, 16'd44354, 16'd49135, 16'd29478, 16'd39878, 16'd33290, 16'd24607, 16'd28696, 16'd47801, 16'd1862, 16'd19821, 16'd64683, 16'd42810});
	test_expansion(128'hc1c71428ef74ff5e99bd6b1acda79630, {16'd40910, 16'd3633, 16'd40928, 16'd43065, 16'd56416, 16'd59560, 16'd49672, 16'd39604, 16'd44800, 16'd39774, 16'd44168, 16'd32681, 16'd16242, 16'd57863, 16'd11764, 16'd22141, 16'd45886, 16'd7632, 16'd53972, 16'd50236, 16'd1115, 16'd26372, 16'd43413, 16'd7182, 16'd110, 16'd23462});
	test_expansion(128'h2a39d56fbec1bff606f2a8ee9a76e5e4, {16'd21716, 16'd4521, 16'd18466, 16'd44231, 16'd58492, 16'd43837, 16'd25313, 16'd58354, 16'd39502, 16'd62345, 16'd26683, 16'd24957, 16'd24947, 16'd16511, 16'd43748, 16'd56470, 16'd59478, 16'd19516, 16'd48350, 16'd35868, 16'd65108, 16'd54491, 16'd56431, 16'd57746, 16'd59653, 16'd24644});
	test_expansion(128'hed1c3e9212d619317296052ed2f21983, {16'd35685, 16'd57523, 16'd56154, 16'd15261, 16'd10672, 16'd13970, 16'd43634, 16'd30074, 16'd46333, 16'd46975, 16'd39369, 16'd19061, 16'd619, 16'd17237, 16'd7472, 16'd62791, 16'd43854, 16'd34375, 16'd60361, 16'd2596, 16'd1802, 16'd3130, 16'd7318, 16'd43272, 16'd43081, 16'd24021});
	test_expansion(128'h398e21a8a27e67f627a65ee84b3a984a, {16'd51321, 16'd43949, 16'd34183, 16'd10915, 16'd10221, 16'd32169, 16'd26392, 16'd61388, 16'd52691, 16'd24121, 16'd21014, 16'd1738, 16'd64676, 16'd65463, 16'd25844, 16'd51029, 16'd40803, 16'd36971, 16'd24318, 16'd20008, 16'd41512, 16'd35392, 16'd2377, 16'd49722, 16'd18067, 16'd13974});
	test_expansion(128'hde55acf14f46e4ea584ca567736d00c7, {16'd32187, 16'd36482, 16'd43163, 16'd34019, 16'd63024, 16'd54951, 16'd58264, 16'd53772, 16'd50325, 16'd50883, 16'd40534, 16'd40728, 16'd20424, 16'd26022, 16'd61258, 16'd4535, 16'd15499, 16'd47482, 16'd19492, 16'd49760, 16'd22143, 16'd33420, 16'd25539, 16'd18088, 16'd47376, 16'd7649});
	test_expansion(128'h147212a21e3d613e8c9ff1550c49cefd, {16'd50574, 16'd26583, 16'd23580, 16'd13171, 16'd64781, 16'd43273, 16'd24326, 16'd14855, 16'd27551, 16'd34149, 16'd62466, 16'd44568, 16'd61661, 16'd45793, 16'd33337, 16'd46720, 16'd9991, 16'd54376, 16'd55070, 16'd35015, 16'd50172, 16'd32507, 16'd48850, 16'd8975, 16'd4025, 16'd63754});
	test_expansion(128'h17343cbb1cb1aa1450e3ed47fc9c8d9e, {16'd29411, 16'd14909, 16'd24857, 16'd49739, 16'd50156, 16'd11666, 16'd518, 16'd25413, 16'd29291, 16'd28913, 16'd18641, 16'd34008, 16'd26711, 16'd43558, 16'd14218, 16'd48888, 16'd39542, 16'd60687, 16'd54147, 16'd43324, 16'd47865, 16'd56148, 16'd35212, 16'd48931, 16'd47778, 16'd48666});
	test_expansion(128'hee684045f161ad4dc020a54e0a5a34a6, {16'd36973, 16'd26139, 16'd4407, 16'd25083, 16'd33498, 16'd19358, 16'd51792, 16'd52401, 16'd29139, 16'd61568, 16'd29208, 16'd50039, 16'd20853, 16'd33605, 16'd40276, 16'd62612, 16'd9712, 16'd8671, 16'd42176, 16'd35525, 16'd43725, 16'd2103, 16'd29818, 16'd23878, 16'd8512, 16'd61176});
	test_expansion(128'h925b2adc485ab641b5f34e72970bd020, {16'd55758, 16'd36706, 16'd47008, 16'd6954, 16'd31500, 16'd5090, 16'd7460, 16'd26037, 16'd60320, 16'd10288, 16'd44626, 16'd29646, 16'd12089, 16'd21865, 16'd7139, 16'd3091, 16'd29862, 16'd11042, 16'd7148, 16'd49279, 16'd34037, 16'd12825, 16'd23430, 16'd13568, 16'd59079, 16'd48560});
	test_expansion(128'h67e34b8fc0f7e14a644775dc8e77a04d, {16'd1616, 16'd10818, 16'd20255, 16'd5858, 16'd61246, 16'd20747, 16'd8174, 16'd52198, 16'd4584, 16'd13465, 16'd31633, 16'd35421, 16'd33857, 16'd60700, 16'd50128, 16'd28735, 16'd60971, 16'd3396, 16'd59754, 16'd1780, 16'd3999, 16'd7941, 16'd8801, 16'd37987, 16'd6428, 16'd63172});
	test_expansion(128'h90afa58999b1896a3b2dd7bde63e1d0d, {16'd62397, 16'd43152, 16'd46151, 16'd25978, 16'd19684, 16'd13034, 16'd9116, 16'd14266, 16'd8173, 16'd60348, 16'd45676, 16'd64339, 16'd64954, 16'd6996, 16'd47844, 16'd18618, 16'd63453, 16'd38132, 16'd49858, 16'd28602, 16'd56641, 16'd62955, 16'd7843, 16'd49650, 16'd56231, 16'd29517});
	test_expansion(128'h1166825c83b21bf4f52376663981808c, {16'd49989, 16'd38698, 16'd3812, 16'd56090, 16'd24123, 16'd18125, 16'd57474, 16'd18096, 16'd11300, 16'd42348, 16'd52779, 16'd42042, 16'd17784, 16'd29278, 16'd45164, 16'd41571, 16'd383, 16'd7072, 16'd4325, 16'd59512, 16'd5204, 16'd63545, 16'd4778, 16'd25719, 16'd2334, 16'd63367});
	test_expansion(128'h0f63de67c4f98c05a849c7fa82a2814c, {16'd58622, 16'd19815, 16'd47512, 16'd6240, 16'd45023, 16'd27258, 16'd54790, 16'd60882, 16'd21146, 16'd57312, 16'd18936, 16'd24795, 16'd19312, 16'd34117, 16'd64573, 16'd9175, 16'd42339, 16'd18817, 16'd4570, 16'd51571, 16'd14525, 16'd1565, 16'd14273, 16'd54787, 16'd505, 16'd28192});
	test_expansion(128'haa296472ca8261cc0567b0997ae3755f, {16'd7764, 16'd30382, 16'd55391, 16'd51321, 16'd15086, 16'd14301, 16'd2694, 16'd6001, 16'd53999, 16'd33350, 16'd23680, 16'd120, 16'd9394, 16'd52688, 16'd15167, 16'd52924, 16'd45478, 16'd64863, 16'd39894, 16'd64525, 16'd4295, 16'd3340, 16'd86, 16'd16065, 16'd37873, 16'd23185});
	test_expansion(128'h01bc305a61a98a643e123c62d83b1e71, {16'd57293, 16'd63254, 16'd44335, 16'd31708, 16'd55814, 16'd5348, 16'd63646, 16'd45085, 16'd20977, 16'd4290, 16'd57277, 16'd52520, 16'd63662, 16'd51247, 16'd32542, 16'd37220, 16'd49075, 16'd48479, 16'd39674, 16'd58239, 16'd57483, 16'd58576, 16'd33384, 16'd8485, 16'd29936, 16'd27890});
	test_expansion(128'hd057d20b8fbf7e9472ff412b38269310, {16'd29704, 16'd63733, 16'd45490, 16'd26577, 16'd12976, 16'd53936, 16'd51160, 16'd25081, 16'd34190, 16'd39752, 16'd8914, 16'd4723, 16'd48232, 16'd19258, 16'd10575, 16'd10148, 16'd43219, 16'd59365, 16'd35393, 16'd36310, 16'd26, 16'd26290, 16'd40383, 16'd28251, 16'd38776, 16'd34262});
	test_expansion(128'hfe0462720ba1ac8cf370170427b177ff, {16'd65190, 16'd13224, 16'd53660, 16'd22742, 16'd38709, 16'd49557, 16'd36012, 16'd52195, 16'd2899, 16'd762, 16'd18314, 16'd39862, 16'd39402, 16'd25970, 16'd59038, 16'd34359, 16'd16588, 16'd50019, 16'd36278, 16'd16124, 16'd59354, 16'd12067, 16'd56467, 16'd25817, 16'd16246, 16'd3635});
	test_expansion(128'hd2e75b66f48b900f80b590243c1b31a3, {16'd3481, 16'd22237, 16'd39028, 16'd3289, 16'd10518, 16'd18703, 16'd41542, 16'd15885, 16'd13141, 16'd25379, 16'd3679, 16'd37709, 16'd35888, 16'd52807, 16'd41352, 16'd17495, 16'd40306, 16'd31208, 16'd55817, 16'd51393, 16'd57275, 16'd33633, 16'd10722, 16'd61351, 16'd47405, 16'd23704});
	test_expansion(128'h06a97f0e62b9cce67e4e4c556cf78dd3, {16'd40064, 16'd32993, 16'd45709, 16'd47636, 16'd34772, 16'd60956, 16'd23554, 16'd31710, 16'd57665, 16'd16252, 16'd28748, 16'd41480, 16'd28639, 16'd45746, 16'd45004, 16'd47466, 16'd25861, 16'd60011, 16'd11620, 16'd40014, 16'd1791, 16'd49947, 16'd15904, 16'd9056, 16'd50520, 16'd42166});
	test_expansion(128'hde39a8f14357ffcf11d9fa1d804d175b, {16'd21714, 16'd37229, 16'd59223, 16'd7153, 16'd45411, 16'd64491, 16'd58597, 16'd37581, 16'd37688, 16'd14867, 16'd12829, 16'd2688, 16'd64745, 16'd59564, 16'd56811, 16'd62706, 16'd61946, 16'd26484, 16'd33155, 16'd5511, 16'd11346, 16'd62512, 16'd36983, 16'd34503, 16'd39944, 16'd22013});
	test_expansion(128'h46cf7f1bf38d00a80d60829d95db99ec, {16'd12485, 16'd56432, 16'd13052, 16'd23168, 16'd10105, 16'd63012, 16'd29591, 16'd46203, 16'd14208, 16'd18511, 16'd35718, 16'd22678, 16'd7108, 16'd27473, 16'd45449, 16'd21313, 16'd13719, 16'd14118, 16'd37867, 16'd55615, 16'd1397, 16'd32719, 16'd47139, 16'd64848, 16'd63505, 16'd59754});
	test_expansion(128'hd2ed46c454bdcfb5642f1b2a4f81a353, {16'd24289, 16'd37861, 16'd51014, 16'd14964, 16'd58875, 16'd8356, 16'd41851, 16'd54062, 16'd11063, 16'd27794, 16'd48284, 16'd47219, 16'd33580, 16'd6484, 16'd20149, 16'd3984, 16'd65058, 16'd62946, 16'd39570, 16'd39475, 16'd50033, 16'd59843, 16'd1980, 16'd40109, 16'd56762, 16'd18018});
	test_expansion(128'h9c2ef46dde1670f12cd9cbab095b1660, {16'd61809, 16'd8073, 16'd57128, 16'd18281, 16'd38010, 16'd64144, 16'd47141, 16'd21118, 16'd5363, 16'd29122, 16'd51658, 16'd53531, 16'd24860, 16'd40020, 16'd2954, 16'd18383, 16'd30708, 16'd7806, 16'd65222, 16'd36463, 16'd59918, 16'd7937, 16'd42490, 16'd3077, 16'd27257, 16'd9890});
	test_expansion(128'he51357fb1f762cffd07d10ce0f70c416, {16'd20484, 16'd528, 16'd56883, 16'd46821, 16'd27624, 16'd2992, 16'd13230, 16'd62938, 16'd50325, 16'd60636, 16'd64915, 16'd2648, 16'd58544, 16'd55396, 16'd37667, 16'd44283, 16'd59300, 16'd16542, 16'd18828, 16'd35728, 16'd46799, 16'd13274, 16'd32724, 16'd62319, 16'd26743, 16'd56335});
	test_expansion(128'h45c612654dd8a20efcdb8c204b2b571f, {16'd42406, 16'd59120, 16'd10789, 16'd57039, 16'd53345, 16'd13958, 16'd50058, 16'd19765, 16'd24537, 16'd44113, 16'd28014, 16'd30395, 16'd52907, 16'd57720, 16'd4646, 16'd39991, 16'd46119, 16'd9854, 16'd56535, 16'd65273, 16'd40782, 16'd34079, 16'd5206, 16'd47097, 16'd3652, 16'd53521});
	test_expansion(128'hf37b103c002ade53fdfe2a5e973ffadb, {16'd45593, 16'd64382, 16'd12153, 16'd37137, 16'd37852, 16'd9425, 16'd15147, 16'd31346, 16'd44091, 16'd31803, 16'd5933, 16'd58659, 16'd32567, 16'd19967, 16'd5595, 16'd15727, 16'd34562, 16'd5419, 16'd31865, 16'd25172, 16'd14395, 16'd6185, 16'd60976, 16'd13689, 16'd9617, 16'd59447});
	test_expansion(128'hb7a10fac3dba69221eb4d09854630a74, {16'd3145, 16'd36411, 16'd17207, 16'd3292, 16'd8655, 16'd7021, 16'd49718, 16'd22822, 16'd18466, 16'd36346, 16'd34112, 16'd7986, 16'd56388, 16'd29457, 16'd62646, 16'd61590, 16'd61629, 16'd16834, 16'd1443, 16'd24149, 16'd51297, 16'd32270, 16'd17093, 16'd16153, 16'd24161, 16'd52428});
	test_expansion(128'h98191692f8c109d5e9d628d4bbe9f01d, {16'd26711, 16'd38199, 16'd21620, 16'd5830, 16'd48153, 16'd27130, 16'd58303, 16'd28827, 16'd553, 16'd56172, 16'd36051, 16'd3040, 16'd62613, 16'd45723, 16'd20921, 16'd65191, 16'd41074, 16'd5278, 16'd13670, 16'd54950, 16'd6728, 16'd4445, 16'd61630, 16'd10239, 16'd36345, 16'd47771});
	test_expansion(128'h4e406dd5f1518a64473549d813dd7afb, {16'd27365, 16'd43963, 16'd52308, 16'd14421, 16'd65448, 16'd63558, 16'd20716, 16'd44787, 16'd26166, 16'd58493, 16'd9357, 16'd36058, 16'd23058, 16'd37908, 16'd24119, 16'd31795, 16'd12731, 16'd64549, 16'd56, 16'd63357, 16'd65517, 16'd30605, 16'd17933, 16'd29164, 16'd23718, 16'd2803});
	test_expansion(128'had30f58d9090f99d56a3532093783404, {16'd28361, 16'd20401, 16'd21132, 16'd20470, 16'd15613, 16'd34473, 16'd59030, 16'd14400, 16'd52642, 16'd25900, 16'd16948, 16'd5461, 16'd13172, 16'd33679, 16'd49912, 16'd30957, 16'd13637, 16'd4277, 16'd796, 16'd63053, 16'd5639, 16'd53445, 16'd26037, 16'd9297, 16'd45518, 16'd29185});
	test_expansion(128'h0448c0ade2a99fed4f84521a049f85e2, {16'd39728, 16'd17444, 16'd1789, 16'd12584, 16'd415, 16'd1247, 16'd53088, 16'd40003, 16'd30151, 16'd48551, 16'd25903, 16'd12248, 16'd63953, 16'd29566, 16'd25368, 16'd58002, 16'd65221, 16'd43740, 16'd41448, 16'd62190, 16'd22569, 16'd18464, 16'd26802, 16'd46807, 16'd3392, 16'd62416});
	test_expansion(128'h397cb2afe43cf6191858a53d5cd6deb3, {16'd7612, 16'd41382, 16'd7766, 16'd53476, 16'd61498, 16'd8085, 16'd39064, 16'd64572, 16'd61253, 16'd27952, 16'd51640, 16'd13007, 16'd25702, 16'd62618, 16'd197, 16'd36039, 16'd62044, 16'd56294, 16'd7975, 16'd28260, 16'd36987, 16'd9555, 16'd29160, 16'd18313, 16'd63266, 16'd59732});
	test_expansion(128'hd904a5d8c052526a35230af482d2ab6f, {16'd53251, 16'd33404, 16'd16091, 16'd20977, 16'd20747, 16'd10432, 16'd37623, 16'd27336, 16'd30861, 16'd31133, 16'd28820, 16'd44233, 16'd25097, 16'd49736, 16'd50650, 16'd57373, 16'd36740, 16'd40094, 16'd16232, 16'd4170, 16'd58423, 16'd29337, 16'd14876, 16'd42521, 16'd12273, 16'd63388});
	test_expansion(128'h7b1c256022de29363b6e24f2a1cc7d5f, {16'd44274, 16'd30381, 16'd13639, 16'd43620, 16'd49812, 16'd2249, 16'd32384, 16'd21981, 16'd37122, 16'd62720, 16'd20932, 16'd5294, 16'd45040, 16'd29571, 16'd23663, 16'd65016, 16'd52595, 16'd30305, 16'd61155, 16'd30501, 16'd14289, 16'd46975, 16'd62802, 16'd49579, 16'd44839, 16'd52878});
	test_expansion(128'hcdc5942e5ea64586c4329b18794f5e46, {16'd12385, 16'd52979, 16'd8506, 16'd55653, 16'd17553, 16'd37875, 16'd18465, 16'd64401, 16'd61425, 16'd50609, 16'd29605, 16'd59451, 16'd45843, 16'd59822, 16'd8392, 16'd57320, 16'd56974, 16'd29082, 16'd25918, 16'd9670, 16'd10567, 16'd12643, 16'd55979, 16'd14530, 16'd52437, 16'd50603});
	test_expansion(128'h69cd80471b3cff8df0654bb14c545565, {16'd8874, 16'd54299, 16'd44244, 16'd16820, 16'd21952, 16'd2834, 16'd14037, 16'd53417, 16'd14477, 16'd33199, 16'd12534, 16'd59178, 16'd3511, 16'd37281, 16'd9514, 16'd31112, 16'd10892, 16'd130, 16'd12836, 16'd40834, 16'd30324, 16'd15649, 16'd21079, 16'd7078, 16'd36612, 16'd30320});
	test_expansion(128'he6cce520789a7d36df4db9fe33b75472, {16'd21716, 16'd10504, 16'd46784, 16'd37471, 16'd64769, 16'd23952, 16'd36394, 16'd3967, 16'd13066, 16'd25652, 16'd15701, 16'd59922, 16'd39649, 16'd40397, 16'd55965, 16'd7520, 16'd21417, 16'd42064, 16'd32351, 16'd36784, 16'd64904, 16'd55429, 16'd1323, 16'd49591, 16'd49735, 16'd55169});
	test_expansion(128'h1daefc644a0619e4d5c4bfe688886c4d, {16'd53070, 16'd18614, 16'd49631, 16'd2204, 16'd26331, 16'd30364, 16'd213, 16'd39078, 16'd32284, 16'd50843, 16'd26435, 16'd17425, 16'd42414, 16'd44723, 16'd64976, 16'd44499, 16'd40070, 16'd46104, 16'd15445, 16'd37912, 16'd40411, 16'd63849, 16'd17923, 16'd27165, 16'd53624, 16'd59275});
	test_expansion(128'hd05fb10a45d271ce7c55aaf70d534529, {16'd25082, 16'd32940, 16'd7668, 16'd49002, 16'd9153, 16'd33684, 16'd62080, 16'd63907, 16'd22806, 16'd52759, 16'd6320, 16'd8181, 16'd19467, 16'd64315, 16'd24719, 16'd11974, 16'd57667, 16'd21999, 16'd44734, 16'd36502, 16'd62932, 16'd15372, 16'd23025, 16'd30025, 16'd615, 16'd40854});
	test_expansion(128'h064e65e7e92511cdc171549926dd0339, {16'd52150, 16'd44966, 16'd56087, 16'd20188, 16'd26467, 16'd3076, 16'd65498, 16'd55109, 16'd25496, 16'd52983, 16'd42433, 16'd41613, 16'd64861, 16'd52979, 16'd12390, 16'd47877, 16'd18761, 16'd8347, 16'd54336, 16'd56315, 16'd57033, 16'd2054, 16'd61174, 16'd64322, 16'd61446, 16'd5551});
	test_expansion(128'h79f44f8e3a2e53dbe0dcc7c3dc493323, {16'd26322, 16'd33154, 16'd42980, 16'd8779, 16'd18794, 16'd64556, 16'd24454, 16'd4506, 16'd19744, 16'd26066, 16'd23191, 16'd13017, 16'd16812, 16'd59682, 16'd25904, 16'd16026, 16'd61599, 16'd26842, 16'd53255, 16'd45794, 16'd13726, 16'd24190, 16'd26229, 16'd48952, 16'd2687, 16'd7212});
	test_expansion(128'h4f2e31402ff7204bcef5c382e2df93db, {16'd60644, 16'd20410, 16'd6743, 16'd36997, 16'd14885, 16'd37206, 16'd42173, 16'd56181, 16'd33879, 16'd26142, 16'd43917, 16'd28990, 16'd7515, 16'd31828, 16'd60919, 16'd18905, 16'd58244, 16'd11720, 16'd9653, 16'd56000, 16'd57138, 16'd43300, 16'd36756, 16'd10700, 16'd46770, 16'd65268});
	test_expansion(128'h5777d897ca82d1bf5f1dba7c09780a2c, {16'd4327, 16'd48374, 16'd60684, 16'd62112, 16'd37079, 16'd55140, 16'd10094, 16'd58136, 16'd23300, 16'd1, 16'd55282, 16'd19570, 16'd23270, 16'd12233, 16'd33777, 16'd55477, 16'd55227, 16'd21844, 16'd51648, 16'd18814, 16'd43936, 16'd26850, 16'd47517, 16'd45943, 16'd46006, 16'd55138});
	test_expansion(128'hb1a5b41bbd4985d890ea7c7d57870bf5, {16'd19300, 16'd21189, 16'd37336, 16'd31263, 16'd58534, 16'd61018, 16'd1263, 16'd41842, 16'd37263, 16'd51470, 16'd23601, 16'd7603, 16'd57356, 16'd22587, 16'd20637, 16'd1239, 16'd57187, 16'd32414, 16'd13222, 16'd25576, 16'd63436, 16'd45344, 16'd12599, 16'd52315, 16'd20148, 16'd27119});
	test_expansion(128'h0b277c86d0708b39f41f67363af1e3b0, {16'd24290, 16'd56884, 16'd44404, 16'd58545, 16'd21783, 16'd31198, 16'd38284, 16'd42018, 16'd29748, 16'd25934, 16'd26517, 16'd57684, 16'd64165, 16'd18702, 16'd1218, 16'd3839, 16'd64325, 16'd11141, 16'd13931, 16'd36057, 16'd56636, 16'd15966, 16'd50185, 16'd62799, 16'd57979, 16'd42990});
	test_expansion(128'h49cff067c066a9dcb99b5c0dc062da7d, {16'd42495, 16'd26335, 16'd49775, 16'd37286, 16'd54416, 16'd18651, 16'd16358, 16'd64033, 16'd59226, 16'd3442, 16'd51418, 16'd43059, 16'd36869, 16'd44377, 16'd38762, 16'd31941, 16'd13304, 16'd7295, 16'd15566, 16'd61746, 16'd50027, 16'd54831, 16'd5105, 16'd17496, 16'd44200, 16'd8420});
	test_expansion(128'h3b24b3e6cdd7988b87b7a5f3df0c3db0, {16'd44916, 16'd9534, 16'd44697, 16'd20516, 16'd5034, 16'd63149, 16'd19897, 16'd5653, 16'd23035, 16'd10294, 16'd40372, 16'd50123, 16'd1575, 16'd58702, 16'd28737, 16'd31883, 16'd40646, 16'd60058, 16'd8724, 16'd50612, 16'd51192, 16'd24037, 16'd8117, 16'd18872, 16'd9534, 16'd48907});
	test_expansion(128'h70a1bc978def4a9d23b6b954eafb6a1e, {16'd63337, 16'd24823, 16'd57196, 16'd4857, 16'd60544, 16'd17023, 16'd19950, 16'd46637, 16'd55201, 16'd42916, 16'd8076, 16'd22889, 16'd27310, 16'd56276, 16'd49517, 16'd34414, 16'd29460, 16'd2908, 16'd33355, 16'd33676, 16'd41722, 16'd52842, 16'd4804, 16'd17631, 16'd9709, 16'd21705});
	test_expansion(128'hb45a73a4fb0d1b755305e58a19fe1272, {16'd43667, 16'd17035, 16'd24795, 16'd40516, 16'd25382, 16'd3055, 16'd53118, 16'd43236, 16'd38456, 16'd36769, 16'd56636, 16'd35412, 16'd12613, 16'd26577, 16'd3485, 16'd3105, 16'd28167, 16'd18995, 16'd41439, 16'd1073, 16'd743, 16'd7884, 16'd33352, 16'd10531, 16'd41112, 16'd58319});
	test_expansion(128'h240c5de17deef70fccef1456075656fe, {16'd40885, 16'd29386, 16'd4975, 16'd39612, 16'd7638, 16'd24366, 16'd12803, 16'd54649, 16'd48387, 16'd61231, 16'd64203, 16'd60849, 16'd58201, 16'd24551, 16'd10459, 16'd47492, 16'd54941, 16'd19435, 16'd38153, 16'd10320, 16'd29238, 16'd41139, 16'd27055, 16'd23195, 16'd28643, 16'd57231});
	test_expansion(128'h99254d3548d5423a1feb5e39cb461048, {16'd51067, 16'd25213, 16'd14511, 16'd38324, 16'd30198, 16'd23642, 16'd14377, 16'd30909, 16'd45908, 16'd15588, 16'd28670, 16'd62295, 16'd16734, 16'd34644, 16'd34382, 16'd15063, 16'd5095, 16'd13645, 16'd43731, 16'd29462, 16'd56773, 16'd37004, 16'd49447, 16'd63282, 16'd12388, 16'd17970});
	test_expansion(128'h6f5a1fdca68d630cf4edc7297acc8792, {16'd4492, 16'd43809, 16'd44124, 16'd22378, 16'd28025, 16'd41973, 16'd21734, 16'd23428, 16'd9385, 16'd43544, 16'd19530, 16'd53499, 16'd23293, 16'd39568, 16'd58669, 16'd46292, 16'd6579, 16'd1103, 16'd394, 16'd33609, 16'd20652, 16'd12861, 16'd58708, 16'd48065, 16'd26812, 16'd30640});
	test_expansion(128'h2ddc8c15d89dcc6b7cf085b3c552a0dc, {16'd26881, 16'd48460, 16'd47150, 16'd41523, 16'd45674, 16'd54427, 16'd823, 16'd65070, 16'd8800, 16'd41130, 16'd44851, 16'd62757, 16'd2609, 16'd18172, 16'd62137, 16'd40234, 16'd64384, 16'd24735, 16'd50128, 16'd7848, 16'd58393, 16'd33956, 16'd28819, 16'd33482, 16'd6103, 16'd9758});
	test_expansion(128'h772359d68217106df210da1414079187, {16'd300, 16'd52969, 16'd36325, 16'd41824, 16'd33537, 16'd2382, 16'd49888, 16'd40673, 16'd54217, 16'd58201, 16'd42775, 16'd35018, 16'd64963, 16'd34921, 16'd47265, 16'd38765, 16'd20323, 16'd29176, 16'd47359, 16'd45008, 16'd23672, 16'd48748, 16'd40468, 16'd33829, 16'd23839, 16'd9000});
	test_expansion(128'h25560b139adc8397a93d23f4da1b9633, {16'd3268, 16'd3938, 16'd15211, 16'd7866, 16'd49246, 16'd53704, 16'd7548, 16'd2482, 16'd44345, 16'd22316, 16'd46560, 16'd51710, 16'd48846, 16'd43256, 16'd27537, 16'd26037, 16'd37445, 16'd21630, 16'd22851, 16'd59672, 16'd5000, 16'd32560, 16'd54409, 16'd20427, 16'd10391, 16'd28771});
	test_expansion(128'hda2f90189b99b1113c2dde1148b8b34f, {16'd29953, 16'd61094, 16'd9596, 16'd3397, 16'd45967, 16'd27650, 16'd10550, 16'd18509, 16'd43020, 16'd33995, 16'd20417, 16'd29925, 16'd10610, 16'd63561, 16'd20066, 16'd12442, 16'd39447, 16'd27891, 16'd2961, 16'd56272, 16'd22135, 16'd47417, 16'd57509, 16'd1766, 16'd43013, 16'd24367});
	test_expansion(128'h39de4fe0afbb146b0c61cb74c1606df5, {16'd62682, 16'd39076, 16'd12111, 16'd51073, 16'd55505, 16'd60654, 16'd7832, 16'd57928, 16'd48306, 16'd17613, 16'd6188, 16'd56807, 16'd63697, 16'd56837, 16'd26900, 16'd64477, 16'd22663, 16'd2941, 16'd18064, 16'd44487, 16'd34031, 16'd37699, 16'd55986, 16'd17660, 16'd45010, 16'd9669});
	test_expansion(128'h372bf439daf585ae37d7206d85d56199, {16'd50113, 16'd7327, 16'd22928, 16'd35046, 16'd44616, 16'd11215, 16'd51279, 16'd18750, 16'd62597, 16'd53815, 16'd13346, 16'd37043, 16'd60245, 16'd50657, 16'd30423, 16'd9072, 16'd63116, 16'd54475, 16'd57510, 16'd64325, 16'd59365, 16'd42207, 16'd4797, 16'd62697, 16'd44875, 16'd29673});
	test_expansion(128'h6ec4420f7d1d49d3fee9425f9692b8bc, {16'd29836, 16'd45858, 16'd15032, 16'd8460, 16'd11712, 16'd37580, 16'd32929, 16'd44416, 16'd38374, 16'd4006, 16'd14892, 16'd5281, 16'd12197, 16'd1976, 16'd39039, 16'd22117, 16'd16929, 16'd22587, 16'd38413, 16'd42433, 16'd19599, 16'd36059, 16'd22603, 16'd41163, 16'd54216, 16'd45216});
	test_expansion(128'h8b3ed56d566149b7175ede7906947731, {16'd23306, 16'd54096, 16'd24720, 16'd5362, 16'd513, 16'd39826, 16'd20878, 16'd34274, 16'd1864, 16'd59648, 16'd9445, 16'd24645, 16'd7208, 16'd47287, 16'd28353, 16'd62131, 16'd13645, 16'd24732, 16'd37834, 16'd45816, 16'd20443, 16'd59820, 16'd29106, 16'd54282, 16'd4678, 16'd24708});
	test_expansion(128'h208c845ca8c53eea95437dda4907af89, {16'd51268, 16'd9053, 16'd58651, 16'd38837, 16'd64099, 16'd44397, 16'd38376, 16'd28352, 16'd29362, 16'd52896, 16'd59829, 16'd23467, 16'd56154, 16'd44218, 16'd35560, 16'd7434, 16'd57930, 16'd32309, 16'd35614, 16'd53366, 16'd46425, 16'd61372, 16'd52621, 16'd32942, 16'd61149, 16'd678});
	test_expansion(128'he9020a298f6fbcf00986ac4d9d585075, {16'd33645, 16'd10908, 16'd47687, 16'd27411, 16'd31734, 16'd60271, 16'd56077, 16'd5521, 16'd3540, 16'd46497, 16'd56890, 16'd21476, 16'd10953, 16'd24756, 16'd26440, 16'd6128, 16'd2164, 16'd62452, 16'd56740, 16'd36975, 16'd63067, 16'd7414, 16'd32050, 16'd29206, 16'd26382, 16'd58926});
	test_expansion(128'h36ffa13e41c09375946dd23593a58a10, {16'd33547, 16'd24969, 16'd15250, 16'd7348, 16'd54817, 16'd50485, 16'd56480, 16'd25193, 16'd6859, 16'd32754, 16'd9498, 16'd16361, 16'd40546, 16'd13906, 16'd46056, 16'd28888, 16'd19191, 16'd8730, 16'd55852, 16'd27375, 16'd43881, 16'd6568, 16'd9903, 16'd53454, 16'd18144, 16'd461});
	test_expansion(128'hab5cd24911d85d8d9c8ff66b9a963c15, {16'd53248, 16'd41584, 16'd24577, 16'd30039, 16'd31432, 16'd11628, 16'd5011, 16'd39988, 16'd12719, 16'd42156, 16'd7571, 16'd1896, 16'd29847, 16'd12403, 16'd46194, 16'd46258, 16'd51641, 16'd59313, 16'd26353, 16'd570, 16'd1316, 16'd53632, 16'd40435, 16'd10851, 16'd21698, 16'd5024});
	test_expansion(128'h87d5778ff248f813bf6a299e1e1361c7, {16'd45368, 16'd20321, 16'd44561, 16'd16716, 16'd50226, 16'd24703, 16'd61947, 16'd59616, 16'd43304, 16'd41492, 16'd20259, 16'd662, 16'd51751, 16'd45325, 16'd15497, 16'd27484, 16'd62408, 16'd63453, 16'd37361, 16'd51198, 16'd46806, 16'd28656, 16'd3830, 16'd1139, 16'd25110, 16'd36434});
	test_expansion(128'heeba678bbdb3d56102b0729e5a9d10ad, {16'd9844, 16'd32628, 16'd14895, 16'd53424, 16'd64158, 16'd15052, 16'd51928, 16'd3730, 16'd1169, 16'd28027, 16'd10712, 16'd42578, 16'd28700, 16'd22035, 16'd14440, 16'd31466, 16'd947, 16'd40179, 16'd41128, 16'd51123, 16'd40497, 16'd27252, 16'd61038, 16'd39635, 16'd16502, 16'd19415});
	test_expansion(128'h4537588ab7fda8079675ceae1b6ab01f, {16'd27772, 16'd43522, 16'd6905, 16'd50291, 16'd34519, 16'd380, 16'd37216, 16'd61230, 16'd49470, 16'd27023, 16'd15912, 16'd20823, 16'd56086, 16'd53145, 16'd17133, 16'd56195, 16'd62202, 16'd1738, 16'd818, 16'd37867, 16'd21140, 16'd27347, 16'd61129, 16'd15458, 16'd18908, 16'd38995});
	test_expansion(128'h23a1cf33e993481964ee3a6487519d88, {16'd26943, 16'd32516, 16'd6824, 16'd39860, 16'd50145, 16'd7137, 16'd25004, 16'd18311, 16'd7701, 16'd13163, 16'd14115, 16'd54237, 16'd38601, 16'd60567, 16'd18628, 16'd3410, 16'd28744, 16'd45616, 16'd54637, 16'd42313, 16'd33199, 16'd57475, 16'd57428, 16'd3987, 16'd22831, 16'd3118});
	test_expansion(128'h6e81445ae73551e81aba8af793a27233, {16'd15109, 16'd61872, 16'd17226, 16'd197, 16'd898, 16'd31073, 16'd5562, 16'd2498, 16'd18965, 16'd15047, 16'd31164, 16'd22914, 16'd27321, 16'd30899, 16'd54432, 16'd24511, 16'd25189, 16'd23332, 16'd1805, 16'd34441, 16'd50196, 16'd2432, 16'd42748, 16'd420, 16'd44323, 16'd24227});
	test_expansion(128'h0f48fe9b5a476a900fec2c9a4b8e9cba, {16'd22649, 16'd55417, 16'd39205, 16'd40243, 16'd61936, 16'd27123, 16'd16746, 16'd20204, 16'd5591, 16'd64369, 16'd38589, 16'd34247, 16'd47284, 16'd1952, 16'd47291, 16'd49165, 16'd25618, 16'd11932, 16'd29966, 16'd64465, 16'd31533, 16'd48695, 16'd47533, 16'd53281, 16'd64567, 16'd43553});
	test_expansion(128'h436eac96b07f6bbefca7f4ca5cf25917, {16'd32333, 16'd30130, 16'd64707, 16'd35792, 16'd40273, 16'd42738, 16'd13499, 16'd22746, 16'd46165, 16'd13356, 16'd31476, 16'd15461, 16'd31302, 16'd21768, 16'd2363, 16'd39763, 16'd43775, 16'd30158, 16'd26159, 16'd13454, 16'd12795, 16'd34803, 16'd49727, 16'd60842, 16'd47767, 16'd36172});
	test_expansion(128'h69cc2b8ad720d3b9becb5734bd234b17, {16'd49229, 16'd64326, 16'd9103, 16'd27678, 16'd2927, 16'd50698, 16'd16993, 16'd2826, 16'd34458, 16'd26886, 16'd40105, 16'd27777, 16'd40889, 16'd23550, 16'd1655, 16'd42763, 16'd2906, 16'd37053, 16'd46762, 16'd13503, 16'd15145, 16'd9257, 16'd32459, 16'd40189, 16'd26897, 16'd17605});
	test_expansion(128'h1257688141bd244c0882f17c50cc54cd, {16'd10505, 16'd35766, 16'd8957, 16'd12464, 16'd59243, 16'd36608, 16'd7721, 16'd22820, 16'd4518, 16'd64578, 16'd56762, 16'd30912, 16'd24760, 16'd23095, 16'd34448, 16'd24385, 16'd65223, 16'd16271, 16'd62860, 16'd12317, 16'd9961, 16'd60691, 16'd16061, 16'd17269, 16'd26839, 16'd40795});
	test_expansion(128'h0cb4f70800763238005c7d3d2710f1bb, {16'd23189, 16'd9829, 16'd38310, 16'd62590, 16'd23142, 16'd22999, 16'd48256, 16'd50869, 16'd2935, 16'd40556, 16'd52821, 16'd60358, 16'd43246, 16'd62583, 16'd59829, 16'd15046, 16'd17511, 16'd55770, 16'd23444, 16'd55146, 16'd21880, 16'd39432, 16'd59035, 16'd58215, 16'd51468, 16'd9984});
	test_expansion(128'h26a5c35fe39068b1717e940965d820f6, {16'd54642, 16'd58668, 16'd29741, 16'd46561, 16'd33058, 16'd61350, 16'd27519, 16'd24478, 16'd50870, 16'd48921, 16'd48693, 16'd59593, 16'd11884, 16'd43578, 16'd31120, 16'd31572, 16'd42346, 16'd55434, 16'd10973, 16'd34079, 16'd39677, 16'd37347, 16'd61591, 16'd5477, 16'd18520, 16'd21275});
	test_expansion(128'hdb41fed6e2a2740e2674e46282b54006, {16'd52810, 16'd18144, 16'd9185, 16'd54112, 16'd6743, 16'd25194, 16'd29224, 16'd27314, 16'd5092, 16'd62610, 16'd33140, 16'd43982, 16'd63605, 16'd2219, 16'd16566, 16'd49190, 16'd51877, 16'd520, 16'd29382, 16'd37171, 16'd43191, 16'd52289, 16'd3343, 16'd16150, 16'd24472, 16'd6461});
	test_expansion(128'head0e9a7c56160b09692b4d42763251c, {16'd52226, 16'd28935, 16'd55451, 16'd16674, 16'd33616, 16'd33831, 16'd18597, 16'd39367, 16'd34005, 16'd19503, 16'd42176, 16'd65521, 16'd34998, 16'd29222, 16'd42578, 16'd2074, 16'd29451, 16'd4504, 16'd38020, 16'd38224, 16'd5451, 16'd61098, 16'd23410, 16'd51350, 16'd27740, 16'd21353});
	test_expansion(128'h41a04929c333dfa75cc4ed62205325c6, {16'd28543, 16'd20538, 16'd5114, 16'd7299, 16'd7217, 16'd35695, 16'd20079, 16'd65074, 16'd48605, 16'd38021, 16'd48855, 16'd19116, 16'd20695, 16'd35001, 16'd9337, 16'd19799, 16'd36426, 16'd5889, 16'd43700, 16'd44389, 16'd29481, 16'd7499, 16'd31422, 16'd32860, 16'd17277, 16'd10282});
	test_expansion(128'hedfba61f0f787e12d610209b52ce8ae2, {16'd42295, 16'd23983, 16'd63814, 16'd60962, 16'd7970, 16'd27529, 16'd50392, 16'd13729, 16'd10865, 16'd44668, 16'd50548, 16'd54781, 16'd7646, 16'd990, 16'd57093, 16'd14059, 16'd40082, 16'd49842, 16'd61990, 16'd47219, 16'd57483, 16'd41620, 16'd10395, 16'd24067, 16'd39113, 16'd45443});
	test_expansion(128'h40817c27487e2b659bcff106868cfb73, {16'd19160, 16'd62982, 16'd24214, 16'd51993, 16'd9798, 16'd10838, 16'd44888, 16'd31045, 16'd12168, 16'd45990, 16'd60289, 16'd30860, 16'd19353, 16'd52799, 16'd32136, 16'd33579, 16'd16504, 16'd31839, 16'd56229, 16'd13067, 16'd19380, 16'd31202, 16'd29868, 16'd19155, 16'd21748, 16'd50901});
	test_expansion(128'hba3fcd49126f31811a3b1ecbf39a9653, {16'd65363, 16'd58104, 16'd59834, 16'd25393, 16'd4512, 16'd44327, 16'd58762, 16'd39165, 16'd43715, 16'd57953, 16'd15828, 16'd6991, 16'd61729, 16'd39986, 16'd62019, 16'd32450, 16'd3917, 16'd48999, 16'd60578, 16'd48229, 16'd5596, 16'd29090, 16'd19710, 16'd48469, 16'd24142, 16'd26124});
	test_expansion(128'h7d40590e78ee9a774c688765005faf2e, {16'd10970, 16'd49886, 16'd21189, 16'd40858, 16'd23133, 16'd12123, 16'd45012, 16'd55729, 16'd53004, 16'd5375, 16'd50772, 16'd17973, 16'd26323, 16'd47080, 16'd28789, 16'd4435, 16'd48830, 16'd50481, 16'd65358, 16'd18427, 16'd63318, 16'd16433, 16'd52486, 16'd34579, 16'd21675, 16'd31163});
	test_expansion(128'h6e7f3e462f1a360c05137a8bec302eb1, {16'd58388, 16'd9901, 16'd29732, 16'd48714, 16'd16696, 16'd62673, 16'd10470, 16'd27630, 16'd37633, 16'd63096, 16'd46895, 16'd30551, 16'd27905, 16'd2178, 16'd60818, 16'd31125, 16'd34100, 16'd58502, 16'd56164, 16'd60028, 16'd7722, 16'd49170, 16'd46522, 16'd12069, 16'd31403, 16'd13787});
	test_expansion(128'heabc933ca4ae216f02e2236a788a5b35, {16'd52210, 16'd16042, 16'd49343, 16'd40179, 16'd64080, 16'd1674, 16'd18229, 16'd42076, 16'd28684, 16'd32121, 16'd30400, 16'd24433, 16'd41922, 16'd50547, 16'd57894, 16'd25344, 16'd14250, 16'd65034, 16'd57049, 16'd5541, 16'd9268, 16'd12194, 16'd29700, 16'd13910, 16'd36292, 16'd8684});
	test_expansion(128'h73bccbaeae5df4f5334ee944f07217eb, {16'd61928, 16'd52101, 16'd65530, 16'd44337, 16'd44704, 16'd37271, 16'd45069, 16'd20173, 16'd58976, 16'd30514, 16'd24418, 16'd46797, 16'd17694, 16'd49468, 16'd3185, 16'd49323, 16'd65033, 16'd52692, 16'd57173, 16'd10471, 16'd43242, 16'd25700, 16'd5710, 16'd39889, 16'd22524, 16'd57954});
	test_expansion(128'h0fee16eb2714aaccb760047f21368415, {16'd14743, 16'd50446, 16'd61656, 16'd44703, 16'd3174, 16'd40419, 16'd17081, 16'd16592, 16'd45764, 16'd47966, 16'd45586, 16'd39593, 16'd7642, 16'd18794, 16'd58952, 16'd60137, 16'd54178, 16'd13023, 16'd9725, 16'd36524, 16'd30559, 16'd7965, 16'd52979, 16'd39378, 16'd58974, 16'd1885});
	test_expansion(128'h40815de697392812685583ff9cd85881, {16'd27256, 16'd61159, 16'd23198, 16'd61901, 16'd48681, 16'd61696, 16'd11827, 16'd30832, 16'd57084, 16'd30970, 16'd19954, 16'd12656, 16'd52144, 16'd31525, 16'd50648, 16'd21387, 16'd24582, 16'd39433, 16'd62718, 16'd27185, 16'd6208, 16'd9465, 16'd6194, 16'd45327, 16'd42802, 16'd33433});
	test_expansion(128'hc850730e10d2c4e35793eb5bd933d4cb, {16'd30916, 16'd2505, 16'd55451, 16'd41437, 16'd21828, 16'd1621, 16'd36148, 16'd57613, 16'd42296, 16'd21929, 16'd5768, 16'd9940, 16'd36767, 16'd55719, 16'd39467, 16'd56413, 16'd39780, 16'd19014, 16'd36985, 16'd42152, 16'd10655, 16'd11223, 16'd50307, 16'd48063, 16'd315, 16'd64607});
	test_expansion(128'hc5eabb6b7fd1bdea2110ec50793e84a7, {16'd44136, 16'd3201, 16'd49861, 16'd8149, 16'd8821, 16'd34665, 16'd21892, 16'd17803, 16'd11511, 16'd20186, 16'd27457, 16'd19553, 16'd22789, 16'd52753, 16'd9826, 16'd65056, 16'd4875, 16'd57132, 16'd6821, 16'd64409, 16'd42758, 16'd47895, 16'd63413, 16'd53556, 16'd44617, 16'd21548});
	test_expansion(128'h4dfdb704f48b64494fc14f83eddc3af0, {16'd30911, 16'd63957, 16'd43658, 16'd43113, 16'd63015, 16'd33125, 16'd618, 16'd40797, 16'd63470, 16'd12140, 16'd49456, 16'd39193, 16'd45189, 16'd18717, 16'd9302, 16'd16436, 16'd59967, 16'd59588, 16'd12250, 16'd63051, 16'd137, 16'd34993, 16'd46922, 16'd21734, 16'd42050, 16'd58284});
	test_expansion(128'h8ee330bf620652e6823b870312006bee, {16'd4, 16'd8286, 16'd14473, 16'd48470, 16'd30033, 16'd40986, 16'd15724, 16'd693, 16'd35427, 16'd40572, 16'd4935, 16'd1089, 16'd5424, 16'd49990, 16'd7425, 16'd35329, 16'd24994, 16'd28771, 16'd5695, 16'd10448, 16'd47388, 16'd56079, 16'd26928, 16'd19140, 16'd29997, 16'd49130});
	test_expansion(128'h1049722a2ba9f8bf54c4c3cd02aaa1e1, {16'd30104, 16'd16205, 16'd1675, 16'd23783, 16'd26901, 16'd41546, 16'd14010, 16'd61296, 16'd16341, 16'd22719, 16'd4818, 16'd49665, 16'd59916, 16'd31942, 16'd38106, 16'd41150, 16'd5468, 16'd44546, 16'd10752, 16'd56973, 16'd41885, 16'd38893, 16'd4472, 16'd16836, 16'd25961, 16'd22599});
	test_expansion(128'h8da79aae8f65d9a7980f7a294e44e748, {16'd34080, 16'd31218, 16'd49245, 16'd29015, 16'd2871, 16'd64173, 16'd51980, 16'd38097, 16'd55121, 16'd9047, 16'd30617, 16'd180, 16'd8035, 16'd18401, 16'd33665, 16'd40543, 16'd38404, 16'd24421, 16'd22931, 16'd35074, 16'd47072, 16'd39349, 16'd21271, 16'd35741, 16'd44158, 16'd11907});
	test_expansion(128'hf86975dc846a953af1bd00c3cc686ee0, {16'd21591, 16'd12404, 16'd55524, 16'd6105, 16'd51456, 16'd31742, 16'd28938, 16'd53557, 16'd42446, 16'd56051, 16'd5756, 16'd9322, 16'd49634, 16'd55666, 16'd55355, 16'd56058, 16'd63461, 16'd23414, 16'd24622, 16'd25735, 16'd7304, 16'd60226, 16'd45741, 16'd38771, 16'd46056, 16'd43720});
	test_expansion(128'hd2f725f106f9581ff5e2916a31ea4bc6, {16'd43522, 16'd41171, 16'd64819, 16'd15077, 16'd49679, 16'd11076, 16'd1605, 16'd64003, 16'd52471, 16'd55057, 16'd29304, 16'd65005, 16'd56094, 16'd1014, 16'd29551, 16'd34799, 16'd57239, 16'd51640, 16'd8402, 16'd3289, 16'd23458, 16'd39945, 16'd59042, 16'd11529, 16'd14311, 16'd61929});
	test_expansion(128'h59955a7946217eb3d1947796bf4ca91e, {16'd29414, 16'd47396, 16'd40929, 16'd53275, 16'd23727, 16'd7841, 16'd4485, 16'd45036, 16'd8379, 16'd3901, 16'd25727, 16'd52135, 16'd61849, 16'd36992, 16'd51650, 16'd53176, 16'd6604, 16'd63140, 16'd61706, 16'd60712, 16'd22046, 16'd61992, 16'd59836, 16'd8341, 16'd56854, 16'd34648});
	test_expansion(128'hd0cb2f3418c169106405151437479072, {16'd59481, 16'd36386, 16'd8598, 16'd25763, 16'd17672, 16'd58137, 16'd16763, 16'd9389, 16'd26552, 16'd58663, 16'd5246, 16'd19517, 16'd19160, 16'd65233, 16'd40972, 16'd41175, 16'd61379, 16'd22883, 16'd7801, 16'd27989, 16'd64638, 16'd64986, 16'd55904, 16'd57945, 16'd18982, 16'd13005});
	test_expansion(128'ha9cb7c6075f518f549b92c9bc76da8e0, {16'd26478, 16'd10725, 16'd17827, 16'd51558, 16'd60943, 16'd44855, 16'd6777, 16'd37970, 16'd65489, 16'd30252, 16'd23401, 16'd60119, 16'd8890, 16'd47056, 16'd2208, 16'd51378, 16'd42191, 16'd63647, 16'd34506, 16'd41527, 16'd57254, 16'd36280, 16'd5228, 16'd52396, 16'd49846, 16'd11883});
	test_expansion(128'h22675c450dd556e3afe3945a211c948a, {16'd58723, 16'd7802, 16'd59791, 16'd29989, 16'd38522, 16'd53337, 16'd57957, 16'd58288, 16'd38026, 16'd46635, 16'd46957, 16'd23952, 16'd26246, 16'd59349, 16'd35481, 16'd64842, 16'd11342, 16'd58643, 16'd15833, 16'd23743, 16'd46467, 16'd23368, 16'd61281, 16'd29034, 16'd9857, 16'd40143});
	test_expansion(128'hcf72ac249b59b402f91623355534a3fc, {16'd20033, 16'd7194, 16'd21295, 16'd63334, 16'd19591, 16'd33351, 16'd62755, 16'd3126, 16'd43413, 16'd62728, 16'd51238, 16'd17556, 16'd23860, 16'd23462, 16'd28953, 16'd38233, 16'd12826, 16'd2771, 16'd26160, 16'd13475, 16'd4637, 16'd21719, 16'd1013, 16'd36821, 16'd17523, 16'd63572});
	test_expansion(128'h0bb26f57bc7831ac8f559c5d0c208ce3, {16'd59113, 16'd40647, 16'd10, 16'd22502, 16'd50887, 16'd11812, 16'd9127, 16'd27856, 16'd44399, 16'd64754, 16'd53867, 16'd2190, 16'd63615, 16'd11763, 16'd54682, 16'd43349, 16'd64544, 16'd52883, 16'd51162, 16'd14116, 16'd33374, 16'd47439, 16'd48404, 16'd53606, 16'd12600, 16'd27421});
	test_expansion(128'h71ee454da2beb553737906a63e76ac34, {16'd13141, 16'd43281, 16'd36454, 16'd38797, 16'd52123, 16'd40765, 16'd54536, 16'd39157, 16'd39004, 16'd36993, 16'd4399, 16'd23687, 16'd56489, 16'd24614, 16'd44532, 16'd56439, 16'd16849, 16'd63055, 16'd40485, 16'd28230, 16'd48358, 16'd54008, 16'd15403, 16'd35219, 16'd29192, 16'd57940});
	test_expansion(128'h620bc891945fb33a6f37260bb9044f6b, {16'd42355, 16'd19037, 16'd30879, 16'd43208, 16'd57003, 16'd5009, 16'd60688, 16'd41482, 16'd11121, 16'd2233, 16'd10972, 16'd29686, 16'd50920, 16'd13077, 16'd8527, 16'd50349, 16'd60742, 16'd53535, 16'd16218, 16'd65258, 16'd18430, 16'd49462, 16'd5186, 16'd11515, 16'd49143, 16'd18492});
	test_expansion(128'h977bcb7b265c5187f6bd51eb3b6d04f2, {16'd47496, 16'd3950, 16'd1346, 16'd27670, 16'd36868, 16'd49663, 16'd29901, 16'd36768, 16'd32011, 16'd56039, 16'd57282, 16'd8235, 16'd22640, 16'd57353, 16'd64862, 16'd13388, 16'd30257, 16'd9170, 16'd63228, 16'd432, 16'd43431, 16'd32321, 16'd8772, 16'd62393, 16'd47612, 16'd31106});
	test_expansion(128'h5f934a259a96e728580a42b402591732, {16'd49985, 16'd37644, 16'd12998, 16'd33655, 16'd62996, 16'd23488, 16'd47273, 16'd25518, 16'd1333, 16'd65048, 16'd63807, 16'd43188, 16'd1472, 16'd43613, 16'd14562, 16'd23399, 16'd41930, 16'd15256, 16'd60711, 16'd35292, 16'd37892, 16'd26619, 16'd38605, 16'd20334, 16'd33475, 16'd27508});
	test_expansion(128'hb8ca8507fd868e56fa991d94aef2982f, {16'd49930, 16'd58838, 16'd54024, 16'd14215, 16'd43848, 16'd52780, 16'd24509, 16'd314, 16'd10898, 16'd49486, 16'd16788, 16'd50121, 16'd17498, 16'd47738, 16'd50634, 16'd9090, 16'd64163, 16'd26049, 16'd55362, 16'd50994, 16'd61462, 16'd33340, 16'd2668, 16'd164, 16'd40526, 16'd7803});
	test_expansion(128'h80b3645329168716f9900841482f3d66, {16'd26240, 16'd27811, 16'd48701, 16'd65144, 16'd37926, 16'd31898, 16'd42204, 16'd27398, 16'd14322, 16'd55941, 16'd35821, 16'd4905, 16'd50417, 16'd13062, 16'd62683, 16'd63634, 16'd50757, 16'd39222, 16'd33886, 16'd49025, 16'd17065, 16'd8610, 16'd22382, 16'd51779, 16'd59388, 16'd32031});
	test_expansion(128'h0b8e5552b8551913caae147124ee3213, {16'd2229, 16'd56120, 16'd33215, 16'd33705, 16'd50353, 16'd674, 16'd50620, 16'd2851, 16'd31933, 16'd37044, 16'd43641, 16'd18704, 16'd34056, 16'd27274, 16'd41569, 16'd32690, 16'd29163, 16'd2753, 16'd43469, 16'd6101, 16'd3004, 16'd41821, 16'd16053, 16'd12250, 16'd38197, 16'd17808});
	test_expansion(128'h108892c37c3d6a035725541d748825fb, {16'd25251, 16'd33944, 16'd28533, 16'd59943, 16'd34783, 16'd58233, 16'd15781, 16'd50621, 16'd56139, 16'd44256, 16'd58409, 16'd13083, 16'd750, 16'd53584, 16'd22269, 16'd56432, 16'd6061, 16'd4019, 16'd22108, 16'd23649, 16'd37737, 16'd33900, 16'd60277, 16'd59228, 16'd45260, 16'd46673});
	test_expansion(128'h8694bd9e7fd3ecc64ba276a17c367ca2, {16'd33215, 16'd24069, 16'd19768, 16'd11080, 16'd50874, 16'd35387, 16'd1980, 16'd48874, 16'd52343, 16'd9519, 16'd9636, 16'd27489, 16'd28927, 16'd23673, 16'd15280, 16'd29186, 16'd30261, 16'd38766, 16'd42621, 16'd4203, 16'd56415, 16'd1442, 16'd37831, 16'd42406, 16'd56319, 16'd27538});
	test_expansion(128'h09e63d84dffb86821c270a303402bdc8, {16'd62965, 16'd46829, 16'd46650, 16'd47831, 16'd39812, 16'd17566, 16'd63735, 16'd21776, 16'd20624, 16'd9268, 16'd59420, 16'd49866, 16'd14397, 16'd4836, 16'd14170, 16'd11113, 16'd56294, 16'd63817, 16'd44064, 16'd45326, 16'd52613, 16'd61766, 16'd53798, 16'd4776, 16'd11898, 16'd62120});
	test_expansion(128'hbf24825e4f4f12fb3f015740f637c744, {16'd16347, 16'd20413, 16'd2832, 16'd48798, 16'd50550, 16'd49243, 16'd38978, 16'd63969, 16'd51229, 16'd52533, 16'd10028, 16'd51131, 16'd21610, 16'd60003, 16'd51518, 16'd13628, 16'd10818, 16'd41969, 16'd33081, 16'd5043, 16'd38967, 16'd29069, 16'd3167, 16'd38363, 16'd28153, 16'd43571});
	test_expansion(128'h4697b3bb9b50884b04031c0792a94e9d, {16'd30301, 16'd38986, 16'd28737, 16'd13703, 16'd3523, 16'd44783, 16'd57148, 16'd42289, 16'd14071, 16'd57943, 16'd26927, 16'd36142, 16'd10910, 16'd11840, 16'd53151, 16'd23620, 16'd46984, 16'd46460, 16'd43194, 16'd26773, 16'd57339, 16'd13028, 16'd34987, 16'd47656, 16'd62282, 16'd59303});
	test_expansion(128'ha642268e1aa4b12b9f0b2a8d23af0ce7, {16'd36412, 16'd24618, 16'd51821, 16'd63357, 16'd10237, 16'd15478, 16'd35809, 16'd23218, 16'd3323, 16'd14005, 16'd47383, 16'd22785, 16'd43309, 16'd44272, 16'd14352, 16'd30988, 16'd53114, 16'd16393, 16'd60990, 16'd24811, 16'd41205, 16'd3282, 16'd40782, 16'd53848, 16'd8841, 16'd24620});
	test_expansion(128'hd2615a0b3e1dfdc03172289ce04accf7, {16'd53594, 16'd62261, 16'd4742, 16'd17969, 16'd48773, 16'd48202, 16'd32920, 16'd11765, 16'd45587, 16'd57368, 16'd40567, 16'd59218, 16'd63263, 16'd41651, 16'd33704, 16'd20099, 16'd22105, 16'd10885, 16'd59589, 16'd26813, 16'd10653, 16'd24950, 16'd1076, 16'd42166, 16'd40835, 16'd60912});
	test_expansion(128'h2eb5616d8029bfd7558adcf155ad11b0, {16'd15692, 16'd64392, 16'd35193, 16'd41266, 16'd45595, 16'd34557, 16'd59214, 16'd30696, 16'd64790, 16'd48249, 16'd55102, 16'd43614, 16'd43484, 16'd38109, 16'd49477, 16'd32307, 16'd26092, 16'd64547, 16'd39412, 16'd53443, 16'd59404, 16'd59255, 16'd53561, 16'd59190, 16'd59475, 16'd24522});
	test_expansion(128'he9bc71e135c08be334b7294fa1165154, {16'd45809, 16'd14556, 16'd4930, 16'd63773, 16'd8188, 16'd49617, 16'd21, 16'd36705, 16'd55272, 16'd29882, 16'd50409, 16'd52603, 16'd38577, 16'd29053, 16'd12187, 16'd56698, 16'd358, 16'd62985, 16'd20229, 16'd56865, 16'd26963, 16'd40059, 16'd47617, 16'd49264, 16'd45514, 16'd18224});
	test_expansion(128'h85ec8d520b0d6fd4b1658bc18717958d, {16'd44369, 16'd52135, 16'd62229, 16'd30291, 16'd17671, 16'd34220, 16'd7458, 16'd58190, 16'd60399, 16'd47083, 16'd55352, 16'd17414, 16'd7239, 16'd24019, 16'd46660, 16'd16979, 16'd7107, 16'd14334, 16'd20200, 16'd35177, 16'd18809, 16'd63879, 16'd26995, 16'd29876, 16'd46240, 16'd63719});
	test_expansion(128'h1e22f963e85f67b538b2bfd22117c60e, {16'd7803, 16'd21276, 16'd19075, 16'd26632, 16'd26143, 16'd37365, 16'd58226, 16'd9493, 16'd9164, 16'd28109, 16'd505, 16'd58642, 16'd32246, 16'd63563, 16'd36476, 16'd53640, 16'd52398, 16'd29281, 16'd39772, 16'd22720, 16'd48992, 16'd62607, 16'd19224, 16'd3918, 16'd20044, 16'd37093});
	test_expansion(128'hec09b7fcfb903d8a0712dbead8c27ef6, {16'd33442, 16'd57368, 16'd45611, 16'd25998, 16'd43841, 16'd1478, 16'd36016, 16'd1416, 16'd50839, 16'd62809, 16'd38333, 16'd4400, 16'd11703, 16'd17721, 16'd26457, 16'd19608, 16'd45291, 16'd54406, 16'd48765, 16'd22627, 16'd62230, 16'd9165, 16'd37786, 16'd31855, 16'd51583, 16'd8025});
	test_expansion(128'h5051f88f7dcb98a1be179bd6b48cacb1, {16'd46923, 16'd63293, 16'd6310, 16'd7934, 16'd37592, 16'd54758, 16'd50430, 16'd13496, 16'd33625, 16'd48947, 16'd42549, 16'd55906, 16'd59407, 16'd47767, 16'd7807, 16'd59274, 16'd33691, 16'd4302, 16'd8274, 16'd7227, 16'd263, 16'd12116, 16'd40816, 16'd1267, 16'd35512, 16'd38733});
	test_expansion(128'h098c0e4a800bf1d33b4a390a399097a7, {16'd28224, 16'd2337, 16'd37194, 16'd61481, 16'd57941, 16'd48248, 16'd17174, 16'd57806, 16'd30138, 16'd5946, 16'd15757, 16'd37115, 16'd62917, 16'd13049, 16'd9765, 16'd38084, 16'd6736, 16'd48049, 16'd4594, 16'd6159, 16'd51783, 16'd36567, 16'd13185, 16'd13356, 16'd51058, 16'd60042});
	test_expansion(128'h983a522f62f8a7185579f9946058214f, {16'd34175, 16'd726, 16'd16573, 16'd14183, 16'd3348, 16'd17615, 16'd31211, 16'd63936, 16'd41284, 16'd35534, 16'd42443, 16'd35811, 16'd54724, 16'd55003, 16'd43226, 16'd57291, 16'd44311, 16'd37397, 16'd50618, 16'd57053, 16'd22296, 16'd21943, 16'd33115, 16'd30911, 16'd63248, 16'd19277});
	test_expansion(128'h6191c03a2541d17a0d7166161afe85f5, {16'd18303, 16'd50435, 16'd10044, 16'd12148, 16'd3029, 16'd48920, 16'd62137, 16'd54015, 16'd26959, 16'd10567, 16'd15273, 16'd14050, 16'd11318, 16'd451, 16'd58601, 16'd4047, 16'd12787, 16'd32142, 16'd29853, 16'd50249, 16'd32934, 16'd53679, 16'd6067, 16'd18092, 16'd48580, 16'd40028});
	test_expansion(128'hb620298054735d65071f78b40baf8174, {16'd29284, 16'd55735, 16'd12058, 16'd56482, 16'd38864, 16'd36984, 16'd56997, 16'd44002, 16'd32801, 16'd15, 16'd18288, 16'd29077, 16'd34443, 16'd21731, 16'd37829, 16'd45838, 16'd8479, 16'd61086, 16'd22675, 16'd48529, 16'd30741, 16'd46949, 16'd22400, 16'd15808, 16'd58961, 16'd34884});
	test_expansion(128'hf76dd9a3a51aa8246e63630f6bc0682e, {16'd39525, 16'd16431, 16'd26509, 16'd57438, 16'd56650, 16'd63257, 16'd48450, 16'd26206, 16'd26056, 16'd40618, 16'd56616, 16'd32623, 16'd12473, 16'd44868, 16'd50215, 16'd51137, 16'd30937, 16'd8343, 16'd28878, 16'd5356, 16'd10712, 16'd43795, 16'd64386, 16'd22906, 16'd18063, 16'd45947});
	test_expansion(128'h01c7f9f99c98312a40590de1192b1f51, {16'd42431, 16'd50120, 16'd47707, 16'd59422, 16'd4056, 16'd24754, 16'd35643, 16'd44353, 16'd28877, 16'd3672, 16'd32116, 16'd10754, 16'd51635, 16'd51111, 16'd53917, 16'd63452, 16'd63084, 16'd51921, 16'd46707, 16'd18146, 16'd49230, 16'd5676, 16'd4742, 16'd40836, 16'd36258, 16'd4892});
	test_expansion(128'h4ea9e350d92dfb809c129114f2ce225b, {16'd19105, 16'd37094, 16'd25471, 16'd19806, 16'd59699, 16'd51432, 16'd4669, 16'd4456, 16'd54149, 16'd29935, 16'd17114, 16'd13929, 16'd15648, 16'd52292, 16'd36106, 16'd23475, 16'd1692, 16'd5904, 16'd4174, 16'd22896, 16'd43168, 16'd21898, 16'd4266, 16'd23935, 16'd15108, 16'd31648});
	test_expansion(128'hcb1da9d8f4ef33b3eaf7aa1781770ada, {16'd39067, 16'd53634, 16'd47344, 16'd37184, 16'd50323, 16'd40768, 16'd3287, 16'd50611, 16'd29322, 16'd58440, 16'd32892, 16'd34179, 16'd64309, 16'd21212, 16'd18545, 16'd46192, 16'd53259, 16'd34550, 16'd10342, 16'd51567, 16'd56904, 16'd61793, 16'd35728, 16'd42329, 16'd2165, 16'd21326});
	test_expansion(128'hd0344d45bae5ba1fe668a57c00d19530, {16'd35067, 16'd45584, 16'd10769, 16'd52463, 16'd31159, 16'd53932, 16'd33655, 16'd19210, 16'd46816, 16'd5213, 16'd36721, 16'd5058, 16'd15540, 16'd570, 16'd13452, 16'd1128, 16'd5491, 16'd5302, 16'd13681, 16'd12035, 16'd14065, 16'd5274, 16'd15943, 16'd28033, 16'd25561, 16'd5327});
	test_expansion(128'hf9ca7a2903204a54bc61e7060675f7b0, {16'd11576, 16'd58996, 16'd1661, 16'd18639, 16'd57522, 16'd6576, 16'd37547, 16'd18973, 16'd25921, 16'd33245, 16'd594, 16'd27857, 16'd44106, 16'd9863, 16'd18585, 16'd13966, 16'd7453, 16'd56362, 16'd12794, 16'd56398, 16'd14706, 16'd43283, 16'd28858, 16'd49885, 16'd26815, 16'd2890});
	test_expansion(128'h728c601626e2a92bb84293f6f365b215, {16'd59179, 16'd31292, 16'd18529, 16'd8449, 16'd30664, 16'd43044, 16'd60809, 16'd41655, 16'd23272, 16'd12929, 16'd26534, 16'd20764, 16'd41224, 16'd6320, 16'd10682, 16'd7277, 16'd57947, 16'd31606, 16'd51595, 16'd43277, 16'd41102, 16'd39600, 16'd49649, 16'd32752, 16'd37090, 16'd51083});
	test_expansion(128'h28efc9ff54e4cc960a19c4d2b6987bf9, {16'd18777, 16'd4672, 16'd59396, 16'd24274, 16'd21094, 16'd37341, 16'd27148, 16'd7447, 16'd39909, 16'd14419, 16'd53370, 16'd14278, 16'd62970, 16'd306, 16'd49643, 16'd3530, 16'd44061, 16'd64812, 16'd5440, 16'd60080, 16'd6182, 16'd46209, 16'd53846, 16'd37044, 16'd56440, 16'd55596});
	test_expansion(128'hb95d0bcf0d644d3da7e89afd0bd1baa0, {16'd47993, 16'd63724, 16'd50544, 16'd32936, 16'd62549, 16'd54591, 16'd15673, 16'd15653, 16'd29116, 16'd42435, 16'd54460, 16'd32576, 16'd62231, 16'd17758, 16'd27923, 16'd19474, 16'd36174, 16'd3048, 16'd7969, 16'd62723, 16'd1947, 16'd61712, 16'd28137, 16'd14106, 16'd18426, 16'd48226});
	test_expansion(128'h5454b5a5f9d6a8477ba3a5f806fb1a9c, {16'd39705, 16'd63198, 16'd40997, 16'd62593, 16'd11452, 16'd54596, 16'd53329, 16'd65329, 16'd64149, 16'd15909, 16'd33806, 16'd42282, 16'd20502, 16'd23878, 16'd31569, 16'd39566, 16'd8499, 16'd18734, 16'd19366, 16'd53681, 16'd18839, 16'd28084, 16'd9741, 16'd3418, 16'd44053, 16'd51329});
	test_expansion(128'h1bd64fd6c3111d27d047616a7964e636, {16'd14389, 16'd16719, 16'd26816, 16'd34475, 16'd29663, 16'd23662, 16'd64923, 16'd58529, 16'd17802, 16'd49871, 16'd35141, 16'd62000, 16'd43097, 16'd54452, 16'd25822, 16'd16200, 16'd20128, 16'd6468, 16'd55363, 16'd40499, 16'd50217, 16'd54024, 16'd27965, 16'd23287, 16'd16914, 16'd6566});
	test_expansion(128'hb5383649e17bb4b87a1a388f8b8ea57e, {16'd59108, 16'd17227, 16'd26010, 16'd26195, 16'd55301, 16'd45530, 16'd35596, 16'd3163, 16'd62235, 16'd11537, 16'd1484, 16'd30715, 16'd20825, 16'd56820, 16'd4511, 16'd38966, 16'd47693, 16'd64742, 16'd15296, 16'd6953, 16'd13381, 16'd41748, 16'd24819, 16'd24295, 16'd47942, 16'd52738});
	test_expansion(128'ha768c58c3e696d1f563f632ff025ff8b, {16'd11840, 16'd40124, 16'd35234, 16'd15412, 16'd23277, 16'd62353, 16'd27180, 16'd33010, 16'd669, 16'd20181, 16'd6800, 16'd41947, 16'd283, 16'd24082, 16'd21060, 16'd59477, 16'd29514, 16'd59470, 16'd51169, 16'd24164, 16'd31232, 16'd39614, 16'd28146, 16'd52291, 16'd61675, 16'd43195});
	test_expansion(128'h54d54e70649e9254d32432bf0872150a, {16'd32208, 16'd62218, 16'd57358, 16'd64280, 16'd1355, 16'd59935, 16'd27246, 16'd53551, 16'd8362, 16'd31436, 16'd42034, 16'd23018, 16'd12695, 16'd60324, 16'd52106, 16'd61657, 16'd23019, 16'd58947, 16'd30305, 16'd20101, 16'd13673, 16'd57905, 16'd59547, 16'd27225, 16'd48130, 16'd16910});
	test_expansion(128'h92807e77a101a89dceb1db1b839db93c, {16'd55023, 16'd24111, 16'd64341, 16'd47507, 16'd55658, 16'd29706, 16'd36290, 16'd16240, 16'd61552, 16'd836, 16'd32711, 16'd37333, 16'd46558, 16'd43376, 16'd14286, 16'd2223, 16'd32407, 16'd30875, 16'd47529, 16'd15842, 16'd15711, 16'd3399, 16'd37875, 16'd51538, 16'd26979, 16'd51719});
	test_expansion(128'hb878c2f46ee636247d102b42cd7bd023, {16'd57406, 16'd24588, 16'd55017, 16'd8595, 16'd43006, 16'd42072, 16'd47405, 16'd11422, 16'd47787, 16'd9463, 16'd19648, 16'd30447, 16'd28917, 16'd45004, 16'd26316, 16'd41244, 16'd21581, 16'd17027, 16'd12288, 16'd41626, 16'd57883, 16'd15130, 16'd15833, 16'd62811, 16'd53611, 16'd50731});
	test_expansion(128'hfd0feae20a64b1611c532af0f4ecb18b, {16'd57631, 16'd5088, 16'd10291, 16'd28904, 16'd48195, 16'd29178, 16'd18358, 16'd41590, 16'd21846, 16'd12415, 16'd23526, 16'd51521, 16'd5290, 16'd25777, 16'd45949, 16'd32723, 16'd29653, 16'd14694, 16'd28039, 16'd60384, 16'd10119, 16'd29234, 16'd7432, 16'd63711, 16'd44745, 16'd47285});
	test_expansion(128'hb27ab682bfe711ec2b36b3eb95912791, {16'd1850, 16'd23679, 16'd64086, 16'd48989, 16'd58495, 16'd16581, 16'd23900, 16'd48789, 16'd18324, 16'd31330, 16'd30442, 16'd27311, 16'd60303, 16'd22593, 16'd24113, 16'd30539, 16'd57725, 16'd44110, 16'd4672, 16'd17336, 16'd17079, 16'd40638, 16'd22460, 16'd56610, 16'd9346, 16'd61370});
	test_expansion(128'h16c8bb9e5cfbe98420ae5b037d31944b, {16'd42159, 16'd46027, 16'd53027, 16'd26737, 16'd30177, 16'd24367, 16'd2307, 16'd62175, 16'd29666, 16'd61312, 16'd58948, 16'd13399, 16'd61948, 16'd30339, 16'd31552, 16'd62179, 16'd46176, 16'd37044, 16'd19668, 16'd11481, 16'd56220, 16'd55846, 16'd32227, 16'd41492, 16'd4428, 16'd51507});
	test_expansion(128'hfc0520eb8eed9f06c09faff95b29b9a7, {16'd56556, 16'd19719, 16'd53785, 16'd5596, 16'd24941, 16'd54147, 16'd42630, 16'd47334, 16'd56016, 16'd974, 16'd51177, 16'd65343, 16'd37938, 16'd1936, 16'd19876, 16'd54725, 16'd23936, 16'd39632, 16'd64469, 16'd59250, 16'd12057, 16'd50876, 16'd36392, 16'd44912, 16'd11684, 16'd2904});
	test_expansion(128'h4945f5791d756a41fa21c490e3ae46d2, {16'd11717, 16'd7306, 16'd11644, 16'd60091, 16'd2487, 16'd34802, 16'd61623, 16'd62207, 16'd10196, 16'd16840, 16'd32871, 16'd28233, 16'd44724, 16'd26490, 16'd20670, 16'd18531, 16'd40066, 16'd63014, 16'd58624, 16'd10922, 16'd4742, 16'd32850, 16'd58185, 16'd46864, 16'd64042, 16'd36738});
	test_expansion(128'heec88360d637e565c3a046802a7063a4, {16'd22468, 16'd14854, 16'd13019, 16'd31177, 16'd38773, 16'd21294, 16'd63533, 16'd33745, 16'd8766, 16'd41753, 16'd33174, 16'd3362, 16'd44313, 16'd8153, 16'd52043, 16'd35931, 16'd52605, 16'd27470, 16'd2462, 16'd37211, 16'd23397, 16'd11692, 16'd63916, 16'd26052, 16'd40968, 16'd60496});
	test_expansion(128'hc0b0d6ca5b9b2233c938281f787ebfb6, {16'd17296, 16'd37584, 16'd24205, 16'd50004, 16'd51250, 16'd63096, 16'd6775, 16'd52670, 16'd383, 16'd64723, 16'd37975, 16'd16752, 16'd28207, 16'd46758, 16'd23176, 16'd13148, 16'd7955, 16'd26295, 16'd10667, 16'd23071, 16'd12103, 16'd14230, 16'd47310, 16'd25871, 16'd60263, 16'd58300});
	test_expansion(128'h90a0e69a0bf8aed3f9cd73cff9e7aaf0, {16'd1298, 16'd5352, 16'd12827, 16'd51692, 16'd17375, 16'd48757, 16'd48895, 16'd62018, 16'd48102, 16'd24057, 16'd51883, 16'd26693, 16'd9540, 16'd13422, 16'd44701, 16'd3484, 16'd44950, 16'd61151, 16'd30676, 16'd30155, 16'd23057, 16'd45217, 16'd3902, 16'd57332, 16'd20985, 16'd50820});
	test_expansion(128'he3c8a835c1f13502fa482c2e050aa8e7, {16'd38124, 16'd29268, 16'd4873, 16'd54782, 16'd29090, 16'd40255, 16'd10262, 16'd60353, 16'd54162, 16'd13514, 16'd40707, 16'd41947, 16'd50822, 16'd7214, 16'd29740, 16'd710, 16'd4655, 16'd4525, 16'd62139, 16'd4436, 16'd11624, 16'd17844, 16'd29190, 16'd62632, 16'd40083, 16'd26458});
	test_expansion(128'h2b8b896d8d3706a6d75ea9c9a97683e1, {16'd1037, 16'd37516, 16'd3034, 16'd31418, 16'd3934, 16'd9748, 16'd27616, 16'd60422, 16'd58337, 16'd31451, 16'd48159, 16'd64015, 16'd53234, 16'd35590, 16'd38145, 16'd44899, 16'd53543, 16'd21779, 16'd28960, 16'd8277, 16'd41119, 16'd57255, 16'd26919, 16'd23595, 16'd49170, 16'd18926});
	test_expansion(128'hc0587275117b3baf52b63970205d989f, {16'd30082, 16'd18850, 16'd1719, 16'd49701, 16'd41194, 16'd61012, 16'd20260, 16'd24600, 16'd17150, 16'd3563, 16'd48369, 16'd33192, 16'd6904, 16'd19702, 16'd55835, 16'd26402, 16'd58026, 16'd21546, 16'd62230, 16'd3206, 16'd51696, 16'd12713, 16'd35288, 16'd11932, 16'd52161, 16'd33007});
	test_expansion(128'hda4b0eacfc0f06022a869250572bb612, {16'd60771, 16'd26898, 16'd64981, 16'd9935, 16'd16460, 16'd16803, 16'd8006, 16'd19833, 16'd41007, 16'd29849, 16'd33188, 16'd20741, 16'd24037, 16'd48781, 16'd27649, 16'd52024, 16'd31450, 16'd26744, 16'd57494, 16'd3722, 16'd38137, 16'd40876, 16'd51308, 16'd53962, 16'd46288, 16'd42689});
	test_expansion(128'ha9f45b0cf63f393822ba9f51065aafe7, {16'd31883, 16'd48366, 16'd55909, 16'd9435, 16'd31760, 16'd37213, 16'd55978, 16'd46422, 16'd11130, 16'd23206, 16'd28774, 16'd43233, 16'd61008, 16'd44612, 16'd20143, 16'd22603, 16'd45671, 16'd23522, 16'd20424, 16'd13480, 16'd26234, 16'd45016, 16'd35714, 16'd4269, 16'd34664, 16'd35272});
	test_expansion(128'h3c868e7d7093629e258c0462b26a5ab3, {16'd54508, 16'd393, 16'd59352, 16'd23242, 16'd3084, 16'd64039, 16'd37976, 16'd8079, 16'd33648, 16'd20380, 16'd1426, 16'd7590, 16'd25932, 16'd17389, 16'd10665, 16'd52354, 16'd18613, 16'd38057, 16'd53341, 16'd3957, 16'd28098, 16'd30863, 16'd18955, 16'd24639, 16'd22772, 16'd65355});
	test_expansion(128'h823c904c77835abca696f6f2d94f2ec4, {16'd61298, 16'd2508, 16'd54892, 16'd5179, 16'd55048, 16'd38065, 16'd467, 16'd2849, 16'd35553, 16'd29739, 16'd35962, 16'd32136, 16'd59613, 16'd29250, 16'd55519, 16'd55026, 16'd41435, 16'd53842, 16'd49219, 16'd20719, 16'd35018, 16'd25817, 16'd51165, 16'd61925, 16'd32532, 16'd18599});
	test_expansion(128'h8f750dcb777bb8e07a2c2cf3b97a6c32, {16'd38296, 16'd43448, 16'd29540, 16'd65430, 16'd6368, 16'd50220, 16'd6699, 16'd57523, 16'd57931, 16'd55111, 16'd50531, 16'd4187, 16'd50360, 16'd45321, 16'd36135, 16'd54407, 16'd13618, 16'd37452, 16'd8578, 16'd32474, 16'd54407, 16'd61601, 16'd40069, 16'd55493, 16'd2233, 16'd25572});
	test_expansion(128'h0b8f5a6943985c6a5a3f69711e0d5389, {16'd30595, 16'd10491, 16'd11234, 16'd62607, 16'd21394, 16'd313, 16'd61374, 16'd39072, 16'd40991, 16'd42557, 16'd28694, 16'd9285, 16'd12451, 16'd43872, 16'd34908, 16'd42367, 16'd31996, 16'd29842, 16'd58472, 16'd7610, 16'd44632, 16'd50222, 16'd36207, 16'd45699, 16'd52981, 16'd56498});
	test_expansion(128'hc8cab5c4221d452c80c0c10a433e96f2, {16'd29258, 16'd55163, 16'd60179, 16'd57021, 16'd51015, 16'd33188, 16'd3817, 16'd39894, 16'd20229, 16'd29576, 16'd36387, 16'd53460, 16'd49729, 16'd16356, 16'd27284, 16'd63052, 16'd9138, 16'd54207, 16'd36020, 16'd52686, 16'd5115, 16'd40516, 16'd34641, 16'd51195, 16'd58132, 16'd56969});
	test_expansion(128'h4d85facc0528f4d69563b4be562f7a35, {16'd19025, 16'd53578, 16'd34260, 16'd40960, 16'd9103, 16'd39391, 16'd37275, 16'd36824, 16'd50620, 16'd20744, 16'd56319, 16'd29764, 16'd41172, 16'd57733, 16'd56160, 16'd12154, 16'd27102, 16'd15881, 16'd304, 16'd44330, 16'd4608, 16'd10924, 16'd47815, 16'd45691, 16'd11374, 16'd4105});
	test_expansion(128'hc509e0b0de08a93b6d55dc825d55e690, {16'd8692, 16'd64969, 16'd55721, 16'd21428, 16'd18291, 16'd36372, 16'd61850, 16'd27475, 16'd36340, 16'd14058, 16'd40920, 16'd14448, 16'd23883, 16'd25747, 16'd54830, 16'd53653, 16'd61910, 16'd49554, 16'd41399, 16'd45600, 16'd37532, 16'd32653, 16'd16992, 16'd25509, 16'd16602, 16'd28268});
	test_expansion(128'haa729280db52dc906538ffdee3454049, {16'd60535, 16'd30548, 16'd31491, 16'd31433, 16'd6856, 16'd45079, 16'd45402, 16'd58604, 16'd58788, 16'd37961, 16'd39254, 16'd37265, 16'd32182, 16'd7050, 16'd3776, 16'd30141, 16'd37794, 16'd42567, 16'd9820, 16'd58100, 16'd41479, 16'd30197, 16'd59402, 16'd41783, 16'd37341, 16'd56721});
	test_expansion(128'h127049f39fbbb6fe26fc3de13a25c345, {16'd35941, 16'd51294, 16'd38629, 16'd27637, 16'd65001, 16'd46301, 16'd50471, 16'd43089, 16'd32123, 16'd23214, 16'd58095, 16'd672, 16'd49038, 16'd57644, 16'd62036, 16'd63894, 16'd20972, 16'd39614, 16'd42961, 16'd37949, 16'd40184, 16'd17105, 16'd16232, 16'd31710, 16'd22514, 16'd60959});
	test_expansion(128'h4171cb45d6fc2ad18ad219ecdaaad023, {16'd26311, 16'd64839, 16'd35495, 16'd38399, 16'd34405, 16'd4807, 16'd36377, 16'd27883, 16'd17940, 16'd57525, 16'd40198, 16'd60174, 16'd4949, 16'd29812, 16'd46042, 16'd11752, 16'd2454, 16'd45604, 16'd4565, 16'd49712, 16'd36251, 16'd37445, 16'd18616, 16'd13642, 16'd4904, 16'd35868});
	test_expansion(128'hcc897615f4322c979fdf3ef6b292aa67, {16'd2286, 16'd14959, 16'd36117, 16'd29018, 16'd36283, 16'd57999, 16'd926, 16'd31884, 16'd6233, 16'd15770, 16'd63827, 16'd33758, 16'd34945, 16'd25440, 16'd60992, 16'd40348, 16'd49213, 16'd37332, 16'd41106, 16'd12928, 16'd58013, 16'd54430, 16'd58139, 16'd4382, 16'd42864, 16'd2898});
	test_expansion(128'ha0b11de7b3b2e5b5eb1181f659e2df52, {16'd19504, 16'd55791, 16'd7910, 16'd39322, 16'd24544, 16'd63638, 16'd10984, 16'd48705, 16'd14067, 16'd38072, 16'd61567, 16'd38685, 16'd20154, 16'd23300, 16'd54779, 16'd45702, 16'd10464, 16'd8743, 16'd47292, 16'd23047, 16'd62859, 16'd52512, 16'd20391, 16'd3119, 16'd22110, 16'd5925});
	test_expansion(128'h334f8ac1541f2904e9b7a33eae455724, {16'd44939, 16'd62743, 16'd28380, 16'd16091, 16'd40949, 16'd46672, 16'd33427, 16'd27483, 16'd48560, 16'd35524, 16'd8711, 16'd50038, 16'd26855, 16'd17122, 16'd12257, 16'd11278, 16'd35561, 16'd19464, 16'd41276, 16'd12998, 16'd41514, 16'd34591, 16'd26096, 16'd34254, 16'd29022, 16'd58003});
	test_expansion(128'h8863fc2b0f6115a0affb7e45cac97dd1, {16'd55256, 16'd52763, 16'd15422, 16'd22339, 16'd15576, 16'd41352, 16'd3865, 16'd52020, 16'd52575, 16'd54728, 16'd2003, 16'd35308, 16'd907, 16'd61162, 16'd47895, 16'd23197, 16'd18955, 16'd38282, 16'd42064, 16'd6293, 16'd2149, 16'd9908, 16'd32476, 16'd33960, 16'd24053, 16'd17557});
	test_expansion(128'he001aee0aeee6fa37f666215b3ce0d73, {16'd43435, 16'd43494, 16'd2711, 16'd18811, 16'd19516, 16'd26441, 16'd30040, 16'd13981, 16'd35030, 16'd20464, 16'd38498, 16'd17626, 16'd30283, 16'd8946, 16'd29945, 16'd13146, 16'd3029, 16'd32489, 16'd32934, 16'd50705, 16'd10745, 16'd22152, 16'd21164, 16'd38233, 16'd64899, 16'd12418});
	test_expansion(128'h6189e93279658ed6951111a6aa362f9d, {16'd9355, 16'd30120, 16'd17777, 16'd17569, 16'd33206, 16'd5235, 16'd9077, 16'd47373, 16'd4760, 16'd42225, 16'd47405, 16'd47874, 16'd15327, 16'd53861, 16'd56173, 16'd10870, 16'd22917, 16'd34829, 16'd64884, 16'd532, 16'd6007, 16'd10544, 16'd37418, 16'd32708, 16'd52708, 16'd24372});
	test_expansion(128'h385c858c9baca589203ca1bf35c2f634, {16'd33097, 16'd44875, 16'd54030, 16'd22264, 16'd24918, 16'd22940, 16'd23083, 16'd39355, 16'd21805, 16'd54243, 16'd15546, 16'd1916, 16'd52355, 16'd30368, 16'd7017, 16'd48676, 16'd37793, 16'd58732, 16'd48103, 16'd36753, 16'd47794, 16'd46189, 16'd31565, 16'd52435, 16'd30771, 16'd27473});
	test_expansion(128'hf457cb6e83ec9f715ae90a4390da2961, {16'd57573, 16'd35021, 16'd5782, 16'd34649, 16'd10929, 16'd31639, 16'd41083, 16'd9298, 16'd8046, 16'd12039, 16'd39221, 16'd23559, 16'd60394, 16'd37118, 16'd64190, 16'd1865, 16'd14436, 16'd46836, 16'd38320, 16'd48999, 16'd46403, 16'd8568, 16'd13828, 16'd49927, 16'd64479, 16'd45484});
	test_expansion(128'h4cc257abf8df5c2cc7d17c3fc4cd536c, {16'd63599, 16'd34701, 16'd38781, 16'd58267, 16'd13407, 16'd7209, 16'd51393, 16'd22110, 16'd40003, 16'd40098, 16'd26342, 16'd43817, 16'd16661, 16'd50303, 16'd52950, 16'd22002, 16'd10945, 16'd3819, 16'd55659, 16'd32525, 16'd49441, 16'd39928, 16'd10512, 16'd10848, 16'd10954, 16'd26892});
	test_expansion(128'he162250a0e4beb5335342b27692066f1, {16'd46602, 16'd41316, 16'd45033, 16'd37209, 16'd12131, 16'd40145, 16'd30026, 16'd52497, 16'd9177, 16'd32474, 16'd65107, 16'd6397, 16'd29428, 16'd32840, 16'd25445, 16'd53863, 16'd51079, 16'd25236, 16'd25981, 16'd7465, 16'd46629, 16'd47585, 16'd14023, 16'd27072, 16'd34478, 16'd58555});
	test_expansion(128'hd93e5b4091450ea6f496c173025f5a90, {16'd54024, 16'd14197, 16'd23636, 16'd62346, 16'd50928, 16'd47224, 16'd36845, 16'd61046, 16'd64570, 16'd19095, 16'd19222, 16'd52250, 16'd52312, 16'd26702, 16'd30495, 16'd51853, 16'd31375, 16'd51439, 16'd61391, 16'd33973, 16'd13606, 16'd3724, 16'd18597, 16'd58577, 16'd36538, 16'd20423});
	test_expansion(128'h5a6f17b3f4d639d282de83eae80f88b1, {16'd15678, 16'd2683, 16'd6424, 16'd11554, 16'd60617, 16'd40863, 16'd44802, 16'd31270, 16'd31907, 16'd50233, 16'd10762, 16'd21336, 16'd18924, 16'd31081, 16'd10583, 16'd47360, 16'd35778, 16'd11112, 16'd3104, 16'd26668, 16'd30542, 16'd45235, 16'd16775, 16'd51954, 16'd52438, 16'd4717});
	test_expansion(128'hf7e4e9c68c60d612d59a6a3eaf61f444, {16'd22415, 16'd15778, 16'd33627, 16'd50714, 16'd16691, 16'd3726, 16'd5955, 16'd15084, 16'd49706, 16'd45015, 16'd20354, 16'd25112, 16'd62535, 16'd42414, 16'd22190, 16'd58774, 16'd12354, 16'd36827, 16'd31750, 16'd61387, 16'd57794, 16'd23923, 16'd55164, 16'd2657, 16'd47183, 16'd49626});
	test_expansion(128'hbd38836ef985afe5af67931b30efdea4, {16'd45235, 16'd22300, 16'd47996, 16'd59175, 16'd64689, 16'd19697, 16'd15764, 16'd24923, 16'd22204, 16'd16280, 16'd42268, 16'd7440, 16'd32559, 16'd43625, 16'd42591, 16'd6851, 16'd6593, 16'd12037, 16'd31354, 16'd59664, 16'd50789, 16'd18966, 16'd7563, 16'd43642, 16'd25773, 16'd50747});
	test_expansion(128'h9ba246710812c7f8e230035159354041, {16'd4264, 16'd30671, 16'd3921, 16'd54192, 16'd61237, 16'd18307, 16'd11075, 16'd46183, 16'd54838, 16'd34020, 16'd59774, 16'd3557, 16'd32056, 16'd62332, 16'd20242, 16'd34545, 16'd16779, 16'd29102, 16'd25322, 16'd14416, 16'd56939, 16'd52925, 16'd1641, 16'd50480, 16'd17468, 16'd64585});
	test_expansion(128'h50a05072e3bf4059b1276ca2eb764087, {16'd17713, 16'd10317, 16'd5583, 16'd13130, 16'd36783, 16'd45200, 16'd52601, 16'd56705, 16'd17236, 16'd4618, 16'd12404, 16'd58006, 16'd18957, 16'd39567, 16'd1164, 16'd26060, 16'd32684, 16'd63315, 16'd62003, 16'd49022, 16'd55383, 16'd367, 16'd41340, 16'd29321, 16'd63378, 16'd15821});
	test_expansion(128'h5739240a5ae667c23cb534916cdd6f66, {16'd63185, 16'd8070, 16'd21347, 16'd54669, 16'd36743, 16'd48326, 16'd49006, 16'd22405, 16'd45548, 16'd25809, 16'd51615, 16'd52230, 16'd13593, 16'd41996, 16'd49327, 16'd11736, 16'd42989, 16'd43627, 16'd9554, 16'd41898, 16'd60692, 16'd58876, 16'd53842, 16'd59384, 16'd12338, 16'd26035});
	test_expansion(128'h9da4a05f4088d310e9af2cecd4336906, {16'd38058, 16'd20844, 16'd22289, 16'd21241, 16'd8577, 16'd20094, 16'd16742, 16'd54791, 16'd28435, 16'd7112, 16'd51936, 16'd24151, 16'd42443, 16'd15508, 16'd29778, 16'd42235, 16'd45325, 16'd55641, 16'd59437, 16'd51025, 16'd10527, 16'd21113, 16'd16083, 16'd39878, 16'd51411, 16'd25878});
	test_expansion(128'h67768cc30a39989e8f55b20fdf71780a, {16'd8587, 16'd56711, 16'd41072, 16'd8597, 16'd52413, 16'd23197, 16'd36589, 16'd35893, 16'd42056, 16'd18050, 16'd21097, 16'd13877, 16'd3929, 16'd18181, 16'd7848, 16'd13268, 16'd32417, 16'd53834, 16'd9792, 16'd53774, 16'd8341, 16'd18712, 16'd290, 16'd58192, 16'd9508, 16'd61038});
	test_expansion(128'h49d1be2ad6f1e3c5c07339de8290ebaa, {16'd38615, 16'd25826, 16'd4311, 16'd50838, 16'd46586, 16'd37965, 16'd26478, 16'd27062, 16'd41724, 16'd52347, 16'd30455, 16'd46135, 16'd12569, 16'd17187, 16'd42197, 16'd64295, 16'd32742, 16'd41401, 16'd40162, 16'd8162, 16'd58883, 16'd9596, 16'd45515, 16'd37633, 16'd28868, 16'd7725});
	test_expansion(128'hfd948b5547b982b9a6f071fd557d4749, {16'd19277, 16'd125, 16'd43479, 16'd14104, 16'd38899, 16'd41356, 16'd10523, 16'd64346, 16'd26215, 16'd56859, 16'd26389, 16'd57579, 16'd61850, 16'd31024, 16'd40432, 16'd3012, 16'd47480, 16'd23950, 16'd31060, 16'd9045, 16'd26445, 16'd16695, 16'd50392, 16'd61826, 16'd9678, 16'd22482});
	test_expansion(128'hdc5a6a1a4ae3aa8e338363b0fb4cf767, {16'd31858, 16'd50794, 16'd7065, 16'd35295, 16'd26730, 16'd24535, 16'd46920, 16'd17628, 16'd35071, 16'd45689, 16'd9984, 16'd28258, 16'd46827, 16'd16309, 16'd64034, 16'd11844, 16'd30537, 16'd23312, 16'd9795, 16'd33579, 16'd57465, 16'd47663, 16'd38276, 16'd9966, 16'd14398, 16'd16177});
	test_expansion(128'h8c57f3731337d9658534b4735f8581b2, {16'd27849, 16'd45716, 16'd60332, 16'd20906, 16'd33749, 16'd52701, 16'd60839, 16'd11555, 16'd35218, 16'd20844, 16'd20651, 16'd53245, 16'd36356, 16'd54352, 16'd43155, 16'd56029, 16'd24220, 16'd24672, 16'd20267, 16'd26959, 16'd42760, 16'd15017, 16'd53115, 16'd4452, 16'd12216, 16'd58756});
	test_expansion(128'hb343ce35eba223c5c2a68d1123f9bea6, {16'd11991, 16'd60945, 16'd46418, 16'd61190, 16'd29260, 16'd53280, 16'd1594, 16'd59418, 16'd27042, 16'd34187, 16'd5197, 16'd49985, 16'd60859, 16'd13931, 16'd61733, 16'd40823, 16'd43456, 16'd59718, 16'd13667, 16'd56882, 16'd8749, 16'd50597, 16'd6792, 16'd52968, 16'd62866, 16'd16338});
	test_expansion(128'h86b135cd89a1f7521934322d573531e0, {16'd42563, 16'd55777, 16'd56296, 16'd49170, 16'd14280, 16'd46643, 16'd6817, 16'd15003, 16'd2927, 16'd20390, 16'd27639, 16'd32198, 16'd48824, 16'd55150, 16'd14070, 16'd59676, 16'd54241, 16'd64336, 16'd19632, 16'd12121, 16'd17866, 16'd21548, 16'd53672, 16'd10006, 16'd11877, 16'd5222});
	test_expansion(128'h0a40cb64c2da80f0c162d6eb85db0bc5, {16'd37951, 16'd865, 16'd14941, 16'd4586, 16'd3552, 16'd22011, 16'd9900, 16'd47383, 16'd13522, 16'd27011, 16'd36360, 16'd64632, 16'd40548, 16'd49027, 16'd49488, 16'd31284, 16'd29315, 16'd46105, 16'd64475, 16'd43912, 16'd29878, 16'd57508, 16'd2220, 16'd38327, 16'd30385, 16'd26688});
	test_expansion(128'hced5e922e1797e0756e8d3914708a51d, {16'd29782, 16'd28377, 16'd43860, 16'd19026, 16'd65034, 16'd36424, 16'd23074, 16'd28542, 16'd55597, 16'd16793, 16'd15423, 16'd34581, 16'd48334, 16'd10381, 16'd5888, 16'd55548, 16'd34160, 16'd17032, 16'd51948, 16'd5864, 16'd5311, 16'd64754, 16'd45375, 16'd52341, 16'd44786, 16'd2047});
	test_expansion(128'h3732c80297e074413a004dc73ee0fb0b, {16'd31441, 16'd45157, 16'd4518, 16'd22778, 16'd55577, 16'd62002, 16'd37683, 16'd65245, 16'd47054, 16'd64007, 16'd1740, 16'd50101, 16'd3918, 16'd57629, 16'd23892, 16'd15952, 16'd19511, 16'd33006, 16'd38088, 16'd58203, 16'd46155, 16'd43897, 16'd19551, 16'd8680, 16'd2312, 16'd49676});
	test_expansion(128'hf2219993bb4aaae991a83df296e12e71, {16'd61235, 16'd29925, 16'd25128, 16'd45434, 16'd21243, 16'd58480, 16'd49108, 16'd44993, 16'd10890, 16'd64830, 16'd32732, 16'd3820, 16'd51959, 16'd26410, 16'd54083, 16'd24516, 16'd10022, 16'd34196, 16'd54404, 16'd14584, 16'd63566, 16'd14243, 16'd10953, 16'd42238, 16'd43584, 16'd21892});
	test_expansion(128'h5ab08572bc1a38fd537ae98041417f36, {16'd44679, 16'd28824, 16'd10594, 16'd14071, 16'd4145, 16'd12284, 16'd58081, 16'd4446, 16'd20986, 16'd50264, 16'd45690, 16'd35349, 16'd24012, 16'd50035, 16'd49343, 16'd9763, 16'd28295, 16'd44025, 16'd38368, 16'd59229, 16'd526, 16'd40456, 16'd57624, 16'd64263, 16'd34858, 16'd63952});
	test_expansion(128'hf0fb227b855f4888abfb57c865d50d73, {16'd55324, 16'd62537, 16'd13923, 16'd8385, 16'd60134, 16'd34885, 16'd57891, 16'd31593, 16'd27929, 16'd25152, 16'd29561, 16'd45716, 16'd61766, 16'd54203, 16'd7639, 16'd4007, 16'd51088, 16'd4077, 16'd36052, 16'd27221, 16'd16826, 16'd12820, 16'd39641, 16'd59266, 16'd52506, 16'd47634});
	test_expansion(128'h5508ec9be180c3a89ae60e582de15c25, {16'd2055, 16'd38832, 16'd13664, 16'd27068, 16'd41067, 16'd42115, 16'd31927, 16'd56090, 16'd8890, 16'd42428, 16'd6981, 16'd62230, 16'd10482, 16'd22311, 16'd36862, 16'd21380, 16'd17832, 16'd17231, 16'd45170, 16'd60650, 16'd28240, 16'd17943, 16'd29962, 16'd64898, 16'd4978, 16'd16636});
	test_expansion(128'h2416c19041c5f3b2be9c50063f7862c5, {16'd31976, 16'd43117, 16'd23561, 16'd12559, 16'd6276, 16'd32649, 16'd26164, 16'd53647, 16'd59395, 16'd43550, 16'd7517, 16'd58119, 16'd49260, 16'd43548, 16'd64010, 16'd53129, 16'd20527, 16'd59583, 16'd55358, 16'd40391, 16'd29797, 16'd19715, 16'd49047, 16'd47127, 16'd41209, 16'd7311});
	test_expansion(128'h45a5284481b76a408cd1c3311a948d41, {16'd16083, 16'd3245, 16'd17467, 16'd48245, 16'd11636, 16'd58623, 16'd54253, 16'd8546, 16'd61483, 16'd50975, 16'd50073, 16'd34329, 16'd31177, 16'd32730, 16'd16011, 16'd47728, 16'd7496, 16'd22793, 16'd6621, 16'd23527, 16'd16779, 16'd61378, 16'd63549, 16'd1986, 16'd1597, 16'd11116});
	test_expansion(128'hf6cb34b986f072944cd3c93a3ed57802, {16'd47464, 16'd31560, 16'd24035, 16'd22573, 16'd47705, 16'd59514, 16'd54450, 16'd26034, 16'd41903, 16'd51466, 16'd64646, 16'd4065, 16'd64359, 16'd3901, 16'd43343, 16'd17138, 16'd46312, 16'd9393, 16'd12649, 16'd29192, 16'd27230, 16'd18325, 16'd23153, 16'd3564, 16'd47298, 16'd23127});
	test_expansion(128'h7e7e973955f35be7ff493199613d8694, {16'd6039, 16'd2344, 16'd59183, 16'd9231, 16'd51677, 16'd25147, 16'd63625, 16'd30560, 16'd9096, 16'd60396, 16'd16826, 16'd59420, 16'd38987, 16'd18283, 16'd55503, 16'd5419, 16'd62085, 16'd23512, 16'd40464, 16'd42393, 16'd52748, 16'd2088, 16'd62071, 16'd51754, 16'd40035, 16'd40188});
	test_expansion(128'h41286ddf3e2e47e9ef1adea839502f54, {16'd56178, 16'd32129, 16'd16298, 16'd9860, 16'd62973, 16'd49073, 16'd44836, 16'd17134, 16'd60411, 16'd32929, 16'd16926, 16'd242, 16'd23580, 16'd59677, 16'd4896, 16'd12376, 16'd34619, 16'd33501, 16'd6672, 16'd21412, 16'd52113, 16'd45837, 16'd70, 16'd50071, 16'd25286, 16'd64227});
	test_expansion(128'h1f94ae3260277ffd8633200acf163a0c, {16'd36193, 16'd63496, 16'd2250, 16'd44440, 16'd17027, 16'd42298, 16'd8054, 16'd23726, 16'd16905, 16'd15532, 16'd350, 16'd64535, 16'd42400, 16'd38067, 16'd44306, 16'd34988, 16'd48797, 16'd49670, 16'd1668, 16'd3685, 16'd54318, 16'd18372, 16'd17229, 16'd51438, 16'd42533, 16'd166});
	test_expansion(128'ha2572312672e4d8a48e4f56ed0898537, {16'd47930, 16'd13037, 16'd60823, 16'd24036, 16'd58410, 16'd24531, 16'd51839, 16'd27015, 16'd350, 16'd29091, 16'd52527, 16'd62918, 16'd50036, 16'd52352, 16'd50320, 16'd42165, 16'd48654, 16'd55090, 16'd8892, 16'd49005, 16'd3054, 16'd43518, 16'd50392, 16'd34864, 16'd16976, 16'd49185});
	test_expansion(128'h019e5c23962b4d89f66bf4b986d6f9ba, {16'd46605, 16'd47420, 16'd30859, 16'd18834, 16'd55337, 16'd41400, 16'd43357, 16'd13306, 16'd46889, 16'd22529, 16'd2591, 16'd57356, 16'd45072, 16'd22957, 16'd42704, 16'd48067, 16'd35944, 16'd109, 16'd21754, 16'd8658, 16'd64886, 16'd63562, 16'd53052, 16'd18711, 16'd53160, 16'd50606});
	test_expansion(128'h19aa3d2bd8906639c299fdc8e4204e1b, {16'd1583, 16'd13279, 16'd63163, 16'd12750, 16'd59052, 16'd599, 16'd7971, 16'd44579, 16'd5300, 16'd12103, 16'd62879, 16'd19428, 16'd16096, 16'd22483, 16'd45979, 16'd6053, 16'd46136, 16'd8019, 16'd54668, 16'd10269, 16'd6969, 16'd12635, 16'd40894, 16'd43028, 16'd21368, 16'd40117});
	test_expansion(128'hc81f30dd69ce4ed6d8d3664e55264a2b, {16'd18379, 16'd59774, 16'd33738, 16'd20859, 16'd57629, 16'd3485, 16'd25706, 16'd52413, 16'd15614, 16'd6425, 16'd29600, 16'd7918, 16'd9524, 16'd3360, 16'd1334, 16'd27019, 16'd6406, 16'd44583, 16'd32106, 16'd21853, 16'd38696, 16'd36288, 16'd56889, 16'd551, 16'd52154, 16'd18941});
	test_expansion(128'hb01d895c8c7db9e319c6854565b0906e, {16'd62458, 16'd41290, 16'd12646, 16'd34151, 16'd30813, 16'd7507, 16'd18084, 16'd40466, 16'd32916, 16'd49003, 16'd29845, 16'd4311, 16'd14023, 16'd53757, 16'd28493, 16'd8367, 16'd57396, 16'd64351, 16'd47545, 16'd27177, 16'd28427, 16'd65521, 16'd34703, 16'd64354, 16'd56536, 16'd25902});
	test_expansion(128'h32973df925250494050adaee6bcfd12e, {16'd61571, 16'd41497, 16'd51886, 16'd25831, 16'd15832, 16'd32344, 16'd37068, 16'd32697, 16'd53040, 16'd20958, 16'd11038, 16'd46134, 16'd49017, 16'd50004, 16'd25029, 16'd59003, 16'd2165, 16'd17549, 16'd57395, 16'd11662, 16'd54670, 16'd62287, 16'd26428, 16'd6271, 16'd8216, 16'd47641});
	test_expansion(128'h81a791637776841130551276b768f982, {16'd8726, 16'd38485, 16'd37061, 16'd21731, 16'd27705, 16'd32392, 16'd22071, 16'd41375, 16'd39554, 16'd39314, 16'd42473, 16'd23230, 16'd21770, 16'd17048, 16'd20052, 16'd61560, 16'd8161, 16'd19566, 16'd54957, 16'd62002, 16'd56456, 16'd25575, 16'd20546, 16'd59294, 16'd29876, 16'd20501});
	test_expansion(128'hbf1d5f81755cf151a50b8eceef2296f5, {16'd22373, 16'd26304, 16'd57655, 16'd41262, 16'd12445, 16'd25686, 16'd4437, 16'd16006, 16'd25981, 16'd40010, 16'd12666, 16'd26268, 16'd63200, 16'd49086, 16'd9719, 16'd63997, 16'd38760, 16'd7072, 16'd60939, 16'd53058, 16'd37151, 16'd14103, 16'd58289, 16'd27470, 16'd4700, 16'd7000});
	test_expansion(128'ha9fc246242239d24819b4355de85762a, {16'd33210, 16'd48654, 16'd49300, 16'd32181, 16'd42335, 16'd62589, 16'd31518, 16'd11605, 16'd26584, 16'd23614, 16'd24664, 16'd28070, 16'd21327, 16'd63570, 16'd54110, 16'd22355, 16'd36892, 16'd23120, 16'd55762, 16'd52750, 16'd47747, 16'd47712, 16'd1491, 16'd38854, 16'd526, 16'd15747});
	test_expansion(128'h7ef81e55224eea0832030d430fa21c4f, {16'd46736, 16'd23282, 16'd7287, 16'd52819, 16'd52422, 16'd57095, 16'd8691, 16'd45645, 16'd60259, 16'd28989, 16'd770, 16'd36476, 16'd52058, 16'd28549, 16'd46415, 16'd21491, 16'd42914, 16'd38926, 16'd36318, 16'd52896, 16'd29260, 16'd732, 16'd56883, 16'd22608, 16'd24083, 16'd36796});
	test_expansion(128'h3ff2301e3e6ce7f1c07e212057986dd0, {16'd48876, 16'd2456, 16'd7090, 16'd28681, 16'd4728, 16'd63812, 16'd62278, 16'd31216, 16'd37542, 16'd3889, 16'd58760, 16'd48029, 16'd43147, 16'd53175, 16'd41412, 16'd25043, 16'd16163, 16'd4787, 16'd47229, 16'd35698, 16'd65056, 16'd63687, 16'd47657, 16'd17601, 16'd12027, 16'd52393});
	test_expansion(128'ha12b075dbbf0776b14399e9a01390324, {16'd35251, 16'd52945, 16'd18273, 16'd39813, 16'd13992, 16'd10901, 16'd28995, 16'd49483, 16'd44618, 16'd2181, 16'd47176, 16'd30987, 16'd53604, 16'd40981, 16'd45636, 16'd6816, 16'd14120, 16'd33220, 16'd20020, 16'd46183, 16'd13550, 16'd13854, 16'd43077, 16'd12903, 16'd52275, 16'd7046});
	test_expansion(128'h49247100c706abe3e37fbe9d3adbee66, {16'd13684, 16'd48524, 16'd42093, 16'd62255, 16'd37515, 16'd50310, 16'd13100, 16'd34201, 16'd37233, 16'd28350, 16'd35513, 16'd64217, 16'd25058, 16'd51292, 16'd50414, 16'd13085, 16'd61620, 16'd55778, 16'd50638, 16'd48721, 16'd10006, 16'd40189, 16'd33921, 16'd29436, 16'd20771, 16'd6511});
	test_expansion(128'h6624679d52f0d073c3c030cddd3a1c7c, {16'd59134, 16'd4910, 16'd12180, 16'd15931, 16'd11438, 16'd65448, 16'd21909, 16'd56044, 16'd92, 16'd1391, 16'd48802, 16'd26845, 16'd19725, 16'd57385, 16'd57930, 16'd46335, 16'd50182, 16'd62173, 16'd46476, 16'd49240, 16'd47833, 16'd38748, 16'd16882, 16'd26548, 16'd37924, 16'd41847});
	test_expansion(128'h8ea30440b2d92d46d7640606067d9547, {16'd35535, 16'd64031, 16'd5345, 16'd65439, 16'd4147, 16'd22159, 16'd24085, 16'd5693, 16'd3526, 16'd32691, 16'd726, 16'd13066, 16'd40146, 16'd16586, 16'd28662, 16'd55946, 16'd36154, 16'd17021, 16'd1298, 16'd15466, 16'd41988, 16'd35282, 16'd42058, 16'd16247, 16'd426, 16'd16394});
	test_expansion(128'h5e9a3e52ffc7e0239b931185d67d8a53, {16'd26572, 16'd53771, 16'd51217, 16'd45036, 16'd22999, 16'd24354, 16'd50859, 16'd56264, 16'd23093, 16'd47782, 16'd28710, 16'd1408, 16'd26377, 16'd37088, 16'd9179, 16'd34865, 16'd9591, 16'd63666, 16'd9196, 16'd64306, 16'd44641, 16'd43421, 16'd46181, 16'd64704, 16'd53456, 16'd53856});
	test_expansion(128'hd78cc70bbbada5d1a56df77055fa9106, {16'd20813, 16'd692, 16'd15269, 16'd49123, 16'd26301, 16'd29567, 16'd37551, 16'd17989, 16'd668, 16'd17866, 16'd12947, 16'd46784, 16'd35994, 16'd4981, 16'd13763, 16'd4737, 16'd43398, 16'd27344, 16'd18808, 16'd17685, 16'd42152, 16'd51247, 16'd50290, 16'd50566, 16'd57826, 16'd45793});
	test_expansion(128'h7ea44872adf85f48a93a72bd11de89f4, {16'd30498, 16'd45412, 16'd49413, 16'd22340, 16'd15335, 16'd25411, 16'd62455, 16'd55643, 16'd13845, 16'd43736, 16'd45008, 16'd36791, 16'd46438, 16'd7637, 16'd47649, 16'd43716, 16'd57957, 16'd31651, 16'd17931, 16'd33144, 16'd11422, 16'd37310, 16'd50285, 16'd59614, 16'd4584, 16'd9914});
	test_expansion(128'h6e32a04fe3725d0113ea3b9b62a83fcb, {16'd17455, 16'd59169, 16'd15983, 16'd30551, 16'd22846, 16'd30033, 16'd48918, 16'd55925, 16'd49058, 16'd32937, 16'd41870, 16'd41592, 16'd50605, 16'd22702, 16'd47484, 16'd43841, 16'd16913, 16'd6634, 16'd24823, 16'd31981, 16'd55785, 16'd16463, 16'd26060, 16'd43602, 16'd10879, 16'd17645});
	test_expansion(128'h1627a1a35835bd2a63b928baa3d89945, {16'd19431, 16'd41567, 16'd51828, 16'd60593, 16'd23677, 16'd30065, 16'd44029, 16'd31622, 16'd38469, 16'd42711, 16'd35342, 16'd6279, 16'd11212, 16'd35904, 16'd14368, 16'd42667, 16'd20816, 16'd33857, 16'd8306, 16'd1450, 16'd41035, 16'd44023, 16'd41326, 16'd14782, 16'd29741, 16'd6555});
	test_expansion(128'h07c7347db4733ae6da486af508733245, {16'd59403, 16'd62878, 16'd42191, 16'd28235, 16'd53357, 16'd10830, 16'd4032, 16'd8891, 16'd1329, 16'd16813, 16'd16984, 16'd28181, 16'd65037, 16'd18832, 16'd8528, 16'd14920, 16'd24634, 16'd61533, 16'd36895, 16'd17271, 16'd18593, 16'd15994, 16'd53372, 16'd30854, 16'd60714, 16'd27335});
	test_expansion(128'hf0d6d0330cac37da3c1635d37a8bbb4e, {16'd48829, 16'd20064, 16'd43564, 16'd13525, 16'd2051, 16'd59106, 16'd14818, 16'd5141, 16'd49974, 16'd17574, 16'd62637, 16'd15914, 16'd10594, 16'd61198, 16'd8095, 16'd38149, 16'd32868, 16'd10560, 16'd882, 16'd43480, 16'd39681, 16'd35924, 16'd3929, 16'd4071, 16'd42120, 16'd45528});
	test_expansion(128'ha5bfc77a75ac440adae9113c89eea787, {16'd31551, 16'd59397, 16'd59784, 16'd39769, 16'd46681, 16'd23082, 16'd16012, 16'd49558, 16'd30916, 16'd47847, 16'd59801, 16'd35573, 16'd61612, 16'd27510, 16'd62939, 16'd14956, 16'd8141, 16'd45073, 16'd9636, 16'd16426, 16'd52228, 16'd30882, 16'd59213, 16'd5585, 16'd16679, 16'd44307});
	test_expansion(128'h23868a75b75df4ea1d5179b04688e16d, {16'd38445, 16'd27943, 16'd4125, 16'd494, 16'd52775, 16'd41035, 16'd35170, 16'd31081, 16'd23223, 16'd16995, 16'd41043, 16'd10283, 16'd39301, 16'd30037, 16'd37449, 16'd12309, 16'd13067, 16'd62329, 16'd12659, 16'd63174, 16'd14920, 16'd56044, 16'd20358, 16'd5411, 16'd22965, 16'd26974});
	test_expansion(128'hf4e824bda260e8cb0ddd94235a535c01, {16'd39444, 16'd11658, 16'd18589, 16'd19780, 16'd64985, 16'd34596, 16'd44866, 16'd28840, 16'd43242, 16'd29767, 16'd13660, 16'd40329, 16'd2780, 16'd62325, 16'd63380, 16'd20885, 16'd25990, 16'd51274, 16'd50482, 16'd3815, 16'd27941, 16'd9066, 16'd38960, 16'd34283, 16'd33313, 16'd58441});
	test_expansion(128'hd59fd5643bce0f1052875ab01f7dde8f, {16'd25968, 16'd10471, 16'd56812, 16'd3703, 16'd16288, 16'd2370, 16'd16494, 16'd58513, 16'd60300, 16'd19035, 16'd31580, 16'd55623, 16'd19816, 16'd36937, 16'd35873, 16'd49310, 16'd56853, 16'd14559, 16'd18883, 16'd25773, 16'd38139, 16'd48400, 16'd6467, 16'd49744, 16'd52698, 16'd40457});
	test_expansion(128'h9f36dbb264a3c2751744bb0bce466191, {16'd57796, 16'd2908, 16'd17946, 16'd38965, 16'd61955, 16'd34818, 16'd33256, 16'd10636, 16'd27847, 16'd8531, 16'd4680, 16'd5489, 16'd30784, 16'd13850, 16'd56657, 16'd19802, 16'd49344, 16'd1818, 16'd65238, 16'd26356, 16'd25679, 16'd59651, 16'd60264, 16'd14948, 16'd56664, 16'd41264});
	test_expansion(128'he48ad2a5464cd4bad1976e29d18578f7, {16'd42367, 16'd56645, 16'd32200, 16'd55276, 16'd42502, 16'd35995, 16'd65304, 16'd64400, 16'd33134, 16'd16482, 16'd8350, 16'd37725, 16'd8061, 16'd13502, 16'd60737, 16'd17846, 16'd16689, 16'd55393, 16'd25489, 16'd16957, 16'd41635, 16'd7551, 16'd65202, 16'd9250, 16'd57938, 16'd34143});
	test_expansion(128'h54cf1f67889a5dc0f3cf2ee270d76e7e, {16'd16502, 16'd29012, 16'd23947, 16'd62052, 16'd21872, 16'd24860, 16'd16296, 16'd60595, 16'd6059, 16'd25887, 16'd28584, 16'd33988, 16'd64301, 16'd505, 16'd15217, 16'd718, 16'd16031, 16'd63726, 16'd39227, 16'd5657, 16'd29657, 16'd3360, 16'd582, 16'd1186, 16'd21895, 16'd64774});
	test_expansion(128'hab0f44bc4138a2ec7f1121a9b29aa3aa, {16'd51582, 16'd45936, 16'd50341, 16'd8102, 16'd46223, 16'd39753, 16'd55101, 16'd28926, 16'd33086, 16'd13446, 16'd36133, 16'd22694, 16'd42014, 16'd63095, 16'd47438, 16'd10311, 16'd14286, 16'd46104, 16'd34945, 16'd20193, 16'd19210, 16'd54753, 16'd8093, 16'd6360, 16'd8048, 16'd171});
	test_expansion(128'h3b184b8002104026a4cefda6b229d3a0, {16'd42721, 16'd43966, 16'd41818, 16'd63009, 16'd44859, 16'd62337, 16'd62623, 16'd51566, 16'd29211, 16'd29070, 16'd24566, 16'd64332, 16'd59952, 16'd6551, 16'd19414, 16'd13819, 16'd5471, 16'd25275, 16'd23285, 16'd60522, 16'd18578, 16'd13815, 16'd30067, 16'd17321, 16'd61165, 16'd63700});
	test_expansion(128'h6ca1e8e7f654ad444aa86f1c67d85601, {16'd32573, 16'd60279, 16'd28855, 16'd25093, 16'd49853, 16'd23706, 16'd20388, 16'd13006, 16'd56733, 16'd52139, 16'd15201, 16'd33286, 16'd48543, 16'd24199, 16'd21327, 16'd39749, 16'd44612, 16'd2700, 16'd50179, 16'd3757, 16'd21326, 16'd47056, 16'd22950, 16'd63530, 16'd60452, 16'd60868});
	test_expansion(128'hdc5586947b51ab9e600b6fc2c983f66d, {16'd47676, 16'd53481, 16'd36943, 16'd11124, 16'd5182, 16'd46480, 16'd52515, 16'd14841, 16'd25365, 16'd1376, 16'd43827, 16'd22025, 16'd31640, 16'd43792, 16'd24562, 16'd37477, 16'd27940, 16'd7161, 16'd7599, 16'd8699, 16'd54420, 16'd59449, 16'd25870, 16'd8443, 16'd18579, 16'd18343});
	test_expansion(128'h130951c8c8c1b4da7c9b0605e53f421c, {16'd6294, 16'd44384, 16'd54832, 16'd42499, 16'd14525, 16'd6929, 16'd19721, 16'd57596, 16'd39564, 16'd6992, 16'd13564, 16'd8396, 16'd11742, 16'd5074, 16'd31387, 16'd35487, 16'd9080, 16'd50666, 16'd18010, 16'd39749, 16'd61169, 16'd55722, 16'd33818, 16'd47376, 16'd28854, 16'd12412});
	test_expansion(128'h4a4b85d534c91183f6c051b79e6ca74d, {16'd2826, 16'd50620, 16'd47026, 16'd48129, 16'd62060, 16'd2463, 16'd64555, 16'd11785, 16'd45687, 16'd35574, 16'd40272, 16'd19755, 16'd30512, 16'd20801, 16'd26274, 16'd11016, 16'd5783, 16'd19347, 16'd1613, 16'd23495, 16'd19619, 16'd65240, 16'd17187, 16'd27899, 16'd31762, 16'd38887});
	test_expansion(128'h5e3d4f7378c0bffa93b93120c1fe0b10, {16'd40531, 16'd49188, 16'd39691, 16'd35446, 16'd23690, 16'd28077, 16'd63428, 16'd4121, 16'd14677, 16'd31464, 16'd26018, 16'd42453, 16'd47689, 16'd62108, 16'd49824, 16'd64192, 16'd53915, 16'd20736, 16'd23859, 16'd56184, 16'd17901, 16'd24409, 16'd12814, 16'd54835, 16'd23312, 16'd64239});
	test_expansion(128'h8c83c0df22ba257ebe725c189018a212, {16'd46549, 16'd15943, 16'd61350, 16'd55702, 16'd54598, 16'd22339, 16'd13416, 16'd47432, 16'd19125, 16'd33710, 16'd42132, 16'd26098, 16'd3524, 16'd34183, 16'd26613, 16'd46011, 16'd58722, 16'd20458, 16'd63462, 16'd4904, 16'd50389, 16'd33106, 16'd33263, 16'd21204, 16'd24976, 16'd57921});
	test_expansion(128'hc643331d87ea0a421b7542257db756e0, {16'd63746, 16'd9624, 16'd65455, 16'd51840, 16'd57638, 16'd52893, 16'd22900, 16'd25263, 16'd10828, 16'd19120, 16'd38543, 16'd7199, 16'd35178, 16'd1312, 16'd37588, 16'd23952, 16'd54402, 16'd19874, 16'd41056, 16'd1833, 16'd11456, 16'd15246, 16'd52778, 16'd17165, 16'd28664, 16'd27436});
	test_expansion(128'hd4c2b7d270abd7994fcc061a959f129d, {16'd53913, 16'd6844, 16'd45513, 16'd56931, 16'd8499, 16'd20060, 16'd60288, 16'd57055, 16'd13261, 16'd2156, 16'd49696, 16'd1746, 16'd32256, 16'd3073, 16'd15231, 16'd51036, 16'd38877, 16'd40004, 16'd30897, 16'd15959, 16'd16130, 16'd56832, 16'd56104, 16'd48749, 16'd56734, 16'd9804});
	test_expansion(128'hbc57c05d96ca7abc67e7cb7d3113ee3f, {16'd31289, 16'd43412, 16'd9474, 16'd34669, 16'd15049, 16'd7296, 16'd4572, 16'd21481, 16'd42287, 16'd6043, 16'd45742, 16'd999, 16'd51382, 16'd27608, 16'd34602, 16'd49691, 16'd23396, 16'd64198, 16'd32447, 16'd62479, 16'd45196, 16'd35531, 16'd58890, 16'd40366, 16'd9985, 16'd24865});
	test_expansion(128'h5492f441df9ed41ccd351ee32a465d5e, {16'd23908, 16'd3746, 16'd56697, 16'd49538, 16'd3184, 16'd6739, 16'd41322, 16'd5896, 16'd40743, 16'd51351, 16'd36654, 16'd57238, 16'd37075, 16'd61569, 16'd53755, 16'd2999, 16'd24119, 16'd24229, 16'd37689, 16'd45084, 16'd52052, 16'd40033, 16'd20335, 16'd52439, 16'd31845, 16'd44860});
	test_expansion(128'h0878b89e5036f5285b167a05d5dd00f7, {16'd27433, 16'd4596, 16'd26770, 16'd45763, 16'd18520, 16'd56626, 16'd57322, 16'd25768, 16'd20653, 16'd12370, 16'd24421, 16'd41199, 16'd29163, 16'd21060, 16'd24523, 16'd54708, 16'd7422, 16'd29290, 16'd42159, 16'd57470, 16'd33631, 16'd7305, 16'd26629, 16'd63094, 16'd38247, 16'd10854});
	test_expansion(128'h00a30174cc97d6fa60c2b69f9ba3ce2e, {16'd5420, 16'd8137, 16'd14489, 16'd44092, 16'd42711, 16'd16933, 16'd15748, 16'd32487, 16'd23569, 16'd2272, 16'd20974, 16'd46721, 16'd30283, 16'd33758, 16'd47499, 16'd29510, 16'd10480, 16'd34256, 16'd42467, 16'd53499, 16'd35332, 16'd52572, 16'd17260, 16'd28813, 16'd34812, 16'd38753});
	test_expansion(128'h850d1745412aa70735a671bfe9483d31, {16'd4118, 16'd46993, 16'd53986, 16'd19271, 16'd47160, 16'd59903, 16'd47276, 16'd52728, 16'd26338, 16'd44062, 16'd43901, 16'd44646, 16'd23259, 16'd34415, 16'd59950, 16'd34055, 16'd46171, 16'd39361, 16'd46732, 16'd57801, 16'd43643, 16'd36647, 16'd62548, 16'd49222, 16'd62400, 16'd22693});
	test_expansion(128'hcd428bc7698e5be58a4ba67d59e63e2d, {16'd12661, 16'd8797, 16'd9876, 16'd24562, 16'd35150, 16'd38340, 16'd39664, 16'd44703, 16'd39640, 16'd17138, 16'd8640, 16'd64862, 16'd42822, 16'd54171, 16'd46572, 16'd49206, 16'd38687, 16'd54769, 16'd11368, 16'd60911, 16'd59712, 16'd12574, 16'd4460, 16'd54672, 16'd15988, 16'd65125});
	test_expansion(128'h2b8ad6c801f93cf596d53a200ecd0a5c, {16'd50160, 16'd2391, 16'd41225, 16'd65059, 16'd7572, 16'd44621, 16'd19754, 16'd62442, 16'd16957, 16'd64925, 16'd5532, 16'd18067, 16'd38777, 16'd50715, 16'd26544, 16'd2311, 16'd24579, 16'd46076, 16'd18216, 16'd52437, 16'd34807, 16'd36955, 16'd7625, 16'd62936, 16'd47921, 16'd3323});
	test_expansion(128'hdbbd2b59c2750ee342f18352270f24f6, {16'd218, 16'd58655, 16'd15947, 16'd60993, 16'd34700, 16'd34363, 16'd57839, 16'd48647, 16'd64319, 16'd23770, 16'd64035, 16'd27076, 16'd52779, 16'd52712, 16'd32334, 16'd64985, 16'd49629, 16'd15537, 16'd42654, 16'd19236, 16'd18892, 16'd15498, 16'd45670, 16'd59726, 16'd43711, 16'd55197});
	test_expansion(128'hd38aacca926cea0196cbce47b8eab88e, {16'd38965, 16'd13193, 16'd63266, 16'd58148, 16'd45133, 16'd38828, 16'd7498, 16'd7966, 16'd11246, 16'd9683, 16'd13480, 16'd53216, 16'd35973, 16'd34454, 16'd46939, 16'd22640, 16'd32259, 16'd49321, 16'd50759, 16'd50697, 16'd8807, 16'd59182, 16'd30239, 16'd59490, 16'd37660, 16'd14906});
	test_expansion(128'h22a9beb614d1ebae480d1d82544f9fd1, {16'd39997, 16'd61810, 16'd15072, 16'd50273, 16'd45163, 16'd4273, 16'd31666, 16'd31740, 16'd11871, 16'd3336, 16'd1187, 16'd30450, 16'd20916, 16'd53935, 16'd63016, 16'd43373, 16'd33913, 16'd56515, 16'd42583, 16'd5700, 16'd48699, 16'd63947, 16'd9027, 16'd59322, 16'd9947, 16'd19626});
	test_expansion(128'h13c3a62a276cf73dce2b6980f03eac71, {16'd38231, 16'd36770, 16'd57553, 16'd2870, 16'd30102, 16'd23690, 16'd4608, 16'd23935, 16'd48308, 16'd59355, 16'd45004, 16'd60287, 16'd38667, 16'd5974, 16'd23142, 16'd12555, 16'd57806, 16'd41010, 16'd52636, 16'd60251, 16'd21947, 16'd55232, 16'd6411, 16'd1648, 16'd56881, 16'd44454});
	test_expansion(128'h0a790f154542f4950c5209b5c0f054c8, {16'd22374, 16'd36514, 16'd53101, 16'd17278, 16'd9888, 16'd7799, 16'd46487, 16'd57461, 16'd19290, 16'd7281, 16'd12760, 16'd37987, 16'd2720, 16'd25895, 16'd6382, 16'd49615, 16'd45245, 16'd39532, 16'd65299, 16'd17385, 16'd58340, 16'd19695, 16'd65489, 16'd10909, 16'd27543, 16'd18127});
	test_expansion(128'ha0f3c5650a18a94bf7353b77c3beedd7, {16'd44688, 16'd5391, 16'd60407, 16'd16356, 16'd44203, 16'd43285, 16'd30325, 16'd15628, 16'd32700, 16'd38787, 16'd16351, 16'd32650, 16'd35341, 16'd27137, 16'd7877, 16'd10023, 16'd1721, 16'd6005, 16'd64542, 16'd550, 16'd65199, 16'd63339, 16'd24623, 16'd13385, 16'd52360, 16'd25772});
	test_expansion(128'hb8fcc4406f2d37c3e85b4b9dea24f375, {16'd37300, 16'd34296, 16'd16708, 16'd40904, 16'd52334, 16'd25791, 16'd58811, 16'd13886, 16'd14108, 16'd49555, 16'd65237, 16'd27857, 16'd63069, 16'd4753, 16'd63396, 16'd56125, 16'd61479, 16'd56619, 16'd16579, 16'd42853, 16'd55916, 16'd37035, 16'd58870, 16'd27212, 16'd42001, 16'd60311});
	test_expansion(128'hdeecb756d7fcf6d028647fe3cbbfc097, {16'd55397, 16'd20222, 16'd1071, 16'd6351, 16'd62599, 16'd40331, 16'd10290, 16'd23499, 16'd27055, 16'd56302, 16'd22104, 16'd21660, 16'd10119, 16'd8782, 16'd54419, 16'd18083, 16'd55208, 16'd33623, 16'd16109, 16'd61811, 16'd4932, 16'd56775, 16'd21155, 16'd39368, 16'd25858, 16'd11432});
	test_expansion(128'h8d916ccbef5a331fcc746aedfb83af9a, {16'd63254, 16'd22033, 16'd48610, 16'd43806, 16'd10662, 16'd46814, 16'd26483, 16'd26084, 16'd56000, 16'd30754, 16'd8037, 16'd41827, 16'd32990, 16'd16442, 16'd17260, 16'd39829, 16'd13084, 16'd62621, 16'd25008, 16'd35459, 16'd49993, 16'd33942, 16'd18225, 16'd41105, 16'd1090, 16'd38896});
	test_expansion(128'h45aaff42a364f39988d7cef8e2e0248f, {16'd10733, 16'd32260, 16'd41876, 16'd10883, 16'd30974, 16'd57686, 16'd24041, 16'd7845, 16'd23661, 16'd32058, 16'd30382, 16'd17362, 16'd16826, 16'd38888, 16'd28482, 16'd43318, 16'd38478, 16'd20902, 16'd51902, 16'd54736, 16'd49749, 16'd44045, 16'd31473, 16'd35876, 16'd31533, 16'd496});
	test_expansion(128'hd1831c8107598af6f10acce9652ade54, {16'd48577, 16'd35348, 16'd18096, 16'd4838, 16'd1413, 16'd57312, 16'd5980, 16'd28716, 16'd30036, 16'd10255, 16'd54379, 16'd31036, 16'd22451, 16'd16406, 16'd43329, 16'd27840, 16'd19260, 16'd52239, 16'd24132, 16'd63896, 16'd28852, 16'd12017, 16'd38440, 16'd16494, 16'd16253, 16'd43648});
	test_expansion(128'h3dc85f85f244c4df0b561f1b80261e1b, {16'd38307, 16'd34346, 16'd45487, 16'd28172, 16'd1928, 16'd56612, 16'd39211, 16'd52990, 16'd58094, 16'd13149, 16'd19051, 16'd37429, 16'd16315, 16'd7284, 16'd8304, 16'd64253, 16'd45258, 16'd55928, 16'd63033, 16'd41308, 16'd18275, 16'd58718, 16'd20148, 16'd29470, 16'd22003, 16'd39085});
	test_expansion(128'hd39a7da59ff125087b90a5dacd1d1d45, {16'd2951, 16'd9802, 16'd10998, 16'd23893, 16'd22655, 16'd36748, 16'd1473, 16'd60599, 16'd18444, 16'd19650, 16'd62552, 16'd3328, 16'd47853, 16'd3002, 16'd40423, 16'd48236, 16'd10353, 16'd59192, 16'd4107, 16'd11287, 16'd21206, 16'd28539, 16'd12435, 16'd16726, 16'd10891, 16'd62003});
	test_expansion(128'he83ce641fc0ed115a338a9e29e6e3d53, {16'd52272, 16'd3288, 16'd54612, 16'd4713, 16'd40047, 16'd45069, 16'd52807, 16'd36832, 16'd46208, 16'd22962, 16'd26779, 16'd30867, 16'd6495, 16'd18216, 16'd46753, 16'd42938, 16'd3654, 16'd18223, 16'd50037, 16'd31982, 16'd53874, 16'd40622, 16'd33726, 16'd17783, 16'd20327, 16'd27039});
	test_expansion(128'h649c727503f23a5ed92b315d5a55d678, {16'd30968, 16'd4127, 16'd41597, 16'd43781, 16'd61943, 16'd21883, 16'd52903, 16'd37638, 16'd57306, 16'd44485, 16'd57677, 16'd61820, 16'd1347, 16'd45311, 16'd37519, 16'd55753, 16'd3334, 16'd10797, 16'd55712, 16'd29381, 16'd56920, 16'd20482, 16'd52066, 16'd50785, 16'd43723, 16'd55169});
	test_expansion(128'h95a822e17763d6f36145871bdd6b6fb6, {16'd16720, 16'd57600, 16'd40902, 16'd42259, 16'd13318, 16'd10683, 16'd56477, 16'd56897, 16'd9304, 16'd17805, 16'd29884, 16'd39403, 16'd32788, 16'd30815, 16'd22335, 16'd17405, 16'd15417, 16'd62836, 16'd28835, 16'd8403, 16'd20014, 16'd51016, 16'd11901, 16'd13226, 16'd33304, 16'd40414});
	test_expansion(128'h3837a0a6d35d3b0dc878c7e15a568fa4, {16'd45612, 16'd15267, 16'd48737, 16'd63701, 16'd45899, 16'd22405, 16'd1882, 16'd46263, 16'd62173, 16'd21124, 16'd33708, 16'd49547, 16'd50733, 16'd25405, 16'd45517, 16'd10490, 16'd35414, 16'd41209, 16'd39155, 16'd52585, 16'd42556, 16'd9959, 16'd1207, 16'd26869, 16'd51909, 16'd35413});
	test_expansion(128'h1efdd6bc8b9fa60454b7f0c5afbdf9b6, {16'd7583, 16'd41178, 16'd29074, 16'd53980, 16'd30713, 16'd56422, 16'd64499, 16'd64839, 16'd33809, 16'd53454, 16'd11586, 16'd3685, 16'd674, 16'd27701, 16'd26050, 16'd58912, 16'd9342, 16'd27141, 16'd54188, 16'd52764, 16'd18058, 16'd39653, 16'd27561, 16'd17081, 16'd29371, 16'd64213});
	test_expansion(128'h887dcbdc32c66d2e36bc29c67f817578, {16'd27394, 16'd12282, 16'd56368, 16'd25580, 16'd54887, 16'd64936, 16'd34593, 16'd30597, 16'd2676, 16'd39473, 16'd52557, 16'd24123, 16'd4776, 16'd59150, 16'd29781, 16'd52537, 16'd40114, 16'd38157, 16'd51613, 16'd23173, 16'd23151, 16'd6074, 16'd56698, 16'd43221, 16'd38535, 16'd20479});
	test_expansion(128'hc120e3b4bf8fbf2f1af7bd9244e2016b, {16'd41240, 16'd13296, 16'd43071, 16'd10331, 16'd58145, 16'd39060, 16'd46648, 16'd29464, 16'd60321, 16'd45141, 16'd33341, 16'd5016, 16'd31594, 16'd42302, 16'd24876, 16'd43024, 16'd56471, 16'd60435, 16'd39926, 16'd28145, 16'd24262, 16'd12987, 16'd23656, 16'd65090, 16'd21163, 16'd57584});
	test_expansion(128'hf43f3cb840c2b346fcf1152e9539c484, {16'd3768, 16'd40522, 16'd10888, 16'd52791, 16'd9022, 16'd34511, 16'd63597, 16'd41196, 16'd52715, 16'd4712, 16'd46976, 16'd15859, 16'd8082, 16'd58251, 16'd12377, 16'd43207, 16'd10246, 16'd47071, 16'd23531, 16'd49313, 16'd27612, 16'd35557, 16'd54596, 16'd4801, 16'd63056, 16'd2789});
	test_expansion(128'hdf35c8715e268dc218d57c9403ac27b5, {16'd16777, 16'd62290, 16'd40920, 16'd14535, 16'd62612, 16'd44649, 16'd36742, 16'd27064, 16'd29592, 16'd46323, 16'd5741, 16'd56098, 16'd25807, 16'd29298, 16'd8424, 16'd51031, 16'd42095, 16'd64417, 16'd2855, 16'd7393, 16'd44832, 16'd38196, 16'd8140, 16'd28390, 16'd31882, 16'd53147});
	test_expansion(128'h52b0f608098217d2a6dadfeb6e49e830, {16'd12812, 16'd30741, 16'd29456, 16'd23523, 16'd35191, 16'd2011, 16'd39903, 16'd25377, 16'd48952, 16'd62681, 16'd20297, 16'd7844, 16'd58968, 16'd10042, 16'd32818, 16'd54135, 16'd26613, 16'd39796, 16'd42298, 16'd8083, 16'd50278, 16'd41964, 16'd59303, 16'd44805, 16'd12249, 16'd26411});
	test_expansion(128'ha29449cc8e5c32f820e02ac2e2998a13, {16'd52992, 16'd20031, 16'd49003, 16'd21469, 16'd53929, 16'd1154, 16'd46654, 16'd36546, 16'd62762, 16'd24252, 16'd48757, 16'd9632, 16'd56533, 16'd37793, 16'd30679, 16'd9789, 16'd62430, 16'd19875, 16'd33792, 16'd42545, 16'd50299, 16'd6578, 16'd49563, 16'd17984, 16'd4559, 16'd4105});
	test_expansion(128'hc466b74642c9a693c30a1ae49a63a613, {16'd30027, 16'd41549, 16'd27552, 16'd64167, 16'd60908, 16'd50093, 16'd13869, 16'd8908, 16'd17112, 16'd33098, 16'd55749, 16'd64760, 16'd28730, 16'd28677, 16'd8654, 16'd47368, 16'd44010, 16'd31819, 16'd6318, 16'd64559, 16'd5208, 16'd23178, 16'd63091, 16'd12256, 16'd48328, 16'd58484});
	test_expansion(128'h5fed8d167945c166cbb251a396d4f240, {16'd16206, 16'd22310, 16'd64633, 16'd45439, 16'd42529, 16'd65512, 16'd11646, 16'd63163, 16'd46927, 16'd52166, 16'd63813, 16'd11330, 16'd55360, 16'd51439, 16'd24523, 16'd57004, 16'd4806, 16'd64719, 16'd53345, 16'd30493, 16'd47205, 16'd50757, 16'd38520, 16'd63900, 16'd27592, 16'd19917});
	test_expansion(128'h02fc7da497ae0ddc5670065ced2d529d, {16'd59058, 16'd22688, 16'd10785, 16'd3124, 16'd7827, 16'd30171, 16'd27672, 16'd60185, 16'd57111, 16'd16074, 16'd16091, 16'd9691, 16'd35122, 16'd31390, 16'd4771, 16'd5748, 16'd26740, 16'd2473, 16'd61420, 16'd64320, 16'd5221, 16'd22399, 16'd41234, 16'd38520, 16'd28707, 16'd29765});
	test_expansion(128'hbc2709c1d00d23f562ec9592a1ede535, {16'd20850, 16'd45442, 16'd9886, 16'd783, 16'd35708, 16'd2243, 16'd25944, 16'd63985, 16'd48473, 16'd47111, 16'd5991, 16'd52960, 16'd48791, 16'd1550, 16'd50866, 16'd17374, 16'd14133, 16'd19408, 16'd60764, 16'd62289, 16'd43448, 16'd2442, 16'd26817, 16'd36466, 16'd9970, 16'd46750});
	test_expansion(128'h4dcfbb34acc2368ca2b7363da4ffc7e8, {16'd60590, 16'd47127, 16'd12669, 16'd35059, 16'd65115, 16'd8572, 16'd49818, 16'd6607, 16'd46933, 16'd5260, 16'd18571, 16'd54394, 16'd17816, 16'd52902, 16'd53112, 16'd47770, 16'd16055, 16'd1523, 16'd8606, 16'd33968, 16'd21945, 16'd38439, 16'd200, 16'd59208, 16'd38555, 16'd50594});
	test_expansion(128'h478ddaf3d40f5eabdc4d4b51f6f0120d, {16'd51883, 16'd17826, 16'd12387, 16'd48553, 16'd54827, 16'd23992, 16'd25039, 16'd31231, 16'd1943, 16'd50720, 16'd61461, 16'd16533, 16'd14091, 16'd17719, 16'd14949, 16'd16708, 16'd51266, 16'd23669, 16'd13436, 16'd13300, 16'd32943, 16'd49903, 16'd5805, 16'd43071, 16'd60106, 16'd61013});
	test_expansion(128'hd2ac64e8430b2fa9bf88f60c2569de80, {16'd32523, 16'd3684, 16'd16001, 16'd51177, 16'd62454, 16'd48761, 16'd7950, 16'd37447, 16'd30540, 16'd17800, 16'd43563, 16'd57430, 16'd51344, 16'd35275, 16'd5929, 16'd10592, 16'd55678, 16'd21600, 16'd58063, 16'd55162, 16'd57278, 16'd4756, 16'd64020, 16'd49546, 16'd37323, 16'd26981});
	test_expansion(128'h45f7b85925aaaf3aea08704be0bebea6, {16'd11641, 16'd28902, 16'd15184, 16'd26616, 16'd54325, 16'd7307, 16'd61084, 16'd31053, 16'd19063, 16'd50217, 16'd12892, 16'd43446, 16'd57282, 16'd55041, 16'd24702, 16'd9759, 16'd8828, 16'd14742, 16'd40233, 16'd52318, 16'd11514, 16'd815, 16'd51437, 16'd1669, 16'd17283, 16'd64335});
	test_expansion(128'h36dee80fb2bf8f9d58e5ec1465c108b8, {16'd21113, 16'd5319, 16'd31718, 16'd62686, 16'd30142, 16'd21858, 16'd12537, 16'd29691, 16'd34128, 16'd55110, 16'd43134, 16'd36442, 16'd51682, 16'd22604, 16'd27476, 16'd51227, 16'd6767, 16'd51847, 16'd11097, 16'd63731, 16'd13510, 16'd65508, 16'd54170, 16'd912, 16'd31442, 16'd54345});
	test_expansion(128'h95b2f8b7958e702869e8ad6091e7555c, {16'd55372, 16'd64244, 16'd50930, 16'd26409, 16'd42984, 16'd53062, 16'd10044, 16'd36419, 16'd35275, 16'd39064, 16'd38858, 16'd23645, 16'd25104, 16'd14274, 16'd21924, 16'd21092, 16'd3298, 16'd57504, 16'd52274, 16'd3952, 16'd21710, 16'd46877, 16'd45559, 16'd30007, 16'd30175, 16'd63577});
	test_expansion(128'h101ef3c574fe9f616b0a246c452cd732, {16'd18571, 16'd55289, 16'd12875, 16'd20616, 16'd41597, 16'd64718, 16'd49907, 16'd33612, 16'd1033, 16'd25538, 16'd37476, 16'd44755, 16'd23994, 16'd31489, 16'd24810, 16'd11805, 16'd56301, 16'd44041, 16'd40548, 16'd35377, 16'd27088, 16'd19298, 16'd63668, 16'd42327, 16'd4528, 16'd49373});
	test_expansion(128'hf0b3fc7473eb875391c5279b2c3a7872, {16'd47196, 16'd37382, 16'd58166, 16'd19233, 16'd35404, 16'd39778, 16'd34791, 16'd61851, 16'd21235, 16'd36776, 16'd45485, 16'd20213, 16'd55945, 16'd1302, 16'd45615, 16'd17425, 16'd30465, 16'd54303, 16'd45361, 16'd49577, 16'd31779, 16'd54106, 16'd18183, 16'd36783, 16'd27922, 16'd17949});
	test_expansion(128'hf2d18af6fb4462d69b97f9a7f43caa16, {16'd30427, 16'd15301, 16'd1072, 16'd26305, 16'd36073, 16'd64408, 16'd43760, 16'd52727, 16'd63115, 16'd31820, 16'd17394, 16'd6026, 16'd35820, 16'd20498, 16'd28883, 16'd2957, 16'd25543, 16'd49772, 16'd16473, 16'd29627, 16'd60571, 16'd44098, 16'd59137, 16'd21997, 16'd49822, 16'd28080});
	test_expansion(128'hbfb72916c91314747a346964cda34dd4, {16'd22318, 16'd21215, 16'd53299, 16'd10489, 16'd53058, 16'd19924, 16'd36278, 16'd37137, 16'd45154, 16'd49257, 16'd64749, 16'd39943, 16'd28942, 16'd33756, 16'd23751, 16'd63598, 16'd15368, 16'd2261, 16'd14703, 16'd34723, 16'd60834, 16'd38162, 16'd44544, 16'd46201, 16'd63627, 16'd52913});
	test_expansion(128'hd6588c962fb965db765dc6ee0b31c347, {16'd61613, 16'd45392, 16'd55080, 16'd59357, 16'd11545, 16'd57207, 16'd37085, 16'd22472, 16'd52388, 16'd39386, 16'd12190, 16'd48235, 16'd11216, 16'd32765, 16'd20706, 16'd22933, 16'd57954, 16'd23816, 16'd65104, 16'd14038, 16'd61988, 16'd48245, 16'd63440, 16'd32795, 16'd61162, 16'd59812});
	test_expansion(128'hedeff5df84c92d3cdc01821790ee89d3, {16'd14582, 16'd47307, 16'd61357, 16'd16508, 16'd27160, 16'd37881, 16'd26199, 16'd15564, 16'd28990, 16'd28889, 16'd57449, 16'd46247, 16'd59414, 16'd29283, 16'd38737, 16'd43095, 16'd9222, 16'd56520, 16'd30141, 16'd54863, 16'd33612, 16'd47234, 16'd47466, 16'd27133, 16'd38663, 16'd2103});
	test_expansion(128'h4965b0dc19bb9601525281fe39881845, {16'd64838, 16'd41035, 16'd42715, 16'd13119, 16'd5066, 16'd1257, 16'd13248, 16'd4997, 16'd36751, 16'd30406, 16'd44162, 16'd40885, 16'd15718, 16'd26580, 16'd27699, 16'd10247, 16'd46620, 16'd60497, 16'd48003, 16'd38337, 16'd53172, 16'd38374, 16'd64249, 16'd6482, 16'd35318, 16'd7616});
	test_expansion(128'hd875072e518cec6351be87320d3b18e1, {16'd18288, 16'd41593, 16'd35931, 16'd41538, 16'd46894, 16'd53921, 16'd63662, 16'd45633, 16'd43523, 16'd47620, 16'd17228, 16'd51716, 16'd22519, 16'd60131, 16'd32214, 16'd49260, 16'd13009, 16'd28858, 16'd16416, 16'd50875, 16'd3300, 16'd33603, 16'd36829, 16'd4558, 16'd32424, 16'd56491});
	test_expansion(128'h07da6a2e1f89da3d38e8f9803dfd0beb, {16'd53071, 16'd39807, 16'd35604, 16'd33766, 16'd35322, 16'd22731, 16'd18073, 16'd21902, 16'd47446, 16'd36652, 16'd6948, 16'd22545, 16'd42131, 16'd3232, 16'd13613, 16'd37256, 16'd48444, 16'd61740, 16'd1697, 16'd50744, 16'd3062, 16'd43742, 16'd3145, 16'd42651, 16'd29927, 16'd12022});
	test_expansion(128'h07343b60750d3f40069e2db0c3e1e4d3, {16'd49120, 16'd54058, 16'd63401, 16'd10453, 16'd63537, 16'd1259, 16'd60220, 16'd33195, 16'd42999, 16'd45368, 16'd37697, 16'd40401, 16'd16875, 16'd50676, 16'd40783, 16'd22550, 16'd15962, 16'd5772, 16'd5941, 16'd7999, 16'd46077, 16'd15455, 16'd60600, 16'd61645, 16'd58054, 16'd13119});
	test_expansion(128'hc9741338b086bbea94b2f9e07b2fdfd9, {16'd24497, 16'd60362, 16'd59578, 16'd61923, 16'd50999, 16'd10194, 16'd18429, 16'd14831, 16'd43458, 16'd61668, 16'd3041, 16'd44867, 16'd43254, 16'd51427, 16'd18752, 16'd3722, 16'd34868, 16'd14121, 16'd55141, 16'd34791, 16'd60844, 16'd1492, 16'd28430, 16'd43999, 16'd45306, 16'd15122});
	test_expansion(128'h6cbb5a56f72cd27eeccac8103c3855c8, {16'd52852, 16'd45957, 16'd17593, 16'd3614, 16'd14896, 16'd62212, 16'd62485, 16'd19048, 16'd49576, 16'd63925, 16'd63028, 16'd46351, 16'd4357, 16'd8497, 16'd33954, 16'd4537, 16'd15327, 16'd62115, 16'd11955, 16'd62735, 16'd55026, 16'd21935, 16'd32419, 16'd49045, 16'd42422, 16'd49192});
	test_expansion(128'h7e31d0e2523490153d04eeb23a79603d, {16'd17692, 16'd44186, 16'd32275, 16'd41781, 16'd48250, 16'd21154, 16'd29734, 16'd48094, 16'd1915, 16'd43378, 16'd51334, 16'd53794, 16'd18317, 16'd5343, 16'd29082, 16'd62922, 16'd27505, 16'd62843, 16'd42724, 16'd18386, 16'd26737, 16'd34486, 16'd31427, 16'd9331, 16'd13300, 16'd17283});
	test_expansion(128'h266f6534ca6928466254abb7df73f6f1, {16'd7511, 16'd58268, 16'd5187, 16'd57735, 16'd33690, 16'd773, 16'd62375, 16'd56340, 16'd24715, 16'd65034, 16'd9126, 16'd49591, 16'd2575, 16'd45968, 16'd54409, 16'd46008, 16'd7268, 16'd5291, 16'd53250, 16'd3928, 16'd57359, 16'd62044, 16'd32012, 16'd60929, 16'd56108, 16'd59241});
	test_expansion(128'ha02ee9033b9b2a748152df8bbae63f99, {16'd6489, 16'd27187, 16'd33510, 16'd59319, 16'd29828, 16'd62849, 16'd20706, 16'd52484, 16'd2602, 16'd57675, 16'd8062, 16'd37670, 16'd28972, 16'd63875, 16'd1686, 16'd10322, 16'd848, 16'd8278, 16'd40361, 16'd41440, 16'd3425, 16'd31019, 16'd20758, 16'd11326, 16'd50058, 16'd36769});
	test_expansion(128'h19ee78e8bca28d641877dce3bae5722f, {16'd41211, 16'd47816, 16'd38722, 16'd52177, 16'd62594, 16'd42957, 16'd27249, 16'd20825, 16'd63648, 16'd30753, 16'd13819, 16'd44795, 16'd19880, 16'd1145, 16'd25979, 16'd57679, 16'd44561, 16'd36539, 16'd21365, 16'd44030, 16'd60400, 16'd1424, 16'd40156, 16'd14002, 16'd33076, 16'd23103});
	test_expansion(128'hd26dd2ffc9eb2bc163a28112b60569b2, {16'd30842, 16'd35157, 16'd3519, 16'd26893, 16'd62631, 16'd59230, 16'd27021, 16'd17386, 16'd6223, 16'd20582, 16'd62113, 16'd25310, 16'd61033, 16'd28393, 16'd55180, 16'd16628, 16'd21153, 16'd13887, 16'd23553, 16'd9176, 16'd49143, 16'd30401, 16'd47065, 16'd18732, 16'd39406, 16'd45811});
	test_expansion(128'hbdfab7acfc127312141440c7356c098f, {16'd586, 16'd63495, 16'd53733, 16'd28533, 16'd17596, 16'd31938, 16'd45666, 16'd9836, 16'd24238, 16'd30670, 16'd13556, 16'd26031, 16'd10081, 16'd42659, 16'd56847, 16'd6492, 16'd49072, 16'd25439, 16'd31765, 16'd13312, 16'd31217, 16'd8266, 16'd23571, 16'd59869, 16'd45119, 16'd20920});
	test_expansion(128'hf52639d154fea5c53f58b89ef5d878ee, {16'd64406, 16'd12682, 16'd39667, 16'd46727, 16'd64409, 16'd47410, 16'd36060, 16'd41683, 16'd30695, 16'd46097, 16'd2233, 16'd57015, 16'd37440, 16'd28668, 16'd43501, 16'd42408, 16'd3001, 16'd52848, 16'd32817, 16'd27290, 16'd14962, 16'd39047, 16'd11419, 16'd28258, 16'd50633, 16'd54506});
	test_expansion(128'h230d23c20195ff94e6d33f109c8b44a9, {16'd5397, 16'd12174, 16'd10751, 16'd62890, 16'd6180, 16'd9821, 16'd52397, 16'd8332, 16'd64813, 16'd60071, 16'd63412, 16'd40113, 16'd35028, 16'd21696, 16'd12030, 16'd11969, 16'd51503, 16'd56807, 16'd24267, 16'd17574, 16'd49072, 16'd26697, 16'd17717, 16'd10617, 16'd5022, 16'd51373});
	test_expansion(128'h7fbe1112013343895fb548c3897bf78c, {16'd47171, 16'd7506, 16'd24189, 16'd62698, 16'd29855, 16'd6673, 16'd56311, 16'd12790, 16'd58440, 16'd51083, 16'd30580, 16'd21885, 16'd16979, 16'd49231, 16'd12827, 16'd55089, 16'd1846, 16'd41844, 16'd52430, 16'd54557, 16'd38034, 16'd21647, 16'd44062, 16'd20408, 16'd42224, 16'd53931});
	test_expansion(128'ha99f5fff8854678da051de8cfadabd83, {16'd52327, 16'd55229, 16'd41379, 16'd18515, 16'd65392, 16'd19221, 16'd27814, 16'd13768, 16'd31452, 16'd23869, 16'd50421, 16'd39519, 16'd24764, 16'd5351, 16'd38940, 16'd57730, 16'd25449, 16'd7808, 16'd36544, 16'd63742, 16'd38659, 16'd44051, 16'd8506, 16'd47429, 16'd51302, 16'd26707});
	test_expansion(128'hb94a771a45c439b0958efd52f22501fd, {16'd41989, 16'd58637, 16'd38581, 16'd57432, 16'd3785, 16'd29703, 16'd15155, 16'd54709, 16'd26900, 16'd58606, 16'd62523, 16'd10345, 16'd33203, 16'd60731, 16'd7854, 16'd43445, 16'd13566, 16'd27835, 16'd58126, 16'd65085, 16'd52315, 16'd44172, 16'd36932, 16'd63516, 16'd29041, 16'd32772});
	test_expansion(128'h3d57eebe34554c202a602305c5b73fd1, {16'd11462, 16'd1134, 16'd22153, 16'd52139, 16'd2499, 16'd45268, 16'd51148, 16'd27332, 16'd46016, 16'd45515, 16'd45650, 16'd48859, 16'd54727, 16'd21307, 16'd24638, 16'd62011, 16'd53399, 16'd40792, 16'd35149, 16'd40065, 16'd52853, 16'd59065, 16'd11250, 16'd12567, 16'd43172, 16'd35065});
	test_expansion(128'h9763f0bdd01c6ade68ffe6ab99637d41, {16'd35527, 16'd48439, 16'd11032, 16'd65112, 16'd39632, 16'd25822, 16'd11805, 16'd11838, 16'd33787, 16'd63704, 16'd36716, 16'd60855, 16'd63776, 16'd2507, 16'd54571, 16'd58067, 16'd32371, 16'd22695, 16'd32473, 16'd12311, 16'd30391, 16'd9797, 16'd30943, 16'd22879, 16'd23360, 16'd39619});
	test_expansion(128'h0978ea9512abbb6f559aded769d8e663, {16'd9732, 16'd14647, 16'd56179, 16'd13044, 16'd15271, 16'd28776, 16'd7741, 16'd2797, 16'd59736, 16'd31252, 16'd60368, 16'd9120, 16'd22680, 16'd32033, 16'd40000, 16'd65067, 16'd19973, 16'd1620, 16'd29058, 16'd11618, 16'd45371, 16'd31877, 16'd6575, 16'd46582, 16'd42157, 16'd49172});
	test_expansion(128'h0bfedd370d51cc530f8c96efea3a4ef9, {16'd41730, 16'd32536, 16'd11161, 16'd5432, 16'd17468, 16'd63315, 16'd8105, 16'd4060, 16'd26533, 16'd55834, 16'd43547, 16'd62115, 16'd31661, 16'd48046, 16'd58739, 16'd27237, 16'd281, 16'd44969, 16'd22674, 16'd39345, 16'd54488, 16'd45985, 16'd60982, 16'd7640, 16'd16001, 16'd1874});
	test_expansion(128'h5ada18c77e6848022545a080b36ecf94, {16'd4008, 16'd22841, 16'd63635, 16'd58303, 16'd55045, 16'd39766, 16'd62937, 16'd51327, 16'd39345, 16'd26444, 16'd23045, 16'd50847, 16'd40865, 16'd59158, 16'd2054, 16'd33963, 16'd2521, 16'd49419, 16'd46881, 16'd31574, 16'd9789, 16'd59791, 16'd46711, 16'd14137, 16'd62057, 16'd9727});
	test_expansion(128'h7137712abde5ba3954a395d8f8955a4b, {16'd31726, 16'd12877, 16'd27853, 16'd56597, 16'd63378, 16'd57535, 16'd14957, 16'd17849, 16'd38717, 16'd3106, 16'd30465, 16'd57223, 16'd43071, 16'd54148, 16'd37466, 16'd62036, 16'd63551, 16'd2171, 16'd52041, 16'd22048, 16'd51235, 16'd15638, 16'd45982, 16'd50593, 16'd42263, 16'd41532});
	test_expansion(128'h7d403f56622825e05a712d61a696347f, {16'd40983, 16'd64608, 16'd33409, 16'd51981, 16'd26619, 16'd48463, 16'd18674, 16'd32243, 16'd52994, 16'd49488, 16'd24313, 16'd55601, 16'd2195, 16'd16905, 16'd26625, 16'd59369, 16'd31600, 16'd34688, 16'd33376, 16'd30878, 16'd8834, 16'd28189, 16'd60832, 16'd47267, 16'd45459, 16'd8756});
	test_expansion(128'h33afdf6481b1abfd3d226aa4107459e4, {16'd57006, 16'd14980, 16'd33170, 16'd51470, 16'd52323, 16'd10574, 16'd3405, 16'd32229, 16'd10571, 16'd48782, 16'd35262, 16'd43194, 16'd51507, 16'd57310, 16'd57014, 16'd53989, 16'd19709, 16'd44793, 16'd3606, 16'd38837, 16'd42516, 16'd64966, 16'd57788, 16'd9726, 16'd32674, 16'd13258});
	test_expansion(128'h51f3011141a7377671b813634f425896, {16'd34982, 16'd27130, 16'd4475, 16'd36365, 16'd35228, 16'd25465, 16'd25290, 16'd64626, 16'd34990, 16'd49803, 16'd14750, 16'd40383, 16'd3250, 16'd60179, 16'd54144, 16'd14615, 16'd3733, 16'd9158, 16'd15228, 16'd9222, 16'd8884, 16'd12493, 16'd48834, 16'd48137, 16'd47153, 16'd41678});
	test_expansion(128'h0eae47d30ecf0ecb239bf66884d0033a, {16'd61504, 16'd48467, 16'd7756, 16'd13852, 16'd2378, 16'd29680, 16'd62868, 16'd11122, 16'd9180, 16'd56253, 16'd59488, 16'd4891, 16'd54180, 16'd56944, 16'd37360, 16'd47423, 16'd45936, 16'd55689, 16'd55049, 16'd43017, 16'd46360, 16'd19902, 16'd38329, 16'd12196, 16'd41060, 16'd55087});
	test_expansion(128'h792c7d34f262ca3ee3a905f4314051ed, {16'd37859, 16'd12484, 16'd34576, 16'd14941, 16'd48120, 16'd61446, 16'd64036, 16'd42419, 16'd26196, 16'd63705, 16'd41302, 16'd62856, 16'd13000, 16'd35438, 16'd55459, 16'd27353, 16'd37175, 16'd15742, 16'd32137, 16'd64135, 16'd63262, 16'd31621, 16'd37457, 16'd43009, 16'd49113, 16'd11961});
	test_expansion(128'h0befb0a7298f8b14793a68e4ce44f0fd, {16'd56426, 16'd64338, 16'd21481, 16'd54096, 16'd28293, 16'd40955, 16'd37587, 16'd11238, 16'd62620, 16'd48224, 16'd41099, 16'd51759, 16'd34830, 16'd26451, 16'd13357, 16'd41037, 16'd26700, 16'd49973, 16'd47608, 16'd49053, 16'd49814, 16'd2340, 16'd39516, 16'd31605, 16'd62311, 16'd28698});
	test_expansion(128'h5830b209e31186e0e7cfd215d43d5c51, {16'd49744, 16'd28444, 16'd2268, 16'd15286, 16'd56181, 16'd12447, 16'd1776, 16'd39335, 16'd43723, 16'd8345, 16'd48659, 16'd8815, 16'd63581, 16'd11373, 16'd3236, 16'd32740, 16'd38073, 16'd9894, 16'd22432, 16'd48613, 16'd33274, 16'd14056, 16'd16174, 16'd58595, 16'd34894, 16'd47637});
	test_expansion(128'h096735514a56222dc2918c5289b3de51, {16'd6606, 16'd22199, 16'd22549, 16'd37299, 16'd21688, 16'd2717, 16'd63114, 16'd3765, 16'd48916, 16'd29408, 16'd29743, 16'd2491, 16'd21129, 16'd1209, 16'd9104, 16'd19813, 16'd3806, 16'd63449, 16'd9231, 16'd11869, 16'd49831, 16'd17829, 16'd60503, 16'd55090, 16'd32708, 16'd37447});
	test_expansion(128'h2e7b2cf4a7b71287ca43adfad79187c1, {16'd59801, 16'd28172, 16'd43110, 16'd48316, 16'd58710, 16'd10450, 16'd16859, 16'd57853, 16'd40222, 16'd14511, 16'd14230, 16'd9676, 16'd4824, 16'd48380, 16'd57745, 16'd33577, 16'd45517, 16'd59984, 16'd60824, 16'd20255, 16'd47850, 16'd2503, 16'd14485, 16'd22116, 16'd64570, 16'd58881});
	test_expansion(128'ha2cab02818bae320935ab4d944c92053, {16'd22761, 16'd38042, 16'd49023, 16'd9167, 16'd59596, 16'd13434, 16'd4646, 16'd57159, 16'd64791, 16'd10174, 16'd5315, 16'd60884, 16'd26052, 16'd34188, 16'd28906, 16'd28870, 16'd51713, 16'd28773, 16'd7744, 16'd64736, 16'd44267, 16'd31615, 16'd11145, 16'd60856, 16'd64388, 16'd10562});
	test_expansion(128'h491685c8f72661d60fee32f591168f59, {16'd34305, 16'd33698, 16'd48567, 16'd6475, 16'd45862, 16'd56730, 16'd44448, 16'd53065, 16'd29278, 16'd60284, 16'd27703, 16'd63439, 16'd6269, 16'd13406, 16'd30283, 16'd60839, 16'd5280, 16'd62310, 16'd8216, 16'd52411, 16'd46918, 16'd19280, 16'd36007, 16'd35588, 16'd349, 16'd28867});
	test_expansion(128'he543df49bc7e39377f8f5f96f157d211, {16'd55558, 16'd6773, 16'd29519, 16'd45156, 16'd18768, 16'd27305, 16'd40504, 16'd59424, 16'd27087, 16'd9574, 16'd23216, 16'd34428, 16'd63653, 16'd47096, 16'd7608, 16'd17227, 16'd31799, 16'd56256, 16'd32600, 16'd56105, 16'd29951, 16'd33065, 16'd59151, 16'd45468, 16'd35311, 16'd39349});
	test_expansion(128'he8f6d64907976e5033d4362195e833ad, {16'd6874, 16'd25261, 16'd30190, 16'd27653, 16'd60401, 16'd17574, 16'd57039, 16'd11213, 16'd16669, 16'd49182, 16'd18166, 16'd31734, 16'd40750, 16'd19141, 16'd12158, 16'd31395, 16'd62129, 16'd56856, 16'd48313, 16'd47660, 16'd19585, 16'd452, 16'd48044, 16'd27012, 16'd36257, 16'd48168});
	test_expansion(128'h7f7252fa033d54aff236d0adb9696fa0, {16'd31665, 16'd55418, 16'd17781, 16'd35804, 16'd30525, 16'd30578, 16'd19916, 16'd17573, 16'd64714, 16'd47236, 16'd1911, 16'd5514, 16'd42411, 16'd16444, 16'd30095, 16'd5303, 16'd59010, 16'd5419, 16'd1620, 16'd13621, 16'd32420, 16'd61770, 16'd5999, 16'd63615, 16'd28591, 16'd54332});
	test_expansion(128'h6267c782eb46eb0e7b20c140ec332d59, {16'd45747, 16'd47161, 16'd7629, 16'd53428, 16'd63306, 16'd50188, 16'd36420, 16'd46500, 16'd31230, 16'd26785, 16'd3679, 16'd8493, 16'd11201, 16'd30834, 16'd48425, 16'd15099, 16'd27350, 16'd63118, 16'd39315, 16'd57077, 16'd53149, 16'd55829, 16'd22941, 16'd27335, 16'd55589, 16'd48461});
	test_expansion(128'h869ef036b10a443587534d47d9943726, {16'd23854, 16'd3342, 16'd43391, 16'd1602, 16'd18706, 16'd4321, 16'd8153, 16'd15477, 16'd33037, 16'd51002, 16'd37858, 16'd29387, 16'd56300, 16'd9786, 16'd53890, 16'd25163, 16'd46972, 16'd27688, 16'd4173, 16'd12248, 16'd16316, 16'd7859, 16'd17217, 16'd650, 16'd57340, 16'd60870});
	test_expansion(128'hfa3afe3c143af47af2ad63d840d25dcb, {16'd17458, 16'd19645, 16'd17173, 16'd8547, 16'd57464, 16'd33345, 16'd1270, 16'd59365, 16'd15468, 16'd40117, 16'd22347, 16'd16480, 16'd55953, 16'd36625, 16'd46175, 16'd54242, 16'd64645, 16'd10808, 16'd35804, 16'd22866, 16'd418, 16'd14928, 16'd39628, 16'd12681, 16'd60777, 16'd4611});
	test_expansion(128'h3bc9a7b1c6a859d7cb52c5673f975daf, {16'd30299, 16'd1488, 16'd9973, 16'd3818, 16'd36462, 16'd46535, 16'd44429, 16'd34440, 16'd47348, 16'd61081, 16'd28576, 16'd38301, 16'd23631, 16'd19272, 16'd43017, 16'd31853, 16'd56438, 16'd585, 16'd10630, 16'd19899, 16'd53021, 16'd29752, 16'd5255, 16'd13546, 16'd54575, 16'd42720});
	test_expansion(128'h2a637e5a2e03986c16333626f440f463, {16'd63032, 16'd50244, 16'd49973, 16'd12610, 16'd60386, 16'd28985, 16'd24937, 16'd64799, 16'd60214, 16'd53864, 16'd33886, 16'd21124, 16'd29972, 16'd44191, 16'd28526, 16'd5754, 16'd2712, 16'd39325, 16'd43342, 16'd26501, 16'd45640, 16'd41154, 16'd37714, 16'd5447, 16'd57091, 16'd38521});
	test_expansion(128'he14cf3108922b764a0064c642ee5447b, {16'd42947, 16'd131, 16'd44985, 16'd31861, 16'd51572, 16'd50723, 16'd52473, 16'd11839, 16'd17838, 16'd448, 16'd45949, 16'd17730, 16'd7632, 16'd63495, 16'd16678, 16'd49755, 16'd19273, 16'd28164, 16'd17805, 16'd38443, 16'd43055, 16'd38708, 16'd13649, 16'd40554, 16'd47188, 16'd15142});
	test_expansion(128'hf58f090d450832387545033476aeb469, {16'd13970, 16'd9268, 16'd60730, 16'd13864, 16'd9620, 16'd39641, 16'd18506, 16'd17429, 16'd61438, 16'd38062, 16'd18382, 16'd60604, 16'd28199, 16'd12202, 16'd49897, 16'd11738, 16'd14177, 16'd40958, 16'd42553, 16'd22054, 16'd26258, 16'd1612, 16'd37557, 16'd12680, 16'd61304, 16'd9643});
	test_expansion(128'h3b51c5da3bf235aa527c1c05dee8dc7d, {16'd54192, 16'd712, 16'd58548, 16'd35576, 16'd31759, 16'd55700, 16'd18217, 16'd44410, 16'd45039, 16'd60135, 16'd53659, 16'd12811, 16'd36966, 16'd62869, 16'd30944, 16'd28897, 16'd29463, 16'd6952, 16'd53917, 16'd45227, 16'd18314, 16'd46195, 16'd19000, 16'd34208, 16'd35905, 16'd21943});
	test_expansion(128'h678548539c183ff0e7044d2362992e9c, {16'd15330, 16'd5336, 16'd52467, 16'd2072, 16'd64027, 16'd20499, 16'd42252, 16'd18923, 16'd41179, 16'd53594, 16'd61381, 16'd35079, 16'd4191, 16'd20646, 16'd38628, 16'd1153, 16'd2347, 16'd52017, 16'd55842, 16'd49100, 16'd35159, 16'd13303, 16'd56017, 16'd20000, 16'd61929, 16'd59599});
	test_expansion(128'h3338a27c8f9e4bd11b38c5ee7536263e, {16'd3484, 16'd36125, 16'd37029, 16'd40872, 16'd59652, 16'd45128, 16'd23912, 16'd6283, 16'd25521, 16'd34873, 16'd30954, 16'd61105, 16'd13434, 16'd56285, 16'd6689, 16'd63661, 16'd16283, 16'd38346, 16'd44012, 16'd1957, 16'd52130, 16'd1997, 16'd45536, 16'd61799, 16'd37754, 16'd42320});
	test_expansion(128'he36e64a2b932640a0699eafa23f2209f, {16'd52987, 16'd26748, 16'd37452, 16'd35632, 16'd48995, 16'd13766, 16'd49842, 16'd7839, 16'd14082, 16'd3719, 16'd17990, 16'd866, 16'd25712, 16'd9286, 16'd55798, 16'd23412, 16'd11035, 16'd34333, 16'd6077, 16'd13386, 16'd10368, 16'd52057, 16'd52123, 16'd35925, 16'd41000, 16'd6960});
	test_expansion(128'h70c109a6ba271ac3bf74a8d196d4375c, {16'd62001, 16'd2794, 16'd46106, 16'd39106, 16'd10904, 16'd976, 16'd42038, 16'd47996, 16'd64125, 16'd22512, 16'd370, 16'd4474, 16'd5898, 16'd53440, 16'd11275, 16'd62884, 16'd26193, 16'd38429, 16'd7781, 16'd47835, 16'd16459, 16'd2745, 16'd11000, 16'd53717, 16'd44239, 16'd61554});
	test_expansion(128'h821829911d265c3a8a1b3d8ddbd1dbc1, {16'd21795, 16'd12653, 16'd59019, 16'd52882, 16'd34337, 16'd10202, 16'd61131, 16'd36504, 16'd46953, 16'd48191, 16'd4031, 16'd11018, 16'd22919, 16'd53796, 16'd57957, 16'd23349, 16'd32863, 16'd50482, 16'd62623, 16'd55556, 16'd60718, 16'd54147, 16'd61578, 16'd3665, 16'd54194, 16'd33808});
	test_expansion(128'h4eaf98e4d30bc5ea96ea1b121d765cb9, {16'd40652, 16'd44491, 16'd159, 16'd17074, 16'd21613, 16'd44715, 16'd64377, 16'd8282, 16'd3746, 16'd25103, 16'd2509, 16'd53872, 16'd30140, 16'd13252, 16'd7109, 16'd18855, 16'd24751, 16'd32437, 16'd14975, 16'd45845, 16'd4700, 16'd42600, 16'd16089, 16'd44257, 16'd16537, 16'd56048});
	test_expansion(128'hfb5b3f0c1169b7dddce43630ca2e25ca, {16'd63075, 16'd59369, 16'd18776, 16'd29917, 16'd30122, 16'd64976, 16'd24838, 16'd53197, 16'd34261, 16'd58182, 16'd12774, 16'd725, 16'd23069, 16'd18684, 16'd32874, 16'd51236, 16'd54792, 16'd5176, 16'd48281, 16'd26701, 16'd6740, 16'd20105, 16'd14252, 16'd9026, 16'd45554, 16'd5034});
	test_expansion(128'h31b560351d394f9e91fefe6ab12cabc2, {16'd54806, 16'd34406, 16'd27116, 16'd41088, 16'd54486, 16'd9985, 16'd56096, 16'd29224, 16'd4306, 16'd23752, 16'd44444, 16'd64166, 16'd51346, 16'd61497, 16'd13783, 16'd24721, 16'd4444, 16'd25678, 16'd27977, 16'd3652, 16'd30880, 16'd32284, 16'd49617, 16'd9289, 16'd52288, 16'd55408});
	test_expansion(128'hd6bbbc5015828b8fcd074d3442a08858, {16'd50330, 16'd17530, 16'd3431, 16'd19867, 16'd37599, 16'd23476, 16'd1979, 16'd13241, 16'd5557, 16'd12335, 16'd2805, 16'd34094, 16'd58657, 16'd55772, 16'd9779, 16'd15596, 16'd54292, 16'd45887, 16'd42962, 16'd6649, 16'd22364, 16'd16303, 16'd35076, 16'd34905, 16'd28187, 16'd34390});
	test_expansion(128'ha646cb7ab4f17d9f72585a25a57bbb9d, {16'd54975, 16'd19932, 16'd20572, 16'd26557, 16'd34353, 16'd49759, 16'd17053, 16'd15693, 16'd11944, 16'd44596, 16'd2106, 16'd235, 16'd52191, 16'd55022, 16'd21004, 16'd63796, 16'd56819, 16'd13778, 16'd12408, 16'd53481, 16'd48614, 16'd39519, 16'd47509, 16'd49733, 16'd34048, 16'd39368});
	test_expansion(128'hd6be790120ab25d39dec383f3d1d57dc, {16'd47461, 16'd20306, 16'd24009, 16'd53058, 16'd43787, 16'd59764, 16'd43200, 16'd8658, 16'd4324, 16'd25021, 16'd58075, 16'd8857, 16'd9126, 16'd18786, 16'd18324, 16'd52235, 16'd29171, 16'd55300, 16'd4775, 16'd52011, 16'd63519, 16'd8305, 16'd57562, 16'd14245, 16'd32164, 16'd5064});
	test_expansion(128'h123e6bb8ead3968b810cab951a8c7580, {16'd17696, 16'd47010, 16'd52459, 16'd24498, 16'd54104, 16'd23505, 16'd19838, 16'd43180, 16'd6697, 16'd61790, 16'd17438, 16'd7920, 16'd10514, 16'd30138, 16'd37317, 16'd9341, 16'd2661, 16'd32772, 16'd61493, 16'd19599, 16'd17612, 16'd7335, 16'd35645, 16'd56244, 16'd18333, 16'd21198});
	test_expansion(128'hee71f9e8f0264c6792cbd3bdde2780ec, {16'd40262, 16'd47945, 16'd3791, 16'd7769, 16'd52293, 16'd35871, 16'd59929, 16'd51428, 16'd20296, 16'd36664, 16'd273, 16'd40787, 16'd36661, 16'd24834, 16'd24366, 16'd45654, 16'd7629, 16'd40202, 16'd2410, 16'd14852, 16'd16773, 16'd53980, 16'd36204, 16'd61496, 16'd23577, 16'd61514});
	test_expansion(128'h19b5c673f2123580a60c32aed5a65a62, {16'd18359, 16'd64627, 16'd39170, 16'd28544, 16'd34861, 16'd33421, 16'd22306, 16'd39631, 16'd61810, 16'd60402, 16'd63526, 16'd60540, 16'd5701, 16'd45604, 16'd23545, 16'd40650, 16'd4279, 16'd22567, 16'd2580, 16'd35093, 16'd41086, 16'd56185, 16'd21319, 16'd23593, 16'd48700, 16'd47474});
	test_expansion(128'h1239920b064e37aff695b58595920187, {16'd27442, 16'd21962, 16'd42870, 16'd22142, 16'd11231, 16'd64914, 16'd54230, 16'd10148, 16'd24918, 16'd23339, 16'd13926, 16'd46136, 16'd41846, 16'd19573, 16'd57438, 16'd31365, 16'd19969, 16'd39461, 16'd28412, 16'd14785, 16'd34627, 16'd30662, 16'd4932, 16'd1443, 16'd9428, 16'd19256});
	test_expansion(128'hc7bf1f2df1f673392824aad29db1de82, {16'd26184, 16'd65427, 16'd60565, 16'd36792, 16'd32885, 16'd49662, 16'd40554, 16'd57351, 16'd27091, 16'd17077, 16'd44472, 16'd26313, 16'd51523, 16'd53644, 16'd56295, 16'd53781, 16'd33970, 16'd49012, 16'd9211, 16'd58303, 16'd44358, 16'd54222, 16'd57048, 16'd48710, 16'd18754, 16'd22784});
	test_expansion(128'h5db54e4e1307102c02e37d2346a0c58a, {16'd6458, 16'd56224, 16'd34589, 16'd63653, 16'd51228, 16'd60567, 16'd34649, 16'd65409, 16'd12498, 16'd26560, 16'd12803, 16'd45638, 16'd5063, 16'd11686, 16'd62464, 16'd3850, 16'd21204, 16'd33607, 16'd30953, 16'd55869, 16'd31372, 16'd49626, 16'd53828, 16'd26189, 16'd52435, 16'd58285});
	test_expansion(128'h2530d5e1622927ebcebaf95f764efb23, {16'd18908, 16'd58024, 16'd22959, 16'd53910, 16'd58044, 16'd50278, 16'd16445, 16'd7564, 16'd52348, 16'd36067, 16'd13487, 16'd33879, 16'd10768, 16'd54009, 16'd56018, 16'd21173, 16'd12134, 16'd4612, 16'd49952, 16'd33207, 16'd51125, 16'd31588, 16'd24772, 16'd53671, 16'd55938, 16'd42101});
	test_expansion(128'hd512d86a280147b5ced7e420828e2f59, {16'd12352, 16'd7208, 16'd31616, 16'd38335, 16'd63245, 16'd46129, 16'd58063, 16'd27404, 16'd14708, 16'd29214, 16'd62084, 16'd10650, 16'd62409, 16'd14301, 16'd51766, 16'd48513, 16'd58571, 16'd31077, 16'd31784, 16'd153, 16'd33803, 16'd8096, 16'd7139, 16'd59807, 16'd38451, 16'd16509});
	test_expansion(128'hb4f7bb8fc96d0453b4cc3767b8889736, {16'd30251, 16'd20071, 16'd32803, 16'd36720, 16'd8860, 16'd50174, 16'd16876, 16'd24758, 16'd12669, 16'd45844, 16'd64308, 16'd37959, 16'd52143, 16'd20042, 16'd6605, 16'd25854, 16'd46294, 16'd50046, 16'd17474, 16'd19144, 16'd6524, 16'd20337, 16'd50891, 16'd32297, 16'd63496, 16'd25118});
	test_expansion(128'h89f74428f658c790010b717aedcfaffd, {16'd11855, 16'd5252, 16'd42053, 16'd10362, 16'd9749, 16'd5896, 16'd59471, 16'd61866, 16'd1170, 16'd64800, 16'd32073, 16'd60084, 16'd45639, 16'd38335, 16'd49170, 16'd28511, 16'd6653, 16'd15390, 16'd29919, 16'd53694, 16'd37753, 16'd12789, 16'd26093, 16'd39236, 16'd12681, 16'd2366});
	test_expansion(128'h79862200ac9681ccd3d3505e723907e9, {16'd39067, 16'd19436, 16'd24773, 16'd26237, 16'd205, 16'd41435, 16'd52164, 16'd10517, 16'd60317, 16'd3364, 16'd35758, 16'd20615, 16'd61179, 16'd16406, 16'd42121, 16'd24909, 16'd25394, 16'd30283, 16'd38373, 16'd61880, 16'd38646, 16'd60650, 16'd19407, 16'd23708, 16'd40361, 16'd9314});
	test_expansion(128'hf4852588a02002c07e0e47baecae21e4, {16'd4634, 16'd62253, 16'd8588, 16'd17218, 16'd19392, 16'd58952, 16'd39348, 16'd43641, 16'd7387, 16'd59359, 16'd54936, 16'd15076, 16'd10371, 16'd3150, 16'd41139, 16'd22232, 16'd49889, 16'd62302, 16'd27117, 16'd60685, 16'd46353, 16'd8985, 16'd32123, 16'd62932, 16'd37445, 16'd19936});
	test_expansion(128'h55b18ac0964c0e1aab50bb65dc855f86, {16'd4936, 16'd56467, 16'd42154, 16'd45305, 16'd4528, 16'd63740, 16'd41037, 16'd4714, 16'd55636, 16'd46337, 16'd63990, 16'd56168, 16'd48767, 16'd4184, 16'd48124, 16'd51839, 16'd40670, 16'd61685, 16'd7463, 16'd16185, 16'd13916, 16'd28496, 16'd13183, 16'd56826, 16'd10767, 16'd28393});
	test_expansion(128'h24222d18995766aec66547d1b735d079, {16'd39721, 16'd50623, 16'd58253, 16'd20709, 16'd39543, 16'd30194, 16'd59058, 16'd5879, 16'd14141, 16'd29390, 16'd42435, 16'd48139, 16'd28036, 16'd41637, 16'd29001, 16'd3298, 16'd53479, 16'd30454, 16'd49623, 16'd51828, 16'd61313, 16'd30744, 16'd37741, 16'd56284, 16'd56777, 16'd19294});
	test_expansion(128'ha2cd8f2f2ce75cf6503db6c0e6402eb0, {16'd3923, 16'd29428, 16'd31449, 16'd50631, 16'd53673, 16'd20379, 16'd11811, 16'd9170, 16'd23502, 16'd40946, 16'd59153, 16'd25980, 16'd46026, 16'd11349, 16'd22265, 16'd32126, 16'd29626, 16'd16482, 16'd32225, 16'd7999, 16'd9539, 16'd64008, 16'd40570, 16'd24580, 16'd59709, 16'd18310});
	test_expansion(128'h077a3808ad36ae6e767bc86d0d480058, {16'd14703, 16'd42578, 16'd55511, 16'd14637, 16'd58341, 16'd11349, 16'd60666, 16'd22796, 16'd8847, 16'd53702, 16'd44368, 16'd32888, 16'd61385, 16'd688, 16'd20563, 16'd53243, 16'd57850, 16'd9336, 16'd43566, 16'd15506, 16'd29550, 16'd36617, 16'd7608, 16'd2617, 16'd29998, 16'd23017});
	test_expansion(128'h8b75073a4d3071236f7d6b733411f69a, {16'd57848, 16'd65212, 16'd63576, 16'd56639, 16'd46484, 16'd65214, 16'd6470, 16'd60327, 16'd22827, 16'd27066, 16'd17034, 16'd12911, 16'd62462, 16'd54639, 16'd6980, 16'd18172, 16'd23840, 16'd62301, 16'd55448, 16'd60454, 16'd28037, 16'd50990, 16'd54555, 16'd18620, 16'd49063, 16'd3153});
	test_expansion(128'hb7094438e41c37f84a21da227b71239e, {16'd41692, 16'd60163, 16'd39933, 16'd61011, 16'd41384, 16'd46816, 16'd62848, 16'd39308, 16'd25411, 16'd62525, 16'd50944, 16'd27735, 16'd52253, 16'd20288, 16'd37534, 16'd60168, 16'd6701, 16'd20581, 16'd43741, 16'd50201, 16'd42496, 16'd7851, 16'd41542, 16'd13304, 16'd59772, 16'd33160});
	test_expansion(128'h5808385e75f486c3f53173db9290ef5e, {16'd33693, 16'd151, 16'd11940, 16'd34264, 16'd21721, 16'd25334, 16'd41319, 16'd59809, 16'd18294, 16'd41367, 16'd13079, 16'd7497, 16'd8220, 16'd19688, 16'd9382, 16'd2278, 16'd40564, 16'd14087, 16'd46698, 16'd51667, 16'd54553, 16'd59657, 16'd21795, 16'd50182, 16'd6134, 16'd40487});
	test_expansion(128'h38a371f1b2e7834bb79e96b642a18cef, {16'd18883, 16'd65398, 16'd4265, 16'd40844, 16'd29069, 16'd58133, 16'd38383, 16'd49551, 16'd21146, 16'd21426, 16'd49287, 16'd24539, 16'd14929, 16'd61938, 16'd34731, 16'd10817, 16'd25168, 16'd12726, 16'd11040, 16'd42262, 16'd21857, 16'd51952, 16'd6835, 16'd20009, 16'd10206, 16'd29804});
	test_expansion(128'h7e1a284e54c037a934c11920566b36a8, {16'd49394, 16'd32781, 16'd49424, 16'd8142, 16'd5787, 16'd31316, 16'd64819, 16'd57123, 16'd50027, 16'd58648, 16'd48898, 16'd503, 16'd17194, 16'd52597, 16'd26831, 16'd37152, 16'd4258, 16'd20921, 16'd38067, 16'd16629, 16'd36834, 16'd60463, 16'd60546, 16'd54602, 16'd48963, 16'd17926});
	test_expansion(128'hd7f175f280b3519168b85a1484cff79c, {16'd10221, 16'd38839, 16'd5633, 16'd8821, 16'd3424, 16'd9386, 16'd28943, 16'd46322, 16'd55872, 16'd32262, 16'd60262, 16'd52451, 16'd20151, 16'd2707, 16'd57539, 16'd10115, 16'd61027, 16'd1283, 16'd63353, 16'd34232, 16'd57201, 16'd55647, 16'd54328, 16'd14478, 16'd44951, 16'd34346});
	test_expansion(128'hd9f0c567dcf484b16be2cd1ac97ed781, {16'd35324, 16'd61782, 16'd4267, 16'd63407, 16'd29702, 16'd30823, 16'd56054, 16'd17074, 16'd47242, 16'd42184, 16'd46613, 16'd2103, 16'd45929, 16'd21816, 16'd34840, 16'd35105, 16'd9476, 16'd33698, 16'd48798, 16'd21900, 16'd39282, 16'd6087, 16'd51676, 16'd26791, 16'd52926, 16'd5716});
	test_expansion(128'hd6ef82f872657ef15ae3cb2e9a95ab0b, {16'd26199, 16'd24120, 16'd8588, 16'd31662, 16'd60729, 16'd24655, 16'd43307, 16'd35177, 16'd44923, 16'd20974, 16'd27855, 16'd13567, 16'd27307, 16'd62055, 16'd64854, 16'd58084, 16'd40744, 16'd64208, 16'd20588, 16'd44935, 16'd11057, 16'd10430, 16'd56683, 16'd62176, 16'd16155, 16'd14132});
	test_expansion(128'h6401d401c67dcae986c84a10d60f9eaa, {16'd53282, 16'd31612, 16'd48830, 16'd31296, 16'd15884, 16'd42999, 16'd43724, 16'd31174, 16'd60390, 16'd17289, 16'd41745, 16'd5023, 16'd50889, 16'd32634, 16'd8172, 16'd18965, 16'd922, 16'd3520, 16'd57544, 16'd24251, 16'd57863, 16'd34872, 16'd16196, 16'd22873, 16'd61803, 16'd32706});
	test_expansion(128'hc2cbb28a7433f096dcb20941d17b122f, {16'd10831, 16'd20092, 16'd14216, 16'd30469, 16'd36055, 16'd48990, 16'd28081, 16'd4409, 16'd27057, 16'd12440, 16'd32224, 16'd7494, 16'd37273, 16'd60766, 16'd3005, 16'd21908, 16'd41270, 16'd15101, 16'd47240, 16'd14726, 16'd54597, 16'd18294, 16'd35258, 16'd13288, 16'd47369, 16'd34219});
	test_expansion(128'h50c9bf294755b9efb1f5a2f12ad55346, {16'd36302, 16'd49789, 16'd40786, 16'd22667, 16'd49332, 16'd56766, 16'd14885, 16'd15076, 16'd31068, 16'd11854, 16'd38856, 16'd45720, 16'd10255, 16'd64781, 16'd34119, 16'd17659, 16'd25531, 16'd23588, 16'd57850, 16'd29908, 16'd29303, 16'd24181, 16'd37159, 16'd48712, 16'd3414, 16'd47167});
	test_expansion(128'h662eafc7e229c7b6e4e8f44097e5f75c, {16'd17614, 16'd30149, 16'd59847, 16'd23460, 16'd29237, 16'd40737, 16'd37953, 16'd21477, 16'd49519, 16'd21943, 16'd47275, 16'd50503, 16'd34219, 16'd6605, 16'd43262, 16'd36685, 16'd63460, 16'd30014, 16'd32991, 16'd36907, 16'd47743, 16'd26925, 16'd48051, 16'd59797, 16'd19304, 16'd49430});
	test_expansion(128'he0c59aa2a2391d8964e9f6b2ea3e20df, {16'd34695, 16'd65021, 16'd58941, 16'd61310, 16'd63000, 16'd9026, 16'd22736, 16'd25611, 16'd26189, 16'd36905, 16'd41907, 16'd43991, 16'd25947, 16'd43525, 16'd38619, 16'd42464, 16'd35079, 16'd55933, 16'd4271, 16'd1365, 16'd15689, 16'd9838, 16'd50847, 16'd51022, 16'd12584, 16'd21204});
	test_expansion(128'hc1c655715b3b87b2a405f6aeac2a3f4d, {16'd61631, 16'd44700, 16'd55776, 16'd26466, 16'd62351, 16'd47797, 16'd20791, 16'd10844, 16'd6887, 16'd33424, 16'd48712, 16'd49165, 16'd35405, 16'd49446, 16'd10186, 16'd45416, 16'd15892, 16'd7782, 16'd49544, 16'd38118, 16'd12050, 16'd27265, 16'd62693, 16'd1406, 16'd40955, 16'd47435});
	test_expansion(128'h8de7c402190f72c351c88ad74492624c, {16'd57673, 16'd3681, 16'd60300, 16'd58574, 16'd33759, 16'd22045, 16'd14100, 16'd64275, 16'd11033, 16'd12545, 16'd40752, 16'd15733, 16'd10979, 16'd13814, 16'd15587, 16'd52969, 16'd53288, 16'd15547, 16'd6910, 16'd53243, 16'd31922, 16'd64678, 16'd6493, 16'd24835, 16'd33533, 16'd23289});
	test_expansion(128'h433bf7ab5fe42d7d7e46c08cc2b5dad9, {16'd48350, 16'd25840, 16'd46665, 16'd62531, 16'd40291, 16'd62793, 16'd37164, 16'd43814, 16'd54272, 16'd31191, 16'd63037, 16'd46849, 16'd22782, 16'd9276, 16'd4274, 16'd4111, 16'd33057, 16'd48281, 16'd35611, 16'd42085, 16'd37026, 16'd63109, 16'd2443, 16'd17011, 16'd47096, 16'd5602});
	test_expansion(128'h58272a70c78b88d1f9640f90f202f2fc, {16'd9904, 16'd9578, 16'd19946, 16'd43587, 16'd30848, 16'd54462, 16'd38176, 16'd43387, 16'd47010, 16'd49681, 16'd51262, 16'd40765, 16'd26622, 16'd33524, 16'd24040, 16'd14663, 16'd14664, 16'd57447, 16'd30496, 16'd56589, 16'd48931, 16'd239, 16'd29961, 16'd42557, 16'd19362, 16'd51944});
	test_expansion(128'hd66c0101b5dc404f88ab599e148b8ce8, {16'd47001, 16'd32639, 16'd44218, 16'd16282, 16'd44319, 16'd17699, 16'd31034, 16'd23370, 16'd43034, 16'd42030, 16'd43373, 16'd20898, 16'd8200, 16'd3312, 16'd51917, 16'd38340, 16'd13837, 16'd21770, 16'd13081, 16'd60247, 16'd61118, 16'd63095, 16'd30679, 16'd48631, 16'd17589, 16'd385});
	test_expansion(128'hfeb2552170bc191758c9889e42f7e261, {16'd2198, 16'd40120, 16'd26392, 16'd22898, 16'd126, 16'd29323, 16'd1049, 16'd30571, 16'd31666, 16'd20622, 16'd12893, 16'd4975, 16'd49606, 16'd49088, 16'd43025, 16'd27738, 16'd6234, 16'd51256, 16'd5469, 16'd29638, 16'd36145, 16'd11906, 16'd18380, 16'd24389, 16'd58196, 16'd21855});
	test_expansion(128'hca5e7bb82226c1e5990b84159d713085, {16'd19123, 16'd58735, 16'd48451, 16'd61419, 16'd5954, 16'd24562, 16'd1106, 16'd36390, 16'd48506, 16'd43899, 16'd25582, 16'd23091, 16'd23432, 16'd31993, 16'd65009, 16'd38980, 16'd35592, 16'd12929, 16'd44750, 16'd46038, 16'd33683, 16'd65273, 16'd27303, 16'd56004, 16'd43399, 16'd29016});
	test_expansion(128'hb48dab13f0c65832c30d180dbf857d5f, {16'd27682, 16'd8177, 16'd50865, 16'd577, 16'd65094, 16'd24104, 16'd2601, 16'd54985, 16'd16, 16'd34335, 16'd19866, 16'd52277, 16'd7419, 16'd36327, 16'd47143, 16'd26334, 16'd47125, 16'd35730, 16'd59552, 16'd5500, 16'd18587, 16'd35268, 16'd59930, 16'd64132, 16'd58383, 16'd50231});
	test_expansion(128'hc7edd971a3f56607682babfbc0494325, {16'd56692, 16'd15036, 16'd65229, 16'd54158, 16'd45732, 16'd1896, 16'd8158, 16'd17174, 16'd57728, 16'd16503, 16'd62253, 16'd560, 16'd48498, 16'd58094, 16'd7232, 16'd18609, 16'd44420, 16'd2369, 16'd62955, 16'd30920, 16'd33501, 16'd30938, 16'd3245, 16'd28221, 16'd1359, 16'd27231});
	test_expansion(128'h3ac5a37b3ce00238d87dd5914f126b50, {16'd37350, 16'd64617, 16'd22984, 16'd19211, 16'd45235, 16'd45912, 16'd11991, 16'd59477, 16'd25037, 16'd53484, 16'd47644, 16'd36626, 16'd38420, 16'd35165, 16'd57018, 16'd716, 16'd2226, 16'd28110, 16'd57093, 16'd3608, 16'd19627, 16'd58680, 16'd8572, 16'd13483, 16'd25779, 16'd5088});
	test_expansion(128'h1f83ba5c77538eb8ee243f6f27707763, {16'd61535, 16'd47036, 16'd64557, 16'd20237, 16'd16110, 16'd3373, 16'd12695, 16'd11076, 16'd16331, 16'd63440, 16'd23457, 16'd11826, 16'd20970, 16'd50937, 16'd2916, 16'd19329, 16'd2778, 16'd63382, 16'd54563, 16'd49920, 16'd37257, 16'd47684, 16'd57333, 16'd41902, 16'd39385, 16'd35693});
	test_expansion(128'h754a96a6c69c6e2ed2cd8a5d79bc00da, {16'd51542, 16'd40574, 16'd8807, 16'd16761, 16'd33197, 16'd5878, 16'd6936, 16'd28704, 16'd24871, 16'd13964, 16'd39028, 16'd61619, 16'd53885, 16'd8914, 16'd63285, 16'd44774, 16'd15402, 16'd7474, 16'd20918, 16'd2942, 16'd45123, 16'd15380, 16'd41731, 16'd8711, 16'd38651, 16'd46973});
	test_expansion(128'h2d8c26a1327fd495f6b6b03d7bb66015, {16'd25676, 16'd18976, 16'd31387, 16'd54489, 16'd60148, 16'd9180, 16'd40365, 16'd32698, 16'd51013, 16'd4772, 16'd5991, 16'd37648, 16'd48545, 16'd34783, 16'd36693, 16'd34024, 16'd41947, 16'd13721, 16'd25216, 16'd22569, 16'd9730, 16'd40084, 16'd50887, 16'd51950, 16'd7074, 16'd19745});
	test_expansion(128'hd3f631a32055635179d48ffe079c25d4, {16'd10212, 16'd16073, 16'd48010, 16'd41917, 16'd52319, 16'd9657, 16'd63433, 16'd35069, 16'd41408, 16'd54578, 16'd47283, 16'd32385, 16'd16166, 16'd58116, 16'd146, 16'd5419, 16'd35601, 16'd52980, 16'd25594, 16'd38462, 16'd43442, 16'd60011, 16'd40988, 16'd28966, 16'd16813, 16'd33845});
	test_expansion(128'h8c52b6759cf093beecfd8f4995de3058, {16'd43988, 16'd40871, 16'd29589, 16'd14719, 16'd64072, 16'd21883, 16'd60165, 16'd58242, 16'd53930, 16'd12576, 16'd61604, 16'd29340, 16'd61748, 16'd58818, 16'd12183, 16'd12425, 16'd26536, 16'd58826, 16'd56717, 16'd8688, 16'd16199, 16'd1747, 16'd4737, 16'd19898, 16'd24457, 16'd34794});
	test_expansion(128'hb762a21ed4e2b47aee253e81211369d6, {16'd2490, 16'd37708, 16'd65224, 16'd19440, 16'd63514, 16'd21847, 16'd11370, 16'd30411, 16'd44386, 16'd48071, 16'd31444, 16'd37925, 16'd6908, 16'd49365, 16'd50996, 16'd21068, 16'd12505, 16'd25847, 16'd25813, 16'd17744, 16'd6695, 16'd28014, 16'd14622, 16'd16481, 16'd913, 16'd8883});
	test_expansion(128'h9e9eef21c0428e7fd636ae31a5ce1255, {16'd11302, 16'd31635, 16'd47343, 16'd8471, 16'd53107, 16'd33333, 16'd64080, 16'd61552, 16'd62118, 16'd60576, 16'd9345, 16'd57902, 16'd62325, 16'd28871, 16'd25291, 16'd16596, 16'd12334, 16'd26570, 16'd12233, 16'd58887, 16'd30070, 16'd58485, 16'd62307, 16'd7798, 16'd41713, 16'd62848});
	test_expansion(128'h5f67381b632d467956066d5869ad088f, {16'd27367, 16'd47346, 16'd45651, 16'd17148, 16'd50545, 16'd24390, 16'd5209, 16'd31868, 16'd63180, 16'd19456, 16'd11255, 16'd59639, 16'd17233, 16'd14442, 16'd5762, 16'd15213, 16'd51271, 16'd11486, 16'd42192, 16'd18693, 16'd32135, 16'd13859, 16'd40602, 16'd30759, 16'd52197, 16'd41177});
	test_expansion(128'h37b483c2931e11d06f770972c91fba45, {16'd16960, 16'd4907, 16'd36858, 16'd21553, 16'd54536, 16'd22955, 16'd52139, 16'd26321, 16'd9726, 16'd31201, 16'd20155, 16'd30842, 16'd11708, 16'd7291, 16'd16127, 16'd974, 16'd31924, 16'd29426, 16'd48655, 16'd49748, 16'd2703, 16'd28891, 16'd59312, 16'd13916, 16'd40810, 16'd42097});
	test_expansion(128'h8e126c0a07e72a54df32913205a1b74d, {16'd44673, 16'd8112, 16'd22089, 16'd14266, 16'd49806, 16'd50247, 16'd27892, 16'd44647, 16'd25476, 16'd63858, 16'd14256, 16'd7617, 16'd31008, 16'd50125, 16'd42369, 16'd11859, 16'd62900, 16'd724, 16'd38769, 16'd12478, 16'd34354, 16'd12538, 16'd47235, 16'd6781, 16'd43035, 16'd45630});
	test_expansion(128'h8705f5deb3da3caddfd42cad1cc6c6e8, {16'd10501, 16'd52230, 16'd19671, 16'd47942, 16'd59826, 16'd55637, 16'd742, 16'd58905, 16'd39371, 16'd44016, 16'd47702, 16'd40017, 16'd41543, 16'd36051, 16'd13311, 16'd3108, 16'd62003, 16'd22483, 16'd38361, 16'd56187, 16'd8170, 16'd55382, 16'd34390, 16'd10115, 16'd32253, 16'd38244});
	test_expansion(128'h844afb93e879f3098ecda13b6e8732c0, {16'd55421, 16'd4673, 16'd31013, 16'd48472, 16'd63359, 16'd22893, 16'd56231, 16'd9788, 16'd55332, 16'd58899, 16'd32617, 16'd9594, 16'd37058, 16'd57284, 16'd53850, 16'd27426, 16'd56936, 16'd5322, 16'd60954, 16'd59898, 16'd28321, 16'd25915, 16'd35537, 16'd10572, 16'd9831, 16'd6807});
	test_expansion(128'h7853fc736d990af61c03450a9a41dd35, {16'd50170, 16'd8179, 16'd6124, 16'd2012, 16'd61227, 16'd54284, 16'd3492, 16'd44134, 16'd346, 16'd4259, 16'd36382, 16'd59861, 16'd14932, 16'd62811, 16'd3166, 16'd45589, 16'd40027, 16'd6003, 16'd61739, 16'd62477, 16'd25411, 16'd51912, 16'd33332, 16'd23651, 16'd5794, 16'd19078});
	test_expansion(128'hfd19e75d0089d728c36206fa949c4403, {16'd44024, 16'd22406, 16'd29822, 16'd28566, 16'd62385, 16'd25212, 16'd20179, 16'd47555, 16'd41315, 16'd58460, 16'd8854, 16'd22039, 16'd37911, 16'd14595, 16'd62374, 16'd8809, 16'd39140, 16'd31537, 16'd64428, 16'd19156, 16'd24988, 16'd37439, 16'd52869, 16'd30075, 16'd58807, 16'd58062});
	test_expansion(128'h5d3a6a991aa6e5be36f7511b608f7abc, {16'd50460, 16'd33150, 16'd48343, 16'd50667, 16'd51507, 16'd55157, 16'd52616, 16'd44605, 16'd46997, 16'd61291, 16'd747, 16'd10062, 16'd41178, 16'd52987, 16'd16803, 16'd56313, 16'd12207, 16'd2282, 16'd28452, 16'd32969, 16'd11102, 16'd40678, 16'd22681, 16'd10375, 16'd1456, 16'd26759});
	test_expansion(128'h068242cc000ffc795cb83c0702521ec7, {16'd17378, 16'd3927, 16'd12179, 16'd2500, 16'd30722, 16'd48063, 16'd4509, 16'd51380, 16'd28825, 16'd64005, 16'd19528, 16'd38199, 16'd52567, 16'd34365, 16'd22913, 16'd50950, 16'd19727, 16'd40156, 16'd1023, 16'd61301, 16'd18494, 16'd54612, 16'd63726, 16'd29987, 16'd13680, 16'd29997});
	test_expansion(128'h6906474af414ceb2fbc3325cc3e8c580, {16'd19440, 16'd50507, 16'd3654, 16'd28898, 16'd12165, 16'd26691, 16'd22422, 16'd44189, 16'd39616, 16'd26633, 16'd47687, 16'd5167, 16'd18488, 16'd24627, 16'd21242, 16'd47409, 16'd43360, 16'd50826, 16'd36661, 16'd1834, 16'd10319, 16'd29826, 16'd28690, 16'd28214, 16'd24030, 16'd20984});
	test_expansion(128'hb17626a5d793c3fd3982ab9e09ec94bd, {16'd43134, 16'd14397, 16'd36938, 16'd40887, 16'd6679, 16'd30654, 16'd60143, 16'd5973, 16'd40661, 16'd17293, 16'd17077, 16'd12649, 16'd55310, 16'd61201, 16'd43806, 16'd32113, 16'd3791, 16'd58327, 16'd51813, 16'd7576, 16'd59599, 16'd9509, 16'd33803, 16'd6054, 16'd14418, 16'd40602});
	test_expansion(128'hc555fe6c7b348263ad28979ee1571bb4, {16'd33824, 16'd9493, 16'd15650, 16'd11834, 16'd37515, 16'd16848, 16'd35075, 16'd30192, 16'd24110, 16'd16567, 16'd56216, 16'd18736, 16'd50026, 16'd50286, 16'd55740, 16'd7682, 16'd13908, 16'd22181, 16'd58772, 16'd52174, 16'd51748, 16'd8084, 16'd43891, 16'd18037, 16'd41667, 16'd8342});
	test_expansion(128'heeca911587ca6655c0e5c5029abfd288, {16'd42404, 16'd34354, 16'd52620, 16'd48323, 16'd64570, 16'd55218, 16'd5497, 16'd52348, 16'd4755, 16'd40115, 16'd597, 16'd48726, 16'd45573, 16'd37261, 16'd44582, 16'd50457, 16'd10065, 16'd22565, 16'd57615, 16'd61448, 16'd36453, 16'd49900, 16'd13307, 16'd50776, 16'd33958, 16'd56833});
	test_expansion(128'h783e9fa4829404ee5f8dc37742875500, {16'd54668, 16'd51772, 16'd20366, 16'd29409, 16'd62534, 16'd11837, 16'd60500, 16'd26389, 16'd43695, 16'd59477, 16'd51139, 16'd44045, 16'd10689, 16'd35202, 16'd64231, 16'd44745, 16'd26271, 16'd11147, 16'd14092, 16'd54326, 16'd43413, 16'd44671, 16'd60241, 16'd31626, 16'd54709, 16'd8296});
	test_expansion(128'hce9178c556ab0ec6fb6d132935e5d03a, {16'd45612, 16'd55736, 16'd34926, 16'd52220, 16'd47792, 16'd54916, 16'd1998, 16'd28563, 16'd495, 16'd2089, 16'd23048, 16'd15271, 16'd26718, 16'd61458, 16'd51186, 16'd44898, 16'd36050, 16'd62885, 16'd18696, 16'd24660, 16'd29358, 16'd65490, 16'd58139, 16'd41567, 16'd9300, 16'd14441});
	test_expansion(128'h3da8cb9fd70c9a10d1c36d65d00ec05c, {16'd42456, 16'd55109, 16'd50611, 16'd44754, 16'd25639, 16'd2031, 16'd2809, 16'd53183, 16'd29587, 16'd50305, 16'd32684, 16'd34993, 16'd45615, 16'd43182, 16'd62690, 16'd45523, 16'd21478, 16'd54562, 16'd44138, 16'd32680, 16'd5037, 16'd35928, 16'd41964, 16'd11985, 16'd5495, 16'd40689});
	test_expansion(128'hb5ddf534efeb866a509e593024c3d737, {16'd13991, 16'd57507, 16'd53728, 16'd52262, 16'd35801, 16'd6463, 16'd50490, 16'd25697, 16'd38323, 16'd53177, 16'd39714, 16'd32788, 16'd41663, 16'd36666, 16'd22186, 16'd39027, 16'd29928, 16'd10723, 16'd43686, 16'd59417, 16'd42459, 16'd8579, 16'd12222, 16'd3035, 16'd25134, 16'd63778});
	test_expansion(128'h185f75729cd578a77bf7f0d5724e4870, {16'd36369, 16'd28655, 16'd24170, 16'd12680, 16'd62407, 16'd17645, 16'd59988, 16'd21837, 16'd63165, 16'd37581, 16'd50773, 16'd32715, 16'd61569, 16'd51481, 16'd22168, 16'd34922, 16'd38551, 16'd40576, 16'd586, 16'd11233, 16'd37837, 16'd42535, 16'd60961, 16'd2127, 16'd9584, 16'd53312});
	test_expansion(128'h88051e043c5c25db172f34e56e32ca29, {16'd8124, 16'd44678, 16'd2427, 16'd43745, 16'd33124, 16'd7654, 16'd9313, 16'd7689, 16'd58659, 16'd22289, 16'd65197, 16'd19499, 16'd7084, 16'd46419, 16'd7439, 16'd14677, 16'd17649, 16'd42641, 16'd46484, 16'd51821, 16'd25648, 16'd26328, 16'd7526, 16'd10191, 16'd40274, 16'd254});
	test_expansion(128'hac5fc06c1636e857aa7403e72aaeb62c, {16'd6113, 16'd33051, 16'd15222, 16'd5025, 16'd18122, 16'd21508, 16'd48879, 16'd52896, 16'd38264, 16'd5739, 16'd25222, 16'd9642, 16'd62605, 16'd7077, 16'd46636, 16'd40140, 16'd26029, 16'd5623, 16'd45675, 16'd58141, 16'd55349, 16'd59156, 16'd3300, 16'd46343, 16'd60290, 16'd9143});
	test_expansion(128'h3508563414d512f45d1a1b903dcfd63b, {16'd8446, 16'd32331, 16'd34519, 16'd51159, 16'd1968, 16'd2945, 16'd61245, 16'd18464, 16'd38113, 16'd61886, 16'd41251, 16'd57935, 16'd64647, 16'd2680, 16'd51242, 16'd4168, 16'd57182, 16'd21770, 16'd56034, 16'd30658, 16'd9314, 16'd48248, 16'd1155, 16'd62019, 16'd39977, 16'd26238});
	test_expansion(128'hd879d7117e617f990515eea23ca9282d, {16'd62917, 16'd9714, 16'd3728, 16'd62267, 16'd28705, 16'd46740, 16'd41214, 16'd13068, 16'd18859, 16'd41813, 16'd21076, 16'd25651, 16'd53423, 16'd332, 16'd19707, 16'd64369, 16'd58011, 16'd49086, 16'd15277, 16'd17812, 16'd23959, 16'd46615, 16'd11769, 16'd59780, 16'd353, 16'd53318});
	test_expansion(128'hd50bf7ce0f5b9d5e3bbb2b52c98ad0bf, {16'd7919, 16'd30125, 16'd36577, 16'd65037, 16'd1519, 16'd22005, 16'd37394, 16'd5453, 16'd4681, 16'd51389, 16'd46905, 16'd18504, 16'd53621, 16'd10536, 16'd52895, 16'd11334, 16'd10444, 16'd33173, 16'd39132, 16'd62758, 16'd61920, 16'd60452, 16'd18456, 16'd38084, 16'd35247, 16'd40941});
	test_expansion(128'hc51107e6faef8ebac475cec9ddb65829, {16'd62097, 16'd46272, 16'd16810, 16'd64090, 16'd60748, 16'd48026, 16'd6896, 16'd41178, 16'd8303, 16'd20086, 16'd62589, 16'd48719, 16'd12999, 16'd42345, 16'd24700, 16'd49793, 16'd6554, 16'd1495, 16'd18284, 16'd5817, 16'd59815, 16'd28033, 16'd55999, 16'd6360, 16'd45707, 16'd62629});
	test_expansion(128'ha38c8897c411bee3f33f474660fd019d, {16'd44421, 16'd29590, 16'd8758, 16'd52774, 16'd9855, 16'd21378, 16'd47370, 16'd53011, 16'd39254, 16'd61262, 16'd43485, 16'd65405, 16'd40043, 16'd65423, 16'd56440, 16'd60565, 16'd43334, 16'd50032, 16'd36787, 16'd10576, 16'd63169, 16'd40688, 16'd17856, 16'd23867, 16'd21418, 16'd21806});
	test_expansion(128'hf335eb66498f6e09a82d122e76165b06, {16'd20389, 16'd14769, 16'd28965, 16'd9321, 16'd59020, 16'd24262, 16'd3783, 16'd23670, 16'd62118, 16'd45205, 16'd35203, 16'd23188, 16'd45736, 16'd63010, 16'd46503, 16'd3167, 16'd48122, 16'd17412, 16'd63019, 16'd62623, 16'd47816, 16'd11988, 16'd15070, 16'd9989, 16'd32335, 16'd62207});
	test_expansion(128'h796be2029a38302fea772898e4a47513, {16'd56597, 16'd43880, 16'd15424, 16'd30063, 16'd62523, 16'd18184, 16'd22432, 16'd46226, 16'd11561, 16'd1951, 16'd11850, 16'd41070, 16'd62895, 16'd25338, 16'd40106, 16'd59991, 16'd50127, 16'd57796, 16'd46770, 16'd22901, 16'd15531, 16'd25945, 16'd56423, 16'd9718, 16'd55003, 16'd20905});
	test_expansion(128'he850ca1fab10a7768b2ae9caa994c5b1, {16'd22497, 16'd55833, 16'd9743, 16'd58995, 16'd62013, 16'd50748, 16'd50699, 16'd9773, 16'd21623, 16'd18538, 16'd59562, 16'd47529, 16'd43067, 16'd37745, 16'd35348, 16'd8736, 16'd27932, 16'd4371, 16'd34164, 16'd18684, 16'd24276, 16'd43153, 16'd28410, 16'd56133, 16'd7416, 16'd47322});
	test_expansion(128'hd30fb3a308d86640261e7d3d0a581f5c, {16'd28472, 16'd21874, 16'd59811, 16'd18621, 16'd37441, 16'd9446, 16'd26893, 16'd15257, 16'd42908, 16'd43914, 16'd60452, 16'd48836, 16'd26791, 16'd7933, 16'd37949, 16'd51594, 16'd23420, 16'd26210, 16'd48162, 16'd35435, 16'd20268, 16'd21865, 16'd12425, 16'd24619, 16'd9707, 16'd23733});
	test_expansion(128'h12473a904461152dd328d46abf218e62, {16'd27740, 16'd63568, 16'd9225, 16'd14394, 16'd49438, 16'd26707, 16'd51252, 16'd21621, 16'd10142, 16'd17649, 16'd23255, 16'd44144, 16'd63082, 16'd20921, 16'd23609, 16'd48469, 16'd42737, 16'd28640, 16'd5799, 16'd8345, 16'd44109, 16'd39515, 16'd49028, 16'd1546, 16'd38214, 16'd14311});
	test_expansion(128'hcf50deb3fdccf4040d0715f9df47a4d7, {16'd63707, 16'd53049, 16'd10515, 16'd22562, 16'd19934, 16'd21326, 16'd1041, 16'd56783, 16'd6763, 16'd12978, 16'd3917, 16'd38556, 16'd54019, 16'd3406, 16'd32955, 16'd41103, 16'd34091, 16'd37371, 16'd48183, 16'd13708, 16'd24534, 16'd28998, 16'd21731, 16'd20101, 16'd35416, 16'd47490});
	test_expansion(128'h866c46ea95d9beb7a9ad01a9cee28e93, {16'd43968, 16'd46543, 16'd39903, 16'd47032, 16'd8379, 16'd16363, 16'd21823, 16'd7985, 16'd44399, 16'd23042, 16'd43847, 16'd64571, 16'd42486, 16'd47000, 16'd45289, 16'd11159, 16'd10418, 16'd25381, 16'd47854, 16'd18517, 16'd5088, 16'd30380, 16'd28839, 16'd54688, 16'd65483, 16'd31131});
	test_expansion(128'h8f2d8b5db4989e9fd607e5662d2fe1da, {16'd53959, 16'd4460, 16'd7942, 16'd6711, 16'd28857, 16'd35065, 16'd62904, 16'd49548, 16'd40630, 16'd42935, 16'd55891, 16'd24340, 16'd1478, 16'd55068, 16'd37402, 16'd39886, 16'd16918, 16'd13465, 16'd17646, 16'd44094, 16'd43197, 16'd49060, 16'd6595, 16'd32772, 16'd16693, 16'd63928});
	test_expansion(128'hd76dc3c43cd899c7c2d739e9986cec7c, {16'd36875, 16'd63047, 16'd56903, 16'd30812, 16'd14478, 16'd18509, 16'd28768, 16'd23955, 16'd55747, 16'd34536, 16'd14702, 16'd21822, 16'd49994, 16'd7594, 16'd57023, 16'd21268, 16'd14658, 16'd2704, 16'd55072, 16'd5709, 16'd30445, 16'd56351, 16'd64850, 16'd5035, 16'd17873, 16'd7269});
	test_expansion(128'h1de031dc02093f559d773e6f92e7f6fd, {16'd46408, 16'd25088, 16'd29977, 16'd7678, 16'd6663, 16'd10663, 16'd45428, 16'd26786, 16'd58510, 16'd10897, 16'd23523, 16'd20280, 16'd59462, 16'd13708, 16'd63500, 16'd17943, 16'd6856, 16'd44384, 16'd36580, 16'd253, 16'd36462, 16'd11126, 16'd33925, 16'd42703, 16'd19080, 16'd63344});
	test_expansion(128'h4dde530d35ff92becd6e2ca002316c71, {16'd35891, 16'd2203, 16'd20751, 16'd9830, 16'd50420, 16'd45673, 16'd25688, 16'd8792, 16'd62069, 16'd63966, 16'd38714, 16'd32924, 16'd26443, 16'd2764, 16'd59813, 16'd59868, 16'd59363, 16'd63262, 16'd36061, 16'd9000, 16'd24255, 16'd29214, 16'd12047, 16'd28050, 16'd5963, 16'd32384});
	test_expansion(128'h31835e4353449b3236c93d26706156bb, {16'd21624, 16'd27480, 16'd60301, 16'd40494, 16'd42703, 16'd48382, 16'd32658, 16'd24215, 16'd46919, 16'd25224, 16'd38230, 16'd25635, 16'd28804, 16'd27286, 16'd46758, 16'd58952, 16'd23141, 16'd5482, 16'd20167, 16'd49132, 16'd45764, 16'd54059, 16'd50100, 16'd54123, 16'd29507, 16'd24197});
	test_expansion(128'hd527732874a86d6578c46a08ef8e7c35, {16'd20322, 16'd946, 16'd44716, 16'd11016, 16'd125, 16'd10789, 16'd63008, 16'd29893, 16'd19018, 16'd7249, 16'd37556, 16'd59320, 16'd14258, 16'd56875, 16'd21261, 16'd11018, 16'd21796, 16'd53241, 16'd42664, 16'd44443, 16'd33165, 16'd37388, 16'd25802, 16'd21866, 16'd10440, 16'd19806});
	test_expansion(128'h22e7732b5383e3a6d7c95b7cb4451d96, {16'd965, 16'd29483, 16'd46118, 16'd33254, 16'd1539, 16'd15293, 16'd31385, 16'd40699, 16'd31183, 16'd33161, 16'd32803, 16'd28626, 16'd31593, 16'd33384, 16'd25110, 16'd62761, 16'd2476, 16'd16420, 16'd3335, 16'd15147, 16'd21524, 16'd667, 16'd35086, 16'd62611, 16'd48759, 16'd33306});
	test_expansion(128'h6eb827ab730ad801ea6aaebd995ff9dd, {16'd42974, 16'd59571, 16'd30132, 16'd37287, 16'd17178, 16'd8232, 16'd51860, 16'd53833, 16'd48135, 16'd18554, 16'd24753, 16'd39156, 16'd17076, 16'd1365, 16'd25136, 16'd64825, 16'd24598, 16'd20831, 16'd57969, 16'd14975, 16'd8214, 16'd10404, 16'd56469, 16'd48761, 16'd52024, 16'd23981});
	test_expansion(128'h59bc57e075787c311d96e9a5c55deb1c, {16'd30315, 16'd47037, 16'd29152, 16'd24035, 16'd46365, 16'd31598, 16'd32951, 16'd57620, 16'd39793, 16'd34985, 16'd42236, 16'd839, 16'd9675, 16'd2871, 16'd22313, 16'd38368, 16'd29842, 16'd16581, 16'd53740, 16'd28908, 16'd16600, 16'd63986, 16'd63398, 16'd46472, 16'd24904, 16'd46490});
	test_expansion(128'h03b62063474e681d2613ce657b90ea42, {16'd55038, 16'd42825, 16'd16091, 16'd16315, 16'd36347, 16'd62919, 16'd16295, 16'd293, 16'd30589, 16'd44877, 16'd43579, 16'd36720, 16'd59811, 16'd45759, 16'd44215, 16'd18496, 16'd61035, 16'd37498, 16'd31294, 16'd8950, 16'd5432, 16'd2442, 16'd34130, 16'd59319, 16'd1637, 16'd32391});
	test_expansion(128'hba610795a6e3d4abb27b6da544bcd3ca, {16'd64547, 16'd9255, 16'd48736, 16'd12555, 16'd48157, 16'd52475, 16'd23865, 16'd40088, 16'd22072, 16'd5696, 16'd54142, 16'd17364, 16'd18254, 16'd34534, 16'd49599, 16'd42327, 16'd35754, 16'd15544, 16'd17992, 16'd60785, 16'd20408, 16'd12212, 16'd14748, 16'd48548, 16'd4267, 16'd397});
	test_expansion(128'h3aaf84d16a2c4f6d4c9d9829a5b892ca, {16'd15348, 16'd33788, 16'd1983, 16'd19353, 16'd42046, 16'd33358, 16'd2544, 16'd25004, 16'd29541, 16'd43435, 16'd12379, 16'd40124, 16'd5985, 16'd29330, 16'd37302, 16'd8526, 16'd27328, 16'd36891, 16'd7780, 16'd52870, 16'd11962, 16'd32858, 16'd21235, 16'd36276, 16'd47139, 16'd41629});
	test_expansion(128'h1a40ef17694a7a64a6b4c5b32746f1fd, {16'd18850, 16'd10151, 16'd19460, 16'd14581, 16'd60936, 16'd64200, 16'd6786, 16'd33411, 16'd8778, 16'd4002, 16'd28122, 16'd63529, 16'd48296, 16'd4989, 16'd34723, 16'd43591, 16'd27331, 16'd53689, 16'd8417, 16'd21498, 16'd22037, 16'd50673, 16'd31716, 16'd57263, 16'd5460, 16'd60688});
	test_expansion(128'h71688d8eba59cdd83d6e9eb56a43c865, {16'd14995, 16'd348, 16'd59286, 16'd657, 16'd60970, 16'd23153, 16'd8803, 16'd22833, 16'd10378, 16'd5202, 16'd55522, 16'd808, 16'd6535, 16'd2253, 16'd19872, 16'd44865, 16'd63095, 16'd45814, 16'd53662, 16'd28366, 16'd36043, 16'd62260, 16'd3059, 16'd23945, 16'd16633, 16'd3307});
	test_expansion(128'haa1af81bb78f33f522e6c568b6831ca5, {16'd21282, 16'd46540, 16'd58232, 16'd61995, 16'd18078, 16'd17985, 16'd4886, 16'd10356, 16'd29922, 16'd1310, 16'd10627, 16'd4578, 16'd20726, 16'd9525, 16'd10607, 16'd22874, 16'd54653, 16'd59437, 16'd3372, 16'd43307, 16'd31288, 16'd45819, 16'd42738, 16'd7478, 16'd45436, 16'd57627});
	test_expansion(128'hc63b9d96dbe96e0d2c586a0937ebe44b, {16'd3475, 16'd29950, 16'd37392, 16'd56919, 16'd11407, 16'd60099, 16'd63212, 16'd34327, 16'd297, 16'd24288, 16'd39231, 16'd15108, 16'd38299, 16'd42306, 16'd40256, 16'd24525, 16'd48100, 16'd50798, 16'd31801, 16'd49947, 16'd40738, 16'd20011, 16'd15985, 16'd57940, 16'd13938, 16'd20102});
	test_expansion(128'h26c84fa086629a5b46bdf7499269e645, {16'd55513, 16'd14542, 16'd15047, 16'd11137, 16'd2325, 16'd47825, 16'd15441, 16'd43141, 16'd38149, 16'd36618, 16'd51297, 16'd19479, 16'd63124, 16'd21776, 16'd51367, 16'd42650, 16'd30505, 16'd10027, 16'd35147, 16'd15592, 16'd57865, 16'd47373, 16'd13727, 16'd17694, 16'd6938, 16'd59517});
	test_expansion(128'hd42349c153292feb013ad97a7233834b, {16'd6377, 16'd4139, 16'd50201, 16'd35444, 16'd61396, 16'd42654, 16'd25665, 16'd4087, 16'd34617, 16'd1017, 16'd20650, 16'd28752, 16'd17078, 16'd30642, 16'd32139, 16'd20096, 16'd25385, 16'd58028, 16'd30243, 16'd28685, 16'd34388, 16'd35287, 16'd35883, 16'd53275, 16'd23017, 16'd14175});
	test_expansion(128'h5dab25cb460d85c54c6e5888921d777c, {16'd37285, 16'd9655, 16'd38130, 16'd35519, 16'd49345, 16'd51903, 16'd30823, 16'd32948, 16'd60774, 16'd62074, 16'd73, 16'd64012, 16'd18353, 16'd17873, 16'd14388, 16'd33906, 16'd11859, 16'd956, 16'd47321, 16'd34007, 16'd33626, 16'd6855, 16'd20870, 16'd41928, 16'd58434, 16'd44770});
	test_expansion(128'h32155795869c7c3ccf24bdb9c63b34a6, {16'd37880, 16'd11448, 16'd59891, 16'd2916, 16'd13706, 16'd54691, 16'd26109, 16'd65012, 16'd54925, 16'd50709, 16'd65256, 16'd52903, 16'd22011, 16'd46077, 16'd17140, 16'd8235, 16'd39455, 16'd25568, 16'd14560, 16'd10363, 16'd39670, 16'd27490, 16'd57219, 16'd21365, 16'd134, 16'd11000});
	test_expansion(128'hd693fc29a4fc40d4b2630e5b632be9ec, {16'd13863, 16'd33756, 16'd214, 16'd3732, 16'd20146, 16'd5799, 16'd6388, 16'd35759, 16'd11420, 16'd19983, 16'd25836, 16'd49009, 16'd61945, 16'd17282, 16'd30254, 16'd61175, 16'd40839, 16'd54206, 16'd29301, 16'd17821, 16'd52246, 16'd25481, 16'd64534, 16'd26499, 16'd44927, 16'd52412});
	test_expansion(128'h097d65ae1528c07de824406cce6d66ea, {16'd17182, 16'd35164, 16'd45768, 16'd22146, 16'd1180, 16'd36190, 16'd3359, 16'd26066, 16'd65228, 16'd10319, 16'd54977, 16'd34282, 16'd47157, 16'd4650, 16'd5636, 16'd14922, 16'd40943, 16'd23206, 16'd47529, 16'd6295, 16'd4469, 16'd27282, 16'd52867, 16'd22972, 16'd3793, 16'd19189});
	test_expansion(128'h09b3924664a4dd81b2cb50413ccf49fe, {16'd47836, 16'd40843, 16'd1450, 16'd32979, 16'd63344, 16'd32685, 16'd28494, 16'd48471, 16'd34923, 16'd6122, 16'd26814, 16'd49585, 16'd63770, 16'd59861, 16'd57420, 16'd35445, 16'd42527, 16'd25649, 16'd34127, 16'd12054, 16'd12814, 16'd42927, 16'd21333, 16'd8564, 16'd37780, 16'd995});
	test_expansion(128'hb2767f02fc7016f9d2939ab293854f9a, {16'd31945, 16'd26630, 16'd62682, 16'd27106, 16'd35904, 16'd54161, 16'd57789, 16'd33973, 16'd56677, 16'd42477, 16'd59456, 16'd7603, 16'd36107, 16'd13608, 16'd22945, 16'd63809, 16'd61722, 16'd52385, 16'd37859, 16'd57770, 16'd7190, 16'd37583, 16'd11976, 16'd15974, 16'd16845, 16'd27592});
	test_expansion(128'he1ce226460c4af84731f5ce24a4cb070, {16'd40750, 16'd44212, 16'd11849, 16'd6860, 16'd14605, 16'd3047, 16'd54356, 16'd2514, 16'd57006, 16'd27987, 16'd7219, 16'd48450, 16'd32245, 16'd31720, 16'd14751, 16'd24798, 16'd202, 16'd16590, 16'd25159, 16'd48367, 16'd41193, 16'd26220, 16'd2696, 16'd62732, 16'd65233, 16'd20884});
	test_expansion(128'he2ed714571b06e60e6a27427bd6b43dc, {16'd22272, 16'd41747, 16'd42675, 16'd44519, 16'd56662, 16'd7561, 16'd45451, 16'd57476, 16'd56967, 16'd36575, 16'd32032, 16'd33254, 16'd2141, 16'd22247, 16'd12880, 16'd21223, 16'd6599, 16'd35043, 16'd9993, 16'd60140, 16'd28806, 16'd18203, 16'd10384, 16'd28709, 16'd8362, 16'd60559});
	test_expansion(128'hc03be0e7a0058f93f41a2dcad3b6d191, {16'd29573, 16'd38270, 16'd52612, 16'd971, 16'd17256, 16'd62472, 16'd63254, 16'd62073, 16'd29522, 16'd34302, 16'd29632, 16'd34190, 16'd25139, 16'd6463, 16'd28817, 16'd15435, 16'd64921, 16'd2163, 16'd42898, 16'd40835, 16'd22073, 16'd37691, 16'd18008, 16'd26822, 16'd24780, 16'd58113});
	test_expansion(128'h3c476b0805e7281a5f192810e91a0155, {16'd60623, 16'd30270, 16'd45526, 16'd45584, 16'd57176, 16'd18528, 16'd42560, 16'd63333, 16'd51723, 16'd55930, 16'd55940, 16'd22338, 16'd10802, 16'd34344, 16'd27177, 16'd35129, 16'd49112, 16'd57266, 16'd9512, 16'd54763, 16'd15148, 16'd3509, 16'd13188, 16'd60272, 16'd63141, 16'd18504});
	test_expansion(128'hf4b6aee94004d4aa9874529b52ef6f50, {16'd47248, 16'd19707, 16'd10153, 16'd50293, 16'd60885, 16'd43840, 16'd30918, 16'd50499, 16'd47501, 16'd40364, 16'd43464, 16'd65056, 16'd6006, 16'd62038, 16'd51595, 16'd15725, 16'd2833, 16'd28893, 16'd54243, 16'd51954, 16'd62195, 16'd41942, 16'd935, 16'd30058, 16'd19798, 16'd56717});
	test_expansion(128'h7122483359e6e5fa55ba4b815292159c, {16'd17665, 16'd26464, 16'd39730, 16'd10783, 16'd42201, 16'd47461, 16'd12592, 16'd12876, 16'd24008, 16'd60988, 16'd60398, 16'd12268, 16'd57823, 16'd65142, 16'd4400, 16'd8804, 16'd51070, 16'd18399, 16'd3593, 16'd5772, 16'd40656, 16'd61109, 16'd57822, 16'd54154, 16'd40626, 16'd64051});
	test_expansion(128'h9f23c3943392335317d5addb956a03f6, {16'd21004, 16'd9722, 16'd38238, 16'd59874, 16'd13594, 16'd13434, 16'd28617, 16'd35161, 16'd49655, 16'd58472, 16'd65281, 16'd37944, 16'd63766, 16'd30045, 16'd12434, 16'd51333, 16'd63335, 16'd4569, 16'd2744, 16'd420, 16'd48470, 16'd25384, 16'd12160, 16'd43458, 16'd10111, 16'd50800});
	test_expansion(128'h1edcd09f5a946f146ff3cdefbfc83d27, {16'd62364, 16'd42098, 16'd10834, 16'd11381, 16'd32001, 16'd5490, 16'd32130, 16'd26415, 16'd44740, 16'd54422, 16'd1377, 16'd35764, 16'd10661, 16'd47128, 16'd44372, 16'd12500, 16'd35870, 16'd5596, 16'd46236, 16'd9795, 16'd23705, 16'd35512, 16'd55447, 16'd48295, 16'd36915, 16'd39719});
	test_expansion(128'hd39086254678af4e77298cede114eb55, {16'd59410, 16'd23032, 16'd20346, 16'd51016, 16'd6310, 16'd45472, 16'd43129, 16'd47502, 16'd35179, 16'd11651, 16'd32223, 16'd34967, 16'd18780, 16'd49, 16'd45379, 16'd9416, 16'd47259, 16'd54200, 16'd55770, 16'd57878, 16'd64950, 16'd7428, 16'd2407, 16'd37482, 16'd43720, 16'd33206});
	test_expansion(128'h330901664de71a0a829f023f759b867b, {16'd14563, 16'd27685, 16'd23921, 16'd37017, 16'd19029, 16'd29180, 16'd3246, 16'd59125, 16'd1864, 16'd45859, 16'd56763, 16'd5193, 16'd58058, 16'd51123, 16'd51360, 16'd21515, 16'd10818, 16'd56496, 16'd31724, 16'd50515, 16'd59482, 16'd51998, 16'd51392, 16'd12252, 16'd9304, 16'd51917});
	test_expansion(128'h9822cfa632f71f3c46c0619ce9a01279, {16'd53195, 16'd65015, 16'd49875, 16'd13137, 16'd38599, 16'd3102, 16'd19122, 16'd29463, 16'd50860, 16'd21655, 16'd5362, 16'd1189, 16'd7129, 16'd4373, 16'd23926, 16'd6340, 16'd62289, 16'd31749, 16'd32863, 16'd51607, 16'd46756, 16'd30408, 16'd35240, 16'd36946, 16'd14848, 16'd723});
	test_expansion(128'h7858a251c4776ec6d7dc430427bf85b7, {16'd64394, 16'd1656, 16'd54629, 16'd2008, 16'd48973, 16'd5323, 16'd37352, 16'd9091, 16'd31940, 16'd39426, 16'd10959, 16'd64850, 16'd19221, 16'd60801, 16'd12548, 16'd1995, 16'd30111, 16'd62453, 16'd2802, 16'd13249, 16'd25856, 16'd33553, 16'd9917, 16'd37540, 16'd235, 16'd26792});
	test_expansion(128'hf6f310cd727afbc5096aa2e26e3cd5ee, {16'd45251, 16'd26720, 16'd9500, 16'd59136, 16'd51902, 16'd36133, 16'd41817, 16'd34389, 16'd60212, 16'd19211, 16'd3922, 16'd31684, 16'd57367, 16'd14787, 16'd24789, 16'd37994, 16'd47642, 16'd58960, 16'd13765, 16'd41276, 16'd51725, 16'd54665, 16'd19132, 16'd52169, 16'd53578, 16'd23505});
	test_expansion(128'h93d6e7c6a8901c61a6a24e1dedf647d3, {16'd44697, 16'd52902, 16'd18118, 16'd61200, 16'd33873, 16'd39307, 16'd20228, 16'd39290, 16'd20110, 16'd35969, 16'd25378, 16'd16058, 16'd12154, 16'd4751, 16'd31828, 16'd43620, 16'd8044, 16'd17365, 16'd45761, 16'd24821, 16'd26271, 16'd21687, 16'd45860, 16'd46899, 16'd29550, 16'd22787});
	test_expansion(128'hee50d5ac1873ff0fb0697d45187a0a6e, {16'd30089, 16'd49470, 16'd2190, 16'd37736, 16'd43030, 16'd34795, 16'd11614, 16'd8223, 16'd15809, 16'd65392, 16'd23496, 16'd59319, 16'd63219, 16'd15234, 16'd38687, 16'd63137, 16'd546, 16'd12264, 16'd42980, 16'd34328, 16'd39866, 16'd25065, 16'd49384, 16'd59871, 16'd38011, 16'd32176});
	test_expansion(128'h1a46fa9d1734669f434e7d7debf55b19, {16'd32387, 16'd20710, 16'd26938, 16'd10720, 16'd14012, 16'd51061, 16'd50936, 16'd8092, 16'd37525, 16'd42982, 16'd25276, 16'd30189, 16'd3347, 16'd29139, 16'd556, 16'd21070, 16'd8809, 16'd59996, 16'd23638, 16'd62430, 16'd57179, 16'd20658, 16'd64785, 16'd43420, 16'd18722, 16'd6885});
	test_expansion(128'h69abe9222b2841dabb7e43f4ee9f345a, {16'd62781, 16'd41908, 16'd21878, 16'd15885, 16'd21170, 16'd32323, 16'd33233, 16'd37156, 16'd15025, 16'd24313, 16'd61767, 16'd39124, 16'd39040, 16'd51000, 16'd41066, 16'd33784, 16'd45015, 16'd22216, 16'd13814, 16'd15944, 16'd35712, 16'd51618, 16'd1972, 16'd59096, 16'd63872, 16'd29592});
	test_expansion(128'h395011e384af119f939da37f25482410, {16'd12505, 16'd53596, 16'd5878, 16'd22681, 16'd31955, 16'd2246, 16'd27762, 16'd4308, 16'd10051, 16'd11556, 16'd15362, 16'd36191, 16'd2867, 16'd20586, 16'd8244, 16'd23473, 16'd36843, 16'd37583, 16'd13116, 16'd16681, 16'd32611, 16'd31120, 16'd20722, 16'd41714, 16'd39753, 16'd55559});
	test_expansion(128'h4dfcdbbdd753a14fd0e3f1f6ea573f06, {16'd58478, 16'd40375, 16'd48285, 16'd32777, 16'd38719, 16'd57267, 16'd43683, 16'd11045, 16'd8192, 16'd28933, 16'd26411, 16'd40905, 16'd19949, 16'd35983, 16'd64613, 16'd63913, 16'd38000, 16'd36689, 16'd37345, 16'd64955, 16'd42113, 16'd54372, 16'd58836, 16'd64467, 16'd13199, 16'd49212});
	test_expansion(128'hf8ef265f474153ec4aa41e6801537047, {16'd23947, 16'd21033, 16'd4726, 16'd32924, 16'd30665, 16'd38678, 16'd40535, 16'd58277, 16'd64643, 16'd38564, 16'd1048, 16'd3014, 16'd10403, 16'd25248, 16'd18364, 16'd2986, 16'd64536, 16'd19722, 16'd39469, 16'd31898, 16'd40960, 16'd21542, 16'd34636, 16'd57331, 16'd41281, 16'd25078});
	test_expansion(128'had03ca47781b07e2b634724c87ce23e8, {16'd411, 16'd58647, 16'd2742, 16'd62663, 16'd22674, 16'd9491, 16'd59632, 16'd15181, 16'd14435, 16'd30916, 16'd33272, 16'd37665, 16'd32039, 16'd64775, 16'd41743, 16'd8297, 16'd15252, 16'd2484, 16'd35860, 16'd14378, 16'd3055, 16'd61310, 16'd39890, 16'd25380, 16'd45373, 16'd63035});
	test_expansion(128'hde4cadaa35459563ef64f9d8ef44a4a2, {16'd33371, 16'd23781, 16'd19587, 16'd10735, 16'd56269, 16'd18912, 16'd29281, 16'd30098, 16'd38420, 16'd11564, 16'd61628, 16'd48986, 16'd36536, 16'd58605, 16'd10610, 16'd43134, 16'd35459, 16'd60350, 16'd9002, 16'd31015, 16'd7799, 16'd20611, 16'd33847, 16'd24280, 16'd17324, 16'd30458});
	test_expansion(128'h5139556dac9c2ac456b6fdac208e187d, {16'd1856, 16'd52235, 16'd19615, 16'd4018, 16'd2806, 16'd29468, 16'd56107, 16'd49918, 16'd1346, 16'd16394, 16'd1884, 16'd31322, 16'd13519, 16'd54807, 16'd63141, 16'd31803, 16'd19720, 16'd1217, 16'd14455, 16'd58035, 16'd48260, 16'd61598, 16'd52534, 16'd18823, 16'd24685, 16'd25563});
	test_expansion(128'h2c44d466f756a07329c2bf9ebda7cd37, {16'd51305, 16'd982, 16'd29429, 16'd59970, 16'd225, 16'd28318, 16'd1529, 16'd62436, 16'd9165, 16'd29309, 16'd29194, 16'd49539, 16'd9763, 16'd12033, 16'd56493, 16'd36892, 16'd60914, 16'd41964, 16'd15243, 16'd60828, 16'd50472, 16'd13831, 16'd57958, 16'd5801, 16'd27, 16'd16409});
	test_expansion(128'h006d1ac7de7bd8833dac628d32f312d9, {16'd36466, 16'd39389, 16'd14390, 16'd25996, 16'd36691, 16'd59508, 16'd12593, 16'd46766, 16'd1379, 16'd40428, 16'd41148, 16'd46138, 16'd8372, 16'd41569, 16'd23667, 16'd58641, 16'd49530, 16'd56230, 16'd26080, 16'd35909, 16'd31802, 16'd15526, 16'd27413, 16'd27415, 16'd22502, 16'd12269});
	test_expansion(128'h620193dafaeef139caaf1a8add1c1087, {16'd36885, 16'd27816, 16'd3595, 16'd847, 16'd27362, 16'd2921, 16'd61647, 16'd43136, 16'd5893, 16'd63752, 16'd41167, 16'd60204, 16'd21361, 16'd25299, 16'd37821, 16'd65196, 16'd24345, 16'd6959, 16'd55887, 16'd57617, 16'd39867, 16'd65510, 16'd46094, 16'd45450, 16'd48073, 16'd61502});
	test_expansion(128'hac50e906b7e18ccf8157fa8ccd72c879, {16'd64714, 16'd9904, 16'd30834, 16'd3384, 16'd2352, 16'd42376, 16'd12824, 16'd14914, 16'd62196, 16'd8079, 16'd60806, 16'd61478, 16'd42504, 16'd52376, 16'd45113, 16'd62362, 16'd43786, 16'd36567, 16'd47075, 16'd37293, 16'd35763, 16'd9585, 16'd3201, 16'd10684, 16'd65220, 16'd12439});
	test_expansion(128'hc0cc18867ff9140c27eefd36fd2f9960, {16'd880, 16'd51240, 16'd33376, 16'd18857, 16'd23265, 16'd15682, 16'd28062, 16'd60956, 16'd52616, 16'd38902, 16'd21284, 16'd51435, 16'd43758, 16'd9921, 16'd29130, 16'd38389, 16'd29588, 16'd47384, 16'd8770, 16'd24233, 16'd49011, 16'd2790, 16'd8911, 16'd6935, 16'd48948, 16'd43872});
	test_expansion(128'hf862279daad8866c2c40558fadc5a7df, {16'd8333, 16'd8254, 16'd35727, 16'd29227, 16'd64825, 16'd2181, 16'd56837, 16'd34716, 16'd12702, 16'd55076, 16'd33705, 16'd12004, 16'd49820, 16'd3723, 16'd46254, 16'd21788, 16'd35668, 16'd34217, 16'd35701, 16'd52752, 16'd26860, 16'd1250, 16'd39695, 16'd50306, 16'd41329, 16'd1802});
	test_expansion(128'hecb30ef46c30029d6c7c03203b41ce81, {16'd44682, 16'd64090, 16'd43629, 16'd4032, 16'd22157, 16'd8103, 16'd7005, 16'd46589, 16'd35000, 16'd55587, 16'd44354, 16'd12760, 16'd15986, 16'd38620, 16'd38474, 16'd59210, 16'd51617, 16'd5687, 16'd47370, 16'd61597, 16'd48502, 16'd6569, 16'd45884, 16'd41821, 16'd13140, 16'd44846});
	test_expansion(128'h71fb912f01aa5eb8b9f614208ad6a4f6, {16'd24990, 16'd2165, 16'd2328, 16'd29667, 16'd48989, 16'd44822, 16'd34690, 16'd10288, 16'd25074, 16'd43685, 16'd6081, 16'd1505, 16'd39937, 16'd39492, 16'd34648, 16'd54098, 16'd63596, 16'd14441, 16'd39841, 16'd17616, 16'd63915, 16'd27746, 16'd56357, 16'd36657, 16'd21560, 16'd58948});
	test_expansion(128'h825bf19b493a1d5828583c31c0aa1d58, {16'd63163, 16'd64581, 16'd3372, 16'd61092, 16'd44875, 16'd46427, 16'd38523, 16'd2814, 16'd41868, 16'd2570, 16'd63769, 16'd38743, 16'd63614, 16'd49256, 16'd50270, 16'd21026, 16'd2633, 16'd11481, 16'd64507, 16'd14944, 16'd4062, 16'd10398, 16'd3865, 16'd48351, 16'd52946, 16'd30306});
	test_expansion(128'h6458ed5e560947893df219b4157432f3, {16'd27530, 16'd5885, 16'd47715, 16'd26116, 16'd1536, 16'd1128, 16'd2243, 16'd5513, 16'd23481, 16'd39015, 16'd47201, 16'd21524, 16'd53493, 16'd49616, 16'd57460, 16'd39499, 16'd20798, 16'd16857, 16'd7642, 16'd44396, 16'd12356, 16'd43526, 16'd2432, 16'd34967, 16'd4418, 16'd7480});
	test_expansion(128'h2fbaedfb5357708a48505e6ef7454369, {16'd21228, 16'd53787, 16'd44401, 16'd20020, 16'd16483, 16'd63416, 16'd46460, 16'd35912, 16'd23860, 16'd58136, 16'd41794, 16'd5405, 16'd10953, 16'd31494, 16'd61864, 16'd65432, 16'd14841, 16'd32420, 16'd49016, 16'd48952, 16'd15380, 16'd20748, 16'd13159, 16'd27108, 16'd5442, 16'd23200});
	test_expansion(128'h95588091000c630469fa54705c2cac96, {16'd2310, 16'd23528, 16'd63962, 16'd16105, 16'd19111, 16'd35502, 16'd49925, 16'd24820, 16'd37817, 16'd33459, 16'd17232, 16'd21760, 16'd36252, 16'd40770, 16'd31245, 16'd1558, 16'd8444, 16'd45160, 16'd30790, 16'd15911, 16'd42261, 16'd62451, 16'd34126, 16'd60913, 16'd7864, 16'd17019});
	test_expansion(128'hafd70f2e26dd6473ab0259046d983b74, {16'd2312, 16'd26515, 16'd50248, 16'd60417, 16'd32052, 16'd29882, 16'd29872, 16'd59263, 16'd32941, 16'd25126, 16'd383, 16'd25033, 16'd48022, 16'd702, 16'd64447, 16'd35116, 16'd26850, 16'd3839, 16'd63851, 16'd31416, 16'd23883, 16'd65018, 16'd51751, 16'd58071, 16'd13850, 16'd25437});
	test_expansion(128'h4ccec912e6ce15f8bb85b615e3b42ad1, {16'd15718, 16'd50326, 16'd24767, 16'd25587, 16'd5599, 16'd47904, 16'd41776, 16'd40447, 16'd32723, 16'd51657, 16'd8895, 16'd43834, 16'd14883, 16'd3013, 16'd46035, 16'd5356, 16'd36312, 16'd449, 16'd21773, 16'd5826, 16'd10481, 16'd31953, 16'd15942, 16'd33369, 16'd55323, 16'd3906});
	test_expansion(128'h7305edc4419be9bd61b3251f57ca58b6, {16'd1919, 16'd14409, 16'd65391, 16'd36892, 16'd37351, 16'd5076, 16'd19279, 16'd24020, 16'd11662, 16'd12492, 16'd32734, 16'd1069, 16'd9640, 16'd24461, 16'd20017, 16'd7710, 16'd11477, 16'd13061, 16'd32584, 16'd11367, 16'd12509, 16'd50363, 16'd14027, 16'd52727, 16'd35082, 16'd6474});
	test_expansion(128'hb124abed81a96ef5c91700d21874d810, {16'd30089, 16'd50794, 16'd9444, 16'd33565, 16'd32890, 16'd13715, 16'd34806, 16'd52195, 16'd3380, 16'd16201, 16'd44567, 16'd55, 16'd4260, 16'd61576, 16'd46331, 16'd39662, 16'd41920, 16'd60706, 16'd20612, 16'd4770, 16'd1848, 16'd25698, 16'd63015, 16'd25181, 16'd5735, 16'd36358});
	test_expansion(128'h1ed17f9f6a10a288085871e1b5193498, {16'd15449, 16'd6103, 16'd7797, 16'd43397, 16'd65330, 16'd32012, 16'd46095, 16'd55466, 16'd52892, 16'd53864, 16'd16904, 16'd31630, 16'd56830, 16'd20427, 16'd22830, 16'd52166, 16'd55003, 16'd20468, 16'd12000, 16'd919, 16'd62354, 16'd20160, 16'd31214, 16'd1523, 16'd54575, 16'd39676});
	test_expansion(128'ha1d9cbbfd45ad5c567c2738c16dfc628, {16'd58327, 16'd61713, 16'd55162, 16'd14017, 16'd54764, 16'd34272, 16'd63035, 16'd62313, 16'd38837, 16'd11729, 16'd18014, 16'd59377, 16'd2862, 16'd10879, 16'd17248, 16'd26445, 16'd34701, 16'd16790, 16'd51552, 16'd42813, 16'd4105, 16'd61015, 16'd42267, 16'd58710, 16'd42864, 16'd871});
	test_expansion(128'haa5b580de7e917fa98856e55e5adebab, {16'd10212, 16'd40957, 16'd62334, 16'd29402, 16'd60634, 16'd52243, 16'd30559, 16'd24873, 16'd3712, 16'd5857, 16'd8853, 16'd63432, 16'd42601, 16'd57477, 16'd37069, 16'd20252, 16'd49757, 16'd24582, 16'd13974, 16'd31426, 16'd1974, 16'd1324, 16'd25370, 16'd57717, 16'd48499, 16'd53679});
	test_expansion(128'h2e409960df30a8bd8c435e8503b864d2, {16'd35401, 16'd60453, 16'd55443, 16'd5924, 16'd58616, 16'd30398, 16'd54505, 16'd21178, 16'd59606, 16'd53965, 16'd24914, 16'd53226, 16'd65002, 16'd54571, 16'd479, 16'd55765, 16'd6212, 16'd61329, 16'd63557, 16'd41140, 16'd23800, 16'd37047, 16'd7680, 16'd31275, 16'd41412, 16'd45096});
	test_expansion(128'h3f6ccd228b7c97dc7be0f1cd560d0519, {16'd29973, 16'd47132, 16'd9999, 16'd52978, 16'd40423, 16'd58756, 16'd27971, 16'd5052, 16'd19957, 16'd48403, 16'd28338, 16'd10878, 16'd43653, 16'd3150, 16'd7335, 16'd33989, 16'd33369, 16'd64563, 16'd55561, 16'd34267, 16'd14226, 16'd49795, 16'd41886, 16'd37811, 16'd5702, 16'd45451});
	test_expansion(128'h6c4777a486db40f98d5670d0c620b566, {16'd32979, 16'd8446, 16'd8628, 16'd24984, 16'd7853, 16'd16917, 16'd48494, 16'd37436, 16'd58756, 16'd50966, 16'd3722, 16'd21443, 16'd45822, 16'd8992, 16'd29628, 16'd18797, 16'd2925, 16'd3521, 16'd9408, 16'd23033, 16'd23594, 16'd16322, 16'd31270, 16'd28758, 16'd62183, 16'd21761});
	test_expansion(128'h4c7e3568a42b57099ca986672eb8fcd8, {16'd25980, 16'd3118, 16'd3867, 16'd17217, 16'd15920, 16'd18448, 16'd16900, 16'd54679, 16'd15571, 16'd51029, 16'd21297, 16'd1855, 16'd30894, 16'd24154, 16'd47993, 16'd17726, 16'd47810, 16'd30093, 16'd40908, 16'd29119, 16'd60362, 16'd12961, 16'd36061, 16'd22465, 16'd42006, 16'd6829});
	test_expansion(128'h525319440d422a327ec78bcfc590eb79, {16'd24360, 16'd13083, 16'd37816, 16'd51507, 16'd13137, 16'd44760, 16'd24270, 16'd60533, 16'd48495, 16'd4555, 16'd31954, 16'd13444, 16'd35971, 16'd8393, 16'd41075, 16'd45872, 16'd38133, 16'd14851, 16'd44231, 16'd19064, 16'd45812, 16'd20896, 16'd39919, 16'd38726, 16'd13507, 16'd39424});
	test_expansion(128'h5889df355d566face95e67a2820d3050, {16'd16557, 16'd43770, 16'd12247, 16'd52594, 16'd39778, 16'd10031, 16'd12021, 16'd43533, 16'd7662, 16'd42319, 16'd41329, 16'd43082, 16'd30904, 16'd26221, 16'd48204, 16'd49631, 16'd38076, 16'd5748, 16'd9906, 16'd15890, 16'd17350, 16'd53321, 16'd22071, 16'd2756, 16'd50788, 16'd12119});
	test_expansion(128'hd762c22c28ee79bd45b0db02c0ca4089, {16'd14280, 16'd60073, 16'd13559, 16'd35787, 16'd7225, 16'd1885, 16'd54203, 16'd55413, 16'd10962, 16'd15329, 16'd7340, 16'd16029, 16'd43908, 16'd12762, 16'd54728, 16'd54334, 16'd12820, 16'd19806, 16'd51539, 16'd12270, 16'd33229, 16'd62956, 16'd13427, 16'd5360, 16'd62041, 16'd32260});
	test_expansion(128'h9d78e70eac1a641d3b5056cba7ea844e, {16'd22752, 16'd9600, 16'd56413, 16'd52038, 16'd52314, 16'd52382, 16'd41521, 16'd58305, 16'd14631, 16'd61723, 16'd29205, 16'd20563, 16'd46020, 16'd42782, 16'd37822, 16'd65435, 16'd46717, 16'd24462, 16'd25099, 16'd52408, 16'd23032, 16'd4051, 16'd45927, 16'd10292, 16'd38238, 16'd21962});
	test_expansion(128'h85b258dfb9a6944459cfb3c05fe451e4, {16'd23003, 16'd56644, 16'd28327, 16'd42983, 16'd64870, 16'd9861, 16'd61730, 16'd55655, 16'd59364, 16'd22114, 16'd27210, 16'd13824, 16'd39887, 16'd38397, 16'd26301, 16'd46743, 16'd20875, 16'd33626, 16'd25355, 16'd58458, 16'd61573, 16'd9184, 16'd36222, 16'd22428, 16'd2827, 16'd22819});
	test_expansion(128'h835d780cc0b268735bed8f41691cfe0a, {16'd36492, 16'd60102, 16'd39159, 16'd24262, 16'd57741, 16'd65329, 16'd22521, 16'd58873, 16'd23932, 16'd30325, 16'd33268, 16'd6361, 16'd26737, 16'd12671, 16'd7178, 16'd63062, 16'd37413, 16'd60572, 16'd24946, 16'd65037, 16'd55508, 16'd46769, 16'd42900, 16'd57378, 16'd55668, 16'd14169});
	test_expansion(128'h9d95f83d5deec4eb019054e9c586c827, {16'd838, 16'd29911, 16'd41767, 16'd10551, 16'd25953, 16'd26473, 16'd2449, 16'd46418, 16'd42872, 16'd26140, 16'd34531, 16'd25158, 16'd32033, 16'd2061, 16'd20404, 16'd2996, 16'd22510, 16'd14654, 16'd65422, 16'd3691, 16'd28856, 16'd49566, 16'd44876, 16'd42330, 16'd51350, 16'd26487});
	test_expansion(128'h0ff8215bf3aab90b17d8a9caadeb8bbc, {16'd13685, 16'd28242, 16'd6146, 16'd8359, 16'd7466, 16'd32185, 16'd36546, 16'd27469, 16'd1211, 16'd57883, 16'd58332, 16'd62313, 16'd20590, 16'd36134, 16'd61690, 16'd19059, 16'd24283, 16'd52821, 16'd26214, 16'd34315, 16'd11855, 16'd57618, 16'd42412, 16'd32319, 16'd50366, 16'd10138});
	test_expansion(128'h52e2ea50692164f343610fcd427ddff4, {16'd34422, 16'd1145, 16'd42903, 16'd630, 16'd19661, 16'd2902, 16'd54424, 16'd52537, 16'd15104, 16'd55453, 16'd20848, 16'd2776, 16'd22812, 16'd15200, 16'd34714, 16'd38919, 16'd57932, 16'd41094, 16'd5635, 16'd14047, 16'd23689, 16'd22587, 16'd24578, 16'd19201, 16'd13630, 16'd43610});
	test_expansion(128'hb9706a787de607711fa508126ba07dca, {16'd36184, 16'd36224, 16'd1925, 16'd55225, 16'd19572, 16'd32693, 16'd8510, 16'd3476, 16'd53040, 16'd30128, 16'd7326, 16'd39811, 16'd29206, 16'd47789, 16'd60344, 16'd25969, 16'd34930, 16'd38985, 16'd37454, 16'd46885, 16'd2588, 16'd43560, 16'd18583, 16'd7921, 16'd45812, 16'd13407});
	test_expansion(128'h716f4f2cba9e0447b3626dc081dc30b7, {16'd17186, 16'd15668, 16'd26245, 16'd48583, 16'd20629, 16'd59814, 16'd25979, 16'd56177, 16'd23455, 16'd58845, 16'd28990, 16'd30771, 16'd41855, 16'd23485, 16'd21758, 16'd61214, 16'd33575, 16'd15175, 16'd22665, 16'd59073, 16'd30676, 16'd62406, 16'd31216, 16'd51607, 16'd61341, 16'd42702});
	test_expansion(128'h5ae1b27dad17db343a62971f9125b560, {16'd29033, 16'd39620, 16'd53270, 16'd2568, 16'd14970, 16'd15109, 16'd50144, 16'd11371, 16'd42091, 16'd1993, 16'd17848, 16'd3867, 16'd12501, 16'd62994, 16'd43814, 16'd65186, 16'd29619, 16'd54909, 16'd45095, 16'd56382, 16'd51391, 16'd43145, 16'd60506, 16'd20362, 16'd55244, 16'd13270});
	test_expansion(128'h622d0f8459473d36e7dfcd2c6de57d1f, {16'd16335, 16'd37393, 16'd43246, 16'd65532, 16'd59581, 16'd27163, 16'd23203, 16'd8600, 16'd61253, 16'd55923, 16'd28324, 16'd58202, 16'd57387, 16'd42192, 16'd59742, 16'd10788, 16'd47296, 16'd50550, 16'd47977, 16'd51976, 16'd28928, 16'd16477, 16'd35886, 16'd24571, 16'd7390, 16'd61155});
	test_expansion(128'h04b3d32d2c6fec9e8a440b90372a539b, {16'd20839, 16'd52633, 16'd34192, 16'd57729, 16'd52188, 16'd7380, 16'd44442, 16'd28936, 16'd56440, 16'd20372, 16'd42677, 16'd48871, 16'd44829, 16'd40781, 16'd62709, 16'd15385, 16'd55916, 16'd23491, 16'd55435, 16'd20472, 16'd11406, 16'd34089, 16'd61399, 16'd9719, 16'd57695, 16'd25172});
	test_expansion(128'h46d8a92e8b02ddca8727dd13e2639105, {16'd59800, 16'd53706, 16'd10132, 16'd60700, 16'd38684, 16'd3243, 16'd6673, 16'd39402, 16'd55471, 16'd58470, 16'd56074, 16'd50967, 16'd50239, 16'd10225, 16'd5792, 16'd23947, 16'd41517, 16'd53386, 16'd61696, 16'd17725, 16'd36263, 16'd50525, 16'd44451, 16'd51335, 16'd48981, 16'd13580});
	test_expansion(128'hb0dbf8ea15cebe9e769dc078e5f9d669, {16'd61642, 16'd32901, 16'd78, 16'd929, 16'd28910, 16'd42017, 16'd65151, 16'd57830, 16'd32107, 16'd64123, 16'd4628, 16'd45652, 16'd13545, 16'd13660, 16'd4172, 16'd53903, 16'd56053, 16'd3182, 16'd24122, 16'd3948, 16'd31440, 16'd32995, 16'd14397, 16'd15659, 16'd28951, 16'd3705});
	test_expansion(128'h404804b7a0d3d005429b94a48f38fe9a, {16'd64874, 16'd54706, 16'd20131, 16'd62695, 16'd5737, 16'd63625, 16'd50999, 16'd16623, 16'd64634, 16'd1335, 16'd39846, 16'd63008, 16'd27031, 16'd56610, 16'd5176, 16'd11316, 16'd26406, 16'd45488, 16'd46331, 16'd39381, 16'd16697, 16'd62266, 16'd12971, 16'd60026, 16'd49576, 16'd38177});
	test_expansion(128'h9849486b2f21cac1ed193137cb40521e, {16'd33161, 16'd48153, 16'd54888, 16'd2245, 16'd47095, 16'd51253, 16'd58561, 16'd25468, 16'd18671, 16'd22026, 16'd49793, 16'd39397, 16'd33881, 16'd27995, 16'd64637, 16'd24706, 16'd5378, 16'd31756, 16'd3354, 16'd14014, 16'd56313, 16'd36766, 16'd34752, 16'd61953, 16'd7268, 16'd55644});
	test_expansion(128'h825202056e63f0d56a5c88cbaccc2ead, {16'd11464, 16'd64229, 16'd52147, 16'd53153, 16'd10671, 16'd19458, 16'd35359, 16'd46734, 16'd53830, 16'd64774, 16'd3791, 16'd13128, 16'd38325, 16'd39717, 16'd21096, 16'd28040, 16'd56391, 16'd20273, 16'd64710, 16'd50743, 16'd50092, 16'd59736, 16'd29016, 16'd42728, 16'd3597, 16'd41704});
	test_expansion(128'hf854a49473c68e00189f8e895a38e124, {16'd40359, 16'd29026, 16'd19594, 16'd18858, 16'd47350, 16'd48878, 16'd23709, 16'd54514, 16'd39756, 16'd38431, 16'd49903, 16'd28935, 16'd24803, 16'd14725, 16'd54866, 16'd51346, 16'd1612, 16'd54738, 16'd45887, 16'd47806, 16'd25048, 16'd60572, 16'd1346, 16'd13949, 16'd21256, 16'd21562});
	test_expansion(128'h8071395a6e2453c23168ca65d8449ef4, {16'd25766, 16'd47291, 16'd22548, 16'd14752, 16'd52972, 16'd58150, 16'd19085, 16'd101, 16'd28794, 16'd2000, 16'd45000, 16'd11248, 16'd1315, 16'd47900, 16'd9852, 16'd31163, 16'd35942, 16'd28984, 16'd56786, 16'd28938, 16'd57002, 16'd23794, 16'd11848, 16'd11606, 16'd46623, 16'd3968});
	test_expansion(128'h69660d52ff7b1e2352f5e229d4be093a, {16'd21650, 16'd2558, 16'd4722, 16'd54930, 16'd55088, 16'd9679, 16'd34965, 16'd40857, 16'd57090, 16'd2420, 16'd21682, 16'd41591, 16'd43005, 16'd23553, 16'd47106, 16'd62536, 16'd42140, 16'd42197, 16'd48423, 16'd54281, 16'd65412, 16'd27461, 16'd50165, 16'd39717, 16'd27649, 16'd30663});
	test_expansion(128'hcc5e4e3a00fbc7096436eb97b5dd2938, {16'd47254, 16'd18164, 16'd58978, 16'd30576, 16'd23144, 16'd63133, 16'd39354, 16'd16537, 16'd9100, 16'd9048, 16'd16018, 16'd7425, 16'd9543, 16'd42980, 16'd32745, 16'd42410, 16'd58582, 16'd10807, 16'd8683, 16'd37137, 16'd1709, 16'd56662, 16'd25859, 16'd9440, 16'd26765, 16'd7576});
	test_expansion(128'h75397ac6e38cf6c48dd7dcf9e0408702, {16'd13679, 16'd45772, 16'd27620, 16'd7109, 16'd23305, 16'd57213, 16'd54935, 16'd59031, 16'd54380, 16'd16281, 16'd48964, 16'd16650, 16'd48078, 16'd38958, 16'd11616, 16'd21537, 16'd19039, 16'd1517, 16'd3535, 16'd59640, 16'd34930, 16'd50440, 16'd2739, 16'd28549, 16'd38406, 16'd4294});
	test_expansion(128'hc0ae8f11b00f118ea95a4e5bd4d92a6a, {16'd13071, 16'd16381, 16'd51500, 16'd25332, 16'd22467, 16'd25735, 16'd58432, 16'd2318, 16'd18506, 16'd33896, 16'd59829, 16'd34707, 16'd30425, 16'd25178, 16'd31989, 16'd33091, 16'd64081, 16'd17628, 16'd18479, 16'd5566, 16'd62855, 16'd40081, 16'd44839, 16'd55981, 16'd59355, 16'd41437});
	test_expansion(128'h9883a11571c6b15fd34d4a1e04566b51, {16'd48421, 16'd53254, 16'd789, 16'd37930, 16'd44756, 16'd1027, 16'd5075, 16'd7613, 16'd10583, 16'd20054, 16'd28851, 16'd59691, 16'd3767, 16'd31588, 16'd48138, 16'd65065, 16'd33205, 16'd13145, 16'd27657, 16'd37503, 16'd19995, 16'd32923, 16'd33839, 16'd33149, 16'd14758, 16'd20712});
	test_expansion(128'h5688bc2492d4807b7d6fdacd3187a2ea, {16'd58485, 16'd29455, 16'd2236, 16'd16562, 16'd11201, 16'd58283, 16'd6993, 16'd60113, 16'd42741, 16'd11129, 16'd45500, 16'd18846, 16'd34773, 16'd44259, 16'd8731, 16'd18273, 16'd28597, 16'd12746, 16'd36125, 16'd14357, 16'd9531, 16'd23224, 16'd20916, 16'd39182, 16'd24365, 16'd3320});
	test_expansion(128'h79470d99deb6eeb57271e6c67af9a461, {16'd34600, 16'd8770, 16'd62107, 16'd44042, 16'd63152, 16'd42299, 16'd45843, 16'd13406, 16'd31608, 16'd47223, 16'd31093, 16'd55592, 16'd53779, 16'd52591, 16'd64693, 16'd52274, 16'd55051, 16'd24681, 16'd18726, 16'd1533, 16'd54795, 16'd3110, 16'd37764, 16'd61733, 16'd52618, 16'd6427});
	test_expansion(128'h6242bc261ce3bda8c8d371422ccf72b6, {16'd34309, 16'd39885, 16'd36518, 16'd45164, 16'd38579, 16'd15312, 16'd28673, 16'd8315, 16'd16227, 16'd31720, 16'd22364, 16'd8757, 16'd50500, 16'd32684, 16'd23649, 16'd46480, 16'd3095, 16'd51566, 16'd31422, 16'd16078, 16'd58364, 16'd23950, 16'd35688, 16'd37027, 16'd54365, 16'd11522});
	test_expansion(128'h06209c0ff1a2902ecc7740be185f36a0, {16'd30485, 16'd55205, 16'd62671, 16'd22438, 16'd23741, 16'd37841, 16'd58191, 16'd44431, 16'd1943, 16'd29451, 16'd43158, 16'd48820, 16'd53737, 16'd28305, 16'd39151, 16'd13037, 16'd23969, 16'd19298, 16'd37431, 16'd56902, 16'd46453, 16'd65286, 16'd61166, 16'd51359, 16'd25673, 16'd21366});
	test_expansion(128'h99ec0820b6d4fda3a4c1b79e747dd033, {16'd1267, 16'd38006, 16'd28790, 16'd43764, 16'd12246, 16'd10589, 16'd65347, 16'd51762, 16'd61139, 16'd39827, 16'd43532, 16'd54390, 16'd32547, 16'd13540, 16'd51871, 16'd11801, 16'd58793, 16'd44422, 16'd57808, 16'd41469, 16'd42567, 16'd33336, 16'd46235, 16'd60607, 16'd15077, 16'd22998});
	test_expansion(128'h5ff74be5df0d2b2d1cc2744ffc29c52d, {16'd35596, 16'd49925, 16'd21613, 16'd10128, 16'd32915, 16'd25725, 16'd61291, 16'd13223, 16'd19289, 16'd6701, 16'd18106, 16'd2568, 16'd49911, 16'd35401, 16'd64227, 16'd44557, 16'd31508, 16'd36265, 16'd6869, 16'd16345, 16'd7518, 16'd17118, 16'd1182, 16'd65012, 16'd54179, 16'd16303});
	test_expansion(128'hbca054d1e19d31a7145e0e18ddceb4c1, {16'd623, 16'd8291, 16'd23858, 16'd33310, 16'd30999, 16'd5420, 16'd42323, 16'd50510, 16'd16667, 16'd33339, 16'd62127, 16'd21545, 16'd19948, 16'd5062, 16'd7347, 16'd57470, 16'd58750, 16'd17937, 16'd64713, 16'd51633, 16'd7842, 16'd54192, 16'd53209, 16'd54859, 16'd56234, 16'd32199});
	test_expansion(128'h9a6cd24d43f2c8d1e8f30931410adacd, {16'd23541, 16'd60854, 16'd12027, 16'd47815, 16'd46553, 16'd25395, 16'd30347, 16'd1159, 16'd41154, 16'd37176, 16'd58018, 16'd22329, 16'd20100, 16'd39579, 16'd9465, 16'd1056, 16'd33119, 16'd1183, 16'd49910, 16'd50794, 16'd49664, 16'd35988, 16'd26749, 16'd59604, 16'd38770, 16'd6790});
	test_expansion(128'hdd9b9fb652e9924ebf8ae6a308c9a40f, {16'd37699, 16'd51283, 16'd47058, 16'd35817, 16'd28221, 16'd55059, 16'd48983, 16'd22448, 16'd278, 16'd48418, 16'd37421, 16'd31662, 16'd57922, 16'd52155, 16'd42695, 16'd23782, 16'd20995, 16'd44046, 16'd65246, 16'd19430, 16'd57264, 16'd4577, 16'd1646, 16'd61779, 16'd62949, 16'd22451});
	test_expansion(128'h3e263483805f3198ed6b73d86651a0b7, {16'd63691, 16'd64550, 16'd2131, 16'd20919, 16'd9774, 16'd28792, 16'd13284, 16'd61079, 16'd4383, 16'd27295, 16'd55170, 16'd32046, 16'd50385, 16'd42945, 16'd34891, 16'd41448, 16'd47226, 16'd26621, 16'd27528, 16'd48515, 16'd353, 16'd56593, 16'd9807, 16'd8662, 16'd5243, 16'd8499});
	test_expansion(128'hbcc330590a64afd2e292d0196b4ee3c8, {16'd40044, 16'd12541, 16'd62985, 16'd2125, 16'd65071, 16'd49032, 16'd16841, 16'd34015, 16'd13725, 16'd3392, 16'd64962, 16'd5278, 16'd52387, 16'd35427, 16'd14586, 16'd61507, 16'd23762, 16'd59789, 16'd44769, 16'd41102, 16'd4677, 16'd33910, 16'd26312, 16'd10084, 16'd63337, 16'd38218});
	test_expansion(128'h57ad47563ef887ff12f78683a6a6df08, {16'd65238, 16'd27615, 16'd28721, 16'd7996, 16'd40160, 16'd51134, 16'd26261, 16'd5637, 16'd55761, 16'd31228, 16'd29154, 16'd15916, 16'd52586, 16'd1666, 16'd7067, 16'd43510, 16'd16563, 16'd21488, 16'd29568, 16'd36629, 16'd15687, 16'd20402, 16'd62949, 16'd60784, 16'd1451, 16'd11639});
	test_expansion(128'hed78ec0596ea5e23fc81ee18bf831c7b, {16'd18854, 16'd59544, 16'd8164, 16'd46153, 16'd12281, 16'd1433, 16'd44074, 16'd46425, 16'd36143, 16'd32014, 16'd23793, 16'd1759, 16'd10400, 16'd25707, 16'd36552, 16'd25551, 16'd36873, 16'd39217, 16'd64227, 16'd24947, 16'd64340, 16'd51, 16'd43569, 16'd45509, 16'd17116, 16'd54576});
	test_expansion(128'hed2e5b7d05051a8e83ca24e1ac810f8c, {16'd11371, 16'd29932, 16'd40455, 16'd61206, 16'd62750, 16'd9643, 16'd21126, 16'd14380, 16'd24705, 16'd23452, 16'd23062, 16'd49864, 16'd38222, 16'd57417, 16'd15773, 16'd52797, 16'd21877, 16'd10619, 16'd45441, 16'd48764, 16'd63221, 16'd25478, 16'd49546, 16'd21712, 16'd7720, 16'd17231});
	test_expansion(128'h6b75caabd3434751cde1669fe4353d12, {16'd52368, 16'd58069, 16'd53265, 16'd14730, 16'd17236, 16'd14123, 16'd35087, 16'd58454, 16'd32824, 16'd63678, 16'd40564, 16'd38021, 16'd25983, 16'd4644, 16'd51090, 16'd14277, 16'd9323, 16'd59912, 16'd62473, 16'd12074, 16'd22487, 16'd48448, 16'd61597, 16'd51243, 16'd38701, 16'd32144});
	test_expansion(128'h91e5242f770e69446b3202a3a3061401, {16'd18750, 16'd21178, 16'd46464, 16'd22740, 16'd7778, 16'd8712, 16'd7989, 16'd7166, 16'd30181, 16'd42912, 16'd30185, 16'd42857, 16'd6646, 16'd58196, 16'd37678, 16'd7138, 16'd13823, 16'd45703, 16'd62618, 16'd24142, 16'd61794, 16'd33455, 16'd43226, 16'd17373, 16'd63486, 16'd4677});
	test_expansion(128'hfdfc03fe4fd7bd0f5e2b2b677b74acb7, {16'd1710, 16'd51582, 16'd45724, 16'd21988, 16'd10376, 16'd56776, 16'd36479, 16'd18605, 16'd27914, 16'd25703, 16'd1867, 16'd33724, 16'd14574, 16'd26271, 16'd45719, 16'd57274, 16'd49809, 16'd12998, 16'd12544, 16'd35434, 16'd31720, 16'd44148, 16'd56636, 16'd6969, 16'd49612, 16'd25211});
	test_expansion(128'h195125a10f7a1cebaf888339253a04cb, {16'd28982, 16'd48069, 16'd53078, 16'd45819, 16'd54001, 16'd23584, 16'd8507, 16'd12546, 16'd43601, 16'd7060, 16'd43665, 16'd61215, 16'd30741, 16'd17766, 16'd40919, 16'd59357, 16'd23835, 16'd1005, 16'd6687, 16'd41303, 16'd58215, 16'd41998, 16'd14337, 16'd55158, 16'd64095, 16'd49047});
	test_expansion(128'h9e31d0f0a395e0115609b3f74ced3df2, {16'd11910, 16'd55936, 16'd57604, 16'd36148, 16'd44378, 16'd42835, 16'd32226, 16'd26514, 16'd39460, 16'd4795, 16'd42844, 16'd7233, 16'd62687, 16'd56174, 16'd29456, 16'd14726, 16'd17192, 16'd31122, 16'd46520, 16'd23186, 16'd24833, 16'd30234, 16'd27236, 16'd18172, 16'd45418, 16'd14061});
	test_expansion(128'h5dc77336b790a580d1d00ca5df13f9ff, {16'd46210, 16'd10870, 16'd35162, 16'd31193, 16'd33360, 16'd41389, 16'd25814, 16'd36134, 16'd55199, 16'd53477, 16'd41203, 16'd8397, 16'd21371, 16'd30853, 16'd16971, 16'd27592, 16'd60814, 16'd55425, 16'd22181, 16'd41406, 16'd25674, 16'd49986, 16'd47784, 16'd26436, 16'd45108, 16'd14865});
	test_expansion(128'h850bd50095e5293e235d0c991979603d, {16'd20656, 16'd49399, 16'd24064, 16'd45679, 16'd36149, 16'd53192, 16'd7093, 16'd15887, 16'd32723, 16'd23778, 16'd32070, 16'd34521, 16'd6201, 16'd1536, 16'd18214, 16'd35817, 16'd3600, 16'd31942, 16'd53757, 16'd37833, 16'd53701, 16'd10158, 16'd44025, 16'd33126, 16'd60648, 16'd50382});
	test_expansion(128'h291a5a59f3b0dd532730937302ce5291, {16'd39377, 16'd35113, 16'd9262, 16'd37934, 16'd22166, 16'd22163, 16'd44887, 16'd16075, 16'd30667, 16'd64392, 16'd60586, 16'd50628, 16'd2260, 16'd56466, 16'd42599, 16'd27664, 16'd42729, 16'd13007, 16'd48428, 16'd26473, 16'd27361, 16'd33077, 16'd14212, 16'd31701, 16'd36913, 16'd17077});
	test_expansion(128'ha23d9d6037e229fce1d6ad00106e4e63, {16'd13275, 16'd1257, 16'd2598, 16'd5178, 16'd41157, 16'd35573, 16'd52485, 16'd60800, 16'd296, 16'd37254, 16'd470, 16'd4652, 16'd41329, 16'd20330, 16'd24042, 16'd62338, 16'd56391, 16'd51513, 16'd9253, 16'd54429, 16'd44742, 16'd51930, 16'd36079, 16'd15233, 16'd20327, 16'd3620});
	test_expansion(128'h0de17876fdeeae24d329afc7f8df81b9, {16'd52144, 16'd55824, 16'd23097, 16'd38449, 16'd39467, 16'd45210, 16'd54105, 16'd44591, 16'd27421, 16'd61512, 16'd64559, 16'd63919, 16'd2702, 16'd26331, 16'd15777, 16'd23982, 16'd10354, 16'd8005, 16'd24015, 16'd39157, 16'd15716, 16'd60705, 16'd20577, 16'd6763, 16'd45273, 16'd35710});
	test_expansion(128'h8aa9ae6edabfb76f032ec36a96ff5bc9, {16'd49292, 16'd8975, 16'd20046, 16'd12762, 16'd64214, 16'd31416, 16'd27714, 16'd55038, 16'd58928, 16'd18729, 16'd51026, 16'd22299, 16'd32339, 16'd45541, 16'd47280, 16'd8779, 16'd18833, 16'd55624, 16'd11523, 16'd28406, 16'd9441, 16'd27167, 16'd41648, 16'd47665, 16'd10674, 16'd33516});
	test_expansion(128'hc2d4acadb92d1a1fb2f01598d22f68a3, {16'd59273, 16'd16000, 16'd18266, 16'd23136, 16'd65492, 16'd17220, 16'd31303, 16'd49786, 16'd11411, 16'd14737, 16'd37051, 16'd33149, 16'd65388, 16'd52875, 16'd65436, 16'd49471, 16'd27777, 16'd37613, 16'd26162, 16'd51726, 16'd4576, 16'd44825, 16'd52569, 16'd49667, 16'd1428, 16'd56745});
	test_expansion(128'h9dac232ae55138ecf1cc0df3532d6657, {16'd3283, 16'd47662, 16'd41088, 16'd47272, 16'd25164, 16'd13057, 16'd32333, 16'd53372, 16'd57711, 16'd597, 16'd1431, 16'd58218, 16'd50830, 16'd43979, 16'd15564, 16'd44657, 16'd39012, 16'd58919, 16'd38519, 16'd28258, 16'd16833, 16'd36226, 16'd38860, 16'd5434, 16'd57694, 16'd58728});
	test_expansion(128'h7b7e8a90a4b93ca2262f08f4864c65c2, {16'd57402, 16'd35284, 16'd31960, 16'd23783, 16'd20132, 16'd45384, 16'd20236, 16'd18783, 16'd46540, 16'd17264, 16'd28125, 16'd34388, 16'd56980, 16'd36845, 16'd26145, 16'd12058, 16'd44126, 16'd47165, 16'd4116, 16'd35432, 16'd42195, 16'd59563, 16'd3105, 16'd39596, 16'd64949, 16'd8464});
	test_expansion(128'hf9adb4e030bfabc42a6fcb5ae28cbbef, {16'd14961, 16'd29628, 16'd43950, 16'd47585, 16'd35962, 16'd20051, 16'd22496, 16'd9451, 16'd38832, 16'd23706, 16'd60687, 16'd28605, 16'd5921, 16'd38439, 16'd58918, 16'd54803, 16'd23197, 16'd42464, 16'd7698, 16'd58295, 16'd13742, 16'd39051, 16'd16988, 16'd29631, 16'd42407, 16'd53706});
	test_expansion(128'hde0eeb95f37c0d7ccb25e63880b5c06c, {16'd45205, 16'd40595, 16'd47265, 16'd54877, 16'd16435, 16'd49864, 16'd24667, 16'd29317, 16'd24303, 16'd62589, 16'd29097, 16'd8457, 16'd48252, 16'd62116, 16'd55827, 16'd34960, 16'd41013, 16'd65110, 16'd37653, 16'd46430, 16'd7624, 16'd45231, 16'd4730, 16'd14028, 16'd25240, 16'd52234});
	test_expansion(128'he9aa23e792f4bd5b34f030f71eee9ebe, {16'd39107, 16'd64583, 16'd59762, 16'd34697, 16'd43371, 16'd18732, 16'd16227, 16'd25457, 16'd42803, 16'd55948, 16'd48021, 16'd34131, 16'd11149, 16'd11296, 16'd18711, 16'd21727, 16'd21407, 16'd6972, 16'd63478, 16'd25869, 16'd37986, 16'd53718, 16'd64584, 16'd33768, 16'd21566, 16'd36457});
	test_expansion(128'h6d706e8d46e82b69f0f3f4ca1efe3fc0, {16'd35082, 16'd38331, 16'd37785, 16'd33709, 16'd18425, 16'd46254, 16'd45586, 16'd33148, 16'd32526, 16'd46020, 16'd46253, 16'd24271, 16'd10858, 16'd25045, 16'd8444, 16'd39710, 16'd38311, 16'd31254, 16'd17343, 16'd400, 16'd8873, 16'd32635, 16'd65327, 16'd40958, 16'd11775, 16'd34098});
	test_expansion(128'hb606badf1753e97f811118ea8fd67595, {16'd65163, 16'd34689, 16'd51896, 16'd48336, 16'd45470, 16'd58687, 16'd37511, 16'd35997, 16'd31437, 16'd17973, 16'd31133, 16'd33085, 16'd52190, 16'd57432, 16'd10167, 16'd40554, 16'd37004, 16'd55826, 16'd41792, 16'd47684, 16'd38670, 16'd27429, 16'd56174, 16'd46997, 16'd16474, 16'd24272});
	test_expansion(128'h45586b8632bd7db216f92119732f8155, {16'd15264, 16'd62365, 16'd6226, 16'd26848, 16'd25439, 16'd37595, 16'd57712, 16'd25537, 16'd44198, 16'd32836, 16'd30472, 16'd18238, 16'd22308, 16'd29078, 16'd38212, 16'd22472, 16'd5366, 16'd38601, 16'd18571, 16'd46582, 16'd24160, 16'd15955, 16'd48861, 16'd52168, 16'd47994, 16'd46254});
	test_expansion(128'hca8009a07f4468f968cc0cb4140620fc, {16'd44646, 16'd63179, 16'd32286, 16'd35148, 16'd5962, 16'd57691, 16'd41340, 16'd60635, 16'd51094, 16'd7887, 16'd49840, 16'd49727, 16'd57436, 16'd14279, 16'd63274, 16'd32083, 16'd57126, 16'd5657, 16'd55036, 16'd19576, 16'd47655, 16'd19549, 16'd29363, 16'd39688, 16'd6115, 16'd30694});
	test_expansion(128'h48d053f4961fa95d38cc219b3919058c, {16'd41204, 16'd43611, 16'd34992, 16'd21080, 16'd35120, 16'd28083, 16'd8082, 16'd39721, 16'd26509, 16'd37968, 16'd4186, 16'd33648, 16'd56336, 16'd14468, 16'd11392, 16'd42467, 16'd58609, 16'd19687, 16'd51316, 16'd13402, 16'd50564, 16'd43942, 16'd17658, 16'd49336, 16'd9187, 16'd57584});
	test_expansion(128'hbe01e3579836c2d32e5d637fe8e1801b, {16'd57171, 16'd48693, 16'd44151, 16'd4480, 16'd57835, 16'd42500, 16'd51734, 16'd48761, 16'd63116, 16'd23164, 16'd44553, 16'd25596, 16'd27999, 16'd10830, 16'd31592, 16'd17264, 16'd44054, 16'd50520, 16'd15862, 16'd1401, 16'd3064, 16'd11203, 16'd23376, 16'd49173, 16'd17624, 16'd33300});
	test_expansion(128'h64ab824ed252c11a7083e177b2155f86, {16'd11018, 16'd4211, 16'd57432, 16'd54379, 16'd62819, 16'd37908, 16'd52946, 16'd19468, 16'd32156, 16'd23987, 16'd40158, 16'd5402, 16'd55241, 16'd34511, 16'd51109, 16'd20364, 16'd48809, 16'd8353, 16'd35627, 16'd11992, 16'd11212, 16'd55044, 16'd10076, 16'd28676, 16'd13696, 16'd16552});
	test_expansion(128'h71e929c223c4e3826f88b39568f1a50c, {16'd8111, 16'd28357, 16'd10981, 16'd21093, 16'd26922, 16'd25070, 16'd40754, 16'd65147, 16'd58686, 16'd5567, 16'd50210, 16'd64641, 16'd62202, 16'd28838, 16'd43588, 16'd36369, 16'd4912, 16'd51843, 16'd51364, 16'd58544, 16'd3816, 16'd36199, 16'd63725, 16'd14501, 16'd3210, 16'd32883});
	test_expansion(128'h01a7b27b27690bc3c3cc198dbe2e0bd2, {16'd14404, 16'd38183, 16'd146, 16'd60031, 16'd24556, 16'd1626, 16'd3104, 16'd35082, 16'd28116, 16'd51940, 16'd56129, 16'd52727, 16'd19609, 16'd45047, 16'd29988, 16'd22896, 16'd7831, 16'd47132, 16'd32001, 16'd17800, 16'd42559, 16'd19244, 16'd29757, 16'd19448, 16'd28717, 16'd12493});
	test_expansion(128'had7d11fd749115a55c281ad1aad6441f, {16'd31671, 16'd42364, 16'd52122, 16'd59748, 16'd21362, 16'd34868, 16'd30388, 16'd63411, 16'd59399, 16'd2144, 16'd28307, 16'd12175, 16'd55625, 16'd33718, 16'd45151, 16'd27468, 16'd22325, 16'd8768, 16'd7477, 16'd62658, 16'd3154, 16'd46013, 16'd19456, 16'd30215, 16'd62522, 16'd48903});
	test_expansion(128'h7f42f947efc207f08a99023605bbb136, {16'd35609, 16'd29962, 16'd64179, 16'd52697, 16'd50295, 16'd16347, 16'd62937, 16'd9710, 16'd54230, 16'd62306, 16'd60414, 16'd50381, 16'd14915, 16'd12029, 16'd31013, 16'd17047, 16'd27166, 16'd60124, 16'd51287, 16'd20041, 16'd53337, 16'd25820, 16'd5815, 16'd24674, 16'd20417, 16'd21035});
	test_expansion(128'h7f3ff0b82fec4325432b00811e68e2d5, {16'd49614, 16'd14555, 16'd60007, 16'd27510, 16'd51805, 16'd957, 16'd14966, 16'd20347, 16'd60211, 16'd42481, 16'd59962, 16'd37764, 16'd35888, 16'd28726, 16'd52728, 16'd48604, 16'd51572, 16'd56467, 16'd21254, 16'd33603, 16'd55060, 16'd62926, 16'd55141, 16'd47848, 16'd11066, 16'd20101});
	test_expansion(128'h3b0a3bc100a97bbfc72010091e4ac674, {16'd37757, 16'd40826, 16'd7768, 16'd36120, 16'd24904, 16'd39884, 16'd57782, 16'd21969, 16'd55265, 16'd18047, 16'd9607, 16'd21546, 16'd47236, 16'd63653, 16'd8184, 16'd34871, 16'd30438, 16'd3264, 16'd25022, 16'd47922, 16'd47085, 16'd2773, 16'd20572, 16'd6393, 16'd13298, 16'd47363});
	test_expansion(128'h539798c5d429e9781834281498cc2e89, {16'd4345, 16'd20046, 16'd31980, 16'd58362, 16'd30931, 16'd46995, 16'd18986, 16'd49673, 16'd26625, 16'd51366, 16'd16922, 16'd36064, 16'd44651, 16'd28696, 16'd11199, 16'd34420, 16'd22754, 16'd21220, 16'd38034, 16'd43950, 16'd46782, 16'd31985, 16'd2503, 16'd56648, 16'd47054, 16'd1105});
	test_expansion(128'h2eea9fad5350143e0dcb8605960facd0, {16'd52, 16'd25406, 16'd25790, 16'd47281, 16'd44028, 16'd10191, 16'd49311, 16'd1690, 16'd40959, 16'd15961, 16'd4978, 16'd35032, 16'd64194, 16'd46034, 16'd43558, 16'd56429, 16'd55395, 16'd59496, 16'd20170, 16'd51709, 16'd32808, 16'd64780, 16'd32781, 16'd36157, 16'd34044, 16'd14393});
	test_expansion(128'h314a541c667cfa79f18d2e9fc78b976f, {16'd37327, 16'd50052, 16'd44670, 16'd11581, 16'd34796, 16'd5562, 16'd36474, 16'd25974, 16'd50399, 16'd42568, 16'd21954, 16'd33666, 16'd48741, 16'd46503, 16'd47213, 16'd21840, 16'd36959, 16'd54196, 16'd29996, 16'd14335, 16'd2364, 16'd39098, 16'd42638, 16'd35082, 16'd61373, 16'd20430});
	test_expansion(128'hb3eb7211a6de143cb5ede72d76e8f415, {16'd16173, 16'd28012, 16'd1614, 16'd32924, 16'd21464, 16'd51062, 16'd12658, 16'd11148, 16'd42458, 16'd7700, 16'd46498, 16'd18456, 16'd20790, 16'd41763, 16'd46950, 16'd7030, 16'd18514, 16'd6566, 16'd24133, 16'd9712, 16'd46402, 16'd4022, 16'd27078, 16'd54936, 16'd52734, 16'd12830});
	test_expansion(128'h1e90fa7b8ef2a865325350c633c81371, {16'd32687, 16'd54365, 16'd8331, 16'd54365, 16'd51921, 16'd50131, 16'd65067, 16'd64742, 16'd29272, 16'd2957, 16'd31095, 16'd15012, 16'd5702, 16'd33948, 16'd44136, 16'd59680, 16'd46323, 16'd33967, 16'd41900, 16'd32843, 16'd29267, 16'd45969, 16'd35826, 16'd58106, 16'd26854, 16'd33245});
	test_expansion(128'he9aeb08077b9e2c0ab05fb695aaf680f, {16'd50031, 16'd40519, 16'd26479, 16'd64473, 16'd12327, 16'd64974, 16'd50144, 16'd17193, 16'd26214, 16'd35292, 16'd38748, 16'd21092, 16'd14866, 16'd42708, 16'd23187, 16'd2915, 16'd50725, 16'd23064, 16'd26042, 16'd49904, 16'd20225, 16'd18003, 16'd61115, 16'd16707, 16'd64872, 16'd52163});
	test_expansion(128'ha73aa9050efede7c253d8c5f5c7c9ce3, {16'd52987, 16'd64544, 16'd12037, 16'd46170, 16'd41939, 16'd7036, 16'd20958, 16'd50095, 16'd57238, 16'd32750, 16'd36301, 16'd9691, 16'd11473, 16'd38227, 16'd36541, 16'd31608, 16'd61669, 16'd15507, 16'd19122, 16'd23467, 16'd59341, 16'd64804, 16'd40417, 16'd51, 16'd36244, 16'd12897});
	test_expansion(128'hc35dcd233e4b29ae9f72f656033563f1, {16'd41644, 16'd23998, 16'd27490, 16'd9052, 16'd10597, 16'd48431, 16'd49165, 16'd11357, 16'd43835, 16'd53980, 16'd58210, 16'd52787, 16'd50261, 16'd20761, 16'd1762, 16'd38506, 16'd27652, 16'd19722, 16'd56543, 16'd32474, 16'd44977, 16'd22567, 16'd7034, 16'd57640, 16'd9524, 16'd10149});
	test_expansion(128'h4286216c0f540a37e0f09bce35cfe6db, {16'd16990, 16'd51627, 16'd50469, 16'd44165, 16'd13686, 16'd29591, 16'd9172, 16'd43037, 16'd51859, 16'd54507, 16'd30340, 16'd8139, 16'd50803, 16'd30158, 16'd13201, 16'd59546, 16'd52169, 16'd37987, 16'd65527, 16'd40022, 16'd9305, 16'd34740, 16'd9270, 16'd43698, 16'd2954, 16'd65424});
	test_expansion(128'h6be18406f576d78f51400dcd41046049, {16'd63580, 16'd55795, 16'd56132, 16'd45249, 16'd3545, 16'd54064, 16'd28847, 16'd24662, 16'd48012, 16'd14915, 16'd7602, 16'd54033, 16'd55529, 16'd52338, 16'd21445, 16'd64096, 16'd33511, 16'd41981, 16'd42943, 16'd56332, 16'd17064, 16'd49096, 16'd42438, 16'd36042, 16'd48722, 16'd9293});
	test_expansion(128'h7e4bcb738838502e47a78d0fe7d91c4f, {16'd61746, 16'd62761, 16'd50957, 16'd45899, 16'd53680, 16'd2484, 16'd62650, 16'd32435, 16'd62761, 16'd54747, 16'd55009, 16'd15559, 16'd33777, 16'd55731, 16'd12541, 16'd41616, 16'd45297, 16'd55218, 16'd28524, 16'd35571, 16'd28394, 16'd1216, 16'd46506, 16'd4697, 16'd45153, 16'd6193});
	test_expansion(128'hd055738602462acf4dca79db32766a3b, {16'd55367, 16'd42810, 16'd51865, 16'd16208, 16'd29364, 16'd60502, 16'd13643, 16'd32236, 16'd23052, 16'd7237, 16'd27595, 16'd25543, 16'd26474, 16'd54756, 16'd57925, 16'd58572, 16'd20721, 16'd145, 16'd1780, 16'd65385, 16'd51220, 16'd9544, 16'd460, 16'd58842, 16'd14249, 16'd10042});
	test_expansion(128'hd308fd98a9ddd41a358a8dfbeffe4069, {16'd11838, 16'd15621, 16'd37172, 16'd46528, 16'd30758, 16'd33447, 16'd9932, 16'd3159, 16'd57931, 16'd25178, 16'd47766, 16'd42249, 16'd18902, 16'd43383, 16'd60830, 16'd39520, 16'd64924, 16'd15752, 16'd51364, 16'd5910, 16'd20411, 16'd33706, 16'd57468, 16'd62163, 16'd30067, 16'd18138});
	test_expansion(128'h6f4225c9a55fac67d6fb6f8dd9faa739, {16'd10352, 16'd16645, 16'd22161, 16'd32103, 16'd14380, 16'd8221, 16'd12603, 16'd35934, 16'd36121, 16'd55271, 16'd35736, 16'd1463, 16'd25330, 16'd23261, 16'd17519, 16'd51322, 16'd59594, 16'd27234, 16'd11394, 16'd54844, 16'd1679, 16'd37697, 16'd8253, 16'd29302, 16'd1502, 16'd42342});
	test_expansion(128'h4ee4e5cd12aaabc7ff484df96f9377eb, {16'd15136, 16'd3478, 16'd36293, 16'd59313, 16'd46194, 16'd13424, 16'd58463, 16'd16348, 16'd31733, 16'd39709, 16'd55537, 16'd23587, 16'd45739, 16'd43267, 16'd11281, 16'd45384, 16'd49353, 16'd48989, 16'd40153, 16'd15313, 16'd54592, 16'd61305, 16'd8368, 16'd37630, 16'd36215, 16'd7876});
	test_expansion(128'h51fb69cf5553f44c73ecc8681cf0dd6b, {16'd19499, 16'd30431, 16'd2372, 16'd9984, 16'd60402, 16'd20293, 16'd97, 16'd5396, 16'd36305, 16'd10907, 16'd6105, 16'd2513, 16'd20541, 16'd19873, 16'd33091, 16'd7495, 16'd63433, 16'd43081, 16'd583, 16'd23394, 16'd61334, 16'd51763, 16'd18241, 16'd9989, 16'd12146, 16'd28972});
	test_expansion(128'hfb45caedc89cb6c1141499e9c881d686, {16'd12568, 16'd60774, 16'd41103, 16'd50378, 16'd49999, 16'd23462, 16'd26786, 16'd12711, 16'd64865, 16'd14368, 16'd43747, 16'd2518, 16'd40204, 16'd18973, 16'd19099, 16'd51583, 16'd11668, 16'd7830, 16'd37391, 16'd17878, 16'd6273, 16'd10245, 16'd3156, 16'd24851, 16'd52252, 16'd39671});
	test_expansion(128'hd31947c4e1e795f3573bf58de43cabf5, {16'd23325, 16'd56677, 16'd29000, 16'd11804, 16'd53193, 16'd20344, 16'd62666, 16'd2424, 16'd18196, 16'd33528, 16'd30831, 16'd48890, 16'd41865, 16'd43901, 16'd25800, 16'd3300, 16'd19657, 16'd57345, 16'd37216, 16'd56617, 16'd28281, 16'd65060, 16'd11853, 16'd52883, 16'd40111, 16'd8328});
	test_expansion(128'h85a25a71e5cdf13c514fee5ea997c51c, {16'd49714, 16'd52860, 16'd19659, 16'd23598, 16'd32660, 16'd43543, 16'd56372, 16'd17460, 16'd39129, 16'd33996, 16'd26291, 16'd51260, 16'd37283, 16'd46253, 16'd34005, 16'd5492, 16'd59212, 16'd36334, 16'd9779, 16'd40783, 16'd31560, 16'd56489, 16'd7794, 16'd33409, 16'd63098, 16'd62983});
	test_expansion(128'heacc58327281bd1c18173dd01ac0d505, {16'd35099, 16'd17710, 16'd49576, 16'd65396, 16'd32573, 16'd39243, 16'd25345, 16'd23644, 16'd35257, 16'd59814, 16'd45842, 16'd51238, 16'd14967, 16'd17151, 16'd44086, 16'd15322, 16'd58374, 16'd64168, 16'd45464, 16'd56732, 16'd59673, 16'd50091, 16'd63633, 16'd10943, 16'd50692, 16'd34521});
	test_expansion(128'h8290b2a15f8737255d37fce0c7591ed7, {16'd10487, 16'd43237, 16'd58345, 16'd46390, 16'd12387, 16'd8682, 16'd29598, 16'd18176, 16'd26789, 16'd14260, 16'd3660, 16'd4064, 16'd39805, 16'd56050, 16'd2640, 16'd9435, 16'd61699, 16'd53584, 16'd61110, 16'd65225, 16'd59468, 16'd334, 16'd57750, 16'd9401, 16'd40583, 16'd65287});
	test_expansion(128'h9d979f807a1a50826c118044fbb30d14, {16'd32121, 16'd42885, 16'd25962, 16'd16339, 16'd24655, 16'd14781, 16'd13980, 16'd29346, 16'd5464, 16'd43038, 16'd1155, 16'd45222, 16'd50159, 16'd65120, 16'd3740, 16'd28249, 16'd50414, 16'd11698, 16'd18097, 16'd17457, 16'd51127, 16'd18213, 16'd54330, 16'd61390, 16'd57887, 16'd11025});
	test_expansion(128'h88faf91318b0db08e69bc0e98889d92f, {16'd9211, 16'd8876, 16'd28991, 16'd23488, 16'd32200, 16'd9831, 16'd16887, 16'd25610, 16'd40237, 16'd38878, 16'd38607, 16'd41786, 16'd34228, 16'd23015, 16'd62991, 16'd39295, 16'd3530, 16'd20849, 16'd21337, 16'd3987, 16'd38270, 16'd18935, 16'd38565, 16'd5357, 16'd12813, 16'd49000});
	test_expansion(128'h9dba9f7188f138093d57c498a6c3a29c, {16'd32870, 16'd10624, 16'd25210, 16'd48757, 16'd36609, 16'd54940, 16'd10215, 16'd62982, 16'd64948, 16'd45182, 16'd19812, 16'd51500, 16'd2739, 16'd15711, 16'd24589, 16'd24312, 16'd64377, 16'd1546, 16'd10619, 16'd15534, 16'd3776, 16'd64738, 16'd48661, 16'd39201, 16'd24012, 16'd56032});
	test_expansion(128'hd510df3191bcab9a2e6598ccb1879070, {16'd49658, 16'd8649, 16'd29055, 16'd21993, 16'd10448, 16'd43653, 16'd64864, 16'd8909, 16'd12740, 16'd15289, 16'd6726, 16'd6356, 16'd48833, 16'd12314, 16'd53612, 16'd55034, 16'd13578, 16'd61401, 16'd28332, 16'd14111, 16'd10141, 16'd55979, 16'd5179, 16'd48357, 16'd22600, 16'd21583});
	test_expansion(128'h501c93d36a592602f122b539b81fe465, {16'd35917, 16'd11026, 16'd41087, 16'd31000, 16'd62604, 16'd46939, 16'd4972, 16'd29991, 16'd1906, 16'd13518, 16'd11012, 16'd7936, 16'd9041, 16'd31856, 16'd21298, 16'd34329, 16'd39891, 16'd32506, 16'd29506, 16'd13836, 16'd54328, 16'd46082, 16'd9870, 16'd14691, 16'd30293, 16'd63423});
	test_expansion(128'h90cd274015ae21d57c5ef844cc8e3496, {16'd18512, 16'd7971, 16'd23670, 16'd50023, 16'd62994, 16'd56342, 16'd41947, 16'd23049, 16'd56273, 16'd6145, 16'd13461, 16'd30054, 16'd60580, 16'd20657, 16'd37235, 16'd7701, 16'd52501, 16'd16881, 16'd33592, 16'd31989, 16'd44056, 16'd23891, 16'd63961, 16'd59035, 16'd5405, 16'd18180});
	test_expansion(128'h3842b29eebd4b2a931a101bc75f1778c, {16'd40125, 16'd53556, 16'd684, 16'd24899, 16'd38393, 16'd45708, 16'd53240, 16'd49339, 16'd10272, 16'd56800, 16'd29435, 16'd59789, 16'd25795, 16'd12520, 16'd1978, 16'd56825, 16'd42779, 16'd4022, 16'd6869, 16'd14237, 16'd31330, 16'd8604, 16'd56174, 16'd62995, 16'd13414, 16'd35941});
	test_expansion(128'h37d0f5b160ae59684f63c0d4ca45bf9d, {16'd3328, 16'd40586, 16'd29054, 16'd21225, 16'd13979, 16'd16708, 16'd10618, 16'd51331, 16'd4877, 16'd54607, 16'd50025, 16'd50017, 16'd12168, 16'd17873, 16'd38198, 16'd19636, 16'd9547, 16'd57222, 16'd21675, 16'd60752, 16'd29600, 16'd39548, 16'd8783, 16'd3369, 16'd19924, 16'd43181});
	test_expansion(128'h77e6044d00287990a4b230d04c13ffbc, {16'd44560, 16'd26358, 16'd55375, 16'd13335, 16'd64066, 16'd55325, 16'd30981, 16'd28853, 16'd13398, 16'd53514, 16'd15517, 16'd32696, 16'd32269, 16'd63584, 16'd43873, 16'd41971, 16'd57690, 16'd14513, 16'd9554, 16'd26841, 16'd43461, 16'd43946, 16'd49560, 16'd49214, 16'd42682, 16'd55122});
	test_expansion(128'hc99923b2c24d8ea2d675fce89fbcfcca, {16'd57110, 16'd46153, 16'd63, 16'd59913, 16'd5230, 16'd65166, 16'd359, 16'd11041, 16'd1731, 16'd31377, 16'd37161, 16'd29666, 16'd8634, 16'd20012, 16'd43006, 16'd7855, 16'd39827, 16'd33489, 16'd23484, 16'd52791, 16'd60106, 16'd22035, 16'd37207, 16'd17097, 16'd54518, 16'd44951});
	test_expansion(128'h9c71d5b8a4347fc1faea1ff08d51c3e2, {16'd37383, 16'd605, 16'd53998, 16'd60584, 16'd4362, 16'd9218, 16'd24962, 16'd57038, 16'd38941, 16'd29882, 16'd20828, 16'd59256, 16'd1414, 16'd3031, 16'd64998, 16'd60558, 16'd61498, 16'd17688, 16'd23436, 16'd739, 16'd14094, 16'd19545, 16'd62550, 16'd39934, 16'd8087, 16'd47303});
	test_expansion(128'h6dbaccaf946e2321ae7c7fd7809db0a2, {16'd25744, 16'd63271, 16'd2190, 16'd28940, 16'd64248, 16'd23851, 16'd62441, 16'd28361, 16'd62259, 16'd25937, 16'd47220, 16'd41876, 16'd60629, 16'd1092, 16'd53040, 16'd35113, 16'd65167, 16'd32503, 16'd43356, 16'd3061, 16'd37994, 16'd53285, 16'd38008, 16'd48483, 16'd4754, 16'd16427});
	test_expansion(128'h1b7dd9fef420844a5749841365addaf8, {16'd25234, 16'd27205, 16'd3715, 16'd15963, 16'd36107, 16'd37378, 16'd17104, 16'd42324, 16'd39507, 16'd27801, 16'd9193, 16'd13473, 16'd49950, 16'd54797, 16'd22186, 16'd21592, 16'd10520, 16'd41138, 16'd12976, 16'd43014, 16'd14753, 16'd31529, 16'd5728, 16'd30554, 16'd3712, 16'd11726});
	test_expansion(128'h4a4f7a6f36dc951bf4cc5e86d0ae4a3f, {16'd16242, 16'd16225, 16'd24426, 16'd40495, 16'd9607, 16'd54458, 16'd30839, 16'd58286, 16'd62568, 16'd56629, 16'd57183, 16'd5512, 16'd54668, 16'd50746, 16'd57322, 16'd35011, 16'd8940, 16'd11602, 16'd20257, 16'd20789, 16'd27566, 16'd19015, 16'd16247, 16'd20728, 16'd29086, 16'd29684});
	test_expansion(128'h496d6662b79be0ad00c50af642622dc1, {16'd37601, 16'd20415, 16'd62611, 16'd27840, 16'd1707, 16'd19376, 16'd10486, 16'd28401, 16'd7308, 16'd60647, 16'd36708, 16'd26324, 16'd43077, 16'd48589, 16'd12658, 16'd44377, 16'd34089, 16'd28750, 16'd13771, 16'd50318, 16'd9054, 16'd58020, 16'd42107, 16'd59686, 16'd24393, 16'd39910});
	test_expansion(128'hd2947a89d023ba0d67eac6ba1e3e213c, {16'd30556, 16'd12846, 16'd56416, 16'd21110, 16'd53743, 16'd21470, 16'd40536, 16'd52483, 16'd47523, 16'd14383, 16'd52561, 16'd53131, 16'd48140, 16'd16660, 16'd35990, 16'd44910, 16'd30608, 16'd33143, 16'd55538, 16'd32641, 16'd63237, 16'd1325, 16'd5270, 16'd61867, 16'd27486, 16'd3560});
	test_expansion(128'h7ba4915b60fc57c7295d0a54cb0a397b, {16'd59437, 16'd23559, 16'd23937, 16'd9996, 16'd44969, 16'd47031, 16'd7151, 16'd12452, 16'd13005, 16'd1478, 16'd22969, 16'd44312, 16'd16896, 16'd3525, 16'd42339, 16'd58674, 16'd4974, 16'd39248, 16'd29198, 16'd52150, 16'd6652, 16'd41114, 16'd62075, 16'd50861, 16'd15272, 16'd46504});
	test_expansion(128'ha6b0a87e7ccec2045354b1a876667a62, {16'd5067, 16'd35969, 16'd25069, 16'd59706, 16'd30563, 16'd56372, 16'd33199, 16'd45853, 16'd53539, 16'd17674, 16'd44686, 16'd15485, 16'd22404, 16'd34677, 16'd65289, 16'd36547, 16'd62691, 16'd46581, 16'd12064, 16'd10555, 16'd22076, 16'd64579, 16'd2506, 16'd25006, 16'd58673, 16'd37518});
	test_expansion(128'ha4d649c6c4f3a6cbfe6c4177b5496d27, {16'd63441, 16'd42496, 16'd30834, 16'd45586, 16'd32686, 16'd5332, 16'd40716, 16'd25637, 16'd60308, 16'd13608, 16'd2095, 16'd21264, 16'd4721, 16'd27381, 16'd28584, 16'd45926, 16'd23111, 16'd15383, 16'd38391, 16'd37644, 16'd54213, 16'd45487, 16'd55948, 16'd29603, 16'd28371, 16'd649});
	test_expansion(128'h04d533b3252318c54a9da1fda95c93a5, {16'd49903, 16'd5935, 16'd49013, 16'd56296, 16'd27056, 16'd37117, 16'd60013, 16'd16386, 16'd59019, 16'd57386, 16'd15549, 16'd37020, 16'd24481, 16'd53240, 16'd17636, 16'd37230, 16'd37118, 16'd7595, 16'd15817, 16'd31743, 16'd33182, 16'd40736, 16'd15428, 16'd18436, 16'd45211, 16'd10329});
	test_expansion(128'he77842dc268b680001283965b5ed9783, {16'd26120, 16'd58607, 16'd23446, 16'd7012, 16'd50422, 16'd19301, 16'd36109, 16'd55090, 16'd49316, 16'd2665, 16'd52686, 16'd43484, 16'd21042, 16'd37326, 16'd22351, 16'd1924, 16'd9529, 16'd47961, 16'd58579, 16'd16876, 16'd23205, 16'd60855, 16'd43061, 16'd7858, 16'd4626, 16'd5311});
	test_expansion(128'h1bbcc34303d47c1d62d8b2f3ac4f71ef, {16'd1610, 16'd35009, 16'd368, 16'd9356, 16'd58854, 16'd58147, 16'd54727, 16'd50292, 16'd26958, 16'd24937, 16'd52047, 16'd34681, 16'd15747, 16'd28230, 16'd46066, 16'd33116, 16'd31545, 16'd15402, 16'd21243, 16'd30558, 16'd23468, 16'd49069, 16'd60338, 16'd4869, 16'd10050, 16'd24626});
	test_expansion(128'h89d6c08c0b7d825ed43a976c5b30560d, {16'd2084, 16'd11950, 16'd45962, 16'd6863, 16'd31033, 16'd16993, 16'd32207, 16'd2862, 16'd18224, 16'd65141, 16'd29228, 16'd29840, 16'd18923, 16'd32731, 16'd31875, 16'd4946, 16'd7945, 16'd61733, 16'd20711, 16'd19548, 16'd41839, 16'd19308, 16'd53716, 16'd25898, 16'd63049, 16'd31852});
	test_expansion(128'he8513563e9a6ff62548f12f1c2d31333, {16'd1410, 16'd9934, 16'd31825, 16'd57952, 16'd24435, 16'd33140, 16'd32160, 16'd396, 16'd60019, 16'd40269, 16'd61604, 16'd11704, 16'd3917, 16'd2690, 16'd11192, 16'd20923, 16'd36627, 16'd37265, 16'd47629, 16'd22905, 16'd22019, 16'd45590, 16'd2190, 16'd13726, 16'd31788, 16'd15810});
	test_expansion(128'h0b0fcce744d8bd6400f80061e303dc81, {16'd16638, 16'd1847, 16'd31161, 16'd24194, 16'd42512, 16'd52890, 16'd38201, 16'd14828, 16'd9822, 16'd58479, 16'd24418, 16'd15517, 16'd64730, 16'd22733, 16'd52374, 16'd21496, 16'd61718, 16'd38337, 16'd49514, 16'd208, 16'd41222, 16'd4286, 16'd54657, 16'd10973, 16'd17091, 16'd48696});
	test_expansion(128'h6eb6a4bdddaf3cf186b9341704b9df4b, {16'd17171, 16'd38605, 16'd34514, 16'd34641, 16'd18612, 16'd29051, 16'd35275, 16'd57797, 16'd47343, 16'd14932, 16'd5175, 16'd28054, 16'd24194, 16'd11231, 16'd14147, 16'd25500, 16'd10416, 16'd38485, 16'd51218, 16'd57897, 16'd62954, 16'd30644, 16'd41637, 16'd31742, 16'd30141, 16'd43153});
	test_expansion(128'h1eb1b050eefb60b806f8d93b9126ef84, {16'd56425, 16'd25870, 16'd44328, 16'd24406, 16'd26853, 16'd24139, 16'd6046, 16'd29472, 16'd19106, 16'd15931, 16'd50069, 16'd59187, 16'd50297, 16'd54473, 16'd15268, 16'd58094, 16'd8914, 16'd50345, 16'd61221, 16'd50324, 16'd49462, 16'd8270, 16'd8668, 16'd10910, 16'd23629, 16'd58239});
	test_expansion(128'hb7c067c10c3b7c73e14f5a022873478f, {16'd25630, 16'd12909, 16'd50585, 16'd49832, 16'd302, 16'd55869, 16'd50964, 16'd26887, 16'd24578, 16'd39064, 16'd24081, 16'd35061, 16'd40338, 16'd28412, 16'd39998, 16'd7879, 16'd52914, 16'd50284, 16'd32625, 16'd41998, 16'd38796, 16'd9490, 16'd35903, 16'd59559, 16'd61430, 16'd32064});
	test_expansion(128'he4e4ccd5359705db7839d358a1254315, {16'd37284, 16'd19719, 16'd45985, 16'd11050, 16'd115, 16'd54431, 16'd45643, 16'd45689, 16'd42444, 16'd22587, 16'd55347, 16'd15345, 16'd57631, 16'd41678, 16'd45468, 16'd31304, 16'd33434, 16'd62850, 16'd26951, 16'd54579, 16'd41754, 16'd41486, 16'd9894, 16'd41366, 16'd32100, 16'd36862});
	test_expansion(128'hb2975d22e693a9ad14b8f329e9f46082, {16'd2645, 16'd5092, 16'd17877, 16'd39444, 16'd65130, 16'd16135, 16'd45627, 16'd27696, 16'd35368, 16'd37123, 16'd2358, 16'd59261, 16'd3475, 16'd57250, 16'd48779, 16'd26787, 16'd50327, 16'd32032, 16'd38713, 16'd32009, 16'd12216, 16'd63304, 16'd34026, 16'd9738, 16'd50646, 16'd45392});
	test_expansion(128'hd6198804bc126aa640840b9da365a2c5, {16'd6776, 16'd42473, 16'd38091, 16'd53483, 16'd63700, 16'd41480, 16'd10703, 16'd57528, 16'd30569, 16'd57396, 16'd57971, 16'd19070, 16'd40648, 16'd26473, 16'd46971, 16'd33732, 16'd52195, 16'd50605, 16'd33847, 16'd24882, 16'd50432, 16'd24925, 16'd42885, 16'd19547, 16'd24432, 16'd29199});
	test_expansion(128'hc292a727cbf49cdb7fa5b467632a6c23, {16'd28828, 16'd49841, 16'd28161, 16'd5004, 16'd39631, 16'd37885, 16'd44071, 16'd7247, 16'd19497, 16'd11521, 16'd58289, 16'd27804, 16'd58181, 16'd29289, 16'd29968, 16'd300, 16'd34471, 16'd53152, 16'd34514, 16'd1945, 16'd56505, 16'd63486, 16'd39697, 16'd13790, 16'd63284, 16'd27289});
	test_expansion(128'h82876ccac4c68fb1efa67a43f178ba37, {16'd24847, 16'd25299, 16'd6121, 16'd3503, 16'd9742, 16'd12587, 16'd58787, 16'd18849, 16'd49432, 16'd59970, 16'd38590, 16'd11174, 16'd51345, 16'd58824, 16'd5722, 16'd33565, 16'd6375, 16'd45168, 16'd25392, 16'd467, 16'd41121, 16'd58507, 16'd3343, 16'd37610, 16'd9785, 16'd10539});
	test_expansion(128'hc2c2dafd328cd1eb1e0508bca8def22e, {16'd50979, 16'd11907, 16'd931, 16'd65158, 16'd21339, 16'd28336, 16'd25544, 16'd42473, 16'd11093, 16'd43545, 16'd49229, 16'd49995, 16'd29590, 16'd33012, 16'd17133, 16'd59076, 16'd59298, 16'd7024, 16'd10645, 16'd37997, 16'd43944, 16'd57381, 16'd40143, 16'd19144, 16'd40610, 16'd64931});
	test_expansion(128'hb072232f7bebce51c9deec682fbb46f7, {16'd31887, 16'd40829, 16'd24034, 16'd39181, 16'd26862, 16'd3454, 16'd54171, 16'd26966, 16'd52387, 16'd6974, 16'd60257, 16'd54120, 16'd58516, 16'd61619, 16'd31114, 16'd10976, 16'd49519, 16'd36232, 16'd16257, 16'd45587, 16'd205, 16'd46970, 16'd16394, 16'd52415, 16'd33988, 16'd23839});
	test_expansion(128'h62f96dc30d39a7ced17fd5558d907fd1, {16'd22450, 16'd6188, 16'd17270, 16'd17665, 16'd21800, 16'd22556, 16'd26829, 16'd63936, 16'd14196, 16'd19219, 16'd14528, 16'd6410, 16'd21982, 16'd52505, 16'd29426, 16'd10012, 16'd10835, 16'd51051, 16'd22167, 16'd27339, 16'd41320, 16'd36579, 16'd14506, 16'd40168, 16'd15099, 16'd18304});
	test_expansion(128'h48f111385e3a44dc01eb442142c0d0ea, {16'd65280, 16'd8988, 16'd12094, 16'd24171, 16'd7929, 16'd17554, 16'd27396, 16'd20132, 16'd32419, 16'd5575, 16'd26747, 16'd31304, 16'd65319, 16'd34030, 16'd13467, 16'd56724, 16'd18216, 16'd57824, 16'd3505, 16'd4068, 16'd27212, 16'd12329, 16'd23565, 16'd30151, 16'd46731, 16'd8186});
	test_expansion(128'hddb6cd8f74a38f4c31f4b8862de1e3ba, {16'd17143, 16'd7310, 16'd33624, 16'd56919, 16'd14542, 16'd30191, 16'd62454, 16'd40619, 16'd49342, 16'd38872, 16'd40975, 16'd13310, 16'd56258, 16'd22720, 16'd12276, 16'd9704, 16'd43894, 16'd58058, 16'd17789, 16'd56364, 16'd28529, 16'd21273, 16'd49967, 16'd48510, 16'd18501, 16'd50146});
	test_expansion(128'h181bb88bf61d125ca54e0523bd327439, {16'd53956, 16'd2285, 16'd6119, 16'd53060, 16'd55776, 16'd41975, 16'd17615, 16'd18752, 16'd46205, 16'd33580, 16'd27857, 16'd45742, 16'd8213, 16'd30729, 16'd44592, 16'd15086, 16'd9041, 16'd48652, 16'd61580, 16'd26354, 16'd58289, 16'd51592, 16'd59975, 16'd114, 16'd63288, 16'd51697});
	test_expansion(128'hbaad1182ac19a7c1caa69b9c9ef25b72, {16'd27963, 16'd47308, 16'd44346, 16'd42674, 16'd27845, 16'd17166, 16'd15650, 16'd42594, 16'd22310, 16'd32137, 16'd38913, 16'd50311, 16'd48735, 16'd21018, 16'd15686, 16'd35975, 16'd47894, 16'd31620, 16'd56806, 16'd64899, 16'd64571, 16'd19735, 16'd7434, 16'd24929, 16'd4384, 16'd4200});
	test_expansion(128'hd40c94bcef9bf88c682809f004b1e565, {16'd17880, 16'd35641, 16'd2649, 16'd16803, 16'd51414, 16'd6388, 16'd56116, 16'd50931, 16'd42236, 16'd23503, 16'd25767, 16'd23336, 16'd20865, 16'd32475, 16'd8127, 16'd39708, 16'd24335, 16'd59466, 16'd36958, 16'd64881, 16'd59609, 16'd9133, 16'd35501, 16'd47382, 16'd5175, 16'd42547});
	test_expansion(128'h54b9605154992276ab6c8377fb2cc1d9, {16'd8365, 16'd12041, 16'd50616, 16'd56850, 16'd25201, 16'd17017, 16'd42185, 16'd52905, 16'd48761, 16'd28591, 16'd16166, 16'd34177, 16'd40695, 16'd45125, 16'd9816, 16'd50318, 16'd47718, 16'd33039, 16'd22718, 16'd46291, 16'd26520, 16'd47212, 16'd56028, 16'd14143, 16'd22065, 16'd23209});
	test_expansion(128'h4af1de5093be392f199f37f84c03f8df, {16'd38430, 16'd17752, 16'd42771, 16'd43175, 16'd38145, 16'd8424, 16'd15764, 16'd38256, 16'd32082, 16'd28539, 16'd45059, 16'd64237, 16'd65419, 16'd1812, 16'd32154, 16'd25829, 16'd51103, 16'd4758, 16'd9463, 16'd63174, 16'd37758, 16'd25959, 16'd13381, 16'd20909, 16'd52701, 16'd63661});
	test_expansion(128'he0a105e40674b1a358d9a94f3112bba4, {16'd39439, 16'd7436, 16'd19877, 16'd56877, 16'd64766, 16'd49586, 16'd42032, 16'd17465, 16'd55651, 16'd31109, 16'd58125, 16'd25225, 16'd62511, 16'd24162, 16'd3701, 16'd44787, 16'd47441, 16'd785, 16'd28632, 16'd55080, 16'd17154, 16'd61617, 16'd8785, 16'd26080, 16'd28498, 16'd65322});
	test_expansion(128'h678a6339abede9a39ccdefeac4fb071a, {16'd61008, 16'd21086, 16'd5703, 16'd35774, 16'd39321, 16'd11188, 16'd24855, 16'd64860, 16'd17756, 16'd35790, 16'd6144, 16'd31331, 16'd26414, 16'd52352, 16'd55251, 16'd64002, 16'd12140, 16'd9949, 16'd30190, 16'd27251, 16'd59723, 16'd49260, 16'd54924, 16'd42947, 16'd63735, 16'd32673});
	test_expansion(128'hf0f5906358dfe1c55eae8968e821d7f1, {16'd30623, 16'd55789, 16'd17531, 16'd8224, 16'd4756, 16'd6676, 16'd55939, 16'd24183, 16'd45266, 16'd40693, 16'd61918, 16'd40534, 16'd5233, 16'd37377, 16'd31890, 16'd42992, 16'd33655, 16'd19034, 16'd22200, 16'd24742, 16'd49513, 16'd19687, 16'd43848, 16'd38123, 16'd33497, 16'd20063});
	test_expansion(128'h31ed5cac823c3e7a28dd1393f02f7bab, {16'd33528, 16'd5743, 16'd41863, 16'd34502, 16'd28391, 16'd49568, 16'd711, 16'd54580, 16'd55383, 16'd42470, 16'd7956, 16'd26581, 16'd47059, 16'd61428, 16'd18254, 16'd33173, 16'd34741, 16'd54637, 16'd12519, 16'd30764, 16'd18219, 16'd26716, 16'd59942, 16'd45930, 16'd150, 16'd25531});
	test_expansion(128'h05107fd2ed8062ddf1bd54c0fc018c2f, {16'd16212, 16'd25454, 16'd14723, 16'd38852, 16'd54173, 16'd7656, 16'd36573, 16'd22876, 16'd62601, 16'd59524, 16'd22863, 16'd13021, 16'd48791, 16'd50130, 16'd22847, 16'd44213, 16'd56693, 16'd51341, 16'd25727, 16'd7215, 16'd53573, 16'd48544, 16'd4199, 16'd40294, 16'd14573, 16'd37146});
	test_expansion(128'h71348aeba429daa4b879ce08fe26699e, {16'd27223, 16'd56003, 16'd59383, 16'd51693, 16'd39992, 16'd48707, 16'd452, 16'd6551, 16'd27974, 16'd40560, 16'd14733, 16'd25257, 16'd27392, 16'd25872, 16'd55932, 16'd22322, 16'd53423, 16'd24885, 16'd54870, 16'd60650, 16'd30841, 16'd46480, 16'd35623, 16'd21031, 16'd58184, 16'd64316});
	test_expansion(128'h5f3c2993727b52e3ee17f205f515bec6, {16'd21052, 16'd42705, 16'd62320, 16'd15502, 16'd12704, 16'd33538, 16'd23439, 16'd64188, 16'd44960, 16'd25584, 16'd14947, 16'd24731, 16'd23915, 16'd47361, 16'd13935, 16'd24615, 16'd42191, 16'd1471, 16'd46586, 16'd1894, 16'd269, 16'd16434, 16'd29101, 16'd57974, 16'd25896, 16'd625});
	test_expansion(128'h385963a3e3d58028f534894e3eab392f, {16'd59968, 16'd52685, 16'd34018, 16'd31828, 16'd34145, 16'd25659, 16'd4073, 16'd32414, 16'd6602, 16'd6037, 16'd46803, 16'd58542, 16'd10013, 16'd33494, 16'd7170, 16'd181, 16'd58398, 16'd41481, 16'd10073, 16'd6066, 16'd29698, 16'd63693, 16'd25578, 16'd61263, 16'd10157, 16'd15019});
	test_expansion(128'h2f01c5ac32265931019936f38c1b7cd4, {16'd18662, 16'd379, 16'd54785, 16'd51956, 16'd28867, 16'd37336, 16'd50388, 16'd29256, 16'd65130, 16'd41711, 16'd40590, 16'd13062, 16'd61474, 16'd46130, 16'd8074, 16'd8740, 16'd11741, 16'd23813, 16'd23403, 16'd57273, 16'd30799, 16'd15960, 16'd11960, 16'd10055, 16'd16549, 16'd47139});
	test_expansion(128'hc5a4ff5384ccda913d20f65594c9e434, {16'd518, 16'd53497, 16'd51758, 16'd46033, 16'd43517, 16'd41114, 16'd26629, 16'd12271, 16'd50286, 16'd53372, 16'd15211, 16'd27028, 16'd2186, 16'd46632, 16'd40217, 16'd17326, 16'd10423, 16'd1271, 16'd45533, 16'd30895, 16'd38789, 16'd6953, 16'd37224, 16'd37885, 16'd25517, 16'd25828});
	test_expansion(128'h6feb887f6cd9b515a7065af72d3ed824, {16'd22681, 16'd12578, 16'd47746, 16'd47828, 16'd25648, 16'd24987, 16'd4695, 16'd64274, 16'd30931, 16'd43372, 16'd13948, 16'd16471, 16'd15518, 16'd25641, 16'd58298, 16'd24127, 16'd21892, 16'd6760, 16'd10926, 16'd30097, 16'd23493, 16'd28680, 16'd59474, 16'd20902, 16'd52481, 16'd10126});
	test_expansion(128'h71fb3e20c4197b56c5df2d462b910f51, {16'd62072, 16'd20295, 16'd10212, 16'd54862, 16'd21355, 16'd838, 16'd28863, 16'd26721, 16'd29228, 16'd52895, 16'd42231, 16'd46040, 16'd23670, 16'd40916, 16'd20687, 16'd60373, 16'd41918, 16'd17463, 16'd30412, 16'd57194, 16'd29934, 16'd27187, 16'd10809, 16'd13904, 16'd50913, 16'd52148});
	test_expansion(128'hcd8ebbea44d4246e646db6910ab7d1a5, {16'd53632, 16'd64435, 16'd39084, 16'd1059, 16'd55643, 16'd42185, 16'd762, 16'd36237, 16'd30722, 16'd57463, 16'd57041, 16'd14579, 16'd1453, 16'd44549, 16'd56639, 16'd5714, 16'd46895, 16'd5860, 16'd33058, 16'd48509, 16'd4385, 16'd62092, 16'd29875, 16'd22955, 16'd37502, 16'd38879});
	test_expansion(128'h8d47d6d881eac63cc79e6e4b532f1714, {16'd32750, 16'd28811, 16'd56497, 16'd51209, 16'd5984, 16'd36068, 16'd7955, 16'd22372, 16'd3639, 16'd25778, 16'd10915, 16'd7220, 16'd39475, 16'd59136, 16'd42592, 16'd22504, 16'd64948, 16'd3467, 16'd52285, 16'd15642, 16'd59752, 16'd15817, 16'd45858, 16'd48781, 16'd43046, 16'd24047});
	test_expansion(128'h8116f981e8afe9ac7365b7e3995f029f, {16'd1108, 16'd8393, 16'd42490, 16'd39781, 16'd9577, 16'd15878, 16'd56315, 16'd34370, 16'd34745, 16'd51676, 16'd26453, 16'd49152, 16'd29380, 16'd13009, 16'd2059, 16'd25381, 16'd55896, 16'd60776, 16'd30557, 16'd51591, 16'd7431, 16'd53689, 16'd38523, 16'd21753, 16'd55576, 16'd40055});
	test_expansion(128'h9023ee6de3657f6543eae4608a98d456, {16'd6700, 16'd50419, 16'd44820, 16'd24367, 16'd13605, 16'd19228, 16'd59446, 16'd29387, 16'd51507, 16'd55058, 16'd14160, 16'd56946, 16'd38190, 16'd19690, 16'd12349, 16'd10551, 16'd10897, 16'd38968, 16'd22130, 16'd9310, 16'd57920, 16'd23474, 16'd5448, 16'd29094, 16'd61554, 16'd8990});
	test_expansion(128'h895e2dc99b013bb7b568ff17ce17b28e, {16'd29112, 16'd15353, 16'd7580, 16'd13793, 16'd11301, 16'd59553, 16'd18428, 16'd25526, 16'd36504, 16'd2401, 16'd5394, 16'd25630, 16'd13867, 16'd43074, 16'd8295, 16'd6832, 16'd22631, 16'd6836, 16'd10332, 16'd35075, 16'd56931, 16'd41806, 16'd29360, 16'd52234, 16'd16699, 16'd4737});
	test_expansion(128'hb80dc2cf36d90624d7d4b1204f801804, {16'd53073, 16'd1114, 16'd7579, 16'd18826, 16'd58311, 16'd1357, 16'd26700, 16'd45832, 16'd46322, 16'd20918, 16'd37573, 16'd23372, 16'd48205, 16'd26478, 16'd8873, 16'd14542, 16'd26704, 16'd8254, 16'd9644, 16'd43065, 16'd65150, 16'd48192, 16'd58275, 16'd45187, 16'd62763, 16'd47818});
	test_expansion(128'h571e6a0fb392a044817a8417961d7404, {16'd19987, 16'd21614, 16'd38745, 16'd21327, 16'd61158, 16'd6008, 16'd49568, 16'd56988, 16'd19341, 16'd12887, 16'd30610, 16'd31851, 16'd57, 16'd50734, 16'd57276, 16'd56096, 16'd60264, 16'd16181, 16'd15596, 16'd28893, 16'd22741, 16'd36225, 16'd15324, 16'd10496, 16'd20990, 16'd25593});
	test_expansion(128'h986549f8f2b03c60b2c94965b95b3232, {16'd64326, 16'd6737, 16'd33310, 16'd41388, 16'd27488, 16'd51365, 16'd20020, 16'd1804, 16'd20277, 16'd64296, 16'd18343, 16'd28625, 16'd61881, 16'd44341, 16'd13965, 16'd827, 16'd26149, 16'd31508, 16'd57463, 16'd34079, 16'd26441, 16'd44196, 16'd18276, 16'd51369, 16'd42764, 16'd52712});
	test_expansion(128'h5ef0cc77f870d897adeba32dfb49a7c2, {16'd42269, 16'd59146, 16'd50375, 16'd19179, 16'd41472, 16'd601, 16'd23867, 16'd38244, 16'd58022, 16'd14743, 16'd18876, 16'd47022, 16'd33099, 16'd10839, 16'd48785, 16'd43977, 16'd43753, 16'd50951, 16'd18617, 16'd59451, 16'd18016, 16'd30884, 16'd19280, 16'd20381, 16'd20845, 16'd56313});
	test_expansion(128'ha967d650e40b8e0fb97abd1c62e7fa36, {16'd36324, 16'd7739, 16'd31588, 16'd60736, 16'd31957, 16'd1019, 16'd59224, 16'd4507, 16'd9639, 16'd42493, 16'd22863, 16'd33162, 16'd47790, 16'd20787, 16'd3268, 16'd1496, 16'd55434, 16'd35692, 16'd52020, 16'd40490, 16'd12853, 16'd46929, 16'd613, 16'd37688, 16'd14854, 16'd49607});
	test_expansion(128'hcd32bf977bf2f755e3f8c5ed4fd86051, {16'd12687, 16'd12938, 16'd14798, 16'd23639, 16'd57301, 16'd53835, 16'd27110, 16'd42878, 16'd8642, 16'd30053, 16'd58157, 16'd27116, 16'd55893, 16'd9709, 16'd33109, 16'd48327, 16'd17969, 16'd276, 16'd12944, 16'd14254, 16'd54999, 16'd40620, 16'd60535, 16'd27821, 16'd21517, 16'd41514});
	test_expansion(128'hf79e8e82c513286db99b2ad1814e0485, {16'd52518, 16'd33708, 16'd26503, 16'd14286, 16'd65452, 16'd42951, 16'd9138, 16'd37789, 16'd62659, 16'd22650, 16'd11250, 16'd24379, 16'd57997, 16'd3068, 16'd13655, 16'd48026, 16'd51487, 16'd18714, 16'd23592, 16'd41521, 16'd30846, 16'd21282, 16'd49785, 16'd50937, 16'd55114, 16'd5092});
	test_expansion(128'h769cf15c8779e73c50c0c5b0159e8d50, {16'd40991, 16'd8074, 16'd21536, 16'd46268, 16'd52732, 16'd11099, 16'd7810, 16'd45778, 16'd508, 16'd50551, 16'd12599, 16'd40295, 16'd31888, 16'd42351, 16'd19863, 16'd6689, 16'd37360, 16'd20870, 16'd31624, 16'd10400, 16'd1566, 16'd3986, 16'd7725, 16'd41360, 16'd56343, 16'd53920});
	test_expansion(128'heb760e098c1d1e53d60a72ecfcab0600, {16'd47645, 16'd43594, 16'd36709, 16'd2823, 16'd33996, 16'd19955, 16'd32106, 16'd19590, 16'd56827, 16'd41999, 16'd56560, 16'd14520, 16'd36538, 16'd32298, 16'd32491, 16'd16874, 16'd22790, 16'd52099, 16'd22775, 16'd9081, 16'd61074, 16'd60891, 16'd32244, 16'd39162, 16'd46421, 16'd60935});
	test_expansion(128'h5fe4a0e92e6a858439bfa4a2132f5cb7, {16'd39222, 16'd17224, 16'd14018, 16'd54066, 16'd11189, 16'd59435, 16'd3095, 16'd49484, 16'd42164, 16'd56435, 16'd51099, 16'd46237, 16'd59687, 16'd25448, 16'd48164, 16'd53019, 16'd23735, 16'd28104, 16'd28477, 16'd46610, 16'd16790, 16'd36000, 16'd11118, 16'd54800, 16'd3492, 16'd20380});
	test_expansion(128'h53678019f22537d51d69b1e1911c51f5, {16'd53370, 16'd17110, 16'd41262, 16'd40920, 16'd9583, 16'd63121, 16'd2586, 16'd52713, 16'd47414, 16'd62998, 16'd30831, 16'd47090, 16'd38078, 16'd27618, 16'd4883, 16'd35112, 16'd45272, 16'd39354, 16'd32181, 16'd25205, 16'd62212, 16'd57002, 16'd55173, 16'd5662, 16'd7313, 16'd53953});
	test_expansion(128'h777bbf0f6402879dd4db6b241a233e9e, {16'd61611, 16'd40050, 16'd1418, 16'd48386, 16'd14665, 16'd58672, 16'd23584, 16'd31072, 16'd26331, 16'd56602, 16'd64085, 16'd12033, 16'd31105, 16'd22692, 16'd47568, 16'd64848, 16'd35791, 16'd35661, 16'd23506, 16'd49962, 16'd8891, 16'd37926, 16'd33262, 16'd51238, 16'd38246, 16'd17324});
	test_expansion(128'h3fbec085a66a44dbcd8c6deb7f710981, {16'd29900, 16'd4864, 16'd24433, 16'd64322, 16'd23383, 16'd38859, 16'd58960, 16'd48097, 16'd59395, 16'd16906, 16'd47425, 16'd55870, 16'd28751, 16'd23237, 16'd51955, 16'd27510, 16'd6914, 16'd53785, 16'd44858, 16'd61505, 16'd46477, 16'd50103, 16'd3294, 16'd44671, 16'd41531, 16'd62971});
	test_expansion(128'h4d5876a61afe81671afe1c94875d8c00, {16'd6434, 16'd35446, 16'd40414, 16'd4714, 16'd5811, 16'd11561, 16'd61299, 16'd29696, 16'd17056, 16'd47300, 16'd4032, 16'd44036, 16'd45617, 16'd29775, 16'd49270, 16'd48380, 16'd60387, 16'd23296, 16'd20341, 16'd30599, 16'd3817, 16'd47989, 16'd43845, 16'd47457, 16'd50125, 16'd59673});
	test_expansion(128'h6a316a0e96103adc7e58fa4dbbea74b7, {16'd28659, 16'd38953, 16'd30265, 16'd15364, 16'd19003, 16'd28611, 16'd40781, 16'd29390, 16'd57397, 16'd63238, 16'd47269, 16'd65458, 16'd18807, 16'd56851, 16'd7938, 16'd50707, 16'd44335, 16'd29825, 16'd45958, 16'd39194, 16'd31938, 16'd63336, 16'd9815, 16'd25070, 16'd63091, 16'd14565});
	test_expansion(128'h40d37cb5326f26ae95cd469266286a72, {16'd13193, 16'd59294, 16'd24912, 16'd22630, 16'd28755, 16'd8308, 16'd18486, 16'd20282, 16'd42010, 16'd24723, 16'd57868, 16'd48089, 16'd44019, 16'd34950, 16'd25524, 16'd10710, 16'd60133, 16'd4585, 16'd8173, 16'd49904, 16'd19042, 16'd7782, 16'd19189, 16'd16557, 16'd13182, 16'd61761});
	test_expansion(128'h9260e6116a6f9059b6513da92cffb565, {16'd34212, 16'd15533, 16'd20144, 16'd9283, 16'd61374, 16'd39604, 16'd45238, 16'd57558, 16'd14360, 16'd42508, 16'd41206, 16'd6443, 16'd64718, 16'd39569, 16'd12489, 16'd27927, 16'd26165, 16'd19323, 16'd2676, 16'd18318, 16'd27881, 16'd12783, 16'd46293, 16'd44728, 16'd40290, 16'd42872});
	test_expansion(128'haded7d9f03ed157e986d5fd2bef03c40, {16'd17751, 16'd21033, 16'd20505, 16'd5013, 16'd32969, 16'd34125, 16'd36341, 16'd58758, 16'd40135, 16'd47109, 16'd8824, 16'd22783, 16'd43554, 16'd60804, 16'd44266, 16'd40112, 16'd12837, 16'd47649, 16'd31519, 16'd27160, 16'd15954, 16'd62303, 16'd57707, 16'd62572, 16'd27304, 16'd52387});
	test_expansion(128'ha00a900cb2cd4734075de590d432549a, {16'd29182, 16'd10597, 16'd51723, 16'd2279, 16'd38977, 16'd49549, 16'd15934, 16'd37770, 16'd37667, 16'd56536, 16'd12863, 16'd51649, 16'd31977, 16'd60542, 16'd38791, 16'd10381, 16'd54444, 16'd52463, 16'd31090, 16'd49151, 16'd22788, 16'd21863, 16'd45607, 16'd60133, 16'd29227, 16'd41447});
	test_expansion(128'h075107ebbf868d53c9fb517827a56a90, {16'd51239, 16'd62138, 16'd56458, 16'd23950, 16'd30636, 16'd29435, 16'd48360, 16'd40169, 16'd45990, 16'd8446, 16'd38564, 16'd42981, 16'd21316, 16'd30211, 16'd29528, 16'd44916, 16'd21133, 16'd14953, 16'd26221, 16'd45137, 16'd37612, 16'd31625, 16'd5209, 16'd59520, 16'd41611, 16'd49208});
	test_expansion(128'h9a99a1b1b02c013f729c42f5ae2d77f2, {16'd41988, 16'd8372, 16'd4647, 16'd32547, 16'd22570, 16'd38463, 16'd60534, 16'd6553, 16'd29934, 16'd46661, 16'd54814, 16'd39339, 16'd46710, 16'd8074, 16'd61024, 16'd49618, 16'd21053, 16'd42385, 16'd34516, 16'd47238, 16'd42289, 16'd52865, 16'd7427, 16'd60556, 16'd29269, 16'd14814});
	test_expansion(128'h77bb2ac0f8a3598ab5c905d89363a519, {16'd31556, 16'd5550, 16'd40345, 16'd64947, 16'd35899, 16'd27276, 16'd10586, 16'd25493, 16'd7594, 16'd12664, 16'd13287, 16'd53266, 16'd29918, 16'd48117, 16'd54397, 16'd9679, 16'd26279, 16'd1386, 16'd42478, 16'd31964, 16'd55734, 16'd45529, 16'd17760, 16'd18249, 16'd50455, 16'd47473});
	test_expansion(128'h8b71acdcac391ea17a25c3d52d6eae2f, {16'd10341, 16'd1457, 16'd40188, 16'd16738, 16'd32124, 16'd29052, 16'd2048, 16'd23689, 16'd57047, 16'd37877, 16'd59846, 16'd46481, 16'd28061, 16'd45470, 16'd62186, 16'd49265, 16'd42298, 16'd5087, 16'd14939, 16'd55683, 16'd33958, 16'd9885, 16'd41115, 16'd19428, 16'd28222, 16'd59199});
	test_expansion(128'h57ec705c61c3ec65f107e6fe3c99f1b0, {16'd16271, 16'd48895, 16'd54766, 16'd24193, 16'd58703, 16'd29621, 16'd62066, 16'd2971, 16'd42728, 16'd56372, 16'd58539, 16'd44676, 16'd24507, 16'd47656, 16'd15, 16'd49278, 16'd46381, 16'd49179, 16'd18735, 16'd60078, 16'd38064, 16'd44073, 16'd10449, 16'd62721, 16'd42266, 16'd38858});
	test_expansion(128'h29ac84f36e8c5388e4a6f75fbcdb93e5, {16'd16214, 16'd49810, 16'd44575, 16'd15693, 16'd56539, 16'd36913, 16'd33798, 16'd47694, 16'd19211, 16'd47660, 16'd60047, 16'd14989, 16'd30843, 16'd54991, 16'd22134, 16'd56773, 16'd65201, 16'd55035, 16'd56910, 16'd40439, 16'd57715, 16'd23475, 16'd60417, 16'd35668, 16'd54119, 16'd13380});
	test_expansion(128'had049eddd3bb91bc99f799f222d94921, {16'd41405, 16'd32412, 16'd13442, 16'd37962, 16'd13827, 16'd58376, 16'd32357, 16'd26661, 16'd1285, 16'd17398, 16'd30390, 16'd28494, 16'd65334, 16'd47259, 16'd1124, 16'd57734, 16'd42307, 16'd49433, 16'd18017, 16'd14060, 16'd47346, 16'd53486, 16'd61361, 16'd61492, 16'd65310, 16'd4728});
	test_expansion(128'h6a8fb0473cf999567daf1396ce5a40f0, {16'd29130, 16'd53064, 16'd49703, 16'd25333, 16'd3505, 16'd13750, 16'd6097, 16'd10124, 16'd41535, 16'd53900, 16'd53671, 16'd54494, 16'd35098, 16'd20452, 16'd58482, 16'd64744, 16'd28068, 16'd42238, 16'd63436, 16'd31367, 16'd9109, 16'd13820, 16'd9452, 16'd56009, 16'd52915, 16'd2289});
	test_expansion(128'h1fd4d981a94146074e8f6a7a693a9f71, {16'd11455, 16'd29169, 16'd30995, 16'd20411, 16'd16120, 16'd7753, 16'd23270, 16'd59940, 16'd64336, 16'd63830, 16'd41619, 16'd58592, 16'd49540, 16'd973, 16'd34691, 16'd46773, 16'd17873, 16'd8307, 16'd22567, 16'd15629, 16'd26395, 16'd8737, 16'd31327, 16'd17018, 16'd39930, 16'd41616});
	test_expansion(128'h6124e4add67fc848be8b2474773b6825, {16'd10412, 16'd8136, 16'd56218, 16'd9731, 16'd55161, 16'd32522, 16'd45273, 16'd23757, 16'd29036, 16'd11613, 16'd33656, 16'd36051, 16'd23692, 16'd46007, 16'd47292, 16'd40275, 16'd21604, 16'd27564, 16'd42067, 16'd20592, 16'd59777, 16'd55069, 16'd55267, 16'd53770, 16'd22479, 16'd17428});
	test_expansion(128'h64beab39a5100c3adecd7c17ef849d19, {16'd29808, 16'd10774, 16'd62788, 16'd34398, 16'd5277, 16'd4083, 16'd29748, 16'd53301, 16'd61325, 16'd26286, 16'd4446, 16'd59023, 16'd40699, 16'd61299, 16'd16217, 16'd5274, 16'd49346, 16'd49206, 16'd35210, 16'd39672, 16'd51727, 16'd7614, 16'd15060, 16'd231, 16'd39361, 16'd10165});
	test_expansion(128'hc131582685aefb467e63ad519a173600, {16'd7302, 16'd63487, 16'd13825, 16'd7222, 16'd26496, 16'd64177, 16'd18313, 16'd31575, 16'd41468, 16'd10911, 16'd11275, 16'd295, 16'd22257, 16'd48483, 16'd33354, 16'd357, 16'd10906, 16'd40868, 16'd11490, 16'd28944, 16'd11629, 16'd17474, 16'd32042, 16'd58861, 16'd20279, 16'd5831});
	test_expansion(128'hdeec58a42f1266d71caace96ceb2bfe4, {16'd33425, 16'd49278, 16'd23123, 16'd4560, 16'd62345, 16'd46804, 16'd61163, 16'd57844, 16'd15095, 16'd19263, 16'd5148, 16'd42135, 16'd46154, 16'd15566, 16'd42550, 16'd23308, 16'd48437, 16'd366, 16'd44170, 16'd60477, 16'd37182, 16'd63129, 16'd57720, 16'd15226, 16'd30111, 16'd11384});
	test_expansion(128'hdd1175088f602aa5f14fc96e4752a01d, {16'd20434, 16'd51, 16'd41590, 16'd45383, 16'd42471, 16'd51566, 16'd62972, 16'd57710, 16'd64861, 16'd41990, 16'd40765, 16'd35447, 16'd63504, 16'd49259, 16'd26501, 16'd23192, 16'd37373, 16'd49379, 16'd53219, 16'd36821, 16'd46531, 16'd58971, 16'd6025, 16'd60508, 16'd24103, 16'd48981});
	test_expansion(128'h671811b1434087c6a0777d1a138f86e0, {16'd1587, 16'd23452, 16'd35654, 16'd62296, 16'd44368, 16'd54380, 16'd2481, 16'd6909, 16'd29550, 16'd60513, 16'd15562, 16'd7153, 16'd38429, 16'd62032, 16'd65013, 16'd54203, 16'd3617, 16'd51511, 16'd39904, 16'd5730, 16'd27005, 16'd42074, 16'd60718, 16'd63157, 16'd12850, 16'd31742});
	test_expansion(128'h4422741189be4488160027b0d23c5c01, {16'd22041, 16'd41424, 16'd51307, 16'd24383, 16'd25865, 16'd43062, 16'd52340, 16'd23711, 16'd47665, 16'd52192, 16'd31, 16'd42031, 16'd16756, 16'd2480, 16'd40539, 16'd38440, 16'd23126, 16'd65497, 16'd9757, 16'd36744, 16'd12856, 16'd9410, 16'd27474, 16'd20675, 16'd7368, 16'd56074});
	test_expansion(128'he1594832f60249f8b041d7dc556f0e0e, {16'd44734, 16'd21212, 16'd42744, 16'd48505, 16'd6977, 16'd22733, 16'd14806, 16'd16486, 16'd35322, 16'd4740, 16'd65057, 16'd55225, 16'd13396, 16'd26326, 16'd46892, 16'd20827, 16'd4880, 16'd59330, 16'd26337, 16'd11752, 16'd3066, 16'd35752, 16'd21196, 16'd52639, 16'd15631, 16'd41289});
	test_expansion(128'hbc4936a0aa5e0170e84d5431a93bd427, {16'd12245, 16'd35957, 16'd1693, 16'd46220, 16'd12893, 16'd29415, 16'd35012, 16'd30582, 16'd39033, 16'd64021, 16'd40374, 16'd2471, 16'd56049, 16'd43054, 16'd45173, 16'd64334, 16'd19033, 16'd38680, 16'd45446, 16'd9771, 16'd24979, 16'd24288, 16'd33035, 16'd19680, 16'd3526, 16'd27133});
	test_expansion(128'ha3f4555c380340194ffb11c72f22477c, {16'd15134, 16'd11443, 16'd59070, 16'd7312, 16'd31580, 16'd3328, 16'd37703, 16'd13785, 16'd61497, 16'd38634, 16'd26865, 16'd9770, 16'd41958, 16'd45134, 16'd26042, 16'd23298, 16'd27978, 16'd50319, 16'd46961, 16'd52733, 16'd8024, 16'd32558, 16'd47971, 16'd10953, 16'd57185, 16'd33677});
	test_expansion(128'h60e5d204f281f54e9d823897816ee7ef, {16'd63897, 16'd6560, 16'd4923, 16'd53093, 16'd21480, 16'd51327, 16'd9739, 16'd25520, 16'd940, 16'd25240, 16'd41283, 16'd62376, 16'd61493, 16'd16747, 16'd23443, 16'd49941, 16'd9545, 16'd61628, 16'd62123, 16'd17246, 16'd55489, 16'd52334, 16'd2120, 16'd24081, 16'd41338, 16'd6502});
	test_expansion(128'h12b8d00105021f74c772617069a4ae1a, {16'd3716, 16'd51548, 16'd10815, 16'd54687, 16'd4289, 16'd47866, 16'd40538, 16'd21696, 16'd45329, 16'd8009, 16'd39092, 16'd1464, 16'd27511, 16'd14324, 16'd16557, 16'd2395, 16'd64243, 16'd1106, 16'd42578, 16'd12195, 16'd15462, 16'd9030, 16'd5621, 16'd36912, 16'd3515, 16'd32072});
	test_expansion(128'h9f748ceeabdce6b9301ee3243551ab99, {16'd29851, 16'd9510, 16'd13107, 16'd22052, 16'd45753, 16'd18759, 16'd3172, 16'd65379, 16'd8351, 16'd6717, 16'd25822, 16'd40442, 16'd5174, 16'd30618, 16'd777, 16'd28660, 16'd54730, 16'd45868, 16'd19699, 16'd42244, 16'd1283, 16'd41019, 16'd34634, 16'd42320, 16'd48582, 16'd22551});
	test_expansion(128'h522c84bdcd7ebb31731e205ead760412, {16'd57761, 16'd12703, 16'd28041, 16'd33746, 16'd27015, 16'd25661, 16'd31561, 16'd56300, 16'd17122, 16'd44310, 16'd43094, 16'd18708, 16'd35095, 16'd1902, 16'd41795, 16'd18995, 16'd19427, 16'd64859, 16'd48092, 16'd50660, 16'd41443, 16'd50054, 16'd7611, 16'd37888, 16'd32043, 16'd880});
	test_expansion(128'h2e9caa417de765ca4dc879cbecbb8f24, {16'd14028, 16'd24091, 16'd31898, 16'd44301, 16'd31947, 16'd56832, 16'd54945, 16'd22502, 16'd6517, 16'd64116, 16'd533, 16'd44057, 16'd61105, 16'd45744, 16'd2239, 16'd8911, 16'd12306, 16'd39674, 16'd3491, 16'd2598, 16'd32982, 16'd27602, 16'd45132, 16'd56907, 16'd37658, 16'd42977});
	test_expansion(128'h76f216d8ceb12846cedc40d32f883b8d, {16'd49232, 16'd41251, 16'd22209, 16'd49418, 16'd28844, 16'd4393, 16'd7719, 16'd61805, 16'd32642, 16'd64437, 16'd26153, 16'd56933, 16'd44437, 16'd40340, 16'd44516, 16'd51714, 16'd64266, 16'd52931, 16'd558, 16'd37735, 16'd41622, 16'd4222, 16'd19570, 16'd39354, 16'd36221, 16'd8118});
	test_expansion(128'h4f8ac3fa7abd97474f36a73c2608e732, {16'd39085, 16'd40345, 16'd20280, 16'd44460, 16'd1405, 16'd2940, 16'd53822, 16'd2463, 16'd62605, 16'd16185, 16'd10932, 16'd53431, 16'd15436, 16'd33602, 16'd21402, 16'd13050, 16'd39133, 16'd35524, 16'd55147, 16'd14619, 16'd40730, 16'd13709, 16'd2777, 16'd13492, 16'd62991, 16'd30061});
	test_expansion(128'hc48a3976c672cabf001c417330b544c7, {16'd59581, 16'd4700, 16'd30091, 16'd39391, 16'd18498, 16'd8706, 16'd10814, 16'd57549, 16'd11731, 16'd12255, 16'd7437, 16'd2100, 16'd33308, 16'd15199, 16'd49767, 16'd6118, 16'd50435, 16'd26259, 16'd33335, 16'd51819, 16'd37933, 16'd63641, 16'd52933, 16'd3525, 16'd28325, 16'd33858});
	test_expansion(128'h3956fc2c6168cba8a63f6778457841b6, {16'd44651, 16'd19799, 16'd51782, 16'd25353, 16'd59392, 16'd3789, 16'd54424, 16'd21347, 16'd5783, 16'd55013, 16'd59822, 16'd24042, 16'd54913, 16'd60206, 16'd37421, 16'd5259, 16'd8085, 16'd55324, 16'd5727, 16'd13012, 16'd62957, 16'd5640, 16'd6800, 16'd10503, 16'd34659, 16'd53915});
	test_expansion(128'had9b973c3d22be582d16cae730b7458b, {16'd21280, 16'd58970, 16'd22058, 16'd61361, 16'd29135, 16'd52823, 16'd33460, 16'd3843, 16'd22990, 16'd22317, 16'd14883, 16'd56936, 16'd15517, 16'd62962, 16'd4532, 16'd22737, 16'd15927, 16'd15397, 16'd39617, 16'd43519, 16'd2929, 16'd16466, 16'd21198, 16'd63446, 16'd4260, 16'd31317});
	test_expansion(128'hd078b17f7c731028aef4c8187ec73f74, {16'd41328, 16'd28835, 16'd54892, 16'd19654, 16'd6310, 16'd55443, 16'd29755, 16'd7604, 16'd56484, 16'd61082, 16'd1824, 16'd64520, 16'd653, 16'd3222, 16'd3181, 16'd37895, 16'd37024, 16'd22722, 16'd59416, 16'd31893, 16'd34208, 16'd57429, 16'd34153, 16'd57197, 16'd3178, 16'd9599});
	test_expansion(128'h0518caafcd11b488139aba00f95bb68e, {16'd11786, 16'd57756, 16'd34830, 16'd35614, 16'd42425, 16'd15688, 16'd63770, 16'd50363, 16'd3279, 16'd17175, 16'd45491, 16'd58426, 16'd33215, 16'd35642, 16'd46928, 16'd8470, 16'd11301, 16'd42668, 16'd1841, 16'd41703, 16'd6524, 16'd35654, 16'd56031, 16'd46088, 16'd10093, 16'd4216});
	test_expansion(128'he8ec7ee8d249a8f2ad2298029b446343, {16'd30954, 16'd23915, 16'd43013, 16'd35971, 16'd14247, 16'd16144, 16'd70, 16'd31265, 16'd7388, 16'd29752, 16'd1765, 16'd43173, 16'd60411, 16'd451, 16'd7552, 16'd14426, 16'd17056, 16'd58871, 16'd23886, 16'd63216, 16'd17164, 16'd15221, 16'd18964, 16'd32459, 16'd13239, 16'd21412});
	test_expansion(128'h355f593c5bcc6a63480975dbde6bedb2, {16'd60171, 16'd15943, 16'd3904, 16'd42617, 16'd56961, 16'd50933, 16'd65011, 16'd60236, 16'd3254, 16'd43767, 16'd43983, 16'd62103, 16'd61296, 16'd19360, 16'd59730, 16'd699, 16'd58896, 16'd32268, 16'd30292, 16'd47629, 16'd57071, 16'd25871, 16'd53770, 16'd37125, 16'd12689, 16'd25662});
	test_expansion(128'h8085081edc6da1e4a2b8727382aa102f, {16'd61965, 16'd17303, 16'd18309, 16'd41426, 16'd10980, 16'd20899, 16'd7424, 16'd45704, 16'd56570, 16'd44542, 16'd7238, 16'd41905, 16'd29869, 16'd6778, 16'd13630, 16'd40722, 16'd13821, 16'd37509, 16'd31778, 16'd35618, 16'd7545, 16'd37966, 16'd30730, 16'd37257, 16'd22537, 16'd31803});
	test_expansion(128'h986de688439e69480a3ae6eb1b34a373, {16'd47303, 16'd37380, 16'd13282, 16'd40768, 16'd9588, 16'd12859, 16'd4188, 16'd22892, 16'd50853, 16'd36211, 16'd54405, 16'd60317, 16'd48807, 16'd33653, 16'd45412, 16'd35970, 16'd12853, 16'd3642, 16'd39636, 16'd13768, 16'd55407, 16'd11352, 16'd42715, 16'd52615, 16'd39397, 16'd27211});
	test_expansion(128'hecfed50507c110e0895c0ed6f62505e9, {16'd43577, 16'd29661, 16'd26972, 16'd27419, 16'd4486, 16'd64499, 16'd61855, 16'd25268, 16'd58149, 16'd13714, 16'd44506, 16'd18411, 16'd20840, 16'd44076, 16'd45001, 16'd11763, 16'd44128, 16'd42960, 16'd50786, 16'd62916, 16'd4154, 16'd18385, 16'd48071, 16'd16810, 16'd63365, 16'd29313});
	test_expansion(128'hf12118c117f8d8e71535991e44f15711, {16'd39219, 16'd59596, 16'd13507, 16'd21052, 16'd60919, 16'd15753, 16'd58492, 16'd7575, 16'd11064, 16'd55960, 16'd27058, 16'd50493, 16'd57152, 16'd19625, 16'd59387, 16'd50327, 16'd31842, 16'd4305, 16'd19076, 16'd37085, 16'd62941, 16'd64566, 16'd64010, 16'd43008, 16'd24444, 16'd13963});
	test_expansion(128'hcb7511e61f8c3b8fe81fffe90a221e5e, {16'd61024, 16'd18039, 16'd44361, 16'd5087, 16'd29080, 16'd3581, 16'd44393, 16'd43503, 16'd5074, 16'd51321, 16'd46533, 16'd63182, 16'd33631, 16'd47263, 16'd41715, 16'd15933, 16'd17895, 16'd46305, 16'd58428, 16'd4217, 16'd16484, 16'd11301, 16'd39551, 16'd50606, 16'd18302, 16'd20103});
	test_expansion(128'hcf3ccd7aceb2af774f471d17e0cab2c6, {16'd30933, 16'd42613, 16'd21229, 16'd33392, 16'd61183, 16'd29864, 16'd4331, 16'd25906, 16'd17232, 16'd4772, 16'd64656, 16'd8598, 16'd55051, 16'd26124, 16'd49510, 16'd1561, 16'd3473, 16'd34194, 16'd45996, 16'd15608, 16'd42984, 16'd42739, 16'd20097, 16'd24889, 16'd7976, 16'd12836});
	test_expansion(128'h66a8e79fe7943f78dfd9f7b3b593fa1a, {16'd9802, 16'd17609, 16'd10391, 16'd29300, 16'd38991, 16'd46547, 16'd36064, 16'd579, 16'd9653, 16'd10979, 16'd29369, 16'd48133, 16'd25930, 16'd50866, 16'd2167, 16'd41256, 16'd15986, 16'd47375, 16'd49281, 16'd29176, 16'd41087, 16'd14474, 16'd25488, 16'd42748, 16'd61897, 16'd4866});
	test_expansion(128'h41e2e0f046b30426cc323fb878741b6f, {16'd23645, 16'd21796, 16'd6786, 16'd63201, 16'd11738, 16'd15839, 16'd46305, 16'd11175, 16'd24580, 16'd16940, 16'd33255, 16'd14153, 16'd56649, 16'd53460, 16'd57247, 16'd21087, 16'd21809, 16'd64762, 16'd42690, 16'd17613, 16'd45202, 16'd24282, 16'd64608, 16'd2018, 16'd47794, 16'd8780});
	test_expansion(128'h5d1cd7b820a4041d7584b39dd84ed67a, {16'd12755, 16'd19487, 16'd4926, 16'd19492, 16'd32119, 16'd50340, 16'd60395, 16'd51276, 16'd24292, 16'd16503, 16'd17766, 16'd54777, 16'd34466, 16'd61435, 16'd18149, 16'd59169, 16'd64828, 16'd52568, 16'd19346, 16'd4180, 16'd46329, 16'd144, 16'd44211, 16'd44233, 16'd18685, 16'd17501});
	test_expansion(128'hbcd713c7e9c00283e400df4a2669d9a0, {16'd29190, 16'd64701, 16'd2253, 16'd31219, 16'd26887, 16'd2219, 16'd18158, 16'd16545, 16'd2039, 16'd14491, 16'd57127, 16'd7928, 16'd54006, 16'd47824, 16'd41386, 16'd50820, 16'd60713, 16'd61055, 16'd2210, 16'd7100, 16'd53244, 16'd15320, 16'd6096, 16'd30548, 16'd21681, 16'd47517});
	test_expansion(128'h1fd28e630d87da927ebf1bd2d02f769c, {16'd36465, 16'd8478, 16'd29932, 16'd18302, 16'd14044, 16'd26195, 16'd58883, 16'd19649, 16'd47123, 16'd17816, 16'd48493, 16'd20193, 16'd32608, 16'd63037, 16'd18572, 16'd5467, 16'd27254, 16'd9218, 16'd8478, 16'd59827, 16'd15820, 16'd42784, 16'd11243, 16'd51777, 16'd49358, 16'd15502});
	test_expansion(128'h267579c710bf88b4fda5dba4fe64ede3, {16'd16701, 16'd54845, 16'd52979, 16'd18146, 16'd59720, 16'd37477, 16'd57152, 16'd23364, 16'd3634, 16'd25814, 16'd30231, 16'd53508, 16'd18666, 16'd14632, 16'd42352, 16'd54576, 16'd57211, 16'd48597, 16'd45626, 16'd58164, 16'd55903, 16'd40282, 16'd61317, 16'd40124, 16'd21229, 16'd7343});
	test_expansion(128'h5f797e9802680308e02ee8f68b871410, {16'd30553, 16'd18123, 16'd47985, 16'd55888, 16'd37883, 16'd17029, 16'd33639, 16'd50675, 16'd56943, 16'd4577, 16'd5597, 16'd39476, 16'd30459, 16'd13373, 16'd12660, 16'd32615, 16'd1979, 16'd23596, 16'd40088, 16'd34215, 16'd16307, 16'd52128, 16'd32270, 16'd54461, 16'd29668, 16'd11452});
	test_expansion(128'hcb632c761206beaf1f866960ce6876a4, {16'd14640, 16'd5666, 16'd10228, 16'd20017, 16'd32423, 16'd46819, 16'd4731, 16'd37241, 16'd11559, 16'd49656, 16'd5742, 16'd11913, 16'd17808, 16'd21241, 16'd10129, 16'd23310, 16'd3489, 16'd36703, 16'd8265, 16'd56667, 16'd46545, 16'd41563, 16'd19534, 16'd11722, 16'd63836, 16'd43866});
	test_expansion(128'h6edaae79de746d8bfccbeef56049163b, {16'd1105, 16'd46438, 16'd8539, 16'd52414, 16'd292, 16'd42375, 16'd33470, 16'd32194, 16'd52107, 16'd43344, 16'd95, 16'd47286, 16'd41773, 16'd34011, 16'd56477, 16'd62945, 16'd33669, 16'd26319, 16'd35215, 16'd29196, 16'd3855, 16'd47623, 16'd46820, 16'd26300, 16'd4184, 16'd845});
	test_expansion(128'he48bdac739cca4b134ec07636e1b5835, {16'd43805, 16'd65448, 16'd53443, 16'd40309, 16'd20022, 16'd26781, 16'd63938, 16'd7849, 16'd33749, 16'd43966, 16'd53669, 16'd4526, 16'd33579, 16'd42791, 16'd13988, 16'd22611, 16'd44335, 16'd20688, 16'd39948, 16'd14725, 16'd17025, 16'd63075, 16'd64117, 16'd5269, 16'd14629, 16'd9966});
	test_expansion(128'hb6c43fa2b6e71d869b9af01fdcdbd47e, {16'd22885, 16'd26990, 16'd28866, 16'd14063, 16'd51837, 16'd2151, 16'd7731, 16'd7153, 16'd34250, 16'd7642, 16'd48130, 16'd18471, 16'd9727, 16'd49307, 16'd58514, 16'd43739, 16'd22033, 16'd25098, 16'd8649, 16'd50278, 16'd14139, 16'd62310, 16'd40656, 16'd45986, 16'd34738, 16'd47632});
	test_expansion(128'h1c7af46a5f3bc29f9fa6cf2c71a34c43, {16'd61239, 16'd13243, 16'd55266, 16'd18016, 16'd1064, 16'd14374, 16'd56304, 16'd11445, 16'd61150, 16'd3039, 16'd54477, 16'd41000, 16'd52083, 16'd17533, 16'd30058, 16'd32829, 16'd455, 16'd57912, 16'd30873, 16'd43851, 16'd7106, 16'd55903, 16'd58926, 16'd62718, 16'd19247, 16'd16473});
	test_expansion(128'h9c876ef1773369e22d2a63c2d4c47d65, {16'd57046, 16'd15302, 16'd30729, 16'd61498, 16'd8749, 16'd54699, 16'd32965, 16'd41701, 16'd43625, 16'd29712, 16'd40838, 16'd6578, 16'd7181, 16'd34229, 16'd48428, 16'd20623, 16'd42708, 16'd17945, 16'd63218, 16'd50060, 16'd65169, 16'd20885, 16'd12431, 16'd4, 16'd52165, 16'd28663});
	test_expansion(128'h2ce89d79ffbf55d3ced349e364593a97, {16'd38676, 16'd55391, 16'd56228, 16'd65151, 16'd61189, 16'd23246, 16'd41741, 16'd34118, 16'd4049, 16'd50720, 16'd16932, 16'd9271, 16'd58014, 16'd47529, 16'd26230, 16'd48240, 16'd37005, 16'd56573, 16'd3268, 16'd20405, 16'd55602, 16'd25732, 16'd32375, 16'd8066, 16'd47424, 16'd47890});
	test_expansion(128'h04a2a4c0fab8049e472eaccdd44b3948, {16'd55782, 16'd31627, 16'd59995, 16'd29176, 16'd39409, 16'd16513, 16'd63048, 16'd47736, 16'd47628, 16'd34579, 16'd3460, 16'd49804, 16'd22479, 16'd58020, 16'd36590, 16'd10149, 16'd22779, 16'd47236, 16'd29936, 16'd59076, 16'd39934, 16'd52347, 16'd43335, 16'd5199, 16'd30611, 16'd23152});
	test_expansion(128'h8ccd29b4c152e357a38913a471f4f70e, {16'd56610, 16'd10275, 16'd51962, 16'd53618, 16'd6204, 16'd50492, 16'd59157, 16'd41789, 16'd47312, 16'd22536, 16'd37951, 16'd32528, 16'd43998, 16'd4347, 16'd1789, 16'd3997, 16'd29030, 16'd2542, 16'd23420, 16'd62708, 16'd58101, 16'd15716, 16'd26164, 16'd28047, 16'd44072, 16'd28573});
	test_expansion(128'hfc067b78087e203587b20eae9862dcfb, {16'd46663, 16'd23416, 16'd60972, 16'd5101, 16'd23167, 16'd32733, 16'd44191, 16'd6509, 16'd47763, 16'd32959, 16'd18716, 16'd10925, 16'd3865, 16'd40984, 16'd465, 16'd14612, 16'd63700, 16'd15320, 16'd11794, 16'd40807, 16'd47224, 16'd64895, 16'd21173, 16'd27315, 16'd39276, 16'd8266});
	test_expansion(128'h538c1d73f2848290b39bd202b7753d07, {16'd46216, 16'd31999, 16'd37587, 16'd6886, 16'd8046, 16'd27092, 16'd26399, 16'd265, 16'd57139, 16'd63488, 16'd40364, 16'd14876, 16'd50675, 16'd65504, 16'd33775, 16'd58536, 16'd17235, 16'd35092, 16'd554, 16'd9630, 16'd49877, 16'd3246, 16'd49855, 16'd25616, 16'd52092, 16'd44435});
	test_expansion(128'hbcc45e102c72f4e3fff0b9ee3d52e25a, {16'd2134, 16'd39064, 16'd40904, 16'd34928, 16'd32868, 16'd37950, 16'd22632, 16'd21573, 16'd15242, 16'd48245, 16'd49810, 16'd5454, 16'd25992, 16'd44856, 16'd11451, 16'd25280, 16'd40510, 16'd36158, 16'd16857, 16'd12804, 16'd25463, 16'd21832, 16'd32061, 16'd8480, 16'd44658, 16'd55674});
	test_expansion(128'h88e049a31edf40121d5a44d140974553, {16'd20902, 16'd12847, 16'd50616, 16'd17819, 16'd5147, 16'd25720, 16'd11221, 16'd7637, 16'd53322, 16'd28690, 16'd12418, 16'd32335, 16'd28445, 16'd33108, 16'd1495, 16'd60025, 16'd1096, 16'd7056, 16'd21972, 16'd60375, 16'd34248, 16'd63950, 16'd30900, 16'd39639, 16'd9783, 16'd47782});
	test_expansion(128'h5d86f582c7d9d03b35aeded1f909d9d6, {16'd23677, 16'd26052, 16'd42479, 16'd35369, 16'd35211, 16'd17492, 16'd50759, 16'd38302, 16'd13210, 16'd14944, 16'd46650, 16'd1276, 16'd52576, 16'd41166, 16'd47704, 16'd56053, 16'd18377, 16'd39462, 16'd36466, 16'd39259, 16'd29665, 16'd43256, 16'd23754, 16'd58050, 16'd29354, 16'd31834});
	test_expansion(128'h1772dd42ce6978e7cfd1cfca3cc7a61c, {16'd7366, 16'd43585, 16'd3465, 16'd55179, 16'd32122, 16'd42525, 16'd36149, 16'd57394, 16'd2579, 16'd41918, 16'd27207, 16'd64582, 16'd64888, 16'd25332, 16'd19293, 16'd63334, 16'd50315, 16'd5140, 16'd29859, 16'd47976, 16'd3406, 16'd24365, 16'd19093, 16'd62559, 16'd41949, 16'd63630});
	test_expansion(128'ha688b2ee913e1c9c23695edbdc1a1b33, {16'd36976, 16'd56662, 16'd20263, 16'd5022, 16'd62403, 16'd12706, 16'd57909, 16'd50374, 16'd2479, 16'd54136, 16'd19413, 16'd43642, 16'd3236, 16'd3941, 16'd62548, 16'd31591, 16'd4842, 16'd33288, 16'd54073, 16'd15668, 16'd17558, 16'd10920, 16'd50623, 16'd9085, 16'd64748, 16'd7286});
	test_expansion(128'hc1b11ee3c187603a0dc88ed10c62962e, {16'd48005, 16'd27130, 16'd11469, 16'd46828, 16'd34190, 16'd31097, 16'd18232, 16'd60150, 16'd61891, 16'd45368, 16'd4684, 16'd4869, 16'd27037, 16'd55322, 16'd8501, 16'd3622, 16'd47343, 16'd14272, 16'd64330, 16'd41617, 16'd55804, 16'd17907, 16'd6601, 16'd8499, 16'd5286, 16'd6135});
	test_expansion(128'h7ec275324c63d5f607a8bd5b4d9bdd09, {16'd42793, 16'd38079, 16'd44825, 16'd32177, 16'd2073, 16'd64678, 16'd44272, 16'd53582, 16'd10701, 16'd37308, 16'd44594, 16'd32150, 16'd63078, 16'd4146, 16'd40703, 16'd30586, 16'd43019, 16'd32304, 16'd55957, 16'd35827, 16'd5316, 16'd56699, 16'd6591, 16'd24455, 16'd32209, 16'd37530});
	test_expansion(128'hfe0dcfea821861d5bb6336493f7f2bb0, {16'd34288, 16'd62565, 16'd45914, 16'd60717, 16'd31700, 16'd52409, 16'd39116, 16'd32719, 16'd19482, 16'd51532, 16'd8594, 16'd45483, 16'd13409, 16'd18103, 16'd49104, 16'd34069, 16'd22895, 16'd34399, 16'd10011, 16'd62323, 16'd50564, 16'd39222, 16'd9237, 16'd56510, 16'd3610, 16'd38856});
	test_expansion(128'h19115142413778f9cff6d82bf7e90f5c, {16'd40627, 16'd30124, 16'd17413, 16'd57341, 16'd15062, 16'd29574, 16'd4295, 16'd13602, 16'd15798, 16'd27150, 16'd52977, 16'd54933, 16'd47568, 16'd8333, 16'd31004, 16'd33116, 16'd756, 16'd25018, 16'd41884, 16'd6064, 16'd41210, 16'd23643, 16'd45833, 16'd33271, 16'd23946, 16'd33452});
	test_expansion(128'h37f2c87d2922362da159a0ce17c85ee6, {16'd62827, 16'd17491, 16'd9583, 16'd22974, 16'd35351, 16'd5835, 16'd7704, 16'd24231, 16'd40888, 16'd17294, 16'd56230, 16'd26946, 16'd14953, 16'd15735, 16'd37671, 16'd14598, 16'd8660, 16'd10212, 16'd17669, 16'd50447, 16'd29660, 16'd9257, 16'd31054, 16'd7415, 16'd11958, 16'd44606});
	test_expansion(128'h44ff21789c850129934bfc777b769d1b, {16'd16658, 16'd52217, 16'd3315, 16'd61337, 16'd52122, 16'd48638, 16'd3584, 16'd30315, 16'd59328, 16'd34015, 16'd62752, 16'd55196, 16'd50206, 16'd11094, 16'd63345, 16'd65234, 16'd38509, 16'd1608, 16'd8378, 16'd26333, 16'd42057, 16'd18702, 16'd48019, 16'd1478, 16'd26012, 16'd14133});
	test_expansion(128'h47790abc9bab83a8277609eee4704949, {16'd29225, 16'd56866, 16'd36745, 16'd20606, 16'd1258, 16'd4054, 16'd58815, 16'd20523, 16'd27010, 16'd56307, 16'd39661, 16'd60890, 16'd51367, 16'd9711, 16'd45852, 16'd45921, 16'd62624, 16'd32519, 16'd39657, 16'd32264, 16'd4221, 16'd1448, 16'd60218, 16'd8859, 16'd51417, 16'd23757});
	test_expansion(128'h34f22319a1967421a2ed0839ed187e05, {16'd485, 16'd6673, 16'd48824, 16'd31941, 16'd51079, 16'd12475, 16'd24367, 16'd60365, 16'd43261, 16'd57307, 16'd8399, 16'd32135, 16'd3708, 16'd59106, 16'd13237, 16'd60729, 16'd43639, 16'd32349, 16'd3293, 16'd22385, 16'd23861, 16'd57311, 16'd56628, 16'd34535, 16'd13066, 16'd54155});
	test_expansion(128'h1d78e12523c2e35c0cc233b13e8e046e, {16'd17554, 16'd44224, 16'd52210, 16'd41562, 16'd35756, 16'd2778, 16'd47589, 16'd57328, 16'd43240, 16'd56987, 16'd52087, 16'd2273, 16'd39070, 16'd41196, 16'd52925, 16'd40929, 16'd32549, 16'd52563, 16'd33468, 16'd24360, 16'd65260, 16'd15014, 16'd27204, 16'd16304, 16'd33932, 16'd39548});
	test_expansion(128'hdcb48307c249a3d49ea0f2245fbd8d8b, {16'd65331, 16'd54034, 16'd45812, 16'd54303, 16'd31156, 16'd4297, 16'd65176, 16'd17881, 16'd56330, 16'd16017, 16'd5263, 16'd13018, 16'd53091, 16'd58375, 16'd30902, 16'd23944, 16'd11265, 16'd32183, 16'd38931, 16'd27310, 16'd55235, 16'd31839, 16'd36640, 16'd29105, 16'd15644, 16'd37369});
	test_expansion(128'h3536018d4c7cd55dbf9b0fc9b4e5a750, {16'd10402, 16'd41789, 16'd59780, 16'd53916, 16'd34381, 16'd45100, 16'd6022, 16'd51210, 16'd50290, 16'd46947, 16'd39088, 16'd61245, 16'd34541, 16'd14635, 16'd30166, 16'd20449, 16'd61974, 16'd56138, 16'd4899, 16'd29548, 16'd23162, 16'd37116, 16'd12368, 16'd53372, 16'd51758, 16'd16940});
	test_expansion(128'h5f22ac85fcef878db923c50c1cd51b66, {16'd62269, 16'd48003, 16'd12233, 16'd636, 16'd61352, 16'd64311, 16'd38422, 16'd1757, 16'd35562, 16'd6131, 16'd20661, 16'd2966, 16'd14872, 16'd13712, 16'd41421, 16'd18159, 16'd42967, 16'd5423, 16'd48472, 16'd62961, 16'd13438, 16'd35188, 16'd8990, 16'd38428, 16'd50533, 16'd2083});
	test_expansion(128'h1a5bcb845b577e14ae41d9a34a5dc97e, {16'd22786, 16'd1252, 16'd51997, 16'd32832, 16'd22980, 16'd50114, 16'd24194, 16'd30882, 16'd11756, 16'd13169, 16'd16306, 16'd40495, 16'd43605, 16'd48337, 16'd20213, 16'd13883, 16'd43167, 16'd52054, 16'd33165, 16'd63249, 16'd54399, 16'd11301, 16'd22337, 16'd27631, 16'd9806, 16'd15833});
	test_expansion(128'he917413603b43f33907ba89e24ea10b4, {16'd14279, 16'd8583, 16'd3818, 16'd17178, 16'd48914, 16'd41567, 16'd21328, 16'd63125, 16'd20437, 16'd50508, 16'd33749, 16'd54823, 16'd46261, 16'd8360, 16'd26902, 16'd31935, 16'd6490, 16'd44626, 16'd64587, 16'd5080, 16'd55197, 16'd13020, 16'd22776, 16'd166, 16'd4326, 16'd60231});
	test_expansion(128'hd85d00adaa67f4b14258f3f24ba571f9, {16'd34616, 16'd39649, 16'd6058, 16'd58992, 16'd25061, 16'd4067, 16'd40269, 16'd43949, 16'd12513, 16'd42633, 16'd12004, 16'd3648, 16'd4146, 16'd58715, 16'd20323, 16'd5632, 16'd20225, 16'd45929, 16'd29115, 16'd19214, 16'd62957, 16'd63979, 16'd47172, 16'd21883, 16'd65479, 16'd61679});
	test_expansion(128'h340759ba832fdaa250c67550559524a7, {16'd36333, 16'd62742, 16'd21519, 16'd21811, 16'd4009, 16'd29197, 16'd28458, 16'd13920, 16'd9564, 16'd50530, 16'd8906, 16'd8430, 16'd47716, 16'd38120, 16'd30805, 16'd58349, 16'd24676, 16'd22939, 16'd40653, 16'd16311, 16'd59785, 16'd35954, 16'd42214, 16'd28112, 16'd46185, 16'd19541});
	test_expansion(128'h7b08b692d03198552bc6548f1876d7d4, {16'd58568, 16'd46031, 16'd58300, 16'd49571, 16'd43660, 16'd48974, 16'd37756, 16'd6406, 16'd60041, 16'd42464, 16'd44109, 16'd37815, 16'd39085, 16'd51578, 16'd28172, 16'd47642, 16'd22704, 16'd58241, 16'd13699, 16'd1615, 16'd15425, 16'd10227, 16'd48445, 16'd15790, 16'd14625, 16'd17991});
	test_expansion(128'hacecef465b201048bad03a7ee01f5543, {16'd53807, 16'd33241, 16'd16690, 16'd55359, 16'd33079, 16'd13929, 16'd60652, 16'd19195, 16'd54148, 16'd23855, 16'd42766, 16'd50486, 16'd6992, 16'd58979, 16'd3270, 16'd23100, 16'd11598, 16'd59561, 16'd10207, 16'd38802, 16'd1974, 16'd54527, 16'd28454, 16'd58394, 16'd40056, 16'd15691});
	test_expansion(128'h14b50858e3338289a74d5f9f6e1c5b15, {16'd10470, 16'd31695, 16'd21659, 16'd28130, 16'd11435, 16'd7898, 16'd3547, 16'd20306, 16'd6215, 16'd8481, 16'd13376, 16'd15023, 16'd32527, 16'd30112, 16'd1602, 16'd61094, 16'd19034, 16'd59246, 16'd48127, 16'd46108, 16'd64590, 16'd22768, 16'd52184, 16'd53131, 16'd45997, 16'd6493});
	test_expansion(128'h5601b24830fde3b886ca5ad2a4a972a2, {16'd57876, 16'd5129, 16'd35829, 16'd3626, 16'd63626, 16'd22920, 16'd17281, 16'd55554, 16'd60169, 16'd43375, 16'd64890, 16'd47207, 16'd33361, 16'd46740, 16'd30726, 16'd19128, 16'd51075, 16'd36128, 16'd15, 16'd34198, 16'd61056, 16'd15852, 16'd55808, 16'd16279, 16'd33579, 16'd45863});
	test_expansion(128'h72447599e17af3ac18278de69198e398, {16'd19663, 16'd45320, 16'd26640, 16'd52823, 16'd63514, 16'd10749, 16'd39427, 16'd56438, 16'd6944, 16'd37742, 16'd52715, 16'd22316, 16'd57184, 16'd11729, 16'd45142, 16'd11430, 16'd47362, 16'd7992, 16'd14153, 16'd6405, 16'd30940, 16'd48486, 16'd54152, 16'd59101, 16'd61460, 16'd31787});
	test_expansion(128'hd9fb687a9e89ae141e4c3d79b54370d4, {16'd1880, 16'd23662, 16'd64666, 16'd50985, 16'd19304, 16'd9484, 16'd44906, 16'd761, 16'd26943, 16'd37138, 16'd63304, 16'd54786, 16'd41664, 16'd21999, 16'd43780, 16'd50971, 16'd35162, 16'd58185, 16'd8294, 16'd37113, 16'd38720, 16'd51174, 16'd43664, 16'd37071, 16'd38517, 16'd41942});
	test_expansion(128'hf8e9c6788408b56c2fabcbed6c963f9c, {16'd10914, 16'd25900, 16'd40692, 16'd16960, 16'd56719, 16'd26933, 16'd55674, 16'd37492, 16'd44986, 16'd51222, 16'd33553, 16'd51097, 16'd36866, 16'd52636, 16'd42021, 16'd56415, 16'd30330, 16'd17585, 16'd4126, 16'd9563, 16'd41651, 16'd6573, 16'd54623, 16'd63391, 16'd59197, 16'd63571});
	test_expansion(128'he009898b22cdc4c340a9335cd928ccb3, {16'd45525, 16'd44101, 16'd9406, 16'd52517, 16'd30730, 16'd53019, 16'd3045, 16'd54688, 16'd53430, 16'd42575, 16'd64119, 16'd52823, 16'd18039, 16'd32796, 16'd46988, 16'd6438, 16'd11149, 16'd35855, 16'd19146, 16'd36671, 16'd43345, 16'd57971, 16'd2237, 16'd7279, 16'd2996, 16'd21459});
	test_expansion(128'hd5dd4763e41ba914672046cd67a6db0f, {16'd22500, 16'd27381, 16'd55111, 16'd51596, 16'd42900, 16'd30026, 16'd3199, 16'd31404, 16'd21542, 16'd37695, 16'd32714, 16'd47853, 16'd62952, 16'd572, 16'd44097, 16'd16299, 16'd38370, 16'd32557, 16'd30728, 16'd14645, 16'd28443, 16'd35166, 16'd48960, 16'd6792, 16'd60697, 16'd53253});
	test_expansion(128'ha0eb1ccac17759900fb3817db821d88d, {16'd7000, 16'd34778, 16'd19522, 16'd24429, 16'd21856, 16'd17673, 16'd14411, 16'd35248, 16'd44742, 16'd42633, 16'd12652, 16'd31178, 16'd40293, 16'd15950, 16'd24547, 16'd18716, 16'd60607, 16'd56420, 16'd2502, 16'd31922, 16'd42788, 16'd24901, 16'd45662, 16'd49462, 16'd13654, 16'd48848});
	test_expansion(128'hfbef23463d990d691ed2070c887f2152, {16'd63963, 16'd53783, 16'd14230, 16'd275, 16'd22367, 16'd3294, 16'd31352, 16'd15370, 16'd21209, 16'd53080, 16'd29701, 16'd11980, 16'd15841, 16'd34110, 16'd50593, 16'd26619, 16'd26820, 16'd14198, 16'd4722, 16'd53955, 16'd43932, 16'd54733, 16'd45165, 16'd28255, 16'd17761, 16'd12122});
	test_expansion(128'h6a6b5b92f7ed640ea056cabc52da72fe, {16'd17579, 16'd35152, 16'd5890, 16'd52813, 16'd43030, 16'd38911, 16'd22905, 16'd30016, 16'd11260, 16'd51129, 16'd31072, 16'd25429, 16'd63548, 16'd13140, 16'd10346, 16'd43174, 16'd8463, 16'd43187, 16'd43714, 16'd63741, 16'd17488, 16'd49121, 16'd38608, 16'd62125, 16'd41138, 16'd28564});
	test_expansion(128'hcd2847048edbaa87656bf3529c69b1ea, {16'd28574, 16'd52504, 16'd34932, 16'd26141, 16'd33304, 16'd58698, 16'd35464, 16'd50924, 16'd48806, 16'd33428, 16'd52647, 16'd49660, 16'd51253, 16'd42486, 16'd54930, 16'd37588, 16'd42122, 16'd6583, 16'd11477, 16'd9399, 16'd45236, 16'd11019, 16'd24079, 16'd25129, 16'd60719, 16'd39254});
	test_expansion(128'hc5df83c6161688f0c1834d246b628f9d, {16'd20103, 16'd25943, 16'd34745, 16'd47676, 16'd7796, 16'd4538, 16'd63040, 16'd24942, 16'd20077, 16'd14858, 16'd53364, 16'd27806, 16'd63160, 16'd15299, 16'd41676, 16'd23336, 16'd46140, 16'd59153, 16'd3950, 16'd11506, 16'd11937, 16'd45676, 16'd4716, 16'd36320, 16'd6326, 16'd10220});
	test_expansion(128'hb3ad14e39b6fadea7876f4f010741103, {16'd43001, 16'd57783, 16'd38338, 16'd17050, 16'd37505, 16'd64824, 16'd39100, 16'd15614, 16'd63750, 16'd52474, 16'd964, 16'd31220, 16'd44194, 16'd44679, 16'd59725, 16'd7826, 16'd63237, 16'd8997, 16'd46473, 16'd46881, 16'd63601, 16'd41205, 16'd63078, 16'd11591, 16'd35815, 16'd14843});
	test_expansion(128'h03e7a91bccf88759694bfcf963bcb579, {16'd22893, 16'd9154, 16'd7271, 16'd57975, 16'd5279, 16'd25477, 16'd54178, 16'd51838, 16'd50294, 16'd14907, 16'd60428, 16'd59834, 16'd758, 16'd16718, 16'd35434, 16'd13203, 16'd15370, 16'd16725, 16'd35523, 16'd18346, 16'd48021, 16'd61779, 16'd35870, 16'd34175, 16'd63538, 16'd4584});
	test_expansion(128'hcd1d778cf0049156f9d23f14f8258e01, {16'd39690, 16'd54699, 16'd18187, 16'd22500, 16'd58209, 16'd25399, 16'd893, 16'd39202, 16'd3674, 16'd11685, 16'd22823, 16'd46958, 16'd10250, 16'd21566, 16'd11718, 16'd596, 16'd50686, 16'd6422, 16'd447, 16'd25837, 16'd33759, 16'd41846, 16'd15491, 16'd11595, 16'd47530, 16'd38401});
	test_expansion(128'he5df43fd28e1c60c33e8a2a82400b97a, {16'd28360, 16'd42070, 16'd39112, 16'd7513, 16'd54994, 16'd37412, 16'd57721, 16'd32307, 16'd6224, 16'd20238, 16'd48509, 16'd22363, 16'd44414, 16'd55271, 16'd9041, 16'd61728, 16'd57760, 16'd10068, 16'd51524, 16'd25785, 16'd14381, 16'd62153, 16'd40364, 16'd23743, 16'd26485, 16'd58068});
	test_expansion(128'h17e7eefa8fec746779105939f0a4b9d5, {16'd41775, 16'd39967, 16'd16654, 16'd1081, 16'd20208, 16'd25268, 16'd5574, 16'd63275, 16'd58360, 16'd54786, 16'd25981, 16'd44172, 16'd20082, 16'd44822, 16'd59610, 16'd36337, 16'd12351, 16'd56184, 16'd22193, 16'd46398, 16'd63057, 16'd32479, 16'd61278, 16'd26924, 16'd29453, 16'd8673});
	test_expansion(128'hc07fb3156854b4f7f8011940e5e1c696, {16'd4688, 16'd28620, 16'd17459, 16'd12381, 16'd61682, 16'd422, 16'd64397, 16'd50868, 16'd9356, 16'd5061, 16'd40732, 16'd8350, 16'd65140, 16'd61494, 16'd31902, 16'd49911, 16'd36188, 16'd54325, 16'd2765, 16'd46865, 16'd61314, 16'd62523, 16'd41017, 16'd872, 16'd20565, 16'd39730});
	test_expansion(128'h60a543d088c3490387bd860fa88d6c9a, {16'd558, 16'd61328, 16'd58627, 16'd1851, 16'd19700, 16'd62994, 16'd9480, 16'd46543, 16'd51534, 16'd21992, 16'd35510, 16'd56714, 16'd41405, 16'd1698, 16'd7478, 16'd19289, 16'd44682, 16'd21065, 16'd57683, 16'd35763, 16'd42801, 16'd28336, 16'd29655, 16'd35714, 16'd62108, 16'd57516});
	test_expansion(128'he57f2ac579a7941003e87adf1723de76, {16'd22701, 16'd45358, 16'd30972, 16'd9082, 16'd12832, 16'd1100, 16'd5845, 16'd21605, 16'd22838, 16'd61828, 16'd38070, 16'd9475, 16'd8606, 16'd32394, 16'd2634, 16'd10551, 16'd28653, 16'd23228, 16'd20651, 16'd63156, 16'd52503, 16'd1240, 16'd40268, 16'd2548, 16'd55109, 16'd16909});
	test_expansion(128'h740e3563fe20494795edbf830ec202c3, {16'd59251, 16'd59358, 16'd59360, 16'd52558, 16'd8546, 16'd16344, 16'd25631, 16'd52254, 16'd9682, 16'd24369, 16'd22822, 16'd24832, 16'd1027, 16'd35728, 16'd39653, 16'd5266, 16'd10561, 16'd6714, 16'd32703, 16'd40200, 16'd1147, 16'd29235, 16'd46229, 16'd23286, 16'd9807, 16'd36750});
	test_expansion(128'hf8908edfe3d8797556409abc8c928973, {16'd64802, 16'd23476, 16'd30334, 16'd10457, 16'd36885, 16'd49413, 16'd30652, 16'd11324, 16'd23204, 16'd23886, 16'd1705, 16'd50467, 16'd48805, 16'd43766, 16'd13384, 16'd24172, 16'd64762, 16'd48699, 16'd21177, 16'd25148, 16'd29463, 16'd8754, 16'd35766, 16'd48984, 16'd46301, 16'd26355});
	test_expansion(128'h8425c59f589f18cf97d8ab13926259b1, {16'd32208, 16'd32726, 16'd6848, 16'd41764, 16'd23335, 16'd58633, 16'd42177, 16'd3902, 16'd11214, 16'd26959, 16'd33294, 16'd41239, 16'd7112, 16'd32742, 16'd22469, 16'd58955, 16'd63162, 16'd48142, 16'd15647, 16'd17555, 16'd7342, 16'd10607, 16'd20100, 16'd51448, 16'd61314, 16'd8522});
	test_expansion(128'hf46465581db4623382c5094e6691bbf3, {16'd41146, 16'd37729, 16'd23743, 16'd48673, 16'd48671, 16'd1661, 16'd33966, 16'd58093, 16'd33277, 16'd1733, 16'd63379, 16'd46623, 16'd39485, 16'd14910, 16'd42744, 16'd28499, 16'd54404, 16'd36627, 16'd63677, 16'd57192, 16'd5776, 16'd20879, 16'd12, 16'd61116, 16'd19007, 16'd59424});
	test_expansion(128'h13d4630d8e2accba605802055d2ea410, {16'd42742, 16'd41173, 16'd15460, 16'd41152, 16'd39802, 16'd30031, 16'd61916, 16'd58518, 16'd14590, 16'd16415, 16'd3010, 16'd4783, 16'd44851, 16'd61672, 16'd22110, 16'd25180, 16'd1360, 16'd24004, 16'd35520, 16'd8979, 16'd2327, 16'd26539, 16'd53325, 16'd17078, 16'd15637, 16'd12149});
	test_expansion(128'hef003c83ace167e7e1fc00e8151a094d, {16'd40277, 16'd43688, 16'd4687, 16'd54185, 16'd47400, 16'd1565, 16'd53576, 16'd30546, 16'd63074, 16'd64343, 16'd49893, 16'd42500, 16'd49977, 16'd18030, 16'd33486, 16'd10099, 16'd60735, 16'd55127, 16'd31403, 16'd27303, 16'd49148, 16'd13792, 16'd54621, 16'd63876, 16'd51753, 16'd11210});
	test_expansion(128'hb68ea05701b42edcbcc526866f0b3405, {16'd51285, 16'd26800, 16'd11657, 16'd47111, 16'd8092, 16'd1144, 16'd13190, 16'd2042, 16'd8028, 16'd31085, 16'd44996, 16'd15351, 16'd3969, 16'd25415, 16'd38467, 16'd10882, 16'd23370, 16'd8638, 16'd36174, 16'd39191, 16'd39084, 16'd17105, 16'd27896, 16'd29214, 16'd62851, 16'd23333});
	test_expansion(128'hd6cf9ba81d4f6feec862b7a5d5bd2165, {16'd65484, 16'd6206, 16'd46151, 16'd3433, 16'd46146, 16'd38256, 16'd4500, 16'd54943, 16'd30377, 16'd49647, 16'd23530, 16'd59283, 16'd18920, 16'd42068, 16'd15083, 16'd19436, 16'd26801, 16'd41782, 16'd53146, 16'd31345, 16'd20217, 16'd14012, 16'd40408, 16'd6223, 16'd55286, 16'd2643});
	test_expansion(128'h46d2e7b12718be28db0d9659a768248d, {16'd9706, 16'd52283, 16'd3695, 16'd8682, 16'd7261, 16'd18903, 16'd17930, 16'd56627, 16'd60568, 16'd49580, 16'd28441, 16'd55581, 16'd61766, 16'd8926, 16'd30862, 16'd19545, 16'd27016, 16'd5008, 16'd16377, 16'd5853, 16'd9068, 16'd39032, 16'd32904, 16'd39294, 16'd57708, 16'd57267});
	test_expansion(128'h0e1a0139ce686a84947c67c54d86f9d2, {16'd3107, 16'd28323, 16'd15275, 16'd17347, 16'd47509, 16'd41274, 16'd54720, 16'd14961, 16'd28955, 16'd3729, 16'd17478, 16'd27555, 16'd30155, 16'd28263, 16'd50230, 16'd48154, 16'd5588, 16'd48120, 16'd4592, 16'd59288, 16'd11117, 16'd26586, 16'd56211, 16'd64749, 16'd20302, 16'd21393});
	test_expansion(128'h9b95812c0ef1e40b4fefaed562264889, {16'd55607, 16'd32334, 16'd1995, 16'd60825, 16'd48098, 16'd55474, 16'd29847, 16'd53443, 16'd35185, 16'd20657, 16'd58428, 16'd56207, 16'd64688, 16'd46308, 16'd63920, 16'd22184, 16'd53313, 16'd1744, 16'd15318, 16'd36735, 16'd12689, 16'd751, 16'd39217, 16'd1391, 16'd47577, 16'd20687});
	test_expansion(128'he00f34c6f7a84fef8fb9d9b77f8e11b0, {16'd54530, 16'd41329, 16'd20538, 16'd30726, 16'd24362, 16'd16078, 16'd31296, 16'd44877, 16'd57098, 16'd35719, 16'd40531, 16'd11267, 16'd17955, 16'd51535, 16'd13693, 16'd44155, 16'd4358, 16'd17492, 16'd59366, 16'd22723, 16'd32360, 16'd45226, 16'd12907, 16'd52394, 16'd15540, 16'd21172});
	test_expansion(128'h80a2548a45248d9835988ad959086db5, {16'd32774, 16'd7527, 16'd38029, 16'd57788, 16'd39406, 16'd40448, 16'd49540, 16'd8963, 16'd33341, 16'd25183, 16'd37769, 16'd46205, 16'd56584, 16'd8438, 16'd43930, 16'd43072, 16'd28324, 16'd37664, 16'd11369, 16'd21753, 16'd41159, 16'd29489, 16'd19034, 16'd3136, 16'd61939, 16'd30800});
	test_expansion(128'h4c912837ab8ca2f9f9bed9cd4739998b, {16'd63360, 16'd53725, 16'd19624, 16'd62849, 16'd56750, 16'd62669, 16'd17069, 16'd42871, 16'd30873, 16'd14686, 16'd22716, 16'd8386, 16'd67, 16'd11345, 16'd56587, 16'd45015, 16'd14044, 16'd27823, 16'd10232, 16'd55492, 16'd61399, 16'd62380, 16'd53893, 16'd26600, 16'd58355, 16'd1973});
	test_expansion(128'h934bad4ddadf6643ec7d1c8b991815ae, {16'd59433, 16'd49011, 16'd55605, 16'd19383, 16'd33077, 16'd62413, 16'd55179, 16'd18757, 16'd56491, 16'd59334, 16'd45105, 16'd60232, 16'd17565, 16'd6339, 16'd1638, 16'd19818, 16'd17687, 16'd35151, 16'd23051, 16'd32079, 16'd62956, 16'd64598, 16'd32222, 16'd31358, 16'd3935, 16'd55291});
	test_expansion(128'hef7c2e85df4bcb65b9e47e723dbfcd9e, {16'd31413, 16'd55722, 16'd26583, 16'd50590, 16'd55925, 16'd10782, 16'd7151, 16'd30757, 16'd50315, 16'd32726, 16'd47138, 16'd31166, 16'd5778, 16'd37246, 16'd32289, 16'd3102, 16'd58040, 16'd3984, 16'd8045, 16'd26584, 16'd21057, 16'd59145, 16'd43182, 16'd38676, 16'd36881, 16'd54700});
	test_expansion(128'h8269747a6b0f22ecbbf55da5d65a33fe, {16'd51579, 16'd59776, 16'd57924, 16'd36082, 16'd10244, 16'd19398, 16'd14511, 16'd8662, 16'd7342, 16'd37393, 16'd31822, 16'd38, 16'd17381, 16'd45694, 16'd225, 16'd53077, 16'd27022, 16'd8062, 16'd50238, 16'd23385, 16'd39039, 16'd17281, 16'd55797, 16'd39343, 16'd55861, 16'd31357});
	test_expansion(128'h9be41e173465c6e4fec021082c9ee527, {16'd49870, 16'd16448, 16'd56529, 16'd9938, 16'd14854, 16'd38362, 16'd27270, 16'd34936, 16'd45990, 16'd31141, 16'd4980, 16'd58453, 16'd9318, 16'd34939, 16'd18750, 16'd47341, 16'd29587, 16'd40234, 16'd57384, 16'd30494, 16'd58685, 16'd45031, 16'd19009, 16'd32619, 16'd9233, 16'd58439});
	test_expansion(128'h0684f39016cf5f90c48617934a31d2ee, {16'd50213, 16'd56209, 16'd61601, 16'd35291, 16'd8167, 16'd30289, 16'd35433, 16'd34847, 16'd25668, 16'd4458, 16'd64930, 16'd7289, 16'd53165, 16'd48420, 16'd59869, 16'd48659, 16'd55925, 16'd47105, 16'd37983, 16'd2428, 16'd12315, 16'd38439, 16'd33636, 16'd8539, 16'd5131, 16'd36222});
	test_expansion(128'hddf79702abb7d9a1d6d4ba7ae6586432, {16'd18770, 16'd64613, 16'd33907, 16'd14045, 16'd10587, 16'd27171, 16'd1590, 16'd47608, 16'd45875, 16'd19983, 16'd8669, 16'd46253, 16'd64903, 16'd5270, 16'd34981, 16'd57120, 16'd3467, 16'd12978, 16'd14389, 16'd18854, 16'd5637, 16'd50481, 16'd32168, 16'd47394, 16'd32645, 16'd57058});
	test_expansion(128'hdfe443e58a7bf5a44f5df8701cf25ccc, {16'd31282, 16'd26103, 16'd38765, 16'd52079, 16'd64266, 16'd34743, 16'd31069, 16'd34152, 16'd53191, 16'd49402, 16'd30064, 16'd8620, 16'd29211, 16'd33247, 16'd56974, 16'd63885, 16'd37904, 16'd16110, 16'd7535, 16'd13330, 16'd37828, 16'd4699, 16'd26798, 16'd36589, 16'd36853, 16'd39668});
	test_expansion(128'h3b5aa34b31baa4a2a42a0ba441f4d939, {16'd3209, 16'd64604, 16'd42649, 16'd23231, 16'd38956, 16'd57576, 16'd54766, 16'd211, 16'd4301, 16'd15302, 16'd11025, 16'd25360, 16'd30617, 16'd11065, 16'd22426, 16'd45644, 16'd37015, 16'd63819, 16'd51473, 16'd60002, 16'd9056, 16'd34559, 16'd43840, 16'd8504, 16'd7678, 16'd15502});
	test_expansion(128'ha9db986733f64114ceb9f861f68dd891, {16'd33107, 16'd44868, 16'd58520, 16'd29248, 16'd46681, 16'd36068, 16'd40022, 16'd21143, 16'd32180, 16'd12440, 16'd33877, 16'd16040, 16'd47667, 16'd47883, 16'd15850, 16'd20753, 16'd58759, 16'd46387, 16'd2775, 16'd5842, 16'd4232, 16'd60304, 16'd38164, 16'd5500, 16'd52552, 16'd45748});
	test_expansion(128'hc5815e9b187ec620d97d7f70df4eaf78, {16'd45148, 16'd24208, 16'd8412, 16'd57861, 16'd64259, 16'd56754, 16'd19426, 16'd38744, 16'd26160, 16'd44280, 16'd15518, 16'd15630, 16'd9444, 16'd21284, 16'd39195, 16'd25800, 16'd42444, 16'd30745, 16'd25478, 16'd13656, 16'd36802, 16'd6967, 16'd26405, 16'd61876, 16'd57253, 16'd50402});
	test_expansion(128'hee6f00e91586274f1076c7da700e8fd5, {16'd60913, 16'd28351, 16'd53556, 16'd7525, 16'd25111, 16'd46845, 16'd23358, 16'd55612, 16'd5210, 16'd52247, 16'd16512, 16'd58975, 16'd18484, 16'd59818, 16'd38735, 16'd27855, 16'd43944, 16'd42756, 16'd26003, 16'd59543, 16'd53207, 16'd13626, 16'd31293, 16'd12842, 16'd30585, 16'd61473});
	test_expansion(128'h7f1878b6edc54dc7c57234a75bee7f2a, {16'd19535, 16'd53332, 16'd46547, 16'd16483, 16'd57606, 16'd53724, 16'd60994, 16'd2766, 16'd980, 16'd12562, 16'd32331, 16'd11790, 16'd62737, 16'd51827, 16'd40930, 16'd54501, 16'd38481, 16'd48464, 16'd44392, 16'd11717, 16'd2666, 16'd31071, 16'd46169, 16'd44613, 16'd25898, 16'd25910});
	test_expansion(128'hc42b319db334659b05ee1bbfd885ad70, {16'd13198, 16'd49812, 16'd54228, 16'd61791, 16'd7550, 16'd27712, 16'd46898, 16'd37244, 16'd21969, 16'd23584, 16'd34549, 16'd41488, 16'd18346, 16'd7596, 16'd23108, 16'd59766, 16'd29540, 16'd55842, 16'd55828, 16'd61614, 16'd53176, 16'd25848, 16'd33426, 16'd40448, 16'd62821, 16'd42203});
	test_expansion(128'h9d715e3b1db54ffc636c2930c47673c8, {16'd55089, 16'd43718, 16'd12212, 16'd46799, 16'd30302, 16'd13134, 16'd11769, 16'd28045, 16'd35578, 16'd43764, 16'd18172, 16'd33953, 16'd60236, 16'd49535, 16'd32582, 16'd52524, 16'd114, 16'd52059, 16'd59176, 16'd61259, 16'd32139, 16'd40757, 16'd26880, 16'd23764, 16'd44567, 16'd53731});
	test_expansion(128'hf994ac1a6ea0aa725f30cb06e2114c5b, {16'd23377, 16'd16431, 16'd43885, 16'd45658, 16'd17162, 16'd3965, 16'd54590, 16'd1208, 16'd5295, 16'd36577, 16'd58420, 16'd22440, 16'd60321, 16'd26399, 16'd52236, 16'd39245, 16'd63378, 16'd5166, 16'd41046, 16'd35826, 16'd49725, 16'd53175, 16'd11851, 16'd62571, 16'd58636, 16'd60921});
	test_expansion(128'heb7633ec01db41f03bfc0881c18f48c8, {16'd57946, 16'd1059, 16'd33256, 16'd47952, 16'd55536, 16'd38150, 16'd55408, 16'd2529, 16'd58788, 16'd5332, 16'd35452, 16'd62688, 16'd12102, 16'd21304, 16'd46025, 16'd52814, 16'd33884, 16'd11833, 16'd28577, 16'd18704, 16'd63907, 16'd18418, 16'd16403, 16'd30902, 16'd63780, 16'd1202});
	test_expansion(128'h6bf7cfb7ee44b54b557979f7ad1e491f, {16'd18933, 16'd54944, 16'd53698, 16'd53805, 16'd53203, 16'd58379, 16'd60150, 16'd48398, 16'd58888, 16'd30235, 16'd53052, 16'd26030, 16'd560, 16'd22300, 16'd3291, 16'd23594, 16'd10860, 16'd46945, 16'd31107, 16'd7272, 16'd58546, 16'd55697, 16'd36567, 16'd39928, 16'd39386, 16'd27031});
	test_expansion(128'h7a847c86dbb538de0d0305d9811415a8, {16'd54145, 16'd40592, 16'd44154, 16'd593, 16'd63280, 16'd3156, 16'd50879, 16'd51656, 16'd53869, 16'd15489, 16'd6216, 16'd29340, 16'd32614, 16'd60554, 16'd36912, 16'd12648, 16'd40351, 16'd12978, 16'd52753, 16'd38058, 16'd31414, 16'd5946, 16'd57710, 16'd6687, 16'd42872, 16'd33842});
	test_expansion(128'h1582050be66b9d3fd25cacd75339a04e, {16'd25905, 16'd57523, 16'd34339, 16'd37458, 16'd4059, 16'd28290, 16'd53285, 16'd25946, 16'd51227, 16'd28110, 16'd13281, 16'd60888, 16'd1070, 16'd46873, 16'd4965, 16'd44007, 16'd2047, 16'd54190, 16'd50831, 16'd65443, 16'd49652, 16'd21561, 16'd18233, 16'd61815, 16'd36076, 16'd60912});
	test_expansion(128'hc6e7df037f082b035f041c826795167d, {16'd62321, 16'd15456, 16'd40626, 16'd47324, 16'd57775, 16'd14644, 16'd63717, 16'd7786, 16'd45431, 16'd14026, 16'd11067, 16'd5158, 16'd63248, 16'd26467, 16'd61016, 16'd64751, 16'd5326, 16'd51887, 16'd16882, 16'd59276, 16'd46089, 16'd8924, 16'd10701, 16'd40401, 16'd32416, 16'd9097});
	test_expansion(128'h65c043faee270d96f48894d8d76846b2, {16'd17194, 16'd51439, 16'd12455, 16'd8991, 16'd58687, 16'd13198, 16'd51298, 16'd14696, 16'd54788, 16'd1381, 16'd49606, 16'd31642, 16'd40433, 16'd22743, 16'd30504, 16'd12579, 16'd23752, 16'd30135, 16'd8900, 16'd38582, 16'd3613, 16'd18733, 16'd33206, 16'd28789, 16'd30498, 16'd25026});
	test_expansion(128'h94ef4726e9de8dbb3f72668d125a4a0b, {16'd63635, 16'd39335, 16'd10628, 16'd42609, 16'd16361, 16'd33183, 16'd59043, 16'd11140, 16'd51556, 16'd53500, 16'd31096, 16'd51390, 16'd42081, 16'd9759, 16'd63172, 16'd10538, 16'd39335, 16'd53600, 16'd12168, 16'd11820, 16'd61957, 16'd45992, 16'd19026, 16'd32580, 16'd19281, 16'd12892});
	test_expansion(128'hefc9154162f1d8b2cc18bcc053aa92fa, {16'd39626, 16'd1813, 16'd35980, 16'd54443, 16'd31558, 16'd6144, 16'd24699, 16'd20944, 16'd11678, 16'd48853, 16'd27438, 16'd26030, 16'd59130, 16'd41322, 16'd47034, 16'd28901, 16'd11409, 16'd25118, 16'd61554, 16'd44929, 16'd36274, 16'd64633, 16'd49318, 16'd50258, 16'd18077, 16'd49483});
	test_expansion(128'h5861a98f18a6476c5e1016917e3e6dd0, {16'd19917, 16'd10754, 16'd6029, 16'd29026, 16'd47560, 16'd17832, 16'd6986, 16'd35847, 16'd56285, 16'd12447, 16'd8529, 16'd17177, 16'd40900, 16'd8111, 16'd14396, 16'd37232, 16'd25298, 16'd28076, 16'd51628, 16'd42210, 16'd32144, 16'd60366, 16'd20629, 16'd13973, 16'd57875, 16'd29486});
	test_expansion(128'h018f795649d3f1d0d806276eedf6798d, {16'd43532, 16'd60692, 16'd25566, 16'd46614, 16'd6786, 16'd4552, 16'd21038, 16'd37472, 16'd63547, 16'd41469, 16'd16925, 16'd63970, 16'd24832, 16'd57513, 16'd12777, 16'd29754, 16'd39875, 16'd37747, 16'd46174, 16'd64356, 16'd36356, 16'd40522, 16'd52682, 16'd50730, 16'd48880, 16'd19863});
	test_expansion(128'h8b4313d6ce93469c3c0e9ac57eccea0c, {16'd22627, 16'd24811, 16'd55731, 16'd53875, 16'd61185, 16'd4115, 16'd59229, 16'd64798, 16'd59857, 16'd41107, 16'd64614, 16'd26227, 16'd26303, 16'd15968, 16'd12484, 16'd55784, 16'd22567, 16'd1975, 16'd12954, 16'd13577, 16'd13990, 16'd43232, 16'd32976, 16'd6037, 16'd46299, 16'd21633});
	test_expansion(128'h4c56c16e234c0388642ce982a8be6e1d, {16'd43577, 16'd7167, 16'd44444, 16'd10068, 16'd34862, 16'd513, 16'd51956, 16'd17036, 16'd13509, 16'd58981, 16'd53849, 16'd63710, 16'd50816, 16'd57479, 16'd23439, 16'd36247, 16'd39870, 16'd45909, 16'd24155, 16'd1491, 16'd13652, 16'd46840, 16'd39451, 16'd28621, 16'd28204, 16'd40223});
	test_expansion(128'h626804eb7ea73925884c5269ab4c9416, {16'd21956, 16'd64505, 16'd15808, 16'd61331, 16'd30326, 16'd36319, 16'd54676, 16'd20032, 16'd627, 16'd57447, 16'd7136, 16'd56519, 16'd10381, 16'd29678, 16'd39409, 16'd56309, 16'd28802, 16'd44844, 16'd16010, 16'd49691, 16'd37509, 16'd51531, 16'd56588, 16'd634, 16'd58730, 16'd32462});
	test_expansion(128'h47a11c61fa9b6664e43ae903ba72d47e, {16'd59682, 16'd65417, 16'd8058, 16'd48571, 16'd64557, 16'd54210, 16'd45745, 16'd50321, 16'd48335, 16'd51880, 16'd59588, 16'd37611, 16'd35125, 16'd35754, 16'd64759, 16'd21111, 16'd50564, 16'd38598, 16'd25139, 16'd31145, 16'd13267, 16'd61066, 16'd55962, 16'd58831, 16'd29332, 16'd21861});
	test_expansion(128'h32bfecfd0d610f2f9d6ee154030c22b0, {16'd54721, 16'd43281, 16'd23463, 16'd57759, 16'd55281, 16'd18610, 16'd39987, 16'd16150, 16'd36953, 16'd42672, 16'd63805, 16'd31546, 16'd59417, 16'd35768, 16'd3383, 16'd43463, 16'd39817, 16'd33775, 16'd28225, 16'd61987, 16'd30744, 16'd52025, 16'd42216, 16'd39949, 16'd52733, 16'd14758});
	test_expansion(128'hb7f6236f18ab47b5454842dbb251a95d, {16'd32876, 16'd54080, 16'd61928, 16'd20927, 16'd20395, 16'd14805, 16'd57110, 16'd2979, 16'd8538, 16'd38197, 16'd25207, 16'd24093, 16'd52986, 16'd26712, 16'd55987, 16'd6093, 16'd57816, 16'd14221, 16'd62587, 16'd16840, 16'd65200, 16'd43334, 16'd3461, 16'd53664, 16'd52701, 16'd29493});
	test_expansion(128'hc919c57c9c7e4a6162162c3c42878970, {16'd30801, 16'd53188, 16'd40856, 16'd37552, 16'd60776, 16'd9286, 16'd15479, 16'd5597, 16'd3197, 16'd61612, 16'd8065, 16'd33130, 16'd11130, 16'd39048, 16'd21435, 16'd45281, 16'd20479, 16'd56268, 16'd25884, 16'd15308, 16'd56418, 16'd41532, 16'd33584, 16'd20108, 16'd50626, 16'd62373});
	test_expansion(128'hfd4b940982764ab999b44ecb550dc42b, {16'd13746, 16'd18665, 16'd5255, 16'd33548, 16'd32719, 16'd17051, 16'd27602, 16'd10202, 16'd118, 16'd24003, 16'd34264, 16'd63597, 16'd39940, 16'd17231, 16'd55120, 16'd44327, 16'd36014, 16'd36967, 16'd12229, 16'd59021, 16'd2785, 16'd5776, 16'd58001, 16'd1850, 16'd28089, 16'd51224});
	test_expansion(128'h3b00e7a3c13cf2e14fff83a3db4a373f, {16'd34139, 16'd41066, 16'd38934, 16'd48939, 16'd41776, 16'd37347, 16'd6989, 16'd117, 16'd51412, 16'd16700, 16'd4008, 16'd29614, 16'd4689, 16'd63089, 16'd14351, 16'd492, 16'd60601, 16'd53435, 16'd9538, 16'd31632, 16'd10105, 16'd12844, 16'd1725, 16'd4203, 16'd27112, 16'd62754});
	test_expansion(128'h7e099013978281b84713305ccfbb889f, {16'd37711, 16'd11942, 16'd25956, 16'd11651, 16'd31232, 16'd64165, 16'd9233, 16'd45583, 16'd44507, 16'd30452, 16'd5481, 16'd36548, 16'd3916, 16'd20375, 16'd58422, 16'd27341, 16'd50584, 16'd36110, 16'd33127, 16'd32304, 16'd45499, 16'd41239, 16'd10734, 16'd63286, 16'd43709, 16'd32534});
	test_expansion(128'h62d7a3af51ed50b06a767a410e9ccfa2, {16'd18021, 16'd3594, 16'd4049, 16'd58785, 16'd41137, 16'd44014, 16'd10671, 16'd21053, 16'd38154, 16'd2369, 16'd6866, 16'd47179, 16'd54126, 16'd43547, 16'd41236, 16'd21978, 16'd52117, 16'd6955, 16'd12067, 16'd5001, 16'd9686, 16'd38033, 16'd44704, 16'd32385, 16'd38226, 16'd29282});
	test_expansion(128'h3877b7245a9994cd4c5f55036e155143, {16'd13458, 16'd37937, 16'd63927, 16'd13905, 16'd28390, 16'd46147, 16'd12953, 16'd52205, 16'd26433, 16'd30761, 16'd26426, 16'd24604, 16'd6048, 16'd53118, 16'd54697, 16'd8080, 16'd54710, 16'd36637, 16'd52045, 16'd1194, 16'd12998, 16'd22462, 16'd5270, 16'd60770, 16'd34914, 16'd45715});
	test_expansion(128'hca6f4672dc11810c868c1f65bbc18187, {16'd10443, 16'd10469, 16'd57485, 16'd11797, 16'd5678, 16'd46059, 16'd8396, 16'd57416, 16'd44372, 16'd22173, 16'd8393, 16'd33291, 16'd33716, 16'd54011, 16'd49832, 16'd33127, 16'd49822, 16'd835, 16'd51612, 16'd3078, 16'd14679, 16'd28515, 16'd49748, 16'd43662, 16'd8736, 16'd15578});
	test_expansion(128'hc4d586699121519b5efc9bd1bf6061fc, {16'd16842, 16'd18423, 16'd47588, 16'd8710, 16'd9843, 16'd51705, 16'd1160, 16'd47295, 16'd27135, 16'd37716, 16'd50377, 16'd36209, 16'd20350, 16'd37226, 16'd23641, 16'd32826, 16'd19870, 16'd31894, 16'd53789, 16'd51716, 16'd20622, 16'd16648, 16'd48706, 16'd47984, 16'd4714, 16'd17157});
	test_expansion(128'h0170831d2b823b37c6f9c178eac55eed, {16'd49880, 16'd31731, 16'd2725, 16'd18568, 16'd60347, 16'd50940, 16'd18076, 16'd31331, 16'd16857, 16'd14076, 16'd39322, 16'd64955, 16'd20774, 16'd16378, 16'd22920, 16'd60252, 16'd26395, 16'd43156, 16'd20862, 16'd10790, 16'd30471, 16'd55830, 16'd582, 16'd40418, 16'd39220, 16'd18084});
	test_expansion(128'h06707724edec7038e56e00b4bd9bd51f, {16'd7470, 16'd58171, 16'd64841, 16'd5029, 16'd54166, 16'd33757, 16'd12075, 16'd52595, 16'd47433, 16'd34236, 16'd39392, 16'd60890, 16'd32165, 16'd24512, 16'd9738, 16'd61579, 16'd57072, 16'd21982, 16'd44605, 16'd48613, 16'd32414, 16'd61684, 16'd50301, 16'd57684, 16'd33146, 16'd40724});
	test_expansion(128'hba53e9c1fe17fb48ffaa1cb93fcef024, {16'd51936, 16'd50591, 16'd34733, 16'd60323, 16'd25619, 16'd7311, 16'd42681, 16'd53415, 16'd46280, 16'd40041, 16'd64275, 16'd39005, 16'd44384, 16'd52248, 16'd32128, 16'd12746, 16'd7857, 16'd15947, 16'd41063, 16'd23305, 16'd48131, 16'd35099, 16'd16397, 16'd7357, 16'd31628, 16'd10625});
	test_expansion(128'h4d108361e77a05aa935279ff42b7e645, {16'd61057, 16'd52873, 16'd63981, 16'd38985, 16'd54048, 16'd59716, 16'd56936, 16'd10933, 16'd44600, 16'd57959, 16'd64869, 16'd27331, 16'd61645, 16'd47749, 16'd2792, 16'd50528, 16'd12076, 16'd51011, 16'd15794, 16'd49018, 16'd2797, 16'd24703, 16'd40474, 16'd18251, 16'd41393, 16'd35817});
	test_expansion(128'h13f27c2ca63c0e6cdf0469fde7fc22d3, {16'd42293, 16'd15315, 16'd1588, 16'd2250, 16'd41340, 16'd21606, 16'd38250, 16'd4627, 16'd35391, 16'd53111, 16'd23624, 16'd47396, 16'd63216, 16'd3468, 16'd4163, 16'd30601, 16'd21897, 16'd51648, 16'd44592, 16'd60692, 16'd48536, 16'd2747, 16'd15396, 16'd63276, 16'd62905, 16'd50316});
	test_expansion(128'h71ec380405351aafc953f8f78e2a294e, {16'd21652, 16'd52200, 16'd21651, 16'd10720, 16'd51613, 16'd64926, 16'd16470, 16'd60552, 16'd47315, 16'd33413, 16'd50937, 16'd3980, 16'd833, 16'd59008, 16'd40128, 16'd21165, 16'd21010, 16'd54256, 16'd13527, 16'd62481, 16'd51593, 16'd28332, 16'd40874, 16'd34059, 16'd24536, 16'd54088});
	test_expansion(128'hb0ae837d1c4da48580102f4d1f8d270a, {16'd41423, 16'd5750, 16'd53406, 16'd30562, 16'd59302, 16'd10685, 16'd8404, 16'd41814, 16'd17743, 16'd9420, 16'd29166, 16'd37713, 16'd50723, 16'd35739, 16'd17384, 16'd48827, 16'd34029, 16'd10053, 16'd13449, 16'd3048, 16'd18697, 16'd12293, 16'd31961, 16'd38188, 16'd18705, 16'd11362});
	test_expansion(128'h2b95f8feeda7874ae4bd45f028f73dad, {16'd33050, 16'd8324, 16'd30107, 16'd18537, 16'd27650, 16'd37953, 16'd16003, 16'd16458, 16'd60290, 16'd46816, 16'd16924, 16'd5160, 16'd35588, 16'd61004, 16'd24110, 16'd65439, 16'd36613, 16'd28770, 16'd48101, 16'd12852, 16'd39239, 16'd30977, 16'd15787, 16'd13393, 16'd45411, 16'd8950});
	test_expansion(128'h6a095130367ea7e465433531de329ca2, {16'd51275, 16'd34974, 16'd54212, 16'd50982, 16'd22038, 16'd4948, 16'd52966, 16'd21806, 16'd28530, 16'd57132, 16'd44840, 16'd56002, 16'd13524, 16'd42065, 16'd36660, 16'd14496, 16'd31643, 16'd49227, 16'd12157, 16'd58544, 16'd64881, 16'd40657, 16'd31750, 16'd14915, 16'd8283, 16'd49980});
	test_expansion(128'h40332c93f7a889af12ccfdc1d4900d92, {16'd54783, 16'd24559, 16'd25327, 16'd36941, 16'd24128, 16'd30991, 16'd24312, 16'd29245, 16'd65167, 16'd30298, 16'd29387, 16'd16709, 16'd44800, 16'd23287, 16'd49738, 16'd55646, 16'd51892, 16'd34964, 16'd29450, 16'd57032, 16'd58291, 16'd51530, 16'd51798, 16'd46284, 16'd22113, 16'd28054});
	test_expansion(128'hd825f8ef0c9907f1e07edd842b6aa479, {16'd16300, 16'd45012, 16'd62161, 16'd46614, 16'd39118, 16'd33076, 16'd43581, 16'd5330, 16'd10579, 16'd56565, 16'd16866, 16'd49490, 16'd46739, 16'd26751, 16'd29519, 16'd35390, 16'd42729, 16'd9089, 16'd52597, 16'd41761, 16'd43928, 16'd21166, 16'd11864, 16'd13908, 16'd11681, 16'd22238});
	test_expansion(128'h928ebafc0f3e418f503278d9f5f8ac10, {16'd10581, 16'd7525, 16'd9992, 16'd38647, 16'd35807, 16'd39583, 16'd18605, 16'd63963, 16'd9903, 16'd42744, 16'd61540, 16'd61820, 16'd15019, 16'd10612, 16'd50975, 16'd4266, 16'd52200, 16'd3059, 16'd58906, 16'd48477, 16'd18358, 16'd2497, 16'd36253, 16'd43449, 16'd25338, 16'd40075});
	test_expansion(128'h92153de69b4d5229c7580dfbdf7808f4, {16'd682, 16'd62755, 16'd49740, 16'd27441, 16'd32493, 16'd8242, 16'd49301, 16'd45699, 16'd18733, 16'd40375, 16'd51491, 16'd41939, 16'd60451, 16'd13776, 16'd17676, 16'd36868, 16'd55592, 16'd53094, 16'd37350, 16'd19391, 16'd38653, 16'd5840, 16'd1823, 16'd30180, 16'd62471, 16'd32574});
	test_expansion(128'hb69ab959e546c2df126689bca46b60b2, {16'd65213, 16'd26672, 16'd21234, 16'd61144, 16'd52477, 16'd24448, 16'd31492, 16'd52089, 16'd44401, 16'd8531, 16'd32665, 16'd4048, 16'd19793, 16'd59025, 16'd25116, 16'd1202, 16'd60256, 16'd63992, 16'd45212, 16'd46988, 16'd40858, 16'd48131, 16'd24518, 16'd2761, 16'd5541, 16'd45283});
	test_expansion(128'hdadd95b0d983610047599feb36308f34, {16'd21607, 16'd59425, 16'd18339, 16'd41626, 16'd58919, 16'd9108, 16'd36133, 16'd8493, 16'd12025, 16'd56624, 16'd18588, 16'd52886, 16'd9882, 16'd20180, 16'd58476, 16'd62499, 16'd38521, 16'd20592, 16'd45930, 16'd59921, 16'd18456, 16'd34261, 16'd51857, 16'd30160, 16'd7692, 16'd64129});
	test_expansion(128'h0891b082b24f2a8365346c51972e3acd, {16'd57361, 16'd2324, 16'd30798, 16'd9079, 16'd57381, 16'd10679, 16'd58157, 16'd19360, 16'd16788, 16'd47739, 16'd24459, 16'd25632, 16'd19540, 16'd63315, 16'd50840, 16'd26491, 16'd52864, 16'd29990, 16'd10279, 16'd15776, 16'd27354, 16'd16619, 16'd18602, 16'd25511, 16'd4216, 16'd45374});
	test_expansion(128'h8435f362dcaea0c0c70bdf699fd10121, {16'd14872, 16'd56186, 16'd61529, 16'd23090, 16'd48345, 16'd31654, 16'd63263, 16'd13566, 16'd22774, 16'd7754, 16'd39879, 16'd14376, 16'd58838, 16'd40772, 16'd14378, 16'd36180, 16'd39631, 16'd42260, 16'd36788, 16'd39397, 16'd25048, 16'd41508, 16'd8341, 16'd45432, 16'd34104, 16'd6672});
	test_expansion(128'hfb5f09d86b9e90a6a7e62e35dcb95788, {16'd10457, 16'd48418, 16'd19078, 16'd47952, 16'd57489, 16'd17421, 16'd43541, 16'd54464, 16'd49163, 16'd35017, 16'd44681, 16'd56947, 16'd2702, 16'd37870, 16'd25098, 16'd42620, 16'd27418, 16'd46353, 16'd57093, 16'd8968, 16'd55096, 16'd38235, 16'd42358, 16'd48092, 16'd46901, 16'd46560});
	test_expansion(128'h167980155399a01972be811dbad891e2, {16'd35897, 16'd39630, 16'd27167, 16'd11687, 16'd6658, 16'd54426, 16'd29587, 16'd39244, 16'd59775, 16'd62519, 16'd32623, 16'd31802, 16'd9864, 16'd35005, 16'd62451, 16'd51789, 16'd11840, 16'd63135, 16'd15996, 16'd18004, 16'd63872, 16'd34434, 16'd56719, 16'd56863, 16'd62685, 16'd45494});
	test_expansion(128'hf0562f612dccf032358fa7289d739039, {16'd3158, 16'd30767, 16'd36857, 16'd21371, 16'd64245, 16'd25485, 16'd5433, 16'd62333, 16'd55306, 16'd19519, 16'd20591, 16'd34763, 16'd57186, 16'd35051, 16'd65171, 16'd8811, 16'd5489, 16'd30336, 16'd65204, 16'd15905, 16'd56722, 16'd20719, 16'd37954, 16'd15673, 16'd54093, 16'd16219});
	test_expansion(128'h543c95341332c82995ef36d6196d4edd, {16'd29574, 16'd48821, 16'd45564, 16'd25259, 16'd21659, 16'd51274, 16'd971, 16'd385, 16'd25353, 16'd49751, 16'd31614, 16'd54357, 16'd43757, 16'd30094, 16'd63946, 16'd55419, 16'd17152, 16'd42890, 16'd27223, 16'd8495, 16'd64168, 16'd27633, 16'd51820, 16'd53858, 16'd28370, 16'd45873});
	test_expansion(128'haffd66107b92a8a9a69842b2c33e3084, {16'd52942, 16'd53528, 16'd49483, 16'd18765, 16'd28147, 16'd42068, 16'd54931, 16'd23233, 16'd52676, 16'd47729, 16'd1855, 16'd18757, 16'd30586, 16'd30465, 16'd35286, 16'd52052, 16'd55674, 16'd35253, 16'd45319, 16'd57601, 16'd50383, 16'd8655, 16'd7415, 16'd21403, 16'd44623, 16'd34352});
	test_expansion(128'h3ee37401a7bcbc67b905530900fe1011, {16'd56552, 16'd51568, 16'd53407, 16'd16959, 16'd50220, 16'd58040, 16'd65030, 16'd19941, 16'd596, 16'd21799, 16'd29864, 16'd58975, 16'd18565, 16'd29086, 16'd56314, 16'd29807, 16'd776, 16'd51381, 16'd32026, 16'd23824, 16'd49343, 16'd29264, 16'd26466, 16'd55015, 16'd52591, 16'd23720});
	test_expansion(128'hb832e63eb785fb2f2a4370ccaa66c1ce, {16'd13826, 16'd43428, 16'd18429, 16'd11317, 16'd61090, 16'd36446, 16'd45513, 16'd18544, 16'd43629, 16'd46461, 16'd52228, 16'd8697, 16'd11999, 16'd10459, 16'd7426, 16'd61306, 16'd34326, 16'd54480, 16'd59606, 16'd13616, 16'd34744, 16'd31153, 16'd44088, 16'd12030, 16'd61823, 16'd40018});
	test_expansion(128'hfa1ec0122d4a7d394c5729c0113ef2e2, {16'd13289, 16'd9151, 16'd61961, 16'd33123, 16'd26520, 16'd56844, 16'd54816, 16'd28582, 16'd24597, 16'd20749, 16'd46664, 16'd54274, 16'd13600, 16'd45200, 16'd19506, 16'd39515, 16'd46363, 16'd40729, 16'd14918, 16'd63117, 16'd19209, 16'd49558, 16'd45590, 16'd64000, 16'd38073, 16'd21980});
	test_expansion(128'hf46296eabbbd50bd3429ec78bceb6353, {16'd34602, 16'd2374, 16'd37416, 16'd50809, 16'd32483, 16'd58782, 16'd30481, 16'd42315, 16'd60006, 16'd45049, 16'd39783, 16'd18582, 16'd41027, 16'd19318, 16'd32048, 16'd58956, 16'd3126, 16'd60528, 16'd37789, 16'd296, 16'd63483, 16'd42618, 16'd16230, 16'd10587, 16'd37061, 16'd58422});
	test_expansion(128'haa08579ee697394b8bbd4fe06b8d8753, {16'd34589, 16'd14729, 16'd56414, 16'd41941, 16'd4133, 16'd61097, 16'd37512, 16'd60379, 16'd32762, 16'd65529, 16'd19249, 16'd35888, 16'd1405, 16'd58782, 16'd5480, 16'd61512, 16'd26726, 16'd50363, 16'd21419, 16'd34655, 16'd16027, 16'd45277, 16'd22630, 16'd62459, 16'd25074, 16'd62354});
	test_expansion(128'he6257c545d7c6c3487d99d57807e614a, {16'd22584, 16'd40959, 16'd13175, 16'd56462, 16'd6303, 16'd33042, 16'd28852, 16'd15352, 16'd45743, 16'd39106, 16'd30533, 16'd30057, 16'd24769, 16'd9696, 16'd33386, 16'd56023, 16'd55559, 16'd64926, 16'd54198, 16'd262, 16'd38176, 16'd38150, 16'd47140, 16'd34899, 16'd18311, 16'd43350});
	test_expansion(128'hbb085232a020f7faa00ff9269bb9d8e6, {16'd20962, 16'd55549, 16'd61238, 16'd27516, 16'd36434, 16'd13560, 16'd35970, 16'd40854, 16'd62260, 16'd61988, 16'd63354, 16'd47468, 16'd7374, 16'd34998, 16'd8231, 16'd65321, 16'd20492, 16'd3669, 16'd12731, 16'd29984, 16'd21600, 16'd36531, 16'd44, 16'd55212, 16'd39433, 16'd65406});
	test_expansion(128'hc3fc9f3117885b3544c1ec5dcd4e6932, {16'd61777, 16'd11434, 16'd31580, 16'd59289, 16'd8351, 16'd46185, 16'd23504, 16'd10199, 16'd37120, 16'd20313, 16'd2219, 16'd41446, 16'd17225, 16'd1238, 16'd21166, 16'd16264, 16'd44959, 16'd54272, 16'd39729, 16'd27543, 16'd37602, 16'd1422, 16'd55792, 16'd5582, 16'd41887, 16'd47864});
	test_expansion(128'h7479524cb4020d518133a6e7a02d1692, {16'd46631, 16'd50406, 16'd63371, 16'd824, 16'd59611, 16'd53256, 16'd47962, 16'd7612, 16'd20338, 16'd38509, 16'd13742, 16'd49255, 16'd39393, 16'd6079, 16'd35075, 16'd50754, 16'd8712, 16'd4843, 16'd42367, 16'd8747, 16'd12782, 16'd54693, 16'd56220, 16'd609, 16'd38366, 16'd12326});
	test_expansion(128'hb2f6f59dca2103a678d8692360781c5c, {16'd15581, 16'd28014, 16'd14404, 16'd17269, 16'd33125, 16'd47653, 16'd61749, 16'd21335, 16'd46601, 16'd33028, 16'd27015, 16'd16590, 16'd5395, 16'd4191, 16'd14017, 16'd58123, 16'd49990, 16'd48850, 16'd56000, 16'd44709, 16'd7266, 16'd28846, 16'd59110, 16'd9752, 16'd2270, 16'd30900});
	test_expansion(128'h55101820d91bf1c089163e89bb94e62e, {16'd35096, 16'd60526, 16'd22218, 16'd13828, 16'd61432, 16'd21465, 16'd5933, 16'd49299, 16'd11576, 16'd48941, 16'd13227, 16'd29710, 16'd20343, 16'd13203, 16'd59871, 16'd3548, 16'd41932, 16'd60186, 16'd55278, 16'd37725, 16'd59390, 16'd53567, 16'd5085, 16'd10592, 16'd38786, 16'd7942});
	test_expansion(128'hd2a56e8222eee29f7f743fcc93eef822, {16'd27314, 16'd54078, 16'd315, 16'd16658, 16'd33575, 16'd30329, 16'd26445, 16'd17613, 16'd52491, 16'd6835, 16'd57754, 16'd22858, 16'd20108, 16'd57340, 16'd2870, 16'd45345, 16'd40228, 16'd64254, 16'd20833, 16'd36838, 16'd34438, 16'd19376, 16'd20501, 16'd36822, 16'd23110, 16'd42162});
	test_expansion(128'hee2daec12931e067ed99ae49e6ce503b, {16'd21947, 16'd51947, 16'd22419, 16'd40865, 16'd16565, 16'd37395, 16'd36153, 16'd128, 16'd63480, 16'd55446, 16'd29886, 16'd7033, 16'd61873, 16'd65136, 16'd44042, 16'd2770, 16'd4099, 16'd2007, 16'd35649, 16'd48382, 16'd37200, 16'd61814, 16'd21668, 16'd25018, 16'd7146, 16'd52406});
	test_expansion(128'he3661aaf1bde1e6dfc7586bbb6f79aae, {16'd62220, 16'd20479, 16'd405, 16'd35535, 16'd22197, 16'd32474, 16'd32874, 16'd10952, 16'd22936, 16'd26904, 16'd45941, 16'd4204, 16'd18783, 16'd9038, 16'd45457, 16'd10655, 16'd458, 16'd33803, 16'd46385, 16'd14948, 16'd34159, 16'd56840, 16'd56929, 16'd2433, 16'd44326, 16'd5778});
	test_expansion(128'hcef7cc5fc33b1afbf8d6f4151d3be7aa, {16'd23475, 16'd32240, 16'd22641, 16'd33270, 16'd17436, 16'd2007, 16'd12691, 16'd3148, 16'd61704, 16'd11910, 16'd15140, 16'd59307, 16'd30958, 16'd58888, 16'd64244, 16'd9167, 16'd53452, 16'd51653, 16'd21001, 16'd50902, 16'd11097, 16'd46260, 16'd28476, 16'd37703, 16'd61922, 16'd31177});
	test_expansion(128'hd33e00c5f79145f0193c1a7bc8227b70, {16'd5797, 16'd7990, 16'd43746, 16'd39422, 16'd21051, 16'd27938, 16'd42223, 16'd26056, 16'd46126, 16'd4736, 16'd47980, 16'd64129, 16'd15414, 16'd44572, 16'd24643, 16'd18667, 16'd54695, 16'd6230, 16'd5242, 16'd8454, 16'd23354, 16'd34322, 16'd24833, 16'd5680, 16'd27910, 16'd37061});
	test_expansion(128'h6c5e68205d286d01deced802a1594c87, {16'd57777, 16'd45841, 16'd49213, 16'd26245, 16'd40946, 16'd43213, 16'd10976, 16'd27785, 16'd22237, 16'd64513, 16'd1452, 16'd28832, 16'd261, 16'd19479, 16'd9000, 16'd47051, 16'd2029, 16'd6900, 16'd11047, 16'd61242, 16'd42884, 16'd61942, 16'd57776, 16'd35864, 16'd20681, 16'd4451});
	test_expansion(128'h5eb95282961740d3a76381b16cf7d198, {16'd22248, 16'd55923, 16'd1877, 16'd39330, 16'd22937, 16'd2332, 16'd4758, 16'd29730, 16'd224, 16'd41003, 16'd15717, 16'd30742, 16'd62137, 16'd15038, 16'd3490, 16'd57956, 16'd40531, 16'd53752, 16'd20275, 16'd14370, 16'd34948, 16'd28926, 16'd5878, 16'd41010, 16'd22037, 16'd6856});
	test_expansion(128'h84e18a327e803ab84f8f03bead5feb2a, {16'd65449, 16'd19121, 16'd24702, 16'd50940, 16'd38779, 16'd16773, 16'd19056, 16'd62998, 16'd29124, 16'd59958, 16'd7228, 16'd34808, 16'd3493, 16'd24035, 16'd63636, 16'd3347, 16'd2651, 16'd41974, 16'd33958, 16'd31354, 16'd20254, 16'd21156, 16'd45574, 16'd39045, 16'd19293, 16'd7086});
	test_expansion(128'h2fe478a240e30518b1789f9a3200a13b, {16'd50445, 16'd2127, 16'd27875, 16'd57471, 16'd31998, 16'd63535, 16'd54659, 16'd57312, 16'd12649, 16'd50463, 16'd60654, 16'd33112, 16'd61436, 16'd4449, 16'd9351, 16'd17960, 16'd45664, 16'd41047, 16'd34687, 16'd44104, 16'd50470, 16'd5154, 16'd30190, 16'd14193, 16'd9388, 16'd695});
	test_expansion(128'h64e91206864642c96b1b724a82a75402, {16'd12607, 16'd5929, 16'd33783, 16'd4017, 16'd57808, 16'd31277, 16'd37407, 16'd20636, 16'd21580, 16'd5916, 16'd56390, 16'd35209, 16'd34793, 16'd13041, 16'd10404, 16'd33097, 16'd35311, 16'd24479, 16'd10387, 16'd34618, 16'd47633, 16'd61172, 16'd52370, 16'd46512, 16'd49207, 16'd52249});
	test_expansion(128'h6317609d6164bf47f1033a5e8e78d452, {16'd38333, 16'd7493, 16'd51292, 16'd54133, 16'd44011, 16'd17354, 16'd33005, 16'd2953, 16'd64175, 16'd27058, 16'd8602, 16'd26164, 16'd18765, 16'd2767, 16'd22314, 16'd48226, 16'd42579, 16'd29072, 16'd5048, 16'd21629, 16'd50404, 16'd48787, 16'd12120, 16'd50089, 16'd19095, 16'd3452});
	test_expansion(128'ha892d0c2328c2fe4cd62b4bc4c8bded7, {16'd32511, 16'd36557, 16'd21207, 16'd41086, 16'd7260, 16'd45374, 16'd54955, 16'd31737, 16'd8779, 16'd4300, 16'd58661, 16'd33645, 16'd11249, 16'd12829, 16'd22947, 16'd16293, 16'd50131, 16'd24295, 16'd45264, 16'd29500, 16'd26697, 16'd34025, 16'd11532, 16'd54129, 16'd45954, 16'd31195});
	test_expansion(128'h647058d9f850869ef5c7cb0c9aadaefe, {16'd64354, 16'd3332, 16'd7451, 16'd43397, 16'd17448, 16'd56164, 16'd21497, 16'd36356, 16'd44777, 16'd61875, 16'd7152, 16'd39951, 16'd62846, 16'd33894, 16'd28257, 16'd23466, 16'd42724, 16'd18164, 16'd45686, 16'd35535, 16'd26271, 16'd6966, 16'd45700, 16'd50118, 16'd13973, 16'd14737});
	test_expansion(128'hbb52cbf29244665571e7589b8058b2ff, {16'd31471, 16'd26083, 16'd17754, 16'd14319, 16'd1688, 16'd49294, 16'd56418, 16'd5016, 16'd52380, 16'd20356, 16'd39137, 16'd49436, 16'd50981, 16'd11251, 16'd26242, 16'd15480, 16'd59002, 16'd11138, 16'd58603, 16'd41686, 16'd42090, 16'd2505, 16'd8760, 16'd37656, 16'd48976, 16'd25650});
	test_expansion(128'h51057db516df7b3c75ad9794065fd17f, {16'd43059, 16'd5492, 16'd30646, 16'd2853, 16'd46442, 16'd33451, 16'd30872, 16'd58226, 16'd51668, 16'd5474, 16'd4398, 16'd34886, 16'd59429, 16'd55255, 16'd46619, 16'd8588, 16'd4676, 16'd9718, 16'd31289, 16'd7144, 16'd23658, 16'd60702, 16'd25828, 16'd51301, 16'd7621, 16'd41850});
	test_expansion(128'hfff607982953da4f1f21795c1755fdce, {16'd36489, 16'd29476, 16'd10528, 16'd29482, 16'd1623, 16'd32663, 16'd56053, 16'd28312, 16'd50057, 16'd22025, 16'd63508, 16'd59703, 16'd20589, 16'd56397, 16'd34877, 16'd11944, 16'd52632, 16'd48894, 16'd44372, 16'd60459, 16'd15128, 16'd39022, 16'd55613, 16'd43781, 16'd1888, 16'd52438});
	test_expansion(128'h98ee9e20c2ec48e46fe45b20cb7648ba, {16'd30192, 16'd51606, 16'd46831, 16'd25273, 16'd43472, 16'd62136, 16'd17708, 16'd6875, 16'd42648, 16'd11728, 16'd40093, 16'd9195, 16'd47258, 16'd26638, 16'd8797, 16'd57899, 16'd26358, 16'd28122, 16'd62820, 16'd43442, 16'd7929, 16'd13014, 16'd50571, 16'd58176, 16'd59353, 16'd51218});
	test_expansion(128'hdd53b56f3cd13c25b6923a577a69371e, {16'd3453, 16'd15439, 16'd12767, 16'd34886, 16'd62936, 16'd58209, 16'd59328, 16'd63271, 16'd50686, 16'd38234, 16'd40182, 16'd35434, 16'd23582, 16'd21692, 16'd7575, 16'd57568, 16'd170, 16'd35421, 16'd6999, 16'd37118, 16'd26578, 16'd41674, 16'd59827, 16'd3806, 16'd11022, 16'd18014});
	test_expansion(128'h1226af3c75769dbabb8767d511667c42, {16'd44033, 16'd18484, 16'd32371, 16'd18663, 16'd35632, 16'd34613, 16'd46090, 16'd63109, 16'd60604, 16'd57197, 16'd28709, 16'd39801, 16'd22281, 16'd7215, 16'd57080, 16'd24998, 16'd12677, 16'd11487, 16'd44597, 16'd58608, 16'd61694, 16'd13939, 16'd53363, 16'd35990, 16'd42900, 16'd844});
	test_expansion(128'h9642b82e88113a30da9cba9278bd0da5, {16'd42918, 16'd45451, 16'd45809, 16'd30687, 16'd55918, 16'd6819, 16'd65246, 16'd27780, 16'd48490, 16'd7902, 16'd1217, 16'd2787, 16'd18164, 16'd21604, 16'd7222, 16'd62244, 16'd48063, 16'd62941, 16'd23192, 16'd54145, 16'd61822, 16'd44474, 16'd52044, 16'd44635, 16'd63765, 16'd21234});
	test_expansion(128'h0b1df25c40dd2b33e0442b39ddd309aa, {16'd18603, 16'd62385, 16'd51423, 16'd38444, 16'd4079, 16'd58321, 16'd16492, 16'd42768, 16'd31715, 16'd59072, 16'd58583, 16'd46431, 16'd37072, 16'd14625, 16'd8313, 16'd48759, 16'd44986, 16'd61168, 16'd23022, 16'd7582, 16'd2058, 16'd51379, 16'd488, 16'd50645, 16'd54686, 16'd14244});
	test_expansion(128'h78f66b150c8f7c0583707ad881ffaf5c, {16'd55928, 16'd30595, 16'd40006, 16'd23088, 16'd16350, 16'd18512, 16'd35628, 16'd50468, 16'd11035, 16'd8370, 16'd38898, 16'd24158, 16'd47645, 16'd28993, 16'd30975, 16'd613, 16'd2656, 16'd54495, 16'd26917, 16'd357, 16'd28867, 16'd33787, 16'd43117, 16'd11752, 16'd14006, 16'd63433});
	test_expansion(128'h09a4a66367b6ab47535fe50b6bef9a0e, {16'd42386, 16'd22251, 16'd60650, 16'd43194, 16'd4716, 16'd22165, 16'd29384, 16'd14265, 16'd65152, 16'd26832, 16'd8721, 16'd57478, 16'd50987, 16'd17801, 16'd31350, 16'd46467, 16'd52959, 16'd8598, 16'd17747, 16'd17489, 16'd29666, 16'd33070, 16'd48635, 16'd56586, 16'd61666, 16'd2827});
	test_expansion(128'h5b4384d0fad0ae3f0df2b8e3db9f25e1, {16'd26711, 16'd9170, 16'd34489, 16'd11051, 16'd47012, 16'd46152, 16'd64615, 16'd51019, 16'd47070, 16'd51011, 16'd59951, 16'd14536, 16'd16528, 16'd28227, 16'd40784, 16'd63, 16'd641, 16'd61843, 16'd22742, 16'd45161, 16'd523, 16'd61170, 16'd37018, 16'd12958, 16'd4107, 16'd51067});
	test_expansion(128'h361040b19454e00b2bdfcb859ad2e5ec, {16'd54010, 16'd64567, 16'd60169, 16'd60118, 16'd47989, 16'd23948, 16'd44991, 16'd54868, 16'd3449, 16'd39528, 16'd13468, 16'd23145, 16'd40142, 16'd26665, 16'd16015, 16'd55965, 16'd64730, 16'd12795, 16'd47947, 16'd54083, 16'd65336, 16'd40518, 16'd13882, 16'd25494, 16'd18547, 16'd32647});
	test_expansion(128'he08ff24a7bbb8e307a84555a16b26d71, {16'd2490, 16'd45943, 16'd2516, 16'd46574, 16'd16670, 16'd55202, 16'd39296, 16'd11767, 16'd35919, 16'd42362, 16'd32218, 16'd48069, 16'd27968, 16'd14897, 16'd43966, 16'd15510, 16'd27806, 16'd55754, 16'd8070, 16'd15035, 16'd8998, 16'd63205, 16'd28060, 16'd36216, 16'd64098, 16'd6967});
	test_expansion(128'hbf668885b3a4be507af7731b5730bceb, {16'd17117, 16'd40767, 16'd43227, 16'd52678, 16'd7913, 16'd4780, 16'd29342, 16'd29363, 16'd55250, 16'd10789, 16'd42043, 16'd56475, 16'd41247, 16'd11979, 16'd42207, 16'd25173, 16'd24845, 16'd55319, 16'd30377, 16'd17361, 16'd51306, 16'd25400, 16'd27799, 16'd44625, 16'd37172, 16'd39920});
	test_expansion(128'h95b582dec28f15dd5f04075318725087, {16'd56259, 16'd28832, 16'd23968, 16'd2623, 16'd22932, 16'd53636, 16'd54342, 16'd37302, 16'd37262, 16'd49701, 16'd9830, 16'd12247, 16'd37367, 16'd2536, 16'd39021, 16'd23918, 16'd32408, 16'd47264, 16'd61293, 16'd14795, 16'd40122, 16'd45490, 16'd50531, 16'd9804, 16'd6624, 16'd63837});
	test_expansion(128'h5ce561a35187b1058c34652dac70a50e, {16'd64104, 16'd6945, 16'd29462, 16'd42890, 16'd54057, 16'd14973, 16'd57408, 16'd32927, 16'd455, 16'd5979, 16'd40409, 16'd56310, 16'd19648, 16'd53903, 16'd31936, 16'd1146, 16'd16723, 16'd64871, 16'd47375, 16'd53780, 16'd32398, 16'd16180, 16'd60644, 16'd42890, 16'd63702, 16'd37569});
	test_expansion(128'h48975ff2124c6d1e1a4eb7a66864be19, {16'd12718, 16'd19436, 16'd9294, 16'd61405, 16'd36382, 16'd59769, 16'd45486, 16'd41689, 16'd17623, 16'd10926, 16'd22576, 16'd45996, 16'd52390, 16'd55057, 16'd4974, 16'd36171, 16'd53268, 16'd45504, 16'd298, 16'd56529, 16'd45028, 16'd10550, 16'd7846, 16'd44140, 16'd40144, 16'd27257});
	test_expansion(128'he079a01364186373fd27cf07edded9c2, {16'd41172, 16'd21891, 16'd5963, 16'd45173, 16'd1320, 16'd3863, 16'd27579, 16'd33330, 16'd55237, 16'd35169, 16'd10808, 16'd30391, 16'd64830, 16'd16076, 16'd21144, 16'd53651, 16'd23661, 16'd60611, 16'd63624, 16'd64996, 16'd27364, 16'd61398, 16'd33150, 16'd42245, 16'd55315, 16'd21604});
	test_expansion(128'h88bdebddbf1390ae503dc677f46a8bf6, {16'd26030, 16'd31362, 16'd58917, 16'd51755, 16'd63257, 16'd51557, 16'd60008, 16'd3874, 16'd31530, 16'd59723, 16'd44189, 16'd39064, 16'd12042, 16'd53273, 16'd3764, 16'd13581, 16'd15679, 16'd37122, 16'd44411, 16'd58014, 16'd40477, 16'd35176, 16'd61891, 16'd9690, 16'd50929, 16'd24520});
	test_expansion(128'h0c7f0be7e191ff5cd7a3301f1a057ef2, {16'd33548, 16'd39051, 16'd16038, 16'd50760, 16'd26603, 16'd63752, 16'd60306, 16'd7711, 16'd12658, 16'd25394, 16'd46847, 16'd14369, 16'd39788, 16'd41191, 16'd33685, 16'd56288, 16'd2939, 16'd65092, 16'd12448, 16'd7729, 16'd47584, 16'd52831, 16'd13811, 16'd46150, 16'd38818, 16'd27140});
	test_expansion(128'haebce2b0313526e3de5697bcfc411247, {16'd57678, 16'd1130, 16'd16425, 16'd22976, 16'd51415, 16'd48657, 16'd27246, 16'd28179, 16'd55243, 16'd43912, 16'd60958, 16'd358, 16'd34782, 16'd64536, 16'd33962, 16'd57426, 16'd36485, 16'd37781, 16'd44242, 16'd43137, 16'd2279, 16'd48743, 16'd5862, 16'd57654, 16'd20661, 16'd1905});
	test_expansion(128'h18fb2a34118247925143c05d9a1ccabe, {16'd38048, 16'd31528, 16'd15865, 16'd51197, 16'd26039, 16'd21541, 16'd52983, 16'd35991, 16'd55480, 16'd32487, 16'd10816, 16'd17338, 16'd32567, 16'd23490, 16'd38934, 16'd8184, 16'd24624, 16'd49337, 16'd5237, 16'd53070, 16'd20325, 16'd48542, 16'd59857, 16'd14182, 16'd36974, 16'd32879});
	test_expansion(128'he73621f06d24e3d75854691bc6bff62b, {16'd36434, 16'd3448, 16'd11698, 16'd36720, 16'd33724, 16'd55466, 16'd3619, 16'd51060, 16'd37571, 16'd35345, 16'd49016, 16'd53570, 16'd702, 16'd9262, 16'd37668, 16'd36028, 16'd29738, 16'd36867, 16'd64109, 16'd9400, 16'd37110, 16'd3518, 16'd28320, 16'd41520, 16'd33765, 16'd54524});
	test_expansion(128'hc044d6b435522a6954272e1cc0141ff6, {16'd30710, 16'd12270, 16'd16015, 16'd96, 16'd47473, 16'd53265, 16'd36110, 16'd21610, 16'd55603, 16'd490, 16'd56008, 16'd45617, 16'd47354, 16'd45950, 16'd63644, 16'd63348, 16'd64817, 16'd39065, 16'd17713, 16'd3633, 16'd19865, 16'd25009, 16'd51938, 16'd1303, 16'd44006, 16'd28552});
	test_expansion(128'ha5e58bdc241611b0a33b3157d9f8652d, {16'd50787, 16'd61912, 16'd22133, 16'd34102, 16'd64111, 16'd703, 16'd28520, 16'd6166, 16'd2784, 16'd61386, 16'd9830, 16'd63929, 16'd6816, 16'd2943, 16'd2359, 16'd45110, 16'd15516, 16'd39452, 16'd9354, 16'd7794, 16'd29644, 16'd19041, 16'd37969, 16'd52129, 16'd45682, 16'd49252});
	test_expansion(128'h3c1bc6d62561878699c6713fd408a0e2, {16'd10267, 16'd39716, 16'd36739, 16'd16345, 16'd35210, 16'd5125, 16'd26408, 16'd53634, 16'd6568, 16'd23496, 16'd47870, 16'd51287, 16'd37761, 16'd7527, 16'd36338, 16'd11627, 16'd42510, 16'd1447, 16'd44461, 16'd40751, 16'd18017, 16'd27443, 16'd43217, 16'd27929, 16'd6261, 16'd27671});
	test_expansion(128'hf5fac558bb3a59ff7db6bbc4eb308e9e, {16'd2120, 16'd47413, 16'd6496, 16'd13995, 16'd41232, 16'd18954, 16'd62540, 16'd40463, 16'd12492, 16'd54429, 16'd60781, 16'd33503, 16'd21404, 16'd19917, 16'd46888, 16'd13676, 16'd29171, 16'd28065, 16'd56644, 16'd47154, 16'd53430, 16'd45513, 16'd49738, 16'd18041, 16'd39207, 16'd64573});
	test_expansion(128'h76b649c6a0d4942aab2d5e4d0e25a7f1, {16'd10198, 16'd25856, 16'd44431, 16'd16296, 16'd5516, 16'd11251, 16'd57323, 16'd7924, 16'd30843, 16'd13623, 16'd15672, 16'd63001, 16'd29467, 16'd62953, 16'd31601, 16'd25473, 16'd26002, 16'd26193, 16'd41455, 16'd2326, 16'd30629, 16'd29304, 16'd30492, 16'd5352, 16'd2591, 16'd58250});
	test_expansion(128'h25068c0e51772e3f991c4b00bf0c7b71, {16'd11486, 16'd30447, 16'd5197, 16'd42603, 16'd21842, 16'd25145, 16'd13613, 16'd50627, 16'd51103, 16'd33424, 16'd19699, 16'd36643, 16'd30961, 16'd40611, 16'd59833, 16'd58932, 16'd13403, 16'd7322, 16'd64810, 16'd22934, 16'd22998, 16'd47916, 16'd60547, 16'd43294, 16'd10556, 16'd63451});
	test_expansion(128'h652de4c94748a2ac3110e485943a6ce3, {16'd5616, 16'd9588, 16'd33756, 16'd15950, 16'd41892, 16'd17570, 16'd61460, 16'd36534, 16'd16077, 16'd7524, 16'd14903, 16'd64581, 16'd63595, 16'd17174, 16'd38884, 16'd46315, 16'd5007, 16'd729, 16'd40044, 16'd63988, 16'd794, 16'd26802, 16'd58852, 16'd8454, 16'd8681, 16'd25279});
	test_expansion(128'hc3dbc13088546c821545e19977ccb889, {16'd32380, 16'd23520, 16'd43270, 16'd45672, 16'd9824, 16'd61291, 16'd58054, 16'd672, 16'd1962, 16'd37419, 16'd52427, 16'd29012, 16'd45849, 16'd36362, 16'd5497, 16'd26287, 16'd22129, 16'd34117, 16'd35618, 16'd50008, 16'd18698, 16'd24889, 16'd50767, 16'd47250, 16'd29251, 16'd24806});
	test_expansion(128'h47845f46df196aacbde5edb9628a3259, {16'd27045, 16'd164, 16'd20901, 16'd33553, 16'd23082, 16'd28896, 16'd63475, 16'd25408, 16'd46985, 16'd12415, 16'd9913, 16'd31716, 16'd55275, 16'd29617, 16'd45286, 16'd26431, 16'd63259, 16'd40716, 16'd26867, 16'd5506, 16'd37929, 16'd60398, 16'd55187, 16'd31376, 16'd26989, 16'd29998});
	test_expansion(128'hda27a548b1857069ef64559177ee23d5, {16'd3741, 16'd1456, 16'd15356, 16'd1314, 16'd2128, 16'd27602, 16'd62262, 16'd46228, 16'd15440, 16'd22316, 16'd25034, 16'd11482, 16'd14979, 16'd21332, 16'd56256, 16'd24087, 16'd32288, 16'd57147, 16'd27991, 16'd17747, 16'd1602, 16'd14028, 16'd13935, 16'd27829, 16'd64244, 16'd19924});
	test_expansion(128'hb28582ac2be0b864cb753701dc2ad916, {16'd56467, 16'd24864, 16'd39756, 16'd59913, 16'd22269, 16'd8175, 16'd6666, 16'd10411, 16'd46778, 16'd17166, 16'd8433, 16'd1131, 16'd57932, 16'd28349, 16'd28832, 16'd44663, 16'd12022, 16'd39524, 16'd31488, 16'd54358, 16'd31847, 16'd8025, 16'd59005, 16'd39083, 16'd39931, 16'd65189});
	test_expansion(128'h93a4cea7031978c2d1f4da1301143d99, {16'd16014, 16'd43428, 16'd38932, 16'd50076, 16'd2508, 16'd46597, 16'd39388, 16'd42920, 16'd43364, 16'd45823, 16'd34448, 16'd52592, 16'd64503, 16'd43440, 16'd54960, 16'd55860, 16'd32458, 16'd27393, 16'd50396, 16'd17374, 16'd60750, 16'd10851, 16'd17402, 16'd55136, 16'd37602, 16'd52435});
	test_expansion(128'hdc1212475723030f6cf733698d181f27, {16'd22955, 16'd38072, 16'd21216, 16'd21057, 16'd50125, 16'd8896, 16'd61275, 16'd15300, 16'd26755, 16'd40265, 16'd46615, 16'd48037, 16'd37224, 16'd51720, 16'd51063, 16'd58219, 16'd29205, 16'd36351, 16'd52186, 16'd40342, 16'd12284, 16'd40774, 16'd48902, 16'd56226, 16'd17594, 16'd39256});
	test_expansion(128'hcf415fdd834958a924b2c70292c5ed7c, {16'd40352, 16'd64907, 16'd52164, 16'd25671, 16'd4050, 16'd37015, 16'd7878, 16'd9804, 16'd17547, 16'd23714, 16'd38943, 16'd25984, 16'd19357, 16'd25682, 16'd17324, 16'd59479, 16'd29206, 16'd5933, 16'd56868, 16'd57394, 16'd42603, 16'd57853, 16'd10125, 16'd35093, 16'd20887, 16'd5044});
	test_expansion(128'h377810a14385cb283aa649e9902558ec, {16'd13107, 16'd2780, 16'd22038, 16'd42726, 16'd40879, 16'd11711, 16'd24875, 16'd32784, 16'd54130, 16'd58689, 16'd46958, 16'd53125, 16'd37889, 16'd51794, 16'd30891, 16'd42609, 16'd53808, 16'd10798, 16'd15406, 16'd36396, 16'd39107, 16'd63872, 16'd12113, 16'd47154, 16'd63943, 16'd3684});
	test_expansion(128'h9be4b7376018a986b05456a7e2e42c60, {16'd4479, 16'd19450, 16'd32582, 16'd22060, 16'd19684, 16'd12824, 16'd32218, 16'd15465, 16'd40948, 16'd36456, 16'd46800, 16'd31089, 16'd13770, 16'd16001, 16'd28035, 16'd32505, 16'd26072, 16'd28891, 16'd65172, 16'd21460, 16'd61903, 16'd28246, 16'd54254, 16'd51061, 16'd6864, 16'd45030});
	test_expansion(128'habc3210215f591976b3d69b47811240c, {16'd28933, 16'd23580, 16'd28549, 16'd34040, 16'd54597, 16'd40212, 16'd43080, 16'd28116, 16'd27220, 16'd1455, 16'd57672, 16'd54596, 16'd38162, 16'd53158, 16'd55526, 16'd40604, 16'd47033, 16'd13468, 16'd7946, 16'd60000, 16'd50468, 16'd54191, 16'd22548, 16'd12466, 16'd14154, 16'd6519});
	test_expansion(128'hc7f7323c7b7b3dfba91f5bd798caec8b, {16'd3880, 16'd14668, 16'd1568, 16'd31899, 16'd28717, 16'd37049, 16'd60761, 16'd16114, 16'd10687, 16'd53197, 16'd11129, 16'd61779, 16'd14856, 16'd34110, 16'd6940, 16'd133, 16'd21882, 16'd20700, 16'd42038, 16'd1750, 16'd45576, 16'd52413, 16'd42066, 16'd47155, 16'd6164, 16'd28894});
	test_expansion(128'h583133091a9097350916e9ce73e40d1d, {16'd10817, 16'd27553, 16'd24089, 16'd56057, 16'd32505, 16'd8267, 16'd46094, 16'd611, 16'd49377, 16'd53559, 16'd16787, 16'd12970, 16'd52873, 16'd40039, 16'd63074, 16'd46430, 16'd65039, 16'd61649, 16'd56597, 16'd13305, 16'd19136, 16'd35341, 16'd65065, 16'd35531, 16'd50698, 16'd60986});
	test_expansion(128'hd991060b08a8a30762511e2ed5473e4b, {16'd47257, 16'd58396, 16'd60810, 16'd31014, 16'd27605, 16'd34249, 16'd22310, 16'd16426, 16'd37429, 16'd37277, 16'd10618, 16'd17398, 16'd30627, 16'd31824, 16'd61355, 16'd25477, 16'd10194, 16'd25876, 16'd62970, 16'd48418, 16'd11851, 16'd41439, 16'd16684, 16'd18198, 16'd25050, 16'd12067});
	test_expansion(128'heaf9bcc5058cb501637336c1a6184c5c, {16'd10725, 16'd5425, 16'd13334, 16'd39265, 16'd4244, 16'd17772, 16'd60624, 16'd46019, 16'd49078, 16'd63951, 16'd42705, 16'd18132, 16'd11074, 16'd23736, 16'd36098, 16'd48926, 16'd54337, 16'd59580, 16'd37796, 16'd46226, 16'd14665, 16'd62774, 16'd47112, 16'd30467, 16'd43476, 16'd25633});
	test_expansion(128'hab209e67d987c4b423e656a6a290c612, {16'd5898, 16'd18756, 16'd58998, 16'd23423, 16'd38139, 16'd64975, 16'd58797, 16'd35678, 16'd53977, 16'd33701, 16'd7677, 16'd27541, 16'd28030, 16'd41837, 16'd20647, 16'd4082, 16'd35268, 16'd40105, 16'd40660, 16'd38124, 16'd9778, 16'd38545, 16'd32500, 16'd57025, 16'd11226, 16'd62884});
	test_expansion(128'h1c8a8aff6fcbcdf3d7863332b1ca1c32, {16'd23866, 16'd906, 16'd12395, 16'd25706, 16'd65373, 16'd54093, 16'd55792, 16'd39279, 16'd16815, 16'd4031, 16'd58681, 16'd43928, 16'd34741, 16'd21644, 16'd27973, 16'd25788, 16'd19333, 16'd52984, 16'd21031, 16'd18512, 16'd8245, 16'd27735, 16'd51781, 16'd10230, 16'd25386, 16'd25522});
	test_expansion(128'hc0a5168f546b0fd1e5d4acb41418a752, {16'd42162, 16'd57445, 16'd57130, 16'd9167, 16'd502, 16'd58425, 16'd55907, 16'd39792, 16'd53226, 16'd42844, 16'd56849, 16'd46283, 16'd17873, 16'd44253, 16'd41026, 16'd36442, 16'd9186, 16'd24799, 16'd28054, 16'd26789, 16'd10946, 16'd28022, 16'd39368, 16'd63429, 16'd56689, 16'd35174});
	test_expansion(128'h05f4be14fb55cfb34d59680a79b1d7c6, {16'd29374, 16'd43990, 16'd62400, 16'd53526, 16'd46801, 16'd46956, 16'd23747, 16'd33786, 16'd24001, 16'd54910, 16'd10784, 16'd45880, 16'd54460, 16'd38704, 16'd20298, 16'd21821, 16'd37469, 16'd11036, 16'd12898, 16'd21338, 16'd15202, 16'd1633, 16'd15027, 16'd59770, 16'd58812, 16'd52636});
	test_expansion(128'hf3346beb67e185690ec327e84d26ab54, {16'd1804, 16'd37016, 16'd1220, 16'd21885, 16'd48399, 16'd23035, 16'd26723, 16'd9388, 16'd62022, 16'd26615, 16'd52689, 16'd11731, 16'd24795, 16'd51629, 16'd22258, 16'd16375, 16'd33489, 16'd50974, 16'd6848, 16'd45465, 16'd52892, 16'd33132, 16'd13064, 16'd27751, 16'd6651, 16'd5680});
	test_expansion(128'ha1cf2996c9f2bd4cedd189659727c15e, {16'd56741, 16'd28726, 16'd22469, 16'd3781, 16'd32173, 16'd4496, 16'd24317, 16'd19942, 16'd27089, 16'd33127, 16'd15486, 16'd49455, 16'd48740, 16'd13927, 16'd22295, 16'd7739, 16'd53974, 16'd9853, 16'd61408, 16'd22348, 16'd27515, 16'd1955, 16'd42339, 16'd8434, 16'd39821, 16'd38215});
	test_expansion(128'hcbfeeb5a6e785e81fc7cc269d7d03e09, {16'd52822, 16'd8185, 16'd53418, 16'd59612, 16'd35882, 16'd51974, 16'd61095, 16'd13302, 16'd47289, 16'd28865, 16'd56845, 16'd28222, 16'd55648, 16'd65014, 16'd53254, 16'd51090, 16'd27377, 16'd47395, 16'd10372, 16'd64421, 16'd17358, 16'd12760, 16'd65072, 16'd1722, 16'd4150, 16'd47038});
	test_expansion(128'h8cbad5967f3e5abd72bb244a0ab1a409, {16'd51100, 16'd36152, 16'd21814, 16'd44310, 16'd3111, 16'd7822, 16'd19906, 16'd12954, 16'd28479, 16'd61744, 16'd32788, 16'd3932, 16'd4703, 16'd31931, 16'd15504, 16'd50676, 16'd53230, 16'd24616, 16'd37208, 16'd25558, 16'd29517, 16'd8735, 16'd46130, 16'd43670, 16'd18999, 16'd37581});
	test_expansion(128'h57fe4f769ba8866157851c42450c1971, {16'd30537, 16'd50410, 16'd53339, 16'd55907, 16'd19489, 16'd8046, 16'd37960, 16'd60854, 16'd54439, 16'd38487, 16'd43053, 16'd64011, 16'd217, 16'd11711, 16'd42386, 16'd6179, 16'd18337, 16'd60123, 16'd59128, 16'd48905, 16'd4031, 16'd6754, 16'd53041, 16'd18209, 16'd21580, 16'd50909});
	test_expansion(128'h39189d80c121d1e73e29e8428eec7ecc, {16'd14014, 16'd35141, 16'd14730, 16'd33456, 16'd44512, 16'd39991, 16'd22480, 16'd39197, 16'd56392, 16'd59393, 16'd50230, 16'd59144, 16'd19603, 16'd7608, 16'd21941, 16'd64873, 16'd28137, 16'd7007, 16'd45692, 16'd26020, 16'd43027, 16'd5834, 16'd16252, 16'd8688, 16'd47075, 16'd48771});
	test_expansion(128'h0a9d441e731d0ee400a3e823a4ea9bb9, {16'd63246, 16'd5110, 16'd41899, 16'd52106, 16'd43013, 16'd10970, 16'd16975, 16'd15755, 16'd6824, 16'd14023, 16'd30351, 16'd30322, 16'd15516, 16'd28209, 16'd27323, 16'd64806, 16'd6299, 16'd55103, 16'd62106, 16'd58631, 16'd15494, 16'd34622, 16'd6903, 16'd19646, 16'd49935, 16'd31599});
	test_expansion(128'hc415834c532eb5cf3da3544bf1c40344, {16'd55697, 16'd39810, 16'd27578, 16'd53565, 16'd20351, 16'd35193, 16'd8910, 16'd45392, 16'd52003, 16'd33562, 16'd53285, 16'd55821, 16'd48503, 16'd20702, 16'd49681, 16'd37813, 16'd8883, 16'd12116, 16'd50038, 16'd3412, 16'd34454, 16'd36678, 16'd34068, 16'd36601, 16'd28557, 16'd54893});
	test_expansion(128'h7f867307c05af7e8c2e8aebe591607d0, {16'd34144, 16'd3983, 16'd41875, 16'd39931, 16'd34741, 16'd12429, 16'd42040, 16'd63912, 16'd35503, 16'd9252, 16'd22288, 16'd657, 16'd20648, 16'd22067, 16'd14929, 16'd49664, 16'd64251, 16'd54131, 16'd19837, 16'd53559, 16'd20996, 16'd55980, 16'd62896, 16'd61136, 16'd4164, 16'd52890});
	test_expansion(128'ha0c65488c052659be2f9a598373989c9, {16'd9686, 16'd19908, 16'd613, 16'd22702, 16'd22068, 16'd63883, 16'd37335, 16'd6215, 16'd63873, 16'd49018, 16'd57245, 16'd33932, 16'd59237, 16'd64364, 16'd63404, 16'd64995, 16'd12300, 16'd15777, 16'd49346, 16'd20455, 16'd4024, 16'd37991, 16'd48479, 16'd14332, 16'd14127, 16'd12413});
	test_expansion(128'h4353ec64148e9a09be5831811610f08d, {16'd38772, 16'd15711, 16'd44261, 16'd29597, 16'd14431, 16'd56683, 16'd10455, 16'd44824, 16'd43557, 16'd12496, 16'd30063, 16'd10924, 16'd4622, 16'd25501, 16'd20703, 16'd58256, 16'd59601, 16'd42089, 16'd35746, 16'd14682, 16'd12821, 16'd54798, 16'd54746, 16'd45029, 16'd58349, 16'd7971});
	test_expansion(128'h2ec8afae50fe35bb978a1f234fd21c3a, {16'd8365, 16'd62639, 16'd8246, 16'd10046, 16'd29595, 16'd22353, 16'd54014, 16'd56318, 16'd21198, 16'd22181, 16'd31828, 16'd60946, 16'd33851, 16'd22748, 16'd49271, 16'd9183, 16'd56978, 16'd21519, 16'd60846, 16'd29677, 16'd51274, 16'd7858, 16'd35814, 16'd37288, 16'd40698, 16'd64291});
	test_expansion(128'h02703028ced6a8974cb5bbdecaae86fc, {16'd24655, 16'd58358, 16'd58755, 16'd60754, 16'd11769, 16'd46051, 16'd61312, 16'd22215, 16'd27317, 16'd4144, 16'd8292, 16'd45651, 16'd41954, 16'd58707, 16'd27246, 16'd12794, 16'd57165, 16'd62374, 16'd13842, 16'd13710, 16'd56966, 16'd57327, 16'd15543, 16'd49808, 16'd23078, 16'd54492});
	test_expansion(128'h018004316b01798c8417e9e2c10c0841, {16'd53311, 16'd12683, 16'd8143, 16'd63086, 16'd380, 16'd13901, 16'd30001, 16'd36108, 16'd35712, 16'd35313, 16'd21578, 16'd43115, 16'd40, 16'd28122, 16'd29028, 16'd16792, 16'd8727, 16'd48280, 16'd10611, 16'd8172, 16'd13665, 16'd25982, 16'd3672, 16'd393, 16'd58401, 16'd53539});
	test_expansion(128'h22dc1b438785fdc3ed80cc276427259e, {16'd8745, 16'd4932, 16'd21429, 16'd42040, 16'd19794, 16'd13050, 16'd10087, 16'd3398, 16'd42505, 16'd13167, 16'd3554, 16'd47520, 16'd20404, 16'd20767, 16'd18303, 16'd24871, 16'd4653, 16'd21356, 16'd48989, 16'd55026, 16'd41086, 16'd27876, 16'd33559, 16'd38635, 16'd56192, 16'd16669});
	test_expansion(128'hb955530c7a473162f27a7a88fc3175d0, {16'd32491, 16'd60303, 16'd24592, 16'd38286, 16'd57461, 16'd55409, 16'd27143, 16'd45596, 16'd45022, 16'd54400, 16'd62385, 16'd496, 16'd47901, 16'd25398, 16'd54500, 16'd55847, 16'd28860, 16'd30217, 16'd27774, 16'd62750, 16'd32171, 16'd40850, 16'd57041, 16'd34296, 16'd13238, 16'd58469});
	test_expansion(128'h82b7296c5d1de67698715071b5356403, {16'd45917, 16'd55444, 16'd42034, 16'd34365, 16'd14005, 16'd30554, 16'd8959, 16'd52880, 16'd17463, 16'd7539, 16'd34765, 16'd40257, 16'd8459, 16'd50874, 16'd11395, 16'd42335, 16'd21888, 16'd30281, 16'd39088, 16'd19092, 16'd25788, 16'd52165, 16'd55195, 16'd49426, 16'd2366, 16'd18150});
	test_expansion(128'hf7e8d08763e702f5c43d8e82fc1c770a, {16'd52551, 16'd57546, 16'd52444, 16'd34830, 16'd54063, 16'd59415, 16'd49261, 16'd15859, 16'd3165, 16'd12360, 16'd55317, 16'd32996, 16'd16235, 16'd34889, 16'd38649, 16'd47803, 16'd36846, 16'd24158, 16'd50246, 16'd22373, 16'd12561, 16'd14296, 16'd27850, 16'd33193, 16'd24101, 16'd8330});
	test_expansion(128'h96b60ae7b553ffc51006ce7b2e17faba, {16'd33452, 16'd8625, 16'd14642, 16'd40149, 16'd47948, 16'd33692, 16'd1174, 16'd47173, 16'd42762, 16'd11492, 16'd64358, 16'd47764, 16'd29510, 16'd32625, 16'd31244, 16'd29291, 16'd17759, 16'd35773, 16'd35216, 16'd49380, 16'd843, 16'd49671, 16'd10302, 16'd51918, 16'd33695, 16'd36497});
	test_expansion(128'hf83c292d9ae55fe7c7747b64956fff55, {16'd5894, 16'd47633, 16'd55215, 16'd12179, 16'd54156, 16'd65213, 16'd9142, 16'd9080, 16'd48989, 16'd59640, 16'd50356, 16'd63724, 16'd10763, 16'd55633, 16'd22761, 16'd56833, 16'd23697, 16'd59603, 16'd28099, 16'd41762, 16'd49253, 16'd20925, 16'd3364, 16'd9025, 16'd37152, 16'd1643});
	test_expansion(128'h47d5e93a96f9ed62e40a871eaf638a73, {16'd49597, 16'd52964, 16'd58322, 16'd31941, 16'd8400, 16'd21640, 16'd38011, 16'd42131, 16'd57601, 16'd58913, 16'd62741, 16'd38060, 16'd7365, 16'd21055, 16'd39401, 16'd24218, 16'd34237, 16'd19918, 16'd60281, 16'd61023, 16'd33728, 16'd61754, 16'd58411, 16'd19321, 16'd53381, 16'd65530});
	test_expansion(128'hea3943137a490cfd2f98969a51fcea99, {16'd47279, 16'd37012, 16'd22948, 16'd19163, 16'd44111, 16'd16367, 16'd10290, 16'd64947, 16'd46075, 16'd45566, 16'd7203, 16'd22858, 16'd13959, 16'd61446, 16'd63320, 16'd9195, 16'd15175, 16'd29334, 16'd506, 16'd43075, 16'd18975, 16'd25999, 16'd43056, 16'd9404, 16'd3718, 16'd49151});
	test_expansion(128'h1d97468993d715ae4bc64311cb20b947, {16'd53816, 16'd32617, 16'd8604, 16'd31385, 16'd53139, 16'd57204, 16'd9220, 16'd23707, 16'd53702, 16'd31120, 16'd29366, 16'd21148, 16'd54170, 16'd22039, 16'd36634, 16'd41918, 16'd9710, 16'd4388, 16'd63957, 16'd45022, 16'd63694, 16'd35983, 16'd19528, 16'd8583, 16'd21858, 16'd38168});
	test_expansion(128'ha82bf0a5764e4fd090fcb47fa7232e7e, {16'd56539, 16'd58436, 16'd43722, 16'd28982, 16'd11285, 16'd58360, 16'd56024, 16'd4064, 16'd50400, 16'd42, 16'd9807, 16'd4975, 16'd38958, 16'd9500, 16'd18308, 16'd51170, 16'd59319, 16'd11757, 16'd52969, 16'd18103, 16'd44588, 16'd27543, 16'd32479, 16'd25922, 16'd26704, 16'd30824});
	test_expansion(128'h4e8283ca4878a1c9a6977c76363d8a84, {16'd30023, 16'd11591, 16'd62003, 16'd3602, 16'd24376, 16'd29246, 16'd39942, 16'd57496, 16'd728, 16'd45308, 16'd12136, 16'd42160, 16'd31057, 16'd49026, 16'd40045, 16'd36470, 16'd10113, 16'd9918, 16'd47197, 16'd36893, 16'd62933, 16'd54877, 16'd18625, 16'd41028, 16'd5561, 16'd17371});
	test_expansion(128'hf795865a89e4df906daffdfe12874e82, {16'd6935, 16'd20792, 16'd22220, 16'd61290, 16'd10726, 16'd205, 16'd36664, 16'd26911, 16'd32513, 16'd46225, 16'd62441, 16'd49897, 16'd63001, 16'd55062, 16'd26175, 16'd23626, 16'd40359, 16'd54709, 16'd18060, 16'd11536, 16'd45595, 16'd55629, 16'd59062, 16'd34634, 16'd39892, 16'd32450});
	test_expansion(128'he02db3aa2d5d0d5a502bc3aeaa35c8b5, {16'd65374, 16'd52617, 16'd15127, 16'd15055, 16'd47795, 16'd17739, 16'd61326, 16'd18058, 16'd45465, 16'd54917, 16'd47288, 16'd63336, 16'd43368, 16'd41420, 16'd8950, 16'd51388, 16'd22109, 16'd38668, 16'd20538, 16'd51458, 16'd51888, 16'd53075, 16'd9004, 16'd20601, 16'd5786, 16'd36343});
	test_expansion(128'h51a0ed85fe1593f6bf08293e9fb7754d, {16'd9687, 16'd35207, 16'd52656, 16'd245, 16'd25234, 16'd19142, 16'd17016, 16'd23336, 16'd38388, 16'd26178, 16'd48902, 16'd35291, 16'd36011, 16'd49987, 16'd16314, 16'd37253, 16'd10007, 16'd38076, 16'd10054, 16'd23582, 16'd63442, 16'd35371, 16'd61603, 16'd17283, 16'd61006, 16'd53030});
	test_expansion(128'h9dd8636a3433b3d028781359fb7ba13d, {16'd50654, 16'd63098, 16'd577, 16'd60468, 16'd3343, 16'd18221, 16'd48175, 16'd19587, 16'd63382, 16'd8960, 16'd25660, 16'd60585, 16'd36942, 16'd65215, 16'd60312, 16'd43587, 16'd42267, 16'd25724, 16'd7053, 16'd41129, 16'd13919, 16'd33300, 16'd25423, 16'd5676, 16'd9869, 16'd36916});
	test_expansion(128'h2da8d55d8034698ffd8c2ec702dc488c, {16'd2417, 16'd42364, 16'd48406, 16'd9240, 16'd55619, 16'd54632, 16'd47822, 16'd45842, 16'd45195, 16'd37995, 16'd8436, 16'd20751, 16'd22818, 16'd33361, 16'd47431, 16'd10069, 16'd61965, 16'd54310, 16'd61339, 16'd61613, 16'd10982, 16'd24725, 16'd26846, 16'd56546, 16'd1976, 16'd55656});
	test_expansion(128'h51336cad55f2e41fe2278f330c7ab707, {16'd41686, 16'd6399, 16'd4941, 16'd11214, 16'd860, 16'd42479, 16'd5888, 16'd49061, 16'd56161, 16'd23533, 16'd53479, 16'd13890, 16'd28469, 16'd32549, 16'd43395, 16'd60899, 16'd45347, 16'd8598, 16'd41882, 16'd13939, 16'd52736, 16'd48942, 16'd58648, 16'd55991, 16'd53339, 16'd64303});
	test_expansion(128'hd63774bd8eaa3a9e6595208b6c67d3ca, {16'd38510, 16'd48675, 16'd13927, 16'd63305, 16'd21513, 16'd41181, 16'd16059, 16'd4896, 16'd34816, 16'd17633, 16'd18149, 16'd24240, 16'd47092, 16'd22029, 16'd56510, 16'd49948, 16'd51356, 16'd39882, 16'd20299, 16'd10554, 16'd63758, 16'd34486, 16'd21401, 16'd41531, 16'd28981, 16'd41246});
	test_expansion(128'h6cdc915b7f60912c666dd057c8ce5a84, {16'd63218, 16'd45394, 16'd54410, 16'd14347, 16'd14363, 16'd22480, 16'd57395, 16'd48345, 16'd15636, 16'd7691, 16'd23424, 16'd16337, 16'd46487, 16'd47090, 16'd45393, 16'd44591, 16'd29180, 16'd17453, 16'd35, 16'd54139, 16'd11818, 16'd47002, 16'd41795, 16'd3324, 16'd54142, 16'd28064});
	test_expansion(128'ha65f45a0946c2cef828bcbd11f5f0b23, {16'd65333, 16'd28345, 16'd33875, 16'd65365, 16'd47962, 16'd22624, 16'd62402, 16'd21130, 16'd19793, 16'd16709, 16'd11551, 16'd16445, 16'd50651, 16'd59520, 16'd36392, 16'd44432, 16'd19771, 16'd18643, 16'd2635, 16'd23904, 16'd11635, 16'd32530, 16'd19467, 16'd42197, 16'd41425, 16'd37714});
	test_expansion(128'h2d94299620b9443281bc0560b44a3892, {16'd33736, 16'd27008, 16'd21112, 16'd49623, 16'd8144, 16'd4481, 16'd2381, 16'd61723, 16'd13482, 16'd12806, 16'd8094, 16'd55399, 16'd57267, 16'd60222, 16'd52561, 16'd41935, 16'd25772, 16'd21126, 16'd41280, 16'd48949, 16'd19742, 16'd31846, 16'd25274, 16'd65198, 16'd26584, 16'd7345});
	test_expansion(128'h5a33b1b60eaec0cec2d7f13fab344b3e, {16'd51035, 16'd17440, 16'd6962, 16'd40763, 16'd26430, 16'd16423, 16'd20324, 16'd50947, 16'd20269, 16'd17075, 16'd55319, 16'd61820, 16'd36133, 16'd25889, 16'd27895, 16'd20342, 16'd18416, 16'd2608, 16'd22429, 16'd44721, 16'd39387, 16'd7510, 16'd15279, 16'd7200, 16'd6151, 16'd15018});
	test_expansion(128'h1588b4fbc83100cf187dbc06ede45660, {16'd44641, 16'd55349, 16'd39756, 16'd10800, 16'd41055, 16'd29412, 16'd39129, 16'd37235, 16'd26072, 16'd32941, 16'd13968, 16'd8759, 16'd42357, 16'd34455, 16'd45120, 16'd48926, 16'd9556, 16'd32885, 16'd15123, 16'd53788, 16'd57956, 16'd63572, 16'd26934, 16'd23869, 16'd30003, 16'd33550});
	test_expansion(128'hac8dc77d15b5c3f1e6cc7a16932d049b, {16'd64839, 16'd44559, 16'd61633, 16'd12612, 16'd45963, 16'd7954, 16'd14543, 16'd41033, 16'd51936, 16'd9494, 16'd19905, 16'd25085, 16'd26081, 16'd18960, 16'd34982, 16'd40042, 16'd40946, 16'd27248, 16'd57234, 16'd21351, 16'd10560, 16'd30128, 16'd49961, 16'd21083, 16'd37534, 16'd174});
	test_expansion(128'hc4c8a349fbbac7b95d35cf6d0bda837d, {16'd10813, 16'd14483, 16'd31617, 16'd40257, 16'd6622, 16'd16043, 16'd56426, 16'd63725, 16'd1870, 16'd21687, 16'd55494, 16'd16448, 16'd48551, 16'd1538, 16'd38304, 16'd13130, 16'd16720, 16'd41544, 16'd2596, 16'd30351, 16'd17799, 16'd17705, 16'd52396, 16'd53200, 16'd40215, 16'd63764});
	test_expansion(128'hb39f5b8d30bb679994462cff1c70c2d2, {16'd12799, 16'd3486, 16'd8443, 16'd10505, 16'd45794, 16'd55755, 16'd36566, 16'd26144, 16'd10272, 16'd44643, 16'd27739, 16'd28446, 16'd19828, 16'd31004, 16'd19031, 16'd7569, 16'd29983, 16'd14349, 16'd38733, 16'd22278, 16'd3418, 16'd35602, 16'd7578, 16'd54922, 16'd44775, 16'd50134});
	test_expansion(128'h840ed831c328c848d97c274d48c04188, {16'd41231, 16'd13540, 16'd54226, 16'd43034, 16'd24574, 16'd4404, 16'd27643, 16'd56583, 16'd29780, 16'd31442, 16'd19080, 16'd13342, 16'd22462, 16'd3145, 16'd16936, 16'd25126, 16'd8570, 16'd14132, 16'd49337, 16'd40416, 16'd169, 16'd33209, 16'd7741, 16'd12833, 16'd10078, 16'd43904});
	test_expansion(128'h9d6b01c630c7820cf22c181c9e593f32, {16'd9244, 16'd46682, 16'd22142, 16'd23461, 16'd52940, 16'd30521, 16'd8291, 16'd51161, 16'd63540, 16'd2210, 16'd43282, 16'd3153, 16'd62024, 16'd62556, 16'd49519, 16'd12601, 16'd48899, 16'd56969, 16'd38639, 16'd53525, 16'd53616, 16'd24046, 16'd54742, 16'd42167, 16'd60867, 16'd9595});
	test_expansion(128'h6e7dc2c2eaa417abf69c28768cf2360f, {16'd60261, 16'd13698, 16'd40148, 16'd9648, 16'd15914, 16'd7229, 16'd27429, 16'd17236, 16'd29935, 16'd45707, 16'd55889, 16'd42317, 16'd44512, 16'd49822, 16'd39973, 16'd12046, 16'd61206, 16'd10056, 16'd35958, 16'd18129, 16'd18072, 16'd59584, 16'd37467, 16'd26968, 16'd47259, 16'd37070});
	test_expansion(128'he0aa86d9ff416f442657666d11a57be0, {16'd19637, 16'd47669, 16'd40173, 16'd8224, 16'd33742, 16'd23605, 16'd35011, 16'd3799, 16'd9902, 16'd62443, 16'd54490, 16'd29664, 16'd37379, 16'd11248, 16'd65435, 16'd47522, 16'd57723, 16'd41269, 16'd4348, 16'd39666, 16'd7721, 16'd31437, 16'd19110, 16'd56829, 16'd25894, 16'd56277});
	test_expansion(128'h071684a6ad41069f1e675c307542b9a1, {16'd39221, 16'd11863, 16'd56608, 16'd50030, 16'd40691, 16'd33712, 16'd41254, 16'd46654, 16'd55180, 16'd2952, 16'd26090, 16'd33445, 16'd18034, 16'd11033, 16'd20638, 16'd43007, 16'd61467, 16'd59747, 16'd15463, 16'd9373, 16'd5619, 16'd27205, 16'd1242, 16'd64002, 16'd5566, 16'd17128});
	test_expansion(128'h678ec97f196d5112d13a87225bcad030, {16'd51097, 16'd11044, 16'd6294, 16'd63634, 16'd24355, 16'd46267, 16'd61784, 16'd31147, 16'd34878, 16'd41928, 16'd29669, 16'd16077, 16'd21260, 16'd13137, 16'd46446, 16'd49802, 16'd14743, 16'd16212, 16'd10518, 16'd65402, 16'd52354, 16'd40130, 16'd29318, 16'd6253, 16'd1322, 16'd556});
	test_expansion(128'h136bb86196ae6424f4fcb549b50fbe0e, {16'd49076, 16'd4305, 16'd60319, 16'd60247, 16'd63286, 16'd36606, 16'd31695, 16'd57815, 16'd5574, 16'd58615, 16'd28536, 16'd12894, 16'd47040, 16'd26171, 16'd28162, 16'd29149, 16'd34036, 16'd41586, 16'd7536, 16'd45610, 16'd6956, 16'd58269, 16'd63495, 16'd22088, 16'd62929, 16'd9163});
	test_expansion(128'h02d355bb0c5ebc53d69fc537f8bbb829, {16'd38017, 16'd43274, 16'd14532, 16'd14096, 16'd19943, 16'd10340, 16'd19369, 16'd55240, 16'd48758, 16'd63401, 16'd15310, 16'd30230, 16'd51484, 16'd8072, 16'd46534, 16'd22199, 16'd29415, 16'd21690, 16'd16156, 16'd34443, 16'd25715, 16'd47894, 16'd62658, 16'd63313, 16'd65034, 16'd44697});
	test_expansion(128'h6cba516a1796a664e4400cb55dd95302, {16'd63451, 16'd42613, 16'd12690, 16'd45792, 16'd45177, 16'd43217, 16'd48871, 16'd33945, 16'd43137, 16'd651, 16'd33714, 16'd15807, 16'd30758, 16'd20190, 16'd8675, 16'd23959, 16'd43969, 16'd36149, 16'd59577, 16'd33813, 16'd55938, 16'd35934, 16'd38436, 16'd31929, 16'd60476, 16'd14779});
	test_expansion(128'hbaf51614e32a842156ec8fd63e679fc9, {16'd16709, 16'd44835, 16'd62604, 16'd37264, 16'd52853, 16'd4579, 16'd43105, 16'd62051, 16'd11277, 16'd61438, 16'd23242, 16'd24234, 16'd21747, 16'd55258, 16'd28623, 16'd21618, 16'd65229, 16'd30747, 16'd1081, 16'd52546, 16'd53260, 16'd29884, 16'd26979, 16'd20424, 16'd55882, 16'd57948});
	test_expansion(128'h41886fd4ab6f38998ea24e8556a21b3e, {16'd49590, 16'd50561, 16'd3998, 16'd63176, 16'd13524, 16'd39030, 16'd4333, 16'd14930, 16'd23960, 16'd55001, 16'd31853, 16'd42572, 16'd30095, 16'd30965, 16'd20034, 16'd10051, 16'd62064, 16'd36115, 16'd14310, 16'd13983, 16'd26623, 16'd48879, 16'd11749, 16'd47393, 16'd25839, 16'd50320});
	test_expansion(128'hde60d86f44fdf87e5a6bf08f80162dc1, {16'd30952, 16'd56909, 16'd44765, 16'd28284, 16'd6989, 16'd9488, 16'd14126, 16'd11863, 16'd21152, 16'd17184, 16'd35621, 16'd1703, 16'd22647, 16'd44391, 16'd33676, 16'd10068, 16'd29959, 16'd11021, 16'd47725, 16'd25820, 16'd18942, 16'd25771, 16'd47822, 16'd34073, 16'd18960, 16'd48843});
	test_expansion(128'hf268e003efacf81656d96439f3054cff, {16'd33838, 16'd50806, 16'd49891, 16'd60979, 16'd28898, 16'd14439, 16'd47164, 16'd46100, 16'd47019, 16'd22914, 16'd15186, 16'd16417, 16'd44696, 16'd54088, 16'd29091, 16'd56112, 16'd12069, 16'd62260, 16'd52866, 16'd25054, 16'd21010, 16'd25377, 16'd52087, 16'd41074, 16'd4075, 16'd64464});
	test_expansion(128'hee9fd52b2549c0a7046509b60a7da224, {16'd49877, 16'd23263, 16'd46055, 16'd57256, 16'd65174, 16'd9700, 16'd54822, 16'd23654, 16'd19079, 16'd45160, 16'd3334, 16'd38800, 16'd64540, 16'd53724, 16'd61116, 16'd60088, 16'd26500, 16'd2280, 16'd37427, 16'd12466, 16'd1163, 16'd4677, 16'd28722, 16'd64033, 16'd20332, 16'd2193});
	test_expansion(128'h2a2b6703ddb231bbcb8bd7fb705d5cc2, {16'd23032, 16'd37673, 16'd44780, 16'd7528, 16'd59308, 16'd24300, 16'd54034, 16'd37565, 16'd59999, 16'd28979, 16'd39428, 16'd52934, 16'd64358, 16'd33924, 16'd12975, 16'd27126, 16'd18546, 16'd57628, 16'd22677, 16'd9857, 16'd4972, 16'd58967, 16'd37985, 16'd12015, 16'd19719, 16'd13391});
	test_expansion(128'h8a50caa3fbf679851d4a2bb6f028ddaa, {16'd57341, 16'd15251, 16'd36355, 16'd38042, 16'd57165, 16'd38968, 16'd14842, 16'd7748, 16'd27262, 16'd43882, 16'd14676, 16'd59368, 16'd4935, 16'd5161, 16'd63828, 16'd28269, 16'd52246, 16'd65426, 16'd29287, 16'd64133, 16'd33205, 16'd33175, 16'd45171, 16'd10265, 16'd36094, 16'd29350});
	test_expansion(128'h2237e4378f33ee7ebe410cbdc57a9994, {16'd14058, 16'd22754, 16'd40818, 16'd21033, 16'd33034, 16'd27535, 16'd61097, 16'd1776, 16'd41860, 16'd54616, 16'd20427, 16'd24991, 16'd55299, 16'd59951, 16'd4733, 16'd15664, 16'd260, 16'd51409, 16'd4122, 16'd25098, 16'd62198, 16'd45692, 16'd8231, 16'd47577, 16'd62105, 16'd23876});
	test_expansion(128'h73c41724477c9e3cf565d637955f0e7f, {16'd26949, 16'd5152, 16'd26219, 16'd55831, 16'd61568, 16'd51046, 16'd51794, 16'd17120, 16'd49635, 16'd42582, 16'd29208, 16'd50609, 16'd52665, 16'd10914, 16'd41506, 16'd56896, 16'd45786, 16'd36154, 16'd61495, 16'd40944, 16'd9510, 16'd22618, 16'd9128, 16'd41437, 16'd65054, 16'd60345});
	test_expansion(128'h9e04b779a949bc43dee878c8ed7c1ddc, {16'd34689, 16'd56706, 16'd1593, 16'd7755, 16'd22836, 16'd7771, 16'd35556, 16'd42414, 16'd40234, 16'd12332, 16'd28898, 16'd48181, 16'd20621, 16'd45632, 16'd6819, 16'd31054, 16'd62466, 16'd64582, 16'd6081, 16'd45239, 16'd3308, 16'd42812, 16'd20126, 16'd44952, 16'd39793, 16'd52716});
	test_expansion(128'he78472b4108e0db400c3ffbca16a00d9, {16'd13637, 16'd15318, 16'd2403, 16'd1879, 16'd15296, 16'd14036, 16'd23160, 16'd49622, 16'd61248, 16'd41275, 16'd38378, 16'd9008, 16'd36212, 16'd18011, 16'd50155, 16'd5031, 16'd58260, 16'd11047, 16'd19263, 16'd57158, 16'd21263, 16'd4110, 16'd28346, 16'd3704, 16'd41444, 16'd33607});
	test_expansion(128'hb08e0cf79c02aebdcbfa8c3a5d048d5e, {16'd62690, 16'd22705, 16'd29315, 16'd50520, 16'd44517, 16'd48770, 16'd954, 16'd37014, 16'd33590, 16'd21458, 16'd44555, 16'd44487, 16'd12684, 16'd51959, 16'd12903, 16'd26075, 16'd16016, 16'd47806, 16'd64706, 16'd29528, 16'd23422, 16'd32088, 16'd21395, 16'd55599, 16'd56945, 16'd41812});
	test_expansion(128'hf08b76fd57ea7e97d6c6aa47f4907bb9, {16'd20275, 16'd63845, 16'd12513, 16'd21057, 16'd28183, 16'd57514, 16'd17178, 16'd6293, 16'd730, 16'd29570, 16'd60349, 16'd38630, 16'd35520, 16'd15801, 16'd25060, 16'd41846, 16'd4676, 16'd39524, 16'd60143, 16'd16811, 16'd43976, 16'd60902, 16'd42225, 16'd33769, 16'd7121, 16'd5980});
	test_expansion(128'hd3f96f5dd803c72502606a7ec163eb47, {16'd32926, 16'd61856, 16'd54932, 16'd3511, 16'd54048, 16'd24381, 16'd53695, 16'd19882, 16'd4970, 16'd3016, 16'd23160, 16'd60959, 16'd54613, 16'd54133, 16'd14594, 16'd5111, 16'd52051, 16'd13462, 16'd51786, 16'd57195, 16'd53924, 16'd374, 16'd29133, 16'd63610, 16'd50406, 16'd25628});
	test_expansion(128'h8964300e98ba2e2a18e952b68a16cfc5, {16'd17376, 16'd64857, 16'd55614, 16'd16831, 16'd38136, 16'd37505, 16'd58048, 16'd37457, 16'd57998, 16'd24628, 16'd46978, 16'd53799, 16'd22020, 16'd22824, 16'd27214, 16'd25517, 16'd17485, 16'd38000, 16'd14521, 16'd18170, 16'd29258, 16'd62343, 16'd43198, 16'd27278, 16'd58973, 16'd28799});
	test_expansion(128'h8f3fe25cb5490d31fafdfe14a6bc2d60, {16'd48070, 16'd59025, 16'd44566, 16'd10340, 16'd3278, 16'd59511, 16'd5480, 16'd60700, 16'd13179, 16'd29088, 16'd21621, 16'd161, 16'd23445, 16'd7628, 16'd51808, 16'd8892, 16'd35374, 16'd29841, 16'd1696, 16'd60582, 16'd31628, 16'd29467, 16'd61569, 16'd51674, 16'd23842, 16'd18482});
	test_expansion(128'hd8ef7645422974b25742e70bf12092c2, {16'd33040, 16'd40185, 16'd22261, 16'd32549, 16'd176, 16'd11451, 16'd56086, 16'd58380, 16'd2101, 16'd1426, 16'd45880, 16'd34526, 16'd4308, 16'd29181, 16'd55180, 16'd48932, 16'd35015, 16'd18988, 16'd32631, 16'd664, 16'd34484, 16'd29916, 16'd42068, 16'd48188, 16'd36497, 16'd40394});
	test_expansion(128'hb8c38dc24fcd5fe685094213fdb15f93, {16'd5748, 16'd49570, 16'd64287, 16'd39795, 16'd60173, 16'd30775, 16'd53032, 16'd8989, 16'd6964, 16'd56170, 16'd52104, 16'd18315, 16'd64090, 16'd55456, 16'd42593, 16'd31472, 16'd13856, 16'd22337, 16'd64983, 16'd18301, 16'd56008, 16'd6119, 16'd5932, 16'd48900, 16'd16676, 16'd31536});
	test_expansion(128'h604d7252cfee0619a6917070eceb6f3e, {16'd49934, 16'd24472, 16'd31198, 16'd32662, 16'd35378, 16'd38893, 16'd10097, 16'd29817, 16'd32774, 16'd14215, 16'd47629, 16'd19582, 16'd2909, 16'd19848, 16'd64286, 16'd23614, 16'd59194, 16'd23841, 16'd5925, 16'd1185, 16'd28100, 16'd30781, 16'd5710, 16'd16051, 16'd33388, 16'd17971});
	test_expansion(128'h7b246190ba3126ef5f9f191ddba927e3, {16'd36626, 16'd50015, 16'd438, 16'd23586, 16'd15374, 16'd7875, 16'd23049, 16'd56938, 16'd59299, 16'd42473, 16'd6647, 16'd18037, 16'd18733, 16'd270, 16'd3816, 16'd55326, 16'd38973, 16'd8123, 16'd40033, 16'd51639, 16'd5960, 16'd62753, 16'd27673, 16'd5477, 16'd5140, 16'd10891});
	test_expansion(128'h8b5f5d20417a863596d7cf5ed7ebf97c, {16'd41481, 16'd62814, 16'd47911, 16'd15514, 16'd63499, 16'd63477, 16'd24567, 16'd31811, 16'd49910, 16'd7523, 16'd37447, 16'd45978, 16'd58005, 16'd64377, 16'd31042, 16'd19706, 16'd40396, 16'd36014, 16'd42441, 16'd55916, 16'd58525, 16'd44677, 16'd48785, 16'd23277, 16'd47200, 16'd29726});
	test_expansion(128'haf145054235796573c382ab05f1bf066, {16'd43785, 16'd19804, 16'd29525, 16'd10797, 16'd54292, 16'd20988, 16'd29701, 16'd3656, 16'd30059, 16'd11733, 16'd63406, 16'd64336, 16'd30002, 16'd10137, 16'd48343, 16'd15056, 16'd12680, 16'd47726, 16'd52693, 16'd6577, 16'd36685, 16'd42719, 16'd19647, 16'd46526, 16'd30847, 16'd30622});
	test_expansion(128'hbd433a10573d64c5af1afccda242f4ef, {16'd59501, 16'd25024, 16'd39640, 16'd42522, 16'd46220, 16'd42555, 16'd65467, 16'd40283, 16'd27594, 16'd17097, 16'd49518, 16'd37965, 16'd13978, 16'd61782, 16'd21765, 16'd49426, 16'd34164, 16'd48089, 16'd8841, 16'd8246, 16'd37445, 16'd22439, 16'd36, 16'd29448, 16'd50916, 16'd42703});
	test_expansion(128'hf689c5649d32bc1177d877fb4f2aa208, {16'd19793, 16'd42640, 16'd60589, 16'd28975, 16'd51788, 16'd44082, 16'd58669, 16'd18333, 16'd25581, 16'd5791, 16'd7849, 16'd47943, 16'd18079, 16'd1941, 16'd51688, 16'd39275, 16'd8119, 16'd2887, 16'd47686, 16'd22675, 16'd716, 16'd12984, 16'd44496, 16'd23080, 16'd46712, 16'd50849});
	test_expansion(128'h010b6fa0be167e9cd12f14f5075b4dd3, {16'd14264, 16'd16254, 16'd12707, 16'd32364, 16'd51012, 16'd36011, 16'd53629, 16'd38176, 16'd57214, 16'd5421, 16'd47116, 16'd29068, 16'd59090, 16'd58081, 16'd26663, 16'd13344, 16'd23143, 16'd39807, 16'd46361, 16'd35236, 16'd33221, 16'd15174, 16'd13157, 16'd23162, 16'd30117, 16'd43448});
	test_expansion(128'h9781dffea9c5aeaf980c7500722e3490, {16'd5798, 16'd21845, 16'd51657, 16'd11391, 16'd912, 16'd50344, 16'd35987, 16'd57635, 16'd25362, 16'd3345, 16'd29544, 16'd11585, 16'd41522, 16'd63704, 16'd42439, 16'd38797, 16'd32336, 16'd63061, 16'd43335, 16'd3226, 16'd40040, 16'd23665, 16'd1230, 16'd15921, 16'd35813, 16'd27729});
	test_expansion(128'h6c9f664586521d7cf87500fccb8be7af, {16'd65484, 16'd2436, 16'd31466, 16'd17294, 16'd54979, 16'd710, 16'd41088, 16'd41434, 16'd27429, 16'd2078, 16'd9530, 16'd13455, 16'd57367, 16'd11085, 16'd31387, 16'd14497, 16'd46629, 16'd19617, 16'd11328, 16'd47061, 16'd9003, 16'd42307, 16'd48424, 16'd33012, 16'd57523, 16'd48440});
	test_expansion(128'hcc6cf2b0ccfbfa21568e6ef6c648b50d, {16'd56887, 16'd19726, 16'd8591, 16'd37099, 16'd56440, 16'd3055, 16'd21453, 16'd56845, 16'd34384, 16'd27216, 16'd22778, 16'd1424, 16'd28962, 16'd20983, 16'd40525, 16'd64714, 16'd57590, 16'd403, 16'd26665, 16'd11043, 16'd8016, 16'd29041, 16'd59254, 16'd36182, 16'd18245, 16'd8913});
	test_expansion(128'h2460484cdffe34f57e23881698129bf8, {16'd35643, 16'd3770, 16'd21061, 16'd41856, 16'd4408, 16'd635, 16'd11236, 16'd39479, 16'd21249, 16'd47731, 16'd32684, 16'd42799, 16'd10328, 16'd43073, 16'd23004, 16'd64134, 16'd15171, 16'd50009, 16'd29236, 16'd13090, 16'd22227, 16'd9541, 16'd40703, 16'd16884, 16'd63539, 16'd50584});
	test_expansion(128'h735f0f07399a34332501aa4c6dd76d8f, {16'd6431, 16'd19535, 16'd7432, 16'd30655, 16'd20173, 16'd20371, 16'd34414, 16'd13851, 16'd8120, 16'd51737, 16'd6253, 16'd43371, 16'd1769, 16'd46955, 16'd36127, 16'd25481, 16'd64005, 16'd56684, 16'd11939, 16'd10989, 16'd25456, 16'd47092, 16'd34212, 16'd2735, 16'd39744, 16'd55662});
	test_expansion(128'hc8df3f24d345ebd0c8f55a13e82e270c, {16'd30098, 16'd22237, 16'd10897, 16'd42308, 16'd27198, 16'd28275, 16'd63517, 16'd30349, 16'd8148, 16'd7433, 16'd58077, 16'd57786, 16'd7167, 16'd19533, 16'd33988, 16'd58925, 16'd60055, 16'd41930, 16'd56714, 16'd61994, 16'd7072, 16'd51887, 16'd13920, 16'd42139, 16'd61000, 16'd31954});
	test_expansion(128'h91ab238cc5a8c5e46893b1ccc02560e6, {16'd50036, 16'd40886, 16'd30477, 16'd27558, 16'd24602, 16'd3138, 16'd12012, 16'd24710, 16'd5941, 16'd63028, 16'd57174, 16'd4284, 16'd36263, 16'd16439, 16'd37190, 16'd62777, 16'd49045, 16'd30183, 16'd57411, 16'd51777, 16'd8824, 16'd24383, 16'd716, 16'd50255, 16'd58274, 16'd36768});
	test_expansion(128'hd9bad66bcd2bf338f75acf54115c3c99, {16'd43322, 16'd51317, 16'd13884, 16'd53892, 16'd50645, 16'd36356, 16'd11081, 16'd60770, 16'd33681, 16'd23747, 16'd29395, 16'd14374, 16'd34216, 16'd8404, 16'd47684, 16'd4465, 16'd6025, 16'd47760, 16'd19528, 16'd9727, 16'd13450, 16'd49199, 16'd49450, 16'd50235, 16'd52486, 16'd38696});
	test_expansion(128'h4a964925be661f7f9722fb87a4645e5a, {16'd20384, 16'd25618, 16'd55182, 16'd16867, 16'd40686, 16'd7054, 16'd46914, 16'd2933, 16'd51259, 16'd33575, 16'd35533, 16'd2164, 16'd13033, 16'd46613, 16'd29247, 16'd52404, 16'd20418, 16'd64228, 16'd17534, 16'd50401, 16'd39781, 16'd50045, 16'd48755, 16'd51075, 16'd22266, 16'd26289});
	test_expansion(128'h7036903fff4289099cbbb03dc4f1e62a, {16'd17915, 16'd50879, 16'd33428, 16'd13444, 16'd54224, 16'd34374, 16'd10107, 16'd26388, 16'd42624, 16'd22291, 16'd46035, 16'd60583, 16'd15240, 16'd43312, 16'd32595, 16'd38248, 16'd25373, 16'd57600, 16'd18698, 16'd41040, 16'd20966, 16'd63119, 16'd34629, 16'd42575, 16'd61762, 16'd8773});
	test_expansion(128'h5cddeeebcc91ed564d3cbc72951cbb3f, {16'd25905, 16'd1026, 16'd54664, 16'd37833, 16'd53524, 16'd21771, 16'd51414, 16'd15716, 16'd60332, 16'd43031, 16'd2368, 16'd43612, 16'd1805, 16'd31988, 16'd841, 16'd39687, 16'd45778, 16'd52094, 16'd24008, 16'd16866, 16'd55868, 16'd25120, 16'd63031, 16'd16880, 16'd23866, 16'd7607});
	test_expansion(128'h3cc2d4a10d4e420c04c82cd1eabc8060, {16'd23686, 16'd24464, 16'd13402, 16'd17078, 16'd30955, 16'd18759, 16'd47631, 16'd14528, 16'd22181, 16'd4982, 16'd34134, 16'd33440, 16'd19567, 16'd38179, 16'd16212, 16'd18104, 16'd22635, 16'd22290, 16'd48592, 16'd8861, 16'd17667, 16'd60861, 16'd8149, 16'd62624, 16'd9, 16'd19891});
	test_expansion(128'h19b86177f1201b3b41e7e5fdfe484c98, {16'd51466, 16'd33055, 16'd56294, 16'd17670, 16'd14063, 16'd9822, 16'd58397, 16'd19784, 16'd33467, 16'd60015, 16'd18908, 16'd37417, 16'd65004, 16'd12972, 16'd14905, 16'd62412, 16'd38499, 16'd25251, 16'd20044, 16'd63989, 16'd55729, 16'd50754, 16'd55010, 16'd39817, 16'd61674, 16'd26982});
	test_expansion(128'h21c9fb95361ce308c4084342761f1c56, {16'd3717, 16'd32556, 16'd2338, 16'd31443, 16'd3650, 16'd16548, 16'd29169, 16'd55707, 16'd10841, 16'd46827, 16'd566, 16'd36471, 16'd17797, 16'd65495, 16'd7573, 16'd14057, 16'd47450, 16'd28027, 16'd39013, 16'd39602, 16'd30160, 16'd54811, 16'd64180, 16'd35201, 16'd909, 16'd63659});
	test_expansion(128'hed39c0d5cfc6fb1c8ff232b3b0bdd81d, {16'd17939, 16'd3, 16'd46700, 16'd33490, 16'd11962, 16'd38540, 16'd32886, 16'd37201, 16'd47692, 16'd44233, 16'd45815, 16'd41250, 16'd18652, 16'd21040, 16'd55672, 16'd23745, 16'd52421, 16'd49568, 16'd29141, 16'd14515, 16'd14288, 16'd27459, 16'd48249, 16'd10717, 16'd17854, 16'd55371});
	test_expansion(128'h464f3e00c0f4cce8107d73ee45750173, {16'd34831, 16'd60268, 16'd30385, 16'd50452, 16'd14273, 16'd35292, 16'd26984, 16'd47611, 16'd9393, 16'd11673, 16'd47524, 16'd63132, 16'd57431, 16'd24611, 16'd60517, 16'd10497, 16'd45723, 16'd28841, 16'd16856, 16'd31017, 16'd5827, 16'd31997, 16'd3, 16'd44157, 16'd39628, 16'd26016});
	test_expansion(128'hb56b94e288bd9ebe6deff0cbe4c34fcf, {16'd5862, 16'd21735, 16'd20834, 16'd7130, 16'd22370, 16'd62632, 16'd48929, 16'd32677, 16'd4765, 16'd31405, 16'd49651, 16'd36957, 16'd14616, 16'd15985, 16'd57801, 16'd47656, 16'd53488, 16'd47787, 16'd62083, 16'd13551, 16'd33933, 16'd47532, 16'd20218, 16'd16804, 16'd11215, 16'd30146});
	test_expansion(128'heaa2a2a2eb18740d7fb7603b89b176f9, {16'd1707, 16'd33320, 16'd9195, 16'd60695, 16'd55941, 16'd18618, 16'd60918, 16'd35615, 16'd7446, 16'd7, 16'd53084, 16'd12070, 16'd63311, 16'd9415, 16'd21589, 16'd10906, 16'd2722, 16'd39441, 16'd2538, 16'd11385, 16'd31566, 16'd1401, 16'd42812, 16'd40475, 16'd57903, 16'd37843});
	test_expansion(128'ha85574abaab7a9a558618b840ffc5807, {16'd177, 16'd33747, 16'd40139, 16'd24452, 16'd10579, 16'd51127, 16'd53388, 16'd53629, 16'd58162, 16'd61488, 16'd27669, 16'd52560, 16'd14879, 16'd25975, 16'd49835, 16'd64523, 16'd41773, 16'd58152, 16'd43541, 16'd37240, 16'd53274, 16'd24838, 16'd35509, 16'd56407, 16'd62525, 16'd7082});
	test_expansion(128'h1edd06e17024f5aaf53404518451d3a2, {16'd34916, 16'd7555, 16'd51424, 16'd65070, 16'd50241, 16'd57853, 16'd30297, 16'd24114, 16'd16785, 16'd6946, 16'd2218, 16'd40764, 16'd40703, 16'd29656, 16'd64321, 16'd29830, 16'd59851, 16'd26664, 16'd17583, 16'd53378, 16'd31664, 16'd36786, 16'd23602, 16'd50018, 16'd53766, 16'd28536});
	test_expansion(128'h943cfb5e11bf58637229d9f334a35b4c, {16'd42802, 16'd30511, 16'd41797, 16'd6524, 16'd8949, 16'd57854, 16'd58548, 16'd53380, 16'd14197, 16'd40922, 16'd3055, 16'd20492, 16'd24478, 16'd19525, 16'd38528, 16'd51166, 16'd55742, 16'd37299, 16'd28180, 16'd29372, 16'd62190, 16'd24901, 16'd64316, 16'd28615, 16'd26825, 16'd40420});
	test_expansion(128'h27d3579a949a764909070200ac67ae33, {16'd7693, 16'd60459, 16'd11184, 16'd59612, 16'd45982, 16'd56557, 16'd11352, 16'd1693, 16'd27108, 16'd33725, 16'd7176, 16'd42269, 16'd1634, 16'd39268, 16'd44213, 16'd30613, 16'd56747, 16'd47144, 16'd2392, 16'd2697, 16'd27104, 16'd62128, 16'd55729, 16'd30480, 16'd28114, 16'd17604});
	test_expansion(128'h3eee02166a5bb6da3d09a37427ebd79d, {16'd39320, 16'd13093, 16'd47527, 16'd6660, 16'd54487, 16'd20524, 16'd54606, 16'd55576, 16'd8338, 16'd16940, 16'd52672, 16'd30044, 16'd55565, 16'd22631, 16'd47902, 16'd11675, 16'd23972, 16'd6082, 16'd45566, 16'd52060, 16'd29753, 16'd3654, 16'd647, 16'd58520, 16'd60584, 16'd9107});
	test_expansion(128'h9b83e4b52d024d955368904d8dd5b5fa, {16'd43205, 16'd34555, 16'd36944, 16'd3002, 16'd18303, 16'd8707, 16'd18234, 16'd39095, 16'd35440, 16'd21861, 16'd39202, 16'd34766, 16'd33002, 16'd1196, 16'd50537, 16'd36088, 16'd11443, 16'd10605, 16'd46473, 16'd60977, 16'd33679, 16'd58547, 16'd38649, 16'd29602, 16'd51850, 16'd29436});
	test_expansion(128'he0edea2035a96095151578081f04e6de, {16'd8926, 16'd44664, 16'd27605, 16'd52962, 16'd16034, 16'd620, 16'd33042, 16'd14563, 16'd44933, 16'd41404, 16'd49376, 16'd29320, 16'd5735, 16'd28345, 16'd64062, 16'd31115, 16'd19844, 16'd13456, 16'd37662, 16'd62009, 16'd15986, 16'd5650, 16'd22283, 16'd40224, 16'd10373, 16'd13305});
	test_expansion(128'hb98ae727a483fea8cc6d81d8f65c3d18, {16'd645, 16'd61007, 16'd36429, 16'd14286, 16'd65249, 16'd39549, 16'd58102, 16'd17430, 16'd47880, 16'd32548, 16'd14000, 16'd21976, 16'd41103, 16'd26998, 16'd32528, 16'd34077, 16'd14061, 16'd37096, 16'd10709, 16'd29543, 16'd49820, 16'd27624, 16'd12909, 16'd27589, 16'd59559, 16'd55123});
	test_expansion(128'h4f9101039cd5b9bf923659b491954208, {16'd51939, 16'd51801, 16'd42581, 16'd41881, 16'd17396, 16'd22674, 16'd42366, 16'd36477, 16'd23480, 16'd65510, 16'd14192, 16'd52599, 16'd44350, 16'd40135, 16'd63414, 16'd38469, 16'd1711, 16'd49147, 16'd51692, 16'd20759, 16'd23120, 16'd19575, 16'd55478, 16'd8011, 16'd30423, 16'd22128});
	test_expansion(128'hb341e6cb88de61708a5f371ba8afe51c, {16'd53010, 16'd65448, 16'd44169, 16'd9783, 16'd48317, 16'd59371, 16'd27869, 16'd43795, 16'd51017, 16'd36341, 16'd46517, 16'd56359, 16'd25933, 16'd682, 16'd16187, 16'd41438, 16'd17314, 16'd41058, 16'd60611, 16'd295, 16'd10049, 16'd6059, 16'd30969, 16'd4911, 16'd7187, 16'd47782});
	test_expansion(128'h8134313984cb60196f8d9b60fc779e82, {16'd11996, 16'd44737, 16'd42385, 16'd20857, 16'd54045, 16'd29978, 16'd64031, 16'd24106, 16'd27586, 16'd20707, 16'd63784, 16'd38212, 16'd63228, 16'd59648, 16'd24915, 16'd21573, 16'd28764, 16'd32215, 16'd9332, 16'd63294, 16'd39076, 16'd35060, 16'd32062, 16'd47695, 16'd7114, 16'd37757});
	test_expansion(128'hccfbb6fa22411b0d28a9b903e826136b, {16'd64215, 16'd46121, 16'd30628, 16'd60097, 16'd58849, 16'd39963, 16'd65281, 16'd10286, 16'd47099, 16'd56912, 16'd28735, 16'd51834, 16'd26088, 16'd26179, 16'd3658, 16'd9972, 16'd14507, 16'd25646, 16'd21685, 16'd43376, 16'd33199, 16'd59877, 16'd1987, 16'd41031, 16'd34486, 16'd23311});
	test_expansion(128'hb762f10dd15b39253e4db8af31772d09, {16'd35593, 16'd6462, 16'd47458, 16'd4633, 16'd56259, 16'd43707, 16'd7024, 16'd49706, 16'd4171, 16'd14559, 16'd4485, 16'd60174, 16'd20818, 16'd12613, 16'd13797, 16'd31843, 16'd58134, 16'd47692, 16'd28961, 16'd14975, 16'd43141, 16'd7078, 16'd53750, 16'd28835, 16'd3331, 16'd13067});
	test_expansion(128'hbfdd10104a96cd68cbe92ce360517627, {16'd21288, 16'd52848, 16'd36320, 16'd52123, 16'd78, 16'd10109, 16'd19444, 16'd19425, 16'd8396, 16'd45444, 16'd11618, 16'd63430, 16'd23645, 16'd63034, 16'd159, 16'd41966, 16'd24568, 16'd46815, 16'd21592, 16'd57803, 16'd50939, 16'd21797, 16'd21329, 16'd52590, 16'd55557, 16'd63757});
	test_expansion(128'h069a591ea6ea1ffcb42d2906bf4900d2, {16'd32385, 16'd45727, 16'd5159, 16'd48462, 16'd31957, 16'd32999, 16'd48333, 16'd900, 16'd65070, 16'd64814, 16'd14036, 16'd7040, 16'd4463, 16'd24595, 16'd9668, 16'd12822, 16'd22758, 16'd24295, 16'd44393, 16'd37506, 16'd23375, 16'd1420, 16'd34916, 16'd8184, 16'd29945, 16'd9146});
	test_expansion(128'h899704e18edfa72a802ee32e92a770b2, {16'd5589, 16'd48161, 16'd39773, 16'd2545, 16'd33712, 16'd5476, 16'd30288, 16'd10967, 16'd55069, 16'd17268, 16'd30636, 16'd14195, 16'd37375, 16'd6305, 16'd63847, 16'd33549, 16'd52796, 16'd492, 16'd62901, 16'd63742, 16'd34867, 16'd14588, 16'd11054, 16'd23371, 16'd46668, 16'd34179});
	test_expansion(128'hfff2daf3e4a25f8362277bf64ca8a6f1, {16'd2340, 16'd32374, 16'd54900, 16'd54199, 16'd33572, 16'd40782, 16'd1224, 16'd33563, 16'd20929, 16'd29587, 16'd40034, 16'd18172, 16'd9350, 16'd56799, 16'd25355, 16'd46518, 16'd31843, 16'd44788, 16'd34019, 16'd10150, 16'd56629, 16'd7727, 16'd13194, 16'd50142, 16'd12554, 16'd25115});
	test_expansion(128'h159472cec16666c33de7fc6160305ada, {16'd47475, 16'd8584, 16'd51054, 16'd45570, 16'd53523, 16'd60162, 16'd19461, 16'd62279, 16'd45679, 16'd13592, 16'd45818, 16'd57324, 16'd32621, 16'd6743, 16'd31725, 16'd29491, 16'd24363, 16'd17904, 16'd16406, 16'd58426, 16'd42129, 16'd3934, 16'd38475, 16'd31728, 16'd39784, 16'd40316});
	test_expansion(128'hcdda1a9b47f053a590290fee71c0b09e, {16'd56313, 16'd33406, 16'd28857, 16'd9785, 16'd23069, 16'd12812, 16'd59573, 16'd25020, 16'd53372, 16'd21298, 16'd33585, 16'd7529, 16'd22919, 16'd62626, 16'd38897, 16'd41860, 16'd36754, 16'd12435, 16'd65098, 16'd56422, 16'd4447, 16'd65461, 16'd3459, 16'd59847, 16'd3960, 16'd64537});
	test_expansion(128'h5d3377bfa83938f64581cff295c70eb3, {16'd20834, 16'd43831, 16'd21178, 16'd11778, 16'd5056, 16'd23517, 16'd21703, 16'd40844, 16'd26641, 16'd29146, 16'd24517, 16'd25689, 16'd26075, 16'd39682, 16'd38131, 16'd49670, 16'd62576, 16'd37051, 16'd9569, 16'd56102, 16'd59251, 16'd16432, 16'd64825, 16'd56802, 16'd41931, 16'd5762});
	test_expansion(128'hff775219683d00756b5449e53817896c, {16'd3399, 16'd55702, 16'd34845, 16'd11822, 16'd23179, 16'd27584, 16'd25088, 16'd33145, 16'd21421, 16'd2195, 16'd1133, 16'd1390, 16'd31318, 16'd14032, 16'd14541, 16'd49437, 16'd4283, 16'd62807, 16'd3662, 16'd33395, 16'd20023, 16'd23747, 16'd48350, 16'd649, 16'd11939, 16'd46983});
	test_expansion(128'h8404bcab8da292d01188c3ea258804fe, {16'd44900, 16'd18210, 16'd62985, 16'd48384, 16'd349, 16'd60111, 16'd15894, 16'd46354, 16'd65230, 16'd25371, 16'd22849, 16'd29006, 16'd40984, 16'd1146, 16'd59597, 16'd25038, 16'd21231, 16'd3437, 16'd2537, 16'd63839, 16'd19348, 16'd15920, 16'd24011, 16'd12394, 16'd63291, 16'd30348});
	test_expansion(128'hef4b1561547395759007689c1e20e6d1, {16'd51743, 16'd40192, 16'd32297, 16'd54342, 16'd20635, 16'd34450, 16'd19802, 16'd32236, 16'd2276, 16'd17558, 16'd50950, 16'd42751, 16'd48706, 16'd16209, 16'd244, 16'd23128, 16'd23206, 16'd2174, 16'd16210, 16'd29605, 16'd41800, 16'd37274, 16'd158, 16'd17543, 16'd32813, 16'd58470});
	test_expansion(128'h590f3f42af0b99ee31886a5b84a1946e, {16'd49034, 16'd44529, 16'd11030, 16'd34181, 16'd41610, 16'd33107, 16'd1822, 16'd28388, 16'd32961, 16'd50338, 16'd38291, 16'd52551, 16'd63425, 16'd18684, 16'd3214, 16'd2061, 16'd54811, 16'd17592, 16'd28089, 16'd57765, 16'd54775, 16'd8312, 16'd14698, 16'd64861, 16'd51070, 16'd10889});
	test_expansion(128'hffe5c147e1538e5d50a39fd674dadb59, {16'd29530, 16'd16576, 16'd15892, 16'd45795, 16'd43693, 16'd50294, 16'd33251, 16'd17403, 16'd31174, 16'd1479, 16'd19884, 16'd54320, 16'd42524, 16'd24172, 16'd29338, 16'd72, 16'd15282, 16'd8848, 16'd18256, 16'd40320, 16'd61779, 16'd40409, 16'd51305, 16'd5554, 16'd54596, 16'd15028});
	test_expansion(128'h5b82fb1d2d64482ac3ef0a55466c54e5, {16'd15833, 16'd14716, 16'd23826, 16'd5137, 16'd31466, 16'd48174, 16'd31512, 16'd5613, 16'd41626, 16'd50416, 16'd27537, 16'd14237, 16'd41673, 16'd31308, 16'd56747, 16'd58604, 16'd37257, 16'd47248, 16'd46446, 16'd14224, 16'd64820, 16'd4872, 16'd60694, 16'd15101, 16'd60895, 16'd51978});
	test_expansion(128'h1f8159f3910807956f2d4bb61771b5b0, {16'd24366, 16'd10560, 16'd14319, 16'd35383, 16'd42199, 16'd63967, 16'd34988, 16'd60069, 16'd31768, 16'd44569, 16'd8583, 16'd4346, 16'd64071, 16'd15973, 16'd6711, 16'd45972, 16'd41364, 16'd62960, 16'd53681, 16'd1488, 16'd47172, 16'd48788, 16'd46655, 16'd5908, 16'd31722, 16'd3706});
	test_expansion(128'h780f92118b963e52c0968815dfb53ed0, {16'd60924, 16'd45034, 16'd59819, 16'd26212, 16'd29398, 16'd21856, 16'd47344, 16'd61726, 16'd31958, 16'd42670, 16'd36520, 16'd48282, 16'd63524, 16'd37071, 16'd24733, 16'd1205, 16'd35908, 16'd38028, 16'd33206, 16'd10760, 16'd48915, 16'd25494, 16'd54570, 16'd23413, 16'd15351, 16'd26011});
	test_expansion(128'ha86ae319bd29e220f30b184be05d155a, {16'd48590, 16'd7363, 16'd15467, 16'd3024, 16'd54991, 16'd7340, 16'd18859, 16'd57370, 16'd25307, 16'd21650, 16'd50759, 16'd30760, 16'd8641, 16'd51460, 16'd12791, 16'd24097, 16'd16464, 16'd47404, 16'd53281, 16'd12540, 16'd40596, 16'd49915, 16'd6012, 16'd4652, 16'd53826, 16'd30563});
	test_expansion(128'h105fca3736e16af957b679e62aa12d5f, {16'd30767, 16'd45132, 16'd64305, 16'd58209, 16'd39451, 16'd18101, 16'd24333, 16'd63999, 16'd18232, 16'd18461, 16'd35489, 16'd15136, 16'd40200, 16'd55229, 16'd47456, 16'd39319, 16'd4399, 16'd63361, 16'd9283, 16'd47212, 16'd3011, 16'd58391, 16'd23393, 16'd61840, 16'd23642, 16'd47992});
	test_expansion(128'h6ba17eebb9de298071fbde17dc3a42c6, {16'd1504, 16'd21330, 16'd20395, 16'd58561, 16'd24932, 16'd7990, 16'd53872, 16'd17178, 16'd43545, 16'd11584, 16'd39543, 16'd58706, 16'd44783, 16'd14223, 16'd43939, 16'd23846, 16'd24473, 16'd56634, 16'd50975, 16'd7433, 16'd25372, 16'd44128, 16'd20202, 16'd22453, 16'd3910, 16'd15468});
	test_expansion(128'hb276431f86fab1cbcc41fed2c78b873b, {16'd56450, 16'd31980, 16'd43844, 16'd16108, 16'd14151, 16'd26845, 16'd41054, 16'd32933, 16'd39266, 16'd38860, 16'd22550, 16'd8770, 16'd39061, 16'd412, 16'd24031, 16'd42993, 16'd49145, 16'd10441, 16'd37924, 16'd19204, 16'd5609, 16'd52699, 16'd4314, 16'd62897, 16'd59081, 16'd52479});
	test_expansion(128'hf46612966f8cd06fc0d930f414bda7be, {16'd23178, 16'd57827, 16'd20147, 16'd13620, 16'd11957, 16'd35146, 16'd2676, 16'd44366, 16'd36632, 16'd15317, 16'd1806, 16'd7074, 16'd48608, 16'd44086, 16'd24861, 16'd54650, 16'd63230, 16'd245, 16'd64553, 16'd33474, 16'd23782, 16'd59722, 16'd59477, 16'd2567, 16'd26446, 16'd59132});
	test_expansion(128'hdaa2cc2f6e05f7a3c342c77fe443acc1, {16'd39968, 16'd526, 16'd52626, 16'd35930, 16'd51896, 16'd62811, 16'd51634, 16'd25930, 16'd52941, 16'd8411, 16'd33494, 16'd142, 16'd55762, 16'd64417, 16'd49648, 16'd49982, 16'd2220, 16'd52707, 16'd42550, 16'd52133, 16'd51163, 16'd20406, 16'd7872, 16'd43081, 16'd59217, 16'd54946});
	test_expansion(128'h0c750e6b4d37295fcd45626d5d6ab899, {16'd8969, 16'd112, 16'd16847, 16'd2365, 16'd10521, 16'd54242, 16'd39948, 16'd54270, 16'd8678, 16'd33529, 16'd56555, 16'd64866, 16'd26847, 16'd14228, 16'd38057, 16'd61957, 16'd40950, 16'd7340, 16'd29515, 16'd9355, 16'd4552, 16'd52932, 16'd55664, 16'd30273, 16'd65207, 16'd57011});
	test_expansion(128'h8131fe1991ae77b52dfb9a9bc1a62a94, {16'd16779, 16'd44917, 16'd21099, 16'd1233, 16'd11068, 16'd62174, 16'd65490, 16'd27463, 16'd64392, 16'd22759, 16'd52222, 16'd8713, 16'd50805, 16'd35701, 16'd1832, 16'd15153, 16'd31500, 16'd32121, 16'd47790, 16'd35773, 16'd40056, 16'd38800, 16'd42628, 16'd18774, 16'd50447, 16'd20833});
	test_expansion(128'hec6d4db0515faadc149dc51332e3716d, {16'd33511, 16'd25701, 16'd28724, 16'd21699, 16'd18811, 16'd40677, 16'd57955, 16'd27294, 16'd10380, 16'd19923, 16'd25206, 16'd47090, 16'd34261, 16'd18741, 16'd8373, 16'd16574, 16'd52711, 16'd43258, 16'd4241, 16'd31534, 16'd64334, 16'd11778, 16'd42450, 16'd18769, 16'd57615, 16'd18038});
	test_expansion(128'h03d250bac5e346afd58cd2f685ab42e0, {16'd38255, 16'd30075, 16'd63364, 16'd6291, 16'd43892, 16'd13632, 16'd37201, 16'd44965, 16'd58921, 16'd7496, 16'd40217, 16'd26317, 16'd53820, 16'd51899, 16'd58858, 16'd8441, 16'd9530, 16'd21273, 16'd1905, 16'd17780, 16'd64746, 16'd33352, 16'd21951, 16'd32568, 16'd28137, 16'd17208});
	test_expansion(128'h10c72a33f40ba639c94cf23c43799a08, {16'd21408, 16'd35164, 16'd44964, 16'd48061, 16'd21263, 16'd26804, 16'd43487, 16'd18564, 16'd54173, 16'd51658, 16'd58024, 16'd38842, 16'd63865, 16'd25177, 16'd39745, 16'd49644, 16'd15300, 16'd51493, 16'd36922, 16'd16738, 16'd21999, 16'd51134, 16'd47068, 16'd31689, 16'd25368, 16'd31855});
	test_expansion(128'he46b483655a89d44747f29fe65b26b8b, {16'd57137, 16'd38049, 16'd62419, 16'd31811, 16'd3497, 16'd4231, 16'd9212, 16'd56172, 16'd506, 16'd10933, 16'd31259, 16'd56641, 16'd10095, 16'd38750, 16'd60789, 16'd13394, 16'd32674, 16'd18714, 16'd37398, 16'd9284, 16'd63860, 16'd19497, 16'd48107, 16'd27200, 16'd55803, 16'd4095});
	test_expansion(128'h85cb4830b8c290ab03eaab8ac5715fd4, {16'd3626, 16'd52740, 16'd31278, 16'd44222, 16'd38408, 16'd43094, 16'd19845, 16'd30642, 16'd19362, 16'd49620, 16'd61667, 16'd19425, 16'd45073, 16'd62282, 16'd21926, 16'd25867, 16'd54634, 16'd12898, 16'd51712, 16'd57444, 16'd2922, 16'd10700, 16'd62705, 16'd9261, 16'd62900, 16'd36386});
	test_expansion(128'h4151f6adaf3ec76f5b124365861d1db9, {16'd24242, 16'd8615, 16'd12832, 16'd59614, 16'd29959, 16'd1797, 16'd51752, 16'd32413, 16'd57428, 16'd30141, 16'd37321, 16'd30278, 16'd29682, 16'd31901, 16'd3259, 16'd54943, 16'd22834, 16'd10734, 16'd49856, 16'd26650, 16'd14062, 16'd21728, 16'd7523, 16'd18366, 16'd47771, 16'd2306});
	test_expansion(128'hc7550e58d72d25360f21f321305cdb3d, {16'd27174, 16'd19232, 16'd15356, 16'd5921, 16'd59872, 16'd11912, 16'd3751, 16'd46813, 16'd62285, 16'd22063, 16'd27003, 16'd41713, 16'd49165, 16'd10933, 16'd35835, 16'd28506, 16'd34387, 16'd22417, 16'd34288, 16'd62297, 16'd41077, 16'd43631, 16'd8969, 16'd42823, 16'd4961, 16'd12306});
	test_expansion(128'h79d6199f57c7a8dae0cadf6b48d9ba87, {16'd36365, 16'd18072, 16'd52189, 16'd9354, 16'd672, 16'd43235, 16'd9044, 16'd23124, 16'd1763, 16'd30600, 16'd20420, 16'd34585, 16'd40715, 16'd57753, 16'd64097, 16'd24306, 16'd45633, 16'd52765, 16'd27614, 16'd35919, 16'd17885, 16'd31442, 16'd20962, 16'd6930, 16'd61988, 16'd30827});
	test_expansion(128'he155e04766357b4415d3ea73504d8fdc, {16'd40835, 16'd11037, 16'd33494, 16'd8170, 16'd62861, 16'd14446, 16'd19961, 16'd43992, 16'd62864, 16'd10300, 16'd2019, 16'd45463, 16'd23769, 16'd42779, 16'd25453, 16'd47948, 16'd30776, 16'd1954, 16'd22800, 16'd38383, 16'd12381, 16'd12506, 16'd10017, 16'd61747, 16'd21525, 16'd9024});
	test_expansion(128'h5d3c44ce3e2ea30b125de1b9bb349059, {16'd1181, 16'd62004, 16'd26458, 16'd62021, 16'd35522, 16'd19120, 16'd44014, 16'd39787, 16'd64655, 16'd31949, 16'd9302, 16'd59460, 16'd36415, 16'd16151, 16'd4354, 16'd37748, 16'd64335, 16'd55145, 16'd5558, 16'd23768, 16'd39167, 16'd8314, 16'd34897, 16'd51336, 16'd31464, 16'd62319});
	test_expansion(128'h8b7ae682b4b049e955d79f4f2df28541, {16'd11255, 16'd15121, 16'd13502, 16'd11879, 16'd33712, 16'd38293, 16'd54701, 16'd5574, 16'd38710, 16'd53797, 16'd4257, 16'd43682, 16'd20951, 16'd40182, 16'd64608, 16'd38200, 16'd22388, 16'd17597, 16'd28745, 16'd11806, 16'd53978, 16'd3323, 16'd62785, 16'd24832, 16'd40383, 16'd21484});
	test_expansion(128'h0e87e02705656bacc1bd03924723c4ba, {16'd37352, 16'd57002, 16'd51177, 16'd3228, 16'd59232, 16'd50282, 16'd34266, 16'd1589, 16'd4315, 16'd57654, 16'd43856, 16'd15024, 16'd38802, 16'd38595, 16'd7703, 16'd44492, 16'd32468, 16'd55027, 16'd46872, 16'd55574, 16'd42383, 16'd14902, 16'd50637, 16'd53509, 16'd61896, 16'd61945});
	test_expansion(128'h60d01eea8837025be1f7c598b20c7998, {16'd24231, 16'd64044, 16'd38921, 16'd45402, 16'd23956, 16'd57855, 16'd29694, 16'd56686, 16'd61141, 16'd5585, 16'd1237, 16'd48674, 16'd60284, 16'd48272, 16'd10408, 16'd12614, 16'd60590, 16'd25329, 16'd45223, 16'd44286, 16'd24120, 16'd16877, 16'd62838, 16'd21814, 16'd22333, 16'd46585});
	test_expansion(128'h0db272b59ab85981a9a4a011ff884826, {16'd57062, 16'd9846, 16'd32698, 16'd7552, 16'd37972, 16'd47739, 16'd36864, 16'd42356, 16'd32192, 16'd58456, 16'd25767, 16'd57364, 16'd44284, 16'd44900, 16'd10266, 16'd1796, 16'd41702, 16'd28462, 16'd55925, 16'd13674, 16'd51805, 16'd44959, 16'd17437, 16'd35893, 16'd60780, 16'd63274});
	test_expansion(128'h629f56721f356442af4cf3a5059b9426, {16'd21269, 16'd39244, 16'd56790, 16'd54435, 16'd30201, 16'd3977, 16'd32316, 16'd53880, 16'd23687, 16'd64132, 16'd59963, 16'd15641, 16'd46050, 16'd5757, 16'd34140, 16'd58409, 16'd16672, 16'd8105, 16'd53664, 16'd45051, 16'd19962, 16'd26704, 16'd10260, 16'd47789, 16'd36294, 16'd13487});
	test_expansion(128'h83a2d64ae56336a63e1d1f9743076a56, {16'd53507, 16'd7094, 16'd35269, 16'd40906, 16'd14982, 16'd28565, 16'd37983, 16'd29171, 16'd54769, 16'd16479, 16'd12623, 16'd45958, 16'd65083, 16'd44576, 16'd37236, 16'd61056, 16'd23433, 16'd33298, 16'd7688, 16'd869, 16'd61630, 16'd56953, 16'd16157, 16'd24749, 16'd39925, 16'd2273});
	test_expansion(128'he338e141e96d591721a7dff48758b358, {16'd60107, 16'd42277, 16'd45218, 16'd296, 16'd29614, 16'd18747, 16'd52225, 16'd27931, 16'd12668, 16'd17700, 16'd51531, 16'd44964, 16'd56827, 16'd12307, 16'd21880, 16'd28369, 16'd59180, 16'd61056, 16'd64373, 16'd19612, 16'd36537, 16'd13709, 16'd34889, 16'd8680, 16'd42690, 16'd60976});
	test_expansion(128'hbdef45c6391ca76cb160e732a51c87dd, {16'd48325, 16'd6757, 16'd54719, 16'd42207, 16'd21326, 16'd62870, 16'd54243, 16'd31944, 16'd23783, 16'd28094, 16'd46554, 16'd13511, 16'd27141, 16'd52834, 16'd46720, 16'd54945, 16'd18104, 16'd63739, 16'd28930, 16'd6539, 16'd16968, 16'd11135, 16'd43943, 16'd12561, 16'd27855, 16'd41768});
	test_expansion(128'h82855fe5953557ff5541b51194bffef7, {16'd9675, 16'd32429, 16'd30849, 16'd58065, 16'd5253, 16'd34696, 16'd8773, 16'd36757, 16'd7997, 16'd48649, 16'd47749, 16'd1228, 16'd4551, 16'd38786, 16'd3285, 16'd44015, 16'd21461, 16'd3777, 16'd55042, 16'd64593, 16'd54967, 16'd22465, 16'd39314, 16'd62393, 16'd55436, 16'd22058});
	test_expansion(128'hb715d81b0c6944cc05f8489fa11e2c1a, {16'd28475, 16'd64782, 16'd61489, 16'd56365, 16'd17691, 16'd59868, 16'd5651, 16'd15385, 16'd4029, 16'd10055, 16'd27775, 16'd7918, 16'd54186, 16'd24398, 16'd25750, 16'd27431, 16'd45624, 16'd54232, 16'd26147, 16'd17496, 16'd3387, 16'd52369, 16'd6766, 16'd52324, 16'd12564, 16'd50663});
	test_expansion(128'h05a257588a42f04015cd39b2e4230254, {16'd44239, 16'd12788, 16'd1783, 16'd44792, 16'd16117, 16'd22758, 16'd27874, 16'd25924, 16'd15775, 16'd63137, 16'd8770, 16'd64340, 16'd57414, 16'd6043, 16'd54682, 16'd54780, 16'd8960, 16'd48897, 16'd29169, 16'd45963, 16'd4316, 16'd57537, 16'd15802, 16'd38676, 16'd31574, 16'd32918});
	test_expansion(128'h5f220029f92e552d516c1415f199b472, {16'd3455, 16'd12608, 16'd24794, 16'd21233, 16'd20072, 16'd14647, 16'd58185, 16'd11653, 16'd27541, 16'd21843, 16'd40090, 16'd53711, 16'd6549, 16'd4998, 16'd13504, 16'd5150, 16'd48137, 16'd38914, 16'd36620, 16'd45407, 16'd37727, 16'd41906, 16'd25862, 16'd17262, 16'd65445, 16'd28654});
	test_expansion(128'hd1dd09bfc2a861adacbfa724dc01ddbc, {16'd36958, 16'd28240, 16'd12268, 16'd32219, 16'd40526, 16'd54297, 16'd27435, 16'd22039, 16'd46405, 16'd55377, 16'd56108, 16'd27857, 16'd45771, 16'd2949, 16'd65413, 16'd13032, 16'd15438, 16'd28701, 16'd32756, 16'd21500, 16'd9831, 16'd31455, 16'd29796, 16'd23877, 16'd6401, 16'd49488});
	test_expansion(128'h6c5660e2a7cee0a941ec341d692431d2, {16'd64571, 16'd42804, 16'd32038, 16'd29652, 16'd52260, 16'd29036, 16'd22433, 16'd57768, 16'd8120, 16'd62696, 16'd28345, 16'd10472, 16'd533, 16'd36798, 16'd30377, 16'd33134, 16'd65043, 16'd45870, 16'd37043, 16'd44351, 16'd14920, 16'd31030, 16'd5130, 16'd34919, 16'd5825, 16'd38478});
	test_expansion(128'hf10f87bddbe4870f71e03a0724d6ae8f, {16'd34437, 16'd52889, 16'd54500, 16'd40357, 16'd64818, 16'd25528, 16'd8546, 16'd9265, 16'd48992, 16'd31837, 16'd18640, 16'd49365, 16'd10991, 16'd3772, 16'd34460, 16'd2040, 16'd34880, 16'd49541, 16'd1928, 16'd40059, 16'd13591, 16'd46548, 16'd33763, 16'd55169, 16'd17679, 16'd17606});
	test_expansion(128'h132cb92b6927a85cc2a880a35535b217, {16'd40825, 16'd50082, 16'd11338, 16'd57784, 16'd60267, 16'd7573, 16'd14209, 16'd15229, 16'd39928, 16'd61855, 16'd52751, 16'd32848, 16'd21428, 16'd2003, 16'd44941, 16'd40545, 16'd31372, 16'd55548, 16'd29658, 16'd32266, 16'd48934, 16'd57580, 16'd20721, 16'd11091, 16'd7571, 16'd49853});
	test_expansion(128'hff4f684dd33bd925122960b2e3a519e5, {16'd1236, 16'd47031, 16'd62444, 16'd9434, 16'd35058, 16'd7816, 16'd4053, 16'd2677, 16'd56779, 16'd46264, 16'd5865, 16'd39659, 16'd25050, 16'd48192, 16'd56227, 16'd53142, 16'd4627, 16'd3349, 16'd36234, 16'd4897, 16'd59959, 16'd27893, 16'd31937, 16'd26957, 16'd29618, 16'd47439});
	test_expansion(128'h79983c04b2be6cfe8b547118acba296a, {16'd50562, 16'd24569, 16'd10281, 16'd25949, 16'd16332, 16'd14756, 16'd47830, 16'd50132, 16'd14395, 16'd43817, 16'd11355, 16'd28682, 16'd19572, 16'd59182, 16'd6320, 16'd6813, 16'd34837, 16'd60241, 16'd46784, 16'd46698, 16'd24516, 16'd37011, 16'd32479, 16'd14131, 16'd62270, 16'd18311});
	test_expansion(128'h4612fef66eb879cd6d116acaf5b504d1, {16'd59565, 16'd8094, 16'd4590, 16'd23992, 16'd24279, 16'd55533, 16'd23904, 16'd17632, 16'd51095, 16'd47627, 16'd48853, 16'd42312, 16'd55236, 16'd60531, 16'd20401, 16'd56483, 16'd60483, 16'd53430, 16'd34498, 16'd65143, 16'd8412, 16'd13879, 16'd44850, 16'd56421, 16'd29795, 16'd8594});
	test_expansion(128'h7e751043f77c25a6f17488584ff850cf, {16'd60068, 16'd64707, 16'd40336, 16'd34392, 16'd15716, 16'd44558, 16'd47461, 16'd43851, 16'd10155, 16'd63484, 16'd36785, 16'd4548, 16'd32069, 16'd26322, 16'd32587, 16'd1252, 16'd30761, 16'd60070, 16'd11106, 16'd61215, 16'd24505, 16'd18673, 16'd40539, 16'd31967, 16'd18936, 16'd838});
	test_expansion(128'hdb726bf13652944e5497a2fffd3ddf37, {16'd31209, 16'd59281, 16'd13032, 16'd31533, 16'd9397, 16'd5623, 16'd46447, 16'd56939, 16'd62810, 16'd1507, 16'd38017, 16'd32597, 16'd26596, 16'd31028, 16'd54919, 16'd39883, 16'd55650, 16'd45405, 16'd38535, 16'd25528, 16'd54155, 16'd8280, 16'd21336, 16'd52329, 16'd22516, 16'd52607});
	test_expansion(128'hb881aa65f9a09774232b7fd38329b477, {16'd56637, 16'd31491, 16'd32128, 16'd22196, 16'd38894, 16'd61612, 16'd14869, 16'd61549, 16'd9734, 16'd8151, 16'd36110, 16'd41290, 16'd44406, 16'd39941, 16'd26758, 16'd56557, 16'd23877, 16'd20141, 16'd61844, 16'd18982, 16'd10620, 16'd1978, 16'd3750, 16'd47441, 16'd62820, 16'd48476});
	test_expansion(128'hbcea9e259e6a938465088471b0ccbdd7, {16'd8163, 16'd16036, 16'd53316, 16'd27117, 16'd58234, 16'd54966, 16'd5452, 16'd31705, 16'd11901, 16'd26172, 16'd16635, 16'd8558, 16'd44467, 16'd37603, 16'd27238, 16'd31494, 16'd30565, 16'd62832, 16'd17710, 16'd64433, 16'd42006, 16'd36012, 16'd62763, 16'd40909, 16'd10814, 16'd52814});
	test_expansion(128'h892b9accce9e30b58aa6db2f89da9b42, {16'd18822, 16'd40092, 16'd32437, 16'd53324, 16'd13760, 16'd29475, 16'd34489, 16'd64652, 16'd58513, 16'd30331, 16'd38694, 16'd36250, 16'd18994, 16'd40493, 16'd57485, 16'd40770, 16'd60667, 16'd313, 16'd41158, 16'd5928, 16'd52793, 16'd60553, 16'd15403, 16'd9481, 16'd40373, 16'd29832});
	test_expansion(128'h2f9126a71b6b404da289105d45bfeef1, {16'd65275, 16'd7338, 16'd51790, 16'd37243, 16'd26420, 16'd9468, 16'd46475, 16'd31819, 16'd6552, 16'd64451, 16'd32710, 16'd46021, 16'd33343, 16'd20639, 16'd7679, 16'd16704, 16'd56099, 16'd27592, 16'd3789, 16'd4710, 16'd40636, 16'd24607, 16'd56038, 16'd45824, 16'd61931, 16'd41683});
	test_expansion(128'h9282b1fbd0d16f199c6a2298e3983afc, {16'd45107, 16'd15044, 16'd63279, 16'd28803, 16'd16419, 16'd54940, 16'd23297, 16'd7105, 16'd55857, 16'd8090, 16'd41160, 16'd22634, 16'd52833, 16'd28169, 16'd59224, 16'd40304, 16'd39994, 16'd13216, 16'd2680, 16'd46967, 16'd55449, 16'd19668, 16'd20299, 16'd8311, 16'd7244, 16'd57483});
	test_expansion(128'h6db213e08066a720aaab60395233261f, {16'd31042, 16'd50894, 16'd5642, 16'd22451, 16'd31171, 16'd1157, 16'd38363, 16'd25330, 16'd5035, 16'd31886, 16'd61429, 16'd44540, 16'd38052, 16'd15213, 16'd22933, 16'd35607, 16'd1842, 16'd55690, 16'd14336, 16'd28709, 16'd9395, 16'd3293, 16'd9680, 16'd847, 16'd49701, 16'd8186});
	test_expansion(128'hb5ad76a8fc66649b8b9d33321d784b83, {16'd15241, 16'd61918, 16'd13610, 16'd64608, 16'd54373, 16'd9665, 16'd11299, 16'd35562, 16'd20625, 16'd64306, 16'd63630, 16'd23432, 16'd34369, 16'd45870, 16'd31576, 16'd30460, 16'd59975, 16'd24830, 16'd19362, 16'd32559, 16'd29700, 16'd47622, 16'd38192, 16'd14483, 16'd12456, 16'd40531});
	test_expansion(128'h86ef8fde41404c5401526347d88097ea, {16'd13208, 16'd38989, 16'd26490, 16'd60334, 16'd17801, 16'd2623, 16'd12765, 16'd154, 16'd60990, 16'd42033, 16'd27290, 16'd5935, 16'd56204, 16'd9971, 16'd16051, 16'd1226, 16'd28520, 16'd64444, 16'd43807, 16'd39479, 16'd61923, 16'd36985, 16'd210, 16'd7911, 16'd12953, 16'd19972});
	test_expansion(128'h433f82764ff0fd7b30c294f00619ee22, {16'd31535, 16'd30926, 16'd29776, 16'd13267, 16'd6173, 16'd6546, 16'd40428, 16'd17938, 16'd26135, 16'd47172, 16'd47481, 16'd57264, 16'd45202, 16'd15664, 16'd43834, 16'd26740, 16'd55253, 16'd33730, 16'd51208, 16'd23795, 16'd11391, 16'd11275, 16'd15040, 16'd14415, 16'd6518, 16'd41279});
	test_expansion(128'hf7e2601d9099ec3e97ee827b0799d167, {16'd23263, 16'd58948, 16'd29768, 16'd61949, 16'd42835, 16'd567, 16'd15419, 16'd37796, 16'd28818, 16'd11940, 16'd9136, 16'd8806, 16'd4560, 16'd58284, 16'd62494, 16'd17458, 16'd19547, 16'd59965, 16'd46637, 16'd43539, 16'd27322, 16'd19876, 16'd24171, 16'd31175, 16'd12940, 16'd12960});
	test_expansion(128'h5d5676aedc98222c5af5071d5c2e1136, {16'd4167, 16'd32145, 16'd61814, 16'd4911, 16'd16967, 16'd51840, 16'd3942, 16'd33788, 16'd49747, 16'd34978, 16'd53290, 16'd64616, 16'd2810, 16'd43479, 16'd31954, 16'd53924, 16'd55602, 16'd50251, 16'd29309, 16'd592, 16'd50222, 16'd9459, 16'd63102, 16'd42618, 16'd51340, 16'd4615});
	test_expansion(128'haf65102bfc617f6ce54d43c443ad70fa, {16'd29350, 16'd33414, 16'd60866, 16'd3565, 16'd56271, 16'd19383, 16'd3473, 16'd792, 16'd6249, 16'd13162, 16'd45627, 16'd28530, 16'd57493, 16'd33289, 16'd8796, 16'd35792, 16'd51574, 16'd40151, 16'd59881, 16'd39950, 16'd57396, 16'd14417, 16'd33361, 16'd39968, 16'd60057, 16'd21167});
	test_expansion(128'h7977249a2c0d39f385804249db5c130f, {16'd58849, 16'd51518, 16'd43663, 16'd16743, 16'd8312, 16'd28644, 16'd25337, 16'd20354, 16'd20623, 16'd32747, 16'd43241, 16'd13236, 16'd16606, 16'd24473, 16'd50088, 16'd22974, 16'd21125, 16'd63846, 16'd26785, 16'd42787, 16'd7334, 16'd1081, 16'd28398, 16'd23761, 16'd52055, 16'd515});
	test_expansion(128'h7f96869a959a5fbdd86a2f261cad4639, {16'd26842, 16'd1294, 16'd16021, 16'd11633, 16'd11935, 16'd62477, 16'd31377, 16'd35035, 16'd42637, 16'd23421, 16'd8211, 16'd5426, 16'd25713, 16'd32076, 16'd34486, 16'd45106, 16'd54292, 16'd27382, 16'd14271, 16'd46756, 16'd36813, 16'd28851, 16'd4805, 16'd8967, 16'd45529, 16'd8286});
	test_expansion(128'h0a78ba5173af52d250d3870059252bb5, {16'd2946, 16'd11523, 16'd43690, 16'd51431, 16'd65039, 16'd41411, 16'd47268, 16'd35788, 16'd28151, 16'd60434, 16'd55816, 16'd1629, 16'd5233, 16'd9533, 16'd39666, 16'd28313, 16'd25010, 16'd22706, 16'd44898, 16'd52929, 16'd25827, 16'd23670, 16'd23238, 16'd370, 16'd57222, 16'd39410});
	test_expansion(128'hb25e142126e0581132a85a91d6cab521, {16'd10387, 16'd18694, 16'd61127, 16'd31312, 16'd21611, 16'd27415, 16'd4891, 16'd47337, 16'd45946, 16'd49747, 16'd41388, 16'd21631, 16'd43096, 16'd31031, 16'd37791, 16'd50259, 16'd534, 16'd20659, 16'd32178, 16'd42571, 16'd25909, 16'd29714, 16'd16619, 16'd15137, 16'd38156, 16'd4849});
	test_expansion(128'h0181e5977233de605a78165eccc213e5, {16'd45914, 16'd50008, 16'd53500, 16'd56383, 16'd10731, 16'd22968, 16'd39879, 16'd18858, 16'd41598, 16'd3655, 16'd24275, 16'd30443, 16'd48870, 16'd45671, 16'd56071, 16'd17705, 16'd29449, 16'd62031, 16'd33453, 16'd13678, 16'd4362, 16'd36215, 16'd56431, 16'd57223, 16'd1876, 16'd18928});
	test_expansion(128'h45e40f527edb10b7b3f39edf861e4bdd, {16'd46637, 16'd10027, 16'd1959, 16'd54, 16'd15982, 16'd56755, 16'd53102, 16'd19388, 16'd42378, 16'd53650, 16'd53069, 16'd55268, 16'd6246, 16'd11575, 16'd40851, 16'd29025, 16'd2855, 16'd43813, 16'd16520, 16'd38780, 16'd61009, 16'd41260, 16'd55562, 16'd39311, 16'd54338, 16'd63243});
	test_expansion(128'h85ebd81e01833730c91720f60533cff0, {16'd41653, 16'd11067, 16'd46993, 16'd35471, 16'd2618, 16'd9638, 16'd60804, 16'd17017, 16'd53374, 16'd59681, 16'd10721, 16'd26417, 16'd34848, 16'd53311, 16'd41237, 16'd40831, 16'd26680, 16'd48318, 16'd10334, 16'd62200, 16'd20673, 16'd34369, 16'd5262, 16'd21220, 16'd28974, 16'd60485});
	test_expansion(128'hbbea7ed5d200bbf7cfde217c24b2efc1, {16'd371, 16'd56705, 16'd6784, 16'd59173, 16'd54118, 16'd11152, 16'd50040, 16'd26704, 16'd19379, 16'd18461, 16'd26577, 16'd8817, 16'd999, 16'd56246, 16'd24510, 16'd45478, 16'd34278, 16'd42937, 16'd7542, 16'd37514, 16'd25865, 16'd33283, 16'd50774, 16'd2005, 16'd22762, 16'd22014});
	test_expansion(128'h31c72e190b5856a30b383e873c710ce4, {16'd46901, 16'd46241, 16'd2658, 16'd58407, 16'd65405, 16'd46371, 16'd25197, 16'd34838, 16'd31441, 16'd12218, 16'd32472, 16'd3863, 16'd46808, 16'd10435, 16'd27123, 16'd32799, 16'd32587, 16'd55657, 16'd58995, 16'd40567, 16'd59417, 16'd30126, 16'd37166, 16'd45844, 16'd40200, 16'd26506});
	test_expansion(128'hb1e1fabe0d5d26339ff3fd6007bd85e2, {16'd54269, 16'd5374, 16'd65069, 16'd45559, 16'd61203, 16'd6234, 16'd28122, 16'd6556, 16'd44154, 16'd44989, 16'd58564, 16'd4610, 16'd58012, 16'd31016, 16'd16594, 16'd8382, 16'd52309, 16'd1283, 16'd45186, 16'd41524, 16'd3044, 16'd37310, 16'd39282, 16'd37133, 16'd60642, 16'd62165});
	test_expansion(128'h804453692a432527869b97bb85f5e31e, {16'd42207, 16'd49290, 16'd6133, 16'd3171, 16'd40351, 16'd20942, 16'd13349, 16'd61737, 16'd46704, 16'd25966, 16'd5762, 16'd31050, 16'd4451, 16'd34493, 16'd41201, 16'd7213, 16'd47216, 16'd3562, 16'd29655, 16'd15763, 16'd14203, 16'd25613, 16'd10294, 16'd21336, 16'd23162, 16'd58881});
	test_expansion(128'h39f594b96bfd515c4b6466a11b817e94, {16'd30385, 16'd61830, 16'd25405, 16'd36300, 16'd63408, 16'd25968, 16'd34340, 16'd7593, 16'd15414, 16'd60966, 16'd53150, 16'd46936, 16'd8681, 16'd45266, 16'd18780, 16'd29502, 16'd13166, 16'd5829, 16'd50442, 16'd16397, 16'd62986, 16'd28986, 16'd17977, 16'd57691, 16'd29776, 16'd52345});
	test_expansion(128'hde711edb93072d3306f30945da92e409, {16'd61618, 16'd1846, 16'd33095, 16'd2176, 16'd56235, 16'd46323, 16'd18092, 16'd15607, 16'd53382, 16'd27018, 16'd42972, 16'd16587, 16'd34931, 16'd51689, 16'd23165, 16'd33090, 16'd39190, 16'd16028, 16'd31465, 16'd30111, 16'd1353, 16'd33091, 16'd44128, 16'd21316, 16'd9602, 16'd31347});
	test_expansion(128'hcbce7167e6f1eb5a61dd702b84c4af51, {16'd57206, 16'd13811, 16'd41067, 16'd38070, 16'd10877, 16'd35722, 16'd17342, 16'd7000, 16'd28265, 16'd6265, 16'd1678, 16'd1671, 16'd23474, 16'd30021, 16'd32389, 16'd14667, 16'd35984, 16'd35677, 16'd16196, 16'd42232, 16'd43640, 16'd9357, 16'd62902, 16'd48460, 16'd57004, 16'd1817});
	test_expansion(128'hee8899198ee837eda9b9a97576f2d023, {16'd44563, 16'd51987, 16'd24280, 16'd745, 16'd59331, 16'd23151, 16'd42563, 16'd31113, 16'd13515, 16'd22791, 16'd12104, 16'd62001, 16'd37808, 16'd53493, 16'd53454, 16'd12119, 16'd2990, 16'd9494, 16'd4568, 16'd10421, 16'd46150, 16'd36607, 16'd4610, 16'd55603, 16'd54170, 16'd43188});
	test_expansion(128'hb4ba1311c8c6d07115baa2665bb4cd87, {16'd65034, 16'd61358, 16'd652, 16'd44811, 16'd62676, 16'd52762, 16'd44214, 16'd25027, 16'd40770, 16'd45310, 16'd9403, 16'd7145, 16'd19529, 16'd42021, 16'd39192, 16'd13671, 16'd51401, 16'd45563, 16'd11317, 16'd38211, 16'd49467, 16'd55960, 16'd39894, 16'd33091, 16'd47416, 16'd65088});
	test_expansion(128'h6add579fbaef58b72817f90ae9b2d6e6, {16'd25958, 16'd24516, 16'd5969, 16'd30729, 16'd27038, 16'd63448, 16'd44861, 16'd62667, 16'd48644, 16'd53480, 16'd9104, 16'd57885, 16'd33770, 16'd32747, 16'd44781, 16'd26283, 16'd8913, 16'd54637, 16'd7671, 16'd45331, 16'd43503, 16'd51745, 16'd57945, 16'd64080, 16'd45166, 16'd7995});
	test_expansion(128'ha2828cecf496b24b8082978e05f53f12, {16'd51167, 16'd40432, 16'd51478, 16'd19129, 16'd19853, 16'd43202, 16'd18992, 16'd19708, 16'd22199, 16'd18495, 16'd52420, 16'd22825, 16'd54718, 16'd24750, 16'd8871, 16'd23357, 16'd18579, 16'd61334, 16'd9464, 16'd10723, 16'd65076, 16'd61073, 16'd26572, 16'd12764, 16'd42585, 16'd153});
	test_expansion(128'h3e995ded6df50107ba3dca71bc696638, {16'd18914, 16'd24090, 16'd9945, 16'd59920, 16'd41308, 16'd53475, 16'd12562, 16'd439, 16'd11843, 16'd29347, 16'd36395, 16'd23938, 16'd15454, 16'd6617, 16'd44778, 16'd26617, 16'd55272, 16'd18113, 16'd21792, 16'd49673, 16'd62778, 16'd27417, 16'd59113, 16'd1155, 16'd36352, 16'd32140});
	test_expansion(128'hdbbd840bf781bd0f59b436882a297413, {16'd61645, 16'd17743, 16'd42956, 16'd62038, 16'd54026, 16'd55357, 16'd25352, 16'd14776, 16'd16758, 16'd41909, 16'd1982, 16'd55826, 16'd59303, 16'd8280, 16'd40045, 16'd49441, 16'd31909, 16'd63125, 16'd61191, 16'd42747, 16'd7285, 16'd43600, 16'd42183, 16'd53377, 16'd9962, 16'd41287});
	test_expansion(128'hd87ccf5410452647f6c169191932d088, {16'd5846, 16'd42652, 16'd54144, 16'd64958, 16'd48468, 16'd15826, 16'd2025, 16'd53056, 16'd60846, 16'd8669, 16'd58950, 16'd12785, 16'd62034, 16'd25610, 16'd8818, 16'd44575, 16'd42975, 16'd59515, 16'd58239, 16'd6118, 16'd3186, 16'd52373, 16'd26610, 16'd5890, 16'd6464, 16'd9544});
	test_expansion(128'hd8018a63304920a3f9fba4c55dd7d226, {16'd62756, 16'd46760, 16'd61753, 16'd46126, 16'd7301, 16'd22741, 16'd8302, 16'd10524, 16'd5571, 16'd19503, 16'd62412, 16'd37976, 16'd21307, 16'd61226, 16'd50418, 16'd47915, 16'd35504, 16'd43673, 16'd38548, 16'd35376, 16'd613, 16'd796, 16'd33675, 16'd14676, 16'd37070, 16'd8426});
	test_expansion(128'hf7b8d7107555ec01558807552619202d, {16'd38483, 16'd48704, 16'd220, 16'd40977, 16'd59824, 16'd537, 16'd945, 16'd52879, 16'd4162, 16'd3743, 16'd33647, 16'd85, 16'd51716, 16'd17714, 16'd53187, 16'd41065, 16'd45378, 16'd18025, 16'd52297, 16'd41811, 16'd46501, 16'd21249, 16'd43669, 16'd20693, 16'd31478, 16'd50977});
	test_expansion(128'h4db69707f509ea1ed6577b1b3a8a0dde, {16'd92, 16'd21191, 16'd57078, 16'd60077, 16'd28592, 16'd40365, 16'd44488, 16'd31225, 16'd34979, 16'd3641, 16'd48310, 16'd59727, 16'd40750, 16'd37335, 16'd20571, 16'd10649, 16'd15159, 16'd22523, 16'd7434, 16'd12672, 16'd42317, 16'd43669, 16'd60131, 16'd26163, 16'd27657, 16'd17892});
	test_expansion(128'h0af182246e5fcca1a13daa8e886b27d7, {16'd28030, 16'd33489, 16'd56341, 16'd21696, 16'd19923, 16'd31748, 16'd29639, 16'd27974, 16'd59976, 16'd13046, 16'd11031, 16'd23954, 16'd12631, 16'd16689, 16'd49599, 16'd55774, 16'd27920, 16'd55493, 16'd33974, 16'd36584, 16'd10037, 16'd36470, 16'd43323, 16'd38804, 16'd23656, 16'd29459});
	test_expansion(128'hf66a74f8b4a66f5ad3aafc465a119d14, {16'd56036, 16'd64799, 16'd49430, 16'd13981, 16'd48177, 16'd41536, 16'd53329, 16'd55401, 16'd12284, 16'd10513, 16'd299, 16'd42358, 16'd30302, 16'd44739, 16'd6437, 16'd46633, 16'd14562, 16'd52207, 16'd34707, 16'd60337, 16'd54821, 16'd32785, 16'd353, 16'd21720, 16'd54979, 16'd11490});
	test_expansion(128'h4d57a8abbf7f4c5d2985df73f8d74d7f, {16'd32809, 16'd43798, 16'd58595, 16'd55776, 16'd36944, 16'd479, 16'd40061, 16'd20556, 16'd62432, 16'd33294, 16'd21311, 16'd42991, 16'd23955, 16'd12047, 16'd52420, 16'd16458, 16'd29413, 16'd33352, 16'd11533, 16'd25646, 16'd5544, 16'd33946, 16'd42367, 16'd15090, 16'd65345, 16'd45384});
	test_expansion(128'h6cb445db9aec2d9acf382c5156694831, {16'd18415, 16'd25740, 16'd2629, 16'd36610, 16'd47084, 16'd21200, 16'd7013, 16'd29404, 16'd37207, 16'd28207, 16'd49973, 16'd2519, 16'd25210, 16'd36537, 16'd45839, 16'd33794, 16'd35840, 16'd24356, 16'd37756, 16'd51796, 16'd43209, 16'd54067, 16'd56795, 16'd37294, 16'd51139, 16'd30716});
	test_expansion(128'hebca2097a7c437777f83b39c6b6c44b5, {16'd16797, 16'd27758, 16'd38410, 16'd48760, 16'd63628, 16'd47309, 16'd58545, 16'd60533, 16'd44619, 16'd25842, 16'd64566, 16'd58729, 16'd18, 16'd65403, 16'd15194, 16'd40556, 16'd9574, 16'd58179, 16'd33068, 16'd21356, 16'd57666, 16'd6379, 16'd6917, 16'd41075, 16'd63040, 16'd29271});
	test_expansion(128'h6dfd796643575013aa99c70890989b82, {16'd44627, 16'd18589, 16'd27827, 16'd41519, 16'd55442, 16'd12341, 16'd33422, 16'd11067, 16'd46871, 16'd11738, 16'd51577, 16'd34110, 16'd61649, 16'd30962, 16'd49357, 16'd35697, 16'd7139, 16'd61161, 16'd2889, 16'd35097, 16'd44703, 16'd34355, 16'd24783, 16'd8865, 16'd40801, 16'd17836});
	test_expansion(128'h4ba9afd51b99b8fdca3b9153de0975d2, {16'd38245, 16'd65377, 16'd26575, 16'd36387, 16'd18535, 16'd29001, 16'd58969, 16'd15085, 16'd56344, 16'd49099, 16'd40223, 16'd34727, 16'd53185, 16'd63048, 16'd41729, 16'd16030, 16'd15789, 16'd12290, 16'd24116, 16'd4390, 16'd43891, 16'd44449, 16'd59282, 16'd24530, 16'd51790, 16'd38166});
	test_expansion(128'h2cb316f39d8ca0a54782bb43ce36dbdf, {16'd6350, 16'd40706, 16'd59280, 16'd52983, 16'd45590, 16'd33869, 16'd64573, 16'd31532, 16'd31180, 16'd63380, 16'd47644, 16'd62661, 16'd41097, 16'd1443, 16'd62588, 16'd54135, 16'd8405, 16'd64682, 16'd19764, 16'd65424, 16'd39308, 16'd60357, 16'd23737, 16'd1530, 16'd57696, 16'd47225});
	test_expansion(128'h717e5c2695916461f46c595b72c87029, {16'd57859, 16'd15520, 16'd5583, 16'd62816, 16'd36167, 16'd11273, 16'd10226, 16'd21740, 16'd33862, 16'd4405, 16'd37958, 16'd40242, 16'd5465, 16'd4947, 16'd24446, 16'd25378, 16'd19970, 16'd3085, 16'd63909, 16'd33635, 16'd38534, 16'd37229, 16'd5221, 16'd33308, 16'd49856, 16'd41923});
	test_expansion(128'h574e38e2191e3712a947211ee6c7daf1, {16'd61773, 16'd17488, 16'd48381, 16'd28807, 16'd54269, 16'd23774, 16'd9950, 16'd44223, 16'd58334, 16'd38814, 16'd57458, 16'd51890, 16'd51157, 16'd50930, 16'd46329, 16'd60471, 16'd56116, 16'd4381, 16'd25017, 16'd48888, 16'd18527, 16'd33586, 16'd12058, 16'd49981, 16'd28363, 16'd42409});
	test_expansion(128'hfce5a0d08aba8cdf8c6b9deba44c6aea, {16'd25240, 16'd12004, 16'd6341, 16'd15659, 16'd1215, 16'd21422, 16'd34827, 16'd10785, 16'd12866, 16'd40522, 16'd25742, 16'd27805, 16'd60182, 16'd3301, 16'd36889, 16'd39015, 16'd15036, 16'd54347, 16'd47841, 16'd51141, 16'd20183, 16'd34895, 16'd26166, 16'd34563, 16'd24152, 16'd52772});
	test_expansion(128'h1b7981164336f36951edaeccdeedce7d, {16'd35188, 16'd30716, 16'd48545, 16'd19132, 16'd47243, 16'd42653, 16'd24387, 16'd56058, 16'd25277, 16'd36709, 16'd55429, 16'd44628, 16'd31461, 16'd9386, 16'd23255, 16'd11086, 16'd63643, 16'd25034, 16'd50323, 16'd22857, 16'd44677, 16'd42196, 16'd27835, 16'd3796, 16'd22394, 16'd59064});
	test_expansion(128'hff4c51525c15f1c34a323a012c6b5b6a, {16'd49498, 16'd59463, 16'd55449, 16'd50851, 16'd21894, 16'd14079, 16'd37562, 16'd41486, 16'd40175, 16'd8422, 16'd46305, 16'd50956, 16'd10623, 16'd37250, 16'd21494, 16'd1606, 16'd62791, 16'd3212, 16'd48062, 16'd35931, 16'd21818, 16'd53927, 16'd1375, 16'd43871, 16'd55755, 16'd54945});
	test_expansion(128'hcce71d7520404dcfdd4b717e33961f35, {16'd41096, 16'd45772, 16'd18125, 16'd17026, 16'd13725, 16'd23246, 16'd54182, 16'd43568, 16'd49153, 16'd48856, 16'd6912, 16'd62721, 16'd57889, 16'd52457, 16'd4086, 16'd62932, 16'd62159, 16'd16457, 16'd40772, 16'd33945, 16'd62670, 16'd36464, 16'd51016, 16'd32096, 16'd9759, 16'd4914});
	test_expansion(128'h7b0d4ae895cc97fae3dcd574954ae808, {16'd34154, 16'd60410, 16'd14213, 16'd22878, 16'd39156, 16'd33251, 16'd43695, 16'd38409, 16'd37095, 16'd43649, 16'd28327, 16'd19511, 16'd30217, 16'd8018, 16'd16298, 16'd56764, 16'd52444, 16'd16519, 16'd52971, 16'd17083, 16'd30316, 16'd6394, 16'd7064, 16'd1456, 16'd27100, 16'd44419});
	test_expansion(128'h2896387e1f75d2c5aab789641474335c, {16'd47344, 16'd21409, 16'd16194, 16'd597, 16'd15531, 16'd26107, 16'd55145, 16'd30291, 16'd8958, 16'd24783, 16'd51453, 16'd23821, 16'd57040, 16'd3979, 16'd37137, 16'd54738, 16'd41126, 16'd42253, 16'd8082, 16'd33148, 16'd8314, 16'd12930, 16'd26605, 16'd939, 16'd23543, 16'd3315});
	test_expansion(128'h13531487e1e1aa025518cfbe6f4a5427, {16'd18758, 16'd44533, 16'd36802, 16'd54162, 16'd40943, 16'd18695, 16'd33262, 16'd55593, 16'd26271, 16'd24042, 16'd1456, 16'd46486, 16'd1066, 16'd12722, 16'd48891, 16'd28899, 16'd16247, 16'd5375, 16'd63811, 16'd64154, 16'd61562, 16'd24726, 16'd47445, 16'd21386, 16'd5839, 16'd54001});
	test_expansion(128'h41bfe8cabc139217c66c29581dc02ca3, {16'd61212, 16'd22072, 16'd5611, 16'd41493, 16'd46294, 16'd58590, 16'd2071, 16'd7858, 16'd13243, 16'd53780, 16'd65422, 16'd20239, 16'd21779, 16'd30842, 16'd59071, 16'd9202, 16'd38939, 16'd24821, 16'd49383, 16'd9812, 16'd45027, 16'd16559, 16'd4643, 16'd58183, 16'd35881, 16'd10454});
	test_expansion(128'h4b3599525edbd28fd8040f932f4afb6b, {16'd34584, 16'd39931, 16'd59460, 16'd16757, 16'd26365, 16'd55942, 16'd4355, 16'd45980, 16'd51626, 16'd23614, 16'd26930, 16'd6978, 16'd14996, 16'd38576, 16'd45805, 16'd19130, 16'd29625, 16'd30636, 16'd15490, 16'd43718, 16'd32342, 16'd38498, 16'd28253, 16'd36886, 16'd29152, 16'd46507});
	test_expansion(128'h01f60f04bc73a8dffd587772b0fa3131, {16'd39334, 16'd8606, 16'd41964, 16'd30190, 16'd23334, 16'd14978, 16'd35982, 16'd62436, 16'd44523, 16'd40253, 16'd15596, 16'd1175, 16'd21134, 16'd24739, 16'd24573, 16'd63576, 16'd51782, 16'd19953, 16'd15737, 16'd17827, 16'd62069, 16'd53646, 16'd43572, 16'd28389, 16'd541, 16'd17978});
	test_expansion(128'h1c7a2d38e6346da5dae5b94b7485bf43, {16'd24050, 16'd45374, 16'd16045, 16'd1087, 16'd47100, 16'd6772, 16'd60618, 16'd37303, 16'd44135, 16'd39756, 16'd5799, 16'd61194, 16'd12430, 16'd61333, 16'd46783, 16'd48434, 16'd35753, 16'd59381, 16'd58129, 16'd32751, 16'd44818, 16'd20304, 16'd1716, 16'd23383, 16'd39159, 16'd60942});
	test_expansion(128'hdd1e37858312e8a01576b8ae9a191d31, {16'd24575, 16'd23632, 16'd24074, 16'd41176, 16'd17820, 16'd64520, 16'd38012, 16'd65493, 16'd47327, 16'd6986, 16'd19171, 16'd28607, 16'd49136, 16'd24460, 16'd40789, 16'd40676, 16'd16412, 16'd38878, 16'd37694, 16'd58772, 16'd37808, 16'd42817, 16'd7576, 16'd37308, 16'd27936, 16'd47533});
	test_expansion(128'hca9620db9b379e675e06b5ec20a7d5ca, {16'd52693, 16'd28300, 16'd9474, 16'd18696, 16'd47705, 16'd24335, 16'd64525, 16'd15310, 16'd32789, 16'd57114, 16'd57042, 16'd57887, 16'd59877, 16'd56466, 16'd15339, 16'd37071, 16'd53890, 16'd40953, 16'd35759, 16'd52307, 16'd27592, 16'd37866, 16'd16769, 16'd64056, 16'd14841, 16'd32661});
	test_expansion(128'h83fd5b406ba041e701bf1bf3af02fbed, {16'd6745, 16'd46752, 16'd20092, 16'd56474, 16'd13191, 16'd24142, 16'd26654, 16'd3686, 16'd52605, 16'd37771, 16'd49650, 16'd10932, 16'd60916, 16'd48712, 16'd44571, 16'd39361, 16'd47326, 16'd21872, 16'd2662, 16'd44014, 16'd1030, 16'd21409, 16'd59777, 16'd18016, 16'd31403, 16'd58085});
	test_expansion(128'h8b6356628996f16babd1482c2febd259, {16'd18943, 16'd28976, 16'd44546, 16'd35571, 16'd52605, 16'd4734, 16'd23774, 16'd45175, 16'd57413, 16'd37715, 16'd2388, 16'd53575, 16'd34922, 16'd32365, 16'd30204, 16'd19911, 16'd6150, 16'd32235, 16'd14381, 16'd19003, 16'd50730, 16'd50662, 16'd5201, 16'd16510, 16'd37955, 16'd65080});
	test_expansion(128'he5df60c9a699a89a7e598b8d5b924e44, {16'd13597, 16'd11953, 16'd5439, 16'd57368, 16'd16884, 16'd9508, 16'd55538, 16'd57240, 16'd62626, 16'd16606, 16'd1976, 16'd41135, 16'd3802, 16'd50843, 16'd41143, 16'd6381, 16'd46295, 16'd52888, 16'd36587, 16'd35763, 16'd28753, 16'd33667, 16'd42189, 16'd12690, 16'd3459, 16'd16365});
	test_expansion(128'hda90f927baa7e7bf0323275efad20454, {16'd5489, 16'd18261, 16'd23338, 16'd43548, 16'd3760, 16'd53980, 16'd3873, 16'd2547, 16'd30770, 16'd32506, 16'd30519, 16'd40818, 16'd53444, 16'd25658, 16'd25472, 16'd47036, 16'd13600, 16'd40438, 16'd10744, 16'd46028, 16'd43566, 16'd52419, 16'd64793, 16'd2887, 16'd10995, 16'd45890});
	test_expansion(128'ha38440e700cbb73e5151ed2de8ed8287, {16'd27860, 16'd42689, 16'd13428, 16'd48487, 16'd20432, 16'd49154, 16'd3876, 16'd46810, 16'd2267, 16'd59346, 16'd15518, 16'd21445, 16'd23744, 16'd63304, 16'd3791, 16'd40572, 16'd35619, 16'd54309, 16'd52293, 16'd53793, 16'd15998, 16'd44539, 16'd9181, 16'd5525, 16'd43941, 16'd59251});
	test_expansion(128'ha79ad828cd2594a6c3c28f4fc720ae04, {16'd26439, 16'd27219, 16'd43841, 16'd36712, 16'd32713, 16'd36928, 16'd48144, 16'd2132, 16'd65416, 16'd9347, 16'd17055, 16'd41296, 16'd32696, 16'd13787, 16'd43186, 16'd23995, 16'd50102, 16'd16791, 16'd53562, 16'd55903, 16'd173, 16'd58695, 16'd39508, 16'd2991, 16'd11039, 16'd56247});
	test_expansion(128'h16da3be08deac341921e19a206cc2849, {16'd8605, 16'd61252, 16'd43333, 16'd11554, 16'd44942, 16'd53416, 16'd46935, 16'd53667, 16'd62817, 16'd26, 16'd56411, 16'd62516, 16'd43306, 16'd7148, 16'd28102, 16'd50324, 16'd36485, 16'd41024, 16'd55629, 16'd38202, 16'd62751, 16'd610, 16'd28807, 16'd53615, 16'd43748, 16'd27732});
	test_expansion(128'h79b6aafc2b507af81faff72bdf64558b, {16'd10177, 16'd56879, 16'd24572, 16'd64705, 16'd34371, 16'd33940, 16'd35931, 16'd45227, 16'd33383, 16'd37408, 16'd23849, 16'd64353, 16'd25472, 16'd1868, 16'd62155, 16'd2442, 16'd14402, 16'd17104, 16'd51275, 16'd39133, 16'd43837, 16'd4458, 16'd32900, 16'd31135, 16'd49884, 16'd1261});
	test_expansion(128'hed9f7429b8054b3bf59d69d80b1d95d9, {16'd32995, 16'd30217, 16'd37132, 16'd53313, 16'd40734, 16'd38243, 16'd38898, 16'd30372, 16'd27264, 16'd7333, 16'd56931, 16'd65485, 16'd35713, 16'd45158, 16'd7286, 16'd52593, 16'd53331, 16'd14634, 16'd34679, 16'd36093, 16'd7299, 16'd64369, 16'd2412, 16'd40306, 16'd62915, 16'd16265});
	test_expansion(128'hae7336cbe8e9c16556ea9c8b763602bc, {16'd33150, 16'd35721, 16'd1028, 16'd36803, 16'd48579, 16'd40537, 16'd24607, 16'd25329, 16'd19342, 16'd14274, 16'd14132, 16'd43953, 16'd34101, 16'd65095, 16'd41503, 16'd18676, 16'd9197, 16'd52332, 16'd47824, 16'd13313, 16'd42633, 16'd45568, 16'd7330, 16'd25747, 16'd22923, 16'd51142});
	test_expansion(128'h02e5ee1f6c5b64e80a2780b6ce369c77, {16'd50933, 16'd14666, 16'd9776, 16'd53090, 16'd48991, 16'd2412, 16'd52583, 16'd47309, 16'd39199, 16'd27759, 16'd4133, 16'd41278, 16'd59409, 16'd45970, 16'd3383, 16'd53421, 16'd38210, 16'd5830, 16'd39617, 16'd63147, 16'd41567, 16'd61293, 16'd31818, 16'd38358, 16'd2724, 16'd63585});
	test_expansion(128'h3296e4a11c7238449e0a5d1e5bb41f15, {16'd2002, 16'd49288, 16'd30804, 16'd7086, 16'd55941, 16'd26632, 16'd19611, 16'd2201, 16'd57555, 16'd4959, 16'd53919, 16'd48418, 16'd49583, 16'd21629, 16'd39511, 16'd22191, 16'd28473, 16'd11140, 16'd2444, 16'd14416, 16'd20144, 16'd14487, 16'd62161, 16'd54130, 16'd17319, 16'd28279});
	test_expansion(128'hfd23ed6fe87b666f58d20aa2d9d16fc5, {16'd27232, 16'd47682, 16'd4466, 16'd13355, 16'd58986, 16'd24528, 16'd54467, 16'd58051, 16'd62689, 16'd54199, 16'd63166, 16'd58151, 16'd62709, 16'd2715, 16'd21119, 16'd62655, 16'd64206, 16'd12184, 16'd36323, 16'd21917, 16'd3979, 16'd52563, 16'd30042, 16'd63555, 16'd33523, 16'd48170});
	test_expansion(128'h2deaea9283bb0e912985db8eb182edaa, {16'd2508, 16'd19231, 16'd41487, 16'd36839, 16'd13954, 16'd43201, 16'd63388, 16'd19919, 16'd458, 16'd16344, 16'd58553, 16'd8266, 16'd28883, 16'd63621, 16'd31500, 16'd7380, 16'd58257, 16'd9181, 16'd32175, 16'd44862, 16'd31814, 16'd47341, 16'd41835, 16'd40884, 16'd8374, 16'd23057});
	test_expansion(128'h6b9f176e0f30607d336135d3231f280f, {16'd19788, 16'd50919, 16'd44112, 16'd12410, 16'd47267, 16'd12139, 16'd13306, 16'd56307, 16'd53398, 16'd7487, 16'd47870, 16'd46329, 16'd2664, 16'd37882, 16'd15395, 16'd61280, 16'd11787, 16'd33174, 16'd18854, 16'd46411, 16'd15390, 16'd60516, 16'd24174, 16'd18231, 16'd18997, 16'd35893});
	test_expansion(128'h59d18ade4b14e883492db54c8f86dbf8, {16'd11387, 16'd11204, 16'd16485, 16'd29637, 16'd45831, 16'd1126, 16'd59509, 16'd44497, 16'd49030, 16'd37606, 16'd47343, 16'd12635, 16'd10414, 16'd40809, 16'd65299, 16'd311, 16'd12029, 16'd11762, 16'd54007, 16'd18164, 16'd48300, 16'd38222, 16'd57717, 16'd33427, 16'd17160, 16'd35860});
	test_expansion(128'h061051d0b1867cf967ae2bdb95831fdd, {16'd51092, 16'd53746, 16'd50982, 16'd48957, 16'd40728, 16'd11649, 16'd51421, 16'd46191, 16'd57692, 16'd45044, 16'd64370, 16'd31947, 16'd10175, 16'd35585, 16'd52154, 16'd41191, 16'd15694, 16'd8288, 16'd12428, 16'd46538, 16'd33180, 16'd30264, 16'd58262, 16'd19030, 16'd13507, 16'd12944});
	test_expansion(128'h9207334a2e5e737ab44aeaa0bf7ea4d9, {16'd25290, 16'd56478, 16'd13176, 16'd46638, 16'd63213, 16'd34717, 16'd27522, 16'd63200, 16'd19512, 16'd32143, 16'd43278, 16'd15453, 16'd52463, 16'd23515, 16'd21524, 16'd56022, 16'd43164, 16'd20160, 16'd1537, 16'd60556, 16'd56918, 16'd21320, 16'd48939, 16'd828, 16'd11709, 16'd55686});
	test_expansion(128'hee08e61f779a7f42fb376ac774352354, {16'd56097, 16'd40546, 16'd43512, 16'd62385, 16'd27324, 16'd57951, 16'd46484, 16'd23930, 16'd27204, 16'd35605, 16'd15644, 16'd63515, 16'd62945, 16'd3681, 16'd22836, 16'd500, 16'd23145, 16'd45563, 16'd63554, 16'd36306, 16'd24293, 16'd41252, 16'd47155, 16'd37723, 16'd43781, 16'd53852});
	test_expansion(128'h4aa1d9ea6ac7fe29df83a168440a9561, {16'd31913, 16'd53454, 16'd34486, 16'd25955, 16'd18690, 16'd43137, 16'd2822, 16'd6885, 16'd4558, 16'd42938, 16'd30061, 16'd5199, 16'd57589, 16'd55081, 16'd46158, 16'd16919, 16'd44696, 16'd43427, 16'd30282, 16'd53552, 16'd38410, 16'd3815, 16'd36036, 16'd52669, 16'd63644, 16'd54990});
	test_expansion(128'h3224c2608c94bf825e3600b466cfe24b, {16'd52000, 16'd6822, 16'd47600, 16'd56486, 16'd44219, 16'd23005, 16'd32910, 16'd20631, 16'd4874, 16'd19429, 16'd15910, 16'd17848, 16'd9795, 16'd46255, 16'd1767, 16'd57552, 16'd36262, 16'd47195, 16'd17282, 16'd15649, 16'd32868, 16'd26520, 16'd48414, 16'd34623, 16'd58799, 16'd11004});
	test_expansion(128'hf4db4c545555ceacd62b94e43c741ead, {16'd32627, 16'd52364, 16'd59831, 16'd31120, 16'd683, 16'd50631, 16'd57550, 16'd63980, 16'd57446, 16'd13658, 16'd63131, 16'd10121, 16'd14506, 16'd3773, 16'd55955, 16'd17591, 16'd49973, 16'd42085, 16'd7344, 16'd59988, 16'd54109, 16'd14500, 16'd43668, 16'd18735, 16'd38622, 16'd26949});
	test_expansion(128'ha5074add04d312ab9e7d82998ce59246, {16'd19257, 16'd54201, 16'd45844, 16'd30830, 16'd64322, 16'd10909, 16'd44636, 16'd25159, 16'd58921, 16'd29410, 16'd38842, 16'd63350, 16'd623, 16'd54411, 16'd928, 16'd50279, 16'd33986, 16'd15723, 16'd16874, 16'd19409, 16'd55618, 16'd62351, 16'd11318, 16'd47920, 16'd29080, 16'd61122});
	test_expansion(128'h7ef7ae48aca461c1df3431030c29345d, {16'd1810, 16'd57705, 16'd60142, 16'd18960, 16'd8879, 16'd53203, 16'd31647, 16'd43015, 16'd28920, 16'd19973, 16'd63611, 16'd2242, 16'd28873, 16'd18286, 16'd35186, 16'd19420, 16'd37530, 16'd57788, 16'd31902, 16'd2281, 16'd22205, 16'd6010, 16'd36652, 16'd50952, 16'd37541, 16'd13119});
	test_expansion(128'h9a7aa434c62f1ded7766ac812ba1ef3c, {16'd57506, 16'd10469, 16'd9988, 16'd49921, 16'd40693, 16'd337, 16'd63061, 16'd51156, 16'd48189, 16'd43520, 16'd6372, 16'd14021, 16'd51338, 16'd50152, 16'd43837, 16'd26791, 16'd40497, 16'd49689, 16'd30203, 16'd3659, 16'd13246, 16'd23206, 16'd52622, 16'd47582, 16'd58290, 16'd16568});
	test_expansion(128'h03b38a92cfdbef3620d0a7c2cd64539a, {16'd41614, 16'd15191, 16'd39825, 16'd24886, 16'd60460, 16'd18101, 16'd23955, 16'd12246, 16'd22142, 16'd9965, 16'd47037, 16'd25840, 16'd45881, 16'd16387, 16'd16238, 16'd51849, 16'd54470, 16'd14751, 16'd35597, 16'd60744, 16'd15742, 16'd686, 16'd64823, 16'd40609, 16'd55547, 16'd48009});
	test_expansion(128'h67ab87d7b84ddc0e2e2dfa96eaf5c0f1, {16'd281, 16'd52067, 16'd38447, 16'd52577, 16'd44462, 16'd22495, 16'd3175, 16'd55212, 16'd28473, 16'd59836, 16'd15132, 16'd7278, 16'd37541, 16'd63732, 16'd15365, 16'd56007, 16'd16732, 16'd61467, 16'd48826, 16'd14688, 16'd56484, 16'd46067, 16'd4629, 16'd56420, 16'd50727, 16'd4014});
	test_expansion(128'h2713d2071031a1f083bdf8570dc1c4ed, {16'd1176, 16'd6781, 16'd22125, 16'd51490, 16'd22970, 16'd29289, 16'd45546, 16'd47350, 16'd61040, 16'd11823, 16'd56271, 16'd22776, 16'd42281, 16'd25701, 16'd48583, 16'd3618, 16'd15023, 16'd17033, 16'd1098, 16'd53569, 16'd1149, 16'd50511, 16'd60746, 16'd5930, 16'd23754, 16'd61663});
	test_expansion(128'h15aea783fddbc62ac7c2e1a49b309e1c, {16'd17801, 16'd16131, 16'd38514, 16'd9932, 16'd63009, 16'd28391, 16'd54410, 16'd53742, 16'd19509, 16'd4374, 16'd48189, 16'd37263, 16'd18914, 16'd65039, 16'd16161, 16'd51378, 16'd35664, 16'd49312, 16'd41732, 16'd16677, 16'd40023, 16'd57944, 16'd37723, 16'd22965, 16'd29771, 16'd60547});
	test_expansion(128'h7e805ee45a5d706afab025419b26511c, {16'd61843, 16'd37554, 16'd10101, 16'd24652, 16'd49179, 16'd53222, 16'd14764, 16'd56350, 16'd18925, 16'd16841, 16'd60206, 16'd34670, 16'd14993, 16'd10349, 16'd53352, 16'd61801, 16'd43861, 16'd59397, 16'd31271, 16'd53137, 16'd1156, 16'd44141, 16'd53819, 16'd28390, 16'd8612, 16'd15248});
	test_expansion(128'hf49273d8a397c91b4afcd7b2c863fabd, {16'd59758, 16'd1702, 16'd34504, 16'd50873, 16'd23799, 16'd52881, 16'd14039, 16'd44595, 16'd18802, 16'd48841, 16'd43804, 16'd49222, 16'd41513, 16'd8690, 16'd30902, 16'd61091, 16'd15717, 16'd12205, 16'd56133, 16'd44996, 16'd49657, 16'd18850, 16'd38151, 16'd57112, 16'd10839, 16'd61944});
	test_expansion(128'hf473a2310e5a1096b884b6eb1106c233, {16'd63245, 16'd21000, 16'd5231, 16'd1455, 16'd55532, 16'd26996, 16'd28155, 16'd23333, 16'd57412, 16'd29415, 16'd63800, 16'd29721, 16'd51810, 16'd33698, 16'd22834, 16'd545, 16'd28480, 16'd5957, 16'd6983, 16'd48529, 16'd5417, 16'd39366, 16'd18721, 16'd40214, 16'd48017, 16'd64909});
	test_expansion(128'h14d7da34b06712d2110e1b6963ab422b, {16'd358, 16'd14874, 16'd7135, 16'd34182, 16'd32555, 16'd57930, 16'd12540, 16'd23072, 16'd57807, 16'd7759, 16'd61922, 16'd42340, 16'd52415, 16'd43990, 16'd51331, 16'd59439, 16'd39257, 16'd48267, 16'd30746, 16'd52989, 16'd2102, 16'd48770, 16'd4123, 16'd10996, 16'd755, 16'd63711});
	test_expansion(128'ha25328e01e02c75fc843844dd95d442e, {16'd38603, 16'd58287, 16'd8678, 16'd59801, 16'd36418, 16'd12717, 16'd58685, 16'd32695, 16'd19944, 16'd64411, 16'd5482, 16'd62000, 16'd57920, 16'd32785, 16'd15330, 16'd2325, 16'd54857, 16'd61702, 16'd16599, 16'd3557, 16'd53267, 16'd6750, 16'd42118, 16'd42476, 16'd30311, 16'd38627});
	test_expansion(128'h1cfd87c1e037a5826fa6ed128a0661f1, {16'd43247, 16'd18303, 16'd22262, 16'd16009, 16'd49834, 16'd59443, 16'd9431, 16'd19159, 16'd32050, 16'd31813, 16'd12003, 16'd1562, 16'd39940, 16'd62387, 16'd44355, 16'd31416, 16'd13891, 16'd62443, 16'd31893, 16'd38322, 16'd23141, 16'd7642, 16'd51923, 16'd12051, 16'd46743, 16'd2438});
	test_expansion(128'ha71cff091054f07cc9538b0274c358ef, {16'd37891, 16'd48184, 16'd2775, 16'd63110, 16'd23325, 16'd55627, 16'd18273, 16'd42265, 16'd8415, 16'd59656, 16'd28179, 16'd31786, 16'd18119, 16'd16323, 16'd15366, 16'd14147, 16'd24274, 16'd11633, 16'd8291, 16'd48602, 16'd54019, 16'd10519, 16'd8444, 16'd61629, 16'd60501, 16'd64799});
	test_expansion(128'h3ba4ae6d2d6bea8201971d6f9b3b1b61, {16'd41934, 16'd34115, 16'd26614, 16'd9656, 16'd30095, 16'd51969, 16'd8561, 16'd58210, 16'd47953, 16'd1303, 16'd21381, 16'd41153, 16'd48101, 16'd61149, 16'd18264, 16'd19278, 16'd4050, 16'd42897, 16'd17868, 16'd3132, 16'd3419, 16'd45547, 16'd2584, 16'd17486, 16'd59817, 16'd15339});
	test_expansion(128'h1d2cfd73793b0e606b25e6d979c52e32, {16'd5734, 16'd32996, 16'd54968, 16'd23580, 16'd33119, 16'd64629, 16'd26191, 16'd17679, 16'd43651, 16'd15348, 16'd31118, 16'd51773, 16'd27780, 16'd985, 16'd55841, 16'd27804, 16'd22544, 16'd54081, 16'd59137, 16'd43981, 16'd57255, 16'd61660, 16'd7242, 16'd35796, 16'd14975, 16'd7268});
	test_expansion(128'he4fd383a2095a4e951d04947edb3aa63, {16'd25933, 16'd4090, 16'd14054, 16'd58070, 16'd21067, 16'd63769, 16'd26681, 16'd39274, 16'd39374, 16'd10035, 16'd48428, 16'd45765, 16'd30321, 16'd10111, 16'd53495, 16'd46497, 16'd53311, 16'd3885, 16'd23486, 16'd40668, 16'd39837, 16'd57125, 16'd65343, 16'd26426, 16'd25422, 16'd19039});
	test_expansion(128'h717f6bbb77fe9ba0a61bb9ed4b466e82, {16'd31389, 16'd34197, 16'd31591, 16'd47556, 16'd44056, 16'd44842, 16'd58442, 16'd42928, 16'd27383, 16'd10527, 16'd18717, 16'd15362, 16'd29137, 16'd38937, 16'd31468, 16'd21284, 16'd9772, 16'd47506, 16'd15164, 16'd40606, 16'd10994, 16'd32759, 16'd36291, 16'd8699, 16'd61168, 16'd43253});
	test_expansion(128'hf8adb7f19e9c1e70a9026ceee26c5b5f, {16'd28990, 16'd59605, 16'd29340, 16'd28903, 16'd8580, 16'd57684, 16'd31044, 16'd30978, 16'd49582, 16'd20366, 16'd60282, 16'd6210, 16'd31061, 16'd53435, 16'd14948, 16'd50029, 16'd19351, 16'd55656, 16'd28588, 16'd35414, 16'd47105, 16'd51751, 16'd28278, 16'd18184, 16'd45179, 16'd8682});
	test_expansion(128'h99f1f26639058b32a8cd6267e14b4f53, {16'd281, 16'd25869, 16'd20309, 16'd34196, 16'd35496, 16'd24155, 16'd41084, 16'd18576, 16'd25772, 16'd44397, 16'd20573, 16'd46264, 16'd4017, 16'd18888, 16'd50375, 16'd56230, 16'd26137, 16'd61778, 16'd58448, 16'd27252, 16'd14763, 16'd6059, 16'd29233, 16'd51494, 16'd1935, 16'd36073});
	test_expansion(128'h2639d514d14588278fa0c09c0ef23c0a, {16'd60151, 16'd22925, 16'd27219, 16'd24356, 16'd7595, 16'd33254, 16'd60741, 16'd52057, 16'd37226, 16'd36824, 16'd44460, 16'd57997, 16'd783, 16'd5664, 16'd41363, 16'd35936, 16'd56887, 16'd29598, 16'd10134, 16'd2094, 16'd28987, 16'd53658, 16'd39953, 16'd6967, 16'd43671, 16'd21257});
	test_expansion(128'hed0201b56af68bb2522981ac27222c99, {16'd12721, 16'd38502, 16'd21980, 16'd5963, 16'd32754, 16'd50540, 16'd50688, 16'd25463, 16'd36323, 16'd38124, 16'd35967, 16'd33317, 16'd3926, 16'd34991, 16'd19154, 16'd4495, 16'd51208, 16'd7441, 16'd39995, 16'd38826, 16'd15243, 16'd15228, 16'd16196, 16'd29943, 16'd49995, 16'd43727});
	test_expansion(128'h2c36ccfe70ea5e1071842e6ad85124df, {16'd10834, 16'd50270, 16'd46456, 16'd38710, 16'd20731, 16'd2324, 16'd64265, 16'd17342, 16'd47093, 16'd7874, 16'd17170, 16'd60933, 16'd53063, 16'd21044, 16'd11433, 16'd58682, 16'd31232, 16'd63996, 16'd35024, 16'd38643, 16'd63264, 16'd53526, 16'd31868, 16'd13650, 16'd38446, 16'd38058});
	test_expansion(128'h3ff0c25041bc4ae62edfed7f6f956832, {16'd37147, 16'd22625, 16'd56795, 16'd57371, 16'd62793, 16'd2421, 16'd16644, 16'd9539, 16'd57549, 16'd46975, 16'd32857, 16'd21807, 16'd15689, 16'd64039, 16'd38196, 16'd37378, 16'd47289, 16'd29723, 16'd65503, 16'd14500, 16'd1366, 16'd56216, 16'd42371, 16'd26260, 16'd36869, 16'd15395});
	test_expansion(128'h980dca81720d82140fd3d3a927fc1786, {16'd41969, 16'd51695, 16'd29063, 16'd42820, 16'd61275, 16'd5387, 16'd44231, 16'd54995, 16'd32191, 16'd55126, 16'd14672, 16'd28349, 16'd29409, 16'd24884, 16'd2228, 16'd32402, 16'd55749, 16'd64582, 16'd30742, 16'd43991, 16'd32748, 16'd25101, 16'd27240, 16'd59629, 16'd1283, 16'd41401});
	test_expansion(128'ha5b5b9829127881f04595ec5b78b1ea4, {16'd8743, 16'd51582, 16'd46549, 16'd61553, 16'd13452, 16'd10395, 16'd49962, 16'd64766, 16'd32516, 16'd25775, 16'd9602, 16'd42216, 16'd59793, 16'd31190, 16'd55680, 16'd24541, 16'd28484, 16'd15103, 16'd27921, 16'd51962, 16'd37892, 16'd45919, 16'd44232, 16'd32988, 16'd5928, 16'd10765});
	test_expansion(128'hfb49211d0131e3e523c39e26c0cf5f23, {16'd39077, 16'd19279, 16'd46413, 16'd45684, 16'd24862, 16'd15040, 16'd28884, 16'd24912, 16'd35227, 16'd21539, 16'd26923, 16'd19579, 16'd21826, 16'd42782, 16'd8076, 16'd62545, 16'd29176, 16'd55699, 16'd57044, 16'd35607, 16'd63084, 16'd59757, 16'd13384, 16'd29708, 16'd53207, 16'd14034});
	test_expansion(128'hc376a8438cbb278edbd5f20b27cf8cb9, {16'd2348, 16'd37480, 16'd52093, 16'd13878, 16'd46638, 16'd9086, 16'd9675, 16'd59598, 16'd51496, 16'd20697, 16'd61044, 16'd29470, 16'd42229, 16'd24562, 16'd30374, 16'd22607, 16'd1716, 16'd5939, 16'd46248, 16'd23080, 16'd46457, 16'd16012, 16'd19854, 16'd33534, 16'd62764, 16'd50974});
	test_expansion(128'h79b8d8d1ef01f831bf980a87caa5dc7f, {16'd10814, 16'd25296, 16'd60763, 16'd5327, 16'd44665, 16'd7329, 16'd36482, 16'd62729, 16'd55053, 16'd57498, 16'd10689, 16'd45548, 16'd7703, 16'd63789, 16'd55330, 16'd25297, 16'd58466, 16'd58443, 16'd41238, 16'd47525, 16'd8856, 16'd63293, 16'd18047, 16'd32488, 16'd43616, 16'd9532});
	test_expansion(128'h3680ea03bfa6466c59046982a0bb1944, {16'd48098, 16'd26340, 16'd16610, 16'd13775, 16'd171, 16'd55794, 16'd36885, 16'd11942, 16'd3245, 16'd31777, 16'd18981, 16'd25201, 16'd51372, 16'd33707, 16'd44900, 16'd1916, 16'd9048, 16'd628, 16'd1752, 16'd3373, 16'd38576, 16'd26635, 16'd14424, 16'd43046, 16'd50043, 16'd31431});
	test_expansion(128'hbf90591e83fffc004f88ec6bba1ce48a, {16'd9270, 16'd42869, 16'd3641, 16'd58463, 16'd9412, 16'd13473, 16'd42383, 16'd38957, 16'd1784, 16'd44489, 16'd38698, 16'd34069, 16'd46338, 16'd63147, 16'd8998, 16'd20548, 16'd8694, 16'd21140, 16'd1710, 16'd27621, 16'd23762, 16'd63374, 16'd40225, 16'd31758, 16'd37808, 16'd61307});
	test_expansion(128'hbe55249f6595aab6f779af39f25349fe, {16'd63627, 16'd53650, 16'd7759, 16'd37337, 16'd31837, 16'd27651, 16'd17372, 16'd32333, 16'd30059, 16'd41280, 16'd17568, 16'd18599, 16'd49815, 16'd3382, 16'd49817, 16'd2534, 16'd55150, 16'd9036, 16'd55435, 16'd42848, 16'd35020, 16'd18408, 16'd52501, 16'd18876, 16'd1489, 16'd36102});
	test_expansion(128'h80a02c26027303b3539b570309dd027b, {16'd15252, 16'd9574, 16'd9583, 16'd45642, 16'd51825, 16'd22698, 16'd29545, 16'd52905, 16'd25161, 16'd31272, 16'd35830, 16'd64000, 16'd25920, 16'd30782, 16'd56024, 16'd64713, 16'd26166, 16'd46355, 16'd38054, 16'd1977, 16'd3260, 16'd13881, 16'd14773, 16'd39421, 16'd7797, 16'd23178});
	test_expansion(128'h26c991f4395c063ca806c81a3089cf31, {16'd30210, 16'd46428, 16'd57364, 16'd29613, 16'd42875, 16'd37310, 16'd39619, 16'd61854, 16'd20904, 16'd40372, 16'd56424, 16'd55063, 16'd45060, 16'd21447, 16'd37457, 16'd62503, 16'd59231, 16'd16041, 16'd64479, 16'd56348, 16'd3589, 16'd40765, 16'd22375, 16'd18110, 16'd4086, 16'd33748});
	test_expansion(128'h82acd3d1d8fb8d88e03a495c4be5e454, {16'd40853, 16'd27947, 16'd41203, 16'd11530, 16'd13026, 16'd11050, 16'd23703, 16'd59940, 16'd9502, 16'd2525, 16'd46201, 16'd39712, 16'd38357, 16'd31456, 16'd46461, 16'd31029, 16'd56743, 16'd41457, 16'd14722, 16'd26041, 16'd11263, 16'd44381, 16'd49836, 16'd42003, 16'd2259, 16'd48199});
	test_expansion(128'hd9aa7fa973167a8c9d171bd9480fdee8, {16'd33909, 16'd24554, 16'd47793, 16'd40930, 16'd32583, 16'd13597, 16'd63241, 16'd20251, 16'd40041, 16'd60897, 16'd13286, 16'd1244, 16'd23593, 16'd20575, 16'd18823, 16'd37730, 16'd18474, 16'd36771, 16'd63093, 16'd60085, 16'd62487, 16'd32348, 16'd40537, 16'd42474, 16'd24902, 16'd18083});
	test_expansion(128'h763fc558a2744f2f7ff9ef1935732099, {16'd38879, 16'd43303, 16'd14285, 16'd57920, 16'd18745, 16'd20286, 16'd38853, 16'd64063, 16'd23310, 16'd47670, 16'd12307, 16'd46277, 16'd36630, 16'd64806, 16'd39919, 16'd57683, 16'd46345, 16'd42888, 16'd55712, 16'd54300, 16'd14457, 16'd52244, 16'd40377, 16'd41915, 16'd3580, 16'd927});
	test_expansion(128'h8fbf71d91f90755d96011a70b7686933, {16'd46438, 16'd12396, 16'd1655, 16'd12936, 16'd35873, 16'd57316, 16'd539, 16'd8307, 16'd17651, 16'd31226, 16'd20330, 16'd63110, 16'd39474, 16'd48880, 16'd47443, 16'd31169, 16'd60512, 16'd45206, 16'd33900, 16'd58867, 16'd49248, 16'd37604, 16'd50433, 16'd27766, 16'd65122, 16'd35298});
	test_expansion(128'h9c2d64f15a4afd33cf7e2a1e6acf4acc, {16'd63912, 16'd53870, 16'd51289, 16'd20367, 16'd25802, 16'd53028, 16'd63497, 16'd54662, 16'd9404, 16'd65114, 16'd55513, 16'd755, 16'd7960, 16'd51596, 16'd41943, 16'd18062, 16'd1031, 16'd38738, 16'd2126, 16'd17741, 16'd39072, 16'd54546, 16'd53196, 16'd1277, 16'd13925, 16'd62433});
	test_expansion(128'h9a82db20d08ce34c7605f69f9a4528b1, {16'd42929, 16'd8478, 16'd17516, 16'd9547, 16'd32918, 16'd58956, 16'd64821, 16'd22935, 16'd30281, 16'd24625, 16'd27914, 16'd46150, 16'd59433, 16'd38506, 16'd4569, 16'd50549, 16'd49161, 16'd46039, 16'd13599, 16'd32285, 16'd47207, 16'd38788, 16'd38576, 16'd31374, 16'd24794, 16'd30367});
	test_expansion(128'h2bb249752296719b0fd42fdb9e063969, {16'd6962, 16'd64942, 16'd45534, 16'd16245, 16'd42593, 16'd57319, 16'd18479, 16'd59595, 16'd29353, 16'd3014, 16'd52071, 16'd33529, 16'd5621, 16'd63498, 16'd52299, 16'd62974, 16'd17962, 16'd30343, 16'd52459, 16'd27083, 16'd59566, 16'd47802, 16'd52385, 16'd26916, 16'd51650, 16'd62776});
	test_expansion(128'h39849bb843dd732db182cbe341dd2abb, {16'd46131, 16'd24360, 16'd59838, 16'd46080, 16'd56614, 16'd15688, 16'd61600, 16'd55494, 16'd61634, 16'd51777, 16'd10608, 16'd32802, 16'd3090, 16'd58887, 16'd8126, 16'd51176, 16'd2604, 16'd12809, 16'd45298, 16'd9906, 16'd44199, 16'd54279, 16'd52914, 16'd15495, 16'd52406, 16'd9926});
	test_expansion(128'h5a74da6d66e4d3cb5ee3848f45309e14, {16'd47728, 16'd19073, 16'd28169, 16'd46471, 16'd416, 16'd16161, 16'd34388, 16'd59472, 16'd16139, 16'd1044, 16'd4895, 16'd35530, 16'd12652, 16'd6705, 16'd1868, 16'd39993, 16'd35785, 16'd12084, 16'd20978, 16'd40270, 16'd40376, 16'd50, 16'd20, 16'd1335, 16'd263, 16'd12575});
	test_expansion(128'hd7357c1a14c1561d3bce89b177f35448, {16'd47963, 16'd40623, 16'd24267, 16'd14383, 16'd61327, 16'd27609, 16'd49642, 16'd61562, 16'd52835, 16'd32711, 16'd8446, 16'd2839, 16'd12122, 16'd54112, 16'd17651, 16'd47362, 16'd7083, 16'd38419, 16'd35622, 16'd35109, 16'd63146, 16'd51572, 16'd8952, 16'd44037, 16'd17209, 16'd23960});
	test_expansion(128'h295aa85c8afe5fe43bef6a0c963efdd0, {16'd34394, 16'd14046, 16'd1145, 16'd39094, 16'd16028, 16'd27788, 16'd4563, 16'd49223, 16'd5060, 16'd19495, 16'd24372, 16'd35272, 16'd44066, 16'd53483, 16'd22361, 16'd53941, 16'd37007, 16'd15595, 16'd48350, 16'd43855, 16'd53280, 16'd21809, 16'd39284, 16'd712, 16'd60103, 16'd5539});
	test_expansion(128'h2c93d15cfec8e59c4935e7c4096d7df0, {16'd6265, 16'd57234, 16'd356, 16'd59156, 16'd34238, 16'd63365, 16'd33452, 16'd40555, 16'd10709, 16'd11387, 16'd60715, 16'd34788, 16'd6279, 16'd5902, 16'd23550, 16'd1542, 16'd64463, 16'd26966, 16'd21586, 16'd30388, 16'd42139, 16'd58853, 16'd56145, 16'd58493, 16'd11064, 16'd40073});
	test_expansion(128'h1b436790e24c90e100ae5d2eab9a928c, {16'd18054, 16'd35120, 16'd40962, 16'd22246, 16'd53304, 16'd2896, 16'd45543, 16'd8938, 16'd58977, 16'd35687, 16'd65290, 16'd6789, 16'd42990, 16'd8721, 16'd10007, 16'd6619, 16'd51957, 16'd31883, 16'd28031, 16'd24488, 16'd62316, 16'd41390, 16'd27594, 16'd30787, 16'd27435, 16'd40296});
	test_expansion(128'h2418c26e8b3f144a122cdb11ef7f370d, {16'd39004, 16'd17674, 16'd20074, 16'd43371, 16'd64201, 16'd1009, 16'd27456, 16'd45563, 16'd57768, 16'd34980, 16'd39955, 16'd25189, 16'd3858, 16'd2876, 16'd58444, 16'd43701, 16'd17966, 16'd61854, 16'd18375, 16'd18950, 16'd17220, 16'd655, 16'd8632, 16'd45584, 16'd48270, 16'd7598});
	test_expansion(128'h14a69cedd5f6b0ae937b032b06cab822, {16'd65417, 16'd51811, 16'd12061, 16'd48072, 16'd28256, 16'd12346, 16'd34911, 16'd57377, 16'd7288, 16'd12137, 16'd24367, 16'd63419, 16'd3406, 16'd303, 16'd54941, 16'd12588, 16'd62968, 16'd38798, 16'd14916, 16'd64790, 16'd50349, 16'd49991, 16'd46026, 16'd47284, 16'd10706, 16'd24191});
	test_expansion(128'h49aca9aca662add19a2cab65e53ec36f, {16'd14293, 16'd2581, 16'd37724, 16'd12121, 16'd24780, 16'd26902, 16'd58009, 16'd5247, 16'd24244, 16'd55929, 16'd15258, 16'd41882, 16'd60792, 16'd61691, 16'd33852, 16'd7791, 16'd4854, 16'd23678, 16'd11566, 16'd6576, 16'd31764, 16'd40763, 16'd55710, 16'd19665, 16'd45750, 16'd14689});
	test_expansion(128'h89c3e366739914832ca51ea782efcf35, {16'd58393, 16'd32499, 16'd23920, 16'd26593, 16'd10860, 16'd60044, 16'd40853, 16'd40837, 16'd7956, 16'd18908, 16'd32329, 16'd53977, 16'd32380, 16'd49609, 16'd21471, 16'd30874, 16'd60657, 16'd45619, 16'd42036, 16'd22821, 16'd18649, 16'd35557, 16'd21624, 16'd15858, 16'd49111, 16'd44655});
	test_expansion(128'h9067ea6ba6fc61a1e5f63f16571899d7, {16'd42424, 16'd32468, 16'd46702, 16'd3926, 16'd16618, 16'd45162, 16'd17338, 16'd16079, 16'd40474, 16'd20339, 16'd6981, 16'd61420, 16'd48236, 16'd3146, 16'd45372, 16'd27978, 16'd43680, 16'd3165, 16'd24273, 16'd13929, 16'd27163, 16'd14269, 16'd47287, 16'd21279, 16'd61447, 16'd46741});
	test_expansion(128'hf64055f1e6e0241a843c23a872b9e877, {16'd27520, 16'd31893, 16'd50181, 16'd65030, 16'd1086, 16'd54451, 16'd52399, 16'd21440, 16'd52251, 16'd4720, 16'd44495, 16'd59012, 16'd55974, 16'd42830, 16'd36087, 16'd34484, 16'd48576, 16'd46146, 16'd42339, 16'd52177, 16'd20128, 16'd13035, 16'd23729, 16'd21402, 16'd50405, 16'd28895});
	test_expansion(128'ha347eb0d65bae98fd07b1e2deff1a658, {16'd32441, 16'd40418, 16'd38891, 16'd54546, 16'd3979, 16'd19604, 16'd53911, 16'd14758, 16'd24234, 16'd2615, 16'd20241, 16'd45959, 16'd56933, 16'd53677, 16'd27353, 16'd14631, 16'd10726, 16'd4439, 16'd2947, 16'd8604, 16'd32953, 16'd38488, 16'd58428, 16'd62445, 16'd49860, 16'd52815});
	test_expansion(128'ha360c7f183aa97773b5f6b582f515a65, {16'd21349, 16'd61231, 16'd64134, 16'd61547, 16'd55036, 16'd32964, 16'd21906, 16'd43904, 16'd37327, 16'd21574, 16'd3899, 16'd38313, 16'd2779, 16'd52593, 16'd3218, 16'd30362, 16'd22858, 16'd14191, 16'd20315, 16'd55137, 16'd25210, 16'd45530, 16'd25786, 16'd24002, 16'd60643, 16'd56666});
	test_expansion(128'h1d165d20dc2530e2c82852f900f29a0a, {16'd25747, 16'd4488, 16'd40612, 16'd37780, 16'd50113, 16'd43512, 16'd27181, 16'd1802, 16'd22343, 16'd13288, 16'd4559, 16'd36316, 16'd38437, 16'd49645, 16'd28695, 16'd18794, 16'd36934, 16'd49439, 16'd28292, 16'd7977, 16'd64814, 16'd54415, 16'd45879, 16'd18912, 16'd52848, 16'd59352});
	test_expansion(128'hdae200664b708772552a735e98a6e844, {16'd27439, 16'd43877, 16'd11649, 16'd56853, 16'd43742, 16'd22581, 16'd45440, 16'd63866, 16'd14970, 16'd14940, 16'd19630, 16'd27690, 16'd1299, 16'd26549, 16'd7842, 16'd47292, 16'd49234, 16'd7961, 16'd49942, 16'd62274, 16'd53389, 16'd45548, 16'd43185, 16'd20434, 16'd43770, 16'd5606});
	test_expansion(128'ha3f654a364a4ec266dcc1c780e1b7f79, {16'd11397, 16'd11607, 16'd8806, 16'd31994, 16'd59230, 16'd48108, 16'd20007, 16'd15571, 16'd44985, 16'd10067, 16'd32379, 16'd44165, 16'd38467, 16'd54528, 16'd21156, 16'd59708, 16'd28985, 16'd15882, 16'd32340, 16'd35870, 16'd57823, 16'd24270, 16'd32952, 16'd25871, 16'd3670, 16'd17863});
	test_expansion(128'ha6692f2806eb8427f9cc6672674ce2ab, {16'd65060, 16'd36235, 16'd60757, 16'd47128, 16'd16885, 16'd36761, 16'd29077, 16'd10206, 16'd56485, 16'd59361, 16'd60312, 16'd39537, 16'd23878, 16'd8494, 16'd12982, 16'd45692, 16'd28156, 16'd11665, 16'd352, 16'd6435, 16'd10036, 16'd20121, 16'd36311, 16'd21529, 16'd34913, 16'd42594});
	test_expansion(128'h88b123c9c59f6cc149b2175822999f75, {16'd41786, 16'd55479, 16'd29905, 16'd25251, 16'd36012, 16'd51902, 16'd17139, 16'd48015, 16'd13360, 16'd499, 16'd22284, 16'd45086, 16'd16304, 16'd44778, 16'd1092, 16'd54477, 16'd23130, 16'd29504, 16'd30713, 16'd58918, 16'd60959, 16'd54227, 16'd38273, 16'd61365, 16'd31098, 16'd47221});
	test_expansion(128'h4a994d16df29341134edd406ff64ece9, {16'd4623, 16'd32186, 16'd23889, 16'd10398, 16'd14645, 16'd9838, 16'd9351, 16'd16116, 16'd45642, 16'd340, 16'd60178, 16'd63374, 16'd23873, 16'd58687, 16'd57856, 16'd30992, 16'd3032, 16'd19199, 16'd21399, 16'd8637, 16'd29712, 16'd22570, 16'd3822, 16'd9318, 16'd7011, 16'd40628});
	test_expansion(128'h37dfdc4ecf747738ce22a4643490fbd3, {16'd26963, 16'd40209, 16'd59485, 16'd47926, 16'd14053, 16'd51956, 16'd53472, 16'd13935, 16'd37069, 16'd21937, 16'd59403, 16'd39440, 16'd10759, 16'd25890, 16'd36789, 16'd28637, 16'd47211, 16'd12004, 16'd55607, 16'd20707, 16'd56480, 16'd6893, 16'd47817, 16'd50685, 16'd39353, 16'd9349});
	test_expansion(128'h9e7068b052383ffb1210768d8bc9ac07, {16'd59658, 16'd713, 16'd42900, 16'd25476, 16'd61780, 16'd109, 16'd27505, 16'd23852, 16'd30278, 16'd22906, 16'd45384, 16'd10738, 16'd26325, 16'd6680, 16'd17010, 16'd21516, 16'd6063, 16'd10443, 16'd40517, 16'd53792, 16'd3705, 16'd28348, 16'd15155, 16'd55984, 16'd2702, 16'd17580});
	test_expansion(128'h348b79c9e8dd90ea64a3d8cc0bb9110e, {16'd2497, 16'd48582, 16'd32186, 16'd42379, 16'd21118, 16'd14724, 16'd13945, 16'd55560, 16'd48466, 16'd11923, 16'd51512, 16'd51477, 16'd51332, 16'd43598, 16'd38159, 16'd47171, 16'd575, 16'd4482, 16'd15520, 16'd14011, 16'd18922, 16'd41868, 16'd14252, 16'd14819, 16'd50843, 16'd10757});
	test_expansion(128'hd041174155797b306349b094273f5391, {16'd32812, 16'd51512, 16'd52346, 16'd60280, 16'd6599, 16'd9927, 16'd63707, 16'd65434, 16'd32895, 16'd26520, 16'd60965, 16'd19761, 16'd18797, 16'd16588, 16'd42007, 16'd63168, 16'd46992, 16'd48041, 16'd21061, 16'd43415, 16'd26269, 16'd53162, 16'd49845, 16'd34612, 16'd8133, 16'd52058});
	test_expansion(128'hd9c19b279efda3f4a1ff1f85d937f379, {16'd52115, 16'd16719, 16'd63167, 16'd6671, 16'd13732, 16'd15095, 16'd1750, 16'd4279, 16'd3963, 16'd17726, 16'd37606, 16'd18371, 16'd57817, 16'd64000, 16'd64163, 16'd45316, 16'd50460, 16'd15931, 16'd14048, 16'd31569, 16'd28962, 16'd61165, 16'd4038, 16'd1579, 16'd49052, 16'd53510});
	test_expansion(128'h0c0ff3d4a72e7c655f66be5ae902ed07, {16'd47455, 16'd35253, 16'd27708, 16'd54465, 16'd57989, 16'd13721, 16'd4324, 16'd12221, 16'd23290, 16'd20269, 16'd23407, 16'd52998, 16'd27704, 16'd34703, 16'd30056, 16'd64441, 16'd63809, 16'd48387, 16'd60613, 16'd30456, 16'd63309, 16'd42557, 16'd54979, 16'd3684, 16'd32978, 16'd54373});
	test_expansion(128'h8a3f0c146a2150f54de8b1abee52a226, {16'd39281, 16'd61528, 16'd60750, 16'd37795, 16'd37547, 16'd49279, 16'd41177, 16'd19638, 16'd61083, 16'd61901, 16'd8203, 16'd2075, 16'd21224, 16'd21461, 16'd38870, 16'd21736, 16'd28589, 16'd45199, 16'd58741, 16'd64569, 16'd64026, 16'd11379, 16'd35022, 16'd45447, 16'd18317, 16'd6581});
	test_expansion(128'h53c80ab0d97c0b71a2cb96adcd01fdd3, {16'd59375, 16'd40617, 16'd7850, 16'd61954, 16'd46733, 16'd18585, 16'd31338, 16'd48414, 16'd24749, 16'd46544, 16'd23750, 16'd61607, 16'd54909, 16'd5354, 16'd62144, 16'd37050, 16'd59805, 16'd8232, 16'd14841, 16'd41882, 16'd23798, 16'd22545, 16'd33099, 16'd65098, 16'd32634, 16'd56329});
	test_expansion(128'h5732f0b048b287a48dba8068a07a9be1, {16'd23695, 16'd19172, 16'd4536, 16'd34417, 16'd26434, 16'd4570, 16'd50700, 16'd49418, 16'd14089, 16'd11497, 16'd50094, 16'd46694, 16'd31684, 16'd44493, 16'd18582, 16'd42296, 16'd64251, 16'd35648, 16'd61529, 16'd28008, 16'd50276, 16'd23561, 16'd59796, 16'd7502, 16'd64305, 16'd3030});
	test_expansion(128'h2821d4189ea82731a0ba29fb0083dea0, {16'd9944, 16'd46032, 16'd59813, 16'd59256, 16'd56276, 16'd43991, 16'd64522, 16'd56125, 16'd46041, 16'd3976, 16'd34803, 16'd22424, 16'd18722, 16'd63414, 16'd42665, 16'd3856, 16'd14369, 16'd25806, 16'd58090, 16'd52006, 16'd30356, 16'd63504, 16'd56621, 16'd56450, 16'd47854, 16'd31754});
	test_expansion(128'h2d3d59f7ed09d4f1e49142640afe6d0f, {16'd9712, 16'd1572, 16'd5998, 16'd34916, 16'd34074, 16'd46165, 16'd33076, 16'd25370, 16'd13847, 16'd35705, 16'd64833, 16'd1586, 16'd50264, 16'd31646, 16'd58139, 16'd19933, 16'd57576, 16'd37361, 16'd14795, 16'd14137, 16'd31165, 16'd59965, 16'd5488, 16'd35545, 16'd35643, 16'd362});
	test_expansion(128'h44af475ea70a9e69a8c4da4ce0e09355, {16'd61472, 16'd31794, 16'd20353, 16'd23092, 16'd1301, 16'd36625, 16'd42825, 16'd54456, 16'd11886, 16'd54811, 16'd38205, 16'd50145, 16'd9619, 16'd3027, 16'd40716, 16'd13021, 16'd51866, 16'd3665, 16'd55388, 16'd23209, 16'd15168, 16'd39530, 16'd21366, 16'd27898, 16'd65357, 16'd10589});
	test_expansion(128'hc29003b881d0ed95c717b8ac9e77266d, {16'd57548, 16'd39304, 16'd63557, 16'd26340, 16'd60709, 16'd60360, 16'd43324, 16'd28019, 16'd45428, 16'd56303, 16'd15999, 16'd62300, 16'd212, 16'd25339, 16'd33661, 16'd23118, 16'd14703, 16'd28317, 16'd23882, 16'd10357, 16'd59723, 16'd17132, 16'd32385, 16'd53834, 16'd39809, 16'd16209});
	test_expansion(128'hf7be184d87b4626af6746e4169c27c8d, {16'd42845, 16'd29930, 16'd1943, 16'd47266, 16'd41159, 16'd22866, 16'd62454, 16'd4704, 16'd24206, 16'd27275, 16'd60045, 16'd61009, 16'd5940, 16'd56398, 16'd25554, 16'd56742, 16'd29660, 16'd32677, 16'd53631, 16'd6102, 16'd9500, 16'd33465, 16'd29658, 16'd16082, 16'd529, 16'd5899});
	test_expansion(128'hbba342f36424e1953335e52df3328548, {16'd58030, 16'd42231, 16'd24775, 16'd7413, 16'd20101, 16'd51055, 16'd14285, 16'd33532, 16'd21797, 16'd32798, 16'd59928, 16'd3200, 16'd47645, 16'd27621, 16'd1019, 16'd63989, 16'd54336, 16'd40980, 16'd31186, 16'd6763, 16'd62989, 16'd62840, 16'd32239, 16'd38596, 16'd27187, 16'd2817});
	test_expansion(128'hff9cdb202cad2e87604d4252ec89d05b, {16'd59547, 16'd34049, 16'd45084, 16'd48685, 16'd42734, 16'd14341, 16'd44892, 16'd57260, 16'd50295, 16'd17803, 16'd43449, 16'd2059, 16'd41024, 16'd38758, 16'd15189, 16'd1093, 16'd15949, 16'd46530, 16'd63809, 16'd17071, 16'd34460, 16'd19965, 16'd12294, 16'd2410, 16'd36892, 16'd6052});
	test_expansion(128'h7629d3c36b549ec4a8973cd3dc0ee1fa, {16'd51941, 16'd40014, 16'd5726, 16'd17707, 16'd23541, 16'd5411, 16'd30824, 16'd57434, 16'd15349, 16'd3981, 16'd21997, 16'd11557, 16'd21341, 16'd16258, 16'd64730, 16'd51307, 16'd38314, 16'd57438, 16'd47821, 16'd34938, 16'd34758, 16'd30352, 16'd64638, 16'd58550, 16'd19294, 16'd2310});
	test_expansion(128'hf1b1459ea9c0177e09b51495360e41ed, {16'd24558, 16'd28139, 16'd61887, 16'd13115, 16'd9306, 16'd1670, 16'd39972, 16'd8722, 16'd46297, 16'd2497, 16'd61990, 16'd3434, 16'd24883, 16'd37906, 16'd43680, 16'd29300, 16'd63965, 16'd56306, 16'd35116, 16'd39488, 16'd28851, 16'd34931, 16'd37706, 16'd46090, 16'd50876, 16'd7867});
	test_expansion(128'h23b2a9cea9282ae30824442a7749f396, {16'd21817, 16'd43688, 16'd4117, 16'd40335, 16'd17908, 16'd10653, 16'd61564, 16'd46859, 16'd50357, 16'd53478, 16'd12076, 16'd19496, 16'd52005, 16'd53194, 16'd27939, 16'd5877, 16'd63789, 16'd50249, 16'd63624, 16'd64315, 16'd47970, 16'd15450, 16'd17345, 16'd53681, 16'd39724, 16'd1944});
	test_expansion(128'h162a692478071e69e6ec580fb6d0609d, {16'd36986, 16'd11042, 16'd60271, 16'd24762, 16'd50567, 16'd3987, 16'd7171, 16'd20704, 16'd13918, 16'd50453, 16'd31412, 16'd14712, 16'd41345, 16'd53578, 16'd23745, 16'd42219, 16'd35102, 16'd52852, 16'd40984, 16'd61075, 16'd4506, 16'd17952, 16'd60336, 16'd65145, 16'd2412, 16'd46487});
	test_expansion(128'h0bb08aec948f3eeca77542ef74ea911f, {16'd9677, 16'd139, 16'd129, 16'd56815, 16'd51628, 16'd7147, 16'd51823, 16'd34342, 16'd43555, 16'd280, 16'd15761, 16'd31945, 16'd42031, 16'd60526, 16'd53718, 16'd29027, 16'd50203, 16'd1307, 16'd61886, 16'd12978, 16'd63957, 16'd17184, 16'd42223, 16'd27231, 16'd28050, 16'd43540});
	test_expansion(128'h648592d8ca60339fb9690d8318743260, {16'd13255, 16'd38121, 16'd61227, 16'd15925, 16'd18895, 16'd26885, 16'd31093, 16'd30496, 16'd45891, 16'd31158, 16'd43818, 16'd3994, 16'd18022, 16'd14243, 16'd43716, 16'd28561, 16'd56490, 16'd52493, 16'd32168, 16'd30090, 16'd35005, 16'd45459, 16'd33529, 16'd43785, 16'd41499, 16'd13303});
	test_expansion(128'h8bb57301314336234e3a6e1527adda8d, {16'd56326, 16'd19738, 16'd57538, 16'd13034, 16'd727, 16'd18604, 16'd65335, 16'd41148, 16'd32460, 16'd62575, 16'd60397, 16'd31033, 16'd5741, 16'd5908, 16'd38945, 16'd37904, 16'd6913, 16'd47966, 16'd63160, 16'd51318, 16'd51530, 16'd23179, 16'd55957, 16'd16484, 16'd40887, 16'd48781});
	test_expansion(128'hb27a6d26e8232ea9a91e3310486a4117, {16'd41110, 16'd22119, 16'd21427, 16'd24586, 16'd34328, 16'd42834, 16'd16503, 16'd13737, 16'd12157, 16'd37839, 16'd14624, 16'd4820, 16'd61616, 16'd62701, 16'd10341, 16'd60526, 16'd28309, 16'd45238, 16'd61660, 16'd33576, 16'd40396, 16'd7665, 16'd37931, 16'd4662, 16'd49145, 16'd33409});
	test_expansion(128'hd35648fecad38f25b7b8620fd7d9a086, {16'd2050, 16'd23965, 16'd14504, 16'd4304, 16'd1648, 16'd44938, 16'd46880, 16'd45991, 16'd46477, 16'd23318, 16'd63902, 16'd35844, 16'd53856, 16'd714, 16'd6155, 16'd61037, 16'd8963, 16'd50400, 16'd9340, 16'd38567, 16'd64764, 16'd34831, 16'd6058, 16'd17621, 16'd56560, 16'd5091});
	test_expansion(128'h8f487e9a4eef787c3956d751e612021d, {16'd43109, 16'd35981, 16'd18244, 16'd19830, 16'd18517, 16'd3779, 16'd11255, 16'd43198, 16'd33373, 16'd21688, 16'd64121, 16'd15099, 16'd4620, 16'd8347, 16'd26529, 16'd59386, 16'd38844, 16'd16493, 16'd27812, 16'd28482, 16'd5265, 16'd23879, 16'd42968, 16'd421, 16'd18112, 16'd17777});
	test_expansion(128'h9b35c137369e2681de8345a77965fb13, {16'd51549, 16'd54212, 16'd24918, 16'd34224, 16'd18062, 16'd9188, 16'd14919, 16'd20918, 16'd34904, 16'd33330, 16'd65243, 16'd26166, 16'd33365, 16'd59528, 16'd65234, 16'd31826, 16'd39803, 16'd43222, 16'd58384, 16'd52776, 16'd3206, 16'd25725, 16'd42361, 16'd54622, 16'd10382, 16'd25875});
	test_expansion(128'h15b373b281d39f528fecfbb9cad33f2c, {16'd8489, 16'd2334, 16'd754, 16'd18028, 16'd39100, 16'd8095, 16'd60213, 16'd30616, 16'd22363, 16'd41096, 16'd61447, 16'd48807, 16'd45825, 16'd56481, 16'd64784, 16'd33781, 16'd49460, 16'd15071, 16'd861, 16'd34861, 16'd28933, 16'd16684, 16'd57994, 16'd65369, 16'd26381, 16'd787});
	test_expansion(128'hff668018a26c8f6fc412700864afc196, {16'd5899, 16'd55085, 16'd8787, 16'd47479, 16'd28578, 16'd42610, 16'd14504, 16'd60635, 16'd14274, 16'd48404, 16'd54001, 16'd37097, 16'd50936, 16'd37712, 16'd30183, 16'd57635, 16'd6012, 16'd54332, 16'd38784, 16'd41100, 16'd47253, 16'd36174, 16'd2601, 16'd12802, 16'd44193, 16'd22117});
	test_expansion(128'ha37991ed605ec0c06411ec7e5033caa4, {16'd8162, 16'd28868, 16'd33657, 16'd49739, 16'd34411, 16'd64846, 16'd33186, 16'd25958, 16'd9196, 16'd9205, 16'd1733, 16'd48259, 16'd3027, 16'd21504, 16'd60535, 16'd14970, 16'd52194, 16'd28572, 16'd852, 16'd25677, 16'd39282, 16'd33813, 16'd58297, 16'd3030, 16'd41434, 16'd22771});
	test_expansion(128'hc5d34f67bedad1b9280bab4fcde53305, {16'd51805, 16'd2504, 16'd46137, 16'd59706, 16'd8589, 16'd53269, 16'd37349, 16'd57538, 16'd27157, 16'd47617, 16'd21883, 16'd64881, 16'd33615, 16'd22449, 16'd22549, 16'd45813, 16'd1848, 16'd23732, 16'd52750, 16'd51918, 16'd26165, 16'd49983, 16'd36467, 16'd14560, 16'd52064, 16'd29270});
	test_expansion(128'h3b5a10284fa6803e789ee60c10f89fe6, {16'd40709, 16'd5338, 16'd54554, 16'd52917, 16'd27818, 16'd52853, 16'd41076, 16'd61937, 16'd34632, 16'd55177, 16'd47843, 16'd10137, 16'd61533, 16'd4169, 16'd54415, 16'd5707, 16'd31122, 16'd61468, 16'd14855, 16'd36846, 16'd43295, 16'd963, 16'd41095, 16'd52482, 16'd29687, 16'd49046});
	test_expansion(128'hbb32af4d4b368e0591a2fdcc4ecb26a5, {16'd23638, 16'd36280, 16'd43882, 16'd5623, 16'd25980, 16'd28531, 16'd58145, 16'd40191, 16'd11608, 16'd57575, 16'd9800, 16'd20481, 16'd61499, 16'd5891, 16'd3184, 16'd33471, 16'd36800, 16'd59076, 16'd31374, 16'd57381, 16'd2948, 16'd34238, 16'd48613, 16'd28062, 16'd35602, 16'd50741});
	test_expansion(128'h6cffeaa2b40b7f1f9376a0623b6be392, {16'd48482, 16'd3973, 16'd22793, 16'd47649, 16'd18017, 16'd36965, 16'd14584, 16'd50768, 16'd39838, 16'd1972, 16'd17790, 16'd42457, 16'd55751, 16'd56653, 16'd16889, 16'd21117, 16'd12618, 16'd55670, 16'd29874, 16'd44405, 16'd37337, 16'd55171, 16'd12849, 16'd45316, 16'd64764, 16'd42097});
	test_expansion(128'he63bfe193aface0d5fc7a84ace30147c, {16'd18161, 16'd4242, 16'd41871, 16'd25399, 16'd45011, 16'd42293, 16'd60833, 16'd14615, 16'd31930, 16'd26319, 16'd15521, 16'd38906, 16'd7763, 16'd7998, 16'd55565, 16'd25614, 16'd39364, 16'd49540, 16'd62261, 16'd50058, 16'd11910, 16'd56184, 16'd51040, 16'd33658, 16'd32289, 16'd53194});
	test_expansion(128'hd4c6a5868b9fb062d3cc832b85ae3923, {16'd22009, 16'd54015, 16'd56235, 16'd19396, 16'd38802, 16'd4569, 16'd31322, 16'd50556, 16'd9929, 16'd29585, 16'd27901, 16'd62417, 16'd17361, 16'd23310, 16'd39121, 16'd37880, 16'd4134, 16'd28204, 16'd15310, 16'd18545, 16'd41633, 16'd49071, 16'd57779, 16'd60566, 16'd47103, 16'd55455});
	test_expansion(128'hc37ddf5d4e1c94fdb92bb9f2f6718f0f, {16'd57181, 16'd44767, 16'd22995, 16'd9567, 16'd31148, 16'd22025, 16'd10077, 16'd11032, 16'd42044, 16'd11640, 16'd38103, 16'd55547, 16'd749, 16'd5851, 16'd14309, 16'd35690, 16'd58443, 16'd13196, 16'd23222, 16'd38461, 16'd10761, 16'd47032, 16'd28664, 16'd6691, 16'd4629, 16'd54363});
	test_expansion(128'h1de18dd913782ea838cb88fde7e563ef, {16'd33865, 16'd50494, 16'd21288, 16'd2998, 16'd22130, 16'd9628, 16'd44718, 16'd60168, 16'd58126, 16'd8737, 16'd64535, 16'd31349, 16'd41815, 16'd18609, 16'd2308, 16'd36326, 16'd30957, 16'd13604, 16'd53288, 16'd4947, 16'd28798, 16'd700, 16'd33885, 16'd21490, 16'd34784, 16'd25053});
	test_expansion(128'h8b8b17b6c1c8c9993270033a42aaca45, {16'd25799, 16'd48200, 16'd3641, 16'd4852, 16'd17642, 16'd5936, 16'd3030, 16'd50310, 16'd62962, 16'd10284, 16'd63924, 16'd9438, 16'd10988, 16'd18320, 16'd59077, 16'd62587, 16'd46810, 16'd3926, 16'd35822, 16'd37483, 16'd51638, 16'd20023, 16'd37004, 16'd56361, 16'd55332, 16'd25710});
	test_expansion(128'hdcf1dad29ee602dcc024469ca752826c, {16'd42404, 16'd40906, 16'd14488, 16'd46250, 16'd3881, 16'd15480, 16'd9102, 16'd1376, 16'd46922, 16'd19442, 16'd62921, 16'd9525, 16'd46160, 16'd25001, 16'd9112, 16'd34003, 16'd58630, 16'd54819, 16'd62056, 16'd29104, 16'd23054, 16'd65034, 16'd52246, 16'd41409, 16'd16605, 16'd37558});
	test_expansion(128'h3c66763744493fb802e7d895d73c50e5, {16'd52163, 16'd53150, 16'd1250, 16'd37094, 16'd46623, 16'd46539, 16'd64350, 16'd10967, 16'd51920, 16'd4284, 16'd9480, 16'd26734, 16'd30362, 16'd11455, 16'd62792, 16'd15481, 16'd53221, 16'd28975, 16'd35458, 16'd50557, 16'd8149, 16'd14204, 16'd19607, 16'd57741, 16'd6943, 16'd56375});
	test_expansion(128'h831fcabfe17a89f21b4502e1d840f9b8, {16'd62901, 16'd21473, 16'd23381, 16'd12421, 16'd46999, 16'd50327, 16'd35495, 16'd29189, 16'd12444, 16'd10604, 16'd42468, 16'd4681, 16'd55426, 16'd18570, 16'd14051, 16'd62646, 16'd6744, 16'd54458, 16'd29281, 16'd21842, 16'd16709, 16'd376, 16'd47652, 16'd55242, 16'd24007, 16'd63150});
	test_expansion(128'h04d94149d25432fe65f84fb2d5f4240d, {16'd739, 16'd11115, 16'd55232, 16'd21677, 16'd31828, 16'd39590, 16'd25279, 16'd58750, 16'd13250, 16'd7870, 16'd24110, 16'd57550, 16'd13310, 16'd18347, 16'd46946, 16'd55311, 16'd12403, 16'd28720, 16'd63852, 16'd24236, 16'd5929, 16'd30214, 16'd5700, 16'd64638, 16'd40476, 16'd27034});
	test_expansion(128'hff131e80dff375891d127fb3a7c4387b, {16'd50278, 16'd21975, 16'd62551, 16'd1012, 16'd33961, 16'd61149, 16'd42633, 16'd27153, 16'd14697, 16'd52731, 16'd42968, 16'd13301, 16'd9361, 16'd9983, 16'd27635, 16'd34046, 16'd19805, 16'd1022, 16'd64034, 16'd12473, 16'd28640, 16'd3554, 16'd25802, 16'd26005, 16'd17024, 16'd1825});
	test_expansion(128'h453739899b9f0774e7d476ec790573dc, {16'd9516, 16'd7959, 16'd39985, 16'd30096, 16'd30686, 16'd26575, 16'd35532, 16'd5657, 16'd15642, 16'd4689, 16'd37618, 16'd57233, 16'd6513, 16'd2651, 16'd16438, 16'd36594, 16'd46208, 16'd26744, 16'd6066, 16'd32438, 16'd24606, 16'd53934, 16'd2380, 16'd39307, 16'd19405, 16'd17847});
	test_expansion(128'h8c2b7581515878efd8909f4bc2d8202a, {16'd60867, 16'd13304, 16'd379, 16'd61395, 16'd32552, 16'd3414, 16'd47922, 16'd19977, 16'd39378, 16'd50116, 16'd13453, 16'd9188, 16'd26929, 16'd10510, 16'd49348, 16'd39944, 16'd21615, 16'd6262, 16'd34111, 16'd18067, 16'd5736, 16'd42040, 16'd23202, 16'd23247, 16'd43279, 16'd41164});
	test_expansion(128'hba505a71caadd7b2eb9c1595f3c0679f, {16'd45563, 16'd41076, 16'd41445, 16'd22916, 16'd38968, 16'd52658, 16'd24734, 16'd62046, 16'd47475, 16'd48035, 16'd36455, 16'd3135, 16'd17374, 16'd32077, 16'd5037, 16'd14327, 16'd56634, 16'd38744, 16'd32618, 16'd12550, 16'd45385, 16'd34645, 16'd31149, 16'd9808, 16'd33153, 16'd34544});
	test_expansion(128'hc3b47a0705642a5d70f9dcb68bf08364, {16'd15564, 16'd15775, 16'd16925, 16'd62796, 16'd17446, 16'd25004, 16'd13734, 16'd61796, 16'd9041, 16'd33649, 16'd63226, 16'd23351, 16'd63574, 16'd9080, 16'd18427, 16'd50829, 16'd52766, 16'd48327, 16'd46781, 16'd21030, 16'd21817, 16'd56041, 16'd50720, 16'd2134, 16'd17415, 16'd9653});
	test_expansion(128'h74aae879e71bf0a8144cf7f77f47bf7e, {16'd46888, 16'd55659, 16'd58391, 16'd10815, 16'd40221, 16'd41175, 16'd8021, 16'd6250, 16'd34617, 16'd34010, 16'd48882, 16'd13986, 16'd29248, 16'd9778, 16'd28509, 16'd53334, 16'd10278, 16'd35035, 16'd8920, 16'd48295, 16'd22214, 16'd16237, 16'd4394, 16'd29808, 16'd1919, 16'd28420});
	test_expansion(128'h8724a3f7577d505db25ec6c59ff6531d, {16'd53156, 16'd38610, 16'd7447, 16'd1379, 16'd8120, 16'd14266, 16'd53657, 16'd35761, 16'd7252, 16'd4402, 16'd52199, 16'd30613, 16'd3228, 16'd54010, 16'd63202, 16'd37062, 16'd39226, 16'd60489, 16'd29188, 16'd33406, 16'd52795, 16'd2237, 16'd41443, 16'd5674, 16'd4928, 16'd29033});
	test_expansion(128'hfa5f921c06f7ece18c0ca7564cc370f8, {16'd7632, 16'd62489, 16'd30175, 16'd13580, 16'd27246, 16'd4972, 16'd32291, 16'd5182, 16'd42674, 16'd45235, 16'd30473, 16'd15498, 16'd8136, 16'd21798, 16'd17873, 16'd25074, 16'd42739, 16'd37152, 16'd45174, 16'd36963, 16'd60165, 16'd27300, 16'd19874, 16'd11779, 16'd34876, 16'd358});
	test_expansion(128'h036173eb6f3276b846339a601731910a, {16'd14628, 16'd10831, 16'd49386, 16'd35112, 16'd15591, 16'd45765, 16'd64110, 16'd30936, 16'd57558, 16'd48062, 16'd22814, 16'd32860, 16'd55422, 16'd988, 16'd8725, 16'd32299, 16'd23933, 16'd4401, 16'd52598, 16'd28303, 16'd37619, 16'd32544, 16'd46179, 16'd53118, 16'd36031, 16'd24015});
	test_expansion(128'h394e1c88e6107d326a14e5448fd244f4, {16'd65103, 16'd59227, 16'd56912, 16'd29842, 16'd41131, 16'd28174, 16'd37137, 16'd51013, 16'd55815, 16'd22868, 16'd31325, 16'd43162, 16'd64117, 16'd29581, 16'd48183, 16'd24104, 16'd18894, 16'd59522, 16'd22500, 16'd32122, 16'd47647, 16'd10214, 16'd63681, 16'd20158, 16'd23704, 16'd50219});
	test_expansion(128'h9f47630a9dcd5d310c9ee5c949ce474e, {16'd35635, 16'd49243, 16'd23503, 16'd33036, 16'd681, 16'd20441, 16'd32513, 16'd46542, 16'd13623, 16'd25130, 16'd19361, 16'd16928, 16'd9054, 16'd3248, 16'd39801, 16'd41850, 16'd53736, 16'd45235, 16'd31439, 16'd54349, 16'd61567, 16'd27276, 16'd42607, 16'd8241, 16'd24765, 16'd53502});
	test_expansion(128'h8bfc63d382cd9ff2bf3ab6e1835c3dbf, {16'd13346, 16'd54786, 16'd56203, 16'd49198, 16'd5689, 16'd1740, 16'd6028, 16'd55161, 16'd17840, 16'd17044, 16'd7766, 16'd32716, 16'd37373, 16'd2061, 16'd15998, 16'd40880, 16'd48400, 16'd18873, 16'd44351, 16'd31854, 16'd50746, 16'd63018, 16'd56763, 16'd31038, 16'd33416, 16'd54203});
	test_expansion(128'hd12c40c60da178a289ffc25d30e836a6, {16'd512, 16'd4232, 16'd12617, 16'd16115, 16'd46765, 16'd41333, 16'd63570, 16'd41106, 16'd30353, 16'd54555, 16'd9339, 16'd44513, 16'd29641, 16'd51430, 16'd42438, 16'd6221, 16'd61777, 16'd28698, 16'd19167, 16'd17610, 16'd11994, 16'd4084, 16'd16325, 16'd31863, 16'd35848, 16'd20466});
	test_expansion(128'h41e3872f6a637ea324714896bd10133f, {16'd64286, 16'd1735, 16'd60187, 16'd25162, 16'd34686, 16'd29432, 16'd6050, 16'd4223, 16'd29075, 16'd8209, 16'd35035, 16'd39035, 16'd18670, 16'd29907, 16'd60422, 16'd14917, 16'd24918, 16'd54668, 16'd36529, 16'd24386, 16'd26331, 16'd33120, 16'd16584, 16'd32435, 16'd33742, 16'd44219});
	test_expansion(128'hb216740f558fb55795281fcd6e3b3a79, {16'd24933, 16'd20989, 16'd10079, 16'd33337, 16'd13816, 16'd28150, 16'd61645, 16'd22303, 16'd3902, 16'd2448, 16'd1483, 16'd44449, 16'd19663, 16'd38636, 16'd47406, 16'd5963, 16'd63775, 16'd55727, 16'd35354, 16'd7015, 16'd61309, 16'd30873, 16'd53424, 16'd61767, 16'd30796, 16'd44719});
	test_expansion(128'h895adbbc9633e5617f491e184b355c5f, {16'd416, 16'd30636, 16'd17982, 16'd61695, 16'd16211, 16'd34440, 16'd12738, 16'd32473, 16'd47982, 16'd15216, 16'd14530, 16'd46708, 16'd51738, 16'd32586, 16'd24068, 16'd33537, 16'd12122, 16'd44355, 16'd14442, 16'd34884, 16'd47250, 16'd1577, 16'd40782, 16'd39375, 16'd37065, 16'd58722});
	test_expansion(128'hf7e529f05cd86106db21584f3af969ba, {16'd20284, 16'd60881, 16'd31528, 16'd8177, 16'd1156, 16'd47633, 16'd39380, 16'd62542, 16'd63653, 16'd2618, 16'd13474, 16'd5807, 16'd60312, 16'd1574, 16'd58095, 16'd15753, 16'd49416, 16'd12087, 16'd30986, 16'd63477, 16'd22924, 16'd29738, 16'd6153, 16'd23528, 16'd58424, 16'd62513});
	test_expansion(128'h29dac8490f7df9fa38a07ee4b9ec9422, {16'd6223, 16'd6107, 16'd15781, 16'd45078, 16'd23351, 16'd50777, 16'd47213, 16'd50835, 16'd20275, 16'd36074, 16'd49959, 16'd58213, 16'd5415, 16'd47905, 16'd22832, 16'd20838, 16'd5562, 16'd25349, 16'd13805, 16'd24229, 16'd18554, 16'd29428, 16'd63405, 16'd13339, 16'd49640, 16'd35499});
	test_expansion(128'h140b540a34d2df08013f85e7f746a122, {16'd3777, 16'd14554, 16'd632, 16'd38069, 16'd9469, 16'd55045, 16'd27596, 16'd17906, 16'd59450, 16'd55254, 16'd50462, 16'd13346, 16'd35832, 16'd53562, 16'd22134, 16'd4517, 16'd60374, 16'd19427, 16'd25200, 16'd13650, 16'd15206, 16'd22939, 16'd23557, 16'd52900, 16'd12366, 16'd1885});
	test_expansion(128'h78caa5f26bcb163b19a7130154fe6558, {16'd9056, 16'd9400, 16'd54296, 16'd4801, 16'd36196, 16'd4438, 16'd41619, 16'd15874, 16'd24943, 16'd27458, 16'd38598, 16'd49097, 16'd43286, 16'd51665, 16'd46656, 16'd25483, 16'd57260, 16'd10237, 16'd50254, 16'd60909, 16'd22230, 16'd40631, 16'd36421, 16'd57701, 16'd13133, 16'd35768});
	test_expansion(128'hb0658fb33b1901b1f57e7bb6a60f3a7d, {16'd25110, 16'd49555, 16'd59991, 16'd9989, 16'd8997, 16'd41601, 16'd63248, 16'd26062, 16'd4476, 16'd15635, 16'd61137, 16'd4560, 16'd39438, 16'd21853, 16'd45315, 16'd14546, 16'd30780, 16'd47252, 16'd58085, 16'd59086, 16'd42265, 16'd42430, 16'd58825, 16'd63253, 16'd8975, 16'd41684});
	test_expansion(128'h9d6f641807f688f0f6d94397b206d138, {16'd48502, 16'd3986, 16'd62383, 16'd46673, 16'd10672, 16'd42779, 16'd24959, 16'd7913, 16'd59684, 16'd7864, 16'd37427, 16'd56272, 16'd23429, 16'd16128, 16'd60596, 16'd16835, 16'd30215, 16'd6176, 16'd3206, 16'd19594, 16'd34441, 16'd50632, 16'd37652, 16'd4999, 16'd10041, 16'd7822});
	test_expansion(128'h747c473ff8c4496add10b98b38b3e8b2, {16'd44006, 16'd24151, 16'd6997, 16'd49119, 16'd9560, 16'd34251, 16'd20368, 16'd37792, 16'd25976, 16'd35013, 16'd24238, 16'd48917, 16'd37384, 16'd34621, 16'd59814, 16'd51089, 16'd30222, 16'd59661, 16'd21616, 16'd1746, 16'd17285, 16'd10843, 16'd52386, 16'd21154, 16'd39430, 16'd15889});
	test_expansion(128'h135a9da331808fdd157688b41eef8104, {16'd12130, 16'd60459, 16'd37044, 16'd45624, 16'd38212, 16'd35920, 16'd42929, 16'd45414, 16'd42090, 16'd33175, 16'd42357, 16'd50494, 16'd42044, 16'd51197, 16'd45562, 16'd41054, 16'd3249, 16'd30482, 16'd16819, 16'd50826, 16'd23311, 16'd32760, 16'd40244, 16'd205, 16'd56145, 16'd21150});
	test_expansion(128'he9d473d1e6f64f189e6d53d54040020e, {16'd64320, 16'd21176, 16'd39506, 16'd22155, 16'd31338, 16'd64197, 16'd51362, 16'd39435, 16'd35577, 16'd38810, 16'd46703, 16'd15170, 16'd47891, 16'd18907, 16'd45910, 16'd23166, 16'd63016, 16'd21274, 16'd51383, 16'd27845, 16'd1220, 16'd65184, 16'd1850, 16'd41940, 16'd16025, 16'd12982});
	test_expansion(128'he4eb7a89f40b8756d57d9d125986e753, {16'd11934, 16'd64842, 16'd27033, 16'd4914, 16'd3366, 16'd26916, 16'd9524, 16'd12706, 16'd3970, 16'd65229, 16'd52083, 16'd35079, 16'd6378, 16'd3313, 16'd13456, 16'd31010, 16'd46794, 16'd34590, 16'd14640, 16'd29574, 16'd27702, 16'd58591, 16'd12549, 16'd2017, 16'd48060, 16'd45256});
	test_expansion(128'hded0cc24b4e356d04a227f54adeba8ca, {16'd39555, 16'd3672, 16'd42578, 16'd53804, 16'd24236, 16'd45197, 16'd51996, 16'd29200, 16'd12655, 16'd31385, 16'd1853, 16'd29675, 16'd50050, 16'd5282, 16'd12682, 16'd47683, 16'd17351, 16'd20036, 16'd39114, 16'd23204, 16'd64917, 16'd60079, 16'd32152, 16'd42960, 16'd24413, 16'd57809});
	test_expansion(128'hf4133316bf674097361f74fb7d887e75, {16'd44848, 16'd64894, 16'd24510, 16'd26154, 16'd35492, 16'd19129, 16'd58952, 16'd5884, 16'd23616, 16'd46123, 16'd52933, 16'd18516, 16'd106, 16'd52900, 16'd23503, 16'd59106, 16'd23465, 16'd60248, 16'd2153, 16'd50983, 16'd12674, 16'd58464, 16'd17436, 16'd36869, 16'd49249, 16'd49888});
	test_expansion(128'h073e899e9b495d2c53ba2b8f3dcdd50e, {16'd18118, 16'd14289, 16'd21774, 16'd28101, 16'd61126, 16'd31752, 16'd31080, 16'd10485, 16'd7567, 16'd24052, 16'd8394, 16'd39773, 16'd7377, 16'd65007, 16'd64608, 16'd22739, 16'd35227, 16'd35498, 16'd30541, 16'd31155, 16'd64642, 16'd30062, 16'd6676, 16'd13717, 16'd887, 16'd9117});
	test_expansion(128'hc78872b394f1ca300b90c6b19438fbdb, {16'd19669, 16'd17087, 16'd19646, 16'd38794, 16'd51806, 16'd52302, 16'd29042, 16'd55108, 16'd4851, 16'd49446, 16'd17789, 16'd43813, 16'd24747, 16'd11258, 16'd36858, 16'd12036, 16'd65487, 16'd58361, 16'd45753, 16'd58424, 16'd58853, 16'd57058, 16'd11132, 16'd54618, 16'd48843, 16'd27094});
	test_expansion(128'haea0824ace72d3e1e5cc22246faeda0c, {16'd3910, 16'd20255, 16'd45148, 16'd56330, 16'd11975, 16'd11391, 16'd54171, 16'd6862, 16'd56314, 16'd1412, 16'd39630, 16'd32952, 16'd64409, 16'd24473, 16'd6361, 16'd1019, 16'd24359, 16'd62652, 16'd53918, 16'd47524, 16'd44470, 16'd3046, 16'd49823, 16'd44094, 16'd6149, 16'd46687});
	test_expansion(128'hd5ade93f2f548930a34fbf6e1037cbeb, {16'd33603, 16'd59655, 16'd31488, 16'd33421, 16'd49918, 16'd57816, 16'd11179, 16'd39597, 16'd57697, 16'd27416, 16'd25772, 16'd42947, 16'd35730, 16'd2842, 16'd60515, 16'd17276, 16'd2774, 16'd51814, 16'd24286, 16'd42773, 16'd47939, 16'd56615, 16'd15167, 16'd11555, 16'd57208, 16'd37093});
	test_expansion(128'hb55f88ff0fb9e1c29b6c268484a7b47e, {16'd10461, 16'd61418, 16'd59398, 16'd38584, 16'd52652, 16'd17792, 16'd30211, 16'd40851, 16'd15595, 16'd13611, 16'd4820, 16'd548, 16'd63381, 16'd57298, 16'd35084, 16'd21305, 16'd40536, 16'd44078, 16'd25972, 16'd57929, 16'd22013, 16'd62952, 16'd29735, 16'd9404, 16'd1495, 16'd12355});
	test_expansion(128'h2b92b02b119f5932147d0fc458b1aaf0, {16'd17934, 16'd50998, 16'd2876, 16'd12243, 16'd30450, 16'd9773, 16'd61864, 16'd47192, 16'd332, 16'd60582, 16'd7670, 16'd49084, 16'd21300, 16'd18933, 16'd35591, 16'd30809, 16'd65178, 16'd47614, 16'd1262, 16'd19872, 16'd38533, 16'd34921, 16'd36639, 16'd5018, 16'd60414, 16'd14324});
	test_expansion(128'h055029ee00a44eec9253e175652730ac, {16'd15094, 16'd57318, 16'd19885, 16'd10728, 16'd36624, 16'd54848, 16'd5248, 16'd7995, 16'd40119, 16'd35378, 16'd2240, 16'd19338, 16'd51177, 16'd26153, 16'd17792, 16'd1887, 16'd44980, 16'd53473, 16'd49052, 16'd29691, 16'd19651, 16'd14729, 16'd36106, 16'd61034, 16'd8798, 16'd29009});
	test_expansion(128'h7a2fcd5ecf0955b4b71ded7f7a8401f4, {16'd41305, 16'd57083, 16'd53506, 16'd14391, 16'd46726, 16'd7694, 16'd15894, 16'd12762, 16'd47144, 16'd29247, 16'd33684, 16'd6632, 16'd42824, 16'd25034, 16'd37086, 16'd29139, 16'd2088, 16'd31961, 16'd50592, 16'd52837, 16'd9514, 16'd38907, 16'd443, 16'd12752, 16'd51624, 16'd47360});
	test_expansion(128'h431d5279182f9b165aa9b7acf73bf249, {16'd56823, 16'd48932, 16'd17776, 16'd46368, 16'd38966, 16'd28685, 16'd21754, 16'd56941, 16'd33132, 16'd253, 16'd57904, 16'd48392, 16'd5851, 16'd7511, 16'd50648, 16'd20281, 16'd23021, 16'd10416, 16'd36724, 16'd43126, 16'd13411, 16'd12780, 16'd30268, 16'd25815, 16'd25124, 16'd31521});
	test_expansion(128'hc753284d53febaba9ebbedc6bc045cef, {16'd34543, 16'd50180, 16'd44833, 16'd25726, 16'd44661, 16'd40720, 16'd14922, 16'd47884, 16'd47608, 16'd65156, 16'd21675, 16'd9203, 16'd7775, 16'd47409, 16'd6970, 16'd20257, 16'd62770, 16'd30266, 16'd50800, 16'd52193, 16'd31731, 16'd6302, 16'd65174, 16'd38076, 16'd20642, 16'd45263});
	test_expansion(128'h6d0615ca358cc9984d07a622f2180d02, {16'd38269, 16'd29424, 16'd27091, 16'd2799, 16'd3930, 16'd35583, 16'd5634, 16'd28447, 16'd64697, 16'd13797, 16'd10888, 16'd13700, 16'd56132, 16'd7313, 16'd11960, 16'd36162, 16'd61869, 16'd65327, 16'd20732, 16'd20557, 16'd21848, 16'd44916, 16'd25204, 16'd48815, 16'd40341, 16'd30632});
	test_expansion(128'ha79b2997982311f9d8f58b63aa753ab8, {16'd23324, 16'd53092, 16'd16169, 16'd24129, 16'd5403, 16'd44425, 16'd42482, 16'd34653, 16'd36523, 16'd28709, 16'd36257, 16'd5041, 16'd62159, 16'd1866, 16'd53650, 16'd58324, 16'd2920, 16'd17351, 16'd9905, 16'd27127, 16'd20210, 16'd4739, 16'd62205, 16'd55058, 16'd43338, 16'd50148});
	test_expansion(128'hdf5ef206ab863e90a7c9b939d1317361, {16'd37046, 16'd11321, 16'd50428, 16'd32020, 16'd7542, 16'd16528, 16'd49228, 16'd41283, 16'd19838, 16'd12764, 16'd40073, 16'd10858, 16'd44653, 16'd44793, 16'd54616, 16'd27567, 16'd52659, 16'd12890, 16'd33926, 16'd59143, 16'd62508, 16'd8740, 16'd42346, 16'd62436, 16'd42854, 16'd46035});
	test_expansion(128'h5650b58e4c5293743ef3adcb4bcec7e5, {16'd25646, 16'd39578, 16'd10172, 16'd11709, 16'd31103, 16'd38443, 16'd17262, 16'd11529, 16'd22694, 16'd17570, 16'd39426, 16'd18036, 16'd47676, 16'd50391, 16'd18307, 16'd42350, 16'd43342, 16'd21929, 16'd29920, 16'd37946, 16'd43160, 16'd13924, 16'd50433, 16'd11280, 16'd6131, 16'd43747});
	test_expansion(128'h10f9334c66c8827b6da04cfdec66fa64, {16'd34804, 16'd51727, 16'd60704, 16'd51643, 16'd15944, 16'd8480, 16'd12342, 16'd7591, 16'd55245, 16'd35955, 16'd45720, 16'd29274, 16'd56703, 16'd50876, 16'd18806, 16'd47426, 16'd4462, 16'd37146, 16'd60006, 16'd24466, 16'd2411, 16'd13709, 16'd8004, 16'd1121, 16'd41267, 16'd13620});
	test_expansion(128'h1e389055c7bbc4e49da70ae4031a08b1, {16'd64605, 16'd21091, 16'd5619, 16'd44562, 16'd13058, 16'd49525, 16'd24328, 16'd2329, 16'd665, 16'd17957, 16'd57861, 16'd11505, 16'd22350, 16'd61655, 16'd17592, 16'd27137, 16'd50746, 16'd28231, 16'd23254, 16'd56617, 16'd61479, 16'd4024, 16'd21598, 16'd47143, 16'd55128, 16'd6449});
	test_expansion(128'h3e21862b7fbacfb69c5d6ad7b37b0726, {16'd23980, 16'd52560, 16'd39499, 16'd20062, 16'd14522, 16'd17272, 16'd43522, 16'd21202, 16'd34940, 16'd64209, 16'd38100, 16'd37455, 16'd34566, 16'd20631, 16'd34847, 16'd44848, 16'd36006, 16'd2697, 16'd1791, 16'd2293, 16'd59133, 16'd90, 16'd55846, 16'd44234, 16'd45122, 16'd37224});
	test_expansion(128'h92cbdebc5470e87cd5b54bc35a842796, {16'd35086, 16'd8849, 16'd35175, 16'd54168, 16'd57354, 16'd8140, 16'd62337, 16'd59354, 16'd392, 16'd56513, 16'd7157, 16'd28675, 16'd5747, 16'd60530, 16'd24046, 16'd26695, 16'd50015, 16'd22808, 16'd33876, 16'd45534, 16'd30650, 16'd40427, 16'd9750, 16'd140, 16'd1907, 16'd52219});
	test_expansion(128'h0f39c0b13a694323f9cd22fe906d7b99, {16'd25296, 16'd48973, 16'd49067, 16'd21625, 16'd46257, 16'd9743, 16'd8480, 16'd59770, 16'd51465, 16'd33132, 16'd11104, 16'd8514, 16'd16655, 16'd29988, 16'd27691, 16'd7286, 16'd24059, 16'd5004, 16'd49061, 16'd63553, 16'd60999, 16'd5758, 16'd31922, 16'd42150, 16'd61791, 16'd31129});
	test_expansion(128'ha19b62de48d7fa12d7c32f60e924913b, {16'd42733, 16'd6846, 16'd60660, 16'd11718, 16'd15824, 16'd56930, 16'd19490, 16'd51660, 16'd33213, 16'd23780, 16'd37820, 16'd48327, 16'd53807, 16'd56447, 16'd23459, 16'd44657, 16'd33751, 16'd2736, 16'd24123, 16'd51711, 16'd4813, 16'd32259, 16'd53729, 16'd54728, 16'd36984, 16'd34546});
	test_expansion(128'ha75ba8a8a84f47bd5b3ad79d9e821d38, {16'd52310, 16'd43607, 16'd17554, 16'd14970, 16'd61202, 16'd46598, 16'd289, 16'd45965, 16'd23517, 16'd43425, 16'd50764, 16'd63276, 16'd8419, 16'd59258, 16'd47055, 16'd37647, 16'd39524, 16'd14283, 16'd54676, 16'd30332, 16'd50266, 16'd2934, 16'd50653, 16'd749, 16'd25754, 16'd42412});
	test_expansion(128'hfda5f72b50525b97c5c8b8eecd2f71e4, {16'd62220, 16'd51630, 16'd51417, 16'd23147, 16'd33711, 16'd13801, 16'd13331, 16'd65522, 16'd158, 16'd22857, 16'd37312, 16'd11341, 16'd30622, 16'd65064, 16'd8400, 16'd64134, 16'd15491, 16'd3076, 16'd38932, 16'd35692, 16'd64160, 16'd21796, 16'd3300, 16'd11534, 16'd51432, 16'd19306});
	test_expansion(128'h17fb688cadae2cfec39c71fb44d7f94f, {16'd2350, 16'd27034, 16'd9232, 16'd38739, 16'd37489, 16'd56808, 16'd57492, 16'd25485, 16'd46384, 16'd13087, 16'd19855, 16'd31538, 16'd38559, 16'd61090, 16'd13767, 16'd17720, 16'd36387, 16'd53571, 16'd7186, 16'd27670, 16'd45740, 16'd3929, 16'd27999, 16'd45448, 16'd48455, 16'd13168});
	test_expansion(128'hfff228109cbbdaca105ffcf5483d8c6a, {16'd25658, 16'd45971, 16'd7016, 16'd30481, 16'd53196, 16'd42534, 16'd16829, 16'd22391, 16'd64910, 16'd9017, 16'd18333, 16'd24468, 16'd3947, 16'd26350, 16'd33855, 16'd11907, 16'd34790, 16'd42314, 16'd53675, 16'd50742, 16'd28753, 16'd16594, 16'd54278, 16'd43905, 16'd17536, 16'd64471});
	test_expansion(128'h9b52e5b4758027b61555de39b891b2d1, {16'd17406, 16'd64820, 16'd53780, 16'd59796, 16'd20897, 16'd33386, 16'd57845, 16'd51506, 16'd62565, 16'd37580, 16'd57643, 16'd16449, 16'd63006, 16'd45311, 16'd24610, 16'd23744, 16'd35804, 16'd49219, 16'd60137, 16'd33338, 16'd17766, 16'd44636, 16'd64869, 16'd38054, 16'd44664, 16'd857});
	test_expansion(128'h84ec6e0c02e92a0c67283741577107c2, {16'd47330, 16'd29595, 16'd24558, 16'd32054, 16'd44130, 16'd5077, 16'd14202, 16'd33637, 16'd44872, 16'd5578, 16'd15446, 16'd16089, 16'd37114, 16'd18220, 16'd24879, 16'd57198, 16'd894, 16'd1701, 16'd31391, 16'd22071, 16'd14476, 16'd42031, 16'd58914, 16'd63850, 16'd30507, 16'd22588});
	test_expansion(128'he22a7c53e362df4eaf2747ead21643fd, {16'd26993, 16'd40222, 16'd47829, 16'd11916, 16'd8404, 16'd7346, 16'd20522, 16'd40931, 16'd61729, 16'd48865, 16'd60454, 16'd5760, 16'd63091, 16'd54796, 16'd35934, 16'd45642, 16'd47146, 16'd13534, 16'd11140, 16'd26374, 16'd43053, 16'd9777, 16'd31730, 16'd18947, 16'd42312, 16'd36364});
	test_expansion(128'h8ccae1722abd5772652d37cb205d7565, {16'd46998, 16'd17333, 16'd48295, 16'd52863, 16'd31520, 16'd37642, 16'd21943, 16'd39545, 16'd65081, 16'd61671, 16'd35986, 16'd19806, 16'd45972, 16'd34607, 16'd13574, 16'd2239, 16'd52927, 16'd16555, 16'd33216, 16'd34832, 16'd60737, 16'd23451, 16'd3682, 16'd51808, 16'd51104, 16'd36174});
	test_expansion(128'h7b1378027e35759a85a2e3d7941fe714, {16'd14194, 16'd31473, 16'd7649, 16'd62788, 16'd19631, 16'd10539, 16'd42729, 16'd17344, 16'd17795, 16'd51349, 16'd62924, 16'd15864, 16'd47777, 16'd22968, 16'd1316, 16'd38341, 16'd51300, 16'd26701, 16'd13858, 16'd6518, 16'd24978, 16'd64014, 16'd597, 16'd40444, 16'd37936, 16'd3753});
	test_expansion(128'hd7ccfa80911f6e33f4cf171b32309b9b, {16'd64691, 16'd25530, 16'd9491, 16'd40829, 16'd62356, 16'd55416, 16'd1467, 16'd20134, 16'd32969, 16'd54675, 16'd10364, 16'd37085, 16'd8221, 16'd13725, 16'd15737, 16'd31484, 16'd36342, 16'd31687, 16'd18274, 16'd49986, 16'd56836, 16'd32669, 16'd45163, 16'd37168, 16'd21152, 16'd65412});
	test_expansion(128'h1ece6c90191e1e24e16e972de2aca395, {16'd42668, 16'd29921, 16'd40239, 16'd35694, 16'd6686, 16'd48439, 16'd40505, 16'd21630, 16'd31453, 16'd19511, 16'd41578, 16'd29697, 16'd2639, 16'd59903, 16'd53219, 16'd33582, 16'd22936, 16'd9129, 16'd32481, 16'd60956, 16'd49455, 16'd25718, 16'd8888, 16'd50844, 16'd5382, 16'd9362});
	test_expansion(128'heafff5d5dde702a90eaba3e1ae3c0fb0, {16'd58840, 16'd3180, 16'd7486, 16'd63171, 16'd36187, 16'd50069, 16'd52303, 16'd56507, 16'd41162, 16'd12732, 16'd53275, 16'd8581, 16'd55242, 16'd49776, 16'd3222, 16'd14784, 16'd28035, 16'd43180, 16'd50590, 16'd22507, 16'd52550, 16'd45333, 16'd56030, 16'd24487, 16'd2817, 16'd42762});
	test_expansion(128'h5320a240b456e06f28f6aebde6abb7f6, {16'd11011, 16'd15330, 16'd18830, 16'd50791, 16'd56329, 16'd31893, 16'd56050, 16'd61984, 16'd29305, 16'd48272, 16'd13164, 16'd62571, 16'd8995, 16'd62157, 16'd23676, 16'd60929, 16'd5336, 16'd30486, 16'd36227, 16'd26897, 16'd43208, 16'd36458, 16'd60330, 16'd13589, 16'd20685, 16'd58811});
	test_expansion(128'hb045ee4003a8fcc6d9e7b04234064ec8, {16'd44943, 16'd41912, 16'd1679, 16'd42343, 16'd38290, 16'd40667, 16'd26717, 16'd6843, 16'd15989, 16'd23785, 16'd14642, 16'd10236, 16'd9065, 16'd51051, 16'd32492, 16'd2425, 16'd42167, 16'd37243, 16'd25515, 16'd55751, 16'd37002, 16'd64501, 16'd1421, 16'd65051, 16'd32519, 16'd58570});
	test_expansion(128'hea05c5d3c16c5d0b04cbfe56f774f31d, {16'd14117, 16'd109, 16'd40314, 16'd30994, 16'd12566, 16'd26087, 16'd48410, 16'd12920, 16'd21086, 16'd15517, 16'd56022, 16'd8156, 16'd11784, 16'd45058, 16'd18884, 16'd63208, 16'd11340, 16'd7411, 16'd8772, 16'd23193, 16'd50655, 16'd55634, 16'd20417, 16'd46683, 16'd20966, 16'd28434});
	test_expansion(128'h96b955e58642b06228dac1000c9e2720, {16'd16470, 16'd17570, 16'd62645, 16'd52315, 16'd30842, 16'd54302, 16'd14668, 16'd25516, 16'd56, 16'd21198, 16'd56953, 16'd41383, 16'd6065, 16'd14590, 16'd26292, 16'd44621, 16'd22850, 16'd34075, 16'd3612, 16'd58753, 16'd56081, 16'd18825, 16'd46950, 16'd50768, 16'd17181, 16'd22452});
	test_expansion(128'h8270969c9c84197d0e7468e786ff1f2d, {16'd55485, 16'd11004, 16'd55921, 16'd3391, 16'd41020, 16'd23443, 16'd20050, 16'd14994, 16'd3208, 16'd38667, 16'd30310, 16'd12486, 16'd49374, 16'd15616, 16'd37349, 16'd47047, 16'd8084, 16'd35335, 16'd7808, 16'd49293, 16'd34869, 16'd24761, 16'd42151, 16'd59003, 16'd14345, 16'd2670});
	test_expansion(128'h0a1b63d8a912b5f09f527fd5f66db82a, {16'd42922, 16'd40742, 16'd20535, 16'd41360, 16'd21860, 16'd17790, 16'd55287, 16'd46705, 16'd62637, 16'd43834, 16'd17639, 16'd25035, 16'd51570, 16'd19610, 16'd21106, 16'd30231, 16'd24471, 16'd35966, 16'd28379, 16'd13112, 16'd48766, 16'd57721, 16'd64542, 16'd9427, 16'd27202, 16'd29825});
	test_expansion(128'h196fdf53c6eb9dee28b381f6af6ac4cc, {16'd26440, 16'd58112, 16'd31205, 16'd32348, 16'd49712, 16'd21969, 16'd40828, 16'd49969, 16'd12251, 16'd3444, 16'd43802, 16'd39343, 16'd41712, 16'd41596, 16'd61266, 16'd21125, 16'd125, 16'd33567, 16'd29933, 16'd40124, 16'd14536, 16'd41472, 16'd5786, 16'd39623, 16'd46411, 16'd22824});
	test_expansion(128'h4f04eea63dfa300875a294b0f85a3d6e, {16'd3114, 16'd9290, 16'd5975, 16'd47940, 16'd48168, 16'd54273, 16'd62738, 16'd30006, 16'd49212, 16'd5392, 16'd47299, 16'd61785, 16'd20795, 16'd41575, 16'd39991, 16'd41419, 16'd25255, 16'd7727, 16'd7020, 16'd54106, 16'd49814, 16'd9602, 16'd13338, 16'd56264, 16'd40788, 16'd27027});
	test_expansion(128'h8eb519022849c6107041b2cc76f18b69, {16'd44128, 16'd34168, 16'd12953, 16'd53978, 16'd20558, 16'd1187, 16'd12207, 16'd49627, 16'd24595, 16'd2037, 16'd29052, 16'd58246, 16'd28802, 16'd47794, 16'd22464, 16'd60477, 16'd13810, 16'd48623, 16'd49175, 16'd5881, 16'd49494, 16'd34350, 16'd7341, 16'd17034, 16'd12702, 16'd45620});
	test_expansion(128'h5c3d0898b5262644959bb2ac59d1c74f, {16'd36379, 16'd34961, 16'd57468, 16'd47470, 16'd14078, 16'd16909, 16'd23466, 16'd57107, 16'd19835, 16'd33195, 16'd42846, 16'd59438, 16'd28455, 16'd60766, 16'd37554, 16'd38688, 16'd53114, 16'd60034, 16'd25542, 16'd15227, 16'd10954, 16'd49244, 16'd63431, 16'd50791, 16'd28420, 16'd51808});
	test_expansion(128'h679a14b31fc92681e581cbec9b996be3, {16'd46603, 16'd1661, 16'd243, 16'd29741, 16'd61982, 16'd45414, 16'd46270, 16'd27947, 16'd30629, 16'd14013, 16'd52662, 16'd38033, 16'd56049, 16'd33869, 16'd55929, 16'd3180, 16'd40108, 16'd44358, 16'd24178, 16'd53321, 16'd8336, 16'd63113, 16'd55319, 16'd17652, 16'd35865, 16'd58448});
	test_expansion(128'h37b75f207dec48d9e04b156b7b5c73c6, {16'd33951, 16'd16487, 16'd60372, 16'd47522, 16'd40112, 16'd8584, 16'd6097, 16'd26208, 16'd32389, 16'd35472, 16'd25931, 16'd24393, 16'd51086, 16'd29848, 16'd47082, 16'd8078, 16'd61696, 16'd22172, 16'd40648, 16'd29504, 16'd22548, 16'd8534, 16'd63999, 16'd60811, 16'd10791, 16'd40393});
	test_expansion(128'h321c9751e3236d24c37a34ebe1182450, {16'd21958, 16'd9369, 16'd19475, 16'd43775, 16'd49705, 16'd57209, 16'd40704, 16'd27572, 16'd36302, 16'd28056, 16'd43108, 16'd28434, 16'd38330, 16'd54617, 16'd65113, 16'd21147, 16'd42887, 16'd23367, 16'd23144, 16'd41484, 16'd37105, 16'd9968, 16'd12991, 16'd40693, 16'd8611, 16'd41193});
	test_expansion(128'ha279d39eeb2495912709768b5220e6f7, {16'd173, 16'd5710, 16'd2968, 16'd17831, 16'd57521, 16'd50495, 16'd43809, 16'd20046, 16'd53873, 16'd46985, 16'd22646, 16'd15021, 16'd56148, 16'd26593, 16'd7109, 16'd50287, 16'd26969, 16'd23161, 16'd204, 16'd40223, 16'd10972, 16'd50336, 16'd17135, 16'd844, 16'd46056, 16'd15672});
	test_expansion(128'he34f39c79896fb07b8670fe8fad91f11, {16'd48727, 16'd35711, 16'd56000, 16'd22162, 16'd27083, 16'd29519, 16'd21925, 16'd13968, 16'd6702, 16'd7070, 16'd38510, 16'd53623, 16'd12072, 16'd53948, 16'd6710, 16'd43334, 16'd10102, 16'd15660, 16'd13142, 16'd53040, 16'd17963, 16'd36915, 16'd14254, 16'd32825, 16'd53091, 16'd39652});
	test_expansion(128'ha85b28707cee61e177af7a636bf92205, {16'd22063, 16'd60936, 16'd44308, 16'd32631, 16'd6016, 16'd46480, 16'd19340, 16'd25356, 16'd45307, 16'd3308, 16'd48921, 16'd4270, 16'd51137, 16'd1087, 16'd39000, 16'd21956, 16'd64395, 16'd29692, 16'd46950, 16'd448, 16'd46772, 16'd21659, 16'd46129, 16'd42267, 16'd23842, 16'd45811});
	test_expansion(128'he9965825d2bfad215a74aee033ac678a, {16'd62608, 16'd47104, 16'd14500, 16'd43115, 16'd16689, 16'd16000, 16'd62777, 16'd59603, 16'd4784, 16'd6365, 16'd52173, 16'd11429, 16'd12799, 16'd871, 16'd8243, 16'd56557, 16'd19665, 16'd47220, 16'd37814, 16'd7217, 16'd3679, 16'd31421, 16'd42281, 16'd10474, 16'd43039, 16'd64610});
	test_expansion(128'hb18ff27a2b5eab0925d7bc0d484f5f23, {16'd3899, 16'd8521, 16'd12225, 16'd54236, 16'd36901, 16'd37562, 16'd26723, 16'd15369, 16'd18269, 16'd52377, 16'd41987, 16'd9321, 16'd43943, 16'd31659, 16'd17635, 16'd47689, 16'd20413, 16'd6423, 16'd26958, 16'd49281, 16'd28371, 16'd7787, 16'd8725, 16'd24034, 16'd23330, 16'd62492});
	test_expansion(128'h16b8ce091bb78acb15efe01db9c060a9, {16'd60661, 16'd24431, 16'd25005, 16'd41769, 16'd8235, 16'd10624, 16'd18903, 16'd55878, 16'd45043, 16'd46151, 16'd36633, 16'd7459, 16'd32125, 16'd8604, 16'd2532, 16'd4740, 16'd48464, 16'd21239, 16'd31440, 16'd43877, 16'd26693, 16'd48649, 16'd5991, 16'd37837, 16'd25426, 16'd824});
	test_expansion(128'h8e98ee5f725957e9a35505e4767a01dd, {16'd61842, 16'd51795, 16'd14513, 16'd31135, 16'd42629, 16'd20507, 16'd16526, 16'd46855, 16'd10724, 16'd1605, 16'd13037, 16'd47246, 16'd43756, 16'd51444, 16'd59267, 16'd2716, 16'd37364, 16'd43110, 16'd26402, 16'd37106, 16'd43821, 16'd44199, 16'd38753, 16'd13796, 16'd35437, 16'd4595});
	test_expansion(128'hfac7f36ca9fb694452ffd19ddc930a80, {16'd27975, 16'd21766, 16'd36161, 16'd25785, 16'd29881, 16'd52512, 16'd61005, 16'd62689, 16'd29144, 16'd23351, 16'd21997, 16'd58963, 16'd38289, 16'd7081, 16'd51635, 16'd21223, 16'd35161, 16'd38547, 16'd3977, 16'd38438, 16'd40199, 16'd54311, 16'd40642, 16'd6159, 16'd29858, 16'd8592});
	test_expansion(128'hb543b2f5371a52206796cecd119fcaa5, {16'd561, 16'd51120, 16'd13945, 16'd3991, 16'd10812, 16'd22444, 16'd51912, 16'd42402, 16'd27562, 16'd4959, 16'd63479, 16'd44425, 16'd29662, 16'd22864, 16'd44827, 16'd39401, 16'd30113, 16'd53535, 16'd12362, 16'd2567, 16'd51000, 16'd61541, 16'd43656, 16'd65502, 16'd56478, 16'd5049});
	test_expansion(128'h9659e43624b7d36fd637938a439ba880, {16'd39115, 16'd56031, 16'd58899, 16'd40512, 16'd39621, 16'd51346, 16'd31295, 16'd51340, 16'd12578, 16'd45288, 16'd4496, 16'd21353, 16'd20840, 16'd60886, 16'd62327, 16'd30696, 16'd31507, 16'd22387, 16'd46214, 16'd53615, 16'd14805, 16'd11587, 16'd31044, 16'd9978, 16'd21001, 16'd29759});
	test_expansion(128'h7f633648e3d77e8be78180504fe7f5f1, {16'd34015, 16'd8156, 16'd46674, 16'd37855, 16'd50784, 16'd63416, 16'd42780, 16'd63497, 16'd1850, 16'd39181, 16'd51810, 16'd32308, 16'd19271, 16'd26637, 16'd50733, 16'd20416, 16'd24251, 16'd43917, 16'd35901, 16'd10237, 16'd25701, 16'd37382, 16'd38353, 16'd3346, 16'd9821, 16'd3026});
	test_expansion(128'h82f8207962c05ec8b04bec0de27c8315, {16'd31036, 16'd848, 16'd2722, 16'd45342, 16'd34887, 16'd42073, 16'd31185, 16'd20272, 16'd30661, 16'd61122, 16'd389, 16'd33879, 16'd3445, 16'd5898, 16'd20000, 16'd8157, 16'd45228, 16'd34230, 16'd22777, 16'd30110, 16'd41688, 16'd36356, 16'd44685, 16'd33952, 16'd1641, 16'd23956});
	test_expansion(128'h77cfe4e6ce06e20800a6b7e961e4e1b8, {16'd4555, 16'd58127, 16'd41221, 16'd27503, 16'd39318, 16'd5029, 16'd46931, 16'd43772, 16'd58497, 16'd64650, 16'd35906, 16'd8012, 16'd842, 16'd5760, 16'd54307, 16'd60853, 16'd8410, 16'd62163, 16'd50414, 16'd45273, 16'd11882, 16'd49169, 16'd38475, 16'd24276, 16'd41397, 16'd39274});
	test_expansion(128'h90cfde926c888628e59a8ec09fdf0803, {16'd24532, 16'd34819, 16'd9240, 16'd37723, 16'd61741, 16'd2143, 16'd48216, 16'd40201, 16'd62612, 16'd33538, 16'd39369, 16'd15436, 16'd40258, 16'd15858, 16'd54752, 16'd30997, 16'd9324, 16'd32065, 16'd358, 16'd23465, 16'd11171, 16'd49248, 16'd58393, 16'd33024, 16'd49200, 16'd54780});
	test_expansion(128'hdf0ba7b40082afceb704ca2015c2c376, {16'd16198, 16'd106, 16'd32857, 16'd1403, 16'd13761, 16'd59948, 16'd11735, 16'd39853, 16'd28033, 16'd50556, 16'd10111, 16'd12380, 16'd52413, 16'd1836, 16'd56912, 16'd39263, 16'd35830, 16'd32612, 16'd60913, 16'd55589, 16'd51871, 16'd61442, 16'd50977, 16'd45020, 16'd58907, 16'd36453});
	test_expansion(128'hff7ee6f215db8ca114a1eada046141fc, {16'd40778, 16'd5333, 16'd29223, 16'd6858, 16'd47620, 16'd12407, 16'd28298, 16'd929, 16'd51150, 16'd33070, 16'd4144, 16'd31099, 16'd12751, 16'd28636, 16'd39356, 16'd19754, 16'd125, 16'd37400, 16'd59691, 16'd21823, 16'd6764, 16'd53340, 16'd13239, 16'd28844, 16'd15764, 16'd49538});
	test_expansion(128'hd816790706018d47714cb1b757292800, {16'd29310, 16'd10402, 16'd64729, 16'd65019, 16'd39498, 16'd19880, 16'd60843, 16'd13074, 16'd39008, 16'd13378, 16'd63439, 16'd42926, 16'd35155, 16'd37404, 16'd59803, 16'd10352, 16'd20725, 16'd42780, 16'd59751, 16'd46446, 16'd42655, 16'd64645, 16'd10927, 16'd33670, 16'd11919, 16'd42550});
	test_expansion(128'h04ff528ca6ac6c4d6c68cc82d247370a, {16'd62191, 16'd4278, 16'd58126, 16'd22742, 16'd21805, 16'd41330, 16'd59909, 16'd24720, 16'd61280, 16'd31634, 16'd41753, 16'd18970, 16'd49537, 16'd16655, 16'd540, 16'd9771, 16'd9679, 16'd52319, 16'd52229, 16'd16060, 16'd6612, 16'd31172, 16'd60781, 16'd12384, 16'd61251, 16'd64028});
	test_expansion(128'hb144258a9366687a58982426a10dfdb9, {16'd49055, 16'd41781, 16'd12628, 16'd4100, 16'd49896, 16'd60727, 16'd17585, 16'd31906, 16'd58242, 16'd10919, 16'd62582, 16'd39727, 16'd22770, 16'd23848, 16'd51000, 16'd61470, 16'd11639, 16'd14851, 16'd51114, 16'd40029, 16'd61230, 16'd57413, 16'd48752, 16'd8964, 16'd4249, 16'd53212});
	test_expansion(128'hd74236036ddb62654d75bc66c06eacbc, {16'd18029, 16'd38888, 16'd51049, 16'd58740, 16'd52518, 16'd56461, 16'd62167, 16'd31614, 16'd56809, 16'd3803, 16'd56214, 16'd38656, 16'd4196, 16'd36933, 16'd19981, 16'd33342, 16'd37195, 16'd9739, 16'd849, 16'd43355, 16'd58521, 16'd28045, 16'd55520, 16'd24746, 16'd10995, 16'd56695});
	test_expansion(128'he2aca46fadbedfb568b883b9a93efa2a, {16'd41372, 16'd45226, 16'd64964, 16'd41694, 16'd7189, 16'd24292, 16'd57718, 16'd11741, 16'd24810, 16'd2875, 16'd61775, 16'd40926, 16'd44397, 16'd61032, 16'd45749, 16'd39834, 16'd4681, 16'd13972, 16'd2397, 16'd64984, 16'd56288, 16'd61627, 16'd6672, 16'd8968, 16'd36247, 16'd26883});
	test_expansion(128'h2de06690fe8638d8ed0f3b7ad612b3e9, {16'd46865, 16'd28057, 16'd23893, 16'd64159, 16'd30364, 16'd39588, 16'd43835, 16'd61287, 16'd2220, 16'd54541, 16'd35797, 16'd21247, 16'd14295, 16'd46297, 16'd50072, 16'd58975, 16'd20899, 16'd3148, 16'd22741, 16'd9811, 16'd5725, 16'd13126, 16'd39338, 16'd64370, 16'd30618, 16'd29658});
	test_expansion(128'h880ed4621a1435da8a6ef678dfe7d8ee, {16'd57246, 16'd22900, 16'd1509, 16'd25210, 16'd27900, 16'd5438, 16'd21314, 16'd48511, 16'd55929, 16'd44655, 16'd31983, 16'd60062, 16'd10814, 16'd19517, 16'd34014, 16'd8226, 16'd56837, 16'd54557, 16'd32530, 16'd64033, 16'd48290, 16'd52236, 16'd54468, 16'd34609, 16'd63847, 16'd21783});
	test_expansion(128'hcbf6c1b5d2992b89ec94817f937e9acb, {16'd29990, 16'd61482, 16'd27858, 16'd42414, 16'd9538, 16'd37539, 16'd27697, 16'd46888, 16'd28163, 16'd38270, 16'd45940, 16'd18809, 16'd56959, 16'd32598, 16'd58000, 16'd12443, 16'd4549, 16'd14605, 16'd18795, 16'd6051, 16'd26653, 16'd46671, 16'd43823, 16'd817, 16'd64610, 16'd10814});
	test_expansion(128'hf1abc64739fbe2676d4fe82f1ff11fc3, {16'd9934, 16'd16623, 16'd58287, 16'd23426, 16'd33794, 16'd3323, 16'd31401, 16'd53941, 16'd21074, 16'd10701, 16'd59297, 16'd32323, 16'd10983, 16'd17580, 16'd6495, 16'd34357, 16'd29779, 16'd62119, 16'd50081, 16'd32883, 16'd35530, 16'd55656, 16'd60356, 16'd65261, 16'd64193, 16'd46533});
	test_expansion(128'h8102052f86057ec146f7dc3a4cf94eca, {16'd45562, 16'd40676, 16'd8346, 16'd42435, 16'd36513, 16'd28863, 16'd56742, 16'd30983, 16'd63319, 16'd21822, 16'd40532, 16'd50986, 16'd37511, 16'd57489, 16'd58020, 16'd7362, 16'd19971, 16'd20341, 16'd13829, 16'd27546, 16'd7276, 16'd15781, 16'd16246, 16'd15166, 16'd43932, 16'd32133});
	test_expansion(128'h8c06201c3e1f2de21b764731714d8cc1, {16'd36832, 16'd59075, 16'd13885, 16'd14677, 16'd52852, 16'd24415, 16'd871, 16'd31276, 16'd46409, 16'd19146, 16'd32041, 16'd21780, 16'd39114, 16'd18015, 16'd47800, 16'd22746, 16'd11874, 16'd47733, 16'd45339, 16'd43111, 16'd13519, 16'd58708, 16'd40418, 16'd6846, 16'd65277, 16'd28181});
	test_expansion(128'h84ce6f5021e921898572969ddc2fb1e3, {16'd25963, 16'd20740, 16'd51976, 16'd36017, 16'd16525, 16'd62449, 16'd9092, 16'd52852, 16'd19345, 16'd8585, 16'd3379, 16'd49189, 16'd22201, 16'd17006, 16'd37937, 16'd29923, 16'd20829, 16'd28066, 16'd8914, 16'd24760, 16'd40980, 16'd23047, 16'd57149, 16'd40856, 16'd61312, 16'd2029});
	test_expansion(128'h029ec57994fbd99c7203fe7b6ef10a46, {16'd4081, 16'd51870, 16'd24231, 16'd16027, 16'd53863, 16'd6731, 16'd51509, 16'd31916, 16'd31866, 16'd10384, 16'd56449, 16'd64759, 16'd51008, 16'd1977, 16'd4192, 16'd36664, 16'd26576, 16'd28374, 16'd51859, 16'd41829, 16'd56801, 16'd28254, 16'd17316, 16'd11268, 16'd13521, 16'd46536});
	test_expansion(128'h913cad22ac4ddd5e4799963bf8e54ca8, {16'd35552, 16'd42592, 16'd31155, 16'd25443, 16'd44452, 16'd31098, 16'd54296, 16'd53740, 16'd26171, 16'd40229, 16'd31491, 16'd15569, 16'd58941, 16'd10176, 16'd33233, 16'd25536, 16'd65007, 16'd34532, 16'd16871, 16'd30112, 16'd5164, 16'd13619, 16'd37369, 16'd62584, 16'd42519, 16'd4944});
	test_expansion(128'h986a46e044898b199971ce1ecf9c46fa, {16'd61271, 16'd38645, 16'd2618, 16'd54435, 16'd5368, 16'd5127, 16'd52025, 16'd3312, 16'd35518, 16'd39492, 16'd4844, 16'd15662, 16'd58101, 16'd1218, 16'd35353, 16'd39237, 16'd26089, 16'd39539, 16'd40341, 16'd31416, 16'd8185, 16'd65406, 16'd55578, 16'd20348, 16'd53852, 16'd13162});
	test_expansion(128'h61e5eff519d1f686822e7ccf02a021ed, {16'd57293, 16'd13428, 16'd31163, 16'd28568, 16'd51602, 16'd47640, 16'd59810, 16'd47571, 16'd55247, 16'd18992, 16'd13522, 16'd16973, 16'd56604, 16'd8547, 16'd46137, 16'd15623, 16'd23286, 16'd28411, 16'd16844, 16'd31337, 16'd51069, 16'd56253, 16'd62, 16'd6622, 16'd19103, 16'd20102});
	test_expansion(128'hb203cc9f5b7163be4e014396e08f6a00, {16'd6349, 16'd48809, 16'd54908, 16'd58092, 16'd58530, 16'd34119, 16'd64749, 16'd25406, 16'd48079, 16'd1925, 16'd30970, 16'd42153, 16'd39272, 16'd47034, 16'd32461, 16'd15824, 16'd45988, 16'd7145, 16'd44361, 16'd7690, 16'd8440, 16'd62941, 16'd54260, 16'd1490, 16'd19239, 16'd29935});
	test_expansion(128'hf780f2f07b55cef46855672010f14d27, {16'd37331, 16'd54873, 16'd13010, 16'd6318, 16'd53152, 16'd7530, 16'd20450, 16'd42337, 16'd34575, 16'd43707, 16'd43160, 16'd10574, 16'd3136, 16'd13280, 16'd7272, 16'd24496, 16'd63111, 16'd27292, 16'd53088, 16'd38120, 16'd12879, 16'd41072, 16'd866, 16'd5672, 16'd11036, 16'd1306});
	test_expansion(128'h3ad52222bf006c40bcc27319992f526c, {16'd51431, 16'd53829, 16'd27688, 16'd51691, 16'd28160, 16'd45592, 16'd58879, 16'd58816, 16'd32343, 16'd18435, 16'd2072, 16'd43669, 16'd7629, 16'd8765, 16'd62673, 16'd39685, 16'd29675, 16'd44969, 16'd15606, 16'd34929, 16'd25588, 16'd40461, 16'd39703, 16'd31876, 16'd1050, 16'd4957});
	test_expansion(128'h7b2439016181b11dc103afbb15387cd4, {16'd45648, 16'd8099, 16'd22018, 16'd8616, 16'd35373, 16'd14341, 16'd12527, 16'd13987, 16'd199, 16'd36967, 16'd54174, 16'd61441, 16'd14680, 16'd32591, 16'd11684, 16'd21896, 16'd33226, 16'd34812, 16'd7194, 16'd16873, 16'd56445, 16'd48606, 16'd2090, 16'd3270, 16'd61907, 16'd48657});
	test_expansion(128'h0afbe91f0d538e2fecf15f212f6f1014, {16'd15713, 16'd54275, 16'd25059, 16'd29406, 16'd46085, 16'd60302, 16'd40672, 16'd6593, 16'd7615, 16'd62409, 16'd57557, 16'd24904, 16'd43487, 16'd23652, 16'd15289, 16'd6818, 16'd49759, 16'd51178, 16'd6826, 16'd17061, 16'd48429, 16'd50512, 16'd53623, 16'd40389, 16'd16148, 16'd28248});
	test_expansion(128'hafa413e7fabf5925d71ba1eea401601f, {16'd45669, 16'd7836, 16'd55706, 16'd28637, 16'd22219, 16'd53695, 16'd16820, 16'd55029, 16'd30296, 16'd58545, 16'd8312, 16'd3564, 16'd29501, 16'd29971, 16'd16611, 16'd37795, 16'd49771, 16'd37000, 16'd9345, 16'd3849, 16'd52539, 16'd21426, 16'd59900, 16'd58520, 16'd10421, 16'd3319});
	test_expansion(128'ha20b0ed1e649719d7388244f08b56c38, {16'd3133, 16'd30914, 16'd24036, 16'd60283, 16'd12770, 16'd17522, 16'd49394, 16'd53811, 16'd26507, 16'd63800, 16'd704, 16'd58648, 16'd16047, 16'd48231, 16'd52131, 16'd17222, 16'd57904, 16'd6415, 16'd14161, 16'd27815, 16'd24296, 16'd32913, 16'd47094, 16'd662, 16'd54625, 16'd45547});
	test_expansion(128'h7aadd7d4ee587b70086641c8fde3cc47, {16'd27791, 16'd17835, 16'd65377, 16'd45081, 16'd19242, 16'd15131, 16'd49871, 16'd48190, 16'd26754, 16'd57962, 16'd33170, 16'd63284, 16'd18880, 16'd44158, 16'd58344, 16'd34700, 16'd10615, 16'd20358, 16'd30600, 16'd21230, 16'd62921, 16'd25005, 16'd23973, 16'd27044, 16'd7325, 16'd7258});
	test_expansion(128'hee3c53c4c628628dffdb32edc9d3e488, {16'd32715, 16'd34099, 16'd27236, 16'd40688, 16'd50562, 16'd58085, 16'd27631, 16'd40150, 16'd11491, 16'd29189, 16'd18962, 16'd18168, 16'd58342, 16'd34593, 16'd10538, 16'd7806, 16'd43285, 16'd33940, 16'd33937, 16'd2234, 16'd19423, 16'd42243, 16'd1624, 16'd14184, 16'd3664, 16'd22631});
	test_expansion(128'h54a5bd7211acb651b7ae145e7cb360a8, {16'd50726, 16'd38665, 16'd42239, 16'd25101, 16'd34859, 16'd26082, 16'd10346, 16'd46868, 16'd63117, 16'd47561, 16'd44411, 16'd61015, 16'd45447, 16'd35005, 16'd9586, 16'd22005, 16'd55356, 16'd19102, 16'd19509, 16'd50778, 16'd26028, 16'd3174, 16'd49707, 16'd12006, 16'd11650, 16'd31770});
	test_expansion(128'hd1601e0c2891052d5878b1e29fbf0303, {16'd30751, 16'd40507, 16'd15233, 16'd17232, 16'd7930, 16'd32231, 16'd62037, 16'd64655, 16'd696, 16'd24551, 16'd23496, 16'd55158, 16'd12360, 16'd35241, 16'd17682, 16'd29990, 16'd58666, 16'd24051, 16'd33906, 16'd34734, 16'd29175, 16'd26452, 16'd65248, 16'd32213, 16'd35272, 16'd55198});
	test_expansion(128'h5bc4fe809964432268c7570d7f888f7e, {16'd54567, 16'd26015, 16'd30175, 16'd1181, 16'd18066, 16'd7691, 16'd36760, 16'd26955, 16'd41734, 16'd43773, 16'd8840, 16'd23647, 16'd33861, 16'd25751, 16'd2259, 16'd48015, 16'd60272, 16'd25371, 16'd21263, 16'd27281, 16'd49391, 16'd16751, 16'd30550, 16'd2944, 16'd41953, 16'd11215});
	test_expansion(128'hcd6f2834dfefb5a7c89d4bbd966344cb, {16'd44468, 16'd23907, 16'd60824, 16'd23043, 16'd44329, 16'd63514, 16'd6663, 16'd23798, 16'd51582, 16'd46971, 16'd18244, 16'd61221, 16'd62497, 16'd8190, 16'd46109, 16'd58630, 16'd33101, 16'd15481, 16'd35646, 16'd30852, 16'd54763, 16'd54701, 16'd6882, 16'd54044, 16'd42085, 16'd34929});
	test_expansion(128'h588b018a98d458406a58e7652648c8e3, {16'd17220, 16'd44196, 16'd64343, 16'd19146, 16'd59811, 16'd642, 16'd57960, 16'd45346, 16'd2569, 16'd9256, 16'd35484, 16'd40036, 16'd63883, 16'd16280, 16'd11239, 16'd51213, 16'd7347, 16'd45094, 16'd21456, 16'd44598, 16'd10693, 16'd63285, 16'd42784, 16'd55253, 16'd22623, 16'd8774});
	test_expansion(128'h62b2dd4b37d175588aade2094f527d9b, {16'd23876, 16'd39741, 16'd14068, 16'd59779, 16'd16992, 16'd5503, 16'd61622, 16'd22805, 16'd37328, 16'd9019, 16'd26044, 16'd61234, 16'd19975, 16'd10334, 16'd47445, 16'd41356, 16'd23309, 16'd22168, 16'd54962, 16'd1602, 16'd4775, 16'd15876, 16'd30350, 16'd24619, 16'd16982, 16'd9318});
	test_expansion(128'hf0f881112b9ad2e41da3b2e47d23c11c, {16'd61379, 16'd33179, 16'd16064, 16'd48704, 16'd30800, 16'd29235, 16'd40139, 16'd1569, 16'd61251, 16'd56761, 16'd44417, 16'd30612, 16'd57369, 16'd24617, 16'd40168, 16'd19443, 16'd37044, 16'd62973, 16'd17781, 16'd2145, 16'd4813, 16'd55790, 16'd8790, 16'd18001, 16'd14165, 16'd18499});
	test_expansion(128'h27cbece21975080ffc29bf8afbd7ee48, {16'd55105, 16'd31949, 16'd5557, 16'd55507, 16'd702, 16'd16251, 16'd60650, 16'd53741, 16'd58358, 16'd34912, 16'd25242, 16'd57717, 16'd55940, 16'd31770, 16'd5974, 16'd33017, 16'd36534, 16'd2862, 16'd19245, 16'd16364, 16'd47757, 16'd54847, 16'd17408, 16'd40550, 16'd40290, 16'd37970});
	test_expansion(128'hebde4b1159fec9a7ed4dfc379ec347a8, {16'd38801, 16'd31515, 16'd1417, 16'd19808, 16'd51702, 16'd15274, 16'd31202, 16'd55647, 16'd43067, 16'd26257, 16'd13812, 16'd8684, 16'd52245, 16'd55536, 16'd34993, 16'd3549, 16'd8454, 16'd9438, 16'd11426, 16'd58757, 16'd11537, 16'd61543, 16'd63632, 16'd60889, 16'd58793, 16'd48754});
	test_expansion(128'h4fbca04a22e222d0455569da8594fc7b, {16'd59540, 16'd26877, 16'd21161, 16'd44487, 16'd49900, 16'd17856, 16'd35109, 16'd25219, 16'd36083, 16'd18576, 16'd12956, 16'd29208, 16'd27782, 16'd48302, 16'd54509, 16'd13365, 16'd13431, 16'd21477, 16'd13239, 16'd34574, 16'd32177, 16'd1879, 16'd59358, 16'd9117, 16'd55869, 16'd53192});
	test_expansion(128'h30c8d36f7f3ae25c74bcad248e2fac84, {16'd17607, 16'd58245, 16'd45876, 16'd35023, 16'd55743, 16'd7619, 16'd25991, 16'd58941, 16'd62455, 16'd17065, 16'd24076, 16'd1288, 16'd48065, 16'd5825, 16'd4498, 16'd116, 16'd800, 16'd63676, 16'd59756, 16'd2307, 16'd25174, 16'd13677, 16'd27084, 16'd55781, 16'd45629, 16'd18779});
	test_expansion(128'ha573e60fb933f53ad4a658d8c13d207d, {16'd46063, 16'd15891, 16'd20356, 16'd6231, 16'd14574, 16'd9342, 16'd56046, 16'd33458, 16'd46237, 16'd7710, 16'd58645, 16'd13731, 16'd45643, 16'd10228, 16'd62093, 16'd47703, 16'd60334, 16'd32982, 16'd61448, 16'd16076, 16'd46866, 16'd47242, 16'd43393, 16'd14243, 16'd33887, 16'd50748});
	test_expansion(128'ha5bf4c9f78076cba08054a9f61db31e8, {16'd56021, 16'd3018, 16'd63969, 16'd57443, 16'd60771, 16'd63906, 16'd47909, 16'd64182, 16'd27562, 16'd869, 16'd44554, 16'd14982, 16'd29558, 16'd59364, 16'd2644, 16'd36597, 16'd46621, 16'd46840, 16'd61304, 16'd32240, 16'd38937, 16'd8384, 16'd15031, 16'd6035, 16'd16800, 16'd35667});
	test_expansion(128'ha6d89bf59ae750ee67ea88ac2e6e36f5, {16'd33233, 16'd16636, 16'd8630, 16'd63175, 16'd24609, 16'd31921, 16'd53016, 16'd56539, 16'd45599, 16'd308, 16'd55338, 16'd10647, 16'd13786, 16'd16338, 16'd28819, 16'd37665, 16'd40664, 16'd22906, 16'd44628, 16'd5780, 16'd9504, 16'd25542, 16'd50072, 16'd20783, 16'd52909, 16'd41640});
	test_expansion(128'hd091e6853e3f788998529ab2bdfa2806, {16'd18027, 16'd39864, 16'd44029, 16'd42028, 16'd50680, 16'd50670, 16'd1615, 16'd18606, 16'd58031, 16'd45040, 16'd39052, 16'd43181, 16'd22613, 16'd45246, 16'd59532, 16'd52497, 16'd17775, 16'd59243, 16'd38034, 16'd19897, 16'd40264, 16'd61507, 16'd45805, 16'd9731, 16'd30502, 16'd36890});
	test_expansion(128'he61909275da3ac2454885cd921522b25, {16'd57274, 16'd12177, 16'd50334, 16'd8862, 16'd31709, 16'd37322, 16'd54168, 16'd34734, 16'd65262, 16'd56245, 16'd6953, 16'd2944, 16'd476, 16'd30387, 16'd13578, 16'd34587, 16'd58247, 16'd19238, 16'd11538, 16'd13771, 16'd26078, 16'd5250, 16'd13556, 16'd49892, 16'd5686, 16'd7356});
	test_expansion(128'he8d922d2c4580d39d62340e11f3cffcd, {16'd23283, 16'd28640, 16'd29993, 16'd9955, 16'd62294, 16'd37197, 16'd41803, 16'd45959, 16'd27915, 16'd3733, 16'd13415, 16'd35002, 16'd16379, 16'd8141, 16'd64977, 16'd13935, 16'd59028, 16'd51373, 16'd33110, 16'd5236, 16'd57348, 16'd62166, 16'd16017, 16'd3868, 16'd49868, 16'd36954});
	test_expansion(128'hdf758a7c7b9b17c204a63932d60eb361, {16'd41174, 16'd28266, 16'd29571, 16'd12313, 16'd30212, 16'd21026, 16'd39614, 16'd21507, 16'd42425, 16'd16093, 16'd44421, 16'd10017, 16'd13595, 16'd40610, 16'd13602, 16'd24452, 16'd43883, 16'd44634, 16'd30856, 16'd16939, 16'd38331, 16'd11698, 16'd11765, 16'd47303, 16'd28238, 16'd33641});
	test_expansion(128'hc3073ddc3aef16483636aaed7f4b3edb, {16'd530, 16'd32044, 16'd23302, 16'd40476, 16'd59377, 16'd58679, 16'd4492, 16'd46905, 16'd53713, 16'd3439, 16'd41830, 16'd15279, 16'd477, 16'd32217, 16'd33522, 16'd19224, 16'd34612, 16'd13705, 16'd1729, 16'd63330, 16'd53874, 16'd31301, 16'd63413, 16'd32775, 16'd7957, 16'd11975});
	test_expansion(128'h3e48f695ff79cc845467f70aa64ae499, {16'd21486, 16'd56558, 16'd18865, 16'd18181, 16'd34797, 16'd31450, 16'd49972, 16'd50140, 16'd54114, 16'd55073, 16'd49656, 16'd48598, 16'd4990, 16'd51532, 16'd40878, 16'd17987, 16'd24100, 16'd36998, 16'd20837, 16'd45190, 16'd45189, 16'd31094, 16'd48533, 16'd55764, 16'd6694, 16'd20590});
	test_expansion(128'h0262b0edb2339d5992c68c4068db7965, {16'd42378, 16'd8047, 16'd8642, 16'd52420, 16'd28696, 16'd13719, 16'd9118, 16'd8714, 16'd30805, 16'd64889, 16'd17004, 16'd19116, 16'd40631, 16'd33244, 16'd41752, 16'd39938, 16'd5907, 16'd55985, 16'd57757, 16'd40838, 16'd48934, 16'd5690, 16'd997, 16'd5737, 16'd58335, 16'd3884});
	test_expansion(128'h667e488580b33a19ada37ccf243ad9ff, {16'd23475, 16'd53334, 16'd23512, 16'd55651, 16'd54697, 16'd54746, 16'd36121, 16'd37960, 16'd18950, 16'd37536, 16'd10915, 16'd17087, 16'd54068, 16'd60965, 16'd45297, 16'd19081, 16'd53225, 16'd39768, 16'd12960, 16'd65529, 16'd41643, 16'd52058, 16'd7941, 16'd8149, 16'd44598, 16'd46838});
	test_expansion(128'h218ace6dee1bb0feae5fdba439d7cd85, {16'd29682, 16'd4756, 16'd21411, 16'd59306, 16'd33670, 16'd15646, 16'd62044, 16'd16118, 16'd22798, 16'd17045, 16'd5247, 16'd43536, 16'd22851, 16'd48429, 16'd2315, 16'd14565, 16'd12533, 16'd6897, 16'd4060, 16'd37030, 16'd29402, 16'd49281, 16'd64102, 16'd34351, 16'd55549, 16'd18397});
	test_expansion(128'h0de319df35dfedb6c1644036ba7a623d, {16'd24279, 16'd15168, 16'd13134, 16'd32409, 16'd51128, 16'd50837, 16'd2320, 16'd63193, 16'd2539, 16'd16912, 16'd14741, 16'd33806, 16'd31043, 16'd17683, 16'd32879, 16'd50224, 16'd24358, 16'd53899, 16'd31339, 16'd8039, 16'd39184, 16'd56688, 16'd4223, 16'd56139, 16'd55713, 16'd24263});
	test_expansion(128'h87bcdfda53ab9fd987477c7ae1e135e8, {16'd63977, 16'd27345, 16'd45301, 16'd6095, 16'd37877, 16'd22254, 16'd57095, 16'd56134, 16'd63834, 16'd3991, 16'd13554, 16'd39899, 16'd30761, 16'd14357, 16'd9840, 16'd26548, 16'd14554, 16'd4305, 16'd28581, 16'd44953, 16'd25327, 16'd45538, 16'd52675, 16'd43964, 16'd809, 16'd8455});
	test_expansion(128'h59aaba32ae87f0f8a2b0bf13082d979a, {16'd9804, 16'd23863, 16'd48236, 16'd24552, 16'd60395, 16'd50925, 16'd61957, 16'd22633, 16'd9518, 16'd12512, 16'd62078, 16'd48967, 16'd12175, 16'd11142, 16'd59988, 16'd13347, 16'd62271, 16'd55914, 16'd5591, 16'd12687, 16'd33812, 16'd26008, 16'd27248, 16'd39653, 16'd30357, 16'd167});
	test_expansion(128'hbeaee838aaf6d31fd5a9a1520a539e77, {16'd1434, 16'd26050, 16'd48178, 16'd15184, 16'd25277, 16'd61119, 16'd36451, 16'd28730, 16'd30127, 16'd55124, 16'd16516, 16'd12051, 16'd10149, 16'd51757, 16'd21510, 16'd40103, 16'd56266, 16'd26878, 16'd1416, 16'd16212, 16'd31072, 16'd3213, 16'd24228, 16'd62314, 16'd59578, 16'd45141});
	test_expansion(128'h009416fd0b8aaf5afaa19ca8320d3f70, {16'd46020, 16'd26164, 16'd9776, 16'd29110, 16'd11, 16'd35252, 16'd48656, 16'd33891, 16'd23838, 16'd59164, 16'd13894, 16'd8829, 16'd64278, 16'd7784, 16'd51696, 16'd21682, 16'd45365, 16'd35134, 16'd35302, 16'd34241, 16'd44801, 16'd51415, 16'd33630, 16'd19727, 16'd61164, 16'd7181});
	test_expansion(128'h0ab81d60b76743f9b18196fc15de9334, {16'd19761, 16'd50816, 16'd10306, 16'd14162, 16'd62706, 16'd25011, 16'd32891, 16'd32942, 16'd6655, 16'd64778, 16'd43009, 16'd56462, 16'd23750, 16'd58648, 16'd33371, 16'd61166, 16'd11072, 16'd16472, 16'd35696, 16'd767, 16'd6634, 16'd40490, 16'd31979, 16'd43856, 16'd22233, 16'd18773});
	test_expansion(128'ha90dcd6b8153a5fd930d37c627d5842f, {16'd28527, 16'd35641, 16'd43390, 16'd57673, 16'd40991, 16'd55539, 16'd13554, 16'd26010, 16'd63222, 16'd4125, 16'd57786, 16'd5030, 16'd32029, 16'd65534, 16'd35266, 16'd30010, 16'd17055, 16'd10610, 16'd8473, 16'd48112, 16'd26770, 16'd45004, 16'd59279, 16'd28432, 16'd10907, 16'd14903});
	test_expansion(128'hb7e93ac540a0969a56564a5fa9cbeaa9, {16'd41961, 16'd58585, 16'd31278, 16'd15705, 16'd6827, 16'd53149, 16'd47379, 16'd24706, 16'd37137, 16'd34784, 16'd48916, 16'd45208, 16'd50094, 16'd31711, 16'd59869, 16'd23655, 16'd23853, 16'd64865, 16'd11915, 16'd20411, 16'd7575, 16'd6637, 16'd5670, 16'd58645, 16'd54100, 16'd34798});
	test_expansion(128'h88706103caf6d9fb939a747202b7e383, {16'd24264, 16'd60518, 16'd52768, 16'd24998, 16'd29985, 16'd46756, 16'd56812, 16'd52612, 16'd13987, 16'd33978, 16'd14821, 16'd36588, 16'd7543, 16'd31015, 16'd9539, 16'd57488, 16'd7059, 16'd3958, 16'd29529, 16'd35970, 16'd47819, 16'd4824, 16'd21989, 16'd59413, 16'd47769, 16'd1959});
	test_expansion(128'h04fe561eca09f425daee1b4ee440d6a3, {16'd6387, 16'd3946, 16'd8796, 16'd17491, 16'd41247, 16'd63308, 16'd51508, 16'd1735, 16'd5589, 16'd20514, 16'd38868, 16'd37434, 16'd30045, 16'd44716, 16'd46802, 16'd18690, 16'd19426, 16'd37411, 16'd42170, 16'd8265, 16'd40556, 16'd7917, 16'd50693, 16'd9885, 16'd43434, 16'd27611});
	test_expansion(128'ha8d7a8235c761734d67c4bc540cc5091, {16'd15089, 16'd11704, 16'd2470, 16'd15177, 16'd4096, 16'd50946, 16'd59840, 16'd12951, 16'd12902, 16'd57544, 16'd60880, 16'd31092, 16'd8674, 16'd7116, 16'd38956, 16'd2128, 16'd19847, 16'd27581, 16'd50350, 16'd62700, 16'd238, 16'd13370, 16'd20686, 16'd64509, 16'd6594, 16'd65165});
	test_expansion(128'hf9a3c094966b03c394192531e0e23807, {16'd8201, 16'd48194, 16'd2553, 16'd35664, 16'd39561, 16'd17748, 16'd56248, 16'd28880, 16'd46908, 16'd26508, 16'd60930, 16'd20158, 16'd50819, 16'd10995, 16'd45626, 16'd15782, 16'd49826, 16'd53534, 16'd64752, 16'd7477, 16'd30481, 16'd46874, 16'd57259, 16'd34113, 16'd29210, 16'd51380});
	test_expansion(128'h3992a2ac23d11bf8be4cf21785d7e873, {16'd6950, 16'd42369, 16'd17841, 16'd53718, 16'd63661, 16'd23773, 16'd64053, 16'd48903, 16'd26718, 16'd53823, 16'd6743, 16'd14107, 16'd33605, 16'd17573, 16'd41342, 16'd19032, 16'd47159, 16'd42226, 16'd16194, 16'd16523, 16'd33048, 16'd22367, 16'd64997, 16'd26477, 16'd54671, 16'd62819});
	test_expansion(128'ha04b9ac62679699511093973610a3a93, {16'd6548, 16'd27213, 16'd11408, 16'd47077, 16'd38356, 16'd39466, 16'd19047, 16'd12817, 16'd10052, 16'd57803, 16'd2833, 16'd40723, 16'd55838, 16'd18816, 16'd3070, 16'd42882, 16'd26453, 16'd28611, 16'd61918, 16'd57246, 16'd1485, 16'd20155, 16'd52277, 16'd34154, 16'd2326, 16'd20939});
	test_expansion(128'h03dc8ae5c3cffb597b3b0614aedc42c5, {16'd43081, 16'd60593, 16'd3883, 16'd53350, 16'd54704, 16'd3451, 16'd13470, 16'd1005, 16'd12693, 16'd1062, 16'd34961, 16'd4135, 16'd13940, 16'd1669, 16'd48663, 16'd41099, 16'd45894, 16'd37954, 16'd14923, 16'd42516, 16'd47126, 16'd47105, 16'd29905, 16'd21940, 16'd51598, 16'd59056});
	test_expansion(128'h8840dba5f78f1c0f7d12a5398bc5823c, {16'd19449, 16'd48554, 16'd32905, 16'd25709, 16'd5160, 16'd34261, 16'd43836, 16'd48749, 16'd54044, 16'd64530, 16'd47081, 16'd1648, 16'd63767, 16'd32709, 16'd37795, 16'd25461, 16'd42481, 16'd35604, 16'd44713, 16'd30529, 16'd22866, 16'd12294, 16'd27641, 16'd2920, 16'd47006, 16'd21252});
	test_expansion(128'h5ec0f6b9ac7c95a626cea90b8b53ef6c, {16'd32352, 16'd11868, 16'd62734, 16'd4329, 16'd46696, 16'd8022, 16'd59936, 16'd44425, 16'd41228, 16'd63911, 16'd49678, 16'd20890, 16'd16419, 16'd40892, 16'd58956, 16'd12865, 16'd25002, 16'd36713, 16'd17393, 16'd61447, 16'd8539, 16'd241, 16'd22959, 16'd37782, 16'd62136, 16'd27988});
	test_expansion(128'hd182e29ac4c031477763af95652b40d4, {16'd20428, 16'd42850, 16'd56510, 16'd14444, 16'd7160, 16'd26044, 16'd3413, 16'd325, 16'd43, 16'd10925, 16'd6853, 16'd2252, 16'd16438, 16'd34345, 16'd62848, 16'd58979, 16'd49225, 16'd7942, 16'd24102, 16'd57929, 16'd45420, 16'd22399, 16'd22860, 16'd28038, 16'd7588, 16'd13102});
	test_expansion(128'ha2069c4cc5ccd62080880d7317d1e6ba, {16'd5597, 16'd50162, 16'd28047, 16'd20638, 16'd47305, 16'd62957, 16'd37928, 16'd64531, 16'd24049, 16'd23995, 16'd56924, 16'd27541, 16'd40122, 16'd53853, 16'd40543, 16'd36703, 16'd63145, 16'd37250, 16'd41182, 16'd13518, 16'd1975, 16'd24364, 16'd64640, 16'd49342, 16'd1595, 16'd64450});
	test_expansion(128'ha07f44303acbb26349d3385843a06b67, {16'd15946, 16'd3379, 16'd56724, 16'd31870, 16'd33349, 16'd37054, 16'd4298, 16'd46651, 16'd47653, 16'd4464, 16'd27879, 16'd32431, 16'd42285, 16'd48612, 16'd2303, 16'd64653, 16'd38271, 16'd58976, 16'd59173, 16'd29027, 16'd26746, 16'd37993, 16'd17793, 16'd44964, 16'd11406, 16'd14373});
	test_expansion(128'hd0cc56050539e9a388a9f81fec42017a, {16'd41653, 16'd16028, 16'd45226, 16'd47415, 16'd5921, 16'd58796, 16'd6786, 16'd14383, 16'd49410, 16'd15468, 16'd11731, 16'd43859, 16'd65221, 16'd1051, 16'd43453, 16'd10542, 16'd4393, 16'd51577, 16'd15123, 16'd17999, 16'd18401, 16'd28930, 16'd40114, 16'd23092, 16'd52755, 16'd41316});
	test_expansion(128'h6c33c2d1fee356f6b6f571091d7b84a3, {16'd14474, 16'd62910, 16'd51305, 16'd16468, 16'd23448, 16'd9088, 16'd35468, 16'd46541, 16'd18900, 16'd56876, 16'd19983, 16'd53298, 16'd49709, 16'd47505, 16'd54051, 16'd63374, 16'd39556, 16'd1868, 16'd49075, 16'd2681, 16'd58755, 16'd50308, 16'd37607, 16'd9964, 16'd1095, 16'd44227});
	test_expansion(128'he17807e6a96bb3faec8e6c587f2d8748, {16'd5112, 16'd44260, 16'd18836, 16'd3024, 16'd13453, 16'd47583, 16'd20953, 16'd46258, 16'd43118, 16'd41243, 16'd18263, 16'd46718, 16'd6808, 16'd25821, 16'd51791, 16'd53109, 16'd12863, 16'd10448, 16'd52641, 16'd21158, 16'd44843, 16'd4072, 16'd46583, 16'd4671, 16'd32470, 16'd26782});
	test_expansion(128'hdaa4adce14937a3cd20a250bebd8f657, {16'd29806, 16'd46586, 16'd36892, 16'd41456, 16'd28446, 16'd56901, 16'd53175, 16'd52373, 16'd38279, 16'd44332, 16'd22878, 16'd22816, 16'd50794, 16'd52833, 16'd23113, 16'd33910, 16'd2844, 16'd15708, 16'd45115, 16'd57205, 16'd24130, 16'd30712, 16'd31815, 16'd51647, 16'd22210, 16'd12636});
	test_expansion(128'h8120615a47f8766d84b0460274ffa1b6, {16'd61398, 16'd20786, 16'd40736, 16'd3970, 16'd29660, 16'd4077, 16'd19593, 16'd23663, 16'd21849, 16'd17160, 16'd35682, 16'd63090, 16'd46655, 16'd39920, 16'd5149, 16'd20923, 16'd28949, 16'd1841, 16'd19451, 16'd10478, 16'd34850, 16'd17754, 16'd52588, 16'd36796, 16'd47687, 16'd25876});
	test_expansion(128'h86592bfb70ac2811979489f188fee32f, {16'd30315, 16'd12407, 16'd60388, 16'd33054, 16'd5109, 16'd58275, 16'd64338, 16'd17929, 16'd60214, 16'd42510, 16'd4507, 16'd57042, 16'd25919, 16'd11314, 16'd62626, 16'd36219, 16'd36747, 16'd61143, 16'd59184, 16'd27118, 16'd45366, 16'd5422, 16'd21144, 16'd37311, 16'd647, 16'd28757});
	test_expansion(128'h987c35db6e49983f91a941e64449815a, {16'd57919, 16'd51391, 16'd36685, 16'd11707, 16'd16759, 16'd31055, 16'd50129, 16'd22779, 16'd9526, 16'd58699, 16'd36065, 16'd10613, 16'd31368, 16'd45169, 16'd5135, 16'd18733, 16'd40046, 16'd52583, 16'd2502, 16'd32930, 16'd28240, 16'd52161, 16'd19419, 16'd53855, 16'd52677, 16'd26980});
	test_expansion(128'h79d9dd2d7c0eddc3f44d70d7aabc10b0, {16'd59123, 16'd52106, 16'd4527, 16'd32527, 16'd56367, 16'd3846, 16'd24571, 16'd3644, 16'd64702, 16'd49909, 16'd9313, 16'd56619, 16'd36855, 16'd58539, 16'd63306, 16'd52182, 16'd46356, 16'd59268, 16'd61324, 16'd32723, 16'd10059, 16'd37005, 16'd24797, 16'd48308, 16'd33749, 16'd41148});
	test_expansion(128'h7fa0a7df4110aa45dd6a1a3692c3fcb7, {16'd9084, 16'd24976, 16'd8962, 16'd24483, 16'd25415, 16'd53287, 16'd34015, 16'd26061, 16'd50655, 16'd60006, 16'd33260, 16'd49981, 16'd19523, 16'd15727, 16'd21980, 16'd6784, 16'd21974, 16'd18878, 16'd16042, 16'd46592, 16'd35425, 16'd59467, 16'd30980, 16'd60491, 16'd58074, 16'd56357});
	test_expansion(128'ha781717d23f30d577bc218bc807f37a3, {16'd63631, 16'd13360, 16'd59777, 16'd29782, 16'd25323, 16'd56589, 16'd52333, 16'd39719, 16'd35447, 16'd17033, 16'd37102, 16'd25549, 16'd48345, 16'd58066, 16'd27483, 16'd62315, 16'd10296, 16'd47859, 16'd35338, 16'd63194, 16'd3519, 16'd59541, 16'd50020, 16'd6367, 16'd22174, 16'd30479});
	test_expansion(128'h7dbf0c06025d157d44a871e2f335eed2, {16'd53579, 16'd58332, 16'd3289, 16'd56606, 16'd13762, 16'd52707, 16'd26284, 16'd52471, 16'd34411, 16'd62874, 16'd12399, 16'd45460, 16'd38580, 16'd45758, 16'd56861, 16'd3930, 16'd60307, 16'd65086, 16'd29832, 16'd54207, 16'd26995, 16'd14063, 16'd18078, 16'd48183, 16'd16711, 16'd11343});
	test_expansion(128'hec69f834d777e3ad70453b994dcc0449, {16'd51493, 16'd50509, 16'd46245, 16'd59056, 16'd6441, 16'd5533, 16'd18244, 16'd3164, 16'd9196, 16'd44588, 16'd26971, 16'd18389, 16'd64222, 16'd9545, 16'd63590, 16'd31126, 16'd6229, 16'd15034, 16'd56543, 16'd42795, 16'd59734, 16'd4293, 16'd48290, 16'd42470, 16'd19669, 16'd7781});
	test_expansion(128'hddb0ad2f05f67ac7292465dc2ea5c448, {16'd48320, 16'd60100, 16'd25588, 16'd12951, 16'd17002, 16'd54726, 16'd5435, 16'd27060, 16'd34725, 16'd42605, 16'd49915, 16'd59224, 16'd3071, 16'd57487, 16'd23170, 16'd43464, 16'd25780, 16'd21364, 16'd52219, 16'd32896, 16'd1731, 16'd43902, 16'd1679, 16'd49140, 16'd15323, 16'd44077});
	test_expansion(128'h5bf721b10cde2bd690f2df7578b2ff1f, {16'd31439, 16'd322, 16'd36530, 16'd5013, 16'd38050, 16'd45561, 16'd5076, 16'd27994, 16'd52053, 16'd42921, 16'd37688, 16'd52975, 16'd32505, 16'd10962, 16'd14999, 16'd65194, 16'd31934, 16'd4313, 16'd4455, 16'd33134, 16'd22852, 16'd39701, 16'd13114, 16'd46236, 16'd19766, 16'd4020});
	test_expansion(128'h39c9d3d77438a8874d79ef7b22de1e20, {16'd25781, 16'd29672, 16'd52055, 16'd47724, 16'd43416, 16'd16430, 16'd47683, 16'd24911, 16'd63143, 16'd40048, 16'd20836, 16'd54203, 16'd20654, 16'd53214, 16'd43791, 16'd39973, 16'd1928, 16'd43084, 16'd28238, 16'd48325, 16'd44571, 16'd19673, 16'd17334, 16'd39702, 16'd50042, 16'd60463});
	test_expansion(128'hd4bf6759a3b5ef300aa6c4a2d7d8c99b, {16'd47722, 16'd61825, 16'd2071, 16'd60158, 16'd31696, 16'd61898, 16'd45277, 16'd21820, 16'd36102, 16'd44339, 16'd22606, 16'd23295, 16'd44033, 16'd20845, 16'd12131, 16'd34207, 16'd49644, 16'd56768, 16'd670, 16'd18548, 16'd41110, 16'd33811, 16'd15656, 16'd44609, 16'd35065, 16'd20985});
	test_expansion(128'h7ebcdbfcc7fa1c73a416c9f50f4a0e35, {16'd51244, 16'd32344, 16'd61114, 16'd42908, 16'd27658, 16'd50406, 16'd61660, 16'd34111, 16'd33143, 16'd40523, 16'd22228, 16'd53062, 16'd55050, 16'd45016, 16'd11961, 16'd42520, 16'd41111, 16'd43156, 16'd1883, 16'd37133, 16'd53612, 16'd5437, 16'd5860, 16'd1569, 16'd14503, 16'd25457});
	test_expansion(128'hac54a6a9087338be7723e9f3d0bc15d0, {16'd48156, 16'd45091, 16'd961, 16'd50115, 16'd11137, 16'd27238, 16'd52923, 16'd58743, 16'd62569, 16'd3220, 16'd19083, 16'd63626, 16'd16724, 16'd57692, 16'd12864, 16'd38569, 16'd18361, 16'd32123, 16'd19737, 16'd50024, 16'd51108, 16'd20570, 16'd36242, 16'd30196, 16'd54277, 16'd10538});
	test_expansion(128'haeac1d36ab27d671376e35e5d9650b2c, {16'd61561, 16'd32133, 16'd24630, 16'd45864, 16'd17283, 16'd63896, 16'd17993, 16'd25707, 16'd9383, 16'd65368, 16'd11349, 16'd49756, 16'd5093, 16'd25675, 16'd62729, 16'd41935, 16'd63439, 16'd41091, 16'd54572, 16'd9934, 16'd57288, 16'd49152, 16'd42764, 16'd32561, 16'd28981, 16'd28696});
	test_expansion(128'h3b4a2a149d45f85d3d1d3d8b3de1acc5, {16'd62744, 16'd39930, 16'd57923, 16'd54255, 16'd43254, 16'd40055, 16'd29874, 16'd52767, 16'd52278, 16'd50742, 16'd15810, 16'd32133, 16'd14834, 16'd58569, 16'd28674, 16'd41312, 16'd52184, 16'd21058, 16'd45182, 16'd12229, 16'd34010, 16'd35317, 16'd28812, 16'd17769, 16'd62096, 16'd38808});
	test_expansion(128'h2df8da0d006a4aa94d8f648cec3ac593, {16'd50586, 16'd46597, 16'd11254, 16'd24423, 16'd7611, 16'd64616, 16'd40230, 16'd54908, 16'd63325, 16'd8117, 16'd1129, 16'd55796, 16'd51992, 16'd45775, 16'd41409, 16'd43858, 16'd26525, 16'd19416, 16'd35560, 16'd41434, 16'd33281, 16'd17307, 16'd57489, 16'd28482, 16'd17865, 16'd29193});
	test_expansion(128'hcf769dce12b797daf87cd61e96510485, {16'd14655, 16'd47515, 16'd15100, 16'd39478, 16'd15840, 16'd27837, 16'd30627, 16'd52323, 16'd17213, 16'd62771, 16'd9331, 16'd41658, 16'd794, 16'd15625, 16'd25340, 16'd34426, 16'd48501, 16'd44458, 16'd37644, 16'd59836, 16'd3606, 16'd4460, 16'd56917, 16'd14626, 16'd47383, 16'd13922});
	test_expansion(128'ha8f43e7ffdd1c163cdf09e6a97c44053, {16'd2172, 16'd31755, 16'd45429, 16'd46696, 16'd28778, 16'd11638, 16'd41864, 16'd28970, 16'd21393, 16'd39353, 16'd12178, 16'd18085, 16'd2780, 16'd15853, 16'd34989, 16'd58075, 16'd18423, 16'd20562, 16'd45972, 16'd43535, 16'd2903, 16'd16448, 16'd28215, 16'd15056, 16'd23123, 16'd40916});
	test_expansion(128'h69ce0e3e8ea2c25649d1becec59e4175, {16'd16711, 16'd32510, 16'd62748, 16'd52128, 16'd4548, 16'd42610, 16'd22571, 16'd50521, 16'd51554, 16'd61185, 16'd43922, 16'd25596, 16'd28864, 16'd49080, 16'd15616, 16'd58860, 16'd35443, 16'd32675, 16'd11958, 16'd13642, 16'd8422, 16'd56400, 16'd31984, 16'd48726, 16'd19131, 16'd52152});
	test_expansion(128'h8fdf4ad7f214d9d6bbdda7a20f673ffd, {16'd363, 16'd26618, 16'd13008, 16'd4278, 16'd11637, 16'd54290, 16'd19035, 16'd680, 16'd31242, 16'd28106, 16'd2671, 16'd28554, 16'd43624, 16'd54547, 16'd59726, 16'd50888, 16'd51714, 16'd50810, 16'd42021, 16'd32741, 16'd39569, 16'd65466, 16'd21219, 16'd63204, 16'd16286, 16'd51778});
	test_expansion(128'h13a1c5867ca3d492facbcda991539033, {16'd37984, 16'd22445, 16'd16960, 16'd17869, 16'd15797, 16'd39059, 16'd56465, 16'd16984, 16'd28210, 16'd57021, 16'd9229, 16'd28852, 16'd21783, 16'd9022, 16'd47247, 16'd36707, 16'd10192, 16'd26538, 16'd11873, 16'd57723, 16'd54974, 16'd1654, 16'd56617, 16'd38707, 16'd42512, 16'd33719});
	test_expansion(128'h0d8ea5a45f13ad26297eb83ebc0c2408, {16'd59626, 16'd3828, 16'd22878, 16'd56954, 16'd22770, 16'd31481, 16'd31543, 16'd59750, 16'd47599, 16'd36002, 16'd18250, 16'd32953, 16'd24821, 16'd65104, 16'd43409, 16'd12832, 16'd42103, 16'd32598, 16'd29699, 16'd8889, 16'd55055, 16'd22935, 16'd16020, 16'd45524, 16'd6844, 16'd62702});
	test_expansion(128'h844cf788d685bd7d8240cb05f1f5e0b9, {16'd8037, 16'd40996, 16'd5368, 16'd45224, 16'd34000, 16'd61154, 16'd5443, 16'd5777, 16'd64528, 16'd65475, 16'd55175, 16'd62312, 16'd36019, 16'd13321, 16'd48930, 16'd58672, 16'd43629, 16'd27926, 16'd32688, 16'd3068, 16'd64116, 16'd7348, 16'd29244, 16'd40017, 16'd13408, 16'd18154});
	test_expansion(128'hf5c6d66bfb15d9a58f4b4f3cb84b8894, {16'd15731, 16'd7331, 16'd17408, 16'd34609, 16'd53983, 16'd14190, 16'd20798, 16'd10724, 16'd24222, 16'd61512, 16'd20012, 16'd48936, 16'd54584, 16'd61897, 16'd19579, 16'd8940, 16'd50586, 16'd22363, 16'd45177, 16'd24780, 16'd57123, 16'd43067, 16'd30199, 16'd60580, 16'd42751, 16'd39972});
	test_expansion(128'h5594ce41add402ca1a3e67aa35d5b89a, {16'd40343, 16'd61887, 16'd34364, 16'd55344, 16'd21507, 16'd45239, 16'd17062, 16'd55712, 16'd31030, 16'd25660, 16'd62844, 16'd3913, 16'd18453, 16'd19515, 16'd17465, 16'd36441, 16'd10479, 16'd6600, 16'd20450, 16'd49113, 16'd37024, 16'd7560, 16'd46392, 16'd55135, 16'd55695, 16'd32704});
	test_expansion(128'h24964932b2498155cdfbc170bb3a2365, {16'd39305, 16'd36105, 16'd51908, 16'd63382, 16'd18133, 16'd54615, 16'd23812, 16'd3611, 16'd2517, 16'd57472, 16'd24517, 16'd54493, 16'd34692, 16'd33250, 16'd41717, 16'd26658, 16'd50259, 16'd60306, 16'd38214, 16'd55028, 16'd42320, 16'd49660, 16'd61359, 16'd5978, 16'd52708, 16'd58547});
	test_expansion(128'hd458f885c218da7cfb863ec0c074d1f6, {16'd12175, 16'd19795, 16'd63426, 16'd27708, 16'd32351, 16'd12673, 16'd50034, 16'd5031, 16'd50116, 16'd55522, 16'd29863, 16'd53439, 16'd14377, 16'd41838, 16'd47723, 16'd53169, 16'd60243, 16'd15859, 16'd30402, 16'd1603, 16'd5732, 16'd28785, 16'd60752, 16'd44132, 16'd30027, 16'd36058});
	test_expansion(128'h177323604b731736a00010e781c787f6, {16'd1792, 16'd13461, 16'd43467, 16'd22605, 16'd53802, 16'd18972, 16'd41421, 16'd35851, 16'd25901, 16'd22093, 16'd8602, 16'd3227, 16'd25592, 16'd28679, 16'd1939, 16'd14480, 16'd12696, 16'd62276, 16'd2202, 16'd4956, 16'd41127, 16'd47782, 16'd44441, 16'd3926, 16'd32687, 16'd16212});
	test_expansion(128'h3062815cb23089b56b7f9782214c1b66, {16'd27044, 16'd14848, 16'd24025, 16'd10486, 16'd29522, 16'd7047, 16'd25116, 16'd19934, 16'd10006, 16'd5275, 16'd6328, 16'd58753, 16'd62000, 16'd17188, 16'd37631, 16'd40700, 16'd64174, 16'd22746, 16'd36405, 16'd62977, 16'd34836, 16'd65021, 16'd15873, 16'd13597, 16'd18565, 16'd40464});
	test_expansion(128'h9490ac9dcf6eaf13df9e2c0e6635a153, {16'd58937, 16'd51982, 16'd18633, 16'd1239, 16'd64940, 16'd12138, 16'd43519, 16'd33348, 16'd37116, 16'd52348, 16'd42215, 16'd9118, 16'd61220, 16'd63416, 16'd13262, 16'd29696, 16'd60210, 16'd8174, 16'd33506, 16'd61303, 16'd17830, 16'd51117, 16'd26013, 16'd54141, 16'd60876, 16'd15219});
	test_expansion(128'hdbbc620d1b28b3560721118218b1aa67, {16'd23465, 16'd34595, 16'd6754, 16'd1512, 16'd49570, 16'd16192, 16'd11436, 16'd28330, 16'd11010, 16'd47361, 16'd60000, 16'd26654, 16'd55159, 16'd46164, 16'd61705, 16'd51463, 16'd51361, 16'd36516, 16'd9342, 16'd7721, 16'd23342, 16'd9720, 16'd23861, 16'd17623, 16'd4182, 16'd56595});
	test_expansion(128'h96d98744404d953757d4cfbfecdaaa06, {16'd10809, 16'd425, 16'd17342, 16'd31503, 16'd50968, 16'd42768, 16'd19218, 16'd61151, 16'd60052, 16'd9866, 16'd49718, 16'd36724, 16'd59382, 16'd13826, 16'd1825, 16'd14253, 16'd86, 16'd25715, 16'd8637, 16'd12431, 16'd38158, 16'd26142, 16'd42741, 16'd62155, 16'd11812, 16'd28670});
	test_expansion(128'h8dc0e19d903a76024fc175fd7c69899d, {16'd8217, 16'd33248, 16'd8153, 16'd41377, 16'd30531, 16'd12302, 16'd23827, 16'd50604, 16'd22760, 16'd56807, 16'd50509, 16'd65289, 16'd38513, 16'd14304, 16'd41661, 16'd19185, 16'd25971, 16'd26048, 16'd26730, 16'd39633, 16'd20787, 16'd54653, 16'd39534, 16'd16960, 16'd13727, 16'd64750});
	test_expansion(128'h86e30b0ef968d3e33ae8b832aea2ec81, {16'd56509, 16'd17280, 16'd29266, 16'd7061, 16'd17277, 16'd1563, 16'd55492, 16'd26076, 16'd31299, 16'd42734, 16'd42571, 16'd23620, 16'd33771, 16'd2123, 16'd48576, 16'd21890, 16'd18882, 16'd41172, 16'd28063, 16'd52438, 16'd22619, 16'd63906, 16'd28582, 16'd12221, 16'd58818, 16'd43438});
	test_expansion(128'h6c80d533cc04867d66e10c5dd155e6cd, {16'd44890, 16'd37506, 16'd44937, 16'd23710, 16'd42007, 16'd23174, 16'd13605, 16'd48342, 16'd8932, 16'd13214, 16'd22008, 16'd13649, 16'd28972, 16'd6481, 16'd22844, 16'd44717, 16'd9288, 16'd63185, 16'd38156, 16'd59916, 16'd5755, 16'd8644, 16'd30734, 16'd15711, 16'd52367, 16'd12047});
	test_expansion(128'he716f97dd52810e5dfd626567c7d7a2b, {16'd3751, 16'd45484, 16'd47848, 16'd27065, 16'd34508, 16'd38889, 16'd11430, 16'd37994, 16'd6900, 16'd4341, 16'd53568, 16'd14426, 16'd38671, 16'd363, 16'd8691, 16'd31407, 16'd63567, 16'd53199, 16'd52830, 16'd7019, 16'd57248, 16'd47667, 16'd50388, 16'd43519, 16'd51659, 16'd11619});
	test_expansion(128'hbcd453482ff6356a6405023355c33277, {16'd15366, 16'd48002, 16'd63951, 16'd28661, 16'd12571, 16'd23850, 16'd2136, 16'd1650, 16'd44126, 16'd9936, 16'd49610, 16'd61032, 16'd11439, 16'd56262, 16'd55528, 16'd25306, 16'd57561, 16'd42799, 16'd44000, 16'd48835, 16'd22913, 16'd5578, 16'd9285, 16'd60711, 16'd61699, 16'd51233});
	test_expansion(128'h5654745a7c4fc769b8150ed1c34edc7b, {16'd64372, 16'd18771, 16'd13304, 16'd23031, 16'd53734, 16'd49968, 16'd39793, 16'd51488, 16'd4826, 16'd1169, 16'd41520, 16'd6164, 16'd36246, 16'd63952, 16'd18699, 16'd60035, 16'd41492, 16'd57556, 16'd77, 16'd1363, 16'd63865, 16'd51505, 16'd32689, 16'd11726, 16'd61587, 16'd53226});
	test_expansion(128'hb5830d86c10a4d844ba2bd48a83a95eb, {16'd51941, 16'd27570, 16'd33009, 16'd56261, 16'd15711, 16'd62719, 16'd47906, 16'd60051, 16'd55159, 16'd31999, 16'd4030, 16'd53124, 16'd27511, 16'd62093, 16'd18842, 16'd39482, 16'd16834, 16'd8595, 16'd37448, 16'd27680, 16'd1274, 16'd51834, 16'd61817, 16'd65431, 16'd9600, 16'd8774});
	test_expansion(128'h27f721851e8781e6dd98b836f8fa30d0, {16'd17451, 16'd47521, 16'd48637, 16'd29737, 16'd27231, 16'd1327, 16'd29452, 16'd57150, 16'd33383, 16'd57088, 16'd60838, 16'd11560, 16'd26172, 16'd64108, 16'd28969, 16'd9669, 16'd3062, 16'd40018, 16'd42511, 16'd3414, 16'd59302, 16'd45429, 16'd33374, 16'd64263, 16'd29197, 16'd6465});
	test_expansion(128'he0ddd44e6162b8a2cedcfa91b640d374, {16'd49611, 16'd47088, 16'd34420, 16'd23672, 16'd4416, 16'd43617, 16'd47018, 16'd43969, 16'd1321, 16'd29258, 16'd36872, 16'd65135, 16'd34207, 16'd55853, 16'd61262, 16'd43042, 16'd4041, 16'd27920, 16'd41824, 16'd60468, 16'd31746, 16'd7366, 16'd32542, 16'd54157, 16'd59124, 16'd47929});
	test_expansion(128'h0a75689aa11e89cd02e4be90987a1edb, {16'd41196, 16'd11342, 16'd17849, 16'd33190, 16'd36685, 16'd40217, 16'd20728, 16'd60196, 16'd47730, 16'd4254, 16'd9501, 16'd32220, 16'd23323, 16'd25417, 16'd5860, 16'd46007, 16'd65464, 16'd49951, 16'd59621, 16'd63980, 16'd17229, 16'd51357, 16'd53867, 16'd53873, 16'd14963, 16'd29364});
	test_expansion(128'h77ae41b422b6bece5a5803517904ff07, {16'd22822, 16'd53634, 16'd29372, 16'd23122, 16'd50376, 16'd17551, 16'd43624, 16'd57887, 16'd44787, 16'd8573, 16'd27556, 16'd13048, 16'd28573, 16'd727, 16'd34419, 16'd3205, 16'd27780, 16'd58032, 16'd11448, 16'd55527, 16'd21847, 16'd13752, 16'd46820, 16'd40997, 16'd55759, 16'd26111});
	test_expansion(128'hefc76d910a87a629d296a285055af458, {16'd4393, 16'd62767, 16'd28222, 16'd6466, 16'd759, 16'd56487, 16'd10169, 16'd19369, 16'd22631, 16'd12780, 16'd26870, 16'd61354, 16'd7949, 16'd48022, 16'd24021, 16'd38291, 16'd8248, 16'd11861, 16'd56822, 16'd41061, 16'd20236, 16'd58482, 16'd3655, 16'd39667, 16'd47053, 16'd12495});
	test_expansion(128'hd1fe0b67fcab683a5743bb1470c12050, {16'd18844, 16'd42350, 16'd19453, 16'd64056, 16'd14705, 16'd64067, 16'd51819, 16'd25137, 16'd8686, 16'd27162, 16'd8022, 16'd2120, 16'd53220, 16'd14684, 16'd27649, 16'd44824, 16'd16812, 16'd3764, 16'd28079, 16'd14975, 16'd11881, 16'd34129, 16'd32920, 16'd45674, 16'd32756, 16'd48751});
	test_expansion(128'h52ffc1875404645d9908a9fe1c36a758, {16'd65283, 16'd54330, 16'd50610, 16'd58966, 16'd41555, 16'd14992, 16'd8311, 16'd54121, 16'd49513, 16'd45856, 16'd22965, 16'd19306, 16'd23450, 16'd23008, 16'd10568, 16'd61418, 16'd16864, 16'd60574, 16'd13196, 16'd47365, 16'd1862, 16'd1480, 16'd60622, 16'd64515, 16'd65125, 16'd9046});
	test_expansion(128'h8d69c82394c487711f24e8110ce34c07, {16'd39410, 16'd15825, 16'd40595, 16'd37659, 16'd49230, 16'd65499, 16'd13871, 16'd23651, 16'd12975, 16'd43244, 16'd33596, 16'd64909, 16'd5928, 16'd21461, 16'd20583, 16'd5205, 16'd60820, 16'd22943, 16'd64721, 16'd14752, 16'd9914, 16'd15730, 16'd33608, 16'd63743, 16'd2319, 16'd33224});
	test_expansion(128'h54fc18ac41be861ec7c46b0475d0f3d7, {16'd1176, 16'd30135, 16'd46614, 16'd9442, 16'd58723, 16'd30123, 16'd36541, 16'd44962, 16'd45515, 16'd25335, 16'd53947, 16'd54253, 16'd10155, 16'd58898, 16'd57016, 16'd31104, 16'd46431, 16'd49151, 16'd2936, 16'd61111, 16'd2906, 16'd27144, 16'd52679, 16'd34598, 16'd52681, 16'd24309});
	test_expansion(128'ha6b9fb5f9003db3f077df175e6952e9b, {16'd61969, 16'd43413, 16'd59770, 16'd13260, 16'd48258, 16'd26123, 16'd63107, 16'd14400, 16'd46276, 16'd22583, 16'd51484, 16'd40960, 16'd7333, 16'd51519, 16'd31468, 16'd41397, 16'd35828, 16'd32652, 16'd21692, 16'd47937, 16'd47876, 16'd22903, 16'd33022, 16'd13451, 16'd57269, 16'd30053});
	test_expansion(128'hcb2f12e35dabb84d89c716d27eb071a1, {16'd44597, 16'd58036, 16'd55341, 16'd52045, 16'd25239, 16'd37626, 16'd36916, 16'd18306, 16'd48918, 16'd19006, 16'd9545, 16'd25389, 16'd61920, 16'd20488, 16'd55427, 16'd9604, 16'd31425, 16'd50373, 16'd39890, 16'd33387, 16'd42062, 16'd35468, 16'd26653, 16'd5071, 16'd5343, 16'd42301});
	test_expansion(128'hba70bdf134bd45a778fb8e5e3f13ebf4, {16'd7710, 16'd56173, 16'd49232, 16'd36771, 16'd12307, 16'd25858, 16'd44013, 16'd13946, 16'd48813, 16'd34189, 16'd38825, 16'd26326, 16'd42871, 16'd34822, 16'd17975, 16'd2782, 16'd62175, 16'd24605, 16'd58839, 16'd33970, 16'd28522, 16'd792, 16'd14157, 16'd23250, 16'd53994, 16'd44325});
	test_expansion(128'h2598f9cc2187cec6a7e3c638f2cb9fe1, {16'd37944, 16'd8103, 16'd58035, 16'd27375, 16'd1910, 16'd38119, 16'd24402, 16'd42766, 16'd57940, 16'd39300, 16'd56168, 16'd9840, 16'd40180, 16'd31529, 16'd1993, 16'd17086, 16'd3035, 16'd9167, 16'd4596, 16'd49393, 16'd20001, 16'd13234, 16'd8235, 16'd59343, 16'd5293, 16'd20975});
	test_expansion(128'h2a2fdd17f71d690378185b3661e14837, {16'd16502, 16'd52050, 16'd60278, 16'd5745, 16'd32412, 16'd54304, 16'd43855, 16'd59679, 16'd52915, 16'd37393, 16'd34263, 16'd57893, 16'd58316, 16'd11629, 16'd63017, 16'd50333, 16'd16054, 16'd44160, 16'd34600, 16'd24471, 16'd20716, 16'd38511, 16'd36039, 16'd28215, 16'd56233, 16'd37380});
	test_expansion(128'h5cec28dfeabd3fa95c1c8fe448229698, {16'd40300, 16'd57911, 16'd50796, 16'd63301, 16'd22312, 16'd51270, 16'd18590, 16'd20923, 16'd18502, 16'd57294, 16'd21278, 16'd17111, 16'd4201, 16'd4548, 16'd14210, 16'd6349, 16'd39556, 16'd8080, 16'd57547, 16'd12216, 16'd45020, 16'd1639, 16'd59409, 16'd40022, 16'd57483, 16'd50819});
	test_expansion(128'h8228c65d8670c5dc67f1167d35495ffa, {16'd26249, 16'd60742, 16'd36678, 16'd21923, 16'd29237, 16'd1360, 16'd19612, 16'd52749, 16'd31115, 16'd50058, 16'd49967, 16'd25956, 16'd57786, 16'd61428, 16'd10057, 16'd22096, 16'd13572, 16'd30150, 16'd9364, 16'd55049, 16'd41372, 16'd49756, 16'd22049, 16'd8859, 16'd48459, 16'd64999});
	test_expansion(128'h91cc1893e1d9a8af1339b8893cf7b3d8, {16'd17633, 16'd63703, 16'd25766, 16'd55731, 16'd22242, 16'd60996, 16'd28316, 16'd50664, 16'd7857, 16'd20004, 16'd60254, 16'd55286, 16'd42348, 16'd24809, 16'd53736, 16'd28532, 16'd2993, 16'd27524, 16'd34638, 16'd46696, 16'd45612, 16'd27603, 16'd53538, 16'd10805, 16'd21612, 16'd44376});
	test_expansion(128'h95e11da45adbba01ae90db86fff7460d, {16'd63497, 16'd44077, 16'd63957, 16'd4678, 16'd5661, 16'd40288, 16'd43879, 16'd37357, 16'd8680, 16'd8304, 16'd14040, 16'd41197, 16'd7987, 16'd20965, 16'd8160, 16'd8114, 16'd45276, 16'd59593, 16'd2477, 16'd7000, 16'd10951, 16'd35163, 16'd56274, 16'd49697, 16'd44865, 16'd57166});
	test_expansion(128'h7dd1f329ab2008b80ac878f033801638, {16'd18521, 16'd33223, 16'd53887, 16'd58893, 16'd23111, 16'd22124, 16'd44955, 16'd38977, 16'd6638, 16'd34957, 16'd692, 16'd57608, 16'd50268, 16'd300, 16'd15115, 16'd57952, 16'd41338, 16'd16183, 16'd37758, 16'd57467, 16'd54768, 16'd59274, 16'd49722, 16'd16183, 16'd19578, 16'd58697});
	test_expansion(128'h2c1946603572f14afcf8bf88456c593f, {16'd19590, 16'd13101, 16'd41591, 16'd685, 16'd7183, 16'd58059, 16'd50681, 16'd40592, 16'd58630, 16'd65038, 16'd55698, 16'd14909, 16'd55123, 16'd23030, 16'd9907, 16'd61698, 16'd41797, 16'd3298, 16'd7362, 16'd1686, 16'd52346, 16'd52644, 16'd17702, 16'd58008, 16'd3238, 16'd63940});
	test_expansion(128'h9cfe2a0d94cc47c0242becf49f093fd8, {16'd50297, 16'd36144, 16'd4148, 16'd3959, 16'd51076, 16'd8347, 16'd53337, 16'd12257, 16'd25464, 16'd58688, 16'd23033, 16'd57794, 16'd21659, 16'd3471, 16'd31674, 16'd24256, 16'd56527, 16'd17520, 16'd8275, 16'd5662, 16'd27796, 16'd7095, 16'd667, 16'd59746, 16'd17407, 16'd34556});
	test_expansion(128'haa3287fa28bcd7ce544f03402827d3e8, {16'd26625, 16'd5467, 16'd53232, 16'd15215, 16'd26256, 16'd14884, 16'd59873, 16'd22021, 16'd29290, 16'd32664, 16'd10835, 16'd12991, 16'd46788, 16'd64224, 16'd17100, 16'd32478, 16'd47556, 16'd22784, 16'd48611, 16'd33642, 16'd54468, 16'd31757, 16'd22889, 16'd10489, 16'd24106, 16'd53154});
	test_expansion(128'hae11e1ea24a5a310c4dbbb10e890b16d, {16'd2283, 16'd49557, 16'd5394, 16'd6572, 16'd34207, 16'd51291, 16'd28277, 16'd31800, 16'd35547, 16'd7408, 16'd29917, 16'd39063, 16'd49108, 16'd57927, 16'd728, 16'd19986, 16'd48477, 16'd34894, 16'd37814, 16'd48726, 16'd17965, 16'd12914, 16'd31190, 16'd43750, 16'd52706, 16'd51967});
	test_expansion(128'h2d1505fcc357e55edce2bf0189e65836, {16'd36581, 16'd33611, 16'd15058, 16'd60775, 16'd55177, 16'd1631, 16'd39243, 16'd61826, 16'd13780, 16'd55842, 16'd56235, 16'd59887, 16'd22181, 16'd19020, 16'd35864, 16'd38916, 16'd28363, 16'd56716, 16'd3806, 16'd21126, 16'd6881, 16'd38646, 16'd15845, 16'd55850, 16'd5440, 16'd13069});
	test_expansion(128'h96215a8419a8eb42fd9a807a5cf4ce6a, {16'd44227, 16'd44329, 16'd10018, 16'd38445, 16'd38849, 16'd24559, 16'd48183, 16'd25744, 16'd42688, 16'd3260, 16'd27558, 16'd23593, 16'd38151, 16'd1460, 16'd52532, 16'd3357, 16'd20194, 16'd22479, 16'd5946, 16'd2387, 16'd10983, 16'd47869, 16'd58947, 16'd2189, 16'd64366, 16'd60208});
	test_expansion(128'h790ae1f99eb21e019bdf220fd28d91c3, {16'd48797, 16'd46905, 16'd4309, 16'd56955, 16'd31691, 16'd28389, 16'd21435, 16'd59706, 16'd45207, 16'd14464, 16'd24527, 16'd48795, 16'd44865, 16'd31586, 16'd39193, 16'd55652, 16'd4431, 16'd60384, 16'd26817, 16'd38684, 16'd762, 16'd58424, 16'd65447, 16'd26998, 16'd23369, 16'd58905});
	test_expansion(128'h1da6025fed28318a1f6c38f4a6be321e, {16'd23030, 16'd14418, 16'd46454, 16'd55131, 16'd31553, 16'd46312, 16'd8545, 16'd49504, 16'd58154, 16'd37256, 16'd21717, 16'd1377, 16'd7360, 16'd43620, 16'd33033, 16'd7608, 16'd3950, 16'd54997, 16'd10304, 16'd20202, 16'd30264, 16'd19165, 16'd46932, 16'd14329, 16'd11433, 16'd23086});
	test_expansion(128'h0da1cdaae577b487ad9a5343ca46844d, {16'd14740, 16'd53703, 16'd63848, 16'd15705, 16'd38316, 16'd56157, 16'd20256, 16'd31703, 16'd7050, 16'd2552, 16'd62548, 16'd51898, 16'd41043, 16'd40334, 16'd48421, 16'd9201, 16'd32654, 16'd31363, 16'd11189, 16'd57388, 16'd30202, 16'd31492, 16'd61548, 16'd40111, 16'd23202, 16'd41582});
	test_expansion(128'hdf1fbe4f183c86c85ba86e7f393b8659, {16'd64361, 16'd13658, 16'd19941, 16'd41590, 16'd48894, 16'd10029, 16'd3961, 16'd7962, 16'd62997, 16'd15564, 16'd46334, 16'd53842, 16'd24253, 16'd40158, 16'd2974, 16'd51221, 16'd142, 16'd61201, 16'd12715, 16'd51402, 16'd22873, 16'd2919, 16'd24757, 16'd3174, 16'd59376, 16'd13441});
	test_expansion(128'h485f5c6ed692ae7e87a468388dabc054, {16'd64977, 16'd387, 16'd18761, 16'd14288, 16'd36907, 16'd45993, 16'd4355, 16'd25912, 16'd48625, 16'd39023, 16'd63502, 16'd28679, 16'd12745, 16'd56640, 16'd42354, 16'd53285, 16'd64240, 16'd51031, 16'd4177, 16'd62883, 16'd25529, 16'd18978, 16'd59106, 16'd54369, 16'd8603, 16'd42063});
	test_expansion(128'h2bfa76e1f2b55a03bec04c017d7cd4fc, {16'd57490, 16'd39798, 16'd53426, 16'd53719, 16'd10522, 16'd44993, 16'd12982, 16'd39182, 16'd3606, 16'd32371, 16'd19958, 16'd53246, 16'd12446, 16'd8913, 16'd24658, 16'd39796, 16'd23652, 16'd38478, 16'd7519, 16'd59915, 16'd30316, 16'd33825, 16'd46102, 16'd56468, 16'd38909, 16'd54077});
	test_expansion(128'h7d2233744c443843ea6f80fa122a4ffd, {16'd61757, 16'd31279, 16'd52895, 16'd64901, 16'd20484, 16'd40956, 16'd6993, 16'd11258, 16'd12439, 16'd8143, 16'd50808, 16'd45741, 16'd43828, 16'd30593, 16'd52885, 16'd52070, 16'd11133, 16'd6397, 16'd29884, 16'd15077, 16'd51277, 16'd39664, 16'd50420, 16'd42133, 16'd36494, 16'd60240});
	test_expansion(128'hf6eeeaae63850c80ecdd27274463e3ab, {16'd24446, 16'd40703, 16'd59933, 16'd52580, 16'd59120, 16'd36187, 16'd64815, 16'd51950, 16'd45986, 16'd57765, 16'd6159, 16'd26389, 16'd18178, 16'd40805, 16'd21745, 16'd46346, 16'd2612, 16'd3074, 16'd3108, 16'd32482, 16'd1912, 16'd53657, 16'd60969, 16'd54117, 16'd10729, 16'd52873});
	test_expansion(128'h42dcd6db9c4e85d9ee6f143c714b6e00, {16'd2200, 16'd38383, 16'd21251, 16'd59177, 16'd35401, 16'd42551, 16'd39260, 16'd42368, 16'd3971, 16'd39123, 16'd62451, 16'd18414, 16'd10341, 16'd21542, 16'd33501, 16'd7372, 16'd33060, 16'd7440, 16'd32234, 16'd18665, 16'd62183, 16'd10659, 16'd51735, 16'd6107, 16'd51236, 16'd9468});
	test_expansion(128'h6b88f78f40587843014f5ec644fd925a, {16'd31524, 16'd31737, 16'd58891, 16'd6578, 16'd12520, 16'd43112, 16'd44990, 16'd4031, 16'd25730, 16'd12591, 16'd36222, 16'd32842, 16'd3670, 16'd54164, 16'd39592, 16'd7908, 16'd58741, 16'd57795, 16'd11814, 16'd61201, 16'd5289, 16'd54173, 16'd40698, 16'd25072, 16'd31644, 16'd36735});
	test_expansion(128'h8885d1b9fdcda6f96eac6349ccc5f40f, {16'd53956, 16'd54205, 16'd23399, 16'd20672, 16'd54429, 16'd25520, 16'd44814, 16'd7679, 16'd4848, 16'd4031, 16'd5357, 16'd11300, 16'd29666, 16'd11200, 16'd12326, 16'd38452, 16'd49448, 16'd35463, 16'd49320, 16'd33849, 16'd46462, 16'd53911, 16'd22646, 16'd14480, 16'd19367, 16'd10187});
	test_expansion(128'he71733c281342a6019ea706dbc4660d3, {16'd26145, 16'd20901, 16'd20777, 16'd12673, 16'd55619, 16'd9985, 16'd9111, 16'd29, 16'd19824, 16'd45624, 16'd19625, 16'd62658, 16'd63952, 16'd6182, 16'd60637, 16'd42065, 16'd52833, 16'd23137, 16'd40509, 16'd29479, 16'd3077, 16'd19777, 16'd47140, 16'd14023, 16'd36525, 16'd54775});
	test_expansion(128'hcf105ff09ff362a2503961a3d0851ba8, {16'd34512, 16'd52421, 16'd30403, 16'd1799, 16'd26579, 16'd56559, 16'd64115, 16'd60973, 16'd44476, 16'd44838, 16'd21581, 16'd17925, 16'd61613, 16'd64435, 16'd48720, 16'd1550, 16'd33507, 16'd1920, 16'd14671, 16'd38427, 16'd8356, 16'd31386, 16'd56794, 16'd42287, 16'd31078, 16'd43582});
	test_expansion(128'hde1471391999d740d9fd4406b8feab1c, {16'd22435, 16'd28831, 16'd40186, 16'd9009, 16'd57896, 16'd10752, 16'd51958, 16'd44711, 16'd19322, 16'd57495, 16'd54972, 16'd6886, 16'd53753, 16'd3702, 16'd49780, 16'd10658, 16'd41129, 16'd51400, 16'd22240, 16'd18594, 16'd31064, 16'd13877, 16'd26862, 16'd31023, 16'd60231, 16'd63150});
	test_expansion(128'h49c559f0672b11bf82e5f6adecb6c130, {16'd47260, 16'd30923, 16'd5505, 16'd21850, 16'd43668, 16'd57986, 16'd52885, 16'd59924, 16'd64402, 16'd27803, 16'd33849, 16'd44858, 16'd20018, 16'd3038, 16'd11284, 16'd19430, 16'd42357, 16'd47853, 16'd8782, 16'd16492, 16'd56832, 16'd46573, 16'd10568, 16'd7002, 16'd3996, 16'd64994});
	test_expansion(128'hcd5ff015a27ce766a2edcaa341a2efe9, {16'd60979, 16'd65338, 16'd26020, 16'd12035, 16'd7547, 16'd63057, 16'd28999, 16'd37814, 16'd3632, 16'd19624, 16'd20460, 16'd10691, 16'd60334, 16'd25647, 16'd18844, 16'd13862, 16'd54451, 16'd55573, 16'd60335, 16'd48656, 16'd14559, 16'd10275, 16'd64020, 16'd29244, 16'd40386, 16'd42861});
	test_expansion(128'h0a7d4e2b60f166a503658da58811c9f7, {16'd54148, 16'd42458, 16'd18480, 16'd51787, 16'd65250, 16'd37923, 16'd37054, 16'd18961, 16'd7246, 16'd33129, 16'd40687, 16'd60176, 16'd52894, 16'd62124, 16'd41939, 16'd6566, 16'd38128, 16'd34295, 16'd53766, 16'd62118, 16'd6645, 16'd2770, 16'd13943, 16'd21237, 16'd13069, 16'd1328});
	test_expansion(128'h47ee03b5e62536bcc1779061c254d354, {16'd40119, 16'd64965, 16'd39555, 16'd12423, 16'd61225, 16'd46380, 16'd33480, 16'd46486, 16'd23134, 16'd27898, 16'd43484, 16'd63798, 16'd56456, 16'd56841, 16'd13052, 16'd47928, 16'd658, 16'd64864, 16'd13934, 16'd34655, 16'd24390, 16'd62736, 16'd25089, 16'd6672, 16'd59932, 16'd65326});
	test_expansion(128'h666fd02215c44c57cc7add339f2e5ea5, {16'd37724, 16'd26365, 16'd64035, 16'd4806, 16'd3644, 16'd43468, 16'd52779, 16'd54183, 16'd9391, 16'd6617, 16'd57330, 16'd20031, 16'd61870, 16'd46390, 16'd60538, 16'd1454, 16'd28588, 16'd47038, 16'd10465, 16'd44677, 16'd20183, 16'd45375, 16'd20574, 16'd26483, 16'd19330, 16'd63874});
	test_expansion(128'he6c7791c1d4fd2bfdb976549cecd2d8e, {16'd53361, 16'd40324, 16'd52295, 16'd16537, 16'd41933, 16'd509, 16'd17495, 16'd20990, 16'd65261, 16'd63136, 16'd20116, 16'd11376, 16'd39501, 16'd55338, 16'd8580, 16'd8191, 16'd28560, 16'd21649, 16'd65200, 16'd57887, 16'd7552, 16'd17651, 16'd10867, 16'd21988, 16'd14116, 16'd48741});
	test_expansion(128'h80d774504aadb8d89deb2addb6fec442, {16'd17433, 16'd33450, 16'd31428, 16'd7380, 16'd10305, 16'd13328, 16'd59721, 16'd35461, 16'd47250, 16'd22646, 16'd12310, 16'd39161, 16'd57455, 16'd24105, 16'd406, 16'd19898, 16'd15819, 16'd23601, 16'd61752, 16'd34641, 16'd22636, 16'd60071, 16'd47147, 16'd36985, 16'd3118, 16'd44235});
	test_expansion(128'h0e790aabc42b592d10ef878fb4710be0, {16'd10605, 16'd61731, 16'd626, 16'd1830, 16'd60013, 16'd44244, 16'd35644, 16'd8789, 16'd63987, 16'd57174, 16'd13271, 16'd4039, 16'd25908, 16'd27124, 16'd58353, 16'd59844, 16'd16972, 16'd48748, 16'd18992, 16'd46755, 16'd50060, 16'd3256, 16'd58014, 16'd7778, 16'd49145, 16'd57474});
	test_expansion(128'h414068e40cd754e78b22f76c418bc7e8, {16'd35207, 16'd50931, 16'd58249, 16'd62165, 16'd53544, 16'd57565, 16'd24408, 16'd20885, 16'd24277, 16'd48841, 16'd3402, 16'd17057, 16'd5874, 16'd63832, 16'd39051, 16'd56981, 16'd51899, 16'd2282, 16'd34929, 16'd52826, 16'd37713, 16'd61728, 16'd1028, 16'd13921, 16'd21882, 16'd21771});
	test_expansion(128'hfe4c18a7170e422853d71f6172749f32, {16'd37470, 16'd20924, 16'd7878, 16'd58320, 16'd2428, 16'd51526, 16'd14681, 16'd60892, 16'd16383, 16'd19890, 16'd25717, 16'd45396, 16'd65066, 16'd38362, 16'd62509, 16'd61202, 16'd41314, 16'd3984, 16'd12855, 16'd38962, 16'd16951, 16'd30166, 16'd25613, 16'd44163, 16'd59518, 16'd50526});
	test_expansion(128'haca27e2be34e0b9695634fea026ac5c0, {16'd18480, 16'd21395, 16'd38692, 16'd52466, 16'd40177, 16'd55821, 16'd36668, 16'd24150, 16'd27633, 16'd38828, 16'd13461, 16'd1198, 16'd44908, 16'd39526, 16'd23426, 16'd62362, 16'd47198, 16'd34562, 16'd3092, 16'd38342, 16'd56607, 16'd24795, 16'd589, 16'd46810, 16'd51853, 16'd62816});
	test_expansion(128'h26d3e1a1f5a345cc572ca83946b73dbb, {16'd54066, 16'd10013, 16'd16140, 16'd63934, 16'd42235, 16'd429, 16'd16210, 16'd63811, 16'd18090, 16'd52274, 16'd6682, 16'd37916, 16'd6170, 16'd59853, 16'd12209, 16'd56595, 16'd41387, 16'd50634, 16'd25205, 16'd60892, 16'd46284, 16'd20493, 16'd40195, 16'd46579, 16'd32110, 16'd56950});
	test_expansion(128'h7c0d4a66f378bef2daa56c22b78665a6, {16'd42122, 16'd29535, 16'd22150, 16'd56462, 16'd38396, 16'd9817, 16'd9057, 16'd18874, 16'd2158, 16'd4988, 16'd25521, 16'd55236, 16'd7699, 16'd16977, 16'd19229, 16'd41930, 16'd41074, 16'd40471, 16'd18143, 16'd64365, 16'd33847, 16'd6162, 16'd52594, 16'd50648, 16'd34173, 16'd59136});
	test_expansion(128'h74c5963cd76c3026d38382b129034dd6, {16'd47525, 16'd60662, 16'd12216, 16'd42831, 16'd37801, 16'd11344, 16'd61419, 16'd8370, 16'd18339, 16'd64979, 16'd56424, 16'd23684, 16'd39979, 16'd21433, 16'd19307, 16'd63147, 16'd14613, 16'd46964, 16'd33483, 16'd49677, 16'd5078, 16'd3432, 16'd35697, 16'd2104, 16'd35069, 16'd42908});
	test_expansion(128'h6ebef5737e03003624a994b4b5296306, {16'd41236, 16'd60867, 16'd29284, 16'd38648, 16'd1134, 16'd36071, 16'd12352, 16'd14150, 16'd44521, 16'd45433, 16'd26551, 16'd62177, 16'd45589, 16'd13466, 16'd15443, 16'd5095, 16'd54196, 16'd38633, 16'd16630, 16'd37526, 16'd63573, 16'd53394, 16'd35679, 16'd40542, 16'd18245, 16'd39698});
	test_expansion(128'h6e94afce2ac8a3ced885d0197ba1c2fc, {16'd61683, 16'd10893, 16'd55224, 16'd51248, 16'd59217, 16'd30660, 16'd43975, 16'd15120, 16'd38386, 16'd54480, 16'd15601, 16'd4209, 16'd58403, 16'd27098, 16'd34915, 16'd17245, 16'd25105, 16'd44056, 16'd46541, 16'd32941, 16'd7051, 16'd11483, 16'd42133, 16'd58389, 16'd36486, 16'd1302});
	test_expansion(128'hd2a0abbcec83a5944090aff61a739b85, {16'd27657, 16'd59501, 16'd17834, 16'd2302, 16'd22529, 16'd14123, 16'd14580, 16'd34727, 16'd26205, 16'd24375, 16'd22038, 16'd57945, 16'd10838, 16'd61303, 16'd32858, 16'd29761, 16'd46214, 16'd46750, 16'd22112, 16'd49895, 16'd47179, 16'd21288, 16'd3633, 16'd42380, 16'd17312, 16'd14399});
	test_expansion(128'ha715cf6e11f8ae4da1f3c21d79c661f2, {16'd9895, 16'd24609, 16'd2671, 16'd63746, 16'd18299, 16'd52158, 16'd11405, 16'd22421, 16'd49498, 16'd58432, 16'd20400, 16'd8491, 16'd20985, 16'd9137, 16'd41705, 16'd32224, 16'd3120, 16'd52340, 16'd9528, 16'd16228, 16'd1087, 16'd20589, 16'd58141, 16'd55377, 16'd4077, 16'd54521});
	test_expansion(128'h0a5962e2ca8d72a4c9a540fd2b27f47e, {16'd10343, 16'd62706, 16'd37815, 16'd43854, 16'd30492, 16'd5321, 16'd11621, 16'd57187, 16'd15599, 16'd52663, 16'd28622, 16'd4821, 16'd2674, 16'd45596, 16'd59653, 16'd4938, 16'd60374, 16'd7234, 16'd58699, 16'd43240, 16'd20385, 16'd57904, 16'd12772, 16'd15003, 16'd39777, 16'd9046});
	test_expansion(128'h2ff11db2a543639638965588c9e7cee4, {16'd53214, 16'd20039, 16'd63281, 16'd24421, 16'd10439, 16'd63222, 16'd26050, 16'd19548, 16'd27283, 16'd58564, 16'd287, 16'd13958, 16'd28453, 16'd48044, 16'd15147, 16'd63674, 16'd3293, 16'd35510, 16'd41530, 16'd55118, 16'd24997, 16'd8723, 16'd19102, 16'd13133, 16'd45067, 16'd56851});
	test_expansion(128'he41ee2a81dced2bf08da3a000125fcca, {16'd14298, 16'd25255, 16'd11366, 16'd12259, 16'd30495, 16'd38724, 16'd15719, 16'd22732, 16'd35282, 16'd19117, 16'd65366, 16'd11674, 16'd22016, 16'd4233, 16'd25753, 16'd8621, 16'd59993, 16'd39974, 16'd17700, 16'd22973, 16'd61808, 16'd35340, 16'd45728, 16'd34500, 16'd21454, 16'd4971});
	test_expansion(128'hdcd8466ec7bd075fec460e1855c5ec80, {16'd11484, 16'd46655, 16'd23180, 16'd25567, 16'd14823, 16'd28350, 16'd33959, 16'd33742, 16'd9051, 16'd50435, 16'd39665, 16'd22056, 16'd26198, 16'd53201, 16'd49873, 16'd46741, 16'd6787, 16'd44208, 16'd27293, 16'd5473, 16'd14027, 16'd28503, 16'd19078, 16'd64537, 16'd47601, 16'd20962});
	test_expansion(128'hf552dd6fcfe30bae5feb742c4f07ebf9, {16'd31862, 16'd62819, 16'd35140, 16'd3412, 16'd27111, 16'd7038, 16'd3282, 16'd9414, 16'd11923, 16'd2496, 16'd2794, 16'd34338, 16'd32158, 16'd30341, 16'd43796, 16'd5135, 16'd55489, 16'd10799, 16'd37530, 16'd21409, 16'd25621, 16'd64758, 16'd36722, 16'd55205, 16'd2661, 16'd18205});
	test_expansion(128'h4ec503cb1a7a3a664a9d8cdade887377, {16'd65219, 16'd47039, 16'd42300, 16'd11978, 16'd53504, 16'd18424, 16'd9804, 16'd60154, 16'd39949, 16'd23715, 16'd39301, 16'd44421, 16'd28604, 16'd23222, 16'd30216, 16'd32661, 16'd38218, 16'd55187, 16'd35954, 16'd14553, 16'd40102, 16'd44510, 16'd6748, 16'd48273, 16'd25630, 16'd6879});
	test_expansion(128'h41ca9c602518e20df7b2ec2e8ddad802, {16'd20030, 16'd17839, 16'd38796, 16'd14544, 16'd48248, 16'd58634, 16'd27824, 16'd10053, 16'd26685, 16'd54410, 16'd6114, 16'd25832, 16'd29002, 16'd14242, 16'd34213, 16'd23616, 16'd60273, 16'd62304, 16'd44280, 16'd32683, 16'd52104, 16'd20268, 16'd13236, 16'd65036, 16'd60106, 16'd36361});
	test_expansion(128'h64325bf5ccc71ccb8953b985e84c95d9, {16'd6541, 16'd49819, 16'd11378, 16'd40413, 16'd48832, 16'd4037, 16'd9012, 16'd167, 16'd37463, 16'd42572, 16'd43883, 16'd11075, 16'd53949, 16'd48140, 16'd25176, 16'd9844, 16'd21608, 16'd42243, 16'd4508, 16'd7558, 16'd7743, 16'd26522, 16'd23626, 16'd31994, 16'd54829, 16'd23245});
	test_expansion(128'hb0e904183ce75d817c402dccaa0b469e, {16'd63734, 16'd41323, 16'd60070, 16'd55123, 16'd27876, 16'd62744, 16'd23532, 16'd17454, 16'd38301, 16'd38290, 16'd17953, 16'd37624, 16'd59226, 16'd24956, 16'd27200, 16'd25353, 16'd40727, 16'd19481, 16'd368, 16'd11834, 16'd809, 16'd33594, 16'd4877, 16'd30356, 16'd3900, 16'd40646});
	test_expansion(128'h1992bba85743dadc8cc0044038a69c80, {16'd47626, 16'd6504, 16'd22817, 16'd33519, 16'd45318, 16'd61190, 16'd32502, 16'd8937, 16'd31230, 16'd415, 16'd53605, 16'd46751, 16'd53914, 16'd51964, 16'd23997, 16'd50712, 16'd22748, 16'd57637, 16'd53378, 16'd8260, 16'd20385, 16'd12079, 16'd18454, 16'd25075, 16'd40691, 16'd57081});
	test_expansion(128'h8d6feb23dae3b2b31d163ccbe483398c, {16'd17779, 16'd43117, 16'd21353, 16'd9321, 16'd62136, 16'd24891, 16'd17357, 16'd37480, 16'd35499, 16'd18696, 16'd22159, 16'd37459, 16'd49539, 16'd47356, 16'd5716, 16'd33978, 16'd36020, 16'd28144, 16'd39905, 16'd29563, 16'd2078, 16'd63510, 16'd45493, 16'd63075, 16'd57549, 16'd31943});
	test_expansion(128'h17ba4071c8cca169171c3a1c943760bf, {16'd33399, 16'd21447, 16'd51885, 16'd58131, 16'd31192, 16'd58727, 16'd10829, 16'd15721, 16'd4801, 16'd64491, 16'd16803, 16'd10661, 16'd32094, 16'd48778, 16'd20461, 16'd39754, 16'd53155, 16'd39956, 16'd46819, 16'd45563, 16'd4118, 16'd64757, 16'd3218, 16'd13790, 16'd57565, 16'd11865});
	test_expansion(128'h9810cb1f011cb173c24b83877ab23210, {16'd64044, 16'd31679, 16'd4705, 16'd54908, 16'd21536, 16'd21746, 16'd56942, 16'd48285, 16'd17392, 16'd49094, 16'd35133, 16'd9292, 16'd46941, 16'd54960, 16'd35526, 16'd47959, 16'd40988, 16'd64129, 16'd12615, 16'd34607, 16'd2338, 16'd49403, 16'd22070, 16'd24667, 16'd8644, 16'd52847});
	test_expansion(128'h5bd519c7de358e0838e34d4931b7c256, {16'd37586, 16'd23667, 16'd31763, 16'd32736, 16'd33918, 16'd28998, 16'd14656, 16'd50211, 16'd43204, 16'd47616, 16'd43674, 16'd37771, 16'd33776, 16'd42715, 16'd12450, 16'd31657, 16'd44556, 16'd21278, 16'd6414, 16'd36845, 16'd26034, 16'd736, 16'd11216, 16'd24509, 16'd26465, 16'd51557});
	test_expansion(128'hee74154973ab7c32d6a35b689a7d6cf9, {16'd41260, 16'd46430, 16'd28036, 16'd17543, 16'd65323, 16'd6244, 16'd52463, 16'd11769, 16'd55966, 16'd125, 16'd37415, 16'd49454, 16'd1639, 16'd45152, 16'd10285, 16'd9868, 16'd53561, 16'd1472, 16'd13697, 16'd64804, 16'd35080, 16'd13011, 16'd48511, 16'd35767, 16'd33695, 16'd22017});
	test_expansion(128'h01349cb7c957b1a4021bde56617ce421, {16'd53233, 16'd23710, 16'd13307, 16'd46182, 16'd12491, 16'd35706, 16'd12168, 16'd40697, 16'd17059, 16'd49750, 16'd32989, 16'd57296, 16'd34939, 16'd52758, 16'd9119, 16'd32633, 16'd56494, 16'd21903, 16'd42183, 16'd247, 16'd35687, 16'd24454, 16'd26571, 16'd40483, 16'd21017, 16'd44851});
	test_expansion(128'hc41fff41c855f5bc2f10977ea00d56aa, {16'd43825, 16'd22716, 16'd691, 16'd12015, 16'd56925, 16'd1165, 16'd47130, 16'd18945, 16'd6175, 16'd53174, 16'd29994, 16'd65137, 16'd38643, 16'd13109, 16'd37293, 16'd29943, 16'd13397, 16'd56749, 16'd6415, 16'd61760, 16'd64557, 16'd10565, 16'd56773, 16'd11451, 16'd54272, 16'd42767});
	test_expansion(128'ha3ef0b466e78568c864744e462a24fa8, {16'd1947, 16'd24499, 16'd10691, 16'd21571, 16'd3313, 16'd52826, 16'd38895, 16'd44047, 16'd17150, 16'd56191, 16'd7114, 16'd42390, 16'd10262, 16'd45259, 16'd39256, 16'd57869, 16'd57825, 16'd56173, 16'd24524, 16'd57911, 16'd33536, 16'd50501, 16'd30998, 16'd48559, 16'd26592, 16'd49123});
	test_expansion(128'h190d53c652f7a4909d35384f70f2bdec, {16'd18864, 16'd28587, 16'd5805, 16'd8963, 16'd14126, 16'd17546, 16'd44321, 16'd2208, 16'd10771, 16'd41871, 16'd11597, 16'd5891, 16'd15313, 16'd30645, 16'd21890, 16'd44204, 16'd51560, 16'd44008, 16'd55341, 16'd32059, 16'd63016, 16'd19945, 16'd61157, 16'd35830, 16'd23892, 16'd2801});
	test_expansion(128'h4e15ae5f4e7951fe7efefd27096fb266, {16'd48434, 16'd65250, 16'd17284, 16'd43044, 16'd21692, 16'd12821, 16'd61115, 16'd2822, 16'd35906, 16'd50131, 16'd11028, 16'd7641, 16'd3831, 16'd44405, 16'd46717, 16'd1802, 16'd12593, 16'd2939, 16'd8613, 16'd43994, 16'd60757, 16'd42541, 16'd61570, 16'd65163, 16'd47690, 16'd15548});
	test_expansion(128'hea8ed7cf1a7fc177a5030b1ba222374d, {16'd6952, 16'd29602, 16'd16525, 16'd6285, 16'd56517, 16'd32490, 16'd1398, 16'd64854, 16'd57057, 16'd33729, 16'd39725, 16'd33613, 16'd20038, 16'd52764, 16'd54484, 16'd27128, 16'd18101, 16'd54462, 16'd3711, 16'd25362, 16'd62604, 16'd58309, 16'd59113, 16'd41132, 16'd56048, 16'd23511});
	test_expansion(128'h90795638b02aea8bfc7d82d4293261cd, {16'd36139, 16'd41826, 16'd28143, 16'd45468, 16'd13582, 16'd42191, 16'd46347, 16'd18841, 16'd45563, 16'd64134, 16'd44090, 16'd36576, 16'd64252, 16'd33407, 16'd19147, 16'd37615, 16'd25507, 16'd47441, 16'd25305, 16'd29231, 16'd12032, 16'd29029, 16'd48374, 16'd40145, 16'd10964, 16'd1495});
	test_expansion(128'h588dd3cfe097c3f82b586cea53bc3b84, {16'd33930, 16'd35918, 16'd17244, 16'd11633, 16'd58903, 16'd43395, 16'd4248, 16'd37285, 16'd27980, 16'd56677, 16'd50352, 16'd57187, 16'd38232, 16'd489, 16'd53715, 16'd31457, 16'd1770, 16'd46992, 16'd8171, 16'd65247, 16'd24748, 16'd43621, 16'd849, 16'd57497, 16'd55482, 16'd39636});
	test_expansion(128'h989642fcf19508ae06392941f30a56e2, {16'd34003, 16'd60737, 16'd828, 16'd28555, 16'd52603, 16'd28506, 16'd62752, 16'd42568, 16'd37219, 16'd48854, 16'd64463, 16'd59392, 16'd44467, 16'd44517, 16'd52307, 16'd64875, 16'd56156, 16'd49989, 16'd31869, 16'd15436, 16'd62650, 16'd22918, 16'd13870, 16'd27412, 16'd37172, 16'd25956});
	test_expansion(128'he9f8d82ee65ec48c173e9d295e43771f, {16'd57086, 16'd17752, 16'd32543, 16'd26705, 16'd63335, 16'd12879, 16'd63304, 16'd46956, 16'd5306, 16'd20334, 16'd14838, 16'd16446, 16'd32977, 16'd61637, 16'd55161, 16'd32099, 16'd10703, 16'd53113, 16'd43215, 16'd26074, 16'd53174, 16'd17892, 16'd48870, 16'd32190, 16'd41612, 16'd26976});
	test_expansion(128'h7f914bedb2ecd37d1522840a4c34ba1b, {16'd31180, 16'd36279, 16'd53172, 16'd24118, 16'd18884, 16'd37011, 16'd22174, 16'd36165, 16'd31397, 16'd7510, 16'd10182, 16'd64070, 16'd4329, 16'd15684, 16'd47098, 16'd14957, 16'd11793, 16'd2034, 16'd48625, 16'd51298, 16'd37795, 16'd24677, 16'd48315, 16'd58637, 16'd45967, 16'd52804});
	test_expansion(128'h1ad97d1326423a09abbd4ce6cb6a7f0e, {16'd39127, 16'd26081, 16'd59031, 16'd22307, 16'd18142, 16'd3734, 16'd46103, 16'd8797, 16'd13568, 16'd22475, 16'd62238, 16'd322, 16'd43464, 16'd47241, 16'd43, 16'd17008, 16'd38623, 16'd43208, 16'd52651, 16'd42478, 16'd51464, 16'd4830, 16'd50898, 16'd14296, 16'd3471, 16'd46325});
	test_expansion(128'hfb6552eb11685085341a2f9021d588cd, {16'd32750, 16'd13893, 16'd15036, 16'd42685, 16'd47339, 16'd35653, 16'd4342, 16'd32893, 16'd25629, 16'd62606, 16'd25635, 16'd36437, 16'd52995, 16'd2994, 16'd63033, 16'd40953, 16'd36582, 16'd22647, 16'd42177, 16'd33211, 16'd33355, 16'd33016, 16'd21120, 16'd6411, 16'd16289, 16'd30800});
	test_expansion(128'hf8111fda3a8b816da8aabd5e0c97b6ff, {16'd10812, 16'd48673, 16'd46283, 16'd15645, 16'd13240, 16'd32646, 16'd38857, 16'd5847, 16'd10659, 16'd8925, 16'd48583, 16'd48160, 16'd43952, 16'd14881, 16'd25503, 16'd35030, 16'd31224, 16'd56810, 16'd1331, 16'd30776, 16'd8435, 16'd38470, 16'd22009, 16'd8169, 16'd61268, 16'd38702});
	test_expansion(128'h08bf4f35e7ae110ce4c6a85ba588075a, {16'd34761, 16'd51461, 16'd4421, 16'd22481, 16'd62795, 16'd44584, 16'd3286, 16'd28718, 16'd17285, 16'd58472, 16'd40441, 16'd1662, 16'd821, 16'd45466, 16'd8375, 16'd47117, 16'd6528, 16'd18380, 16'd9394, 16'd53984, 16'd2411, 16'd52911, 16'd38221, 16'd26436, 16'd42691, 16'd33558});
	test_expansion(128'h05d7a4723cbc91d2738342001ac6a9a1, {16'd27835, 16'd48146, 16'd4204, 16'd28074, 16'd20211, 16'd55972, 16'd9119, 16'd84, 16'd12164, 16'd36408, 16'd4378, 16'd63322, 16'd3901, 16'd20175, 16'd36496, 16'd5542, 16'd35480, 16'd3157, 16'd56508, 16'd30884, 16'd13683, 16'd46496, 16'd63569, 16'd30206, 16'd22257, 16'd37762});
	test_expansion(128'h074fb202c1875b50ed003cf477982629, {16'd59143, 16'd22914, 16'd39729, 16'd65385, 16'd10421, 16'd44531, 16'd26310, 16'd57699, 16'd55263, 16'd8666, 16'd34560, 16'd41487, 16'd58606, 16'd21320, 16'd60656, 16'd48311, 16'd42834, 16'd3593, 16'd44150, 16'd2824, 16'd795, 16'd29046, 16'd2470, 16'd9878, 16'd19485, 16'd1065});
	test_expansion(128'h6c153481e3dd627420cad2922085c85f, {16'd21663, 16'd37058, 16'd22376, 16'd16304, 16'd58912, 16'd42692, 16'd30430, 16'd39849, 16'd29888, 16'd41299, 16'd11476, 16'd14341, 16'd62094, 16'd62845, 16'd46158, 16'd56454, 16'd19165, 16'd42883, 16'd13656, 16'd26751, 16'd4104, 16'd58188, 16'd63514, 16'd2514, 16'd5903, 16'd3258});
	test_expansion(128'h514d00d272743403507306a0d293949b, {16'd10022, 16'd56944, 16'd29128, 16'd34481, 16'd25873, 16'd22844, 16'd64293, 16'd53519, 16'd3173, 16'd28127, 16'd34746, 16'd28215, 16'd55385, 16'd27318, 16'd11470, 16'd28909, 16'd51216, 16'd1942, 16'd47547, 16'd4895, 16'd59888, 16'd53875, 16'd21584, 16'd29700, 16'd10459, 16'd5853});
	test_expansion(128'hf82e991a5f9e80854482bee045eaa63a, {16'd20337, 16'd43961, 16'd62222, 16'd52455, 16'd32454, 16'd56742, 16'd45152, 16'd18264, 16'd60531, 16'd29550, 16'd27471, 16'd47839, 16'd26862, 16'd21402, 16'd59833, 16'd34848, 16'd39987, 16'd57184, 16'd20987, 16'd22100, 16'd28287, 16'd1381, 16'd43870, 16'd6321, 16'd34302, 16'd28822});
	test_expansion(128'h89539e53c80bcf1f4b54efb9ba723e3b, {16'd13666, 16'd55905, 16'd29477, 16'd22937, 16'd58979, 16'd61292, 16'd33157, 16'd5917, 16'd33615, 16'd20383, 16'd58269, 16'd45472, 16'd23142, 16'd48192, 16'd17790, 16'd41817, 16'd31531, 16'd12437, 16'd22780, 16'd34507, 16'd63855, 16'd63988, 16'd17995, 16'd57042, 16'd9774, 16'd54620});
	test_expansion(128'ha0448e85a1bbea1b8f49155d02a434e9, {16'd59446, 16'd29322, 16'd48687, 16'd42664, 16'd33880, 16'd50142, 16'd47552, 16'd51719, 16'd52822, 16'd54181, 16'd49461, 16'd25836, 16'd61343, 16'd12092, 16'd12990, 16'd42832, 16'd27037, 16'd49613, 16'd26775, 16'd5410, 16'd57267, 16'd29630, 16'd28504, 16'd13517, 16'd21346, 16'd53639});
	test_expansion(128'h1b00fb4416a8ce182a9ef8f89d2480d6, {16'd61732, 16'd13258, 16'd59922, 16'd56161, 16'd39138, 16'd7795, 16'd20829, 16'd37653, 16'd7617, 16'd44590, 16'd30500, 16'd10209, 16'd3512, 16'd54384, 16'd54214, 16'd51669, 16'd63506, 16'd53677, 16'd62610, 16'd54686, 16'd18285, 16'd27978, 16'd3896, 16'd3570, 16'd55037, 16'd61897});
	test_expansion(128'h155f4447207e89fc5c208deaf659850f, {16'd20835, 16'd13946, 16'd2505, 16'd52038, 16'd8751, 16'd29078, 16'd64064, 16'd43599, 16'd50791, 16'd5355, 16'd9183, 16'd5274, 16'd21905, 16'd37738, 16'd30025, 16'd28649, 16'd64579, 16'd56674, 16'd18642, 16'd43493, 16'd21526, 16'd54163, 16'd42553, 16'd25929, 16'd60157, 16'd6879});
	test_expansion(128'h8a6d2d8887e60e06dd567156334c55a4, {16'd59735, 16'd39089, 16'd31241, 16'd25273, 16'd27628, 16'd60070, 16'd7851, 16'd18822, 16'd62144, 16'd56668, 16'd36148, 16'd3008, 16'd55934, 16'd34423, 16'd11693, 16'd43974, 16'd15477, 16'd54093, 16'd64962, 16'd60120, 16'd44073, 16'd12604, 16'd58158, 16'd47050, 16'd27387, 16'd47786});
	test_expansion(128'h5cc19cf03ecdfaedd3696c64b77908b7, {16'd50437, 16'd14538, 16'd47770, 16'd42025, 16'd33579, 16'd10112, 16'd10243, 16'd28994, 16'd39430, 16'd26362, 16'd6008, 16'd31657, 16'd53115, 16'd4341, 16'd45023, 16'd2804, 16'd51036, 16'd40778, 16'd63947, 16'd61441, 16'd28675, 16'd8235, 16'd1710, 16'd8862, 16'd8529, 16'd5367});
	test_expansion(128'hd8046b5b2e7aca354c7f25774f64c362, {16'd35599, 16'd50934, 16'd15916, 16'd44974, 16'd34459, 16'd13761, 16'd31859, 16'd1740, 16'd35221, 16'd16465, 16'd52024, 16'd18967, 16'd9839, 16'd39289, 16'd28706, 16'd51700, 16'd62427, 16'd62025, 16'd39252, 16'd43881, 16'd56690, 16'd49614, 16'd6830, 16'd16616, 16'd9192, 16'd44669});
	test_expansion(128'hba120d6dd04718380b0b26d9fca4bb11, {16'd36505, 16'd55592, 16'd34106, 16'd7877, 16'd34457, 16'd11141, 16'd15038, 16'd50030, 16'd38882, 16'd29032, 16'd31812, 16'd36303, 16'd6279, 16'd31096, 16'd47124, 16'd36555, 16'd27256, 16'd46296, 16'd60488, 16'd37007, 16'd4727, 16'd56287, 16'd41583, 16'd60921, 16'd39257, 16'd2245});
	test_expansion(128'h224a8342e0e97efaef5f939dbbf25253, {16'd49268, 16'd54167, 16'd31678, 16'd52481, 16'd8947, 16'd5072, 16'd53267, 16'd4875, 16'd49723, 16'd54100, 16'd1383, 16'd51799, 16'd42653, 16'd29517, 16'd33936, 16'd8087, 16'd31138, 16'd61304, 16'd49454, 16'd63969, 16'd17587, 16'd52889, 16'd19229, 16'd53147, 16'd21431, 16'd59341});
	test_expansion(128'h653318ded4deb17374d2feafb1969761, {16'd10183, 16'd16121, 16'd24175, 16'd62039, 16'd55266, 16'd54829, 16'd29957, 16'd62357, 16'd65177, 16'd38264, 16'd23106, 16'd18231, 16'd24463, 16'd46961, 16'd50760, 16'd2317, 16'd37409, 16'd21539, 16'd51571, 16'd43253, 16'd54820, 16'd35516, 16'd29586, 16'd3840, 16'd15827, 16'd48417});
	test_expansion(128'h695b5cf9187ac614bc8e75f2a4dacc36, {16'd6148, 16'd36426, 16'd11675, 16'd47995, 16'd15468, 16'd1072, 16'd55625, 16'd16802, 16'd39414, 16'd51346, 16'd47458, 16'd18218, 16'd29487, 16'd21678, 16'd40901, 16'd27668, 16'd63453, 16'd6386, 16'd60319, 16'd9037, 16'd34971, 16'd27832, 16'd1213, 16'd21032, 16'd27223, 16'd19619});
	test_expansion(128'h13421ed49038f9ef2eafb0e4dfbcc0f6, {16'd1928, 16'd51142, 16'd60867, 16'd56376, 16'd19477, 16'd6410, 16'd64313, 16'd49774, 16'd48917, 16'd61771, 16'd56382, 16'd50321, 16'd49095, 16'd59612, 16'd31036, 16'd26467, 16'd31062, 16'd9248, 16'd54188, 16'd30654, 16'd30753, 16'd36314, 16'd53552, 16'd41981, 16'd29638, 16'd31501});
	test_expansion(128'hd0e2a6091124cee416edbed226a0241b, {16'd56551, 16'd53202, 16'd54026, 16'd16650, 16'd10970, 16'd59378, 16'd63869, 16'd20834, 16'd45180, 16'd5844, 16'd17197, 16'd57773, 16'd15484, 16'd28661, 16'd42716, 16'd50907, 16'd38926, 16'd27312, 16'd63969, 16'd35113, 16'd5056, 16'd19084, 16'd672, 16'd41874, 16'd11994, 16'd13140});
	test_expansion(128'hce1baf3f8542923a555f544ef3d3f59c, {16'd57549, 16'd32924, 16'd23550, 16'd52208, 16'd50561, 16'd2282, 16'd12539, 16'd12487, 16'd19545, 16'd60207, 16'd26882, 16'd17111, 16'd6796, 16'd53262, 16'd32546, 16'd12899, 16'd59574, 16'd21432, 16'd20275, 16'd10998, 16'd9727, 16'd53446, 16'd19109, 16'd62655, 16'd1071, 16'd25999});
	test_expansion(128'h1d207cff2d1fe0bf904ccd9670574ba1, {16'd23814, 16'd54541, 16'd20700, 16'd54040, 16'd43291, 16'd54680, 16'd17606, 16'd35509, 16'd40079, 16'd50031, 16'd55058, 16'd8815, 16'd24495, 16'd53125, 16'd64598, 16'd65380, 16'd63669, 16'd54916, 16'd34067, 16'd34277, 16'd36232, 16'd13082, 16'd42573, 16'd27565, 16'd18969, 16'd48722});
	test_expansion(128'hc4379c4a41175e5da46d39649e7d8593, {16'd60782, 16'd25758, 16'd26412, 16'd25678, 16'd63833, 16'd43330, 16'd28833, 16'd18486, 16'd5112, 16'd62024, 16'd11965, 16'd37153, 16'd15969, 16'd58324, 16'd14392, 16'd43269, 16'd27171, 16'd40998, 16'd55278, 16'd32388, 16'd51686, 16'd8319, 16'd1792, 16'd9208, 16'd49156, 16'd37457});
	test_expansion(128'h2e2720f3446536c02f0e054f5f14e7d9, {16'd47933, 16'd47862, 16'd58796, 16'd39701, 16'd12911, 16'd17535, 16'd763, 16'd16394, 16'd47556, 16'd56179, 16'd45003, 16'd29922, 16'd17449, 16'd10011, 16'd52, 16'd6313, 16'd41391, 16'd28979, 16'd31430, 16'd53073, 16'd35139, 16'd11661, 16'd14747, 16'd26179, 16'd22557, 16'd2638});
	test_expansion(128'hd1073cee51c598d5fb379acdac5448fe, {16'd34736, 16'd48499, 16'd25540, 16'd15209, 16'd30667, 16'd56702, 16'd12968, 16'd2712, 16'd43662, 16'd55350, 16'd60480, 16'd2617, 16'd3788, 16'd10786, 16'd40712, 16'd14457, 16'd34753, 16'd36394, 16'd17073, 16'd33472, 16'd60890, 16'd36430, 16'd59528, 16'd30010, 16'd55576, 16'd25816});
	test_expansion(128'he991a78336cefea5641aa1c6e777c9d7, {16'd55595, 16'd14881, 16'd38800, 16'd43945, 16'd44164, 16'd4031, 16'd62628, 16'd13575, 16'd24815, 16'd27432, 16'd51995, 16'd5922, 16'd35048, 16'd32780, 16'd52128, 16'd79, 16'd3058, 16'd24363, 16'd26710, 16'd49095, 16'd63996, 16'd45672, 16'd48736, 16'd54434, 16'd59555, 16'd36512});
	test_expansion(128'h853b5f0beee12d74102eb8d65735cfcb, {16'd62706, 16'd9750, 16'd65067, 16'd4311, 16'd51834, 16'd41417, 16'd62801, 16'd16649, 16'd34938, 16'd63166, 16'd7311, 16'd61633, 16'd45365, 16'd39919, 16'd16779, 16'd7113, 16'd5209, 16'd5418, 16'd57493, 16'd41961, 16'd60052, 16'd13274, 16'd30007, 16'd51616, 16'd50245, 16'd9188});
	test_expansion(128'ha9bc28d36cfd892f86742ce4a043b5e9, {16'd10648, 16'd47522, 16'd17178, 16'd33817, 16'd44762, 16'd4238, 16'd62870, 16'd13383, 16'd55747, 16'd35052, 16'd62821, 16'd49272, 16'd3908, 16'd4073, 16'd4252, 16'd7892, 16'd46874, 16'd32610, 16'd63682, 16'd57904, 16'd57000, 16'd40089, 16'd7, 16'd44687, 16'd61842, 16'd48569});
	test_expansion(128'hdfe6d8d00c210e81d4bf6f970f0abec7, {16'd7133, 16'd33461, 16'd14254, 16'd50346, 16'd32634, 16'd28158, 16'd42124, 16'd19651, 16'd20027, 16'd32494, 16'd53376, 16'd50765, 16'd9424, 16'd21805, 16'd31032, 16'd17327, 16'd3325, 16'd50874, 16'd39537, 16'd61231, 16'd59667, 16'd20535, 16'd48211, 16'd8507, 16'd56216, 16'd37902});
	test_expansion(128'ha0153885b4b251fe80203d393b6474ac, {16'd37988, 16'd56468, 16'd54458, 16'd28438, 16'd36148, 16'd46000, 16'd17279, 16'd20038, 16'd31939, 16'd27982, 16'd38538, 16'd62345, 16'd56707, 16'd12995, 16'd49570, 16'd37963, 16'd65049, 16'd64199, 16'd47943, 16'd41264, 16'd34849, 16'd62242, 16'd57221, 16'd8777, 16'd33513, 16'd22824});
	test_expansion(128'h448ab82be59dbfa1de6a8c84536c9053, {16'd53279, 16'd40200, 16'd6567, 16'd50758, 16'd1676, 16'd47531, 16'd9905, 16'd866, 16'd54108, 16'd9059, 16'd29068, 16'd21567, 16'd11465, 16'd1275, 16'd5863, 16'd6907, 16'd46530, 16'd13480, 16'd14003, 16'd44010, 16'd6764, 16'd45340, 16'd59440, 16'd14877, 16'd55363, 16'd64825});
	test_expansion(128'h5c074046ba2269e1f1f9ef4094ba9e3d, {16'd10888, 16'd42976, 16'd41603, 16'd13453, 16'd35795, 16'd27508, 16'd61895, 16'd32612, 16'd14618, 16'd32620, 16'd65118, 16'd27914, 16'd28885, 16'd34268, 16'd62591, 16'd1927, 16'd25924, 16'd58540, 16'd40110, 16'd57604, 16'd40075, 16'd23570, 16'd48162, 16'd42678, 16'd37850, 16'd10324});
	test_expansion(128'h0a3ada652ffdfba9b78d662e69d0a1c8, {16'd35275, 16'd41536, 16'd49391, 16'd24654, 16'd47322, 16'd30716, 16'd15868, 16'd57899, 16'd52556, 16'd13840, 16'd4449, 16'd1577, 16'd27094, 16'd23226, 16'd37418, 16'd65028, 16'd516, 16'd27447, 16'd59765, 16'd10299, 16'd65122, 16'd61457, 16'd5826, 16'd3280, 16'd63830, 16'd7913});
	test_expansion(128'hec4267a7a422993dac0cbfe98f738a13, {16'd30520, 16'd45699, 16'd57459, 16'd26422, 16'd45516, 16'd29385, 16'd7627, 16'd32270, 16'd42169, 16'd33606, 16'd31572, 16'd21101, 16'd26018, 16'd52460, 16'd52549, 16'd2659, 16'd18653, 16'd15944, 16'd22597, 16'd5650, 16'd23112, 16'd44285, 16'd5227, 16'd43946, 16'd43000, 16'd36602});
	test_expansion(128'h1e1e2d06c5d5e3a8e159f0ffcca94f00, {16'd11201, 16'd57040, 16'd35779, 16'd12165, 16'd32003, 16'd27818, 16'd57875, 16'd39223, 16'd19796, 16'd54136, 16'd2627, 16'd6800, 16'd19416, 16'd12008, 16'd15994, 16'd12849, 16'd62607, 16'd46492, 16'd8704, 16'd58074, 16'd46259, 16'd31934, 16'd23333, 16'd22530, 16'd20087, 16'd23663});
	test_expansion(128'h14018a02a420b1bc75920b79d3358754, {16'd63209, 16'd33305, 16'd9712, 16'd50017, 16'd47670, 16'd34229, 16'd60070, 16'd6112, 16'd10818, 16'd16836, 16'd62963, 16'd13801, 16'd5387, 16'd18755, 16'd6147, 16'd20903, 16'd17847, 16'd29284, 16'd54732, 16'd40398, 16'd2102, 16'd60354, 16'd44326, 16'd62071, 16'd15005, 16'd45902});
	test_expansion(128'h7fead7383eb8113ccab74e2b25f3d6bf, {16'd15077, 16'd19695, 16'd27266, 16'd13617, 16'd16998, 16'd53767, 16'd34479, 16'd816, 16'd36618, 16'd38534, 16'd32626, 16'd7927, 16'd1186, 16'd12208, 16'd36710, 16'd58745, 16'd37275, 16'd51462, 16'd3874, 16'd43487, 16'd64400, 16'd12080, 16'd4450, 16'd29517, 16'd31586, 16'd54181});
	test_expansion(128'had8526690ca5bdd4b25f8b1a7a522692, {16'd34607, 16'd62658, 16'd7192, 16'd50024, 16'd31446, 16'd13795, 16'd57974, 16'd41040, 16'd63251, 16'd16130, 16'd12676, 16'd34104, 16'd45188, 16'd24797, 16'd11665, 16'd24019, 16'd43357, 16'd1403, 16'd35918, 16'd53263, 16'd7659, 16'd55097, 16'd23011, 16'd40716, 16'd24305, 16'd25594});
	test_expansion(128'h210d3c13c79fb5551c9fb6442f7267f8, {16'd50135, 16'd56358, 16'd14941, 16'd33678, 16'd4544, 16'd8322, 16'd16074, 16'd54601, 16'd20924, 16'd12385, 16'd58417, 16'd42420, 16'd15948, 16'd47613, 16'd55887, 16'd12543, 16'd18203, 16'd19693, 16'd53962, 16'd58791, 16'd48063, 16'd41311, 16'd14951, 16'd9226, 16'd7408, 16'd15197});
	test_expansion(128'ha1dd6b3252d5f8cc4df917560f34d8f1, {16'd57592, 16'd16424, 16'd22816, 16'd30228, 16'd28242, 16'd10462, 16'd20165, 16'd28122, 16'd6124, 16'd65516, 16'd64308, 16'd63513, 16'd26203, 16'd42746, 16'd35392, 16'd52530, 16'd11535, 16'd46538, 16'd47607, 16'd54206, 16'd41512, 16'd6165, 16'd24451, 16'd60820, 16'd15595, 16'd57291});
	test_expansion(128'h1a17ef50133d7668c83625fc23c5fa42, {16'd13468, 16'd13414, 16'd52562, 16'd16316, 16'd33329, 16'd53781, 16'd11162, 16'd21072, 16'd37898, 16'd53824, 16'd64849, 16'd38897, 16'd24691, 16'd5086, 16'd51684, 16'd55140, 16'd53825, 16'd7443, 16'd26, 16'd61716, 16'd39312, 16'd59581, 16'd4463, 16'd9730, 16'd39109, 16'd53891});
	test_expansion(128'h35e9c2bc8bc7013ae8ecdfa9a2963273, {16'd65120, 16'd493, 16'd15206, 16'd11171, 16'd26383, 16'd39372, 16'd11424, 16'd41264, 16'd38732, 16'd51182, 16'd5339, 16'd41006, 16'd31956, 16'd59657, 16'd16581, 16'd47732, 16'd42693, 16'd17555, 16'd42343, 16'd61785, 16'd23266, 16'd15688, 16'd53599, 16'd52006, 16'd41553, 16'd36874});
	test_expansion(128'hcad046106a3cbe744217af4512032140, {16'd53982, 16'd10881, 16'd35751, 16'd60057, 16'd19224, 16'd9035, 16'd25262, 16'd23152, 16'd35178, 16'd13755, 16'd18225, 16'd56192, 16'd47763, 16'd34208, 16'd40609, 16'd30607, 16'd26596, 16'd38037, 16'd49714, 16'd6321, 16'd58317, 16'd34889, 16'd52545, 16'd83, 16'd3000, 16'd817});
	test_expansion(128'h8ab7e286d22ee6d9914cd259bc30750d, {16'd14028, 16'd19573, 16'd1543, 16'd4070, 16'd5106, 16'd50278, 16'd3412, 16'd1356, 16'd20629, 16'd28761, 16'd38267, 16'd15460, 16'd47242, 16'd11343, 16'd27653, 16'd26260, 16'd55297, 16'd35009, 16'd29522, 16'd60113, 16'd64349, 16'd19081, 16'd36195, 16'd65282, 16'd18073, 16'd58404});
	test_expansion(128'h1c152827846126b80fc8897f6aa08828, {16'd49626, 16'd7157, 16'd55513, 16'd47799, 16'd33827, 16'd52569, 16'd9999, 16'd19499, 16'd10080, 16'd14943, 16'd62930, 16'd35525, 16'd35238, 16'd37053, 16'd37814, 16'd58933, 16'd48305, 16'd38771, 16'd7907, 16'd47484, 16'd16191, 16'd42673, 16'd59816, 16'd56508, 16'd11714, 16'd22457});
	test_expansion(128'hba5661015107228655b4e8303c7a264e, {16'd12502, 16'd41885, 16'd29350, 16'd31626, 16'd43737, 16'd50129, 16'd29337, 16'd35171, 16'd58047, 16'd37520, 16'd44842, 16'd33097, 16'd4258, 16'd28916, 16'd24971, 16'd63765, 16'd50710, 16'd55340, 16'd52109, 16'd3842, 16'd48730, 16'd60430, 16'd54696, 16'd29442, 16'd3782, 16'd8006});
	test_expansion(128'h76abe9fbcd8a9ca37ef9383ce99ba843, {16'd3783, 16'd54047, 16'd31208, 16'd26326, 16'd57542, 16'd49461, 16'd48545, 16'd28478, 16'd25814, 16'd63087, 16'd64657, 16'd20843, 16'd47735, 16'd27686, 16'd45852, 16'd61649, 16'd37126, 16'd37672, 16'd46142, 16'd14748, 16'd12653, 16'd63064, 16'd5991, 16'd60440, 16'd19977, 16'd55788});
	test_expansion(128'h3c1526cb30a4dc180994bb064f22e522, {16'd55750, 16'd2621, 16'd49848, 16'd63015, 16'd50684, 16'd50939, 16'd51421, 16'd55545, 16'd31270, 16'd13144, 16'd44547, 16'd46114, 16'd18786, 16'd29309, 16'd16396, 16'd29545, 16'd47613, 16'd27353, 16'd6255, 16'd13608, 16'd35871, 16'd3313, 16'd59327, 16'd29320, 16'd64281, 16'd15604});
	test_expansion(128'hbe17adb3944db9096567b70dace435ae, {16'd1266, 16'd36943, 16'd54156, 16'd64966, 16'd11719, 16'd58287, 16'd27729, 16'd35896, 16'd23751, 16'd59884, 16'd2197, 16'd32427, 16'd24667, 16'd31786, 16'd12369, 16'd9934, 16'd44660, 16'd32728, 16'd16489, 16'd2473, 16'd13121, 16'd59478, 16'd58372, 16'd3550, 16'd51382, 16'd18944});
	test_expansion(128'h53df5b64fa44e075181d02fedae0e416, {16'd10611, 16'd37717, 16'd57939, 16'd38870, 16'd35204, 16'd8853, 16'd4066, 16'd7984, 16'd40754, 16'd35214, 16'd2012, 16'd43620, 16'd20164, 16'd55203, 16'd3928, 16'd29771, 16'd21595, 16'd50194, 16'd41974, 16'd61028, 16'd19903, 16'd64306, 16'd61988, 16'd64667, 16'd4537, 16'd31719});
	test_expansion(128'h401033bfffaf56cf2f0028019c0d7eb6, {16'd52753, 16'd2020, 16'd47495, 16'd29198, 16'd47906, 16'd14383, 16'd55763, 16'd43453, 16'd42679, 16'd26273, 16'd45604, 16'd64436, 16'd48134, 16'd11454, 16'd34912, 16'd40208, 16'd14468, 16'd5190, 16'd43606, 16'd13907, 16'd37449, 16'd13381, 16'd65374, 16'd47529, 16'd36343, 16'd22072});
	test_expansion(128'h128f0d8a0e93ff6fba442e3a5836f197, {16'd6084, 16'd7449, 16'd41941, 16'd59435, 16'd25415, 16'd60651, 16'd62028, 16'd11084, 16'd558, 16'd36481, 16'd44217, 16'd4929, 16'd60479, 16'd59747, 16'd53882, 16'd64324, 16'd55554, 16'd46629, 16'd7787, 16'd8958, 16'd22667, 16'd64542, 16'd5418, 16'd35947, 16'd42089, 16'd26006});
	test_expansion(128'hce4c70abacb080e20d2ddb76514af35b, {16'd53917, 16'd10332, 16'd4544, 16'd9171, 16'd9287, 16'd53283, 16'd38812, 16'd27846, 16'd27296, 16'd10242, 16'd4563, 16'd32239, 16'd17974, 16'd44640, 16'd6418, 16'd15493, 16'd45426, 16'd49136, 16'd49256, 16'd15713, 16'd36833, 16'd8957, 16'd62706, 16'd2846, 16'd39230, 16'd12928});
	test_expansion(128'hae244f867d7ed00f73f38fa61ad4552f, {16'd8606, 16'd56350, 16'd33312, 16'd27330, 16'd32498, 16'd6117, 16'd27168, 16'd56894, 16'd14264, 16'd53107, 16'd45702, 16'd34895, 16'd55835, 16'd17860, 16'd45823, 16'd7201, 16'd27904, 16'd36656, 16'd62726, 16'd47244, 16'd32590, 16'd20903, 16'd47255, 16'd17255, 16'd1632, 16'd40219});
	test_expansion(128'he4d099f02fda27adad5b99ef424872ff, {16'd15794, 16'd45675, 16'd60914, 16'd55717, 16'd33527, 16'd35856, 16'd9743, 16'd13592, 16'd48371, 16'd31754, 16'd10061, 16'd5768, 16'd53114, 16'd39912, 16'd51297, 16'd51529, 16'd48924, 16'd64630, 16'd61167, 16'd62799, 16'd25789, 16'd18043, 16'd51790, 16'd14905, 16'd16530, 16'd10707});
	test_expansion(128'hcd0b09ed7d76619b2413cba334967610, {16'd11379, 16'd35217, 16'd48738, 16'd35900, 16'd27116, 16'd33201, 16'd8398, 16'd42472, 16'd61435, 16'd51730, 16'd49129, 16'd60641, 16'd23275, 16'd40922, 16'd1182, 16'd6721, 16'd441, 16'd51593, 16'd46508, 16'd31696, 16'd57609, 16'd22722, 16'd2884, 16'd43621, 16'd21830, 16'd61616});
	test_expansion(128'h745861a5eaf505943cdf5293ad3ed5cf, {16'd12674, 16'd9190, 16'd14490, 16'd49443, 16'd29143, 16'd27657, 16'd39514, 16'd57147, 16'd33072, 16'd7010, 16'd4884, 16'd38860, 16'd25676, 16'd38585, 16'd25034, 16'd58940, 16'd31872, 16'd24835, 16'd33886, 16'd45427, 16'd17475, 16'd57388, 16'd55398, 16'd1867, 16'd23358, 16'd49245});
	test_expansion(128'h309d5eb9db7314285a448a6152364468, {16'd56483, 16'd26970, 16'd43197, 16'd57304, 16'd18749, 16'd19809, 16'd44205, 16'd4543, 16'd55648, 16'd58466, 16'd51466, 16'd1850, 16'd33762, 16'd20474, 16'd62620, 16'd8088, 16'd6659, 16'd9182, 16'd52545, 16'd37064, 16'd39689, 16'd23695, 16'd37165, 16'd28637, 16'd14933, 16'd25057});
	test_expansion(128'h7889f1214ae40df9d4bcfa02829fbb64, {16'd9229, 16'd55740, 16'd10028, 16'd60595, 16'd3737, 16'd16182, 16'd22577, 16'd14130, 16'd29455, 16'd11192, 16'd8444, 16'd10849, 16'd43225, 16'd12754, 16'd63157, 16'd20834, 16'd27859, 16'd60740, 16'd33316, 16'd55080, 16'd27462, 16'd55693, 16'd31572, 16'd2301, 16'd58033, 16'd63135});
	test_expansion(128'h344fa849ff466722768274f93374e5da, {16'd25560, 16'd30218, 16'd45221, 16'd33909, 16'd12006, 16'd60224, 16'd43425, 16'd7840, 16'd23286, 16'd57649, 16'd51596, 16'd43082, 16'd42822, 16'd35075, 16'd56463, 16'd56461, 16'd16669, 16'd13267, 16'd26129, 16'd4880, 16'd6730, 16'd61510, 16'd14597, 16'd55468, 16'd35221, 16'd9868});
	test_expansion(128'h2aea46e0f1d785e2b00e2f887678e748, {16'd16682, 16'd738, 16'd29838, 16'd29238, 16'd58978, 16'd59600, 16'd40864, 16'd63664, 16'd47306, 16'd45986, 16'd14971, 16'd52793, 16'd1055, 16'd62992, 16'd47975, 16'd29067, 16'd7566, 16'd42506, 16'd35931, 16'd18802, 16'd36113, 16'd5746, 16'd13880, 16'd20885, 16'd63683, 16'd21494});
	test_expansion(128'h9a1ce72202facc37190df0ae98917113, {16'd30398, 16'd53536, 16'd16103, 16'd45727, 16'd5632, 16'd6974, 16'd51252, 16'd38200, 16'd65094, 16'd56818, 16'd35735, 16'd2451, 16'd19461, 16'd16780, 16'd17023, 16'd4720, 16'd59184, 16'd2378, 16'd62955, 16'd1504, 16'd22997, 16'd39566, 16'd20578, 16'd17964, 16'd46078, 16'd48912});
	test_expansion(128'hcef1d408126cbddfad7c03db80826a4b, {16'd65171, 16'd12531, 16'd31224, 16'd15923, 16'd106, 16'd34107, 16'd19968, 16'd3508, 16'd35323, 16'd6262, 16'd27583, 16'd63955, 16'd36367, 16'd53846, 16'd39628, 16'd45071, 16'd18366, 16'd60576, 16'd53993, 16'd22326, 16'd8469, 16'd13994, 16'd15626, 16'd16049, 16'd16856, 16'd61655});
	test_expansion(128'hc1069ac05d1664aaddc2e7c583a304f5, {16'd26309, 16'd4093, 16'd44551, 16'd43245, 16'd29137, 16'd53698, 16'd57500, 16'd44754, 16'd53357, 16'd46760, 16'd14041, 16'd16214, 16'd61721, 16'd9561, 16'd39645, 16'd45840, 16'd11979, 16'd40090, 16'd14139, 16'd47621, 16'd51018, 16'd45542, 16'd17753, 16'd65225, 16'd32470, 16'd61655});
	test_expansion(128'h54c8bc20b1f377ebe1b8a4bba6217d60, {16'd19962, 16'd456, 16'd61511, 16'd19752, 16'd37273, 16'd8376, 16'd4220, 16'd52668, 16'd27549, 16'd49892, 16'd48614, 16'd59524, 16'd52030, 16'd9683, 16'd62886, 16'd10058, 16'd23162, 16'd62649, 16'd29304, 16'd39647, 16'd55642, 16'd45757, 16'd53766, 16'd55336, 16'd29689, 16'd63289});
	test_expansion(128'hed474e0783072547bd99d30ccfa146e5, {16'd52770, 16'd27896, 16'd59284, 16'd62079, 16'd14579, 16'd14183, 16'd3042, 16'd46451, 16'd8923, 16'd10318, 16'd42589, 16'd12017, 16'd910, 16'd7865, 16'd18197, 16'd12647, 16'd26261, 16'd57447, 16'd57097, 16'd38610, 16'd990, 16'd58504, 16'd59866, 16'd27436, 16'd53460, 16'd46481});
	test_expansion(128'hef212b5701e386822d8ed52ee836ace2, {16'd57711, 16'd2881, 16'd45917, 16'd18656, 16'd29510, 16'd18819, 16'd61093, 16'd55153, 16'd45306, 16'd31512, 16'd63328, 16'd48992, 16'd37263, 16'd14992, 16'd17447, 16'd13197, 16'd32550, 16'd8277, 16'd57684, 16'd64428, 16'd9498, 16'd52695, 16'd29896, 16'd55841, 16'd49758, 16'd33951});
	test_expansion(128'h606ab358f29856145fa31b321f732f44, {16'd63814, 16'd26958, 16'd3127, 16'd47245, 16'd56774, 16'd51157, 16'd53962, 16'd33812, 16'd55811, 16'd3305, 16'd5020, 16'd56811, 16'd33064, 16'd39756, 16'd20776, 16'd30249, 16'd17394, 16'd32054, 16'd15918, 16'd27786, 16'd33642, 16'd9228, 16'd19596, 16'd22937, 16'd16032, 16'd33962});
	test_expansion(128'h08ac0a19daed47e9cc527f3925e55eb5, {16'd55648, 16'd2371, 16'd3231, 16'd46535, 16'd36177, 16'd1061, 16'd5382, 16'd18875, 16'd10688, 16'd53330, 16'd33575, 16'd7793, 16'd55624, 16'd13795, 16'd52667, 16'd56702, 16'd16233, 16'd12714, 16'd23266, 16'd18591, 16'd26572, 16'd53767, 16'd58001, 16'd54263, 16'd47888, 16'd9191});
	test_expansion(128'h65b543a43af6dff1d9603584462ae3d9, {16'd61824, 16'd9150, 16'd58540, 16'd34141, 16'd26767, 16'd19920, 16'd14229, 16'd61512, 16'd32464, 16'd4374, 16'd57798, 16'd54670, 16'd14213, 16'd31428, 16'd26180, 16'd46660, 16'd33433, 16'd1657, 16'd35221, 16'd42671, 16'd63929, 16'd34138, 16'd51014, 16'd39144, 16'd4462, 16'd22971});
	test_expansion(128'h87c2a6633347787702de0c251ddcee57, {16'd34471, 16'd50592, 16'd65329, 16'd13166, 16'd37804, 16'd49030, 16'd61947, 16'd60974, 16'd9179, 16'd62088, 16'd48811, 16'd94, 16'd18198, 16'd15465, 16'd36269, 16'd23810, 16'd34662, 16'd30877, 16'd14326, 16'd1507, 16'd50730, 16'd22067, 16'd19568, 16'd43767, 16'd59192, 16'd39180});
	test_expansion(128'h1d58e08fb715edd1af31f2d1ad97643b, {16'd52972, 16'd57810, 16'd63112, 16'd63119, 16'd3751, 16'd26422, 16'd22049, 16'd12532, 16'd41714, 16'd43199, 16'd45401, 16'd2892, 16'd54342, 16'd3423, 16'd2663, 16'd26831, 16'd64016, 16'd3913, 16'd38691, 16'd2827, 16'd4244, 16'd16047, 16'd22716, 16'd31963, 16'd35575, 16'd39336});
	test_expansion(128'hc3d954b2dad0cc8e9debd4a2ebdb5089, {16'd45853, 16'd1904, 16'd3950, 16'd12476, 16'd3361, 16'd48918, 16'd54425, 16'd43481, 16'd45082, 16'd50131, 16'd17703, 16'd1560, 16'd51155, 16'd38288, 16'd6803, 16'd23334, 16'd39866, 16'd63351, 16'd35264, 16'd41832, 16'd45653, 16'd50690, 16'd4407, 16'd53555, 16'd3137, 16'd14482});
	test_expansion(128'h6d44f0c99631796bd3fadc0b3a7bf05f, {16'd57553, 16'd6267, 16'd32236, 16'd65268, 16'd60803, 16'd63945, 16'd27264, 16'd16626, 16'd47182, 16'd54100, 16'd2748, 16'd54391, 16'd36559, 16'd52880, 16'd36227, 16'd40962, 16'd51475, 16'd36943, 16'd53826, 16'd32824, 16'd44094, 16'd27402, 16'd2541, 16'd37765, 16'd9662, 16'd32677});
	test_expansion(128'hbeff9f16fa2fae3ba1c5dc0fc4734a9d, {16'd50978, 16'd40659, 16'd13326, 16'd45707, 16'd61168, 16'd47209, 16'd59928, 16'd13458, 16'd13337, 16'd18607, 16'd29914, 16'd24157, 16'd54008, 16'd20287, 16'd27533, 16'd26992, 16'd6356, 16'd38995, 16'd992, 16'd31715, 16'd53701, 16'd6920, 16'd35942, 16'd62846, 16'd11514, 16'd35028});
	test_expansion(128'h24976a0c86320f8a0f5dc507a4cc80f2, {16'd51440, 16'd49943, 16'd22189, 16'd50636, 16'd35070, 16'd49860, 16'd32, 16'd55397, 16'd13001, 16'd43606, 16'd33444, 16'd9222, 16'd40261, 16'd42859, 16'd41135, 16'd51170, 16'd55659, 16'd38138, 16'd4231, 16'd9926, 16'd33512, 16'd46002, 16'd13280, 16'd25537, 16'd1021, 16'd26091});
	test_expansion(128'h8c86bfcc9484de2c3161dd4d4e0c3363, {16'd51846, 16'd64042, 16'd17410, 16'd34702, 16'd54338, 16'd50210, 16'd59664, 16'd54275, 16'd4293, 16'd58377, 16'd42060, 16'd5443, 16'd57690, 16'd24187, 16'd43685, 16'd64210, 16'd22617, 16'd2893, 16'd15073, 16'd39921, 16'd46642, 16'd9886, 16'd6633, 16'd25188, 16'd58646, 16'd9970});
	test_expansion(128'h33bc0164bbf0e94457d4a5406e811c76, {16'd75, 16'd63476, 16'd30873, 16'd65300, 16'd9940, 16'd17663, 16'd27992, 16'd2242, 16'd24664, 16'd42031, 16'd61498, 16'd6699, 16'd16502, 16'd24864, 16'd2433, 16'd42349, 16'd3532, 16'd9614, 16'd49537, 16'd16419, 16'd39925, 16'd26781, 16'd61208, 16'd55967, 16'd63906, 16'd41011});
	test_expansion(128'h0ecf124e942b1c15e5b05ec9207a7f9f, {16'd52438, 16'd24323, 16'd58786, 16'd12695, 16'd9285, 16'd27703, 16'd15265, 16'd13569, 16'd57206, 16'd23130, 16'd69, 16'd10729, 16'd52759, 16'd49142, 16'd42315, 16'd45196, 16'd62378, 16'd36221, 16'd16711, 16'd45467, 16'd36266, 16'd30348, 16'd8544, 16'd21080, 16'd55424, 16'd56807});
	test_expansion(128'hb85f9aa384b40eaf06b5cf8d585f76b0, {16'd28424, 16'd3435, 16'd63068, 16'd59023, 16'd57169, 16'd877, 16'd27106, 16'd20005, 16'd52388, 16'd45352, 16'd54500, 16'd24577, 16'd44115, 16'd16655, 16'd20267, 16'd39738, 16'd56582, 16'd58817, 16'd6454, 16'd45364, 16'd19024, 16'd8740, 16'd39498, 16'd45831, 16'd24590, 16'd32276});
	test_expansion(128'h35bc38480fdf2e1279d298b0ff03ac9f, {16'd37867, 16'd33552, 16'd60383, 16'd51626, 16'd2692, 16'd22423, 16'd44859, 16'd26247, 16'd59668, 16'd9535, 16'd61622, 16'd16862, 16'd22778, 16'd39649, 16'd40760, 16'd61978, 16'd9402, 16'd44570, 16'd62586, 16'd10945, 16'd18367, 16'd63494, 16'd966, 16'd50013, 16'd11251, 16'd7873});
	test_expansion(128'hd7310361e9902204f9282ce0a618a3de, {16'd35528, 16'd56149, 16'd41017, 16'd61399, 16'd54716, 16'd8761, 16'd38114, 16'd38474, 16'd42906, 16'd44274, 16'd43682, 16'd2756, 16'd48714, 16'd9800, 16'd8445, 16'd34552, 16'd26147, 16'd59299, 16'd58794, 16'd24503, 16'd21907, 16'd64873, 16'd51282, 16'd16692, 16'd21089, 16'd13116});
	test_expansion(128'he3db3b4d0dfb60e39a77d39b28e5efa6, {16'd16138, 16'd46338, 16'd40514, 16'd14272, 16'd50646, 16'd35872, 16'd41302, 16'd43558, 16'd56013, 16'd12758, 16'd13539, 16'd3348, 16'd43312, 16'd51091, 16'd37247, 16'd28852, 16'd51962, 16'd36380, 16'd22561, 16'd60563, 16'd14671, 16'd53478, 16'd16820, 16'd43434, 16'd35177, 16'd28281});
	test_expansion(128'hecedc595433c509c52a4cd8ec59fd139, {16'd56211, 16'd3938, 16'd8148, 16'd5821, 16'd52370, 16'd31281, 16'd64826, 16'd45968, 16'd45348, 16'd42163, 16'd27101, 16'd61534, 16'd57069, 16'd35787, 16'd5353, 16'd34280, 16'd31682, 16'd7079, 16'd7008, 16'd33992, 16'd8266, 16'd42437, 16'd41259, 16'd13676, 16'd55655, 16'd40128});
	test_expansion(128'h0ca406ea8a1d78069a9ff3a5390a045f, {16'd23794, 16'd8444, 16'd42334, 16'd38255, 16'd62052, 16'd55538, 16'd19445, 16'd22057, 16'd13079, 16'd60849, 16'd29733, 16'd22494, 16'd14291, 16'd6023, 16'd26786, 16'd21321, 16'd33737, 16'd32226, 16'd3353, 16'd47411, 16'd28721, 16'd9911, 16'd62149, 16'd51715, 16'd30142, 16'd32459});
	test_expansion(128'hf4eda61903cde5c2a021d78e1a876e9f, {16'd39432, 16'd64232, 16'd38676, 16'd42175, 16'd42443, 16'd20261, 16'd59825, 16'd52057, 16'd51137, 16'd24420, 16'd65031, 16'd12072, 16'd47043, 16'd64567, 16'd46508, 16'd1836, 16'd47500, 16'd55688, 16'd24264, 16'd48703, 16'd61240, 16'd16168, 16'd25919, 16'd43619, 16'd18368, 16'd32183});
	test_expansion(128'hea19cffb713d2b021effb03d1e61ce73, {16'd63046, 16'd63014, 16'd42629, 16'd53477, 16'd32530, 16'd33657, 16'd33787, 16'd42032, 16'd14690, 16'd57659, 16'd51953, 16'd49421, 16'd47521, 16'd22275, 16'd33248, 16'd47999, 16'd41414, 16'd9742, 16'd43497, 16'd22638, 16'd43510, 16'd58833, 16'd58499, 16'd46028, 16'd42393, 16'd44592});
	test_expansion(128'h9f04f2fcbe24f56787c8b3fca7cca4a8, {16'd12088, 16'd24987, 16'd59230, 16'd40400, 16'd24134, 16'd29776, 16'd49008, 16'd29026, 16'd24303, 16'd60187, 16'd5148, 16'd56638, 16'd41161, 16'd36839, 16'd64724, 16'd34602, 16'd47443, 16'd19143, 16'd24130, 16'd41898, 16'd18780, 16'd39410, 16'd64288, 16'd65450, 16'd17804, 16'd60064});
	test_expansion(128'hc2e1d3d29544a6f8ca78e2ec531aec34, {16'd23838, 16'd64562, 16'd60843, 16'd6925, 16'd27912, 16'd49595, 16'd21981, 16'd60544, 16'd51098, 16'd45108, 16'd54738, 16'd47737, 16'd59946, 16'd30412, 16'd64384, 16'd30150, 16'd27130, 16'd46626, 16'd49926, 16'd4263, 16'd34567, 16'd34028, 16'd8814, 16'd7073, 16'd6829, 16'd29267});
	test_expansion(128'h7534ddaac8ab985430297b9f592103a8, {16'd2371, 16'd46181, 16'd33214, 16'd5874, 16'd13695, 16'd8861, 16'd9223, 16'd64514, 16'd16683, 16'd18944, 16'd50714, 16'd31931, 16'd30759, 16'd65462, 16'd2517, 16'd53600, 16'd10121, 16'd39465, 16'd60272, 16'd22787, 16'd49410, 16'd33701, 16'd48921, 16'd55951, 16'd23527, 16'd33203});
	test_expansion(128'h4eec1b28342a16d4e15352dc6b6664b6, {16'd49652, 16'd44087, 16'd58977, 16'd19102, 16'd54733, 16'd11256, 16'd47700, 16'd4324, 16'd37099, 16'd63512, 16'd6456, 16'd24255, 16'd39473, 16'd28375, 16'd65048, 16'd39383, 16'd61719, 16'd18155, 16'd61432, 16'd19968, 16'd14564, 16'd71, 16'd1567, 16'd40571, 16'd15654, 16'd48144});
	test_expansion(128'h084bab2f88fcd4f5637213534342d360, {16'd54543, 16'd43631, 16'd33650, 16'd58514, 16'd51952, 16'd38982, 16'd65093, 16'd41243, 16'd48440, 16'd17145, 16'd58715, 16'd44018, 16'd27936, 16'd47158, 16'd3338, 16'd21954, 16'd32456, 16'd18095, 16'd14742, 16'd9848, 16'd43594, 16'd36512, 16'd20689, 16'd31421, 16'd28369, 16'd52729});
	test_expansion(128'hfca7269527e6328ed9e58f5d4a7e57c3, {16'd39028, 16'd61736, 16'd63826, 16'd49995, 16'd54830, 16'd61304, 16'd60390, 16'd36602, 16'd26842, 16'd51359, 16'd4191, 16'd60079, 16'd47749, 16'd47741, 16'd61024, 16'd19636, 16'd57824, 16'd47452, 16'd53305, 16'd46737, 16'd33758, 16'd9715, 16'd1681, 16'd17839, 16'd11079, 16'd49995});
	test_expansion(128'ha37a554d4b57d0a8987809e77ccec064, {16'd2989, 16'd36917, 16'd24579, 16'd4605, 16'd43736, 16'd59828, 16'd29487, 16'd6897, 16'd34111, 16'd15272, 16'd21770, 16'd10676, 16'd44808, 16'd51660, 16'd29118, 16'd62225, 16'd15635, 16'd24036, 16'd5998, 16'd19269, 16'd46727, 16'd18346, 16'd52736, 16'd19442, 16'd6471, 16'd38078});
	test_expansion(128'h977edfe7c111d4a17e92a3f037dc1cb6, {16'd32793, 16'd5643, 16'd58816, 16'd199, 16'd12942, 16'd35905, 16'd872, 16'd59506, 16'd52748, 16'd13431, 16'd16545, 16'd24918, 16'd11734, 16'd34186, 16'd58456, 16'd41125, 16'd55177, 16'd693, 16'd64858, 16'd61156, 16'd58217, 16'd14329, 16'd59383, 16'd41776, 16'd23832, 16'd18426});
	test_expansion(128'h3bf0dd40415391c2984f7954931ad83e, {16'd48987, 16'd6403, 16'd61960, 16'd5285, 16'd60715, 16'd47516, 16'd56218, 16'd11807, 16'd40719, 16'd48183, 16'd39351, 16'd12034, 16'd56035, 16'd5295, 16'd34794, 16'd31395, 16'd42848, 16'd54954, 16'd25189, 16'd29241, 16'd55829, 16'd43165, 16'd40045, 16'd15628, 16'd40615, 16'd18889});
	test_expansion(128'h558817ca1a4d8073b338d345bc9a78dc, {16'd3721, 16'd60977, 16'd41314, 16'd39443, 16'd60388, 16'd26198, 16'd34428, 16'd26105, 16'd19976, 16'd7250, 16'd20770, 16'd19916, 16'd52403, 16'd52540, 16'd21006, 16'd14605, 16'd47646, 16'd45557, 16'd2636, 16'd52610, 16'd19803, 16'd60958, 16'd45719, 16'd16368, 16'd59815, 16'd47133});
	test_expansion(128'hb2bd4001d7080f7111b7b4da2376ec44, {16'd22930, 16'd58938, 16'd10275, 16'd59400, 16'd40260, 16'd3352, 16'd35225, 16'd44791, 16'd27828, 16'd51074, 16'd49756, 16'd14525, 16'd44324, 16'd34605, 16'd41888, 16'd20937, 16'd14195, 16'd12547, 16'd49012, 16'd22438, 16'd42664, 16'd32158, 16'd26007, 16'd7508, 16'd26113, 16'd9052});
	test_expansion(128'h39427c47dd818dd2404f4825325cb9aa, {16'd10904, 16'd36591, 16'd18799, 16'd11630, 16'd8937, 16'd39067, 16'd33974, 16'd48305, 16'd43957, 16'd23105, 16'd1409, 16'd31517, 16'd57385, 16'd42621, 16'd3000, 16'd24547, 16'd14926, 16'd46978, 16'd19381, 16'd59785, 16'd6, 16'd38660, 16'd5965, 16'd18080, 16'd25298, 16'd85});
	test_expansion(128'hb87e5987a0bbcc1a72c685f15891f96a, {16'd51552, 16'd55422, 16'd49663, 16'd59866, 16'd48379, 16'd9238, 16'd16613, 16'd45718, 16'd20279, 16'd64118, 16'd11578, 16'd26159, 16'd14024, 16'd9135, 16'd10724, 16'd49712, 16'd56338, 16'd10493, 16'd11834, 16'd46878, 16'd45101, 16'd26, 16'd11025, 16'd4052, 16'd39332, 16'd19983});
	test_expansion(128'hb66a7f7d4e6ef50ba2a554fbcd60e1fb, {16'd28657, 16'd42301, 16'd25649, 16'd30625, 16'd8910, 16'd54786, 16'd39546, 16'd58885, 16'd30357, 16'd30191, 16'd48785, 16'd15592, 16'd12592, 16'd56096, 16'd50251, 16'd7924, 16'd19029, 16'd17163, 16'd64703, 16'd6216, 16'd10823, 16'd33985, 16'd16147, 16'd18871, 16'd18582, 16'd23601});
	test_expansion(128'h9b39c99eecbab679b55ba8723eadf33a, {16'd26872, 16'd5683, 16'd2264, 16'd57145, 16'd443, 16'd33509, 16'd18659, 16'd18574, 16'd49886, 16'd36868, 16'd21575, 16'd9270, 16'd51058, 16'd29440, 16'd18617, 16'd48184, 16'd7010, 16'd46831, 16'd16470, 16'd42235, 16'd16408, 16'd59643, 16'd23055, 16'd15524, 16'd1129, 16'd63945});
	test_expansion(128'h7fbd093ef7a9689dfe768d7b9e4cd381, {16'd26316, 16'd10021, 16'd27211, 16'd11330, 16'd54795, 16'd23447, 16'd59026, 16'd37672, 16'd39298, 16'd49364, 16'd108, 16'd64954, 16'd28312, 16'd14005, 16'd63890, 16'd64065, 16'd2868, 16'd14848, 16'd2845, 16'd30711, 16'd18997, 16'd41286, 16'd38463, 16'd11309, 16'd57587, 16'd59258});
	test_expansion(128'h3019f43ec4919b76e122e48ba27b085a, {16'd55263, 16'd11068, 16'd32981, 16'd38731, 16'd26086, 16'd27497, 16'd19625, 16'd33388, 16'd17139, 16'd21398, 16'd2549, 16'd20180, 16'd62101, 16'd12874, 16'd53099, 16'd32272, 16'd9431, 16'd50192, 16'd37672, 16'd26332, 16'd58205, 16'd17603, 16'd24269, 16'd9617, 16'd35262, 16'd1775});
	test_expansion(128'h4ed784ce1401bb214b386f7d9a175b9e, {16'd42926, 16'd22091, 16'd51135, 16'd55727, 16'd23063, 16'd62502, 16'd47658, 16'd50317, 16'd10539, 16'd46971, 16'd16802, 16'd51925, 16'd16590, 16'd27802, 16'd11456, 16'd47430, 16'd18611, 16'd15733, 16'd26907, 16'd52123, 16'd3774, 16'd22361, 16'd2954, 16'd27055, 16'd28490, 16'd2152});
	test_expansion(128'h66e0d52f1672c9bccc773ba4444a30b0, {16'd63712, 16'd3726, 16'd29500, 16'd5572, 16'd23827, 16'd58776, 16'd30948, 16'd55898, 16'd55960, 16'd8750, 16'd40043, 16'd44925, 16'd16996, 16'd53469, 16'd34096, 16'd49304, 16'd58526, 16'd54094, 16'd133, 16'd42927, 16'd28316, 16'd4259, 16'd2026, 16'd23848, 16'd7656, 16'd24905});
	test_expansion(128'hec85af359759cbe5a023fb59424db2cc, {16'd51122, 16'd5497, 16'd52510, 16'd12829, 16'd30321, 16'd58843, 16'd26321, 16'd27422, 16'd21200, 16'd8195, 16'd17738, 16'd44453, 16'd11415, 16'd3902, 16'd31806, 16'd20474, 16'd37549, 16'd55447, 16'd55427, 16'd1223, 16'd44567, 16'd38638, 16'd59740, 16'd4206, 16'd26023, 16'd44473});
	test_expansion(128'he2b914224a53cdc7e77f295a9aa57563, {16'd28552, 16'd55405, 16'd65051, 16'd26377, 16'd16161, 16'd24893, 16'd7023, 16'd3620, 16'd31064, 16'd63035, 16'd30341, 16'd10396, 16'd52804, 16'd31637, 16'd22727, 16'd18906, 16'd15226, 16'd21504, 16'd56624, 16'd58999, 16'd17011, 16'd47580, 16'd54819, 16'd30098, 16'd30010, 16'd21582});
	test_expansion(128'h54f54e079b29741f3b0512e726dcf112, {16'd12722, 16'd9100, 16'd1591, 16'd35610, 16'd43310, 16'd26086, 16'd41903, 16'd26495, 16'd19683, 16'd3942, 16'd48431, 16'd41423, 16'd44489, 16'd5478, 16'd24713, 16'd54928, 16'd60543, 16'd33994, 16'd1925, 16'd6309, 16'd53569, 16'd16973, 16'd28467, 16'd62641, 16'd52295, 16'd52427});
	test_expansion(128'hd9ed1d1117c8952840e10fcf0deb73bd, {16'd30852, 16'd31225, 16'd33279, 16'd60437, 16'd31494, 16'd43541, 16'd43793, 16'd26082, 16'd14224, 16'd1448, 16'd64275, 16'd45220, 16'd7457, 16'd47380, 16'd52879, 16'd64890, 16'd50717, 16'd32503, 16'd35024, 16'd30518, 16'd11385, 16'd21843, 16'd42047, 16'd55299, 16'd23597, 16'd50779});
	test_expansion(128'h6c166d664587099b468aa3cb9c2a17a5, {16'd39339, 16'd3943, 16'd10652, 16'd49064, 16'd52331, 16'd55039, 16'd42375, 16'd29898, 16'd11606, 16'd9191, 16'd47490, 16'd37129, 16'd53395, 16'd51367, 16'd14339, 16'd11223, 16'd20238, 16'd59091, 16'd18226, 16'd21552, 16'd28601, 16'd3409, 16'd48593, 16'd34092, 16'd46588, 16'd5764});
	test_expansion(128'hb44b9752db1527f0ed1dd2571d9328c9, {16'd16677, 16'd27679, 16'd24109, 16'd39172, 16'd56082, 16'd22029, 16'd537, 16'd26425, 16'd32313, 16'd39739, 16'd3330, 16'd52524, 16'd11617, 16'd23462, 16'd9706, 16'd61939, 16'd53209, 16'd39878, 16'd31927, 16'd16872, 16'd14388, 16'd42878, 16'd708, 16'd45278, 16'd62436, 16'd64133});
	test_expansion(128'h255695ba31207b3638542ddc5af607ca, {16'd22238, 16'd36082, 16'd14354, 16'd60653, 16'd8879, 16'd34018, 16'd6869, 16'd35557, 16'd53584, 16'd44057, 16'd35458, 16'd60617, 16'd29525, 16'd28449, 16'd4391, 16'd63280, 16'd49788, 16'd47896, 16'd38565, 16'd3519, 16'd48242, 16'd33248, 16'd43414, 16'd57499, 16'd32427, 16'd51290});
	test_expansion(128'h6805599ebe597f312aa3c7bd84b16552, {16'd56802, 16'd52686, 16'd17561, 16'd31560, 16'd28727, 16'd38761, 16'd64275, 16'd37702, 16'd43713, 16'd3040, 16'd48522, 16'd1814, 16'd33084, 16'd19996, 16'd40289, 16'd42711, 16'd36497, 16'd44888, 16'd31540, 16'd147, 16'd32992, 16'd7103, 16'd16510, 16'd17180, 16'd28532, 16'd61632});
	test_expansion(128'h5a6be17bbb8fa4199fe89e9f84f75633, {16'd29143, 16'd7784, 16'd46232, 16'd975, 16'd10891, 16'd44703, 16'd46663, 16'd44232, 16'd30737, 16'd41103, 16'd11910, 16'd34136, 16'd3381, 16'd36695, 16'd4007, 16'd52774, 16'd1347, 16'd41587, 16'd20569, 16'd33254, 16'd12626, 16'd6993, 16'd23131, 16'd29607, 16'd63356, 16'd4847});
	test_expansion(128'hbb10786aa38982591ccd94fe785cd970, {16'd50808, 16'd64431, 16'd3583, 16'd27014, 16'd60638, 16'd52822, 16'd56144, 16'd19706, 16'd12287, 16'd62901, 16'd17397, 16'd24552, 16'd9346, 16'd12330, 16'd3368, 16'd55808, 16'd31322, 16'd23150, 16'd32281, 16'd40229, 16'd28337, 16'd31611, 16'd31184, 16'd25604, 16'd44861, 16'd63742});
	test_expansion(128'ha71c3b7744e405e2e61be8c81ff805d2, {16'd1962, 16'd28154, 16'd24811, 16'd41495, 16'd14879, 16'd6376, 16'd29856, 16'd17629, 16'd19183, 16'd22804, 16'd2509, 16'd3233, 16'd51937, 16'd16279, 16'd63742, 16'd17119, 16'd45014, 16'd11968, 16'd33253, 16'd49552, 16'd25080, 16'd46918, 16'd28238, 16'd56065, 16'd53788, 16'd15788});
	test_expansion(128'h9aac412d62e413ea51915cd2a54f3e7a, {16'd61641, 16'd14432, 16'd6203, 16'd15329, 16'd42202, 16'd20134, 16'd65532, 16'd16993, 16'd53836, 16'd64697, 16'd3751, 16'd57945, 16'd14527, 16'd15379, 16'd25291, 16'd38683, 16'd21024, 16'd5310, 16'd55386, 16'd11614, 16'd54096, 16'd37113, 16'd29846, 16'd7586, 16'd54954, 16'd45999});
	test_expansion(128'hf0130c0c3c521a1b0eb3c15da1d59017, {16'd23530, 16'd16586, 16'd890, 16'd17730, 16'd46120, 16'd43731, 16'd59148, 16'd38604, 16'd36170, 16'd13253, 16'd19413, 16'd49975, 16'd26581, 16'd21552, 16'd62463, 16'd23435, 16'd26133, 16'd38435, 16'd39185, 16'd56273, 16'd15715, 16'd17173, 16'd13923, 16'd22957, 16'd25220, 16'd19111});
	test_expansion(128'h152919897f6a2ff31943f9255a8e3d8e, {16'd44113, 16'd2736, 16'd62173, 16'd50422, 16'd19133, 16'd61552, 16'd43009, 16'd56579, 16'd33981, 16'd54220, 16'd62068, 16'd12370, 16'd39079, 16'd16078, 16'd18157, 16'd31683, 16'd23569, 16'd36463, 16'd16532, 16'd49992, 16'd659, 16'd44975, 16'd30767, 16'd14390, 16'd47580, 16'd14776});
	test_expansion(128'h7479e96a251fdb35ea9d23b3d327c149, {16'd16153, 16'd59562, 16'd37568, 16'd64120, 16'd32661, 16'd20525, 16'd39524, 16'd58705, 16'd34656, 16'd8174, 16'd13093, 16'd54454, 16'd43725, 16'd44750, 16'd20802, 16'd41855, 16'd23545, 16'd13306, 16'd10041, 16'd39048, 16'd2995, 16'd10463, 16'd42338, 16'd62708, 16'd26325, 16'd18978});
	test_expansion(128'h481f5e9f12b65fcdf2644a28d4377adc, {16'd59349, 16'd44032, 16'd14547, 16'd36382, 16'd35103, 16'd41129, 16'd56385, 16'd31456, 16'd27369, 16'd12702, 16'd57769, 16'd20387, 16'd50363, 16'd39200, 16'd40101, 16'd60012, 16'd9536, 16'd40100, 16'd13305, 16'd6124, 16'd38720, 16'd9546, 16'd26774, 16'd22750, 16'd4440, 16'd7443});
	test_expansion(128'h6b2a198b70da6e8ef98c84824ec01874, {16'd34393, 16'd32874, 16'd34130, 16'd64924, 16'd53991, 16'd23882, 16'd1635, 16'd40351, 16'd23225, 16'd18442, 16'd64533, 16'd14480, 16'd47460, 16'd16219, 16'd36628, 16'd2734, 16'd42313, 16'd29657, 16'd43858, 16'd27065, 16'd8419, 16'd31723, 16'd23154, 16'd15951, 16'd44969, 16'd16091});
	test_expansion(128'h436f1f3973908c0a6cb149af532d5bf0, {16'd34960, 16'd32457, 16'd60536, 16'd29772, 16'd62456, 16'd30828, 16'd38909, 16'd6811, 16'd56572, 16'd28681, 16'd32697, 16'd20321, 16'd12154, 16'd19700, 16'd54002, 16'd59930, 16'd63662, 16'd18305, 16'd62097, 16'd539, 16'd60240, 16'd61686, 16'd32505, 16'd15265, 16'd64402, 16'd22202});
	test_expansion(128'hf96a5b8df3fdf1b7fa73227b979c62e4, {16'd32461, 16'd31345, 16'd60254, 16'd48119, 16'd17783, 16'd31666, 16'd42784, 16'd1911, 16'd49550, 16'd3637, 16'd7017, 16'd20771, 16'd48777, 16'd15877, 16'd16111, 16'd13010, 16'd64930, 16'd41434, 16'd15313, 16'd45063, 16'd17014, 16'd29965, 16'd32974, 16'd13399, 16'd10607, 16'd65298});
	test_expansion(128'h295ccd1f59cc34b2974209dfbd06e2a4, {16'd46242, 16'd3558, 16'd47006, 16'd41336, 16'd48760, 16'd38944, 16'd43196, 16'd17672, 16'd62056, 16'd63756, 16'd45342, 16'd46700, 16'd41001, 16'd18256, 16'd30903, 16'd12098, 16'd9210, 16'd42407, 16'd9657, 16'd64692, 16'd2439, 16'd58411, 16'd57250, 16'd44161, 16'd36226, 16'd28817});
	test_expansion(128'hd7ad3e2173325abe2849298e192d8d9c, {16'd33778, 16'd16527, 16'd6101, 16'd42516, 16'd47114, 16'd9411, 16'd5719, 16'd18457, 16'd32424, 16'd31323, 16'd18344, 16'd41657, 16'd24459, 16'd28464, 16'd41362, 16'd44310, 16'd22303, 16'd31202, 16'd12528, 16'd6906, 16'd20899, 16'd59719, 16'd38410, 16'd1685, 16'd7578, 16'd61527});
	test_expansion(128'h82a3ba20c6798f5835579a4667da8815, {16'd13899, 16'd61056, 16'd39770, 16'd63078, 16'd18648, 16'd62435, 16'd56198, 16'd19402, 16'd682, 16'd5955, 16'd24020, 16'd14138, 16'd6960, 16'd63552, 16'd35228, 16'd4679, 16'd61807, 16'd9406, 16'd43826, 16'd45896, 16'd50690, 16'd10134, 16'd37719, 16'd10110, 16'd62336, 16'd55223});
	test_expansion(128'h36656312bdacd457a0d975655f522637, {16'd64813, 16'd48912, 16'd37925, 16'd34109, 16'd43438, 16'd63425, 16'd28252, 16'd53516, 16'd18920, 16'd51731, 16'd63829, 16'd61111, 16'd24926, 16'd45108, 16'd17476, 16'd24521, 16'd18099, 16'd61425, 16'd1493, 16'd5146, 16'd43888, 16'd24772, 16'd64855, 16'd21950, 16'd14487, 16'd480});
	test_expansion(128'h83358c4f0082304ce62f7423b8037193, {16'd14810, 16'd42799, 16'd58600, 16'd18501, 16'd6475, 16'd14663, 16'd38517, 16'd57707, 16'd48915, 16'd46559, 16'd38615, 16'd47753, 16'd23277, 16'd33996, 16'd11779, 16'd43601, 16'd62790, 16'd514, 16'd54621, 16'd51268, 16'd30318, 16'd13550, 16'd59413, 16'd34673, 16'd18777, 16'd42283});
	test_expansion(128'h928a7e134757d91117b2ebbba164335a, {16'd32047, 16'd43638, 16'd2418, 16'd44440, 16'd2521, 16'd21326, 16'd16434, 16'd8230, 16'd30302, 16'd32755, 16'd14404, 16'd27012, 16'd58955, 16'd39833, 16'd32263, 16'd31694, 16'd41770, 16'd58649, 16'd61237, 16'd56610, 16'd58107, 16'd50925, 16'd13059, 16'd11458, 16'd45557, 16'd10180});
	test_expansion(128'h9f2f8ae9e2946271688b6a67707b46b6, {16'd61014, 16'd53147, 16'd40052, 16'd4185, 16'd8398, 16'd8440, 16'd2227, 16'd37448, 16'd43711, 16'd65184, 16'd18254, 16'd22928, 16'd51498, 16'd26292, 16'd34163, 16'd19358, 16'd56774, 16'd9064, 16'd60075, 16'd57227, 16'd32044, 16'd4108, 16'd33269, 16'd21375, 16'd45284, 16'd6802});
	test_expansion(128'h2ca6cba2ebdce573662d6bb7450771a9, {16'd4246, 16'd32161, 16'd43225, 16'd41316, 16'd63084, 16'd49660, 16'd62864, 16'd242, 16'd30474, 16'd39802, 16'd37602, 16'd35618, 16'd23998, 16'd53035, 16'd32461, 16'd37491, 16'd4437, 16'd2589, 16'd58186, 16'd56899, 16'd62088, 16'd51485, 16'd61538, 16'd47216, 16'd6694, 16'd54372});
	test_expansion(128'h7e2c4dd0ca2e26bd136e7330f001ef58, {16'd28146, 16'd16340, 16'd41014, 16'd22902, 16'd28567, 16'd28921, 16'd5898, 16'd47059, 16'd25297, 16'd4163, 16'd9647, 16'd7125, 16'd19573, 16'd60670, 16'd8749, 16'd63238, 16'd9766, 16'd57383, 16'd36851, 16'd58014, 16'd62051, 16'd50658, 16'd11783, 16'd50412, 16'd50010, 16'd24932});
	test_expansion(128'h3e32cf25863a2f9e1290b0bb19035b11, {16'd53167, 16'd18567, 16'd12263, 16'd8939, 16'd43885, 16'd11161, 16'd54381, 16'd65089, 16'd33270, 16'd9137, 16'd49097, 16'd46182, 16'd17000, 16'd59182, 16'd53753, 16'd12799, 16'd44019, 16'd28191, 16'd35169, 16'd48020, 16'd23604, 16'd37606, 16'd50055, 16'd31206, 16'd40549, 16'd58136});
	test_expansion(128'hb9bad98bf514cf9a443543b1b86256a1, {16'd50656, 16'd6692, 16'd5383, 16'd45495, 16'd64857, 16'd49120, 16'd29164, 16'd43405, 16'd3373, 16'd28274, 16'd13445, 16'd55631, 16'd10604, 16'd18944, 16'd64571, 16'd48927, 16'd38819, 16'd5752, 16'd23148, 16'd3475, 16'd53017, 16'd17363, 16'd56064, 16'd50397, 16'd34379, 16'd25170});
	test_expansion(128'h6141c7cc06fd1779329e1c63b767a3da, {16'd39758, 16'd34269, 16'd6740, 16'd30649, 16'd57346, 16'd3328, 16'd36485, 16'd951, 16'd55359, 16'd13376, 16'd22827, 16'd21004, 16'd35534, 16'd118, 16'd16888, 16'd60774, 16'd20555, 16'd45811, 16'd47577, 16'd21406, 16'd32634, 16'd11553, 16'd49712, 16'd56714, 16'd58351, 16'd45468});
	test_expansion(128'h12c21e1f94c640b63d7ce30f452956a7, {16'd2649, 16'd36093, 16'd21786, 16'd18809, 16'd4887, 16'd10913, 16'd31958, 16'd36264, 16'd14974, 16'd9572, 16'd11571, 16'd18208, 16'd1107, 16'd28425, 16'd48451, 16'd30230, 16'd8531, 16'd43858, 16'd53135, 16'd46654, 16'd55385, 16'd5464, 16'd9760, 16'd33180, 16'd1205, 16'd24949});
	test_expansion(128'h57f3188973b4eddc1f398a20c678e16d, {16'd14713, 16'd20599, 16'd18579, 16'd28825, 16'd8521, 16'd9973, 16'd50104, 16'd17213, 16'd23566, 16'd20120, 16'd49168, 16'd25534, 16'd535, 16'd42893, 16'd1188, 16'd15070, 16'd59515, 16'd33141, 16'd15338, 16'd53053, 16'd63372, 16'd24598, 16'd58774, 16'd49452, 16'd9903, 16'd14618});
	test_expansion(128'hca1694d104e8df7c9fd0d3a21d663f8f, {16'd29125, 16'd21434, 16'd37793, 16'd59830, 16'd36548, 16'd11446, 16'd6644, 16'd29613, 16'd33100, 16'd34534, 16'd53160, 16'd28281, 16'd2388, 16'd5501, 16'd4875, 16'd32120, 16'd54849, 16'd29243, 16'd46458, 16'd49478, 16'd1849, 16'd56504, 16'd44020, 16'd40813, 16'd11708, 16'd34512});
	test_expansion(128'h0db1eb434ee37fdf038a9f61d24e1aac, {16'd45334, 16'd59882, 16'd53072, 16'd34932, 16'd61963, 16'd8683, 16'd49052, 16'd14332, 16'd58035, 16'd58438, 16'd51334, 16'd48473, 16'd804, 16'd33814, 16'd48491, 16'd29534, 16'd43641, 16'd47099, 16'd31402, 16'd15408, 16'd2814, 16'd47423, 16'd12382, 16'd31086, 16'd50877, 16'd48574});
	test_expansion(128'h596129dbd660faafd96c79753606e818, {16'd10458, 16'd14131, 16'd42297, 16'd32856, 16'd3318, 16'd64515, 16'd48379, 16'd1780, 16'd57330, 16'd25013, 16'd250, 16'd29842, 16'd36330, 16'd55726, 16'd43168, 16'd4246, 16'd38752, 16'd53156, 16'd52614, 16'd57894, 16'd43170, 16'd52004, 16'd40890, 16'd32846, 16'd41174, 16'd46648});
	test_expansion(128'hf7c888f1a35bebcba5bc03f93d5329a3, {16'd14847, 16'd54363, 16'd59201, 16'd15188, 16'd15778, 16'd8050, 16'd27241, 16'd61571, 16'd13378, 16'd4588, 16'd43125, 16'd59098, 16'd43505, 16'd31950, 16'd18336, 16'd47350, 16'd20256, 16'd53743, 16'd61619, 16'd20912, 16'd14761, 16'd63235, 16'd17378, 16'd40535, 16'd38098, 16'd14825});
	test_expansion(128'h94cb8e57d06502a433f6ccd3869d9f5a, {16'd38803, 16'd36046, 16'd5936, 16'd37398, 16'd34848, 16'd41537, 16'd11909, 16'd5708, 16'd2130, 16'd32835, 16'd15726, 16'd32972, 16'd55967, 16'd4857, 16'd62659, 16'd35499, 16'd24669, 16'd36511, 16'd35893, 16'd51984, 16'd62200, 16'd4036, 16'd13043, 16'd58716, 16'd27407, 16'd660});
	test_expansion(128'hc5de47cfb1157c71bf2a82fd44fe3303, {16'd9241, 16'd42266, 16'd39317, 16'd10016, 16'd16176, 16'd31959, 16'd61821, 16'd2049, 16'd10474, 16'd7741, 16'd26293, 16'd30124, 16'd34822, 16'd27407, 16'd34085, 16'd60862, 16'd18194, 16'd63155, 16'd60889, 16'd9685, 16'd65448, 16'd15375, 16'd60892, 16'd26802, 16'd13399, 16'd43039});
	test_expansion(128'h4b78aa1f389d5d220366f840cfbb65e6, {16'd15165, 16'd58875, 16'd52781, 16'd4217, 16'd31398, 16'd46706, 16'd36117, 16'd4819, 16'd23715, 16'd14919, 16'd10922, 16'd30749, 16'd42298, 16'd34023, 16'd21977, 16'd58384, 16'd648, 16'd24047, 16'd20569, 16'd37794, 16'd3643, 16'd31868, 16'd12435, 16'd195, 16'd14823, 16'd11806});
	test_expansion(128'hfdbb03452db9043d6c744b39534cada7, {16'd31059, 16'd37184, 16'd18993, 16'd34648, 16'd36421, 16'd61508, 16'd43506, 16'd56741, 16'd49295, 16'd18239, 16'd39075, 16'd1722, 16'd12554, 16'd55523, 16'd62951, 16'd7269, 16'd21702, 16'd57514, 16'd13510, 16'd57391, 16'd4111, 16'd6133, 16'd39463, 16'd54881, 16'd21427, 16'd39996});
	test_expansion(128'h58cce32054ed41b37bdfa6e411ebc3fc, {16'd61751, 16'd15879, 16'd23886, 16'd63680, 16'd53675, 16'd43468, 16'd13865, 16'd39388, 16'd28959, 16'd18984, 16'd32319, 16'd46843, 16'd22960, 16'd24190, 16'd41009, 16'd52869, 16'd20121, 16'd50491, 16'd28771, 16'd1302, 16'd59538, 16'd55148, 16'd46043, 16'd24082, 16'd63520, 16'd56295});
	test_expansion(128'h7a065b78fd66bfde9b4bebba000a1f36, {16'd11283, 16'd39764, 16'd26790, 16'd40095, 16'd20639, 16'd59711, 16'd59656, 16'd52889, 16'd51833, 16'd18648, 16'd27136, 16'd61891, 16'd41406, 16'd28992, 16'd34441, 16'd64920, 16'd49136, 16'd28564, 16'd44148, 16'd3418, 16'd19074, 16'd12601, 16'd12163, 16'd45195, 16'd1813, 16'd6913});
	test_expansion(128'hec4bf645433edab533b00b44c5e016c4, {16'd62027, 16'd33450, 16'd59447, 16'd48434, 16'd55803, 16'd15794, 16'd17223, 16'd17501, 16'd50652, 16'd28901, 16'd1444, 16'd53556, 16'd32288, 16'd20904, 16'd27643, 16'd23196, 16'd61232, 16'd2073, 16'd24501, 16'd40818, 16'd30816, 16'd10508, 16'd38396, 16'd18976, 16'd59778, 16'd30506});
	test_expansion(128'hb0f4be5d0cd61e04a2015ba89afda191, {16'd54891, 16'd29086, 16'd51397, 16'd50141, 16'd16205, 16'd45580, 16'd3880, 16'd21665, 16'd50282, 16'd51133, 16'd51682, 16'd1894, 16'd28660, 16'd8519, 16'd56902, 16'd51434, 16'd57097, 16'd62172, 16'd4198, 16'd44027, 16'd28204, 16'd5517, 16'd49919, 16'd33507, 16'd12357, 16'd9240});
	test_expansion(128'h57064ec01dc0ea20bc3e61805f8c1fb3, {16'd62311, 16'd15647, 16'd16677, 16'd17766, 16'd41881, 16'd16204, 16'd22208, 16'd59367, 16'd31099, 16'd3985, 16'd23201, 16'd40366, 16'd23129, 16'd42170, 16'd55468, 16'd20165, 16'd34157, 16'd33136, 16'd62800, 16'd29461, 16'd30149, 16'd54441, 16'd21218, 16'd31117, 16'd19547, 16'd18525});
	test_expansion(128'h88e6d1c8418cdfd90c2c374c0901d9d1, {16'd23493, 16'd11416, 16'd45167, 16'd26994, 16'd56466, 16'd64968, 16'd11182, 16'd48801, 16'd33083, 16'd26674, 16'd1183, 16'd46984, 16'd9790, 16'd1955, 16'd6597, 16'd41867, 16'd65433, 16'd12838, 16'd8803, 16'd28840, 16'd11088, 16'd38707, 16'd35208, 16'd8037, 16'd37261, 16'd21021});
	test_expansion(128'he9f7ad8b106f9b6fa684d431babc5b05, {16'd35566, 16'd52471, 16'd14884, 16'd13205, 16'd10755, 16'd35366, 16'd45384, 16'd5065, 16'd9811, 16'd21980, 16'd22023, 16'd14299, 16'd3878, 16'd23375, 16'd4526, 16'd43584, 16'd8113, 16'd25491, 16'd48820, 16'd12832, 16'd48225, 16'd44761, 16'd36294, 16'd51203, 16'd28506, 16'd5374});
	test_expansion(128'hfbe57ed644b6574ccb4bb62a6876143d, {16'd5230, 16'd57041, 16'd13370, 16'd41739, 16'd24993, 16'd16026, 16'd57827, 16'd38226, 16'd27470, 16'd11829, 16'd59419, 16'd44232, 16'd54039, 16'd39986, 16'd65420, 16'd20190, 16'd52033, 16'd8905, 16'd34585, 16'd22949, 16'd60580, 16'd15849, 16'd56227, 16'd58415, 16'd20181, 16'd44311});
	test_expansion(128'h46cff32d7dfe1c512cbb66ff2a479bf6, {16'd65463, 16'd42286, 16'd41059, 16'd33336, 16'd14528, 16'd48220, 16'd5479, 16'd11147, 16'd37770, 16'd20587, 16'd35905, 16'd615, 16'd30583, 16'd17163, 16'd2129, 16'd5599, 16'd43259, 16'd60591, 16'd42905, 16'd35785, 16'd55366, 16'd12383, 16'd8738, 16'd47655, 16'd23638, 16'd39083});
	test_expansion(128'h0cc24e778dfe22f93664d818d35edaa9, {16'd30329, 16'd34894, 16'd48090, 16'd3956, 16'd23424, 16'd51437, 16'd11625, 16'd51051, 16'd61092, 16'd64744, 16'd2454, 16'd45501, 16'd6216, 16'd3882, 16'd3343, 16'd28075, 16'd23242, 16'd15190, 16'd30831, 16'd34668, 16'd702, 16'd7976, 16'd5754, 16'd57213, 16'd18985, 16'd1566});
	test_expansion(128'h92b5390a958b82635e75c49515d3a178, {16'd36142, 16'd4123, 16'd39842, 16'd11080, 16'd35891, 16'd8055, 16'd10083, 16'd1442, 16'd48308, 16'd18700, 16'd41802, 16'd47903, 16'd29320, 16'd40927, 16'd19359, 16'd49538, 16'd51897, 16'd27417, 16'd63960, 16'd5188, 16'd240, 16'd47810, 16'd21930, 16'd17498, 16'd50905, 16'd9485});
	test_expansion(128'h43e4fc2c6a40edd0c60a8676de38c031, {16'd46980, 16'd27011, 16'd55580, 16'd32292, 16'd2229, 16'd2559, 16'd27977, 16'd24498, 16'd10301, 16'd35945, 16'd50851, 16'd55273, 16'd28762, 16'd50928, 16'd37726, 16'd11045, 16'd48321, 16'd64043, 16'd47158, 16'd34463, 16'd15750, 16'd44047, 16'd27849, 16'd9437, 16'd5686, 16'd16947});
	test_expansion(128'ha33e4a86a58687439a518afed33451d6, {16'd24692, 16'd6571, 16'd22613, 16'd52230, 16'd59056, 16'd16975, 16'd65254, 16'd63232, 16'd15038, 16'd7664, 16'd36569, 16'd60616, 16'd19584, 16'd10048, 16'd881, 16'd8858, 16'd55573, 16'd24865, 16'd7612, 16'd23598, 16'd46981, 16'd12931, 16'd38305, 16'd5961, 16'd9509, 16'd26758});
	test_expansion(128'h133e7faeb3d2032f028762c844685a1f, {16'd23089, 16'd14480, 16'd58507, 16'd55669, 16'd15948, 16'd15806, 16'd17132, 16'd23079, 16'd22795, 16'd12139, 16'd53165, 16'd54835, 16'd20658, 16'd35975, 16'd36299, 16'd38069, 16'd41906, 16'd24773, 16'd64604, 16'd62116, 16'd22182, 16'd36046, 16'd20470, 16'd19428, 16'd18279, 16'd24587});
	test_expansion(128'h127c417b08b23e9e5fbcc5c6630db52f, {16'd36515, 16'd60415, 16'd26909, 16'd37573, 16'd36540, 16'd57767, 16'd59270, 16'd37119, 16'd5859, 16'd9990, 16'd9711, 16'd64739, 16'd6979, 16'd11993, 16'd30845, 16'd4432, 16'd82, 16'd32383, 16'd3075, 16'd57682, 16'd46775, 16'd46302, 16'd37567, 16'd1564, 16'd45698, 16'd38965});
	test_expansion(128'hf808852fb6cd470d565d4c2159a3580c, {16'd37166, 16'd12111, 16'd2824, 16'd61447, 16'd51827, 16'd6205, 16'd50341, 16'd40369, 16'd11553, 16'd56167, 16'd16486, 16'd63504, 16'd11491, 16'd50648, 16'd37586, 16'd54448, 16'd14219, 16'd43422, 16'd8967, 16'd35361, 16'd1413, 16'd41625, 16'd35407, 16'd65167, 16'd25235, 16'd13467});
	test_expansion(128'h4a76494f45780efd77264f2eb5e95a0d, {16'd38491, 16'd20407, 16'd35795, 16'd29796, 16'd585, 16'd798, 16'd36843, 16'd18396, 16'd51096, 16'd21540, 16'd62831, 16'd40553, 16'd7852, 16'd3087, 16'd11258, 16'd21267, 16'd47070, 16'd41990, 16'd54532, 16'd51337, 16'd62734, 16'd11702, 16'd23478, 16'd16950, 16'd49288, 16'd32266});
	test_expansion(128'hc8bcc2c0fcb028e2108fa95633e0700c, {16'd53159, 16'd22865, 16'd18291, 16'd39492, 16'd44541, 16'd1028, 16'd28570, 16'd4796, 16'd6800, 16'd38903, 16'd14905, 16'd57901, 16'd8721, 16'd6727, 16'd60243, 16'd50344, 16'd1465, 16'd6577, 16'd561, 16'd18282, 16'd61488, 16'd11405, 16'd55025, 16'd60372, 16'd21680, 16'd35982});
	test_expansion(128'h9268d726c986f3f63f8d71857813f1f0, {16'd22747, 16'd11213, 16'd40421, 16'd59554, 16'd22499, 16'd33924, 16'd48078, 16'd348, 16'd18774, 16'd62573, 16'd61834, 16'd29318, 16'd58491, 16'd47041, 16'd46570, 16'd43800, 16'd57217, 16'd63587, 16'd58184, 16'd19900, 16'd9471, 16'd10106, 16'd4616, 16'd38386, 16'd34956, 16'd61298});
	test_expansion(128'ha1bb9acb21d8b08a7120ac8ca20fae23, {16'd17927, 16'd33117, 16'd54763, 16'd35136, 16'd1726, 16'd35801, 16'd7698, 16'd24683, 16'd31606, 16'd10418, 16'd21898, 16'd51001, 16'd43356, 16'd18718, 16'd525, 16'd21545, 16'd57312, 16'd8063, 16'd29370, 16'd4999, 16'd39541, 16'd46356, 16'd22841, 16'd12940, 16'd22165, 16'd35440});
	test_expansion(128'hbdc6e090bce0371d2c41239f9cf37ed0, {16'd52811, 16'd39725, 16'd597, 16'd25862, 16'd19285, 16'd59526, 16'd28669, 16'd35734, 16'd45712, 16'd24079, 16'd16123, 16'd55529, 16'd42388, 16'd46589, 16'd36060, 16'd33033, 16'd47454, 16'd33315, 16'd546, 16'd60464, 16'd48529, 16'd6675, 16'd25496, 16'd39059, 16'd18187, 16'd6346});
	test_expansion(128'h98ba915853fc108bb477bb429d24278a, {16'd47864, 16'd40469, 16'd52981, 16'd27239, 16'd24708, 16'd20874, 16'd2955, 16'd56570, 16'd429, 16'd47681, 16'd7194, 16'd2517, 16'd49484, 16'd6682, 16'd45263, 16'd50404, 16'd9691, 16'd15539, 16'd38140, 16'd54836, 16'd27710, 16'd41966, 16'd17109, 16'd6222, 16'd10207, 16'd13852});
	test_expansion(128'h4b08cc3ed02eff5d6c5a4871a08bc63a, {16'd38161, 16'd56751, 16'd51846, 16'd60698, 16'd14962, 16'd49557, 16'd14998, 16'd13804, 16'd33164, 16'd16350, 16'd1347, 16'd11107, 16'd46346, 16'd49732, 16'd42754, 16'd62071, 16'd1514, 16'd51015, 16'd64273, 16'd56826, 16'd59662, 16'd846, 16'd13355, 16'd37245, 16'd9719, 16'd44823});
	test_expansion(128'h57d12a7589f4e37a147bf90d65d002e7, {16'd151, 16'd52028, 16'd35544, 16'd6530, 16'd43372, 16'd13376, 16'd25759, 16'd64324, 16'd44911, 16'd59820, 16'd27837, 16'd60386, 16'd9561, 16'd20657, 16'd29690, 16'd35547, 16'd30910, 16'd39505, 16'd62009, 16'd41569, 16'd18812, 16'd45359, 16'd43309, 16'd56621, 16'd9624, 16'd14203});
	test_expansion(128'hee6b5968ca1edaddd52cd95d5ed0799f, {16'd4319, 16'd20958, 16'd34452, 16'd56061, 16'd63927, 16'd8226, 16'd8737, 16'd49143, 16'd8734, 16'd42373, 16'd27806, 16'd2761, 16'd24499, 16'd16683, 16'd26767, 16'd55075, 16'd7557, 16'd7838, 16'd16986, 16'd53428, 16'd36092, 16'd51345, 16'd3010, 16'd5610, 16'd18153, 16'd34800});
	test_expansion(128'h8e097c144d1121278a5512742d28e60e, {16'd1249, 16'd19344, 16'd49384, 16'd41469, 16'd8959, 16'd21286, 16'd55450, 16'd21648, 16'd30068, 16'd33488, 16'd338, 16'd47077, 16'd34604, 16'd43306, 16'd7778, 16'd33787, 16'd10742, 16'd54086, 16'd31030, 16'd17474, 16'd28812, 16'd38785, 16'd25156, 16'd33453, 16'd9701, 16'd30127});
	test_expansion(128'h7a067f155dceed454dc7608ac6aa70fe, {16'd37518, 16'd58350, 16'd13584, 16'd38599, 16'd19424, 16'd47154, 16'd59706, 16'd63113, 16'd13992, 16'd42595, 16'd232, 16'd35385, 16'd35210, 16'd5973, 16'd10354, 16'd60686, 16'd34853, 16'd17029, 16'd14011, 16'd19354, 16'd17022, 16'd50920, 16'd42459, 16'd9761, 16'd58855, 16'd51785});
	test_expansion(128'h109f9a50323ffe4e959ab5c6e9aaee88, {16'd40838, 16'd13423, 16'd33648, 16'd37603, 16'd40010, 16'd39858, 16'd10867, 16'd32940, 16'd5982, 16'd57169, 16'd16660, 16'd36386, 16'd31856, 16'd40304, 16'd52964, 16'd43752, 16'd31146, 16'd20292, 16'd44415, 16'd31550, 16'd2823, 16'd16161, 16'd32251, 16'd55451, 16'd51716, 16'd54213});
	test_expansion(128'h8d7689d003f52b0b50fd14f829128e30, {16'd62812, 16'd13252, 16'd56138, 16'd4700, 16'd48961, 16'd2606, 16'd40304, 16'd19949, 16'd24975, 16'd11733, 16'd33643, 16'd57826, 16'd58846, 16'd60191, 16'd18243, 16'd12174, 16'd35546, 16'd53333, 16'd55213, 16'd31419, 16'd7815, 16'd51814, 16'd54905, 16'd10388, 16'd56271, 16'd6579});
	test_expansion(128'h9d866d5fb44f4ed1140901b69253023b, {16'd21923, 16'd1774, 16'd40383, 16'd11789, 16'd22914, 16'd15346, 16'd49811, 16'd14860, 16'd6409, 16'd32656, 16'd42725, 16'd51251, 16'd57066, 16'd654, 16'd6087, 16'd63028, 16'd36566, 16'd16015, 16'd4485, 16'd6760, 16'd33134, 16'd44679, 16'd11429, 16'd6771, 16'd62060, 16'd36398});
	test_expansion(128'hf4873feb17b23008204b1c2d4a14cf0c, {16'd24336, 16'd31935, 16'd20661, 16'd33202, 16'd15475, 16'd18749, 16'd36473, 16'd24877, 16'd9632, 16'd62511, 16'd42935, 16'd5065, 16'd2541, 16'd17758, 16'd1733, 16'd17974, 16'd21449, 16'd38241, 16'd60048, 16'd57342, 16'd41760, 16'd7005, 16'd8218, 16'd40741, 16'd50606, 16'd2914});
	test_expansion(128'h0100d041aa05c67e1a4cbcbccf1cb20c, {16'd33589, 16'd1435, 16'd14072, 16'd3443, 16'd44794, 16'd37049, 16'd45541, 16'd17566, 16'd3898, 16'd54034, 16'd14124, 16'd14206, 16'd10068, 16'd12166, 16'd46525, 16'd18384, 16'd50971, 16'd18838, 16'd22531, 16'd6114, 16'd48170, 16'd6430, 16'd55514, 16'd52296, 16'd51307, 16'd59934});
	test_expansion(128'hfe751126b3615e16424973015430accc, {16'd55010, 16'd52044, 16'd46647, 16'd61607, 16'd54464, 16'd14505, 16'd4420, 16'd41485, 16'd43892, 16'd64297, 16'd2203, 16'd28173, 16'd9792, 16'd22000, 16'd54852, 16'd53228, 16'd29196, 16'd29991, 16'd35425, 16'd11574, 16'd16525, 16'd47746, 16'd19630, 16'd62781, 16'd51598, 16'd62293});
	test_expansion(128'hdd050c6e300eccda907150c46d237ad3, {16'd7917, 16'd57329, 16'd63382, 16'd39181, 16'd45658, 16'd62688, 16'd7737, 16'd23156, 16'd15917, 16'd8302, 16'd37264, 16'd3639, 16'd39180, 16'd10927, 16'd44648, 16'd24816, 16'd46103, 16'd34717, 16'd43184, 16'd60040, 16'd34251, 16'd55023, 16'd12404, 16'd57717, 16'd36403, 16'd35844});
	test_expansion(128'h3cbe3cd6cbfd24c9d61e5f9b74ab9ef6, {16'd56591, 16'd41863, 16'd52250, 16'd64587, 16'd1491, 16'd3780, 16'd4438, 16'd61742, 16'd12014, 16'd38878, 16'd54082, 16'd40467, 16'd38310, 16'd45749, 16'd4734, 16'd63415, 16'd33348, 16'd28764, 16'd11410, 16'd47683, 16'd59438, 16'd18470, 16'd30930, 16'd33369, 16'd56060, 16'd62974});
	test_expansion(128'h579bad2aa3d7de4c9e3c3982f2842c33, {16'd15242, 16'd39781, 16'd4109, 16'd12206, 16'd12216, 16'd58309, 16'd50065, 16'd39896, 16'd23271, 16'd21661, 16'd8243, 16'd32882, 16'd45639, 16'd20951, 16'd2059, 16'd35817, 16'd43961, 16'd23646, 16'd10264, 16'd11469, 16'd46917, 16'd55518, 16'd22704, 16'd248, 16'd33411, 16'd53807});
	test_expansion(128'h80d9e9fb0e4eb0765aa6fa78b71eab21, {16'd27231, 16'd60418, 16'd17815, 16'd29499, 16'd46643, 16'd36880, 16'd49891, 16'd33719, 16'd27901, 16'd42687, 16'd8247, 16'd38681, 16'd47776, 16'd42026, 16'd63385, 16'd5042, 16'd56190, 16'd43568, 16'd51867, 16'd63114, 16'd22263, 16'd48804, 16'd37483, 16'd55675, 16'd60235, 16'd35200});
	test_expansion(128'hf4d7b9ccfe10f351fa3a79814a8b6fbb, {16'd42629, 16'd2365, 16'd27472, 16'd31379, 16'd29184, 16'd26195, 16'd5860, 16'd5705, 16'd1713, 16'd36913, 16'd26517, 16'd98, 16'd26799, 16'd34329, 16'd25239, 16'd30421, 16'd63766, 16'd17556, 16'd60585, 16'd30160, 16'd44255, 16'd52983, 16'd16542, 16'd844, 16'd22375, 16'd46002});
	test_expansion(128'h56461e8a27be55e901b3ea15cd7cdfe5, {16'd51176, 16'd5769, 16'd61716, 16'd33666, 16'd56059, 16'd39544, 16'd8345, 16'd45801, 16'd53157, 16'd35800, 16'd64440, 16'd18436, 16'd56249, 16'd28642, 16'd26792, 16'd42874, 16'd40404, 16'd50422, 16'd57605, 16'd29373, 16'd19306, 16'd22669, 16'd39132, 16'd20684, 16'd21673, 16'd14238});
	test_expansion(128'h5522a196d225cacded7d6f5e1fa33d7c, {16'd26797, 16'd61121, 16'd17814, 16'd41209, 16'd762, 16'd37280, 16'd42399, 16'd61756, 16'd9967, 16'd13826, 16'd11737, 16'd24987, 16'd57275, 16'd26381, 16'd26097, 16'd52239, 16'd8973, 16'd3830, 16'd46094, 16'd6094, 16'd1999, 16'd11678, 16'd34747, 16'd53972, 16'd21745, 16'd33976});
	test_expansion(128'h09b8005bec2e0aa3887b5692b1af5403, {16'd29111, 16'd34660, 16'd37269, 16'd58445, 16'd21346, 16'd45022, 16'd57253, 16'd29872, 16'd35554, 16'd7875, 16'd33277, 16'd33048, 16'd50415, 16'd30921, 16'd3188, 16'd28592, 16'd23422, 16'd21758, 16'd44851, 16'd35301, 16'd57410, 16'd11006, 16'd30521, 16'd18220, 16'd32830, 16'd9593});
	test_expansion(128'h3e99ac2eb46edb689014a5e8f2131e8c, {16'd64279, 16'd173, 16'd13259, 16'd35313, 16'd6747, 16'd2118, 16'd15615, 16'd50922, 16'd65182, 16'd49939, 16'd32925, 16'd60917, 16'd59648, 16'd37093, 16'd19068, 16'd43367, 16'd36352, 16'd59658, 16'd60577, 16'd33299, 16'd30382, 16'd9262, 16'd59941, 16'd9228, 16'd2365, 16'd39559});
	test_expansion(128'hce0c1a87aef9ade1fc6ea4363d643e37, {16'd42676, 16'd51149, 16'd5169, 16'd49320, 16'd9270, 16'd38041, 16'd4707, 16'd33495, 16'd29354, 16'd47672, 16'd9030, 16'd261, 16'd30402, 16'd10766, 16'd24680, 16'd34045, 16'd35894, 16'd37332, 16'd19087, 16'd27580, 16'd30173, 16'd56239, 16'd6389, 16'd15288, 16'd28748, 16'd39544});
	test_expansion(128'h797d916af61f1478a6bf958373f8c293, {16'd50581, 16'd52634, 16'd50194, 16'd56054, 16'd60303, 16'd41687, 16'd10895, 16'd16324, 16'd50948, 16'd34899, 16'd43766, 16'd60512, 16'd58835, 16'd4021, 16'd29222, 16'd15709, 16'd21927, 16'd10309, 16'd25208, 16'd63294, 16'd41854, 16'd27349, 16'd16238, 16'd20291, 16'd59345, 16'd42054});
	test_expansion(128'ha314630d4d8a36cf98c4cd0161e80dfe, {16'd57027, 16'd39731, 16'd23338, 16'd26802, 16'd14697, 16'd2235, 16'd34424, 16'd38295, 16'd16010, 16'd2336, 16'd17688, 16'd34356, 16'd34971, 16'd19190, 16'd42898, 16'd13781, 16'd23095, 16'd33933, 16'd6248, 16'd8432, 16'd5458, 16'd2710, 16'd49553, 16'd42260, 16'd43131, 16'd21164});
	test_expansion(128'h1bf5559f4614c16b0b525162fec7e76f, {16'd58823, 16'd3710, 16'd50136, 16'd18082, 16'd22741, 16'd24544, 16'd33720, 16'd65266, 16'd22115, 16'd36560, 16'd15481, 16'd10070, 16'd56011, 16'd25337, 16'd12975, 16'd51782, 16'd65127, 16'd3135, 16'd24101, 16'd18834, 16'd3067, 16'd4734, 16'd51018, 16'd36682, 16'd35037, 16'd19375});
	test_expansion(128'hb41c77586707c1c707bc1dffc29b43b2, {16'd31903, 16'd59134, 16'd53153, 16'd22340, 16'd25813, 16'd18760, 16'd14320, 16'd14139, 16'd6105, 16'd54465, 16'd40386, 16'd6494, 16'd33317, 16'd25541, 16'd57685, 16'd30676, 16'd45510, 16'd61995, 16'd14649, 16'd20447, 16'd1814, 16'd50078, 16'd12913, 16'd62414, 16'd51663, 16'd4179});
	test_expansion(128'h47fcc654e06c257441553f95f0ad1d41, {16'd54384, 16'd58404, 16'd52731, 16'd58826, 16'd26102, 16'd11904, 16'd34701, 16'd42836, 16'd37709, 16'd3997, 16'd887, 16'd62191, 16'd33514, 16'd24186, 16'd65137, 16'd2463, 16'd60527, 16'd23417, 16'd22152, 16'd55792, 16'd25824, 16'd14478, 16'd51769, 16'd38309, 16'd24776, 16'd43840});
	test_expansion(128'hb878056c464a56c9d6c2434f2a667485, {16'd43764, 16'd20877, 16'd32068, 16'd28784, 16'd35715, 16'd6390, 16'd18539, 16'd18931, 16'd6830, 16'd56005, 16'd36019, 16'd5744, 16'd10360, 16'd55445, 16'd44300, 16'd10747, 16'd45200, 16'd14589, 16'd27415, 16'd12895, 16'd10367, 16'd43107, 16'd39202, 16'd24561, 16'd41530, 16'd56427});
	test_expansion(128'h46a8b1e5e4c567f08ff8cfd27949a6c3, {16'd38541, 16'd43126, 16'd38834, 16'd50495, 16'd8108, 16'd28777, 16'd57847, 16'd40209, 16'd60177, 16'd12770, 16'd52955, 16'd49612, 16'd37090, 16'd3245, 16'd38421, 16'd14907, 16'd41934, 16'd9317, 16'd28550, 16'd64797, 16'd29134, 16'd32591, 16'd33981, 16'd61016, 16'd52146, 16'd34334});
	test_expansion(128'h95b903dd6dfb5680b21771ccb18e375f, {16'd28433, 16'd17557, 16'd28807, 16'd45915, 16'd49599, 16'd27782, 16'd10198, 16'd3475, 16'd8883, 16'd2818, 16'd23471, 16'd37593, 16'd44262, 16'd4486, 16'd8908, 16'd21307, 16'd51578, 16'd49735, 16'd34211, 16'd9687, 16'd53803, 16'd14701, 16'd28447, 16'd4315, 16'd56095, 16'd60080});
	test_expansion(128'h5fac317e9595064a017da45ecadba02c, {16'd5808, 16'd44243, 16'd8863, 16'd63609, 16'd8235, 16'd18042, 16'd47276, 16'd36331, 16'd6165, 16'd48905, 16'd26050, 16'd26475, 16'd37855, 16'd24614, 16'd41683, 16'd21324, 16'd45903, 16'd2849, 16'd17768, 16'd1378, 16'd2883, 16'd20615, 16'd56107, 16'd54544, 16'd59734, 16'd63638});
	test_expansion(128'h5059cf3ebe78b9c4b2a83c45fbb468cc, {16'd18955, 16'd15274, 16'd20828, 16'd60184, 16'd55451, 16'd64545, 16'd3483, 16'd63251, 16'd6335, 16'd27258, 16'd51736, 16'd44077, 16'd25872, 16'd54191, 16'd27664, 16'd57398, 16'd22162, 16'd47452, 16'd3629, 16'd44138, 16'd26511, 16'd44927, 16'd45587, 16'd29316, 16'd56380, 16'd52218});
	test_expansion(128'h4699a77666cb03ae1c448457e58a765c, {16'd6259, 16'd27565, 16'd46640, 16'd13948, 16'd60444, 16'd39132, 16'd32753, 16'd27123, 16'd47134, 16'd4094, 16'd15037, 16'd13756, 16'd46882, 16'd12712, 16'd1048, 16'd16951, 16'd12651, 16'd43325, 16'd43142, 16'd29537, 16'd4760, 16'd43525, 16'd41452, 16'd42074, 16'd62480, 16'd36188});
	test_expansion(128'h662992b41913638f74e50b9d719cc08d, {16'd1883, 16'd16176, 16'd62132, 16'd45193, 16'd21981, 16'd38626, 16'd54285, 16'd55244, 16'd4990, 16'd27876, 16'd2738, 16'd35697, 16'd13805, 16'd38243, 16'd30440, 16'd13962, 16'd5479, 16'd49554, 16'd5937, 16'd15696, 16'd52310, 16'd51355, 16'd15671, 16'd14525, 16'd58034, 16'd60573});
	test_expansion(128'h537a3a62fc83607f1532b47ca491bc60, {16'd45568, 16'd47546, 16'd754, 16'd56140, 16'd16627, 16'd48728, 16'd42557, 16'd61923, 16'd21569, 16'd54472, 16'd40937, 16'd53854, 16'd47990, 16'd11543, 16'd31057, 16'd36561, 16'd10293, 16'd50372, 16'd27259, 16'd59150, 16'd26706, 16'd57996, 16'd61118, 16'd13651, 16'd50709, 16'd55987});
	test_expansion(128'h6fd9f374ec408e424917da81b1eb9132, {16'd34899, 16'd8977, 16'd46477, 16'd41033, 16'd32973, 16'd56445, 16'd62239, 16'd43961, 16'd27302, 16'd39821, 16'd60989, 16'd34202, 16'd39378, 16'd43339, 16'd46910, 16'd56845, 16'd8778, 16'd22530, 16'd24121, 16'd58177, 16'd49458, 16'd47842, 16'd54555, 16'd55238, 16'd19610, 16'd44218});
	test_expansion(128'hbb8e947ff9050f573a4e7fcc55e7eca1, {16'd28034, 16'd35661, 16'd11606, 16'd36676, 16'd2080, 16'd303, 16'd30521, 16'd2349, 16'd14046, 16'd2299, 16'd34225, 16'd29814, 16'd25498, 16'd47450, 16'd39370, 16'd65226, 16'd64786, 16'd48364, 16'd37332, 16'd39892, 16'd50558, 16'd57375, 16'd48228, 16'd642, 16'd34079, 16'd17556});
	test_expansion(128'h708e8c28e671fb50d1f25f760e50d8f6, {16'd46423, 16'd21670, 16'd18356, 16'd43245, 16'd28965, 16'd8617, 16'd23913, 16'd6032, 16'd50316, 16'd51706, 16'd12402, 16'd30218, 16'd64476, 16'd63720, 16'd51471, 16'd43347, 16'd50563, 16'd21927, 16'd19020, 16'd64116, 16'd44365, 16'd56213, 16'd57764, 16'd28545, 16'd22066, 16'd65325});
	test_expansion(128'h3f4d022a6aa4033021185e353d3c428e, {16'd30589, 16'd8953, 16'd56037, 16'd2783, 16'd22152, 16'd1970, 16'd9002, 16'd8785, 16'd57586, 16'd13163, 16'd7334, 16'd3835, 16'd11064, 16'd56511, 16'd7549, 16'd37283, 16'd22806, 16'd10452, 16'd58577, 16'd37430, 16'd1003, 16'd24821, 16'd21550, 16'd16392, 16'd35280, 16'd19853});
	test_expansion(128'hcceef8f0f692568ea4caf82a37531702, {16'd22567, 16'd50954, 16'd24966, 16'd24579, 16'd43209, 16'd63465, 16'd54243, 16'd35043, 16'd2607, 16'd53830, 16'd32190, 16'd17884, 16'd54687, 16'd42978, 16'd9813, 16'd533, 16'd19480, 16'd51231, 16'd10515, 16'd7572, 16'd52202, 16'd62236, 16'd6194, 16'd28718, 16'd36426, 16'd35370});
	test_expansion(128'hf792b84efd2f097f9ff81954bc2f7398, {16'd36216, 16'd32337, 16'd22205, 16'd9965, 16'd34185, 16'd26599, 16'd43582, 16'd17793, 16'd61506, 16'd58186, 16'd41449, 16'd39862, 16'd28464, 16'd4807, 16'd57978, 16'd6428, 16'd506, 16'd60154, 16'd45675, 16'd64085, 16'd40137, 16'd13005, 16'd21361, 16'd13035, 16'd46183, 16'd46336});
	test_expansion(128'h96452f1bf5f42eb30c1acef63c59f12a, {16'd8531, 16'd1383, 16'd27077, 16'd34422, 16'd13535, 16'd50204, 16'd16530, 16'd8383, 16'd32193, 16'd64174, 16'd61428, 16'd22205, 16'd48077, 16'd52105, 16'd44986, 16'd4059, 16'd29992, 16'd61489, 16'd3171, 16'd30762, 16'd59994, 16'd14424, 16'd4981, 16'd24381, 16'd27610, 16'd12626});
	test_expansion(128'h372fb972385a1470ea37845ae75d32ae, {16'd26414, 16'd11495, 16'd26167, 16'd16956, 16'd7941, 16'd10022, 16'd572, 16'd47621, 16'd36544, 16'd52585, 16'd15384, 16'd60552, 16'd11933, 16'd47773, 16'd10675, 16'd24387, 16'd50665, 16'd54395, 16'd62457, 16'd11769, 16'd17455, 16'd52110, 16'd16147, 16'd63205, 16'd13220, 16'd2524});
	test_expansion(128'hc33748a82ad855ea69c2e6667f17f616, {16'd42308, 16'd36686, 16'd56499, 16'd6695, 16'd56529, 16'd39408, 16'd43014, 16'd8847, 16'd27463, 16'd41950, 16'd27025, 16'd29779, 16'd39449, 16'd22017, 16'd61097, 16'd29953, 16'd42211, 16'd51461, 16'd9296, 16'd59475, 16'd59812, 16'd6121, 16'd10072, 16'd42089, 16'd13409, 16'd61088});
	test_expansion(128'h90af1e53b3fb316aa991ec45855ed675, {16'd4704, 16'd4696, 16'd22955, 16'd18271, 16'd3560, 16'd59474, 16'd15992, 16'd52665, 16'd56998, 16'd49012, 16'd52796, 16'd55683, 16'd33200, 16'd49327, 16'd55162, 16'd40976, 16'd2593, 16'd21272, 16'd14794, 16'd9638, 16'd208, 16'd37543, 16'd26522, 16'd48187, 16'd36606, 16'd59174});
	test_expansion(128'hfffd27d61591a0121ad3691544c6ad35, {16'd56317, 16'd49953, 16'd64245, 16'd37322, 16'd43631, 16'd39943, 16'd12573, 16'd44747, 16'd4830, 16'd9671, 16'd1177, 16'd61695, 16'd45796, 16'd59429, 16'd56337, 16'd29887, 16'd3404, 16'd55204, 16'd47387, 16'd19366, 16'd19250, 16'd23643, 16'd26312, 16'd37978, 16'd53957, 16'd17229});
	test_expansion(128'h708ee63be24be89656c0edb9dc56e13a, {16'd4569, 16'd20679, 16'd44922, 16'd35261, 16'd43130, 16'd3606, 16'd26410, 16'd55410, 16'd59806, 16'd46552, 16'd48941, 16'd49822, 16'd33962, 16'd40654, 16'd4670, 16'd33753, 16'd42246, 16'd24070, 16'd429, 16'd8015, 16'd27809, 16'd62156, 16'd24848, 16'd22201, 16'd40953, 16'd24980});
	test_expansion(128'h19a9425a3796f10f8ee6e51610b05c3c, {16'd41442, 16'd42259, 16'd2692, 16'd48380, 16'd20584, 16'd55191, 16'd18520, 16'd24831, 16'd12504, 16'd25070, 16'd17569, 16'd2268, 16'd6083, 16'd51273, 16'd2805, 16'd38787, 16'd16760, 16'd27094, 16'd40130, 16'd8728, 16'd54140, 16'd30719, 16'd36741, 16'd56915, 16'd44912, 16'd38656});
	test_expansion(128'hb6ab5be3b6226d860c3cb18a776e8fb8, {16'd37992, 16'd44193, 16'd65227, 16'd40058, 16'd26110, 16'd32026, 16'd59198, 16'd27763, 16'd27732, 16'd61809, 16'd3371, 16'd540, 16'd38261, 16'd46880, 16'd64342, 16'd14412, 16'd31040, 16'd36295, 16'd22730, 16'd49758, 16'd6398, 16'd47011, 16'd28077, 16'd59633, 16'd58675, 16'd51874});
	test_expansion(128'h59fc4392aa0ff2d329557bfd42be8aa2, {16'd58110, 16'd1675, 16'd30586, 16'd23264, 16'd31911, 16'd28995, 16'd46203, 16'd45995, 16'd53332, 16'd7991, 16'd7904, 16'd61587, 16'd46736, 16'd24410, 16'd34222, 16'd51224, 16'd5974, 16'd61928, 16'd34785, 16'd16291, 16'd1532, 16'd17608, 16'd61247, 16'd22294, 16'd31764, 16'd3833});
	test_expansion(128'h8e8284c64942e47db24929a67751a062, {16'd16033, 16'd23669, 16'd35487, 16'd41122, 16'd43436, 16'd26398, 16'd40586, 16'd65261, 16'd48308, 16'd51059, 16'd40790, 16'd16255, 16'd14753, 16'd38841, 16'd8732, 16'd44010, 16'd29974, 16'd35860, 16'd57671, 16'd51691, 16'd22281, 16'd992, 16'd36283, 16'd61339, 16'd22576, 16'd61938});
	test_expansion(128'hae9bb6d6e3d2bcb265d0308c4870bf27, {16'd20556, 16'd31065, 16'd45853, 16'd47765, 16'd47721, 16'd10746, 16'd46651, 16'd35982, 16'd40110, 16'd26819, 16'd15471, 16'd16371, 16'd35234, 16'd3600, 16'd40187, 16'd34625, 16'd48014, 16'd29415, 16'd35665, 16'd63627, 16'd45489, 16'd48666, 16'd1020, 16'd60405, 16'd18565, 16'd27764});
	test_expansion(128'hbc95d29043a69f3d4d1825b1e9fe76a3, {16'd60512, 16'd52861, 16'd5030, 16'd30071, 16'd62737, 16'd22998, 16'd8603, 16'd29894, 16'd15569, 16'd27830, 16'd4486, 16'd32683, 16'd58272, 16'd28089, 16'd34689, 16'd59022, 16'd14988, 16'd32061, 16'd15886, 16'd13562, 16'd54337, 16'd50532, 16'd43318, 16'd65056, 16'd26393, 16'd19315});
	test_expansion(128'he40ee24b3b601b7a66caf37a2e953297, {16'd57876, 16'd2997, 16'd10656, 16'd47146, 16'd24908, 16'd20229, 16'd43771, 16'd16222, 16'd1425, 16'd24078, 16'd40308, 16'd42274, 16'd37968, 16'd13038, 16'd47677, 16'd44852, 16'd30356, 16'd43969, 16'd16706, 16'd49928, 16'd16363, 16'd34326, 16'd59226, 16'd18797, 16'd2513, 16'd35658});
	test_expansion(128'h655b6a9394a870470b9bb11e4e3a32b7, {16'd2811, 16'd18449, 16'd63110, 16'd60410, 16'd62754, 16'd60593, 16'd49411, 16'd9577, 16'd35094, 16'd22754, 16'd2911, 16'd31369, 16'd53204, 16'd52290, 16'd28473, 16'd11810, 16'd4735, 16'd59345, 16'd64838, 16'd41055, 16'd33681, 16'd37082, 16'd39198, 16'd57679, 16'd45927, 16'd22108});
	test_expansion(128'h8e5e2782764c20fc24770fa3d21160bf, {16'd29425, 16'd33346, 16'd8114, 16'd27438, 16'd26209, 16'd42234, 16'd15737, 16'd9140, 16'd27397, 16'd57581, 16'd3947, 16'd6450, 16'd7591, 16'd27620, 16'd18933, 16'd29259, 16'd2642, 16'd5064, 16'd63054, 16'd53099, 16'd31905, 16'd6933, 16'd49541, 16'd24076, 16'd47594, 16'd58610});
	test_expansion(128'h6b8e983e2148898c6fb259d838c2d99a, {16'd20411, 16'd45111, 16'd30760, 16'd3376, 16'd26821, 16'd38343, 16'd37815, 16'd62544, 16'd20307, 16'd14842, 16'd56824, 16'd32518, 16'd3121, 16'd49080, 16'd49514, 16'd8209, 16'd44902, 16'd35097, 16'd56820, 16'd60840, 16'd38566, 16'd17800, 16'd37176, 16'd5421, 16'd9728, 16'd17621});
	test_expansion(128'h808c90bbb6d0cd8a209b40a51dbe9382, {16'd59596, 16'd49843, 16'd33913, 16'd46750, 16'd30724, 16'd34835, 16'd11969, 16'd29884, 16'd43872, 16'd29553, 16'd30824, 16'd8151, 16'd63914, 16'd53609, 16'd5626, 16'd52163, 16'd310, 16'd50516, 16'd58596, 16'd5986, 16'd57140, 16'd6533, 16'd5217, 16'd41560, 16'd42114, 16'd43233});
	test_expansion(128'h84dd1c79d6ab713efde271079cafff16, {16'd17559, 16'd22526, 16'd9874, 16'd1289, 16'd30193, 16'd60834, 16'd17617, 16'd61272, 16'd26099, 16'd10790, 16'd26147, 16'd29919, 16'd35832, 16'd49461, 16'd2203, 16'd22815, 16'd6664, 16'd57579, 16'd31141, 16'd46608, 16'd41401, 16'd8390, 16'd62898, 16'd12558, 16'd22768, 16'd59855});
	test_expansion(128'h04eb04c5ed3adf2e494d40ce0c517952, {16'd35440, 16'd31695, 16'd43401, 16'd28776, 16'd56336, 16'd11805, 16'd58444, 16'd21313, 16'd58894, 16'd19623, 16'd25292, 16'd2395, 16'd15300, 16'd24217, 16'd39089, 16'd15073, 16'd63095, 16'd64435, 16'd36285, 16'd18083, 16'd64785, 16'd32646, 16'd40023, 16'd52554, 16'd9965, 16'd14575});
	test_expansion(128'hb4ab088ab9fad11cb49c6577173c75f1, {16'd31016, 16'd28684, 16'd17695, 16'd62580, 16'd52492, 16'd52406, 16'd61222, 16'd41438, 16'd38023, 16'd24496, 16'd29629, 16'd9420, 16'd27286, 16'd553, 16'd3735, 16'd65119, 16'd40800, 16'd6319, 16'd60486, 16'd51289, 16'd34616, 16'd55414, 16'd36235, 16'd27115, 16'd35200, 16'd43098});
	test_expansion(128'hb76bf50a5c8c1ff3ce60c4791bde7d53, {16'd36360, 16'd26948, 16'd4889, 16'd6672, 16'd17576, 16'd31431, 16'd24376, 16'd24067, 16'd21727, 16'd32384, 16'd38393, 16'd12884, 16'd61690, 16'd56233, 16'd5468, 16'd43571, 16'd21967, 16'd2924, 16'd61626, 16'd25404, 16'd62788, 16'd44816, 16'd26710, 16'd22495, 16'd44624, 16'd58920});
	test_expansion(128'h9e2787d63074ee24e8f4b2dc9723a20f, {16'd12412, 16'd26801, 16'd2675, 16'd15178, 16'd12031, 16'd43527, 16'd45811, 16'd24105, 16'd776, 16'd12633, 16'd37017, 16'd48025, 16'd33965, 16'd6076, 16'd43546, 16'd32322, 16'd4580, 16'd48441, 16'd878, 16'd7814, 16'd54844, 16'd15656, 16'd27940, 16'd5242, 16'd14899, 16'd16972});
	test_expansion(128'h01d6d0b560e681c0ded172924fc46a0a, {16'd6918, 16'd61983, 16'd5996, 16'd4756, 16'd35902, 16'd123, 16'd2530, 16'd5082, 16'd65047, 16'd45149, 16'd22274, 16'd34539, 16'd13235, 16'd60270, 16'd47619, 16'd58392, 16'd22882, 16'd31627, 16'd63262, 16'd8301, 16'd48509, 16'd51433, 16'd64288, 16'd10942, 16'd58585, 16'd4549});
	test_expansion(128'h5a7def10b21ba9230cc66890b08a28c0, {16'd36083, 16'd35440, 16'd51576, 16'd8815, 16'd31328, 16'd31084, 16'd50281, 16'd27273, 16'd23824, 16'd31694, 16'd45181, 16'd1995, 16'd45781, 16'd44699, 16'd2778, 16'd61636, 16'd26448, 16'd15365, 16'd3443, 16'd63268, 16'd60524, 16'd31339, 16'd732, 16'd27589, 16'd11468, 16'd34827});
	test_expansion(128'h91ab41deebe3be584e6fbd5ab8fe060a, {16'd47424, 16'd49587, 16'd13982, 16'd10341, 16'd63165, 16'd41633, 16'd12516, 16'd39328, 16'd41773, 16'd36050, 16'd48623, 16'd8398, 16'd54475, 16'd25187, 16'd38012, 16'd18679, 16'd38527, 16'd10550, 16'd14129, 16'd7166, 16'd21674, 16'd63732, 16'd33767, 16'd50132, 16'd52713, 16'd40987});
	test_expansion(128'h32453a84d82e8286e37e7647226acd20, {16'd36608, 16'd15511, 16'd31725, 16'd2830, 16'd32329, 16'd12833, 16'd33021, 16'd41687, 16'd58595, 16'd28176, 16'd14826, 16'd44626, 16'd21864, 16'd42698, 16'd53550, 16'd40734, 16'd53444, 16'd47619, 16'd33190, 16'd14127, 16'd37655, 16'd31230, 16'd65190, 16'd28076, 16'd9113, 16'd1088});
	test_expansion(128'he5c45821e4550966bd5cee839522f108, {16'd28308, 16'd6513, 16'd50418, 16'd34143, 16'd38277, 16'd65184, 16'd8002, 16'd49269, 16'd39381, 16'd53846, 16'd51840, 16'd16314, 16'd59898, 16'd13254, 16'd38527, 16'd46241, 16'd6984, 16'd5668, 16'd13727, 16'd36125, 16'd63623, 16'd25179, 16'd58611, 16'd60702, 16'd51916, 16'd14119});
	test_expansion(128'h6182fa0cfb2cdb6278d8f909fe870997, {16'd43886, 16'd49812, 16'd47961, 16'd5874, 16'd51267, 16'd14484, 16'd7212, 16'd12173, 16'd51218, 16'd39106, 16'd39393, 16'd390, 16'd8325, 16'd23263, 16'd24995, 16'd21084, 16'd51793, 16'd7667, 16'd41742, 16'd17577, 16'd23864, 16'd13233, 16'd57027, 16'd21636, 16'd27174, 16'd7586});
	test_expansion(128'he3d764d7bef47a46895243b7b31ef284, {16'd36572, 16'd44519, 16'd39032, 16'd35760, 16'd25615, 16'd1791, 16'd11530, 16'd56091, 16'd999, 16'd37328, 16'd53845, 16'd30123, 16'd62121, 16'd44606, 16'd7466, 16'd58019, 16'd7971, 16'd4303, 16'd60665, 16'd41642, 16'd57268, 16'd48991, 16'd44718, 16'd58063, 16'd20382, 16'd27622});
	test_expansion(128'h44a75e6083be8eb6abc07413e0a93d15, {16'd47334, 16'd4943, 16'd6725, 16'd11526, 16'd44409, 16'd56367, 16'd41114, 16'd56673, 16'd5066, 16'd11791, 16'd24950, 16'd46107, 16'd13557, 16'd62825, 16'd49492, 16'd60428, 16'd57210, 16'd56423, 16'd17437, 16'd59591, 16'd23532, 16'd60618, 16'd52195, 16'd27939, 16'd61109, 16'd8491});
	test_expansion(128'h35aa831c99d06eb652cc5fcb37569f31, {16'd18166, 16'd15572, 16'd15055, 16'd59106, 16'd58170, 16'd62609, 16'd59565, 16'd61736, 16'd41169, 16'd20856, 16'd12254, 16'd52713, 16'd47487, 16'd22030, 16'd64937, 16'd29208, 16'd204, 16'd11567, 16'd21686, 16'd38314, 16'd1424, 16'd51275, 16'd17172, 16'd29766, 16'd6469, 16'd7255});
	test_expansion(128'hdbe6c2dcbf61fd5a18726938b8825a12, {16'd12096, 16'd10563, 16'd2778, 16'd14530, 16'd8569, 16'd4880, 16'd31170, 16'd29212, 16'd39976, 16'd10512, 16'd14194, 16'd55703, 16'd9677, 16'd48626, 16'd29868, 16'd8817, 16'd22847, 16'd26751, 16'd53093, 16'd65360, 16'd39139, 16'd38680, 16'd42776, 16'd2163, 16'd10740, 16'd22826});
	test_expansion(128'h135b0adc90adb4a2433b08c9206f501d, {16'd52064, 16'd48049, 16'd10248, 16'd20507, 16'd63584, 16'd46012, 16'd31134, 16'd30300, 16'd48051, 16'd20438, 16'd15263, 16'd8839, 16'd59319, 16'd9854, 16'd11842, 16'd41587, 16'd24672, 16'd32241, 16'd64980, 16'd32287, 16'd32652, 16'd47658, 16'd3283, 16'd41358, 16'd10541, 16'd15529});
	test_expansion(128'h0c6601f8d34ccf115ed7f326b11c96cb, {16'd23768, 16'd7924, 16'd41549, 16'd418, 16'd42434, 16'd63464, 16'd34814, 16'd31833, 16'd12550, 16'd5051, 16'd49158, 16'd52889, 16'd27327, 16'd23094, 16'd27289, 16'd20977, 16'd35405, 16'd52664, 16'd59872, 16'd62884, 16'd39685, 16'd1522, 16'd2653, 16'd5580, 16'd36878, 16'd61503});
	test_expansion(128'hf0d535d1569e0c1e7ea461e13308ce3d, {16'd25183, 16'd14470, 16'd19942, 16'd61280, 16'd50198, 16'd61262, 16'd58916, 16'd35847, 16'd23088, 16'd53499, 16'd10011, 16'd50884, 16'd55165, 16'd58980, 16'd42687, 16'd4760, 16'd30082, 16'd21728, 16'd56136, 16'd4246, 16'd54589, 16'd43489, 16'd33799, 16'd52940, 16'd42016, 16'd30943});
	test_expansion(128'hdd4d0b4a2c9e35b63ffdfae4b80ccb68, {16'd15605, 16'd2073, 16'd20998, 16'd41373, 16'd57002, 16'd11269, 16'd6977, 16'd33973, 16'd63625, 16'd58507, 16'd23317, 16'd4648, 16'd41066, 16'd8118, 16'd25179, 16'd5116, 16'd2336, 16'd3544, 16'd55161, 16'd602, 16'd52206, 16'd44025, 16'd64748, 16'd65172, 16'd49791, 16'd3036});
	test_expansion(128'h45fb1af1ea7c27e9c84c021596109708, {16'd926, 16'd54145, 16'd22611, 16'd45106, 16'd40179, 16'd26716, 16'd2622, 16'd37410, 16'd1397, 16'd26288, 16'd5960, 16'd41582, 16'd17009, 16'd14349, 16'd4624, 16'd60528, 16'd46441, 16'd9825, 16'd44648, 16'd28013, 16'd26869, 16'd43118, 16'd50525, 16'd1758, 16'd23017, 16'd28742});
	test_expansion(128'ha23ec1482ed46b0e46bedf47708a1a71, {16'd9855, 16'd24628, 16'd15563, 16'd16694, 16'd47997, 16'd17507, 16'd20943, 16'd4695, 16'd10230, 16'd10236, 16'd59949, 16'd33631, 16'd8734, 16'd53055, 16'd60046, 16'd6274, 16'd59736, 16'd29733, 16'd23626, 16'd42864, 16'd27135, 16'd6915, 16'd2631, 16'd26181, 16'd5726, 16'd18536});
	test_expansion(128'hd4db2ef0087f45c97159c66a7deeb46b, {16'd34059, 16'd4424, 16'd8226, 16'd27717, 16'd36347, 16'd19134, 16'd45509, 16'd1006, 16'd36048, 16'd31830, 16'd33873, 16'd9275, 16'd54593, 16'd29817, 16'd47910, 16'd58233, 16'd3593, 16'd28012, 16'd24937, 16'd48816, 16'd9153, 16'd10738, 16'd19560, 16'd18391, 16'd61819, 16'd18672});
	test_expansion(128'h6e0074f8a7bfcc9375e9c3923ac6a7ab, {16'd50797, 16'd50399, 16'd51415, 16'd25387, 16'd19842, 16'd63011, 16'd9712, 16'd54117, 16'd12709, 16'd14702, 16'd7709, 16'd61540, 16'd59887, 16'd45453, 16'd60122, 16'd24297, 16'd55078, 16'd27812, 16'd41386, 16'd57259, 16'd4917, 16'd14497, 16'd6908, 16'd26972, 16'd45906, 16'd62454});
	test_expansion(128'h66499c9e50a383cae2597deb7caf6621, {16'd50155, 16'd53241, 16'd27667, 16'd28107, 16'd4957, 16'd34874, 16'd50075, 16'd12026, 16'd37575, 16'd28779, 16'd30130, 16'd3757, 16'd32496, 16'd55191, 16'd36518, 16'd43752, 16'd52927, 16'd3223, 16'd44990, 16'd28919, 16'd55805, 16'd55005, 16'd14710, 16'd20190, 16'd31877, 16'd9445});
	test_expansion(128'h3d9bbf16d53aa4e9ee6aaf1a7be2b00e, {16'd14560, 16'd56725, 16'd33178, 16'd5958, 16'd38449, 16'd38167, 16'd6124, 16'd55746, 16'd62291, 16'd56228, 16'd22744, 16'd60853, 16'd10007, 16'd36527, 16'd3832, 16'd36461, 16'd54116, 16'd37592, 16'd38399, 16'd8675, 16'd50958, 16'd57893, 16'd230, 16'd34964, 16'd26651, 16'd57666});
	test_expansion(128'h659ec6adc8cb72bb404b38a6ea8d29be, {16'd62219, 16'd8260, 16'd52904, 16'd14378, 16'd54551, 16'd61500, 16'd60797, 16'd28902, 16'd49548, 16'd5655, 16'd15532, 16'd63479, 16'd34386, 16'd38402, 16'd11962, 16'd56751, 16'd28505, 16'd56481, 16'd35886, 16'd25588, 16'd27389, 16'd4667, 16'd38563, 16'd62379, 16'd37985, 16'd32883});
	test_expansion(128'ha8f1b39a0c1815b08d957d334a6fb2cb, {16'd16070, 16'd20273, 16'd40508, 16'd29898, 16'd59135, 16'd649, 16'd7767, 16'd8266, 16'd45942, 16'd55277, 16'd27262, 16'd27067, 16'd58258, 16'd65052, 16'd18114, 16'd63209, 16'd31909, 16'd17669, 16'd45436, 16'd19879, 16'd23028, 16'd10007, 16'd47260, 16'd61030, 16'd1464, 16'd12920});
	test_expansion(128'h42dcbfe87f69c9f5b76d50d7c78bae58, {16'd10270, 16'd1756, 16'd63334, 16'd46345, 16'd39184, 16'd32987, 16'd47048, 16'd64905, 16'd13395, 16'd36744, 16'd24428, 16'd18236, 16'd36718, 16'd24522, 16'd55677, 16'd22085, 16'd49572, 16'd11235, 16'd36030, 16'd38498, 16'd63142, 16'd6002, 16'd27430, 16'd675, 16'd40293, 16'd23313});
	test_expansion(128'hd3c37073b16c8b3b88b4462567c2f1b5, {16'd7056, 16'd54072, 16'd58466, 16'd9160, 16'd11569, 16'd32093, 16'd42428, 16'd52341, 16'd14517, 16'd33132, 16'd63247, 16'd62468, 16'd49232, 16'd3418, 16'd64972, 16'd47957, 16'd12212, 16'd12192, 16'd39520, 16'd42508, 16'd53412, 16'd5571, 16'd14575, 16'd19235, 16'd29189, 16'd55098});
	test_expansion(128'h51b1a8fa5eeab48925fc1ed99be5f217, {16'd22272, 16'd11619, 16'd43659, 16'd51206, 16'd49570, 16'd54207, 16'd1011, 16'd43912, 16'd29131, 16'd39487, 16'd41039, 16'd25972, 16'd37083, 16'd6815, 16'd30784, 16'd43612, 16'd16640, 16'd21091, 16'd51685, 16'd28562, 16'd33370, 16'd42992, 16'd16720, 16'd33147, 16'd26698, 16'd22360});
	test_expansion(128'hc4800e50b9b519165cdd2ae0bbec5c6c, {16'd45160, 16'd43679, 16'd64464, 16'd24095, 16'd54997, 16'd59954, 16'd55966, 16'd27752, 16'd63522, 16'd10441, 16'd12020, 16'd34510, 16'd50765, 16'd29739, 16'd61559, 16'd12995, 16'd8003, 16'd18490, 16'd20050, 16'd47943, 16'd1193, 16'd27915, 16'd9010, 16'd41224, 16'd28691, 16'd42764});
	test_expansion(128'h9296521bc8757d2c391cca5b3beed6fd, {16'd35875, 16'd24926, 16'd54256, 16'd50174, 16'd59073, 16'd7564, 16'd4202, 16'd30819, 16'd33707, 16'd16093, 16'd41637, 16'd41593, 16'd12612, 16'd1320, 16'd13173, 16'd55431, 16'd34266, 16'd53262, 16'd7957, 16'd64737, 16'd42317, 16'd52482, 16'd41928, 16'd19049, 16'd30991, 16'd30634});
	test_expansion(128'hc02a3bc32aab1685e4666e111914de83, {16'd16392, 16'd2928, 16'd56924, 16'd57304, 16'd3354, 16'd41422, 16'd59745, 16'd20843, 16'd18885, 16'd41914, 16'd54654, 16'd50800, 16'd35250, 16'd44031, 16'd1786, 16'd63803, 16'd8148, 16'd9386, 16'd10695, 16'd18770, 16'd15823, 16'd29557, 16'd26542, 16'd28722, 16'd4254, 16'd22031});
	test_expansion(128'h4153bad8b6d965c27c6c89d51ea51160, {16'd8656, 16'd46186, 16'd16703, 16'd60474, 16'd41731, 16'd55923, 16'd24728, 16'd7737, 16'd5893, 16'd3623, 16'd7525, 16'd38929, 16'd55587, 16'd56076, 16'd37023, 16'd22712, 16'd30081, 16'd14314, 16'd15492, 16'd29023, 16'd48046, 16'd12722, 16'd34050, 16'd22748, 16'd29981, 16'd13869});
	test_expansion(128'hd1960ef07d384bb4754c52d69709a234, {16'd61854, 16'd28085, 16'd28441, 16'd24936, 16'd38373, 16'd42147, 16'd19521, 16'd28495, 16'd21802, 16'd20566, 16'd15335, 16'd41828, 16'd50425, 16'd15074, 16'd34541, 16'd5345, 16'd63974, 16'd63850, 16'd3014, 16'd55970, 16'd2437, 16'd29376, 16'd8218, 16'd2136, 16'd30349, 16'd27587});
	test_expansion(128'h12ccb82d19e98a4cab6f7610049513d5, {16'd49470, 16'd22603, 16'd49026, 16'd54300, 16'd28045, 16'd34146, 16'd2123, 16'd37033, 16'd37961, 16'd35163, 16'd48680, 16'd17939, 16'd24430, 16'd45721, 16'd7656, 16'd19250, 16'd58335, 16'd63088, 16'd44067, 16'd55716, 16'd32123, 16'd40804, 16'd33825, 16'd37621, 16'd27911, 16'd33717});
	test_expansion(128'h7ea78a425aac57573dbb2985cca520f0, {16'd42529, 16'd8998, 16'd50089, 16'd51011, 16'd27723, 16'd2327, 16'd28489, 16'd22233, 16'd38375, 16'd51282, 16'd36855, 16'd48928, 16'd45049, 16'd14536, 16'd64417, 16'd26553, 16'd46751, 16'd19794, 16'd53288, 16'd17383, 16'd57402, 16'd25521, 16'd35451, 16'd47106, 16'd14644, 16'd6203});
	test_expansion(128'hf7010bf1a0dab016b8d7cf3e2cb0f095, {16'd36543, 16'd30944, 16'd17740, 16'd44390, 16'd814, 16'd56911, 16'd42306, 16'd9085, 16'd8541, 16'd58440, 16'd58823, 16'd42944, 16'd34386, 16'd26727, 16'd6010, 16'd51487, 16'd20668, 16'd17328, 16'd8479, 16'd29945, 16'd58638, 16'd10652, 16'd38758, 16'd35108, 16'd13451, 16'd40078});
	test_expansion(128'h73cda52b278549c9459ef39a1f0ffd5b, {16'd52170, 16'd22205, 16'd35772, 16'd40505, 16'd5063, 16'd41179, 16'd54966, 16'd47735, 16'd26270, 16'd53254, 16'd44876, 16'd37271, 16'd32796, 16'd46065, 16'd20251, 16'd12699, 16'd45079, 16'd2927, 16'd16804, 16'd56273, 16'd15497, 16'd50743, 16'd4359, 16'd29365, 16'd53153, 16'd27390});
	test_expansion(128'h275b00e0c106fb99f42a0a1d83626499, {16'd48003, 16'd24480, 16'd51907, 16'd14490, 16'd44705, 16'd3070, 16'd11361, 16'd21933, 16'd19939, 16'd62897, 16'd46530, 16'd30817, 16'd17928, 16'd16419, 16'd27026, 16'd30653, 16'd55805, 16'd24088, 16'd32600, 16'd10540, 16'd3358, 16'd60068, 16'd61003, 16'd20566, 16'd34525, 16'd14586});
	test_expansion(128'h428e6e6f22b31c44dfac9bd61c2982de, {16'd23513, 16'd13683, 16'd29772, 16'd20943, 16'd28309, 16'd60085, 16'd21270, 16'd41289, 16'd14760, 16'd20714, 16'd31976, 16'd46884, 16'd24820, 16'd16167, 16'd15028, 16'd36888, 16'd20572, 16'd15439, 16'd63759, 16'd33060, 16'd53223, 16'd5366, 16'd40011, 16'd22930, 16'd24193, 16'd48002});
	test_expansion(128'h97ec14af3d02c90119a982f5407da14a, {16'd11672, 16'd57743, 16'd46954, 16'd58122, 16'd39495, 16'd64121, 16'd33492, 16'd34244, 16'd1408, 16'd42043, 16'd23728, 16'd59679, 16'd52678, 16'd16116, 16'd25530, 16'd51097, 16'd8134, 16'd61398, 16'd14012, 16'd57618, 16'd57897, 16'd37972, 16'd19884, 16'd30826, 16'd40330, 16'd17568});
	test_expansion(128'h1137a91abe6ead54b63402a7b57cb1cd, {16'd21547, 16'd41214, 16'd15320, 16'd58904, 16'd3989, 16'd37747, 16'd301, 16'd49180, 16'd55067, 16'd57168, 16'd630, 16'd22658, 16'd56002, 16'd53830, 16'd37877, 16'd7152, 16'd37458, 16'd24590, 16'd15721, 16'd41806, 16'd46354, 16'd28447, 16'd14557, 16'd30720, 16'd31877, 16'd11223});
	test_expansion(128'he2f8a273a9ee113171c33b68c8ac7761, {16'd65464, 16'd45609, 16'd29636, 16'd5610, 16'd64092, 16'd58007, 16'd5746, 16'd56357, 16'd14966, 16'd2537, 16'd50308, 16'd40696, 16'd2736, 16'd24128, 16'd60499, 16'd19578, 16'd14009, 16'd12003, 16'd56944, 16'd50576, 16'd65525, 16'd36066, 16'd30070, 16'd21131, 16'd58894, 16'd22030});
	test_expansion(128'hf609e167c469059fb78c390f7ba6424b, {16'd62084, 16'd40926, 16'd44094, 16'd8491, 16'd54922, 16'd4291, 16'd59796, 16'd38922, 16'd47972, 16'd51609, 16'd42243, 16'd61404, 16'd1599, 16'd37281, 16'd49166, 16'd55344, 16'd30617, 16'd31995, 16'd36567, 16'd3487, 16'd16529, 16'd59023, 16'd42464, 16'd2223, 16'd60772, 16'd2337});
	test_expansion(128'h01b71b8c8615cec54dfbefe947a364d7, {16'd21794, 16'd27916, 16'd40859, 16'd24964, 16'd23317, 16'd65015, 16'd38302, 16'd14863, 16'd14009, 16'd39775, 16'd51008, 16'd30130, 16'd2397, 16'd32930, 16'd41602, 16'd54177, 16'd4458, 16'd16174, 16'd47294, 16'd58981, 16'd26255, 16'd2635, 16'd58868, 16'd33005, 16'd50026, 16'd25727});
	test_expansion(128'h98ceb95efd7ac18d0b0a51639df07b49, {16'd58746, 16'd3064, 16'd63298, 16'd33142, 16'd19163, 16'd49286, 16'd40766, 16'd14899, 16'd54518, 16'd16101, 16'd33421, 16'd3335, 16'd19496, 16'd19450, 16'd29805, 16'd39907, 16'd23301, 16'd24212, 16'd63640, 16'd22461, 16'd24460, 16'd17163, 16'd45677, 16'd42902, 16'd51000, 16'd13689});
	test_expansion(128'h3587db22a2bcf78448e22f064f7219a6, {16'd7437, 16'd5586, 16'd1686, 16'd5410, 16'd43206, 16'd54950, 16'd5791, 16'd22349, 16'd5027, 16'd13155, 16'd32801, 16'd14113, 16'd16176, 16'd34706, 16'd55067, 16'd38802, 16'd3858, 16'd15462, 16'd25333, 16'd31125, 16'd55615, 16'd8899, 16'd33551, 16'd33975, 16'd19497, 16'd28114});
	test_expansion(128'h0ea1c325bc7fde42104679fa619b9c5e, {16'd35964, 16'd57001, 16'd28257, 16'd12192, 16'd1085, 16'd9744, 16'd19646, 16'd60884, 16'd3712, 16'd41650, 16'd39545, 16'd103, 16'd9267, 16'd57342, 16'd65276, 16'd58803, 16'd53157, 16'd28469, 16'd436, 16'd52138, 16'd44110, 16'd38348, 16'd59041, 16'd3371, 16'd42554, 16'd37810});
	test_expansion(128'ha1ab91e07cc7ba1872b95ebcc0678c49, {16'd25482, 16'd12733, 16'd5723, 16'd6922, 16'd48317, 16'd39716, 16'd4652, 16'd13561, 16'd3788, 16'd55536, 16'd15962, 16'd4467, 16'd2412, 16'd31008, 16'd33934, 16'd56673, 16'd1955, 16'd23042, 16'd52037, 16'd2564, 16'd53193, 16'd64451, 16'd60628, 16'd63743, 16'd43878, 16'd52447});
	test_expansion(128'h1fb76ce48de202f817459a506cf9f439, {16'd65515, 16'd38428, 16'd14829, 16'd59394, 16'd9388, 16'd3477, 16'd43673, 16'd62098, 16'd48840, 16'd58074, 16'd3512, 16'd46047, 16'd50151, 16'd61473, 16'd63458, 16'd44872, 16'd44930, 16'd36986, 16'd43703, 16'd13350, 16'd64747, 16'd1959, 16'd64485, 16'd62034, 16'd41202, 16'd39088});
	test_expansion(128'hacad4429c7a53ae48f72742697e3e874, {16'd55418, 16'd51292, 16'd61518, 16'd56802, 16'd11234, 16'd339, 16'd12452, 16'd36254, 16'd44918, 16'd38573, 16'd27826, 16'd5642, 16'd42236, 16'd2799, 16'd47054, 16'd64268, 16'd48022, 16'd1608, 16'd31882, 16'd58520, 16'd13356, 16'd44691, 16'd34900, 16'd16238, 16'd31570, 16'd22277});
	test_expansion(128'hf4b9390f7c9e201e987f66b6dcf1e3c9, {16'd3975, 16'd37467, 16'd2507, 16'd51724, 16'd11449, 16'd45093, 16'd13780, 16'd3016, 16'd48441, 16'd13646, 16'd20601, 16'd15521, 16'd51464, 16'd12844, 16'd40024, 16'd42108, 16'd48716, 16'd6745, 16'd49734, 16'd23506, 16'd52264, 16'd62180, 16'd33790, 16'd20860, 16'd2208, 16'd42543});
	test_expansion(128'hb411ece6dd901d066ffe815857b9572f, {16'd23257, 16'd28930, 16'd43768, 16'd7803, 16'd5486, 16'd63742, 16'd50002, 16'd42683, 16'd43802, 16'd43133, 16'd42447, 16'd49101, 16'd62597, 16'd12255, 16'd13853, 16'd3051, 16'd56985, 16'd24303, 16'd54090, 16'd48097, 16'd57432, 16'd62465, 16'd26344, 16'd51754, 16'd14945, 16'd34721});
	test_expansion(128'h7c0c4a237992e6331270df52f0e8e6bf, {16'd15341, 16'd12591, 16'd30223, 16'd28719, 16'd27405, 16'd22136, 16'd44352, 16'd39954, 16'd10519, 16'd27926, 16'd46392, 16'd50886, 16'd43141, 16'd31321, 16'd30957, 16'd21707, 16'd43338, 16'd51930, 16'd38797, 16'd63332, 16'd60019, 16'd41552, 16'd38278, 16'd46492, 16'd63436, 16'd9236});
	test_expansion(128'he301953ad2249929d2df14b9f5f8deb6, {16'd49185, 16'd27752, 16'd27451, 16'd65450, 16'd45380, 16'd811, 16'd17555, 16'd34746, 16'd45251, 16'd48502, 16'd14946, 16'd32373, 16'd17905, 16'd45992, 16'd18229, 16'd7128, 16'd6351, 16'd3382, 16'd25765, 16'd22902, 16'd3299, 16'd38845, 16'd53328, 16'd14911, 16'd57388, 16'd26337});
	test_expansion(128'hed72daeaa5cdc2b0037cdfa765f81b2b, {16'd60548, 16'd1337, 16'd24750, 16'd60139, 16'd50319, 16'd53115, 16'd60907, 16'd13614, 16'd28974, 16'd43708, 16'd10463, 16'd57860, 16'd9752, 16'd55079, 16'd55633, 16'd11294, 16'd39005, 16'd15614, 16'd19741, 16'd12827, 16'd25928, 16'd15432, 16'd1169, 16'd9934, 16'd40834, 16'd9537});
	test_expansion(128'h6d975d2b25ce265cd44f4ade4c9d3500, {16'd8470, 16'd15852, 16'd27746, 16'd38306, 16'd57622, 16'd21661, 16'd42900, 16'd11834, 16'd36915, 16'd61859, 16'd11035, 16'd23106, 16'd35034, 16'd13540, 16'd63282, 16'd59316, 16'd33947, 16'd47745, 16'd21310, 16'd32469, 16'd15168, 16'd36295, 16'd25383, 16'd6299, 16'd36335, 16'd61547});
	test_expansion(128'hbcf9d7a746d162072eedac584548f43b, {16'd7037, 16'd52071, 16'd49203, 16'd46462, 16'd21877, 16'd1210, 16'd6918, 16'd60263, 16'd16913, 16'd55836, 16'd27676, 16'd24949, 16'd23702, 16'd59604, 16'd24901, 16'd39439, 16'd34102, 16'd62234, 16'd42731, 16'd47652, 16'd9697, 16'd29771, 16'd16643, 16'd43502, 16'd22357, 16'd48261});
	test_expansion(128'hbe8c7248953af11b7bfe32feb0219f25, {16'd477, 16'd57305, 16'd17725, 16'd41552, 16'd55476, 16'd41864, 16'd62802, 16'd18707, 16'd47456, 16'd30934, 16'd12367, 16'd39909, 16'd149, 16'd63811, 16'd44937, 16'd8896, 16'd7492, 16'd61940, 16'd47313, 16'd44787, 16'd36800, 16'd30733, 16'd32935, 16'd48105, 16'd31712, 16'd25206});
	test_expansion(128'hb345529ebc5ffa7626edee97d03a27ee, {16'd5105, 16'd40981, 16'd53317, 16'd60093, 16'd6210, 16'd630, 16'd58756, 16'd23284, 16'd45478, 16'd54919, 16'd50124, 16'd41370, 16'd27529, 16'd36180, 16'd17119, 16'd27726, 16'd40342, 16'd54758, 16'd58914, 16'd7918, 16'd14445, 16'd21637, 16'd30582, 16'd31397, 16'd48962, 16'd63572});
	test_expansion(128'h9153e174878dc3f203bae2a80a1e6c87, {16'd33784, 16'd40574, 16'd37175, 16'd23810, 16'd29544, 16'd1847, 16'd34095, 16'd28251, 16'd4514, 16'd16400, 16'd12551, 16'd44246, 16'd31802, 16'd29941, 16'd29160, 16'd56285, 16'd55146, 16'd56402, 16'd64149, 16'd28396, 16'd48791, 16'd20664, 16'd8921, 16'd7082, 16'd58664, 16'd20340});
	test_expansion(128'h04b95d5836590afb078fcc34c30d6c55, {16'd61123, 16'd11999, 16'd54494, 16'd22119, 16'd16422, 16'd35152, 16'd48174, 16'd13920, 16'd48172, 16'd65081, 16'd55955, 16'd50442, 16'd3752, 16'd63265, 16'd9651, 16'd1304, 16'd32708, 16'd4765, 16'd6744, 16'd12195, 16'd53140, 16'd26772, 16'd60110, 16'd17464, 16'd62046, 16'd63508});
	test_expansion(128'h101bdca29166989d35dec6fe672c610d, {16'd23742, 16'd40812, 16'd10953, 16'd65486, 16'd56816, 16'd1487, 16'd54181, 16'd45637, 16'd4942, 16'd27663, 16'd65264, 16'd65296, 16'd59056, 16'd59867, 16'd31746, 16'd30362, 16'd9957, 16'd14697, 16'd19870, 16'd52650, 16'd21657, 16'd13021, 16'd5073, 16'd16189, 16'd16230, 16'd32473});
	test_expansion(128'hf6f3dfe26b5271007fb799fd2215cf0a, {16'd56181, 16'd15899, 16'd30702, 16'd25018, 16'd9403, 16'd63358, 16'd19052, 16'd40473, 16'd50080, 16'd54449, 16'd51679, 16'd21615, 16'd28694, 16'd7733, 16'd64258, 16'd56787, 16'd4649, 16'd26772, 16'd19584, 16'd62529, 16'd59508, 16'd6905, 16'd21343, 16'd58481, 16'd47233, 16'd24008});
	test_expansion(128'h3693b0555a9eadef09ddc81f7370a848, {16'd64315, 16'd38579, 16'd31911, 16'd61818, 16'd33697, 16'd2787, 16'd7937, 16'd28800, 16'd19919, 16'd6056, 16'd31881, 16'd23958, 16'd11231, 16'd6506, 16'd44039, 16'd44843, 16'd29438, 16'd16122, 16'd11169, 16'd3616, 16'd37852, 16'd7145, 16'd36263, 16'd61949, 16'd54349, 16'd54746});
	test_expansion(128'h84f2ab2115e0dadf4178251e27dece42, {16'd43752, 16'd44365, 16'd50084, 16'd38683, 16'd17836, 16'd44576, 16'd29064, 16'd26151, 16'd63328, 16'd40025, 16'd33834, 16'd50888, 16'd57852, 16'd51643, 16'd23172, 16'd4692, 16'd12776, 16'd26235, 16'd15487, 16'd58441, 16'd19904, 16'd3267, 16'd26902, 16'd14768, 16'd59853, 16'd59393});
	test_expansion(128'h037a07a2ab003fe0ce9361673727673a, {16'd59542, 16'd54196, 16'd48665, 16'd58501, 16'd25571, 16'd31686, 16'd50922, 16'd49501, 16'd44533, 16'd56796, 16'd7582, 16'd25679, 16'd8362, 16'd15425, 16'd6465, 16'd8548, 16'd20821, 16'd54798, 16'd49432, 16'd23422, 16'd44364, 16'd7066, 16'd28149, 16'd62319, 16'd56450, 16'd18026});
	test_expansion(128'h1850ceab2241d4d07dda1eeefa0a6973, {16'd16917, 16'd7154, 16'd39217, 16'd6003, 16'd30858, 16'd48102, 16'd46539, 16'd1261, 16'd26412, 16'd7160, 16'd43808, 16'd15451, 16'd28575, 16'd15903, 16'd18708, 16'd60368, 16'd15289, 16'd52900, 16'd64050, 16'd55275, 16'd27805, 16'd59466, 16'd62712, 16'd51501, 16'd35719, 16'd40502});
	test_expansion(128'h1f9764c71d8cab0e5afc2c1f9b392be8, {16'd55500, 16'd64646, 16'd26596, 16'd12262, 16'd41594, 16'd624, 16'd41596, 16'd37835, 16'd26952, 16'd22016, 16'd22501, 16'd19153, 16'd62663, 16'd63140, 16'd25905, 16'd36554, 16'd17224, 16'd12070, 16'd52409, 16'd7480, 16'd16631, 16'd9199, 16'd49498, 16'd9760, 16'd38395, 16'd54017});
	test_expansion(128'h4e6a7219198994a1cbee2fd7397ea2f4, {16'd26391, 16'd63210, 16'd56344, 16'd44352, 16'd4349, 16'd31201, 16'd29378, 16'd47259, 16'd7876, 16'd57661, 16'd31162, 16'd25109, 16'd40972, 16'd56203, 16'd25784, 16'd42491, 16'd24205, 16'd54139, 16'd47363, 16'd64688, 16'd54633, 16'd37149, 16'd18897, 16'd42522, 16'd37522, 16'd18754});
	test_expansion(128'hb504a3c4002fd75398584e92d58e5579, {16'd44049, 16'd23232, 16'd35273, 16'd26508, 16'd21170, 16'd32561, 16'd38087, 16'd52130, 16'd32235, 16'd47131, 16'd34875, 16'd47732, 16'd56454, 16'd62171, 16'd61080, 16'd28755, 16'd5734, 16'd28897, 16'd32424, 16'd50838, 16'd3078, 16'd12308, 16'd57680, 16'd20624, 16'd10244, 16'd55912});
	test_expansion(128'h9feb0ac517138b35a57518643412192c, {16'd10576, 16'd50713, 16'd43874, 16'd65127, 16'd46089, 16'd50204, 16'd5780, 16'd39344, 16'd26103, 16'd58394, 16'd51955, 16'd58147, 16'd53012, 16'd39901, 16'd40107, 16'd36737, 16'd41694, 16'd39932, 16'd21698, 16'd32904, 16'd53253, 16'd41356, 16'd1609, 16'd11211, 16'd1401, 16'd49382});
	test_expansion(128'h93349026b936f1d3412e571cb744a405, {16'd19522, 16'd42291, 16'd28915, 16'd34016, 16'd53129, 16'd36254, 16'd62374, 16'd5385, 16'd37427, 16'd55474, 16'd19296, 16'd41840, 16'd44997, 16'd11552, 16'd50746, 16'd50355, 16'd42463, 16'd21653, 16'd39646, 16'd38026, 16'd36546, 16'd49314, 16'd17156, 16'd50886, 16'd5360, 16'd14466});
	test_expansion(128'ha9e8f9d7b3e21cc924b6d242b120123a, {16'd26051, 16'd9268, 16'd53380, 16'd60081, 16'd46804, 16'd40128, 16'd13242, 16'd34518, 16'd12277, 16'd28532, 16'd12016, 16'd15034, 16'd22432, 16'd33054, 16'd17605, 16'd17280, 16'd54323, 16'd24355, 16'd10633, 16'd36549, 16'd52046, 16'd55706, 16'd44860, 16'd24527, 16'd60607, 16'd459});
	test_expansion(128'ha1238c1ac1c95b1eb03dbe68fa0da6f9, {16'd7042, 16'd65377, 16'd28375, 16'd58102, 16'd32351, 16'd29384, 16'd12737, 16'd52443, 16'd5234, 16'd36562, 16'd51725, 16'd23774, 16'd42249, 16'd46473, 16'd56126, 16'd56998, 16'd53176, 16'd30721, 16'd39603, 16'd5294, 16'd12481, 16'd63558, 16'd21084, 16'd54626, 16'd58968, 16'd20328});
	test_expansion(128'h616dd61b94b2154de1eb21898bacdb02, {16'd48374, 16'd37381, 16'd59286, 16'd64327, 16'd23653, 16'd28322, 16'd29236, 16'd21783, 16'd4985, 16'd11376, 16'd44989, 16'd44869, 16'd18026, 16'd51532, 16'd60857, 16'd64913, 16'd18596, 16'd40754, 16'd33864, 16'd62973, 16'd3578, 16'd12514, 16'd37181, 16'd19592, 16'd52707, 16'd21185});
	test_expansion(128'he44ec44a9e89636c8a77d4f6d3269d5e, {16'd57867, 16'd38486, 16'd2528, 16'd56480, 16'd36109, 16'd31493, 16'd52494, 16'd19156, 16'd43482, 16'd31317, 16'd40419, 16'd21416, 16'd39240, 16'd29055, 16'd19936, 16'd10120, 16'd1549, 16'd28971, 16'd31164, 16'd16323, 16'd39920, 16'd2230, 16'd21353, 16'd29371, 16'd51055, 16'd4622});
	test_expansion(128'hb18b826ec8383157498e66b7f3c30180, {16'd30103, 16'd15311, 16'd14051, 16'd4654, 16'd5154, 16'd19071, 16'd43402, 16'd12095, 16'd11168, 16'd11941, 16'd17187, 16'd40727, 16'd25955, 16'd26429, 16'd61582, 16'd38572, 16'd10480, 16'd60766, 16'd3071, 16'd59933, 16'd6152, 16'd1843, 16'd17181, 16'd40589, 16'd168, 16'd20707});
	test_expansion(128'haffa554b309fe74f361df8ae56ae7299, {16'd26712, 16'd57469, 16'd53257, 16'd49128, 16'd58086, 16'd14304, 16'd2249, 16'd10006, 16'd47870, 16'd2713, 16'd49199, 16'd51453, 16'd6526, 16'd31647, 16'd24100, 16'd6232, 16'd21072, 16'd34006, 16'd6386, 16'd52746, 16'd48262, 16'd62997, 16'd13834, 16'd13725, 16'd19237, 16'd2738});
	test_expansion(128'hfc0dab465d818a623fe837e9d0ac7021, {16'd50722, 16'd41791, 16'd25812, 16'd8130, 16'd38662, 16'd37898, 16'd16774, 16'd33869, 16'd64359, 16'd39407, 16'd19768, 16'd7822, 16'd4910, 16'd4001, 16'd38533, 16'd2621, 16'd24132, 16'd12634, 16'd36043, 16'd50295, 16'd10126, 16'd3503, 16'd14037, 16'd14054, 16'd64848, 16'd9559});
	test_expansion(128'h43acf5501108c716b2d55721806525d0, {16'd56547, 16'd28807, 16'd15954, 16'd25921, 16'd43029, 16'd58672, 16'd39785, 16'd55141, 16'd10576, 16'd7477, 16'd55204, 16'd48212, 16'd3076, 16'd56029, 16'd55625, 16'd28631, 16'd3326, 16'd51617, 16'd30180, 16'd40746, 16'd16452, 16'd60137, 16'd49146, 16'd37283, 16'd50401, 16'd57727});
	test_expansion(128'hbc9b5671a3de28db90f0248cb0b6e873, {16'd58857, 16'd42422, 16'd3601, 16'd27194, 16'd3406, 16'd35348, 16'd13435, 16'd1728, 16'd45939, 16'd43693, 16'd61791, 16'd30907, 16'd5045, 16'd6084, 16'd37322, 16'd55657, 16'd35610, 16'd60426, 16'd38145, 16'd13408, 16'd64363, 16'd5919, 16'd7138, 16'd34393, 16'd59725, 16'd43383});
	test_expansion(128'h79a4ae47405d2caa5ee2d33ec8361211, {16'd55404, 16'd59140, 16'd9036, 16'd53603, 16'd47949, 16'd28566, 16'd21649, 16'd48377, 16'd47488, 16'd24030, 16'd64947, 16'd16840, 16'd24079, 16'd16204, 16'd2438, 16'd60548, 16'd7835, 16'd27451, 16'd1013, 16'd4496, 16'd13837, 16'd31168, 16'd33879, 16'd50600, 16'd28755, 16'd12364});
	test_expansion(128'h12f22f4b892695c291df9b94d7783af1, {16'd54823, 16'd44941, 16'd48456, 16'd18208, 16'd58737, 16'd28702, 16'd59932, 16'd25789, 16'd29576, 16'd3327, 16'd30645, 16'd43696, 16'd37548, 16'd53158, 16'd34020, 16'd54216, 16'd16240, 16'd6710, 16'd43137, 16'd22816, 16'd9764, 16'd43049, 16'd65381, 16'd55114, 16'd12430, 16'd47552});
	test_expansion(128'h7ce362223a439d440abe0cc6e5c11207, {16'd798, 16'd63699, 16'd48770, 16'd46728, 16'd25747, 16'd36897, 16'd45610, 16'd19524, 16'd18725, 16'd18294, 16'd24276, 16'd46295, 16'd16030, 16'd42789, 16'd29565, 16'd1605, 16'd20733, 16'd15058, 16'd37332, 16'd64577, 16'd7391, 16'd57563, 16'd14804, 16'd524, 16'd27656, 16'd10387});
	test_expansion(128'h7e9d10499019037a1047d6c1e8ca60b3, {16'd57129, 16'd9538, 16'd42090, 16'd29388, 16'd61051, 16'd27291, 16'd64292, 16'd14450, 16'd13222, 16'd50092, 16'd33321, 16'd22666, 16'd9611, 16'd47970, 16'd13843, 16'd59993, 16'd54914, 16'd31467, 16'd43350, 16'd38746, 16'd4251, 16'd31150, 16'd14885, 16'd7349, 16'd43778, 16'd6106});
	test_expansion(128'h99e8a397ff66e0feb87366d356bacbd0, {16'd32564, 16'd33287, 16'd46838, 16'd59514, 16'd33135, 16'd16558, 16'd31329, 16'd32461, 16'd29694, 16'd3157, 16'd17515, 16'd27110, 16'd27088, 16'd28446, 16'd40768, 16'd23391, 16'd27822, 16'd54180, 16'd26138, 16'd55769, 16'd24982, 16'd30024, 16'd35519, 16'd53166, 16'd45512, 16'd42102});
	test_expansion(128'h93641c2de2bd315ae2ad3ae649ce4dcc, {16'd25177, 16'd49440, 16'd52720, 16'd48020, 16'd7104, 16'd11591, 16'd9570, 16'd34238, 16'd23867, 16'd12639, 16'd18004, 16'd37679, 16'd13041, 16'd52143, 16'd15173, 16'd56919, 16'd20270, 16'd3114, 16'd3776, 16'd57491, 16'd54766, 16'd5128, 16'd4509, 16'd42137, 16'd42401, 16'd10835});
	test_expansion(128'h851aee624b3bd2a6cf5fa865185e9a30, {16'd36325, 16'd16833, 16'd4521, 16'd12842, 16'd44662, 16'd58731, 16'd30854, 16'd39832, 16'd34106, 16'd25748, 16'd42547, 16'd5727, 16'd15200, 16'd1989, 16'd35710, 16'd51481, 16'd45265, 16'd2229, 16'd43084, 16'd22086, 16'd9988, 16'd55547, 16'd40328, 16'd52799, 16'd37524, 16'd62322});
	test_expansion(128'haced59fc701b7837bb0f706a90276024, {16'd52051, 16'd32740, 16'd63812, 16'd21112, 16'd771, 16'd63773, 16'd48102, 16'd49190, 16'd32303, 16'd52406, 16'd62061, 16'd42888, 16'd50644, 16'd18669, 16'd40400, 16'd42809, 16'd10885, 16'd45265, 16'd8532, 16'd44138, 16'd27551, 16'd19135, 16'd22535, 16'd4581, 16'd9472, 16'd37277});
	test_expansion(128'h77d6d0096d24f77db8fb50b0a286b73b, {16'd54586, 16'd52325, 16'd2797, 16'd52486, 16'd18708, 16'd31036, 16'd54160, 16'd33845, 16'd21017, 16'd46239, 16'd53543, 16'd56187, 16'd36824, 16'd32868, 16'd29876, 16'd15067, 16'd53527, 16'd58502, 16'd21066, 16'd8801, 16'd29474, 16'd3219, 16'd35845, 16'd6548, 16'd12626, 16'd18358});
	test_expansion(128'hdf8413b099cf986b5f38dc0edfa5bd03, {16'd8192, 16'd52882, 16'd60030, 16'd15632, 16'd15906, 16'd8244, 16'd62674, 16'd9678, 16'd25272, 16'd46551, 16'd50971, 16'd13550, 16'd25551, 16'd54909, 16'd27560, 16'd20014, 16'd17209, 16'd60047, 16'd18105, 16'd59851, 16'd13883, 16'd7804, 16'd45987, 16'd55637, 16'd44127, 16'd34602});
	test_expansion(128'h9872536bacd2691374f422b0d5f3b9ef, {16'd11809, 16'd23443, 16'd50810, 16'd65332, 16'd34723, 16'd63716, 16'd19858, 16'd1049, 16'd36421, 16'd49694, 16'd41115, 16'd29271, 16'd17121, 16'd46180, 16'd60200, 16'd60640, 16'd33950, 16'd7228, 16'd11995, 16'd69, 16'd49398, 16'd9140, 16'd37889, 16'd10892, 16'd29706, 16'd64273});
	test_expansion(128'h4bab14b3b2312f16ddd12545d12b0213, {16'd6686, 16'd10022, 16'd20930, 16'd26231, 16'd43830, 16'd2613, 16'd58313, 16'd46280, 16'd4599, 16'd5156, 16'd34134, 16'd27366, 16'd17800, 16'd12328, 16'd33729, 16'd48870, 16'd33989, 16'd53733, 16'd39753, 16'd35770, 16'd3333, 16'd13256, 16'd2980, 16'd34623, 16'd55181, 16'd33832});
	test_expansion(128'hcfe76733614f8017a1eec36c1c089a9e, {16'd61417, 16'd5300, 16'd63690, 16'd5971, 16'd47136, 16'd58950, 16'd4425, 16'd48547, 16'd63575, 16'd57836, 16'd22502, 16'd17401, 16'd50478, 16'd28407, 16'd9943, 16'd19849, 16'd27646, 16'd46181, 16'd33877, 16'd8994, 16'd31707, 16'd47576, 16'd21889, 16'd42043, 16'd44817, 16'd28758});
	test_expansion(128'h122b71ae6323b99ce005664bc4bd7e0c, {16'd37298, 16'd44560, 16'd6502, 16'd12574, 16'd19951, 16'd8211, 16'd61121, 16'd2158, 16'd7849, 16'd44281, 16'd31491, 16'd13149, 16'd28722, 16'd27404, 16'd46160, 16'd17562, 16'd28546, 16'd43604, 16'd39550, 16'd43449, 16'd64512, 16'd31236, 16'd39694, 16'd59296, 16'd6826, 16'd30402});
	test_expansion(128'ha1c130937aed68748c68a57dfe6505c9, {16'd43336, 16'd59493, 16'd6480, 16'd22185, 16'd15686, 16'd46768, 16'd25804, 16'd58420, 16'd36399, 16'd37229, 16'd34970, 16'd49703, 16'd30077, 16'd54130, 16'd29579, 16'd10880, 16'd40803, 16'd522, 16'd3053, 16'd59871, 16'd40339, 16'd10316, 16'd37205, 16'd17082, 16'd41010, 16'd30791});
	test_expansion(128'h20e2ab2f784af1ac11b40202eb9e3ec0, {16'd63630, 16'd31627, 16'd13709, 16'd36003, 16'd32976, 16'd54150, 16'd50973, 16'd22110, 16'd42043, 16'd8415, 16'd1691, 16'd10727, 16'd500, 16'd19940, 16'd1008, 16'd4198, 16'd65187, 16'd25937, 16'd64904, 16'd39046, 16'd47499, 16'd5568, 16'd51337, 16'd46490, 16'd60575, 16'd43850});
	test_expansion(128'h3ca2ea605a489aeef190701afa21412a, {16'd880, 16'd61403, 16'd6464, 16'd15919, 16'd62752, 16'd63646, 16'd43437, 16'd59975, 16'd36360, 16'd10896, 16'd48421, 16'd33893, 16'd57347, 16'd45692, 16'd36360, 16'd16162, 16'd30715, 16'd2971, 16'd50819, 16'd42839, 16'd27176, 16'd10531, 16'd28919, 16'd24740, 16'd26215, 16'd38348});
	test_expansion(128'h639dbb5c404ef3eaf3d5f07e15debc6c, {16'd6506, 16'd54805, 16'd62975, 16'd22702, 16'd27891, 16'd61319, 16'd34294, 16'd25582, 16'd43104, 16'd6490, 16'd36786, 16'd4040, 16'd36623, 16'd3399, 16'd50204, 16'd38564, 16'd56422, 16'd40600, 16'd14127, 16'd64754, 16'd31707, 16'd51187, 16'd7247, 16'd45692, 16'd7990, 16'd9059});
	test_expansion(128'hf3539866fd13496dfa01057341adf06d, {16'd52013, 16'd58666, 16'd50507, 16'd41715, 16'd537, 16'd39850, 16'd25305, 16'd60763, 16'd63738, 16'd50256, 16'd21174, 16'd55034, 16'd51185, 16'd1704, 16'd62997, 16'd13785, 16'd58979, 16'd41441, 16'd35032, 16'd55048, 16'd51852, 16'd23491, 16'd20500, 16'd28611, 16'd64805, 16'd31775});
	test_expansion(128'h89941037fc552e446e055576748c7b95, {16'd5482, 16'd30024, 16'd27144, 16'd45717, 16'd49584, 16'd48370, 16'd51769, 16'd21547, 16'd15959, 16'd30688, 16'd64686, 16'd10266, 16'd17057, 16'd35287, 16'd55046, 16'd52336, 16'd21456, 16'd5713, 16'd35889, 16'd15417, 16'd61953, 16'd42097, 16'd44695, 16'd47050, 16'd47344, 16'd55073});
	test_expansion(128'hcc9f5b16e8b0739df57cf1e0f05e8ef4, {16'd45391, 16'd254, 16'd64054, 16'd20877, 16'd17772, 16'd51600, 16'd26722, 16'd5210, 16'd15382, 16'd64402, 16'd37433, 16'd55326, 16'd1864, 16'd14321, 16'd17560, 16'd48093, 16'd31359, 16'd57138, 16'd23250, 16'd39981, 16'd50860, 16'd59700, 16'd62116, 16'd13602, 16'd38157, 16'd9754});
	test_expansion(128'hc7e07e1d49e8292a51590d9c99c8dc84, {16'd31917, 16'd33815, 16'd38127, 16'd64754, 16'd54531, 16'd19624, 16'd31104, 16'd46770, 16'd20501, 16'd62314, 16'd40957, 16'd28805, 16'd8254, 16'd47722, 16'd39982, 16'd53831, 16'd27078, 16'd6675, 16'd34081, 16'd57464, 16'd28440, 16'd31993, 16'd40244, 16'd50164, 16'd13501, 16'd8864});
	test_expansion(128'h802aea8452409673dfba6722f9fbb636, {16'd18518, 16'd8617, 16'd15870, 16'd42503, 16'd23543, 16'd63751, 16'd24787, 16'd36971, 16'd16008, 16'd29402, 16'd56238, 16'd29579, 16'd11364, 16'd43454, 16'd11148, 16'd60031, 16'd11923, 16'd15927, 16'd8791, 16'd44077, 16'd23411, 16'd3656, 16'd44383, 16'd10546, 16'd33300, 16'd18224});
	test_expansion(128'h66d4ff29ad779b69f70e7586ab2dd41c, {16'd16592, 16'd9655, 16'd28335, 16'd42267, 16'd27776, 16'd8069, 16'd63028, 16'd58436, 16'd34395, 16'd34759, 16'd49025, 16'd27396, 16'd24129, 16'd48757, 16'd53856, 16'd2998, 16'd36332, 16'd21150, 16'd46203, 16'd49339, 16'd59558, 16'd46945, 16'd51130, 16'd58252, 16'd61786, 16'd64520});
	test_expansion(128'he241f4e2dbdb765eb22e1728f66f1232, {16'd35616, 16'd38809, 16'd31612, 16'd17428, 16'd23135, 16'd31671, 16'd9508, 16'd53236, 16'd35557, 16'd51393, 16'd25712, 16'd58615, 16'd34078, 16'd16783, 16'd41841, 16'd32439, 16'd56990, 16'd14705, 16'd61544, 16'd27608, 16'd60940, 16'd50325, 16'd13936, 16'd34982, 16'd20015, 16'd45568});
	test_expansion(128'ha8aee3b084c13522a24f96ebc76c9bf7, {16'd39041, 16'd15624, 16'd57645, 16'd21232, 16'd24772, 16'd14406, 16'd20469, 16'd63085, 16'd28931, 16'd54122, 16'd44983, 16'd31216, 16'd10133, 16'd37644, 16'd59082, 16'd20073, 16'd8990, 16'd36937, 16'd50682, 16'd48864, 16'd35115, 16'd41700, 16'd49326, 16'd45334, 16'd58261, 16'd6649});
	test_expansion(128'h160b0615f628f38243353f92fc4f21cd, {16'd22630, 16'd33037, 16'd33170, 16'd46647, 16'd62064, 16'd5955, 16'd35343, 16'd25824, 16'd21758, 16'd35731, 16'd23837, 16'd59814, 16'd16771, 16'd31658, 16'd38472, 16'd15246, 16'd39405, 16'd64588, 16'd33614, 16'd16624, 16'd23232, 16'd22870, 16'd15517, 16'd46079, 16'd27129, 16'd28116});
	test_expansion(128'h170a9b7203e197c3c90767effd3b885a, {16'd1425, 16'd47517, 16'd39361, 16'd34628, 16'd30274, 16'd62081, 16'd5597, 16'd28962, 16'd45278, 16'd63060, 16'd8560, 16'd45274, 16'd61094, 16'd30453, 16'd63513, 16'd63371, 16'd65356, 16'd27144, 16'd47646, 16'd14404, 16'd33235, 16'd1963, 16'd60258, 16'd26085, 16'd3079, 16'd17395});
	test_expansion(128'h73da65dddc2c6069914c4edf08058f7f, {16'd36037, 16'd61292, 16'd63181, 16'd38529, 16'd17747, 16'd35807, 16'd15239, 16'd15863, 16'd56514, 16'd28397, 16'd18539, 16'd37982, 16'd61507, 16'd43940, 16'd44173, 16'd39521, 16'd12742, 16'd2129, 16'd57738, 16'd62912, 16'd18838, 16'd36570, 16'd52428, 16'd52186, 16'd52142, 16'd22714});
	test_expansion(128'hf4fc99b5bd793e184e0f8599a73a499b, {16'd52372, 16'd11025, 16'd18498, 16'd45916, 16'd10146, 16'd3024, 16'd23578, 16'd34447, 16'd52644, 16'd2593, 16'd17357, 16'd55633, 16'd40353, 16'd36012, 16'd34663, 16'd16068, 16'd60995, 16'd5228, 16'd63478, 16'd26237, 16'd63415, 16'd37997, 16'd21619, 16'd61593, 16'd53221, 16'd26392});
	test_expansion(128'h617a27d16132d905155c887f4cb099e8, {16'd11849, 16'd29209, 16'd60684, 16'd29331, 16'd53871, 16'd8021, 16'd19103, 16'd9063, 16'd62885, 16'd12404, 16'd64257, 16'd27578, 16'd38903, 16'd25342, 16'd44748, 16'd13715, 16'd34056, 16'd14903, 16'd52248, 16'd37725, 16'd30097, 16'd29195, 16'd59181, 16'd13065, 16'd11759, 16'd52796});
	test_expansion(128'hef8221b5809314cd0504e7a3deb23112, {16'd33334, 16'd62928, 16'd11273, 16'd48959, 16'd9793, 16'd58752, 16'd16814, 16'd51652, 16'd47798, 16'd57409, 16'd20846, 16'd9914, 16'd45072, 16'd34568, 16'd40225, 16'd57112, 16'd33832, 16'd45261, 16'd1026, 16'd65036, 16'd1717, 16'd14613, 16'd34551, 16'd45708, 16'd65507, 16'd25927});
	test_expansion(128'hafc9b9e9aed71b46b2df8fbeeb123e3b, {16'd51901, 16'd49658, 16'd43614, 16'd4390, 16'd4826, 16'd30369, 16'd49184, 16'd28852, 16'd24042, 16'd56851, 16'd40873, 16'd57407, 16'd43015, 16'd42587, 16'd48559, 16'd59608, 16'd49228, 16'd1558, 16'd54378, 16'd30646, 16'd40501, 16'd19846, 16'd60504, 16'd62322, 16'd32096, 16'd16867});
	test_expansion(128'hb68c1424b719878bf8ed177581827f78, {16'd12442, 16'd29040, 16'd24544, 16'd27253, 16'd5927, 16'd5741, 16'd33875, 16'd18923, 16'd44133, 16'd39678, 16'd56485, 16'd42829, 16'd44316, 16'd6617, 16'd25810, 16'd22820, 16'd7110, 16'd28878, 16'd40179, 16'd6671, 16'd21917, 16'd51214, 16'd46007, 16'd34618, 16'd52860, 16'd21968});
	test_expansion(128'h95d62db21353032e4a5ab1e1e7e1f64a, {16'd41347, 16'd28439, 16'd61738, 16'd3744, 16'd47648, 16'd9399, 16'd30269, 16'd63295, 16'd47878, 16'd39617, 16'd24977, 16'd50361, 16'd50201, 16'd20770, 16'd4777, 16'd15082, 16'd3274, 16'd55862, 16'd32996, 16'd7135, 16'd2416, 16'd45571, 16'd30745, 16'd40771, 16'd60799, 16'd1323});
	test_expansion(128'h24d5b9245227dcbaf700be317954fc76, {16'd17547, 16'd35312, 16'd29158, 16'd54949, 16'd28678, 16'd240, 16'd62324, 16'd45777, 16'd37530, 16'd37805, 16'd12466, 16'd53420, 16'd40915, 16'd20029, 16'd55728, 16'd54666, 16'd29154, 16'd577, 16'd39147, 16'd24606, 16'd18926, 16'd53885, 16'd36271, 16'd9383, 16'd51324, 16'd20257});
	test_expansion(128'h4a26d9108d3d05ec9789783cd2dbff1c, {16'd22911, 16'd43600, 16'd36986, 16'd860, 16'd34560, 16'd11385, 16'd47391, 16'd22775, 16'd41031, 16'd50755, 16'd26163, 16'd28473, 16'd25173, 16'd19871, 16'd65448, 16'd21427, 16'd35928, 16'd27035, 16'd44182, 16'd61183, 16'd58402, 16'd63352, 16'd34700, 16'd42629, 16'd1482, 16'd19356});
	test_expansion(128'hc6476a9267c88aac2c437adaa58ea05a, {16'd767, 16'd61063, 16'd49491, 16'd44824, 16'd45636, 16'd1203, 16'd13632, 16'd14156, 16'd31346, 16'd19234, 16'd20111, 16'd39038, 16'd13763, 16'd37120, 16'd20032, 16'd44844, 16'd42157, 16'd17129, 16'd47560, 16'd52773, 16'd24297, 16'd24594, 16'd19255, 16'd24556, 16'd15313, 16'd58978});
	test_expansion(128'h57f9ba59fd6f54e9c84e4503b0846d5f, {16'd45889, 16'd23630, 16'd31515, 16'd46458, 16'd10317, 16'd36813, 16'd61926, 16'd29479, 16'd7851, 16'd53470, 16'd31456, 16'd65261, 16'd57163, 16'd29467, 16'd19262, 16'd51084, 16'd43867, 16'd29269, 16'd21717, 16'd31869, 16'd44687, 16'd46263, 16'd54259, 16'd4180, 16'd31863, 16'd5525});
	test_expansion(128'haf4c0bec4e7da68e96ab2359f6bc0236, {16'd55963, 16'd54827, 16'd1836, 16'd23878, 16'd49742, 16'd51655, 16'd45261, 16'd41282, 16'd22262, 16'd33607, 16'd15758, 16'd60490, 16'd9995, 16'd60839, 16'd46681, 16'd43596, 16'd12957, 16'd45297, 16'd25495, 16'd2861, 16'd14197, 16'd52396, 16'd54702, 16'd43907, 16'd59635, 16'd18334});
	test_expansion(128'h88a3f6fa944e9f1bd54a7590a07cad60, {16'd46575, 16'd36194, 16'd2129, 16'd2627, 16'd11695, 16'd42854, 16'd39740, 16'd34456, 16'd37715, 16'd32338, 16'd4503, 16'd20353, 16'd62523, 16'd30515, 16'd24178, 16'd48688, 16'd2078, 16'd40106, 16'd19783, 16'd8411, 16'd20501, 16'd23233, 16'd61878, 16'd45079, 16'd26893, 16'd57116});
	test_expansion(128'h483a38da96a95c05ee0fb0b386162438, {16'd2760, 16'd21898, 16'd14599, 16'd4934, 16'd45104, 16'd7222, 16'd3877, 16'd61824, 16'd49167, 16'd29395, 16'd53191, 16'd8437, 16'd14018, 16'd22864, 16'd39358, 16'd14934, 16'd51124, 16'd9969, 16'd35836, 16'd14904, 16'd30959, 16'd13043, 16'd33256, 16'd43309, 16'd42864, 16'd44678});
	test_expansion(128'h1ec4a7922472a7c4caa0244312b83e13, {16'd24547, 16'd20331, 16'd34745, 16'd26231, 16'd23789, 16'd14167, 16'd55117, 16'd20933, 16'd65221, 16'd12283, 16'd15061, 16'd62661, 16'd15824, 16'd23856, 16'd64260, 16'd31883, 16'd46495, 16'd43350, 16'd42242, 16'd34427, 16'd62892, 16'd3317, 16'd4893, 16'd61056, 16'd64709, 16'd42861});
	test_expansion(128'hcb9b9679a6035e5b5288579a44ad2e65, {16'd62569, 16'd266, 16'd36425, 16'd27101, 16'd142, 16'd59566, 16'd45165, 16'd61966, 16'd34586, 16'd45305, 16'd19864, 16'd17044, 16'd17839, 16'd16460, 16'd4999, 16'd16246, 16'd10587, 16'd48866, 16'd42253, 16'd39472, 16'd42273, 16'd51791, 16'd53230, 16'd52957, 16'd29036, 16'd61034});
	test_expansion(128'ha992ab95babcfc85b2283e9748d00aee, {16'd18284, 16'd9046, 16'd44757, 16'd26530, 16'd17219, 16'd2463, 16'd65180, 16'd12338, 16'd25779, 16'd19836, 16'd2138, 16'd21708, 16'd27165, 16'd64436, 16'd15370, 16'd47334, 16'd62397, 16'd12149, 16'd6214, 16'd27188, 16'd41404, 16'd3911, 16'd39351, 16'd28672, 16'd40491, 16'd36516});
	test_expansion(128'h6077307159d40ea5544039ba8c75b2f0, {16'd32305, 16'd57290, 16'd24904, 16'd7947, 16'd60825, 16'd56790, 16'd49978, 16'd7691, 16'd45494, 16'd45146, 16'd53849, 16'd40998, 16'd50154, 16'd38190, 16'd1647, 16'd13455, 16'd53667, 16'd22905, 16'd50945, 16'd60772, 16'd43146, 16'd14394, 16'd23172, 16'd36401, 16'd11345, 16'd58053});
	test_expansion(128'h5b7a6a7def7b4f905e70f21c1757f48b, {16'd49285, 16'd26348, 16'd21065, 16'd36790, 16'd47424, 16'd26342, 16'd51750, 16'd51504, 16'd62783, 16'd29221, 16'd51480, 16'd33116, 16'd53870, 16'd34797, 16'd50469, 16'd53661, 16'd62155, 16'd62488, 16'd8779, 16'd60440, 16'd29714, 16'd48731, 16'd10753, 16'd38807, 16'd27911, 16'd56057});
	test_expansion(128'h9b0ae0c43c85fadd82d2e2c79e05879f, {16'd42631, 16'd46480, 16'd62566, 16'd17921, 16'd63474, 16'd62339, 16'd19461, 16'd10885, 16'd26871, 16'd34549, 16'd65275, 16'd61427, 16'd49213, 16'd36632, 16'd11070, 16'd22490, 16'd20457, 16'd16235, 16'd61218, 16'd65383, 16'd21427, 16'd41872, 16'd36912, 16'd22825, 16'd61868, 16'd1787});
	test_expansion(128'h6b75242884ac529ed155b16dd57dd01c, {16'd45968, 16'd20693, 16'd56952, 16'd30638, 16'd19926, 16'd31523, 16'd52385, 16'd37345, 16'd51939, 16'd5449, 16'd50810, 16'd61646, 16'd17752, 16'd57702, 16'd65338, 16'd41603, 16'd11663, 16'd65532, 16'd59426, 16'd15926, 16'd44936, 16'd28072, 16'd35989, 16'd60925, 16'd47568, 16'd34396});
	test_expansion(128'he3ec818a977462fc5bc22d1eeff451df, {16'd9757, 16'd31774, 16'd47991, 16'd6398, 16'd55465, 16'd53414, 16'd39668, 16'd26193, 16'd11598, 16'd49463, 16'd25772, 16'd26699, 16'd63623, 16'd9504, 16'd25020, 16'd30196, 16'd41905, 16'd1030, 16'd14517, 16'd20094, 16'd6079, 16'd57833, 16'd57693, 16'd45293, 16'd50267, 16'd4050});
	test_expansion(128'hc3cecb2a71999b951f2bd028b1af4d3a, {16'd33717, 16'd59334, 16'd5944, 16'd22211, 16'd35746, 16'd505, 16'd29335, 16'd8904, 16'd60618, 16'd21472, 16'd22848, 16'd65253, 16'd23197, 16'd50545, 16'd9091, 16'd47135, 16'd65127, 16'd62927, 16'd13886, 16'd64948, 16'd61426, 16'd53693, 16'd27626, 16'd29705, 16'd64493, 16'd23560});
	test_expansion(128'h71fc867ca85320ad997dd5a7d77a4acb, {16'd5764, 16'd50189, 16'd1034, 16'd47859, 16'd22169, 16'd60432, 16'd31173, 16'd21585, 16'd13064, 16'd32694, 16'd33686, 16'd43875, 16'd39096, 16'd5643, 16'd9241, 16'd51714, 16'd19845, 16'd51399, 16'd12678, 16'd22508, 16'd10342, 16'd49769, 16'd37499, 16'd27208, 16'd36702, 16'd1549});
	test_expansion(128'hfab9da5f3a5492627e15a599fea10b67, {16'd46596, 16'd27938, 16'd59083, 16'd13187, 16'd33407, 16'd3898, 16'd4419, 16'd217, 16'd60407, 16'd43820, 16'd688, 16'd1350, 16'd25812, 16'd49557, 16'd15437, 16'd20225, 16'd31688, 16'd55593, 16'd41805, 16'd64774, 16'd52585, 16'd43599, 16'd25477, 16'd38866, 16'd25386, 16'd40217});
	test_expansion(128'h39e0e761b6bd877301b4166010ace896, {16'd41241, 16'd13606, 16'd37933, 16'd40179, 16'd20901, 16'd7610, 16'd28099, 16'd49314, 16'd22178, 16'd4754, 16'd60396, 16'd63652, 16'd35968, 16'd36642, 16'd48314, 16'd43201, 16'd12944, 16'd29978, 16'd25378, 16'd46431, 16'd21475, 16'd17610, 16'd32947, 16'd51630, 16'd21514, 16'd7305});
	test_expansion(128'h32ec1042c6ebc0a57425945a109e8590, {16'd13644, 16'd8878, 16'd63763, 16'd40883, 16'd27505, 16'd51628, 16'd59380, 16'd29976, 16'd23791, 16'd53356, 16'd46730, 16'd6818, 16'd40702, 16'd2938, 16'd9113, 16'd64842, 16'd36266, 16'd47978, 16'd27164, 16'd4741, 16'd47374, 16'd47746, 16'd60513, 16'd48134, 16'd65001, 16'd50401});
	test_expansion(128'h0222aadd899db30f33d559da3c8f3401, {16'd43379, 16'd32253, 16'd5638, 16'd19259, 16'd31958, 16'd36013, 16'd11860, 16'd43048, 16'd8827, 16'd44440, 16'd53562, 16'd43485, 16'd43664, 16'd47766, 16'd44493, 16'd15947, 16'd42443, 16'd44502, 16'd44125, 16'd63655, 16'd57531, 16'd15628, 16'd4450, 16'd60079, 16'd61247, 16'd40441});
	test_expansion(128'h1afed1fa189f0a2429ff703340c92528, {16'd17149, 16'd62137, 16'd7714, 16'd53083, 16'd23485, 16'd52378, 16'd25365, 16'd20111, 16'd8672, 16'd65223, 16'd45648, 16'd14089, 16'd37537, 16'd31045, 16'd18684, 16'd60276, 16'd28944, 16'd50393, 16'd41531, 16'd15357, 16'd14127, 16'd40317, 16'd931, 16'd48703, 16'd3701, 16'd26003});
	test_expansion(128'hef2d63946fa4830a7e48b10fec03bb52, {16'd57845, 16'd30831, 16'd6491, 16'd23145, 16'd51649, 16'd47680, 16'd3787, 16'd39107, 16'd36692, 16'd52714, 16'd14884, 16'd3476, 16'd11927, 16'd2026, 16'd13647, 16'd58090, 16'd25695, 16'd60401, 16'd13103, 16'd20453, 16'd37443, 16'd31145, 16'd56090, 16'd55283, 16'd48350, 16'd24531});
	test_expansion(128'hf2324fc4252a5a76a14ff69c3101c5c6, {16'd36568, 16'd40327, 16'd387, 16'd21142, 16'd10723, 16'd59252, 16'd49360, 16'd43989, 16'd31793, 16'd39551, 16'd56246, 16'd18882, 16'd54639, 16'd15589, 16'd30873, 16'd8752, 16'd56842, 16'd920, 16'd32365, 16'd13647, 16'd2756, 16'd60104, 16'd63026, 16'd26182, 16'd57182, 16'd13143});
	test_expansion(128'ha274f8604a775fb124a5f4c1319af638, {16'd32790, 16'd64890, 16'd52926, 16'd9298, 16'd39492, 16'd14860, 16'd50670, 16'd20137, 16'd13561, 16'd24287, 16'd28225, 16'd29179, 16'd24077, 16'd55558, 16'd7654, 16'd22428, 16'd14592, 16'd30194, 16'd6414, 16'd57980, 16'd51967, 16'd35540, 16'd57761, 16'd21295, 16'd1827, 16'd8582});
	test_expansion(128'h58c5b3ab5252f7e47539bcd3cd23fe59, {16'd58006, 16'd38497, 16'd15847, 16'd40475, 16'd29210, 16'd681, 16'd65153, 16'd33588, 16'd61391, 16'd8094, 16'd45774, 16'd63319, 16'd12576, 16'd2549, 16'd58465, 16'd6789, 16'd53251, 16'd26982, 16'd54447, 16'd35187, 16'd46997, 16'd49963, 16'd39366, 16'd8050, 16'd38782, 16'd24859});
	test_expansion(128'h97d86f6fcc00750c2bb570c4b65121a1, {16'd38154, 16'd35568, 16'd47514, 16'd42674, 16'd56498, 16'd4917, 16'd10339, 16'd59561, 16'd31103, 16'd52699, 16'd48431, 16'd6011, 16'd6792, 16'd33668, 16'd3226, 16'd29852, 16'd17853, 16'd21628, 16'd43477, 16'd63227, 16'd64702, 16'd9083, 16'd26906, 16'd30064, 16'd57327, 16'd34185});
	test_expansion(128'h63a176bb8c6176b9cebdc9802629052a, {16'd3099, 16'd44024, 16'd44027, 16'd53377, 16'd37784, 16'd25094, 16'd54950, 16'd35850, 16'd27703, 16'd18558, 16'd57920, 16'd44362, 16'd42435, 16'd26264, 16'd33446, 16'd44021, 16'd37577, 16'd24661, 16'd60761, 16'd14848, 16'd17026, 16'd37806, 16'd58844, 16'd50021, 16'd14599, 16'd47516});
	test_expansion(128'h57ba03ab9e7083d413360060135bd008, {16'd22113, 16'd11620, 16'd43896, 16'd34144, 16'd50974, 16'd5587, 16'd52786, 16'd54706, 16'd19156, 16'd44419, 16'd20269, 16'd30747, 16'd26107, 16'd37497, 16'd2688, 16'd13711, 16'd18330, 16'd35295, 16'd36133, 16'd24513, 16'd49178, 16'd10629, 16'd50749, 16'd43271, 16'd27035, 16'd63282});
	test_expansion(128'hc6ab45ae697122bb779739476c49ab51, {16'd60320, 16'd9077, 16'd17698, 16'd30978, 16'd18834, 16'd5101, 16'd46333, 16'd52602, 16'd34162, 16'd64548, 16'd42425, 16'd32692, 16'd8412, 16'd1784, 16'd2978, 16'd44016, 16'd37620, 16'd4324, 16'd32891, 16'd2563, 16'd50730, 16'd32120, 16'd45530, 16'd4671, 16'd18789, 16'd31679});
	test_expansion(128'h9d6169cab750109f86b2efaf4deaae66, {16'd21296, 16'd23597, 16'd33896, 16'd5761, 16'd13732, 16'd1578, 16'd64502, 16'd12781, 16'd63501, 16'd32274, 16'd53560, 16'd2446, 16'd64778, 16'd56161, 16'd62329, 16'd30426, 16'd27788, 16'd30548, 16'd46303, 16'd33147, 16'd44427, 16'd4445, 16'd16769, 16'd28286, 16'd42489, 16'd36932});
	test_expansion(128'hf6431fafe90b20b550fb7ba07eef7d69, {16'd59764, 16'd1326, 16'd39573, 16'd24811, 16'd7641, 16'd30494, 16'd37195, 16'd6714, 16'd2267, 16'd47329, 16'd22273, 16'd41327, 16'd38664, 16'd45885, 16'd2172, 16'd9631, 16'd21013, 16'd58351, 16'd48140, 16'd64940, 16'd35113, 16'd34171, 16'd21412, 16'd52667, 16'd36293, 16'd17062});
	test_expansion(128'hdcc2cba580244d414c981ca99d4bd2cd, {16'd52198, 16'd63291, 16'd64762, 16'd65198, 16'd53916, 16'd24917, 16'd27626, 16'd16321, 16'd37024, 16'd65180, 16'd23727, 16'd21602, 16'd8948, 16'd61379, 16'd52446, 16'd64196, 16'd19040, 16'd63440, 16'd4167, 16'd2162, 16'd15087, 16'd48968, 16'd10494, 16'd30021, 16'd2446, 16'd63671});
	test_expansion(128'hb805647e2c5d9c4b009d8b50632d6f31, {16'd34045, 16'd65309, 16'd44669, 16'd47114, 16'd24697, 16'd22868, 16'd31360, 16'd22469, 16'd20708, 16'd31187, 16'd33892, 16'd5915, 16'd51777, 16'd6867, 16'd8487, 16'd45617, 16'd12461, 16'd11954, 16'd4245, 16'd10694, 16'd14131, 16'd19903, 16'd10164, 16'd65238, 16'd39368, 16'd63480});
	test_expansion(128'hb99424155e240f60be03cdf1865ce559, {16'd20703, 16'd52030, 16'd42208, 16'd22182, 16'd32534, 16'd38450, 16'd36405, 16'd17273, 16'd8318, 16'd6677, 16'd13441, 16'd33433, 16'd50, 16'd36921, 16'd3462, 16'd7118, 16'd53656, 16'd12665, 16'd3625, 16'd25928, 16'd39598, 16'd24445, 16'd56093, 16'd17898, 16'd8636, 16'd59038});
	test_expansion(128'h059e063aebaace1ba4ee1a772afe3b5c, {16'd31505, 16'd30226, 16'd32943, 16'd3466, 16'd59464, 16'd56836, 16'd53473, 16'd32218, 16'd56055, 16'd16018, 16'd63633, 16'd9222, 16'd18145, 16'd39762, 16'd37634, 16'd20778, 16'd63408, 16'd61886, 16'd42354, 16'd5773, 16'd48688, 16'd2604, 16'd51306, 16'd59216, 16'd49801, 16'd64174});
	test_expansion(128'hf027b9f71ecd6fd0107fdc0fe3788bb3, {16'd5444, 16'd24430, 16'd32369, 16'd27095, 16'd9410, 16'd16425, 16'd10036, 16'd4224, 16'd36237, 16'd21067, 16'd19788, 16'd20883, 16'd32618, 16'd56287, 16'd22394, 16'd30823, 16'd54486, 16'd33351, 16'd65194, 16'd24692, 16'd7609, 16'd54694, 16'd15771, 16'd20659, 16'd782, 16'd9285});
	test_expansion(128'ha238d88114089b7399b79e203d67fd16, {16'd61417, 16'd26834, 16'd36757, 16'd40800, 16'd51441, 16'd20005, 16'd46329, 16'd16162, 16'd43236, 16'd58589, 16'd38731, 16'd32755, 16'd17251, 16'd62688, 16'd9027, 16'd22573, 16'd20636, 16'd62276, 16'd24948, 16'd46197, 16'd8735, 16'd35252, 16'd22794, 16'd32664, 16'd46844, 16'd2367});
	test_expansion(128'h23c1333fd8725fcde116d8d3da9c8a3a, {16'd30237, 16'd3166, 16'd28544, 16'd3094, 16'd11610, 16'd12601, 16'd44347, 16'd42431, 16'd9940, 16'd58107, 16'd55505, 16'd9117, 16'd38246, 16'd43012, 16'd38851, 16'd11059, 16'd64021, 16'd44660, 16'd33649, 16'd25594, 16'd43184, 16'd39867, 16'd5785, 16'd23701, 16'd42997, 16'd62535});
	test_expansion(128'hccbb686e21867c8e34b177d01650b0d5, {16'd36471, 16'd60446, 16'd22384, 16'd32063, 16'd36883, 16'd19607, 16'd60083, 16'd55253, 16'd58476, 16'd15062, 16'd28425, 16'd37542, 16'd16465, 16'd3251, 16'd9279, 16'd15136, 16'd25706, 16'd54352, 16'd1407, 16'd19559, 16'd14478, 16'd13550, 16'd25376, 16'd31701, 16'd26150, 16'd56776});
	test_expansion(128'hc5629a080573f3582e49f84134b0e899, {16'd42408, 16'd44745, 16'd28844, 16'd52240, 16'd26398, 16'd10429, 16'd55546, 16'd8491, 16'd17193, 16'd64398, 16'd31606, 16'd64633, 16'd33192, 16'd27405, 16'd35075, 16'd17238, 16'd47197, 16'd20905, 16'd44663, 16'd36574, 16'd34208, 16'd18398, 16'd6332, 16'd33671, 16'd24209, 16'd41253});
	test_expansion(128'h65bd552f357baa9b1b6e2d7feb5b663a, {16'd42789, 16'd5363, 16'd5199, 16'd31925, 16'd61499, 16'd39726, 16'd37809, 16'd50029, 16'd33424, 16'd53146, 16'd12400, 16'd40371, 16'd49189, 16'd9987, 16'd49962, 16'd39355, 16'd21940, 16'd60354, 16'd4425, 16'd35490, 16'd25326, 16'd21879, 16'd17778, 16'd39821, 16'd49397, 16'd2409});
	test_expansion(128'h9828b18019d22720e465930824218b15, {16'd15634, 16'd21997, 16'd65100, 16'd34369, 16'd53024, 16'd19560, 16'd16446, 16'd29678, 16'd56754, 16'd62520, 16'd59570, 16'd33781, 16'd1882, 16'd38227, 16'd5122, 16'd50946, 16'd93, 16'd47114, 16'd16013, 16'd12472, 16'd7413, 16'd48017, 16'd24189, 16'd20593, 16'd21211, 16'd44328});
	test_expansion(128'h639e8dffc9ce3e162c00d63c59e2828d, {16'd63962, 16'd31512, 16'd12954, 16'd33385, 16'd21351, 16'd54035, 16'd32331, 16'd37658, 16'd27631, 16'd36911, 16'd11194, 16'd58838, 16'd18193, 16'd376, 16'd53769, 16'd50937, 16'd25079, 16'd63055, 16'd43154, 16'd45843, 16'd39550, 16'd23929, 16'd54912, 16'd560, 16'd3852, 16'd59664});
	test_expansion(128'h056f14e630ffe2740e06fd6b4ef69c4e, {16'd33771, 16'd20917, 16'd39826, 16'd41467, 16'd32908, 16'd52801, 16'd47284, 16'd56515, 16'd62480, 16'd30238, 16'd9443, 16'd59036, 16'd63232, 16'd52078, 16'd23481, 16'd8078, 16'd26, 16'd60463, 16'd64998, 16'd62523, 16'd31344, 16'd34553, 16'd9239, 16'd4925, 16'd20825, 16'd57});
	test_expansion(128'h375538491a101c7814de40093653d9ac, {16'd20896, 16'd26664, 16'd55770, 16'd17685, 16'd58242, 16'd25425, 16'd14066, 16'd53728, 16'd31493, 16'd16130, 16'd16087, 16'd19244, 16'd8615, 16'd29056, 16'd30251, 16'd61981, 16'd39443, 16'd42682, 16'd28218, 16'd14297, 16'd24594, 16'd35057, 16'd8624, 16'd54550, 16'd43655, 16'd25889});
	test_expansion(128'h274b26cbba48dd1af238c12bc77080a8, {16'd46873, 16'd17052, 16'd14956, 16'd3826, 16'd3867, 16'd36345, 16'd10198, 16'd16016, 16'd56203, 16'd51930, 16'd4825, 16'd33252, 16'd19946, 16'd49532, 16'd21880, 16'd47729, 16'd38802, 16'd3644, 16'd34533, 16'd60850, 16'd9901, 16'd11614, 16'd35436, 16'd26362, 16'd28128, 16'd6255});
	test_expansion(128'h7962596e2019cfe91d6592275de0e4fe, {16'd23938, 16'd57797, 16'd25003, 16'd56757, 16'd16339, 16'd21237, 16'd16002, 16'd22281, 16'd55433, 16'd31439, 16'd40978, 16'd19198, 16'd47248, 16'd31664, 16'd29509, 16'd48058, 16'd42176, 16'd53686, 16'd30397, 16'd34651, 16'd53104, 16'd44040, 16'd36760, 16'd47301, 16'd63156, 16'd35848});
	test_expansion(128'h1277b276a227364ff455a69798f72ce2, {16'd45245, 16'd10228, 16'd40860, 16'd42175, 16'd2845, 16'd35139, 16'd20693, 16'd20930, 16'd40385, 16'd39108, 16'd12418, 16'd51220, 16'd44329, 16'd63260, 16'd38367, 16'd11889, 16'd49993, 16'd46367, 16'd32100, 16'd36100, 16'd12428, 16'd5908, 16'd16376, 16'd64675, 16'd15850, 16'd47528});
	test_expansion(128'hc972a999a7a30f935cf4fde44000de9c, {16'd44377, 16'd45899, 16'd32601, 16'd56426, 16'd41880, 16'd40915, 16'd23070, 16'd51539, 16'd28981, 16'd20485, 16'd45738, 16'd18548, 16'd26808, 16'd25350, 16'd29958, 16'd16405, 16'd58885, 16'd59310, 16'd43766, 16'd64751, 16'd17517, 16'd5158, 16'd32495, 16'd54113, 16'd14778, 16'd41931});
	test_expansion(128'h236c45ce401f3e8bf98b09ad2ca4b0c9, {16'd6737, 16'd55662, 16'd9568, 16'd8816, 16'd516, 16'd55554, 16'd60976, 16'd25525, 16'd2641, 16'd25304, 16'd36292, 16'd3040, 16'd10954, 16'd19770, 16'd8680, 16'd64881, 16'd46130, 16'd11540, 16'd55494, 16'd12946, 16'd56547, 16'd3407, 16'd55419, 16'd34762, 16'd25324, 16'd61819});
	test_expansion(128'hf005f30b44ff7756b529dd0ab247fb0f, {16'd52383, 16'd22813, 16'd50628, 16'd23449, 16'd35478, 16'd36594, 16'd21532, 16'd31507, 16'd2504, 16'd58972, 16'd30182, 16'd36588, 16'd11239, 16'd7602, 16'd44925, 16'd2206, 16'd2412, 16'd13229, 16'd12707, 16'd36485, 16'd34295, 16'd32523, 16'd29015, 16'd24211, 16'd34560, 16'd24682});
	test_expansion(128'h2dd27be414acc7c0c9da4404c6f3dca1, {16'd36682, 16'd2094, 16'd42082, 16'd14476, 16'd59572, 16'd61373, 16'd38252, 16'd25281, 16'd18602, 16'd53669, 16'd17241, 16'd57511, 16'd43354, 16'd55255, 16'd20666, 16'd27284, 16'd22621, 16'd42785, 16'd11383, 16'd42967, 16'd13293, 16'd49889, 16'd31868, 16'd46523, 16'd27393, 16'd54672});
	test_expansion(128'h30f4597dac8e1e543767933f808d2318, {16'd47984, 16'd34036, 16'd39609, 16'd21901, 16'd11766, 16'd34618, 16'd33436, 16'd8215, 16'd55368, 16'd24224, 16'd30155, 16'd29646, 16'd31232, 16'd40418, 16'd63944, 16'd9759, 16'd39376, 16'd46193, 16'd27695, 16'd42495, 16'd41353, 16'd27659, 16'd148, 16'd27611, 16'd16018, 16'd23789});
	test_expansion(128'hf98665d29c9713cc4d371c297ee8cc12, {16'd2577, 16'd56674, 16'd2026, 16'd10865, 16'd28310, 16'd13758, 16'd18256, 16'd14176, 16'd36129, 16'd53694, 16'd35931, 16'd16608, 16'd14810, 16'd57380, 16'd34031, 16'd38897, 16'd356, 16'd27532, 16'd22151, 16'd64975, 16'd46028, 16'd30996, 16'd4531, 16'd57457, 16'd52860, 16'd31410});
	test_expansion(128'hb60f97173ec3d14a5772dc30420ed29e, {16'd46859, 16'd41568, 16'd45053, 16'd7970, 16'd19718, 16'd45722, 16'd29678, 16'd15379, 16'd64710, 16'd24121, 16'd20386, 16'd21436, 16'd51523, 16'd48475, 16'd21720, 16'd59957, 16'd501, 16'd3993, 16'd39658, 16'd29113, 16'd55188, 16'd43573, 16'd4170, 16'd10034, 16'd3289, 16'd55712});
	test_expansion(128'h8e55742660e65217bf95c8c53e182147, {16'd59355, 16'd60798, 16'd25387, 16'd15052, 16'd55881, 16'd2844, 16'd28437, 16'd5951, 16'd24581, 16'd10740, 16'd40413, 16'd2933, 16'd55983, 16'd164, 16'd48861, 16'd55693, 16'd54656, 16'd7939, 16'd19824, 16'd13150, 16'd30287, 16'd43441, 16'd35318, 16'd7552, 16'd20999, 16'd34080});
	test_expansion(128'he953345d21565c962014b13bc2b59a11, {16'd39508, 16'd54579, 16'd41008, 16'd7681, 16'd41702, 16'd62353, 16'd12069, 16'd56643, 16'd22366, 16'd7699, 16'd10922, 16'd21212, 16'd25496, 16'd65502, 16'd20530, 16'd18502, 16'd12388, 16'd30023, 16'd35909, 16'd38742, 16'd47075, 16'd14319, 16'd61196, 16'd45196, 16'd18679, 16'd13284});
	test_expansion(128'ha54d7015b050c74cb99d2b098f0094f6, {16'd20370, 16'd2588, 16'd50783, 16'd19692, 16'd38614, 16'd1060, 16'd32501, 16'd56510, 16'd19960, 16'd6027, 16'd29079, 16'd40625, 16'd62704, 16'd61346, 16'd58143, 16'd48929, 16'd59488, 16'd28488, 16'd49060, 16'd6589, 16'd5117, 16'd17280, 16'd10590, 16'd11622, 16'd29420, 16'd53055});
	test_expansion(128'h9aef7cc3537602f4995c09d31f66f28f, {16'd24683, 16'd45028, 16'd21850, 16'd6037, 16'd19142, 16'd9863, 16'd24444, 16'd24614, 16'd46425, 16'd44543, 16'd49038, 16'd41426, 16'd37893, 16'd11286, 16'd46377, 16'd13040, 16'd5113, 16'd2744, 16'd22946, 16'd25533, 16'd25927, 16'd34332, 16'd27020, 16'd16230, 16'd33146, 16'd10724});
	test_expansion(128'haf7f554047b907308585cdc5062b741e, {16'd10648, 16'd52638, 16'd46540, 16'd57588, 16'd22127, 16'd18729, 16'd16155, 16'd15532, 16'd20045, 16'd4796, 16'd11917, 16'd29534, 16'd9263, 16'd44821, 16'd49101, 16'd50717, 16'd56023, 16'd31911, 16'd36937, 16'd1276, 16'd3091, 16'd31349, 16'd28714, 16'd62412, 16'd45062, 16'd24589});
	test_expansion(128'ha80e1ab6fb248cfa8240fcd011e1abdd, {16'd28885, 16'd25647, 16'd23612, 16'd60535, 16'd36839, 16'd13399, 16'd52936, 16'd22989, 16'd5818, 16'd552, 16'd60703, 16'd64143, 16'd420, 16'd18906, 16'd15879, 16'd44485, 16'd52916, 16'd31285, 16'd36496, 16'd59825, 16'd58568, 16'd21802, 16'd40525, 16'd15699, 16'd57078, 16'd4773});
	test_expansion(128'h8e6f31fe1cc15f349a5c8e1465927b73, {16'd21040, 16'd29027, 16'd23202, 16'd59640, 16'd23744, 16'd40698, 16'd42700, 16'd40767, 16'd60849, 16'd51912, 16'd15101, 16'd11756, 16'd15910, 16'd10139, 16'd11669, 16'd47223, 16'd42053, 16'd5146, 16'd65025, 16'd43962, 16'd23615, 16'd14944, 16'd62993, 16'd13351, 16'd16735, 16'd64090});
	test_expansion(128'h05a543872427677546799b0c05a27a0c, {16'd64470, 16'd17758, 16'd1813, 16'd63535, 16'd41145, 16'd41520, 16'd42350, 16'd62832, 16'd30650, 16'd56855, 16'd18520, 16'd25065, 16'd19181, 16'd48369, 16'd12074, 16'd39840, 16'd18359, 16'd10593, 16'd34430, 16'd23006, 16'd49022, 16'd28129, 16'd34320, 16'd57095, 16'd60404, 16'd38083});
	test_expansion(128'h78610678a4f8072bb9e9ec6fd8c408ed, {16'd35020, 16'd18637, 16'd39294, 16'd54484, 16'd20353, 16'd15875, 16'd42295, 16'd61062, 16'd32337, 16'd13075, 16'd62923, 16'd34115, 16'd713, 16'd50144, 16'd59392, 16'd32436, 16'd17660, 16'd3017, 16'd23282, 16'd30973, 16'd16473, 16'd53936, 16'd334, 16'd16181, 16'd9955, 16'd58639});
	test_expansion(128'hcfda09aa77ca530357657f24cdd68df8, {16'd8065, 16'd29676, 16'd12447, 16'd54491, 16'd31553, 16'd22510, 16'd13727, 16'd3448, 16'd53993, 16'd21346, 16'd31283, 16'd41489, 16'd33055, 16'd19569, 16'd33937, 16'd62634, 16'd13770, 16'd26866, 16'd7509, 16'd4776, 16'd52822, 16'd48240, 16'd59805, 16'd23371, 16'd28457, 16'd52325});
	test_expansion(128'hf9b5ddff5fa0e9437a0c5147bf3297de, {16'd96, 16'd63572, 16'd37679, 16'd37564, 16'd6942, 16'd12251, 16'd60035, 16'd10014, 16'd10119, 16'd4391, 16'd19586, 16'd4463, 16'd9821, 16'd4614, 16'd52580, 16'd63672, 16'd18639, 16'd32437, 16'd37623, 16'd19033, 16'd57013, 16'd33721, 16'd4242, 16'd59060, 16'd5522, 16'd40273});
	test_expansion(128'h0cc54b78124343b42323290ac0a8300c, {16'd21570, 16'd37744, 16'd9715, 16'd59166, 16'd39682, 16'd13916, 16'd62555, 16'd51427, 16'd22412, 16'd52252, 16'd705, 16'd2056, 16'd62801, 16'd31220, 16'd12468, 16'd22413, 16'd19971, 16'd10090, 16'd42484, 16'd1704, 16'd35229, 16'd61570, 16'd36162, 16'd46951, 16'd64600, 16'd55681});
	test_expansion(128'h4a94cb9909182d1b82c6bf08f2fc6adb, {16'd22500, 16'd31211, 16'd37257, 16'd1916, 16'd32892, 16'd33658, 16'd8656, 16'd2781, 16'd59550, 16'd51043, 16'd31928, 16'd54875, 16'd62765, 16'd21119, 16'd28873, 16'd47419, 16'd63060, 16'd46481, 16'd34376, 16'd19661, 16'd32664, 16'd38472, 16'd33274, 16'd32349, 16'd22064, 16'd7990});
	test_expansion(128'h70914ce6c51af0fdd785296580e3f7d8, {16'd12056, 16'd12050, 16'd58067, 16'd40555, 16'd8429, 16'd21424, 16'd6665, 16'd44590, 16'd49282, 16'd16084, 16'd31796, 16'd56804, 16'd34106, 16'd33627, 16'd50306, 16'd32191, 16'd34332, 16'd31284, 16'd58567, 16'd20504, 16'd63869, 16'd11291, 16'd21905, 16'd49790, 16'd7749, 16'd23888});
	test_expansion(128'h83f95e0859a82d11e478cb52aad3df6b, {16'd59348, 16'd53044, 16'd41830, 16'd38218, 16'd9615, 16'd34092, 16'd65428, 16'd19732, 16'd14368, 16'd20389, 16'd39244, 16'd4863, 16'd45565, 16'd11276, 16'd50641, 16'd30560, 16'd6088, 16'd9630, 16'd26611, 16'd15930, 16'd3570, 16'd57495, 16'd59740, 16'd47814, 16'd34834, 16'd57743});
	test_expansion(128'he8582381218fa00f8566425557288886, {16'd20655, 16'd9787, 16'd41423, 16'd30046, 16'd47734, 16'd54699, 16'd33333, 16'd14118, 16'd44, 16'd59150, 16'd17973, 16'd14074, 16'd34179, 16'd61384, 16'd7097, 16'd57580, 16'd32105, 16'd43046, 16'd56136, 16'd59233, 16'd1254, 16'd32873, 16'd62573, 16'd1758, 16'd34302, 16'd59676});
	test_expansion(128'hd78eca72a5732088b4d541f53ae5e97f, {16'd52579, 16'd46580, 16'd26108, 16'd8853, 16'd17650, 16'd13203, 16'd2332, 16'd58901, 16'd37833, 16'd37388, 16'd19229, 16'd54967, 16'd46943, 16'd37657, 16'd47476, 16'd33420, 16'd64589, 16'd21243, 16'd54133, 16'd29559, 16'd9386, 16'd36532, 16'd46543, 16'd39780, 16'd36080, 16'd59944});
	test_expansion(128'hd46dc10567226ba6da8d879da13e8686, {16'd25775, 16'd40208, 16'd23933, 16'd64596, 16'd26389, 16'd64914, 16'd27474, 16'd35747, 16'd1496, 16'd46863, 16'd54445, 16'd7472, 16'd2055, 16'd34363, 16'd61960, 16'd19331, 16'd60422, 16'd30659, 16'd27917, 16'd16501, 16'd56210, 16'd5697, 16'd5662, 16'd21479, 16'd62389, 16'd55669});
	test_expansion(128'hab8c2dc8e91fb27519f1f4dd32246107, {16'd1530, 16'd61051, 16'd63422, 16'd32521, 16'd35293, 16'd41551, 16'd53350, 16'd1108, 16'd52238, 16'd24324, 16'd5343, 16'd16782, 16'd56543, 16'd61604, 16'd13321, 16'd20195, 16'd32491, 16'd32296, 16'd19056, 16'd60958, 16'd21554, 16'd9356, 16'd36390, 16'd50785, 16'd2432, 16'd5209});
	test_expansion(128'h5ad432c8ea19d2eb90c67489af7198fb, {16'd38673, 16'd44016, 16'd63732, 16'd28986, 16'd47300, 16'd50949, 16'd28857, 16'd17579, 16'd45790, 16'd65131, 16'd26568, 16'd42850, 16'd10682, 16'd58342, 16'd28458, 16'd42088, 16'd3276, 16'd29697, 16'd14300, 16'd8800, 16'd10694, 16'd45799, 16'd17625, 16'd27381, 16'd50545, 16'd60321});
	test_expansion(128'h1884c62535fcdda2c243da4aa9f31e9a, {16'd5699, 16'd3838, 16'd10380, 16'd16142, 16'd62136, 16'd56744, 16'd48652, 16'd20118, 16'd26231, 16'd37345, 16'd14021, 16'd49804, 16'd54094, 16'd21279, 16'd59320, 16'd51967, 16'd64913, 16'd43961, 16'd12277, 16'd14448, 16'd39785, 16'd41262, 16'd16342, 16'd41869, 16'd33636, 16'd31272});
	test_expansion(128'hffed784f4b8aba82ef829a63e950c005, {16'd64571, 16'd25330, 16'd45777, 16'd20703, 16'd46273, 16'd26659, 16'd18778, 16'd2527, 16'd54911, 16'd8594, 16'd19340, 16'd53848, 16'd2936, 16'd51211, 16'd42875, 16'd15364, 16'd23474, 16'd56171, 16'd15638, 16'd9550, 16'd47161, 16'd27697, 16'd34120, 16'd30466, 16'd53501, 16'd2087});
	test_expansion(128'hac11aac26fbc084ca18a06238995dd67, {16'd61835, 16'd20309, 16'd63637, 16'd51989, 16'd48789, 16'd46414, 16'd14406, 16'd22816, 16'd15751, 16'd63666, 16'd32670, 16'd59917, 16'd49375, 16'd19202, 16'd16460, 16'd58435, 16'd49975, 16'd35869, 16'd34707, 16'd25826, 16'd9315, 16'd9027, 16'd6641, 16'd35510, 16'd58685, 16'd41453});
	test_expansion(128'h993424d8e933f9107a61dd85015ab61b, {16'd36119, 16'd39831, 16'd8664, 16'd24234, 16'd55191, 16'd54247, 16'd22047, 16'd17871, 16'd25779, 16'd20928, 16'd28489, 16'd28261, 16'd46544, 16'd7760, 16'd749, 16'd60479, 16'd1194, 16'd17818, 16'd22909, 16'd46402, 16'd62467, 16'd42101, 16'd64744, 16'd17111, 16'd16468, 16'd47926});
	test_expansion(128'hbdef5ae8386116188cb52a1141f0380a, {16'd13604, 16'd22174, 16'd42071, 16'd43806, 16'd56692, 16'd45180, 16'd23964, 16'd5995, 16'd4863, 16'd29943, 16'd31178, 16'd15692, 16'd34764, 16'd33742, 16'd25947, 16'd3219, 16'd14060, 16'd41447, 16'd10542, 16'd265, 16'd6283, 16'd64823, 16'd53594, 16'd62572, 16'd10234, 16'd28077});
	test_expansion(128'h9276ad3431768a4d0822f4489e008ac4, {16'd29341, 16'd57350, 16'd14323, 16'd60002, 16'd9408, 16'd2732, 16'd30294, 16'd53094, 16'd36908, 16'd45945, 16'd45200, 16'd46423, 16'd48331, 16'd61566, 16'd56563, 16'd34673, 16'd19633, 16'd11200, 16'd53894, 16'd49312, 16'd42404, 16'd48566, 16'd7686, 16'd32470, 16'd11941, 16'd49212});
	test_expansion(128'h2d1a6718e05cdabd786a877244f97311, {16'd3038, 16'd55441, 16'd26010, 16'd6486, 16'd62973, 16'd804, 16'd4494, 16'd51629, 16'd58099, 16'd56630, 16'd47316, 16'd38100, 16'd12685, 16'd46577, 16'd8368, 16'd20963, 16'd32294, 16'd26326, 16'd40897, 16'd13283, 16'd15815, 16'd39601, 16'd58340, 16'd54107, 16'd15425, 16'd6005});
	test_expansion(128'h2fe7700cdf9b6bf96cb50be90a24004a, {16'd57718, 16'd3127, 16'd262, 16'd30456, 16'd30595, 16'd9594, 16'd45728, 16'd37736, 16'd44038, 16'd44774, 16'd529, 16'd21299, 16'd48483, 16'd37838, 16'd14255, 16'd65467, 16'd33471, 16'd14938, 16'd10174, 16'd59092, 16'd21196, 16'd50123, 16'd21952, 16'd48031, 16'd8658, 16'd4605});
	test_expansion(128'haca640295e135e570cdd71b896422a48, {16'd31227, 16'd51434, 16'd5807, 16'd57411, 16'd54070, 16'd43024, 16'd28297, 16'd61635, 16'd44482, 16'd44220, 16'd41217, 16'd64160, 16'd64797, 16'd35489, 16'd58296, 16'd46200, 16'd2289, 16'd59080, 16'd43402, 16'd30703, 16'd45769, 16'd11935, 16'd31550, 16'd39744, 16'd37627, 16'd43975});
	test_expansion(128'h162116d339f43efa70d417de99b107fb, {16'd59343, 16'd1568, 16'd31216, 16'd12682, 16'd35570, 16'd20878, 16'd37435, 16'd46911, 16'd20497, 16'd33302, 16'd21607, 16'd14426, 16'd25464, 16'd50232, 16'd13195, 16'd2821, 16'd24469, 16'd64119, 16'd51956, 16'd35413, 16'd25269, 16'd53487, 16'd10922, 16'd57981, 16'd21220, 16'd61721});
	test_expansion(128'h91039781a4ce11239e849702cfb7128e, {16'd52519, 16'd60603, 16'd4902, 16'd44153, 16'd49231, 16'd54702, 16'd61254, 16'd40650, 16'd32279, 16'd3291, 16'd3175, 16'd49139, 16'd46324, 16'd48471, 16'd48543, 16'd30101, 16'd27393, 16'd30931, 16'd41983, 16'd62932, 16'd435, 16'd59056, 16'd3253, 16'd31836, 16'd13672, 16'd19890});
	test_expansion(128'h7ec758c0ed60d31414ac029eaf0b5ca2, {16'd22210, 16'd39543, 16'd56214, 16'd28944, 16'd26237, 16'd59528, 16'd11051, 16'd5093, 16'd12285, 16'd10430, 16'd22819, 16'd15575, 16'd38685, 16'd10240, 16'd37154, 16'd8754, 16'd64171, 16'd30377, 16'd49409, 16'd24291, 16'd57651, 16'd21, 16'd9781, 16'd62689, 16'd35319, 16'd40357});
	test_expansion(128'h6b2370b98c552c9f46097e93fc564700, {16'd39263, 16'd14809, 16'd46681, 16'd11960, 16'd24208, 16'd39821, 16'd57767, 16'd49702, 16'd62369, 16'd38988, 16'd6300, 16'd12025, 16'd33068, 16'd18189, 16'd32628, 16'd3228, 16'd43285, 16'd59002, 16'd63343, 16'd18577, 16'd48678, 16'd17405, 16'd58566, 16'd5147, 16'd63387, 16'd61545});
	test_expansion(128'hac97419dd89366ed90d428d7e0722a10, {16'd584, 16'd9484, 16'd16640, 16'd62518, 16'd15217, 16'd44119, 16'd18200, 16'd6031, 16'd13821, 16'd25561, 16'd30527, 16'd48419, 16'd53303, 16'd42357, 16'd27055, 16'd5470, 16'd21863, 16'd21489, 16'd709, 16'd62517, 16'd10642, 16'd57091, 16'd58402, 16'd22342, 16'd52697, 16'd10975});
	test_expansion(128'hf48778e33004c798c1b3f371090ba24d, {16'd63231, 16'd61602, 16'd46875, 16'd59862, 16'd19125, 16'd38038, 16'd13710, 16'd55423, 16'd63842, 16'd19947, 16'd31279, 16'd49611, 16'd11057, 16'd60407, 16'd38071, 16'd61809, 16'd46894, 16'd8148, 16'd54520, 16'd52757, 16'd16467, 16'd19153, 16'd7529, 16'd12807, 16'd10501, 16'd26696});
	test_expansion(128'h74f983083fdd85d4b38dde6e57223cfc, {16'd62201, 16'd8082, 16'd59887, 16'd34674, 16'd57614, 16'd30622, 16'd57419, 16'd39832, 16'd56503, 16'd64940, 16'd42818, 16'd56420, 16'd41862, 16'd4173, 16'd39661, 16'd9704, 16'd33197, 16'd9943, 16'd27332, 16'd43327, 16'd31484, 16'd10740, 16'd58721, 16'd64566, 16'd24086, 16'd55182});
	test_expansion(128'he05cca31c72aa6628a2e784198b0a4e8, {16'd61099, 16'd7401, 16'd11980, 16'd11313, 16'd3128, 16'd48596, 16'd28800, 16'd2705, 16'd607, 16'd17819, 16'd59092, 16'd16107, 16'd27187, 16'd15440, 16'd44706, 16'd39217, 16'd42845, 16'd12351, 16'd39065, 16'd52878, 16'd19271, 16'd20543, 16'd50254, 16'd4276, 16'd60791, 16'd30740});
	test_expansion(128'hcbef24295fcfc273a19a6f1ec5802f98, {16'd58194, 16'd13135, 16'd46885, 16'd13201, 16'd40555, 16'd4743, 16'd57206, 16'd35303, 16'd26656, 16'd28525, 16'd25157, 16'd52223, 16'd46849, 16'd51905, 16'd9964, 16'd18551, 16'd51480, 16'd8921, 16'd38861, 16'd53696, 16'd44189, 16'd18187, 16'd33557, 16'd53646, 16'd62555, 16'd54501});
	test_expansion(128'he7c2c0496bc00a3f58596524e39dd7f6, {16'd63736, 16'd27748, 16'd45381, 16'd53997, 16'd14374, 16'd6885, 16'd19862, 16'd52258, 16'd39880, 16'd38964, 16'd36469, 16'd2560, 16'd1194, 16'd51732, 16'd4135, 16'd1945, 16'd36170, 16'd30373, 16'd4570, 16'd57933, 16'd14401, 16'd47855, 16'd48948, 16'd39176, 16'd49029, 16'd15329});
	test_expansion(128'he493366841ff5a27e3ab26e07414d3c4, {16'd30279, 16'd47183, 16'd8001, 16'd44136, 16'd11967, 16'd58457, 16'd12749, 16'd21468, 16'd19385, 16'd3253, 16'd5269, 16'd15194, 16'd20177, 16'd57007, 16'd46229, 16'd29119, 16'd41107, 16'd57677, 16'd47949, 16'd46889, 16'd41925, 16'd13239, 16'd31815, 16'd57941, 16'd34628, 16'd3018});
	test_expansion(128'h21f5d192fe79d820ff6214fbdcbce6e8, {16'd60140, 16'd52711, 16'd13399, 16'd21791, 16'd18026, 16'd34539, 16'd15201, 16'd15390, 16'd29140, 16'd33026, 16'd15838, 16'd38264, 16'd5551, 16'd37232, 16'd45658, 16'd11577, 16'd42601, 16'd19905, 16'd25832, 16'd63275, 16'd32382, 16'd3121, 16'd63559, 16'd58784, 16'd41561, 16'd63723});
	test_expansion(128'h9754a25d820b628fcf4b8d7de3ec6267, {16'd32419, 16'd5792, 16'd51194, 16'd11684, 16'd47701, 16'd55139, 16'd8329, 16'd49324, 16'd19368, 16'd64597, 16'd13733, 16'd41442, 16'd44011, 16'd18107, 16'd13543, 16'd3074, 16'd50957, 16'd47112, 16'd43120, 16'd43700, 16'd9441, 16'd34656, 16'd22724, 16'd49105, 16'd50734, 16'd32720});
	test_expansion(128'hfe3f42629b19d93654c70207bab43d01, {16'd45467, 16'd63540, 16'd41656, 16'd64189, 16'd53696, 16'd1859, 16'd34177, 16'd63872, 16'd26703, 16'd29346, 16'd41153, 16'd46886, 16'd23204, 16'd37119, 16'd56592, 16'd33530, 16'd52679, 16'd20622, 16'd15829, 16'd13483, 16'd45882, 16'd28643, 16'd17382, 16'd217, 16'd16525, 16'd58756});
	test_expansion(128'h5c8bb33773661b2c2cc9a7d668682ba5, {16'd64345, 16'd5220, 16'd41374, 16'd16898, 16'd30358, 16'd4756, 16'd15669, 16'd48779, 16'd49571, 16'd14834, 16'd4660, 16'd15052, 16'd58599, 16'd63478, 16'd25963, 16'd29883, 16'd52817, 16'd4637, 16'd1801, 16'd13150, 16'd17796, 16'd52479, 16'd61318, 16'd17807, 16'd54068, 16'd63873});
	test_expansion(128'h3aaa714037c1487360f4b1c428ccc2e6, {16'd55681, 16'd46002, 16'd25965, 16'd29291, 16'd53131, 16'd6701, 16'd44271, 16'd22282, 16'd16685, 16'd35018, 16'd19482, 16'd51900, 16'd1897, 16'd44874, 16'd9805, 16'd4571, 16'd46637, 16'd26666, 16'd49337, 16'd53141, 16'd17694, 16'd20181, 16'd39672, 16'd9588, 16'd13960, 16'd22764});
	test_expansion(128'hdc54e5a598ecfba84d55a07dd435a483, {16'd32087, 16'd47592, 16'd62845, 16'd41755, 16'd7485, 16'd17506, 16'd28989, 16'd47872, 16'd37365, 16'd49298, 16'd8593, 16'd64793, 16'd40217, 16'd29344, 16'd11029, 16'd15633, 16'd23493, 16'd32162, 16'd45591, 16'd31142, 16'd38080, 16'd10904, 16'd28109, 16'd7000, 16'd15592, 16'd46312});
	test_expansion(128'h5343b1193fb096f183a0fa092e5b5137, {16'd48230, 16'd47693, 16'd39197, 16'd40976, 16'd19527, 16'd4492, 16'd28550, 16'd25380, 16'd33807, 16'd52130, 16'd56447, 16'd29629, 16'd44395, 16'd32962, 16'd8659, 16'd63256, 16'd53255, 16'd3540, 16'd31043, 16'd14225, 16'd11498, 16'd33964, 16'd35894, 16'd23889, 16'd46729, 16'd26175});
	test_expansion(128'hc8470606502681d4e8115faeecd43d5b, {16'd40259, 16'd19144, 16'd30107, 16'd39213, 16'd43792, 16'd17657, 16'd4059, 16'd39958, 16'd16372, 16'd52544, 16'd2074, 16'd30825, 16'd21090, 16'd30590, 16'd38280, 16'd23424, 16'd41650, 16'd6876, 16'd65449, 16'd34879, 16'd1328, 16'd31770, 16'd51111, 16'd21285, 16'd63690, 16'd56822});
	test_expansion(128'h08cb8a2b74d9c088641928ef7fc2fd28, {16'd57557, 16'd1223, 16'd58893, 16'd28599, 16'd4018, 16'd42382, 16'd53828, 16'd56786, 16'd18776, 16'd31454, 16'd37185, 16'd26519, 16'd12500, 16'd44988, 16'd24252, 16'd55220, 16'd62102, 16'd64840, 16'd53038, 16'd57732, 16'd26320, 16'd26647, 16'd42022, 16'd55444, 16'd28791, 16'd60074});
	test_expansion(128'hae42c51b95316cb15b675e5288541109, {16'd48729, 16'd45931, 16'd62339, 16'd28234, 16'd54435, 16'd48271, 16'd6218, 16'd54985, 16'd49567, 16'd33495, 16'd29426, 16'd25536, 16'd20205, 16'd5228, 16'd52888, 16'd25858, 16'd17850, 16'd35477, 16'd31747, 16'd53047, 16'd6117, 16'd9265, 16'd55440, 16'd65319, 16'd8535, 16'd46297});
	test_expansion(128'h49406dadd89fdf1de920011ef333e51b, {16'd26011, 16'd58283, 16'd5324, 16'd29993, 16'd42601, 16'd2766, 16'd49087, 16'd41984, 16'd37775, 16'd44312, 16'd53084, 16'd59125, 16'd56402, 16'd35375, 16'd49229, 16'd24363, 16'd31321, 16'd13041, 16'd7429, 16'd61593, 16'd61612, 16'd62970, 16'd31682, 16'd19117, 16'd43732, 16'd13788});
	test_expansion(128'hc2d0e4d3541ca566cce19f32bcc52cb9, {16'd15902, 16'd13578, 16'd20469, 16'd52972, 16'd52518, 16'd60976, 16'd63560, 16'd65175, 16'd22594, 16'd50343, 16'd12532, 16'd14483, 16'd58655, 16'd63559, 16'd31272, 16'd55433, 16'd50077, 16'd17504, 16'd21664, 16'd50816, 16'd5399, 16'd5287, 16'd24142, 16'd46186, 16'd31731, 16'd2451});
	test_expansion(128'h24aacead4c6b1e97e3dfc8cabd0b7011, {16'd35558, 16'd38763, 16'd60163, 16'd41301, 16'd1633, 16'd11013, 16'd13285, 16'd31924, 16'd63986, 16'd54724, 16'd47575, 16'd37692, 16'd54976, 16'd47593, 16'd25323, 16'd2932, 16'd45236, 16'd34588, 16'd54100, 16'd21318, 16'd313, 16'd12854, 16'd15698, 16'd59118, 16'd37531, 16'd11810});
	test_expansion(128'hdf8bca334a190fc207b037e0e14d6b67, {16'd12170, 16'd5341, 16'd27903, 16'd6447, 16'd9629, 16'd49119, 16'd20237, 16'd39329, 16'd29835, 16'd25826, 16'd51112, 16'd54594, 16'd22602, 16'd59481, 16'd62286, 16'd38283, 16'd17300, 16'd9027, 16'd37726, 16'd35381, 16'd29956, 16'd62307, 16'd5802, 16'd50797, 16'd4188, 16'd20268});
	test_expansion(128'hfd00d599032702a10424057ebf22285f, {16'd12414, 16'd4024, 16'd38419, 16'd5712, 16'd20665, 16'd29617, 16'd49276, 16'd47247, 16'd19121, 16'd81, 16'd46685, 16'd50066, 16'd24338, 16'd9229, 16'd9781, 16'd36628, 16'd23990, 16'd18386, 16'd22574, 16'd44059, 16'd7917, 16'd1598, 16'd29253, 16'd31007, 16'd28410, 16'd15412});
	test_expansion(128'h8a1e2821da3c3666d152f14610bf291c, {16'd52460, 16'd42588, 16'd32796, 16'd715, 16'd46215, 16'd57845, 16'd11568, 16'd2521, 16'd48734, 16'd52043, 16'd32070, 16'd48878, 16'd46341, 16'd9366, 16'd28638, 16'd52686, 16'd23960, 16'd39296, 16'd60153, 16'd39530, 16'd42071, 16'd53584, 16'd51015, 16'd52405, 16'd60784, 16'd12584});
	test_expansion(128'h700dc4e9c6b927d94eec65acdf48db95, {16'd51069, 16'd42954, 16'd8704, 16'd17047, 16'd3141, 16'd26481, 16'd24655, 16'd47219, 16'd37054, 16'd42624, 16'd5402, 16'd404, 16'd16188, 16'd16920, 16'd25891, 16'd46240, 16'd13658, 16'd12255, 16'd38685, 16'd14605, 16'd44979, 16'd40714, 16'd53251, 16'd23506, 16'd16616, 16'd37109});
	test_expansion(128'h1455ba0d2f0fe17d27fa96041818989a, {16'd63387, 16'd14969, 16'd38962, 16'd49203, 16'd16311, 16'd50612, 16'd32238, 16'd14517, 16'd13645, 16'd62466, 16'd48448, 16'd55855, 16'd38288, 16'd33308, 16'd41459, 16'd39161, 16'd21414, 16'd57089, 16'd4445, 16'd803, 16'd50383, 16'd52985, 16'd54352, 16'd5221, 16'd55312, 16'd17214});
	test_expansion(128'h1330044a8cc148b5bfc0bcb66ea260c0, {16'd48942, 16'd57330, 16'd10780, 16'd49432, 16'd52837, 16'd49293, 16'd50494, 16'd57962, 16'd61083, 16'd49548, 16'd44228, 16'd9358, 16'd10814, 16'd58588, 16'd43925, 16'd31100, 16'd12913, 16'd34742, 16'd52254, 16'd50269, 16'd22297, 16'd3491, 16'd53635, 16'd21168, 16'd11900, 16'd20618});
	test_expansion(128'h73776cfeddfbe67cb2c03b983823e2e3, {16'd57506, 16'd64724, 16'd26495, 16'd1488, 16'd29537, 16'd4409, 16'd29492, 16'd17570, 16'd27669, 16'd49625, 16'd5698, 16'd21616, 16'd27952, 16'd55080, 16'd23424, 16'd615, 16'd52496, 16'd34293, 16'd11719, 16'd4133, 16'd23534, 16'd47522, 16'd42927, 16'd55754, 16'd42006, 16'd10638});
	test_expansion(128'hf3c6bcdc5ec677d8e3e7f3bc05ec406d, {16'd5397, 16'd20127, 16'd57523, 16'd47873, 16'd14641, 16'd31880, 16'd64667, 16'd4729, 16'd5162, 16'd63812, 16'd48177, 16'd2536, 16'd38191, 16'd889, 16'd53265, 16'd16163, 16'd26898, 16'd30477, 16'd58986, 16'd5222, 16'd21838, 16'd51675, 16'd36394, 16'd64699, 16'd42467, 16'd27843});
	test_expansion(128'h5f9a10b23880e64accfd257a17cfc940, {16'd54887, 16'd60976, 16'd36224, 16'd16618, 16'd45907, 16'd24635, 16'd40182, 16'd26612, 16'd42748, 16'd40824, 16'd29971, 16'd33216, 16'd57807, 16'd9050, 16'd42053, 16'd45170, 16'd26345, 16'd1355, 16'd33847, 16'd47048, 16'd62264, 16'd48256, 16'd41024, 16'd28829, 16'd50383, 16'd59144});
	test_expansion(128'h188b7bc81585246ebbb2e714f36442f0, {16'd5320, 16'd37950, 16'd44627, 16'd15165, 16'd42606, 16'd17815, 16'd1421, 16'd7630, 16'd58631, 16'd5454, 16'd57973, 16'd43251, 16'd51098, 16'd40896, 16'd2055, 16'd37041, 16'd61502, 16'd9334, 16'd43054, 16'd41777, 16'd53297, 16'd40632, 16'd4722, 16'd34335, 16'd8379, 16'd6051});
	test_expansion(128'h67b2bd9b686e830e7d1fee6bb939b1f5, {16'd3014, 16'd32719, 16'd56992, 16'd35854, 16'd8530, 16'd65016, 16'd63978, 16'd24535, 16'd6673, 16'd8521, 16'd13184, 16'd23503, 16'd15628, 16'd5383, 16'd22655, 16'd33578, 16'd33523, 16'd29333, 16'd2766, 16'd45837, 16'd60136, 16'd49025, 16'd35287, 16'd40115, 16'd28359, 16'd46600});
	test_expansion(128'h91cc7c5d0f770f4dc2de76e214457aab, {16'd6917, 16'd63380, 16'd39513, 16'd47139, 16'd63045, 16'd27877, 16'd62201, 16'd62706, 16'd16214, 16'd58006, 16'd65087, 16'd28953, 16'd4688, 16'd60653, 16'd38779, 16'd24981, 16'd11584, 16'd62754, 16'd42647, 16'd54312, 16'd56863, 16'd37939, 16'd20602, 16'd16455, 16'd58587, 16'd9206});
	test_expansion(128'h59c9eb3371911222b59f2c80c5bd867c, {16'd55537, 16'd37520, 16'd15106, 16'd50428, 16'd56495, 16'd54181, 16'd23681, 16'd45291, 16'd44287, 16'd42886, 16'd7506, 16'd49208, 16'd27954, 16'd32923, 16'd34381, 16'd19818, 16'd18128, 16'd31047, 16'd33493, 16'd47596, 16'd3052, 16'd18035, 16'd23764, 16'd46863, 16'd43774, 16'd6626});
	test_expansion(128'h153034a573b1cd841edcb408fbf760dd, {16'd1765, 16'd25172, 16'd45010, 16'd6208, 16'd40972, 16'd63859, 16'd31658, 16'd31439, 16'd34650, 16'd34793, 16'd44741, 16'd33232, 16'd51456, 16'd58633, 16'd57387, 16'd8693, 16'd34307, 16'd53534, 16'd5913, 16'd8741, 16'd22132, 16'd18412, 16'd30839, 16'd58041, 16'd29171, 16'd47298});
	test_expansion(128'hdb1eb3676a8c61f0ed404295040a4e01, {16'd34205, 16'd27657, 16'd33761, 16'd41942, 16'd35994, 16'd9389, 16'd25464, 16'd13087, 16'd57001, 16'd13130, 16'd28525, 16'd12989, 16'd58645, 16'd45524, 16'd2226, 16'd1959, 16'd30318, 16'd19744, 16'd3685, 16'd2683, 16'd18187, 16'd49935, 16'd39748, 16'd17525, 16'd13526, 16'd26651});
	test_expansion(128'hb0e6d38aba53cd27511abb0423b4991e, {16'd15179, 16'd31182, 16'd36238, 16'd18499, 16'd24715, 16'd31063, 16'd25936, 16'd3679, 16'd58084, 16'd43971, 16'd62735, 16'd11414, 16'd59712, 16'd13884, 16'd3982, 16'd62811, 16'd6994, 16'd44003, 16'd3545, 16'd27872, 16'd25042, 16'd56476, 16'd12112, 16'd46939, 16'd20678, 16'd20076});
	test_expansion(128'h23de8d3b50f7642c7b8b615031a71616, {16'd22851, 16'd24289, 16'd8453, 16'd35925, 16'd19367, 16'd58780, 16'd44156, 16'd1979, 16'd59437, 16'd58363, 16'd37667, 16'd22208, 16'd44678, 16'd19979, 16'd24688, 16'd46981, 16'd7095, 16'd36574, 16'd22923, 16'd42905, 16'd55899, 16'd13490, 16'd39479, 16'd5219, 16'd48933, 16'd18785});
	test_expansion(128'h9fd4fee96837b39159b25cc1a36e42b4, {16'd11109, 16'd6331, 16'd30216, 16'd31720, 16'd46980, 16'd56966, 16'd55280, 16'd9291, 16'd52097, 16'd30346, 16'd60563, 16'd48477, 16'd43187, 16'd39516, 16'd621, 16'd36242, 16'd63130, 16'd10214, 16'd46188, 16'd24974, 16'd62997, 16'd39218, 16'd16823, 16'd29399, 16'd27376, 16'd30030});
	test_expansion(128'h2b6493c199005a32605ac30381a32fee, {16'd30648, 16'd28330, 16'd55934, 16'd660, 16'd24358, 16'd435, 16'd13515, 16'd19322, 16'd13873, 16'd47766, 16'd9732, 16'd43144, 16'd1471, 16'd48166, 16'd38592, 16'd27066, 16'd19463, 16'd42318, 16'd48111, 16'd12670, 16'd53959, 16'd11320, 16'd29152, 16'd59436, 16'd20266, 16'd35866});
	test_expansion(128'h6d9db5afb74edfd7d66b08354d8cbf7a, {16'd48734, 16'd58315, 16'd53923, 16'd34188, 16'd25285, 16'd27633, 16'd16706, 16'd23535, 16'd20936, 16'd14892, 16'd57976, 16'd49664, 16'd20405, 16'd41366, 16'd28436, 16'd7374, 16'd11107, 16'd36466, 16'd4408, 16'd22636, 16'd18495, 16'd45620, 16'd26849, 16'd13334, 16'd54407, 16'd44430});
	test_expansion(128'hfd54f9abf93177695208f2d0d4d2fabf, {16'd19437, 16'd17272, 16'd10126, 16'd26164, 16'd11079, 16'd8881, 16'd49571, 16'd22764, 16'd11223, 16'd44095, 16'd57283, 16'd55102, 16'd26925, 16'd56721, 16'd11349, 16'd36911, 16'd53667, 16'd48094, 16'd46004, 16'd45199, 16'd57880, 16'd46761, 16'd54852, 16'd43228, 16'd33754, 16'd16891});
	test_expansion(128'hdd099b736792211d53886e8e01b492e8, {16'd18093, 16'd16481, 16'd2546, 16'd44356, 16'd57043, 16'd18928, 16'd27719, 16'd17153, 16'd28731, 16'd23876, 16'd8926, 16'd4307, 16'd20700, 16'd50014, 16'd5097, 16'd53684, 16'd46170, 16'd51996, 16'd24875, 16'd16646, 16'd28352, 16'd4835, 16'd4602, 16'd57849, 16'd23135, 16'd51095});
	test_expansion(128'hb9ec33c6a37dc7edd548c6b6e6cfda51, {16'd57637, 16'd48944, 16'd33054, 16'd35664, 16'd31228, 16'd17498, 16'd13357, 16'd65414, 16'd65392, 16'd10069, 16'd38410, 16'd32747, 16'd63600, 16'd56420, 16'd4736, 16'd42176, 16'd37723, 16'd60334, 16'd36125, 16'd44248, 16'd40327, 16'd5167, 16'd51155, 16'd58944, 16'd29203, 16'd412});
	test_expansion(128'h3087884fb6ab39eef46e76c6b4b6d45a, {16'd8569, 16'd4594, 16'd54180, 16'd58259, 16'd49538, 16'd21142, 16'd8210, 16'd15394, 16'd61154, 16'd31274, 16'd62158, 16'd52744, 16'd41572, 16'd35281, 16'd20834, 16'd49400, 16'd57415, 16'd51802, 16'd22426, 16'd54078, 16'd9705, 16'd44971, 16'd46595, 16'd62088, 16'd65491, 16'd64407});
	test_expansion(128'h8f2b1f1a44af69d4137e71e6edd59ee4, {16'd15967, 16'd29996, 16'd34218, 16'd31893, 16'd48000, 16'd24064, 16'd64488, 16'd13894, 16'd5603, 16'd62452, 16'd9699, 16'd37097, 16'd50974, 16'd22094, 16'd52757, 16'd23476, 16'd1216, 16'd57337, 16'd42577, 16'd37678, 16'd22712, 16'd48553, 16'd7932, 16'd42734, 16'd54269, 16'd19792});
	test_expansion(128'h0f7cbc262d64c16bc64d6f8706c84c1a, {16'd26196, 16'd20832, 16'd60427, 16'd54776, 16'd38054, 16'd52676, 16'd22104, 16'd10463, 16'd63898, 16'd9478, 16'd44793, 16'd25966, 16'd42609, 16'd4679, 16'd30010, 16'd42729, 16'd11203, 16'd49407, 16'd24363, 16'd64124, 16'd50333, 16'd28666, 16'd5548, 16'd9268, 16'd2646, 16'd11007});
	test_expansion(128'h54d0b210a0944e0f52373502173741f0, {16'd13266, 16'd29906, 16'd16674, 16'd12783, 16'd62028, 16'd43228, 16'd50673, 16'd21157, 16'd3162, 16'd35503, 16'd24969, 16'd14494, 16'd47268, 16'd58371, 16'd39618, 16'd47544, 16'd60068, 16'd36279, 16'd38474, 16'd33312, 16'd23672, 16'd58115, 16'd14603, 16'd56797, 16'd1832, 16'd64430});
	test_expansion(128'h57dd6c53dc1cf6bce34f19583e555019, {16'd51774, 16'd21680, 16'd2302, 16'd49167, 16'd5014, 16'd5734, 16'd18801, 16'd5997, 16'd18107, 16'd7526, 16'd44466, 16'd34292, 16'd5912, 16'd12301, 16'd62041, 16'd2208, 16'd15753, 16'd42250, 16'd2230, 16'd38004, 16'd18846, 16'd35597, 16'd47967, 16'd59911, 16'd59109, 16'd16787});
	test_expansion(128'h4f726051ca1e95547948185f62baab4b, {16'd24990, 16'd52563, 16'd33729, 16'd39159, 16'd45877, 16'd46067, 16'd60737, 16'd20326, 16'd17319, 16'd26190, 16'd49888, 16'd32923, 16'd765, 16'd64857, 16'd56317, 16'd828, 16'd33447, 16'd45144, 16'd31175, 16'd57530, 16'd693, 16'd43382, 16'd12916, 16'd15549, 16'd52676, 16'd61346});
	test_expansion(128'hc1991d54b575c9cd2de33c671be62d36, {16'd59005, 16'd52233, 16'd44969, 16'd21730, 16'd10233, 16'd9906, 16'd55678, 16'd7682, 16'd62305, 16'd38291, 16'd65535, 16'd13193, 16'd30292, 16'd64530, 16'd25712, 16'd0, 16'd62245, 16'd1149, 16'd21243, 16'd194, 16'd3891, 16'd16104, 16'd33882, 16'd28985, 16'd27789, 16'd26096});
	test_expansion(128'h30ec0512f4addc2b11e961497a50e2bd, {16'd3086, 16'd57974, 16'd62014, 16'd64464, 16'd64511, 16'd24789, 16'd59249, 16'd17562, 16'd36412, 16'd33729, 16'd19262, 16'd11561, 16'd16813, 16'd30489, 16'd19957, 16'd51123, 16'd41558, 16'd3421, 16'd43302, 16'd481, 16'd5432, 16'd25099, 16'd38203, 16'd43953, 16'd28257, 16'd58000});
	test_expansion(128'h875acffc391bc43bd4b4820896d558fb, {16'd11858, 16'd60568, 16'd12034, 16'd25558, 16'd48271, 16'd20434, 16'd11445, 16'd63945, 16'd62006, 16'd34183, 16'd56301, 16'd26840, 16'd63129, 16'd19676, 16'd18662, 16'd44280, 16'd53725, 16'd1559, 16'd39853, 16'd27354, 16'd4242, 16'd20420, 16'd24297, 16'd38105, 16'd21637, 16'd43039});
	test_expansion(128'h7e44cb132fbb44ee2e08500f55eed2f5, {16'd22820, 16'd6350, 16'd35496, 16'd20491, 16'd54591, 16'd33825, 16'd21677, 16'd15520, 16'd11441, 16'd62826, 16'd34163, 16'd61559, 16'd44311, 16'd11463, 16'd38424, 16'd7746, 16'd33908, 16'd3515, 16'd34492, 16'd21329, 16'd65409, 16'd53736, 16'd40313, 16'd46823, 16'd9146, 16'd60173});
	test_expansion(128'hb235e80e1f986e1ef05de131fba23080, {16'd26362, 16'd55454, 16'd55088, 16'd29258, 16'd19265, 16'd737, 16'd30864, 16'd22459, 16'd53461, 16'd62344, 16'd29286, 16'd1653, 16'd19236, 16'd46976, 16'd53571, 16'd486, 16'd55192, 16'd41366, 16'd12335, 16'd58247, 16'd58427, 16'd54857, 16'd64204, 16'd28943, 16'd64673, 16'd43497});
	test_expansion(128'h92c32b5a269d45c5ad5016af413c9cae, {16'd57590, 16'd47281, 16'd64139, 16'd57264, 16'd25243, 16'd9022, 16'd63720, 16'd51226, 16'd58242, 16'd19525, 16'd10660, 16'd59617, 16'd13652, 16'd56022, 16'd8625, 16'd45526, 16'd47332, 16'd54782, 16'd19827, 16'd23236, 16'd57293, 16'd61127, 16'd47873, 16'd46831, 16'd41517, 16'd16395});
	test_expansion(128'hb0cd6d091cc4242a83be147f6869ac58, {16'd29022, 16'd52889, 16'd6478, 16'd11958, 16'd39954, 16'd11102, 16'd32545, 16'd24144, 16'd50289, 16'd20820, 16'd2826, 16'd17062, 16'd46238, 16'd36595, 16'd27532, 16'd38323, 16'd60608, 16'd61215, 16'd27802, 16'd41931, 16'd52224, 16'd40326, 16'd39632, 16'd62328, 16'd7220, 16'd26911});
	test_expansion(128'h5cde377b968bb197f638ce8efff803e0, {16'd27552, 16'd55394, 16'd22908, 16'd43760, 16'd59205, 16'd44129, 16'd60687, 16'd32370, 16'd48032, 16'd58436, 16'd58647, 16'd7927, 16'd42431, 16'd9863, 16'd61245, 16'd58247, 16'd48200, 16'd65093, 16'd33941, 16'd11867, 16'd18498, 16'd47164, 16'd49406, 16'd54416, 16'd56699, 16'd50711});
	test_expansion(128'h8362cbda995b269648cc567d83e394ac, {16'd28930, 16'd31329, 16'd41257, 16'd2386, 16'd30866, 16'd25757, 16'd42570, 16'd40692, 16'd41420, 16'd4639, 16'd42440, 16'd62504, 16'd4346, 16'd46846, 16'd33957, 16'd54685, 16'd28851, 16'd34968, 16'd2438, 16'd60922, 16'd30267, 16'd41864, 16'd45210, 16'd2778, 16'd29519, 16'd38916});
	test_expansion(128'h7ed95de84d2677428ec0adeb0acca472, {16'd25356, 16'd44771, 16'd23439, 16'd12661, 16'd35075, 16'd61920, 16'd17484, 16'd38420, 16'd48203, 16'd5082, 16'd8827, 16'd3758, 16'd24643, 16'd63477, 16'd13255, 16'd54469, 16'd52368, 16'd34072, 16'd4429, 16'd30603, 16'd39151, 16'd27979, 16'd21766, 16'd42534, 16'd41184, 16'd18553});
	test_expansion(128'h14b3797a07412c705e8099102bafcfe8, {16'd54324, 16'd58669, 16'd34236, 16'd1508, 16'd25560, 16'd64141, 16'd63095, 16'd59138, 16'd20986, 16'd32847, 16'd60505, 16'd40204, 16'd11251, 16'd58989, 16'd16547, 16'd4757, 16'd19006, 16'd63743, 16'd7600, 16'd8336, 16'd7488, 16'd46995, 16'd14688, 16'd64895, 16'd17136, 16'd22417});
	test_expansion(128'ha16943fa8ddaf6d555af992c5ba95384, {16'd25940, 16'd4578, 16'd48616, 16'd14817, 16'd39550, 16'd61805, 16'd30137, 16'd15184, 16'd23865, 16'd20992, 16'd21245, 16'd41964, 16'd452, 16'd60240, 16'd30899, 16'd8378, 16'd14103, 16'd7151, 16'd47817, 16'd33899, 16'd14869, 16'd56214, 16'd27660, 16'd22582, 16'd10026, 16'd1497});
	test_expansion(128'h2fd853549833e59e7e59c865c31cc71a, {16'd56813, 16'd54878, 16'd24632, 16'd13070, 16'd21393, 16'd44058, 16'd3348, 16'd10294, 16'd17142, 16'd64600, 16'd46311, 16'd19212, 16'd48917, 16'd21647, 16'd15804, 16'd57623, 16'd31132, 16'd47944, 16'd5113, 16'd9146, 16'd30026, 16'd1456, 16'd16463, 16'd59730, 16'd35767, 16'd4934});
	test_expansion(128'h58c678f2edebb66a01642a7ec24bf8d6, {16'd12391, 16'd59688, 16'd38123, 16'd33249, 16'd61572, 16'd27040, 16'd44696, 16'd55717, 16'd31463, 16'd25931, 16'd10307, 16'd45725, 16'd64505, 16'd59884, 16'd15543, 16'd2808, 16'd16176, 16'd35080, 16'd61677, 16'd32593, 16'd12306, 16'd41252, 16'd30195, 16'd8321, 16'd15850, 16'd56062});
	test_expansion(128'h703b65c62989fbfec9da9b4622b82339, {16'd41821, 16'd52479, 16'd33800, 16'd32073, 16'd26173, 16'd9908, 16'd17946, 16'd61584, 16'd25788, 16'd40889, 16'd21422, 16'd30784, 16'd59690, 16'd46149, 16'd63937, 16'd23804, 16'd8209, 16'd7754, 16'd13137, 16'd64144, 16'd44522, 16'd47287, 16'd11654, 16'd63219, 16'd62265, 16'd22481});
	test_expansion(128'h1bed481e677559181bec49c5d8a3b65e, {16'd59863, 16'd5724, 16'd53071, 16'd63485, 16'd76, 16'd23170, 16'd49605, 16'd39739, 16'd56797, 16'd62431, 16'd49267, 16'd45209, 16'd16279, 16'd21918, 16'd51893, 16'd57663, 16'd17933, 16'd55571, 16'd50731, 16'd3647, 16'd47087, 16'd45497, 16'd40307, 16'd53697, 16'd3953, 16'd14098});
	test_expansion(128'h2182d7ada6ef43b173acbdbf69e54815, {16'd57275, 16'd25216, 16'd4563, 16'd28908, 16'd48979, 16'd29882, 16'd51696, 16'd14617, 16'd43196, 16'd50572, 16'd59350, 16'd23040, 16'd33025, 16'd23815, 16'd33749, 16'd38914, 16'd47683, 16'd29069, 16'd33024, 16'd59887, 16'd33642, 16'd48143, 16'd43073, 16'd37487, 16'd1648, 16'd7416});
	test_expansion(128'he1d2a1ca911a8ba02bd9ae9bf3979e9e, {16'd56362, 16'd44728, 16'd27658, 16'd11479, 16'd20186, 16'd15088, 16'd23153, 16'd16541, 16'd27553, 16'd6708, 16'd53284, 16'd39445, 16'd31175, 16'd56608, 16'd31105, 16'd60930, 16'd48005, 16'd29281, 16'd15127, 16'd46755, 16'd6232, 16'd9403, 16'd58837, 16'd1775, 16'd13261, 16'd25054});
	test_expansion(128'h94c785473d2c60f10e0260573fee7f1b, {16'd34885, 16'd61427, 16'd30958, 16'd57591, 16'd25038, 16'd6443, 16'd57991, 16'd10409, 16'd43133, 16'd1384, 16'd36292, 16'd63628, 16'd819, 16'd50024, 16'd40142, 16'd60932, 16'd30251, 16'd8736, 16'd59812, 16'd3969, 16'd36563, 16'd49766, 16'd11912, 16'd27049, 16'd27932, 16'd7957});
	test_expansion(128'hf614c5be68ce4c82369628f0bf962e69, {16'd33041, 16'd2441, 16'd38632, 16'd44034, 16'd31520, 16'd55956, 16'd37285, 16'd50224, 16'd40948, 16'd37554, 16'd14869, 16'd42931, 16'd58490, 16'd25753, 16'd20896, 16'd6229, 16'd2700, 16'd30729, 16'd4357, 16'd38545, 16'd34876, 16'd61082, 16'd37954, 16'd37544, 16'd47333, 16'd25919});
	test_expansion(128'h207017d7359b7cca40ac12e627f8b8cf, {16'd60411, 16'd45962, 16'd50663, 16'd62615, 16'd55027, 16'd29480, 16'd16323, 16'd12716, 16'd27846, 16'd58606, 16'd25342, 16'd16213, 16'd53354, 16'd50858, 16'd1468, 16'd9079, 16'd8042, 16'd41332, 16'd18700, 16'd33334, 16'd36422, 16'd56265, 16'd45016, 16'd46305, 16'd18155, 16'd25106});
	test_expansion(128'hc6334aec0ec67349f4781d7ba916c049, {16'd31311, 16'd3642, 16'd20806, 16'd30289, 16'd7496, 16'd47367, 16'd16951, 16'd38337, 16'd34893, 16'd63998, 16'd40606, 16'd32385, 16'd20322, 16'd27773, 16'd14534, 16'd4192, 16'd52163, 16'd35578, 16'd51706, 16'd18202, 16'd8714, 16'd16341, 16'd53626, 16'd50720, 16'd17763, 16'd14845});
	test_expansion(128'h2c9655821ef1566a5af232a2b6b332be, {16'd38970, 16'd24221, 16'd19453, 16'd43473, 16'd3804, 16'd2285, 16'd65272, 16'd42177, 16'd22898, 16'd49098, 16'd37799, 16'd22156, 16'd41352, 16'd21968, 16'd6635, 16'd21212, 16'd34311, 16'd13832, 16'd52285, 16'd48332, 16'd62133, 16'd39310, 16'd35250, 16'd11617, 16'd53000, 16'd8053});
	test_expansion(128'h7e6a7ecd1ca5ed0f588b73d2a3ef7a22, {16'd54287, 16'd16307, 16'd13425, 16'd64609, 16'd62244, 16'd10862, 16'd31893, 16'd18582, 16'd8159, 16'd23793, 16'd38837, 16'd52083, 16'd42473, 16'd57961, 16'd63762, 16'd4079, 16'd2954, 16'd4439, 16'd47087, 16'd6569, 16'd52165, 16'd50334, 16'd7101, 16'd11159, 16'd27032, 16'd2294});
	test_expansion(128'ha8d28f81fc54d153e396efb009ddbe6f, {16'd55645, 16'd37649, 16'd65234, 16'd50366, 16'd42174, 16'd14922, 16'd32160, 16'd12670, 16'd52587, 16'd37182, 16'd7797, 16'd41840, 16'd11540, 16'd61603, 16'd60633, 16'd40596, 16'd33628, 16'd28587, 16'd5286, 16'd10210, 16'd37618, 16'd19823, 16'd880, 16'd56909, 16'd58485, 16'd40193});
	test_expansion(128'he25063b9ac6d2c452a1ffb967143962c, {16'd4283, 16'd49502, 16'd21865, 16'd20924, 16'd9304, 16'd55463, 16'd17169, 16'd21986, 16'd25746, 16'd48595, 16'd1374, 16'd14511, 16'd15233, 16'd51308, 16'd5505, 16'd63177, 16'd38670, 16'd10720, 16'd25009, 16'd29704, 16'd43457, 16'd8333, 16'd11979, 16'd49769, 16'd28480, 16'd27648});
	test_expansion(128'h6d7a5257c0ffc90d29f9d2ba38d0fa76, {16'd50150, 16'd56874, 16'd42710, 16'd49462, 16'd3730, 16'd43729, 16'd20555, 16'd46265, 16'd20761, 16'd3487, 16'd28482, 16'd28070, 16'd27006, 16'd3759, 16'd65371, 16'd47090, 16'd61113, 16'd54813, 16'd22533, 16'd22568, 16'd38775, 16'd35951, 16'd2335, 16'd64512, 16'd54429, 16'd38919});
	test_expansion(128'h915be67303fb0e2bf4d429c12aa8e0b8, {16'd26226, 16'd32583, 16'd17164, 16'd26645, 16'd45976, 16'd45150, 16'd9929, 16'd62461, 16'd30028, 16'd22558, 16'd18475, 16'd56298, 16'd11013, 16'd8525, 16'd64829, 16'd25733, 16'd56311, 16'd14661, 16'd9519, 16'd51391, 16'd3385, 16'd57237, 16'd45727, 16'd10196, 16'd48326, 16'd395});
	test_expansion(128'hcd01ba4f189bf06acfbf59f176040a56, {16'd22518, 16'd15777, 16'd49566, 16'd48923, 16'd21711, 16'd4673, 16'd27413, 16'd17228, 16'd34985, 16'd56267, 16'd57211, 16'd29124, 16'd20134, 16'd26175, 16'd10153, 16'd62768, 16'd29253, 16'd18246, 16'd57823, 16'd14416, 16'd3945, 16'd28855, 16'd53836, 16'd22237, 16'd7115, 16'd6152});
	test_expansion(128'h6de0bc805da29af85fcc9802a2960f97, {16'd55299, 16'd23975, 16'd62694, 16'd11073, 16'd42246, 16'd27893, 16'd64284, 16'd25743, 16'd48511, 16'd30616, 16'd46255, 16'd50854, 16'd48221, 16'd61142, 16'd63877, 16'd63683, 16'd61914, 16'd8417, 16'd61680, 16'd5502, 16'd15470, 16'd1058, 16'd46414, 16'd23991, 16'd61992, 16'd28074});
	test_expansion(128'hb49cead442930c1456044ffcbad5046a, {16'd60831, 16'd32739, 16'd62988, 16'd47812, 16'd7907, 16'd8538, 16'd53191, 16'd9725, 16'd45415, 16'd32828, 16'd41453, 16'd26587, 16'd38836, 16'd17791, 16'd47682, 16'd14162, 16'd42207, 16'd2573, 16'd54126, 16'd39067, 16'd1188, 16'd37313, 16'd41545, 16'd61393, 16'd46089, 16'd57035});
	test_expansion(128'he65891cf440c8a0962fe73d13fc0f7bf, {16'd63444, 16'd54879, 16'd42746, 16'd3697, 16'd55640, 16'd62625, 16'd46224, 16'd64832, 16'd10858, 16'd16128, 16'd61985, 16'd24866, 16'd50747, 16'd23894, 16'd18383, 16'd37172, 16'd6539, 16'd36184, 16'd9384, 16'd55082, 16'd34451, 16'd18140, 16'd27345, 16'd44377, 16'd27889, 16'd55231});
	test_expansion(128'h982a04213f37f82368a69717a4258a03, {16'd19572, 16'd35631, 16'd51697, 16'd40591, 16'd41707, 16'd51681, 16'd47401, 16'd31902, 16'd26290, 16'd30324, 16'd35850, 16'd8751, 16'd65236, 16'd57254, 16'd60157, 16'd9990, 16'd52556, 16'd14914, 16'd40410, 16'd48766, 16'd55018, 16'd50847, 16'd58160, 16'd25438, 16'd29898, 16'd37501});
	test_expansion(128'h7601fff0b04bd4affe77e70b3c0a0563, {16'd58961, 16'd5783, 16'd18726, 16'd59683, 16'd25196, 16'd35923, 16'd9399, 16'd21378, 16'd20432, 16'd4657, 16'd36693, 16'd46952, 16'd3939, 16'd47647, 16'd55389, 16'd33730, 16'd3610, 16'd39388, 16'd64758, 16'd20230, 16'd29337, 16'd35304, 16'd37474, 16'd46993, 16'd42305, 16'd54264});
	test_expansion(128'h4a1823ac39696d55cdc9a28b0445c52a, {16'd57663, 16'd12841, 16'd36363, 16'd52490, 16'd40792, 16'd55852, 16'd19105, 16'd40938, 16'd56983, 16'd40921, 16'd63631, 16'd41726, 16'd42626, 16'd52624, 16'd35418, 16'd4008, 16'd48275, 16'd45327, 16'd26075, 16'd17980, 16'd32241, 16'd3801, 16'd26128, 16'd6031, 16'd25909, 16'd27783});
	test_expansion(128'h1801c89f27f1bdba21cbbe02c854a218, {16'd65095, 16'd62568, 16'd16385, 16'd51091, 16'd3039, 16'd46196, 16'd40304, 16'd2823, 16'd1295, 16'd43992, 16'd60399, 16'd63246, 16'd57841, 16'd28047, 16'd43416, 16'd25790, 16'd31811, 16'd7138, 16'd58665, 16'd53117, 16'd10922, 16'd38129, 16'd41656, 16'd45712, 16'd53502, 16'd26120});
	test_expansion(128'h90ff2e7a6e8d8e2cefada7e502dd7ab8, {16'd3583, 16'd41920, 16'd36723, 16'd23841, 16'd42408, 16'd63842, 16'd35166, 16'd13748, 16'd24821, 16'd21359, 16'd43405, 16'd17502, 16'd29037, 16'd38600, 16'd60010, 16'd54069, 16'd20685, 16'd11415, 16'd3767, 16'd14868, 16'd33790, 16'd6834, 16'd39893, 16'd58135, 16'd64813, 16'd35178});
	test_expansion(128'ha931fd4a08b620773016fd2f1808b139, {16'd52357, 16'd36950, 16'd41922, 16'd5463, 16'd3391, 16'd28448, 16'd4947, 16'd58393, 16'd11271, 16'd42348, 16'd25799, 16'd22582, 16'd56755, 16'd49231, 16'd28038, 16'd53963, 16'd17251, 16'd45888, 16'd6642, 16'd27907, 16'd64317, 16'd45153, 16'd43488, 16'd31873, 16'd33180, 16'd37584});
	test_expansion(128'hee9be39d83dc0da99bf530fe5b2a2682, {16'd53363, 16'd50413, 16'd20852, 16'd63483, 16'd39783, 16'd5426, 16'd51693, 16'd15994, 16'd17456, 16'd14978, 16'd2390, 16'd8018, 16'd767, 16'd39492, 16'd46472, 16'd26296, 16'd2318, 16'd35629, 16'd63021, 16'd62570, 16'd14270, 16'd2799, 16'd63142, 16'd38660, 16'd60893, 16'd46708});
	test_expansion(128'hf3df7625804c15fc0633450d5078d31a, {16'd760, 16'd40218, 16'd58761, 16'd34617, 16'd48015, 16'd28062, 16'd20182, 16'd18468, 16'd17447, 16'd39302, 16'd46132, 16'd45043, 16'd45508, 16'd52754, 16'd42507, 16'd51941, 16'd47279, 16'd56725, 16'd7770, 16'd4703, 16'd31850, 16'd57468, 16'd45775, 16'd7086, 16'd12109, 16'd50824});
	test_expansion(128'h7c9ef976cf886041cdb4d5b46280ee13, {16'd52332, 16'd62525, 16'd777, 16'd56329, 16'd8388, 16'd29302, 16'd16903, 16'd11289, 16'd25849, 16'd1849, 16'd64471, 16'd43961, 16'd28865, 16'd16888, 16'd58166, 16'd61581, 16'd61635, 16'd46932, 16'd2089, 16'd61971, 16'd43524, 16'd3416, 16'd50269, 16'd33487, 16'd34140, 16'd59321});
	test_expansion(128'h81f9511434890c70e6d6ec1eaca19f6a, {16'd22462, 16'd7931, 16'd2409, 16'd48944, 16'd29205, 16'd25180, 16'd57055, 16'd63500, 16'd50210, 16'd44003, 16'd40106, 16'd55318, 16'd51494, 16'd28372, 16'd60355, 16'd37610, 16'd3715, 16'd30559, 16'd6209, 16'd58404, 16'd65436, 16'd20340, 16'd41246, 16'd63460, 16'd33469, 16'd29826});
	test_expansion(128'h6c3e6fa2a91050a74b1c31c4bb5a23c7, {16'd36523, 16'd56267, 16'd26275, 16'd34426, 16'd6200, 16'd39400, 16'd53554, 16'd61570, 16'd37446, 16'd63455, 16'd60232, 16'd6611, 16'd9572, 16'd14136, 16'd3143, 16'd7954, 16'd37117, 16'd49380, 16'd64792, 16'd56555, 16'd783, 16'd25060, 16'd38034, 16'd42194, 16'd19390, 16'd30243});
	test_expansion(128'h5fd51604c309509d61144887a23718b6, {16'd36987, 16'd7998, 16'd20688, 16'd40463, 16'd53422, 16'd28841, 16'd32157, 16'd22155, 16'd9438, 16'd46696, 16'd48370, 16'd22905, 16'd60437, 16'd54155, 16'd40843, 16'd63814, 16'd50434, 16'd5404, 16'd44244, 16'd1566, 16'd64321, 16'd58931, 16'd50718, 16'd64933, 16'd30908, 16'd41385});
	test_expansion(128'hc15394400cffa074026d129e9c75b4fa, {16'd10596, 16'd54793, 16'd45729, 16'd46447, 16'd17697, 16'd29732, 16'd21875, 16'd24938, 16'd42857, 16'd43975, 16'd9287, 16'd4352, 16'd22377, 16'd62037, 16'd64637, 16'd53431, 16'd27723, 16'd3964, 16'd49431, 16'd28668, 16'd23660, 16'd22609, 16'd15504, 16'd29147, 16'd4015, 16'd54366});
	test_expansion(128'h01d1d4d4ebfdf6a5a3e0be171802cda8, {16'd25227, 16'd43875, 16'd56563, 16'd29764, 16'd8381, 16'd7670, 16'd38934, 16'd43298, 16'd28916, 16'd50006, 16'd62831, 16'd45234, 16'd26836, 16'd40401, 16'd58684, 16'd61072, 16'd38835, 16'd41350, 16'd64799, 16'd44752, 16'd19023, 16'd40330, 16'd2724, 16'd27435, 16'd27784, 16'd22340});
	test_expansion(128'h805d4014355196acf65b2190f0e7caac, {16'd28319, 16'd6608, 16'd3478, 16'd3080, 16'd32771, 16'd31178, 16'd47863, 16'd28546, 16'd59484, 16'd47974, 16'd50842, 16'd4107, 16'd41501, 16'd42838, 16'd48869, 16'd39141, 16'd50635, 16'd45098, 16'd8508, 16'd21919, 16'd18993, 16'd26680, 16'd23917, 16'd2241, 16'd50327, 16'd19490});
	test_expansion(128'hd1b2d99e3f98f548b31eaf6b59ed9b7e, {16'd4356, 16'd14, 16'd20717, 16'd23913, 16'd30516, 16'd41114, 16'd64843, 16'd23202, 16'd178, 16'd41329, 16'd26585, 16'd9466, 16'd17587, 16'd62597, 16'd29755, 16'd15250, 16'd50846, 16'd38806, 16'd26359, 16'd54383, 16'd55420, 16'd39862, 16'd39582, 16'd63116, 16'd8938, 16'd5866});
	test_expansion(128'h2765b1524659d78fd8b0b0dda26c82c9, {16'd30390, 16'd49449, 16'd8214, 16'd48731, 16'd19308, 16'd8993, 16'd60847, 16'd11258, 16'd40787, 16'd5505, 16'd24649, 16'd2080, 16'd51704, 16'd30882, 16'd32103, 16'd28386, 16'd43717, 16'd25815, 16'd45238, 16'd17100, 16'd56559, 16'd33240, 16'd19653, 16'd22796, 16'd60415, 16'd55358});
	test_expansion(128'h69173b5884ea356c6c1a4fc7758b1612, {16'd9634, 16'd48916, 16'd45115, 16'd45455, 16'd63823, 16'd30108, 16'd30177, 16'd62668, 16'd51470, 16'd43578, 16'd33960, 16'd25564, 16'd48086, 16'd29512, 16'd22531, 16'd41049, 16'd28815, 16'd65081, 16'd40592, 16'd7694, 16'd37661, 16'd25183, 16'd65507, 16'd35436, 16'd21669, 16'd14030});
	test_expansion(128'h4546544c6f1c04f7ab9d7a690b713222, {16'd42286, 16'd32652, 16'd64098, 16'd34944, 16'd4557, 16'd10228, 16'd18723, 16'd22835, 16'd34750, 16'd7029, 16'd14249, 16'd34095, 16'd8443, 16'd10367, 16'd12608, 16'd31577, 16'd63379, 16'd34634, 16'd55246, 16'd19348, 16'd28723, 16'd49479, 16'd47387, 16'd8775, 16'd53923, 16'd17916});
	test_expansion(128'h798161f6935ffbb3041f12695d8ea2ac, {16'd58522, 16'd14003, 16'd3011, 16'd24321, 16'd18693, 16'd47236, 16'd20528, 16'd60537, 16'd15534, 16'd28079, 16'd26043, 16'd29505, 16'd27419, 16'd7029, 16'd41937, 16'd21804, 16'd34717, 16'd47308, 16'd25536, 16'd933, 16'd50711, 16'd25152, 16'd34258, 16'd3072, 16'd32529, 16'd7842});
	test_expansion(128'h4c7e87491ec4da2aad2a7388ea0f1ed8, {16'd15596, 16'd39932, 16'd52939, 16'd58318, 16'd3002, 16'd6106, 16'd15367, 16'd52726, 16'd36354, 16'd58328, 16'd16502, 16'd16637, 16'd13108, 16'd49556, 16'd20577, 16'd12241, 16'd42259, 16'd14201, 16'd51377, 16'd33746, 16'd38646, 16'd34914, 16'd8461, 16'd52877, 16'd21882, 16'd61435});
	test_expansion(128'hd8dc9b616e8947e99f98e5da7cae155c, {16'd12339, 16'd31125, 16'd14049, 16'd32727, 16'd64922, 16'd1793, 16'd64457, 16'd17658, 16'd21819, 16'd28748, 16'd54145, 16'd12239, 16'd14138, 16'd63335, 16'd58215, 16'd32932, 16'd53528, 16'd27556, 16'd37828, 16'd8670, 16'd29465, 16'd46795, 16'd14591, 16'd60024, 16'd41979, 16'd6313});
	test_expansion(128'h5fa31a819d4822aac1e8d6f6d1eaaeff, {16'd19049, 16'd54790, 16'd48297, 16'd31628, 16'd13370, 16'd37704, 16'd22782, 16'd29105, 16'd26972, 16'd39839, 16'd29773, 16'd23756, 16'd47392, 16'd20084, 16'd19934, 16'd28351, 16'd59930, 16'd5718, 16'd37303, 16'd46023, 16'd27190, 16'd29063, 16'd41881, 16'd14583, 16'd16979, 16'd62515});
	test_expansion(128'h74c89288f9382116894ed1d621dd4fa6, {16'd49600, 16'd32622, 16'd64233, 16'd56915, 16'd58425, 16'd33842, 16'd4022, 16'd6757, 16'd59266, 16'd45622, 16'd8267, 16'd31700, 16'd20246, 16'd30050, 16'd65215, 16'd46837, 16'd32089, 16'd26442, 16'd34982, 16'd41946, 16'd15022, 16'd31736, 16'd3173, 16'd64297, 16'd11809, 16'd9535});
	test_expansion(128'h30e3f5bfd68513e692a091e9c59dc324, {16'd38083, 16'd40365, 16'd4330, 16'd58921, 16'd63626, 16'd33153, 16'd58564, 16'd46324, 16'd20496, 16'd53064, 16'd13095, 16'd11, 16'd41712, 16'd64534, 16'd59459, 16'd15548, 16'd13635, 16'd43751, 16'd15050, 16'd43171, 16'd31672, 16'd20861, 16'd33795, 16'd55149, 16'd25039, 16'd21187});
	test_expansion(128'h45fee9dfd7318680d0d52d716fddabe3, {16'd8760, 16'd53477, 16'd15948, 16'd2431, 16'd46115, 16'd10274, 16'd7577, 16'd5272, 16'd64657, 16'd13702, 16'd30330, 16'd2812, 16'd49623, 16'd40871, 16'd48857, 16'd56201, 16'd31835, 16'd45210, 16'd27993, 16'd47593, 16'd58607, 16'd40018, 16'd14132, 16'd32672, 16'd52690, 16'd22753});
	test_expansion(128'hfba94af0276c6d6cbb7e73273a2063d6, {16'd10335, 16'd9949, 16'd43132, 16'd49414, 16'd47530, 16'd24060, 16'd35646, 16'd2512, 16'd58476, 16'd5773, 16'd11403, 16'd3882, 16'd7545, 16'd59770, 16'd1796, 16'd52390, 16'd22871, 16'd59271, 16'd18640, 16'd6368, 16'd48843, 16'd21312, 16'd5389, 16'd7161, 16'd19913, 16'd23717});
	test_expansion(128'he25589e984041b8d70dcbc0e485eb78e, {16'd58199, 16'd1215, 16'd46951, 16'd53981, 16'd31822, 16'd63627, 16'd36648, 16'd34211, 16'd10788, 16'd48727, 16'd212, 16'd8169, 16'd17192, 16'd63149, 16'd55255, 16'd38879, 16'd63965, 16'd58912, 16'd27468, 16'd32300, 16'd37820, 16'd22594, 16'd41242, 16'd16652, 16'd19250, 16'd23961});
	test_expansion(128'he695378d521bb6d594b677729720a688, {16'd10686, 16'd53501, 16'd41404, 16'd20115, 16'd16782, 16'd45953, 16'd4782, 16'd13476, 16'd45965, 16'd21304, 16'd62718, 16'd65417, 16'd946, 16'd48644, 16'd13393, 16'd13534, 16'd31209, 16'd34017, 16'd52673, 16'd22990, 16'd4868, 16'd35052, 16'd37871, 16'd3879, 16'd12304, 16'd51246});
	test_expansion(128'h0f21bd79dcccf6a1e76e0b97e13f2e26, {16'd48250, 16'd44109, 16'd3629, 16'd63397, 16'd47286, 16'd23852, 16'd54668, 16'd23668, 16'd17231, 16'd39599, 16'd41309, 16'd41188, 16'd29974, 16'd37202, 16'd34272, 16'd60269, 16'd57909, 16'd15438, 16'd56051, 16'd49371, 16'd14343, 16'd23651, 16'd51117, 16'd15951, 16'd4705, 16'd10424});
	test_expansion(128'h2057f189ba79a22d127af26dbd2f349d, {16'd57031, 16'd24428, 16'd31398, 16'd33636, 16'd27645, 16'd1855, 16'd43929, 16'd51430, 16'd12896, 16'd31494, 16'd50468, 16'd57879, 16'd5246, 16'd37494, 16'd14747, 16'd62197, 16'd27695, 16'd32284, 16'd51531, 16'd11185, 16'd4371, 16'd5505, 16'd41566, 16'd41841, 16'd64175, 16'd42999});
	test_expansion(128'hce8859fb1d4273db42ce948f6d598f2e, {16'd61807, 16'd45383, 16'd48414, 16'd220, 16'd50871, 16'd22563, 16'd45095, 16'd34389, 16'd65196, 16'd15367, 16'd36518, 16'd27438, 16'd63090, 16'd34726, 16'd27049, 16'd63405, 16'd61083, 16'd60829, 16'd22373, 16'd16171, 16'd34295, 16'd56997, 16'd63963, 16'd27498, 16'd38168, 16'd28927});
	test_expansion(128'h8228c1f93348bc251874927117476050, {16'd15718, 16'd3031, 16'd42710, 16'd27042, 16'd41901, 16'd18423, 16'd49760, 16'd48651, 16'd56768, 16'd9920, 16'd48132, 16'd46269, 16'd1653, 16'd54336, 16'd11841, 16'd47991, 16'd23805, 16'd210, 16'd30271, 16'd52991, 16'd28922, 16'd575, 16'd55205, 16'd56173, 16'd7188, 16'd1043});
	test_expansion(128'h32075e317c58587c384bcb0d0bc8e25e, {16'd61538, 16'd34124, 16'd6117, 16'd4842, 16'd24853, 16'd59598, 16'd21430, 16'd17276, 16'd30649, 16'd56403, 16'd3453, 16'd41875, 16'd31051, 16'd20971, 16'd42669, 16'd13288, 16'd27521, 16'd54841, 16'd40516, 16'd13489, 16'd23515, 16'd56792, 16'd14904, 16'd4167, 16'd762, 16'd7011});
	test_expansion(128'h3d0ab81724d53e1c333be1d58b616070, {16'd55972, 16'd47328, 16'd9551, 16'd45609, 16'd22437, 16'd64555, 16'd13439, 16'd36875, 16'd26452, 16'd1641, 16'd39019, 16'd37239, 16'd51451, 16'd44147, 16'd58089, 16'd20916, 16'd44841, 16'd6854, 16'd24773, 16'd59109, 16'd46685, 16'd4114, 16'd62327, 16'd3229, 16'd55477, 16'd38533});
	test_expansion(128'hcbb32506b68ceaeade42491af1a63d38, {16'd40043, 16'd30980, 16'd17353, 16'd21103, 16'd23950, 16'd28771, 16'd48639, 16'd56963, 16'd9517, 16'd42451, 16'd23629, 16'd61632, 16'd11012, 16'd43723, 16'd25167, 16'd8196, 16'd27121, 16'd14765, 16'd40338, 16'd42552, 16'd37732, 16'd14911, 16'd61224, 16'd40844, 16'd50624, 16'd27200});
	test_expansion(128'h7dcc6059cc1070114fb11e261a1d11a3, {16'd31626, 16'd12222, 16'd50255, 16'd30880, 16'd18968, 16'd36275, 16'd47441, 16'd22485, 16'd48494, 16'd24931, 16'd58739, 16'd41759, 16'd55240, 16'd52454, 16'd44759, 16'd62396, 16'd28144, 16'd42635, 16'd19991, 16'd52962, 16'd30895, 16'd28033, 16'd61504, 16'd10192, 16'd46219, 16'd43568});
	test_expansion(128'h186560224bc9c83e4818a0d2136a4026, {16'd43927, 16'd55457, 16'd64243, 16'd35940, 16'd36072, 16'd24502, 16'd2970, 16'd14831, 16'd48415, 16'd55849, 16'd3992, 16'd37522, 16'd16072, 16'd52047, 16'd60065, 16'd19989, 16'd53786, 16'd6848, 16'd34680, 16'd20252, 16'd12666, 16'd44897, 16'd24878, 16'd45819, 16'd34721, 16'd7677});
	test_expansion(128'h3b626098d547aaf286f820c6a4d776cd, {16'd53351, 16'd57521, 16'd9258, 16'd60452, 16'd1975, 16'd14564, 16'd35011, 16'd17286, 16'd47067, 16'd24899, 16'd28225, 16'd16272, 16'd61356, 16'd14164, 16'd63789, 16'd24129, 16'd26114, 16'd65154, 16'd20329, 16'd1606, 16'd13084, 16'd64676, 16'd894, 16'd11528, 16'd23698, 16'd61825});
	test_expansion(128'hfedb5e17cdaa8b5e4230bcd73999f246, {16'd30181, 16'd13073, 16'd17327, 16'd28346, 16'd39537, 16'd48890, 16'd44780, 16'd61182, 16'd32281, 16'd55381, 16'd11712, 16'd41594, 16'd31328, 16'd25968, 16'd56680, 16'd8198, 16'd20186, 16'd20897, 16'd7700, 16'd12978, 16'd7188, 16'd9076, 16'd40339, 16'd26584, 16'd30556, 16'd7971});
	test_expansion(128'h5871985642b0c60ab4cc2405bbbc94d0, {16'd8139, 16'd61585, 16'd46901, 16'd37399, 16'd33594, 16'd52853, 16'd62169, 16'd40931, 16'd52185, 16'd36977, 16'd21875, 16'd27302, 16'd782, 16'd58116, 16'd57193, 16'd39237, 16'd57873, 16'd1004, 16'd32615, 16'd32588, 16'd31114, 16'd2154, 16'd62088, 16'd59882, 16'd34977, 16'd63635});
	test_expansion(128'hb17707a3d93f290f6ed5ff9fcf6f03c0, {16'd4036, 16'd8908, 16'd14498, 16'd19928, 16'd56691, 16'd5704, 16'd32123, 16'd14824, 16'd15262, 16'd24731, 16'd17237, 16'd53907, 16'd39532, 16'd39720, 16'd19886, 16'd55944, 16'd28804, 16'd42503, 16'd9229, 16'd62252, 16'd26488, 16'd47276, 16'd27447, 16'd53790, 16'd48470, 16'd27295});
	test_expansion(128'h4f6377ab24969164a668d301bae29f93, {16'd39869, 16'd60159, 16'd62873, 16'd51260, 16'd4033, 16'd54940, 16'd18121, 16'd35384, 16'd4985, 16'd39269, 16'd59138, 16'd37849, 16'd34460, 16'd45042, 16'd9316, 16'd52080, 16'd35566, 16'd63145, 16'd17594, 16'd16269, 16'd43229, 16'd57182, 16'd42374, 16'd42659, 16'd53454, 16'd60236});
	test_expansion(128'h67642829f9628124ee91bd8fe2b98de3, {16'd59642, 16'd62918, 16'd29922, 16'd10159, 16'd32051, 16'd65405, 16'd17426, 16'd14771, 16'd61687, 16'd22736, 16'd16395, 16'd37539, 16'd27455, 16'd41650, 16'd14414, 16'd32107, 16'd5045, 16'd4869, 16'd31158, 16'd8893, 16'd49244, 16'd26278, 16'd62236, 16'd32450, 16'd22611, 16'd44115});
	test_expansion(128'ha9fc3269084a816d707eb31df8f2e540, {16'd16553, 16'd22144, 16'd11275, 16'd20626, 16'd18253, 16'd13557, 16'd18046, 16'd43022, 16'd32960, 16'd28442, 16'd23284, 16'd51950, 16'd31937, 16'd13180, 16'd3430, 16'd59889, 16'd54539, 16'd2026, 16'd1964, 16'd14060, 16'd21969, 16'd57776, 16'd50801, 16'd439, 16'd57123, 16'd12892});
	test_expansion(128'hccda2807b6607818bd1b9b8db87e4334, {16'd25764, 16'd3944, 16'd62865, 16'd21528, 16'd33012, 16'd24363, 16'd16867, 16'd35177, 16'd16688, 16'd21263, 16'd25976, 16'd1031, 16'd49294, 16'd60672, 16'd4879, 16'd11617, 16'd56515, 16'd4289, 16'd28238, 16'd60974, 16'd26730, 16'd16170, 16'd6997, 16'd23694, 16'd10330, 16'd11249});
	test_expansion(128'hc21816244a3ef8471d3b83396502824d, {16'd53980, 16'd80, 16'd59068, 16'd40676, 16'd59427, 16'd32169, 16'd39083, 16'd27913, 16'd40257, 16'd60745, 16'd61665, 16'd8019, 16'd24247, 16'd31904, 16'd39796, 16'd18293, 16'd22823, 16'd951, 16'd3147, 16'd11229, 16'd25839, 16'd48634, 16'd11800, 16'd57540, 16'd52777, 16'd54845});
	test_expansion(128'h44e2f18ec460fce17f37b0482360239c, {16'd52054, 16'd19375, 16'd32782, 16'd42234, 16'd61142, 16'd14714, 16'd9507, 16'd1973, 16'd53182, 16'd27064, 16'd60785, 16'd26863, 16'd54457, 16'd17662, 16'd31763, 16'd61813, 16'd42713, 16'd3751, 16'd16073, 16'd31690, 16'd618, 16'd44730, 16'd491, 16'd58777, 16'd62129, 16'd24495});
	test_expansion(128'h58c084b306ddd58528ecce7c849df798, {16'd37645, 16'd15534, 16'd50021, 16'd48543, 16'd34252, 16'd3800, 16'd11079, 16'd63724, 16'd56162, 16'd18078, 16'd10677, 16'd57237, 16'd60900, 16'd6215, 16'd30733, 16'd19768, 16'd24888, 16'd46198, 16'd24504, 16'd61727, 16'd65034, 16'd47939, 16'd13712, 16'd62600, 16'd55108, 16'd51564});
	test_expansion(128'h4df1294bc972fadefa0098befcf7ce55, {16'd63434, 16'd7599, 16'd52121, 16'd41547, 16'd30481, 16'd17153, 16'd36467, 16'd709, 16'd35821, 16'd34419, 16'd45360, 16'd14663, 16'd1048, 16'd33919, 16'd13995, 16'd63646, 16'd52539, 16'd60699, 16'd334, 16'd60211, 16'd22393, 16'd25313, 16'd52626, 16'd39212, 16'd57526, 16'd62829});
	test_expansion(128'h6404adc64eafd9cdc4c51c7f915aca9e, {16'd9407, 16'd29837, 16'd23423, 16'd27946, 16'd61194, 16'd37218, 16'd42780, 16'd64311, 16'd38605, 16'd47405, 16'd22711, 16'd51578, 16'd48482, 16'd63400, 16'd44165, 16'd26433, 16'd42908, 16'd5599, 16'd46809, 16'd64708, 16'd58134, 16'd53458, 16'd11835, 16'd40970, 16'd14280, 16'd54150});
	test_expansion(128'h8502774395fc8e8cc25d379d3738ba06, {16'd32442, 16'd4868, 16'd63559, 16'd12629, 16'd61890, 16'd61300, 16'd61536, 16'd26997, 16'd3970, 16'd3992, 16'd5467, 16'd37430, 16'd21930, 16'd15126, 16'd15921, 16'd20894, 16'd60568, 16'd34864, 16'd54603, 16'd17075, 16'd22525, 16'd53813, 16'd38638, 16'd36793, 16'd16490, 16'd33623});
	test_expansion(128'h24a69215f3af07b9fffd38fb1b996ae9, {16'd18823, 16'd6104, 16'd45685, 16'd17371, 16'd30654, 16'd3757, 16'd48807, 16'd44617, 16'd2301, 16'd48990, 16'd37671, 16'd434, 16'd60113, 16'd886, 16'd39843, 16'd37517, 16'd52127, 16'd53851, 16'd24778, 16'd2585, 16'd54283, 16'd16196, 16'd3137, 16'd16536, 16'd1414, 16'd64983});
	test_expansion(128'ha54480daea35697db2c6a0ad29e1212d, {16'd48752, 16'd51838, 16'd42977, 16'd21084, 16'd63124, 16'd10622, 16'd29225, 16'd43916, 16'd57459, 16'd11278, 16'd16010, 16'd52499, 16'd27843, 16'd35009, 16'd45660, 16'd21592, 16'd1301, 16'd39274, 16'd32819, 16'd35089, 16'd29689, 16'd35098, 16'd46808, 16'd58586, 16'd58309, 16'd33613});
	test_expansion(128'h443f95227c3d5d29919898e9a8321ca9, {16'd44202, 16'd49991, 16'd42616, 16'd17052, 16'd16014, 16'd28402, 16'd7269, 16'd33153, 16'd48483, 16'd22356, 16'd59590, 16'd34719, 16'd63855, 16'd18118, 16'd40209, 16'd30130, 16'd58267, 16'd52560, 16'd25099, 16'd43188, 16'd30722, 16'd20046, 16'd42253, 16'd20401, 16'd8655, 16'd49418});
	test_expansion(128'h7c2fce852148c4f43937d4f2ef360570, {16'd24277, 16'd39642, 16'd62035, 16'd6791, 16'd39987, 16'd1665, 16'd22061, 16'd18649, 16'd55344, 16'd51934, 16'd1070, 16'd55043, 16'd40211, 16'd32042, 16'd65146, 16'd46465, 16'd59141, 16'd22958, 16'd21288, 16'd8132, 16'd646, 16'd57818, 16'd26258, 16'd22787, 16'd14478, 16'd51556});
	test_expansion(128'h5b1527773552f42cce984d643913faa0, {16'd6438, 16'd60436, 16'd38841, 16'd28636, 16'd55926, 16'd13608, 16'd10284, 16'd28939, 16'd9315, 16'd20696, 16'd16956, 16'd62544, 16'd48146, 16'd9400, 16'd6653, 16'd20515, 16'd27343, 16'd58556, 16'd54659, 16'd22544, 16'd39615, 16'd15675, 16'd24863, 16'd39508, 16'd18559, 16'd4751});
	test_expansion(128'h63c88804ebf68a457bb6bc016b92c865, {16'd29018, 16'd65500, 16'd1700, 16'd29123, 16'd13041, 16'd60741, 16'd11393, 16'd41740, 16'd4708, 16'd57763, 16'd6262, 16'd2512, 16'd9552, 16'd51303, 16'd43258, 16'd42563, 16'd30985, 16'd61418, 16'd2379, 16'd38, 16'd28189, 16'd26593, 16'd32455, 16'd44305, 16'd33223, 16'd63352});
	test_expansion(128'h091e3061951d4b69f86b69496e94ce7a, {16'd36391, 16'd26778, 16'd28923, 16'd46439, 16'd13375, 16'd6266, 16'd62344, 16'd4859, 16'd62069, 16'd48950, 16'd38315, 16'd342, 16'd14388, 16'd41854, 16'd900, 16'd1221, 16'd64412, 16'd28703, 16'd4710, 16'd64789, 16'd21335, 16'd25255, 16'd21669, 16'd44990, 16'd18765, 16'd12161});
	test_expansion(128'hae3c637ef6c944521df3f66b14908d5c, {16'd1144, 16'd40658, 16'd24963, 16'd20949, 16'd24821, 16'd56554, 16'd46068, 16'd29616, 16'd16088, 16'd20162, 16'd32828, 16'd30484, 16'd38786, 16'd13644, 16'd18327, 16'd9940, 16'd37073, 16'd41577, 16'd39594, 16'd1569, 16'd23835, 16'd12430, 16'd376, 16'd25072, 16'd15909, 16'd58785});
	test_expansion(128'h381c121fca50cb6db8a20075b0f0c53f, {16'd36939, 16'd58311, 16'd13816, 16'd58224, 16'd49266, 16'd50026, 16'd22786, 16'd34112, 16'd40198, 16'd59055, 16'd26062, 16'd54385, 16'd41042, 16'd14606, 16'd48406, 16'd11862, 16'd34048, 16'd47232, 16'd60766, 16'd30348, 16'd38219, 16'd15347, 16'd51791, 16'd22813, 16'd25401, 16'd11695});
	test_expansion(128'h56bde33cf6829bd25d7b433c21e72651, {16'd61073, 16'd13579, 16'd2202, 16'd19471, 16'd46704, 16'd13490, 16'd12571, 16'd47889, 16'd51868, 16'd54228, 16'd35827, 16'd24840, 16'd21118, 16'd44299, 16'd26990, 16'd8459, 16'd21223, 16'd60819, 16'd22228, 16'd15203, 16'd13762, 16'd33945, 16'd8895, 16'd64480, 16'd41282, 16'd43395});
	test_expansion(128'h1a0e9a9aef3850e07b66ca58a7b54928, {16'd57107, 16'd56977, 16'd54382, 16'd3710, 16'd55510, 16'd8998, 16'd45402, 16'd35347, 16'd20972, 16'd20172, 16'd10882, 16'd56606, 16'd25313, 16'd11794, 16'd53824, 16'd60135, 16'd39898, 16'd18080, 16'd361, 16'd48535, 16'd63795, 16'd28524, 16'd38053, 16'd8324, 16'd892, 16'd49230});
	test_expansion(128'h17e3c27bfb653a2134b623d2a99c1708, {16'd44767, 16'd28504, 16'd4090, 16'd49054, 16'd51127, 16'd25908, 16'd20378, 16'd48910, 16'd1280, 16'd19125, 16'd11233, 16'd17883, 16'd30017, 16'd17171, 16'd38721, 16'd34938, 16'd47150, 16'd32439, 16'd18394, 16'd36012, 16'd18536, 16'd36212, 16'd61687, 16'd28924, 16'd43245, 16'd15235});
	test_expansion(128'ha0f5d370b046d54e824ec0fb9abd5f0b, {16'd27301, 16'd28285, 16'd16191, 16'd20523, 16'd32354, 16'd50952, 16'd54167, 16'd56784, 16'd28386, 16'd48511, 16'd64257, 16'd46851, 16'd45550, 16'd40058, 16'd27774, 16'd20462, 16'd18823, 16'd14399, 16'd38973, 16'd52106, 16'd6776, 16'd59521, 16'd38267, 16'd6967, 16'd55596, 16'd46314});
	test_expansion(128'h86db6036546d8072e0ccb5468ea4bd54, {16'd18280, 16'd60811, 16'd878, 16'd33482, 16'd56377, 16'd46611, 16'd54848, 16'd53569, 16'd37142, 16'd32791, 16'd43017, 16'd8378, 16'd45940, 16'd40284, 16'd4788, 16'd40941, 16'd18485, 16'd40453, 16'd5353, 16'd56759, 16'd48736, 16'd38372, 16'd29213, 16'd50854, 16'd19431, 16'd6071});
	test_expansion(128'h5d0ec09d127c7a38f4c6d53a5a341e69, {16'd45686, 16'd64039, 16'd21454, 16'd27167, 16'd23245, 16'd7649, 16'd60747, 16'd44385, 16'd64723, 16'd6307, 16'd9011, 16'd5845, 16'd34537, 16'd31121, 16'd30452, 16'd54477, 16'd33817, 16'd35029, 16'd12413, 16'd60223, 16'd42908, 16'd64407, 16'd17410, 16'd16212, 16'd633, 16'd62661});
	test_expansion(128'hff2efc6ea7504394db03da11c20d3abb, {16'd15912, 16'd13083, 16'd45447, 16'd15580, 16'd24923, 16'd35830, 16'd55603, 16'd36314, 16'd62263, 16'd29002, 16'd55390, 16'd22515, 16'd13956, 16'd6212, 16'd56620, 16'd19082, 16'd19426, 16'd31174, 16'd13991, 16'd14428, 16'd54550, 16'd20276, 16'd8408, 16'd53930, 16'd17328, 16'd37783});
	test_expansion(128'h62697d47a765a18ccd87be62bd213f02, {16'd41883, 16'd38054, 16'd48969, 16'd25571, 16'd10577, 16'd39071, 16'd39094, 16'd26538, 16'd55692, 16'd63764, 16'd3741, 16'd22175, 16'd41679, 16'd30772, 16'd38150, 16'd55059, 16'd19029, 16'd7860, 16'd31973, 16'd13308, 16'd52630, 16'd28051, 16'd21730, 16'd39028, 16'd47116, 16'd64351});
	test_expansion(128'h6779a14e167d4a9e32eee388b1af6b76, {16'd30406, 16'd51078, 16'd48873, 16'd38639, 16'd6983, 16'd3525, 16'd56306, 16'd51897, 16'd41830, 16'd27975, 16'd65518, 16'd26812, 16'd27077, 16'd29786, 16'd12702, 16'd13195, 16'd38276, 16'd34542, 16'd12767, 16'd25838, 16'd42099, 16'd27393, 16'd30458, 16'd53494, 16'd28586, 16'd52644});
	test_expansion(128'h308c28017000438572bbd0354fa31c15, {16'd38375, 16'd39822, 16'd58393, 16'd63325, 16'd44646, 16'd2080, 16'd17717, 16'd49094, 16'd23453, 16'd57116, 16'd3934, 16'd31855, 16'd57292, 16'd7697, 16'd41057, 16'd1980, 16'd62012, 16'd53546, 16'd31278, 16'd22446, 16'd46777, 16'd23257, 16'd56950, 16'd21103, 16'd31789, 16'd41833});
	test_expansion(128'hfc47dad1e8cffc9ae3c7ce994b530f90, {16'd55693, 16'd58614, 16'd12024, 16'd61182, 16'd17255, 16'd13474, 16'd24698, 16'd28794, 16'd37415, 16'd55193, 16'd3376, 16'd58510, 16'd36253, 16'd44929, 16'd10086, 16'd17706, 16'd19665, 16'd64398, 16'd21260, 16'd34127, 16'd26270, 16'd34872, 16'd25093, 16'd15833, 16'd58203, 16'd8639});
	test_expansion(128'h7654e1e70e00e16f0a6f9187f0b4d22f, {16'd2216, 16'd2569, 16'd32475, 16'd46774, 16'd58339, 16'd49224, 16'd25569, 16'd9964, 16'd4787, 16'd45003, 16'd6554, 16'd61549, 16'd40717, 16'd54895, 16'd53658, 16'd64330, 16'd62007, 16'd41617, 16'd52749, 16'd62649, 16'd53253, 16'd46695, 16'd50543, 16'd36785, 16'd63895, 16'd64172});
	test_expansion(128'hbf12207bedeaa9b95b03af0bf40149c8, {16'd43122, 16'd3388, 16'd36745, 16'd11793, 16'd15640, 16'd23208, 16'd39154, 16'd58620, 16'd64791, 16'd4999, 16'd15097, 16'd62660, 16'd39302, 16'd65490, 16'd1784, 16'd18492, 16'd22381, 16'd125, 16'd57026, 16'd30648, 16'd59268, 16'd4693, 16'd5565, 16'd10624, 16'd5010, 16'd7138});
	test_expansion(128'he84454e1e889c9a542baede537ce0b13, {16'd57325, 16'd28450, 16'd5805, 16'd32306, 16'd40686, 16'd30771, 16'd39688, 16'd10670, 16'd14735, 16'd21828, 16'd41725, 16'd53561, 16'd17452, 16'd54015, 16'd57714, 16'd55251, 16'd17578, 16'd50570, 16'd22035, 16'd28860, 16'd27903, 16'd52631, 16'd40093, 16'd16597, 16'd8599, 16'd23978});
	test_expansion(128'ha773b0c17b8e33e38f55f260a7825dd6, {16'd24668, 16'd46318, 16'd18517, 16'd64235, 16'd62603, 16'd51082, 16'd6329, 16'd49321, 16'd33951, 16'd48394, 16'd3912, 16'd54830, 16'd38047, 16'd48639, 16'd24705, 16'd34912, 16'd44059, 16'd2763, 16'd4883, 16'd61721, 16'd49253, 16'd41790, 16'd19225, 16'd28686, 16'd64805, 16'd55059});
	test_expansion(128'h4d9a666f6f2448d92bd2f29509511627, {16'd57570, 16'd1193, 16'd6583, 16'd35795, 16'd65356, 16'd4054, 16'd56640, 16'd49839, 16'd26731, 16'd64142, 16'd16821, 16'd12381, 16'd15405, 16'd39834, 16'd12076, 16'd52585, 16'd5536, 16'd56756, 16'd7508, 16'd29677, 16'd27247, 16'd8856, 16'd26990, 16'd13030, 16'd16714, 16'd28304});
	test_expansion(128'h8f3eae81d84eb63fb0cd33564ff6f8ea, {16'd17676, 16'd27552, 16'd44190, 16'd27389, 16'd5917, 16'd61864, 16'd9697, 16'd14483, 16'd55549, 16'd34826, 16'd45632, 16'd7158, 16'd64125, 16'd43341, 16'd49239, 16'd37152, 16'd6277, 16'd65511, 16'd58969, 16'd13561, 16'd34977, 16'd27927, 16'd6013, 16'd25581, 16'd2894, 16'd33282});
	test_expansion(128'hbdc9a7af9c3bf74c9a788872f03afac9, {16'd24013, 16'd55551, 16'd64762, 16'd37219, 16'd16767, 16'd29988, 16'd49518, 16'd58521, 16'd53035, 16'd34023, 16'd52281, 16'd38438, 16'd1662, 16'd25687, 16'd18918, 16'd14540, 16'd39364, 16'd29434, 16'd1687, 16'd43805, 16'd41576, 16'd46807, 16'd6268, 16'd1580, 16'd41511, 16'd4995});
	test_expansion(128'h3810732a31d98e7a7eef3b4734d10246, {16'd35191, 16'd11647, 16'd52135, 16'd11359, 16'd14218, 16'd57142, 16'd33247, 16'd50256, 16'd8118, 16'd16122, 16'd42094, 16'd37602, 16'd62386, 16'd39990, 16'd39534, 16'd53460, 16'd6511, 16'd50476, 16'd22651, 16'd59729, 16'd30898, 16'd41147, 16'd10078, 16'd15045, 16'd13876, 16'd19557});
	test_expansion(128'h1e4c944d628d0be662c8aa8bf93fb293, {16'd43923, 16'd35575, 16'd35761, 16'd54661, 16'd59055, 16'd53447, 16'd24881, 16'd11728, 16'd32387, 16'd58351, 16'd61086, 16'd15248, 16'd1171, 16'd65000, 16'd51276, 16'd62784, 16'd48622, 16'd30000, 16'd36755, 16'd40469, 16'd29326, 16'd50834, 16'd45197, 16'd40241, 16'd436, 16'd62666});
	test_expansion(128'hb911ede7c0c058f92cfc02573463d51f, {16'd2575, 16'd64369, 16'd35530, 16'd2138, 16'd59956, 16'd13754, 16'd28982, 16'd39848, 16'd17776, 16'd57272, 16'd54100, 16'd4775, 16'd37237, 16'd46045, 16'd24658, 16'd38223, 16'd7012, 16'd32344, 16'd22886, 16'd57222, 16'd58952, 16'd39538, 16'd12424, 16'd53210, 16'd48340, 16'd50499});
	test_expansion(128'hfb0541eb1120e0f5880c72d2bfc1749b, {16'd7463, 16'd54871, 16'd15541, 16'd24209, 16'd56940, 16'd1179, 16'd30749, 16'd3843, 16'd47473, 16'd32890, 16'd27769, 16'd16314, 16'd15866, 16'd45508, 16'd24900, 16'd3246, 16'd7359, 16'd22202, 16'd60437, 16'd63612, 16'd61280, 16'd8338, 16'd28216, 16'd17643, 16'd28648, 16'd41597});
	test_expansion(128'h26c55abd9118bc2e2bda78d343ee493e, {16'd64848, 16'd45529, 16'd6227, 16'd16902, 16'd29039, 16'd15138, 16'd52973, 16'd23066, 16'd36923, 16'd5626, 16'd10112, 16'd6433, 16'd21881, 16'd27951, 16'd30317, 16'd29369, 16'd56858, 16'd47182, 16'd44155, 16'd34865, 16'd1286, 16'd30859, 16'd28694, 16'd5834, 16'd37395, 16'd17145});
	test_expansion(128'h06092cd973f6ffab4ecde0d080a3cd29, {16'd6055, 16'd10965, 16'd15244, 16'd56129, 16'd60872, 16'd47011, 16'd49255, 16'd47374, 16'd52426, 16'd35507, 16'd31311, 16'd29494, 16'd11015, 16'd15585, 16'd49925, 16'd1482, 16'd5422, 16'd53472, 16'd57581, 16'd64798, 16'd4112, 16'd6078, 16'd7357, 16'd9696, 16'd8387, 16'd26900});
	test_expansion(128'h4bc3b70fb773e801c3dee249446e7705, {16'd16745, 16'd53258, 16'd59003, 16'd44939, 16'd13957, 16'd18352, 16'd23873, 16'd2125, 16'd6504, 16'd23839, 16'd22228, 16'd34899, 16'd53249, 16'd6797, 16'd57535, 16'd15219, 16'd15970, 16'd45920, 16'd53114, 16'd12960, 16'd44486, 16'd8593, 16'd36088, 16'd32807, 16'd54570, 16'd64716});
	test_expansion(128'h2b59679e295b9d59b08331b147fbf0a9, {16'd879, 16'd18490, 16'd3173, 16'd28854, 16'd39111, 16'd63304, 16'd39153, 16'd27684, 16'd25086, 16'd25642, 16'd19228, 16'd47908, 16'd57248, 16'd915, 16'd37716, 16'd7418, 16'd15094, 16'd33245, 16'd11479, 16'd26430, 16'd64951, 16'd65439, 16'd1681, 16'd39127, 16'd1619, 16'd3885});
	test_expansion(128'hc10530f056784d168441cd97cc04c300, {16'd47673, 16'd58549, 16'd62428, 16'd2992, 16'd46598, 16'd21169, 16'd29346, 16'd3429, 16'd19700, 16'd31688, 16'd39422, 16'd63982, 16'd31747, 16'd27762, 16'd27357, 16'd3494, 16'd13828, 16'd8892, 16'd40820, 16'd43410, 16'd39956, 16'd5900, 16'd21557, 16'd20736, 16'd12488, 16'd27930});
	test_expansion(128'hf4cbfa90d1d28f7c63ce017cb5b43053, {16'd54296, 16'd29732, 16'd16624, 16'd48833, 16'd64505, 16'd36600, 16'd16816, 16'd18234, 16'd32435, 16'd6485, 16'd8732, 16'd19961, 16'd16034, 16'd65239, 16'd8569, 16'd60840, 16'd12549, 16'd15349, 16'd35384, 16'd48510, 16'd2584, 16'd45703, 16'd55220, 16'd14369, 16'd59569, 16'd45618});
	test_expansion(128'h1936f73f8a93373e6a33238ad36efccc, {16'd3037, 16'd14180, 16'd48408, 16'd37506, 16'd29487, 16'd45666, 16'd1161, 16'd58851, 16'd36606, 16'd3707, 16'd5396, 16'd4991, 16'd42181, 16'd59941, 16'd63582, 16'd42998, 16'd55934, 16'd9729, 16'd34717, 16'd12046, 16'd5601, 16'd44006, 16'd54204, 16'd44195, 16'd24492, 16'd3149});
	test_expansion(128'ha019c9e38c8b4bc4beec9f0c43a746e3, {16'd23646, 16'd50220, 16'd42828, 16'd39256, 16'd10853, 16'd6674, 16'd26709, 16'd18925, 16'd29554, 16'd9650, 16'd49219, 16'd2199, 16'd41216, 16'd46467, 16'd32129, 16'd53260, 16'd19200, 16'd55188, 16'd19538, 16'd60103, 16'd30635, 16'd1619, 16'd17478, 16'd49490, 16'd26886, 16'd46955});
	test_expansion(128'h1f7800e52acc5c754a16e8a606fef417, {16'd6082, 16'd493, 16'd65068, 16'd17208, 16'd12005, 16'd48100, 16'd40519, 16'd51019, 16'd23313, 16'd48334, 16'd32825, 16'd30638, 16'd43999, 16'd36803, 16'd40974, 16'd9675, 16'd10722, 16'd25125, 16'd37860, 16'd35429, 16'd48529, 16'd20643, 16'd38159, 16'd24142, 16'd35113, 16'd48966});
	test_expansion(128'h158d08e853f8eba9b20a9b316d831b79, {16'd6267, 16'd29661, 16'd27824, 16'd53507, 16'd14859, 16'd21319, 16'd51073, 16'd33501, 16'd13632, 16'd62970, 16'd34631, 16'd32713, 16'd29657, 16'd59457, 16'd55978, 16'd26965, 16'd53755, 16'd35735, 16'd6126, 16'd31486, 16'd43081, 16'd62282, 16'd17875, 16'd9378, 16'd51017, 16'd18406});
	test_expansion(128'h13de87ccda1b3b40e95f751a6b5eefd2, {16'd22073, 16'd28017, 16'd36959, 16'd20579, 16'd2837, 16'd2752, 16'd3088, 16'd54250, 16'd39070, 16'd15994, 16'd49398, 16'd58456, 16'd9465, 16'd2903, 16'd55006, 16'd17975, 16'd61954, 16'd37429, 16'd7243, 16'd59424, 16'd6237, 16'd8742, 16'd4429, 16'd57833, 16'd31493, 16'd22476});
	test_expansion(128'h271c4baa8c7090a978684d521f568719, {16'd62069, 16'd4285, 16'd3429, 16'd56021, 16'd64656, 16'd7105, 16'd56489, 16'd22096, 16'd54443, 16'd56709, 16'd4228, 16'd59294, 16'd44556, 16'd24351, 16'd9936, 16'd57598, 16'd27088, 16'd15010, 16'd27585, 16'd11164, 16'd32918, 16'd15277, 16'd17626, 16'd6891, 16'd51834, 16'd43371});
	test_expansion(128'h623b2a4607882c09bfea800c04cd4e39, {16'd38425, 16'd12445, 16'd62841, 16'd11718, 16'd24439, 16'd15246, 16'd43577, 16'd16430, 16'd9254, 16'd62100, 16'd42994, 16'd50899, 16'd51428, 16'd11730, 16'd19343, 16'd23357, 16'd40841, 16'd62660, 16'd31799, 16'd33885, 16'd14065, 16'd35624, 16'd39430, 16'd456, 16'd55551, 16'd18099});
	test_expansion(128'h11b42c3d328e323f1ab1575ab24a10ff, {16'd4220, 16'd23407, 16'd6087, 16'd1309, 16'd49155, 16'd38694, 16'd14609, 16'd4145, 16'd20491, 16'd54010, 16'd28773, 16'd46006, 16'd29888, 16'd63234, 16'd19319, 16'd4600, 16'd16395, 16'd9838, 16'd3902, 16'd61563, 16'd43074, 16'd52686, 16'd9949, 16'd13021, 16'd37986, 16'd7636});
	test_expansion(128'hdca7eea15e66890c5d444c58165fe154, {16'd56699, 16'd30865, 16'd11455, 16'd23675, 16'd29081, 16'd827, 16'd57467, 16'd9363, 16'd16565, 16'd6567, 16'd36147, 16'd57227, 16'd39648, 16'd64395, 16'd41628, 16'd11870, 16'd13062, 16'd6579, 16'd49778, 16'd54352, 16'd23641, 16'd38415, 16'd19590, 16'd15236, 16'd12833, 16'd7192});
	test_expansion(128'h619d84b02a665406406f0f2e82b94edb, {16'd31287, 16'd7557, 16'd7434, 16'd26445, 16'd23341, 16'd45371, 16'd40375, 16'd63663, 16'd37573, 16'd37525, 16'd49213, 16'd14523, 16'd3146, 16'd4989, 16'd13538, 16'd51349, 16'd64022, 16'd48292, 16'd38102, 16'd12015, 16'd19292, 16'd12666, 16'd61322, 16'd12197, 16'd43280, 16'd1441});
	test_expansion(128'hb073cce7192e348e05a080320a1f0906, {16'd26965, 16'd47738, 16'd58040, 16'd20815, 16'd8538, 16'd44834, 16'd56513, 16'd48359, 16'd64389, 16'd36493, 16'd29725, 16'd11945, 16'd43472, 16'd12407, 16'd31349, 16'd31365, 16'd51625, 16'd14891, 16'd19286, 16'd34604, 16'd38831, 16'd42495, 16'd10538, 16'd15244, 16'd52366, 16'd10334});
	test_expansion(128'h57f8ff2870f65824768fe3f104683992, {16'd63511, 16'd31187, 16'd27985, 16'd53381, 16'd34271, 16'd59908, 16'd38665, 16'd42415, 16'd26310, 16'd23355, 16'd38214, 16'd10569, 16'd38660, 16'd33013, 16'd40537, 16'd17798, 16'd60485, 16'd9983, 16'd40701, 16'd52460, 16'd6281, 16'd55958, 16'd33915, 16'd37417, 16'd57634, 16'd39236});
	test_expansion(128'h0ceb8dbf0be059098ea503521b2fe5f1, {16'd60545, 16'd59504, 16'd57508, 16'd41217, 16'd46115, 16'd32599, 16'd31216, 16'd50125, 16'd11076, 16'd43734, 16'd11652, 16'd50555, 16'd58471, 16'd22712, 16'd62656, 16'd50330, 16'd51839, 16'd41614, 16'd8620, 16'd22212, 16'd53143, 16'd57246, 16'd26027, 16'd27983, 16'd49168, 16'd29702});
	test_expansion(128'hed83c6bda02e34f51a39e7bd6808932b, {16'd60204, 16'd53114, 16'd3668, 16'd47983, 16'd5889, 16'd38133, 16'd30344, 16'd22733, 16'd27304, 16'd64226, 16'd30458, 16'd27752, 16'd20674, 16'd63164, 16'd16918, 16'd49452, 16'd64682, 16'd27951, 16'd40010, 16'd5823, 16'd60366, 16'd37557, 16'd4562, 16'd31127, 16'd54281, 16'd33710});
	test_expansion(128'h9d1d2a1dc7eeac15b4a182d4f1f2ce15, {16'd38339, 16'd21089, 16'd12395, 16'd54964, 16'd23618, 16'd38649, 16'd49587, 16'd33343, 16'd37531, 16'd4643, 16'd18249, 16'd60086, 16'd13068, 16'd25159, 16'd705, 16'd35906, 16'd38690, 16'd25241, 16'd59002, 16'd21987, 16'd46781, 16'd31719, 16'd26858, 16'd6501, 16'd25497, 16'd33955});
	test_expansion(128'h2cc659986052a41025e07eacf2d1466f, {16'd11845, 16'd35071, 16'd13045, 16'd63609, 16'd36019, 16'd10622, 16'd32640, 16'd40334, 16'd39269, 16'd38852, 16'd39020, 16'd43975, 16'd55984, 16'd61071, 16'd21867, 16'd7743, 16'd26822, 16'd7449, 16'd13985, 16'd14764, 16'd59528, 16'd48259, 16'd62054, 16'd702, 16'd19714, 16'd21184});
	test_expansion(128'hd24839188ee71b3fe5b6ec2db2a8574f, {16'd46260, 16'd9096, 16'd28792, 16'd27126, 16'd26841, 16'd1353, 16'd47025, 16'd8245, 16'd18490, 16'd29829, 16'd13357, 16'd26716, 16'd23203, 16'd44120, 16'd61759, 16'd4716, 16'd8304, 16'd17898, 16'd8808, 16'd3932, 16'd17379, 16'd10485, 16'd3583, 16'd25458, 16'd3118, 16'd38459});
	test_expansion(128'h1362c77c4983968e10649e5a3303e37e, {16'd50356, 16'd35628, 16'd14743, 16'd21135, 16'd4751, 16'd46737, 16'd57418, 16'd3742, 16'd65168, 16'd16372, 16'd39465, 16'd57551, 16'd20154, 16'd64910, 16'd53714, 16'd104, 16'd18499, 16'd28928, 16'd64180, 16'd47014, 16'd54547, 16'd61061, 16'd7220, 16'd61833, 16'd14037, 16'd46000});
	test_expansion(128'hc8be824c9e84d1df013bce176ebe3b34, {16'd16515, 16'd54636, 16'd22901, 16'd59167, 16'd27245, 16'd28874, 16'd23526, 16'd22390, 16'd47188, 16'd22420, 16'd24852, 16'd5770, 16'd17498, 16'd32073, 16'd22114, 16'd20096, 16'd57100, 16'd13244, 16'd10576, 16'd61164, 16'd19003, 16'd60359, 16'd19212, 16'd38266, 16'd41300, 16'd41541});
	test_expansion(128'h82ad102327407c3c7ad2ec3c4d713a94, {16'd24518, 16'd18585, 16'd63325, 16'd33684, 16'd10573, 16'd33265, 16'd39000, 16'd63317, 16'd52524, 16'd58558, 16'd61367, 16'd58872, 16'd23534, 16'd43009, 16'd62837, 16'd14443, 16'd42317, 16'd19259, 16'd52586, 16'd9833, 16'd26040, 16'd46512, 16'd21378, 16'd10206, 16'd49239, 16'd25452});
	test_expansion(128'h50d985420b51c74065533533a445b419, {16'd58937, 16'd2107, 16'd6871, 16'd31017, 16'd34456, 16'd35119, 16'd30097, 16'd61528, 16'd56283, 16'd29297, 16'd34927, 16'd6042, 16'd14279, 16'd32354, 16'd48654, 16'd29287, 16'd27637, 16'd28112, 16'd16555, 16'd11088, 16'd2044, 16'd2814, 16'd64875, 16'd26718, 16'd11863, 16'd10498});
	test_expansion(128'h4483c3af9d431261a13087d7d3e72a9f, {16'd52675, 16'd57661, 16'd13534, 16'd56663, 16'd53652, 16'd51149, 16'd14747, 16'd48357, 16'd31693, 16'd58325, 16'd46900, 16'd33108, 16'd30226, 16'd17261, 16'd6091, 16'd20130, 16'd30988, 16'd44055, 16'd27429, 16'd16189, 16'd57722, 16'd50692, 16'd35924, 16'd63372, 16'd44023, 16'd18644});
	test_expansion(128'hc9df008fa04d5f7ba00e80780a113f6c, {16'd42586, 16'd21710, 16'd32706, 16'd4934, 16'd8935, 16'd5643, 16'd10343, 16'd65306, 16'd36934, 16'd56675, 16'd38864, 16'd17732, 16'd51548, 16'd54409, 16'd62266, 16'd12345, 16'd20214, 16'd42616, 16'd60169, 16'd53363, 16'd17715, 16'd4670, 16'd42619, 16'd17964, 16'd65120, 16'd34293});
	test_expansion(128'h3405b734f12bc7bbbbd0748a8ad4f23b, {16'd14517, 16'd61510, 16'd20854, 16'd17038, 16'd45264, 16'd19909, 16'd44734, 16'd12929, 16'd9256, 16'd49222, 16'd43054, 16'd12800, 16'd34314, 16'd52251, 16'd20031, 16'd36262, 16'd54881, 16'd62545, 16'd13904, 16'd59814, 16'd17356, 16'd49698, 16'd14115, 16'd39490, 16'd44620, 16'd60594});
	test_expansion(128'h89230e31db6e4229bd87d65ea7735ce4, {16'd15039, 16'd7704, 16'd1119, 16'd19515, 16'd38436, 16'd29426, 16'd61367, 16'd5677, 16'd30529, 16'd38579, 16'd63479, 16'd3492, 16'd47860, 16'd60614, 16'd5979, 16'd23053, 16'd38508, 16'd25624, 16'd34081, 16'd3594, 16'd65517, 16'd10453, 16'd17319, 16'd42723, 16'd6751, 16'd7328});
	test_expansion(128'hc988eaa462cfc381e172fb4b4b6a9812, {16'd21684, 16'd9138, 16'd57052, 16'd21525, 16'd20473, 16'd30989, 16'd51340, 16'd56542, 16'd26977, 16'd49416, 16'd19184, 16'd6531, 16'd52516, 16'd29442, 16'd1961, 16'd63161, 16'd2145, 16'd27798, 16'd8562, 16'd45835, 16'd560, 16'd35341, 16'd54094, 16'd41429, 16'd11291, 16'd42984});
	test_expansion(128'h43e4f0f227fb55b0719ebfd8b89efa20, {16'd51038, 16'd18979, 16'd53211, 16'd1533, 16'd37269, 16'd43173, 16'd49240, 16'd53136, 16'd60952, 16'd35987, 16'd52966, 16'd53162, 16'd14454, 16'd27364, 16'd7079, 16'd62753, 16'd58541, 16'd5127, 16'd23652, 16'd57107, 16'd28838, 16'd47695, 16'd50979, 16'd23085, 16'd19840, 16'd15971});
	test_expansion(128'hc340b18ccaa0263821e54fbbf8242482, {16'd40964, 16'd32638, 16'd32688, 16'd46512, 16'd35443, 16'd56510, 16'd40964, 16'd65231, 16'd7912, 16'd3444, 16'd48863, 16'd43281, 16'd43886, 16'd33886, 16'd64802, 16'd38198, 16'd15266, 16'd54925, 16'd59901, 16'd3887, 16'd27834, 16'd4574, 16'd44239, 16'd39726, 16'd20886, 16'd17056});
	test_expansion(128'h78b64a3dc50848a93bcbd346b7743a28, {16'd36412, 16'd42311, 16'd64060, 16'd8828, 16'd2289, 16'd41438, 16'd36360, 16'd38586, 16'd43593, 16'd46895, 16'd13894, 16'd63099, 16'd26868, 16'd64386, 16'd49617, 16'd61209, 16'd38989, 16'd33188, 16'd35566, 16'd31176, 16'd46706, 16'd45252, 16'd36103, 16'd51373, 16'd2706, 16'd43382});
	test_expansion(128'ha4ef485f9ae0ef3d9f1ba6f0151445bb, {16'd26926, 16'd58897, 16'd51819, 16'd46369, 16'd28631, 16'd34302, 16'd36287, 16'd32603, 16'd30282, 16'd36430, 16'd48302, 16'd49260, 16'd6339, 16'd53069, 16'd4631, 16'd33950, 16'd40985, 16'd41839, 16'd31006, 16'd48877, 16'd20254, 16'd60620, 16'd25536, 16'd34627, 16'd7657, 16'd22981});
	test_expansion(128'h44bd59a05a93165aefc70a9f29b3bcac, {16'd40592, 16'd31250, 16'd33139, 16'd11762, 16'd47837, 16'd31942, 16'd4997, 16'd10475, 16'd11414, 16'd47507, 16'd9121, 16'd35512, 16'd21040, 16'd24576, 16'd20241, 16'd11285, 16'd58977, 16'd19864, 16'd428, 16'd48193, 16'd29529, 16'd11513, 16'd13287, 16'd42877, 16'd58148, 16'd22761});
	test_expansion(128'hb4e82ca152287457b4470fe28ec416fc, {16'd3826, 16'd23414, 16'd8532, 16'd37080, 16'd22488, 16'd27144, 16'd53331, 16'd28757, 16'd5211, 16'd22952, 16'd45907, 16'd40717, 16'd1673, 16'd1269, 16'd61902, 16'd18178, 16'd437, 16'd63994, 16'd21699, 16'd23353, 16'd65107, 16'd5012, 16'd59771, 16'd28120, 16'd56010, 16'd36936});
	test_expansion(128'h4b88d15ccf0deef4357ddb39b47ba621, {16'd30280, 16'd57162, 16'd52443, 16'd15498, 16'd22781, 16'd17590, 16'd25884, 16'd42795, 16'd49982, 16'd45054, 16'd12508, 16'd46745, 16'd23257, 16'd59787, 16'd35974, 16'd26654, 16'd1004, 16'd49154, 16'd3902, 16'd15980, 16'd49383, 16'd64369, 16'd41617, 16'd48132, 16'd41195, 16'd34693});
	test_expansion(128'h25ba45888258e6dc41b3f6c5f2e92a85, {16'd51670, 16'd43183, 16'd9598, 16'd33273, 16'd19533, 16'd41423, 16'd22792, 16'd6368, 16'd15214, 16'd50698, 16'd39239, 16'd64314, 16'd37011, 16'd32403, 16'd2935, 16'd1553, 16'd54938, 16'd13101, 16'd27526, 16'd25046, 16'd13556, 16'd41403, 16'd4106, 16'd38682, 16'd30567, 16'd53322});
	test_expansion(128'hda551178b28bc6fec07c4e0b69a21e7f, {16'd64712, 16'd63380, 16'd27757, 16'd11330, 16'd23544, 16'd25998, 16'd43347, 16'd62983, 16'd49672, 16'd59839, 16'd36035, 16'd1701, 16'd15255, 16'd36017, 16'd30914, 16'd47298, 16'd52626, 16'd41329, 16'd4771, 16'd27197, 16'd28997, 16'd28035, 16'd49911, 16'd1293, 16'd24276, 16'd33517});
	test_expansion(128'he812b8bb60891bb8cdd4205b30ad6191, {16'd34513, 16'd63101, 16'd63877, 16'd8760, 16'd59698, 16'd45390, 16'd52147, 16'd3037, 16'd3265, 16'd26063, 16'd37990, 16'd33511, 16'd53422, 16'd39402, 16'd27180, 16'd59009, 16'd33286, 16'd41705, 16'd20041, 16'd45667, 16'd16783, 16'd50457, 16'd3014, 16'd48268, 16'd32949, 16'd62572});
	test_expansion(128'h92cdc9af59ba241ab8e7a6a41d365bc7, {16'd46555, 16'd35641, 16'd1457, 16'd64457, 16'd60315, 16'd61259, 16'd30686, 16'd41376, 16'd33943, 16'd40044, 16'd1516, 16'd63470, 16'd50114, 16'd20526, 16'd50910, 16'd17526, 16'd36924, 16'd14431, 16'd55754, 16'd43288, 16'd9776, 16'd9719, 16'd59111, 16'd39865, 16'd13169, 16'd518});
	test_expansion(128'h9c27009603b58098691bd719c8005422, {16'd50430, 16'd38601, 16'd3351, 16'd58026, 16'd37058, 16'd25023, 16'd40895, 16'd15275, 16'd30469, 16'd55763, 16'd6052, 16'd26957, 16'd23379, 16'd47717, 16'd48421, 16'd15046, 16'd12421, 16'd20458, 16'd6350, 16'd31736, 16'd9499, 16'd12455, 16'd39961, 16'd17247, 16'd57809, 16'd5146});
	test_expansion(128'h9906076b8bb52f101c6f11c5b8317792, {16'd29455, 16'd48796, 16'd50405, 16'd47772, 16'd9241, 16'd20593, 16'd14966, 16'd20946, 16'd40405, 16'd50752, 16'd40599, 16'd22652, 16'd48547, 16'd5795, 16'd54899, 16'd31016, 16'd25143, 16'd32208, 16'd11432, 16'd29651, 16'd7191, 16'd35211, 16'd956, 16'd64695, 16'd53859, 16'd25637});
	test_expansion(128'h435f2b30fa55fc164669a258ff876fe2, {16'd59299, 16'd35706, 16'd11392, 16'd30709, 16'd17212, 16'd21039, 16'd32446, 16'd21707, 16'd58881, 16'd42810, 16'd47352, 16'd18786, 16'd26110, 16'd21517, 16'd15406, 16'd7094, 16'd10113, 16'd56995, 16'd20671, 16'd60618, 16'd10768, 16'd34852, 16'd834, 16'd63539, 16'd37783, 16'd51996});
	test_expansion(128'h42a4edbe0efad0447da42671367bda29, {16'd44533, 16'd46345, 16'd52804, 16'd34572, 16'd8923, 16'd29854, 16'd37373, 16'd36902, 16'd44886, 16'd20831, 16'd51474, 16'd6108, 16'd25952, 16'd60605, 16'd37121, 16'd24139, 16'd34711, 16'd42245, 16'd5781, 16'd57586, 16'd11280, 16'd13431, 16'd47158, 16'd57049, 16'd60230, 16'd58296});
	test_expansion(128'h439db27d539ef9f8aaa414597b28a96e, {16'd30845, 16'd60783, 16'd24690, 16'd59414, 16'd6347, 16'd24458, 16'd5971, 16'd62659, 16'd64487, 16'd63971, 16'd24132, 16'd52158, 16'd54594, 16'd7185, 16'd12240, 16'd61255, 16'd42010, 16'd45727, 16'd43254, 16'd29128, 16'd35108, 16'd45396, 16'd1540, 16'd43742, 16'd30970, 16'd22284});
	test_expansion(128'hc57db21ce9fb4e41c61adc6a0880611c, {16'd36435, 16'd15937, 16'd19796, 16'd53084, 16'd26964, 16'd30691, 16'd6759, 16'd47825, 16'd43343, 16'd63504, 16'd22507, 16'd53639, 16'd34282, 16'd22762, 16'd60138, 16'd34479, 16'd2913, 16'd13228, 16'd51721, 16'd7269, 16'd9237, 16'd38111, 16'd36405, 16'd61449, 16'd7927, 16'd59264});
	test_expansion(128'hde0ee4eb1027eabdce28c8ca03ddf44c, {16'd30251, 16'd7649, 16'd49083, 16'd8847, 16'd43213, 16'd8670, 16'd60507, 16'd4843, 16'd30576, 16'd27079, 16'd47816, 16'd15006, 16'd6135, 16'd41774, 16'd39787, 16'd41494, 16'd8985, 16'd18553, 16'd60469, 16'd6162, 16'd43504, 16'd17614, 16'd4908, 16'd8539, 16'd52060, 16'd40496});
	test_expansion(128'h540987cded8c6dc8e45a8b60613884c9, {16'd46087, 16'd46533, 16'd29416, 16'd2564, 16'd51400, 16'd43956, 16'd62289, 16'd54369, 16'd20305, 16'd48616, 16'd37390, 16'd33452, 16'd53455, 16'd16029, 16'd46574, 16'd23528, 16'd45611, 16'd57627, 16'd35229, 16'd62137, 16'd8117, 16'd21360, 16'd50465, 16'd33910, 16'd6122, 16'd33241});
	test_expansion(128'h8df9b389b1bc32a57637853c62b14908, {16'd12528, 16'd39233, 16'd375, 16'd31827, 16'd47126, 16'd39685, 16'd61071, 16'd35296, 16'd25229, 16'd35449, 16'd45360, 16'd47184, 16'd12584, 16'd59744, 16'd10259, 16'd81, 16'd9157, 16'd1401, 16'd10320, 16'd18538, 16'd28270, 16'd53164, 16'd57197, 16'd12867, 16'd21635, 16'd15710});
	test_expansion(128'h8bfe16ca7bc3380afda04b6cde146cde, {16'd59700, 16'd42870, 16'd11096, 16'd29629, 16'd46264, 16'd62704, 16'd55282, 16'd12231, 16'd12433, 16'd12250, 16'd54101, 16'd62865, 16'd23064, 16'd40093, 16'd19192, 16'd1960, 16'd53822, 16'd29667, 16'd20194, 16'd1014, 16'd33986, 16'd29882, 16'd61528, 16'd20911, 16'd40973, 16'd12949});
	test_expansion(128'hfb949428eee134ac84fa0d87c5b115f2, {16'd54429, 16'd27355, 16'd28000, 16'd19143, 16'd19965, 16'd21574, 16'd49329, 16'd43621, 16'd30839, 16'd6374, 16'd20105, 16'd26547, 16'd49394, 16'd44358, 16'd49572, 16'd57538, 16'd20624, 16'd50609, 16'd19933, 16'd35695, 16'd2280, 16'd16780, 16'd47374, 16'd16021, 16'd53120, 16'd23214});
	test_expansion(128'h75fa956890adf6c6325268441f929ec7, {16'd43723, 16'd29019, 16'd56166, 16'd21871, 16'd37575, 16'd16939, 16'd30584, 16'd5145, 16'd41641, 16'd19848, 16'd37069, 16'd63088, 16'd63772, 16'd19875, 16'd12946, 16'd25815, 16'd55084, 16'd29957, 16'd589, 16'd5341, 16'd17249, 16'd5534, 16'd21918, 16'd56772, 16'd57841, 16'd23924});
	test_expansion(128'he8196e4973aead5a3d022cd92aaa1a0a, {16'd23260, 16'd62971, 16'd57396, 16'd33264, 16'd58526, 16'd38450, 16'd32703, 16'd31388, 16'd10170, 16'd37839, 16'd32649, 16'd47500, 16'd57825, 16'd35521, 16'd60746, 16'd40628, 16'd6776, 16'd62827, 16'd45383, 16'd24779, 16'd49292, 16'd47679, 16'd913, 16'd17254, 16'd38389, 16'd62981});
	test_expansion(128'hda7f8828c1b854d2b242e766f2a115c6, {16'd54005, 16'd27043, 16'd47173, 16'd58319, 16'd35767, 16'd31724, 16'd62938, 16'd29680, 16'd60719, 16'd27971, 16'd51901, 16'd14250, 16'd31413, 16'd7988, 16'd61961, 16'd15982, 16'd13728, 16'd57782, 16'd30695, 16'd44434, 16'd42681, 16'd41184, 16'd52810, 16'd51119, 16'd4367, 16'd2873});
	test_expansion(128'hbe875a2e83cc78ac992366596caeba46, {16'd15017, 16'd54263, 16'd41992, 16'd7704, 16'd30287, 16'd38796, 16'd23753, 16'd6400, 16'd15645, 16'd2822, 16'd56326, 16'd55274, 16'd51571, 16'd48905, 16'd65208, 16'd33901, 16'd50440, 16'd46842, 16'd59136, 16'd21398, 16'd60499, 16'd9064, 16'd39251, 16'd42415, 16'd47438, 16'd38325});
	test_expansion(128'h775bf445eccd0aaca6439d8174d0a435, {16'd2839, 16'd16749, 16'd57548, 16'd20793, 16'd11692, 16'd64385, 16'd14035, 16'd12338, 16'd64492, 16'd4292, 16'd63381, 16'd7634, 16'd20460, 16'd55709, 16'd45409, 16'd4338, 16'd4797, 16'd62253, 16'd8243, 16'd61914, 16'd64524, 16'd28929, 16'd38790, 16'd42652, 16'd46534, 16'd61560});
	test_expansion(128'h2eb41e22902fa2a2ab618ee0d6c91117, {16'd20856, 16'd44815, 16'd12325, 16'd32422, 16'd12621, 16'd33365, 16'd56495, 16'd64105, 16'd63493, 16'd61051, 16'd23743, 16'd49544, 16'd36065, 16'd49905, 16'd28530, 16'd16113, 16'd48084, 16'd57073, 16'd9213, 16'd44188, 16'd56372, 16'd64387, 16'd40849, 16'd21908, 16'd53573, 16'd33928});
	test_expansion(128'heeb1cc69e5c317091453874c8ce904c2, {16'd6017, 16'd35491, 16'd51447, 16'd10089, 16'd27276, 16'd63157, 16'd58751, 16'd14362, 16'd9425, 16'd5945, 16'd24828, 16'd5851, 16'd573, 16'd57079, 16'd18149, 16'd13301, 16'd23464, 16'd46060, 16'd38029, 16'd62487, 16'd17196, 16'd655, 16'd47553, 16'd63941, 16'd62293, 16'd52628});
	test_expansion(128'h0a27834b72aff2e010134022e6145efb, {16'd56030, 16'd52436, 16'd57868, 16'd26609, 16'd54457, 16'd55551, 16'd34563, 16'd17108, 16'd13081, 16'd10659, 16'd8606, 16'd53322, 16'd9777, 16'd61878, 16'd24011, 16'd18783, 16'd48481, 16'd8677, 16'd15910, 16'd42494, 16'd48510, 16'd1789, 16'd35589, 16'd8292, 16'd9204, 16'd1728});
	test_expansion(128'h7dc613b7ed1cf9c64d91dd916cfc3f37, {16'd9062, 16'd46569, 16'd42012, 16'd16869, 16'd13660, 16'd18317, 16'd35678, 16'd28715, 16'd19362, 16'd48620, 16'd21797, 16'd52521, 16'd42454, 16'd28592, 16'd58143, 16'd40912, 16'd50678, 16'd28195, 16'd56280, 16'd50885, 16'd50550, 16'd4954, 16'd23815, 16'd35751, 16'd12600, 16'd29854});
	test_expansion(128'h6978bfa8288524c4e8405f7af65cd1c2, {16'd8725, 16'd15557, 16'd25932, 16'd38763, 16'd15618, 16'd37482, 16'd60126, 16'd39019, 16'd59475, 16'd13531, 16'd5333, 16'd33072, 16'd25070, 16'd46307, 16'd31900, 16'd6955, 16'd21052, 16'd1667, 16'd29314, 16'd37064, 16'd28813, 16'd32604, 16'd10709, 16'd8032, 16'd18093, 16'd25486});
	test_expansion(128'h310b3828da49602a6c39ad0f15c1a0df, {16'd21952, 16'd25556, 16'd33042, 16'd4970, 16'd39641, 16'd18757, 16'd13849, 16'd38253, 16'd53369, 16'd6872, 16'd43641, 16'd45573, 16'd49285, 16'd64651, 16'd25767, 16'd7613, 16'd34318, 16'd24288, 16'd10839, 16'd52539, 16'd45214, 16'd48413, 16'd24355, 16'd58573, 16'd4421, 16'd18171});
	test_expansion(128'h35c2c993c22b2b84ae0c8e940dd36c3a, {16'd64295, 16'd40609, 16'd55473, 16'd45401, 16'd5001, 16'd56450, 16'd15386, 16'd14877, 16'd39658, 16'd36509, 16'd17523, 16'd17357, 16'd63999, 16'd32595, 16'd5152, 16'd45829, 16'd15090, 16'd32407, 16'd17810, 16'd43413, 16'd10384, 16'd9952, 16'd28760, 16'd7550, 16'd8204, 16'd58016});
	test_expansion(128'ha661eec14c7b669fa1ca1c4ff122e247, {16'd2271, 16'd49893, 16'd38824, 16'd41239, 16'd23043, 16'd62692, 16'd60613, 16'd61805, 16'd26838, 16'd24266, 16'd19855, 16'd48849, 16'd11438, 16'd334, 16'd46366, 16'd60306, 16'd30434, 16'd14253, 16'd34148, 16'd64944, 16'd20643, 16'd63576, 16'd42480, 16'd60574, 16'd19073, 16'd60833});
	test_expansion(128'h718ab03710d13be4bce1c77d818a2682, {16'd23163, 16'd30627, 16'd7318, 16'd3516, 16'd43845, 16'd36119, 16'd7163, 16'd40537, 16'd5159, 16'd28345, 16'd12792, 16'd1129, 16'd28336, 16'd65027, 16'd50754, 16'd27470, 16'd40012, 16'd32479, 16'd64504, 16'd32180, 16'd24648, 16'd53875, 16'd6885, 16'd53219, 16'd50437, 16'd47448});
	test_expansion(128'h7c707feffd34adc8416b2f077d04f1f6, {16'd31313, 16'd54556, 16'd5877, 16'd19145, 16'd16248, 16'd35036, 16'd48887, 16'd40796, 16'd63564, 16'd10635, 16'd18759, 16'd23214, 16'd43289, 16'd27726, 16'd35702, 16'd20229, 16'd45519, 16'd21162, 16'd24715, 16'd64319, 16'd54509, 16'd6730, 16'd40801, 16'd21323, 16'd15606, 16'd25633});
	test_expansion(128'h62c8b46ec25b093964a40be723c8466d, {16'd15201, 16'd63264, 16'd6424, 16'd314, 16'd4500, 16'd5636, 16'd28367, 16'd30522, 16'd14374, 16'd10619, 16'd34243, 16'd32075, 16'd38699, 16'd42743, 16'd33039, 16'd7584, 16'd59159, 16'd50849, 16'd36986, 16'd49417, 16'd38467, 16'd6764, 16'd13112, 16'd3867, 16'd7641, 16'd32632});
	test_expansion(128'he1358fa184cdc61caff3a7d6df259d49, {16'd52157, 16'd12233, 16'd7898, 16'd23673, 16'd63203, 16'd1817, 16'd38710, 16'd48491, 16'd36333, 16'd8739, 16'd41453, 16'd55827, 16'd3183, 16'd60094, 16'd19592, 16'd46152, 16'd18270, 16'd57814, 16'd53274, 16'd57539, 16'd59300, 16'd48417, 16'd39370, 16'd41719, 16'd38122, 16'd31332});
	test_expansion(128'h0782ff52af8340fa6096183e596b72e7, {16'd63400, 16'd16732, 16'd25344, 16'd36921, 16'd43285, 16'd62103, 16'd30322, 16'd24510, 16'd18292, 16'd52073, 16'd46899, 16'd61570, 16'd26259, 16'd58819, 16'd11949, 16'd48268, 16'd32518, 16'd44439, 16'd36342, 16'd12589, 16'd15450, 16'd20236, 16'd32608, 16'd15030, 16'd56538, 16'd41016});
	test_expansion(128'he4954e49bc82d09274933d9171122a26, {16'd2542, 16'd20955, 16'd46716, 16'd36147, 16'd714, 16'd4299, 16'd30970, 16'd30563, 16'd53785, 16'd38209, 16'd22807, 16'd30624, 16'd50958, 16'd32507, 16'd51031, 16'd18054, 16'd4087, 16'd63480, 16'd36625, 16'd9188, 16'd3612, 16'd1045, 16'd46955, 16'd33448, 16'd23086, 16'd40739});
	test_expansion(128'he8b8129e0d077bc751515d7938305fdb, {16'd9715, 16'd626, 16'd38634, 16'd35771, 16'd5342, 16'd38407, 16'd14434, 16'd50283, 16'd37517, 16'd11268, 16'd4912, 16'd34824, 16'd29044, 16'd14010, 16'd39353, 16'd48175, 16'd5543, 16'd57892, 16'd23008, 16'd54539, 16'd25163, 16'd48653, 16'd3059, 16'd49167, 16'd22775, 16'd9800});
	test_expansion(128'h755ffe266f1efa836b74b2bd8406c945, {16'd16770, 16'd4470, 16'd54787, 16'd30293, 16'd59633, 16'd1775, 16'd27256, 16'd20309, 16'd26835, 16'd33237, 16'd5790, 16'd2594, 16'd31789, 16'd5513, 16'd13981, 16'd20868, 16'd27953, 16'd7595, 16'd43456, 16'd64369, 16'd11956, 16'd25081, 16'd38550, 16'd26600, 16'd7814, 16'd54733});
	test_expansion(128'h66c7aacadfd1733afc46bb24c18d00e4, {16'd49642, 16'd47264, 16'd14342, 16'd54999, 16'd60196, 16'd26754, 16'd34247, 16'd13116, 16'd35300, 16'd39789, 16'd64344, 16'd10713, 16'd24376, 16'd62391, 16'd49198, 16'd23150, 16'd57162, 16'd2495, 16'd42996, 16'd27588, 16'd40559, 16'd37569, 16'd26911, 16'd44310, 16'd44451, 16'd14948});
	test_expansion(128'h8253f39ae842b20eec719bb06abe2357, {16'd9146, 16'd9685, 16'd55846, 16'd27035, 16'd35633, 16'd15863, 16'd19789, 16'd20731, 16'd28516, 16'd26559, 16'd8306, 16'd40276, 16'd57089, 16'd54723, 16'd4713, 16'd25327, 16'd11265, 16'd13190, 16'd10792, 16'd63163, 16'd61099, 16'd50125, 16'd36718, 16'd14168, 16'd50902, 16'd62388});
	test_expansion(128'hdf4967816eeb95f75990a4547d834a34, {16'd22028, 16'd59106, 16'd22876, 16'd17974, 16'd9541, 16'd36317, 16'd39434, 16'd11825, 16'd34594, 16'd10255, 16'd32061, 16'd26514, 16'd10485, 16'd20757, 16'd60263, 16'd41976, 16'd28040, 16'd52548, 16'd40057, 16'd64814, 16'd1730, 16'd37758, 16'd36123, 16'd64326, 16'd14295, 16'd30258});
	test_expansion(128'hee3483143abfd1c389d846153966a686, {16'd51391, 16'd9591, 16'd46224, 16'd106, 16'd22800, 16'd63539, 16'd43087, 16'd20468, 16'd18998, 16'd9438, 16'd39886, 16'd27657, 16'd11723, 16'd65166, 16'd25681, 16'd59639, 16'd36266, 16'd13878, 16'd29754, 16'd64982, 16'd51139, 16'd35948, 16'd35178, 16'd27821, 16'd27661, 16'd43153});
	test_expansion(128'ha9b3fd8e23943e8198e1e07a95174f40, {16'd20373, 16'd9466, 16'd34507, 16'd52782, 16'd1604, 16'd62061, 16'd59307, 16'd3900, 16'd41748, 16'd29321, 16'd61498, 16'd27101, 16'd37817, 16'd27172, 16'd33731, 16'd26526, 16'd11844, 16'd30665, 16'd38931, 16'd32151, 16'd40017, 16'd11387, 16'd40565, 16'd8464, 16'd42875, 16'd37745});
	test_expansion(128'h58cc88069215217782a5eee095f17c44, {16'd28047, 16'd32436, 16'd17999, 16'd62628, 16'd33192, 16'd23431, 16'd33727, 16'd15942, 16'd53801, 16'd19163, 16'd44567, 16'd62341, 16'd14999, 16'd29453, 16'd65471, 16'd3432, 16'd62762, 16'd48145, 16'd16303, 16'd48883, 16'd27393, 16'd7301, 16'd43885, 16'd8813, 16'd26251, 16'd5278});
	test_expansion(128'h039d803d2dbfa7c2cffc2384244180ad, {16'd58618, 16'd7986, 16'd7101, 16'd48197, 16'd9442, 16'd40283, 16'd18020, 16'd43861, 16'd7077, 16'd15692, 16'd58456, 16'd21803, 16'd46415, 16'd30818, 16'd44914, 16'd35682, 16'd33279, 16'd7775, 16'd56965, 16'd57219, 16'd7037, 16'd24579, 16'd38815, 16'd55347, 16'd38132, 16'd45709});
	test_expansion(128'he6442eb6ba42dd55e90dcdd5010be864, {16'd58278, 16'd31767, 16'd29997, 16'd38420, 16'd31704, 16'd48468, 16'd55492, 16'd1202, 16'd4162, 16'd14953, 16'd28766, 16'd52738, 16'd9, 16'd10794, 16'd38084, 16'd24481, 16'd23721, 16'd33079, 16'd52531, 16'd15239, 16'd22484, 16'd18505, 16'd37112, 16'd38866, 16'd10979, 16'd53475});
	test_expansion(128'h9c820a86a1723ad099310083a940ebda, {16'd50834, 16'd43921, 16'd56112, 16'd60231, 16'd19372, 16'd44079, 16'd64872, 16'd40856, 16'd25671, 16'd41914, 16'd44719, 16'd46341, 16'd979, 16'd46990, 16'd11474, 16'd49135, 16'd53388, 16'd64983, 16'd44022, 16'd7944, 16'd49054, 16'd39280, 16'd6240, 16'd29573, 16'd58808, 16'd43226});
	test_expansion(128'h2e04158181a1fd4e0d4cb77fb2c1b1a0, {16'd57940, 16'd61094, 16'd59306, 16'd38190, 16'd50892, 16'd6853, 16'd43316, 16'd34609, 16'd2067, 16'd25613, 16'd1924, 16'd45499, 16'd38460, 16'd12370, 16'd48271, 16'd35894, 16'd53427, 16'd39199, 16'd43845, 16'd7, 16'd41745, 16'd15706, 16'd59139, 16'd11705, 16'd15624, 16'd38816});
	test_expansion(128'hd9c5bf169f7b2b26c7b65536bf73f7b2, {16'd52759, 16'd19100, 16'd27515, 16'd19466, 16'd50224, 16'd10423, 16'd56175, 16'd45262, 16'd34553, 16'd38362, 16'd49356, 16'd59001, 16'd2130, 16'd30071, 16'd47503, 16'd45957, 16'd37280, 16'd34495, 16'd45775, 16'd13882, 16'd62636, 16'd17536, 16'd3421, 16'd51193, 16'd31802, 16'd56484});
	test_expansion(128'h3620bf65c366ad4a914b17c57fe339b8, {16'd4212, 16'd37020, 16'd21065, 16'd45805, 16'd18847, 16'd52047, 16'd2605, 16'd52751, 16'd26580, 16'd35386, 16'd64325, 16'd63452, 16'd38337, 16'd61122, 16'd24904, 16'd24021, 16'd12505, 16'd29100, 16'd41041, 16'd43404, 16'd8185, 16'd38929, 16'd59972, 16'd11854, 16'd24928, 16'd11660});
	test_expansion(128'h62f0e7bade3c68e68af087844f73c1cc, {16'd57878, 16'd47054, 16'd3689, 16'd865, 16'd31858, 16'd559, 16'd46743, 16'd26241, 16'd26498, 16'd56820, 16'd51122, 16'd34667, 16'd48852, 16'd51447, 16'd18918, 16'd62832, 16'd5859, 16'd3361, 16'd29577, 16'd46227, 16'd41736, 16'd16401, 16'd47110, 16'd24701, 16'd49761, 16'd44980});
	test_expansion(128'hf127cd0c0102ff3662f0872a4d7e9332, {16'd41408, 16'd14047, 16'd35361, 16'd51718, 16'd56383, 16'd35614, 16'd59052, 16'd28465, 16'd28396, 16'd30546, 16'd26267, 16'd16779, 16'd17122, 16'd13740, 16'd7199, 16'd62577, 16'd49903, 16'd46025, 16'd12176, 16'd10151, 16'd25052, 16'd43002, 16'd8286, 16'd33102, 16'd18140, 16'd22193});
	test_expansion(128'hfc4bbcef54c13fb585da4c4bd33063b6, {16'd31175, 16'd10033, 16'd36110, 16'd1082, 16'd62975, 16'd58358, 16'd20430, 16'd57940, 16'd47015, 16'd28794, 16'd33606, 16'd29849, 16'd49279, 16'd7826, 16'd19511, 16'd60193, 16'd8090, 16'd12105, 16'd7262, 16'd33866, 16'd12045, 16'd21284, 16'd14721, 16'd46831, 16'd15688, 16'd58918});
	test_expansion(128'h7ecc7abc2e00d71fa79e4b63fc6b2599, {16'd38497, 16'd62424, 16'd1682, 16'd46909, 16'd64540, 16'd1404, 16'd24679, 16'd47662, 16'd19402, 16'd53846, 16'd11060, 16'd2566, 16'd50636, 16'd63188, 16'd6846, 16'd6251, 16'd34227, 16'd13989, 16'd13217, 16'd8138, 16'd7904, 16'd36345, 16'd14373, 16'd36629, 16'd46324, 16'd25649});
	test_expansion(128'h1b0d3535c61583943e37a6bfdd536965, {16'd30261, 16'd36886, 16'd60384, 16'd41980, 16'd27604, 16'd59695, 16'd57766, 16'd45168, 16'd54043, 16'd52571, 16'd38829, 16'd50694, 16'd53426, 16'd51713, 16'd5713, 16'd51887, 16'd4243, 16'd29768, 16'd31780, 16'd49977, 16'd28712, 16'd45572, 16'd49272, 16'd58021, 16'd12875, 16'd47748});
	test_expansion(128'h8a3bd57aa9c8988764faa00f44d9d359, {16'd52741, 16'd54874, 16'd15248, 16'd61433, 16'd22342, 16'd42255, 16'd64256, 16'd58443, 16'd24743, 16'd55211, 16'd32945, 16'd19497, 16'd16131, 16'd4632, 16'd25700, 16'd27131, 16'd20603, 16'd13072, 16'd1287, 16'd61560, 16'd40267, 16'd19028, 16'd33963, 16'd12524, 16'd26878, 16'd53578});
	test_expansion(128'hc78adc31dbef423fe6bdb1207deb3d8f, {16'd24768, 16'd29707, 16'd35892, 16'd9764, 16'd20990, 16'd52058, 16'd12411, 16'd39805, 16'd50750, 16'd5098, 16'd4425, 16'd49264, 16'd29095, 16'd21178, 16'd25990, 16'd65445, 16'd39700, 16'd16229, 16'd9058, 16'd48406, 16'd36641, 16'd56940, 16'd64795, 16'd20250, 16'd25570, 16'd7999});
	test_expansion(128'hb4f71dcb94a4c1fcf271012ee2e292eb, {16'd52539, 16'd4841, 16'd47963, 16'd15821, 16'd61710, 16'd599, 16'd52271, 16'd51909, 16'd14212, 16'd1968, 16'd29835, 16'd9021, 16'd8356, 16'd62082, 16'd25010, 16'd30823, 16'd19243, 16'd21756, 16'd41530, 16'd3605, 16'd18722, 16'd58677, 16'd42718, 16'd5978, 16'd61409, 16'd16930});
	test_expansion(128'h0733ed0ecf83355f1c6a744c41c3b452, {16'd21947, 16'd28484, 16'd14364, 16'd28498, 16'd50188, 16'd53171, 16'd33501, 16'd58167, 16'd27158, 16'd41516, 16'd25742, 16'd25834, 16'd6026, 16'd4680, 16'd61721, 16'd49672, 16'd17813, 16'd42280, 16'd49567, 16'd9231, 16'd49105, 16'd2822, 16'd46228, 16'd59222, 16'd2989, 16'd58744});
	test_expansion(128'ha8c13ea7fb869e28a9bc6ceb28189629, {16'd30509, 16'd29216, 16'd18253, 16'd848, 16'd17451, 16'd53955, 16'd17131, 16'd2473, 16'd58479, 16'd46766, 16'd10688, 16'd54020, 16'd63186, 16'd45223, 16'd17681, 16'd16046, 16'd32683, 16'd50806, 16'd37067, 16'd65293, 16'd38227, 16'd34083, 16'd9788, 16'd62846, 16'd18155, 16'd58974});
	test_expansion(128'h38c9d6ba4bc1aad1981fbd3e5f4038ee, {16'd30130, 16'd11743, 16'd13383, 16'd28939, 16'd2659, 16'd36089, 16'd6967, 16'd62949, 16'd29664, 16'd52509, 16'd1256, 16'd9690, 16'd13018, 16'd5526, 16'd25348, 16'd60357, 16'd40102, 16'd4558, 16'd28320, 16'd29840, 16'd21064, 16'd22785, 16'd58502, 16'd16205, 16'd47395, 16'd57780});
	test_expansion(128'hb4ab4f3be39300c91d78f6bd8002f2b2, {16'd33308, 16'd26469, 16'd10077, 16'd27093, 16'd28453, 16'd12918, 16'd55047, 16'd56391, 16'd50335, 16'd46572, 16'd4793, 16'd48780, 16'd15656, 16'd7190, 16'd19630, 16'd12733, 16'd26777, 16'd8089, 16'd23605, 16'd29161, 16'd9869, 16'd36236, 16'd4153, 16'd53479, 16'd57917, 16'd55503});
	test_expansion(128'heacd0f97330c4733ef615f50db945e9b, {16'd40874, 16'd25306, 16'd31051, 16'd42195, 16'd36775, 16'd20734, 16'd59260, 16'd40663, 16'd16656, 16'd23065, 16'd63238, 16'd26707, 16'd2000, 16'd20586, 16'd60110, 16'd2517, 16'd21723, 16'd7679, 16'd30354, 16'd21021, 16'd31764, 16'd43620, 16'd60137, 16'd57886, 16'd29445, 16'd62934});
	test_expansion(128'ha86da1d1a94dfb1a20663f49d68c1152, {16'd7553, 16'd5673, 16'd13549, 16'd10145, 16'd7587, 16'd47775, 16'd38626, 16'd64523, 16'd29426, 16'd38728, 16'd61150, 16'd10934, 16'd1296, 16'd53360, 16'd56966, 16'd61379, 16'd34046, 16'd49903, 16'd38892, 16'd2557, 16'd36189, 16'd13584, 16'd20401, 16'd54464, 16'd51399, 16'd14684});
	test_expansion(128'he306b3e927eaa237f768dbbcab68b3cd, {16'd48683, 16'd20871, 16'd29291, 16'd35835, 16'd7020, 16'd50617, 16'd24210, 16'd45180, 16'd4774, 16'd36578, 16'd12977, 16'd45130, 16'd59306, 16'd27690, 16'd37198, 16'd17954, 16'd42296, 16'd25498, 16'd5087, 16'd44236, 16'd54800, 16'd39571, 16'd35620, 16'd52141, 16'd40458, 16'd5271});
	test_expansion(128'hfa7f5f124cdc05ebcb1d60ce7cf1de9d, {16'd20669, 16'd37517, 16'd30661, 16'd22007, 16'd39402, 16'd57663, 16'd49024, 16'd35428, 16'd47132, 16'd38072, 16'd20913, 16'd59464, 16'd7193, 16'd57032, 16'd24372, 16'd31088, 16'd62670, 16'd11322, 16'd13767, 16'd40583, 16'd12000, 16'd56049, 16'd9514, 16'd11262, 16'd21990, 16'd58453});
	test_expansion(128'h9bb4bb4b6d5e0e7eb8f4cbdf87164716, {16'd14639, 16'd867, 16'd1119, 16'd21842, 16'd17440, 16'd27070, 16'd36286, 16'd60964, 16'd60280, 16'd42158, 16'd62677, 16'd24492, 16'd58480, 16'd56248, 16'd41738, 16'd14254, 16'd30887, 16'd10012, 16'd38872, 16'd22561, 16'd51402, 16'd32349, 16'd38539, 16'd37892, 16'd21228, 16'd64237});
	test_expansion(128'hca1b7970d335b9335cceeed184707051, {16'd18895, 16'd19349, 16'd39403, 16'd16236, 16'd3638, 16'd16084, 16'd41350, 16'd2271, 16'd759, 16'd29918, 16'd50670, 16'd15383, 16'd65280, 16'd44707, 16'd10910, 16'd23263, 16'd41608, 16'd16575, 16'd27728, 16'd31434, 16'd39182, 16'd48846, 16'd49387, 16'd47112, 16'd45929, 16'd4962});
	test_expansion(128'h65c3a3954cd8457852a495eda1ddfdb0, {16'd19383, 16'd38868, 16'd40152, 16'd56053, 16'd63707, 16'd2360, 16'd36310, 16'd58501, 16'd39920, 16'd6323, 16'd22848, 16'd9658, 16'd61704, 16'd10250, 16'd53620, 16'd52684, 16'd60526, 16'd51842, 16'd59274, 16'd6084, 16'd61797, 16'd18549, 16'd41734, 16'd13553, 16'd46207, 16'd54912});
	test_expansion(128'h44d849421ecbbf784a4cb52a085885a4, {16'd46030, 16'd43468, 16'd37630, 16'd19532, 16'd3513, 16'd2005, 16'd6730, 16'd42414, 16'd24437, 16'd34974, 16'd60550, 16'd50785, 16'd3876, 16'd6475, 16'd55052, 16'd20748, 16'd51618, 16'd29014, 16'd18868, 16'd9361, 16'd57081, 16'd32275, 16'd7065, 16'd65210, 16'd59223, 16'd38469});
	test_expansion(128'haca0d9147c1fb7aa96d8e5b999b2d1c0, {16'd35786, 16'd61814, 16'd52376, 16'd11924, 16'd39075, 16'd7375, 16'd12235, 16'd41578, 16'd39393, 16'd4777, 16'd23784, 16'd2905, 16'd42838, 16'd7435, 16'd2154, 16'd43491, 16'd8736, 16'd21057, 16'd39722, 16'd61478, 16'd61190, 16'd12106, 16'd56368, 16'd6658, 16'd9218, 16'd65});
	test_expansion(128'h00123a89fffa89ab30bc6abe712520fa, {16'd16881, 16'd63546, 16'd48666, 16'd41165, 16'd57244, 16'd43902, 16'd12505, 16'd54277, 16'd41150, 16'd56457, 16'd46530, 16'd20485, 16'd52062, 16'd9450, 16'd8331, 16'd20784, 16'd22068, 16'd16097, 16'd17141, 16'd3132, 16'd56577, 16'd10942, 16'd15823, 16'd49180, 16'd44904, 16'd34921});
	test_expansion(128'had60be0b319ccc7219d4b545c0129098, {16'd6282, 16'd25042, 16'd36033, 16'd4381, 16'd29070, 16'd26756, 16'd3250, 16'd27966, 16'd51498, 16'd42749, 16'd26178, 16'd36391, 16'd3286, 16'd64848, 16'd13704, 16'd26325, 16'd11684, 16'd32098, 16'd14094, 16'd3997, 16'd40468, 16'd34907, 16'd38875, 16'd1359, 16'd7736, 16'd52096});
	test_expansion(128'h511f35cbb82f9a444a762a882a004f30, {16'd16840, 16'd10712, 16'd4571, 16'd42413, 16'd22103, 16'd62900, 16'd64847, 16'd60342, 16'd62661, 16'd20328, 16'd38572, 16'd27038, 16'd51117, 16'd43342, 16'd40001, 16'd10154, 16'd37887, 16'd43871, 16'd43237, 16'd43204, 16'd13143, 16'd48381, 16'd11911, 16'd22031, 16'd33296, 16'd57543});
	test_expansion(128'h4dc3b2dea9ee3be0ddd42ea357083f4d, {16'd49965, 16'd33737, 16'd47070, 16'd46208, 16'd62292, 16'd45444, 16'd13750, 16'd29975, 16'd2320, 16'd34471, 16'd36061, 16'd55038, 16'd43458, 16'd48091, 16'd23480, 16'd253, 16'd37434, 16'd13750, 16'd62110, 16'd56358, 16'd34999, 16'd44495, 16'd4806, 16'd24123, 16'd28173, 16'd8732});
	test_expansion(128'h812a42b719e80f926856fa2db84e26cb, {16'd40160, 16'd16571, 16'd53215, 16'd33929, 16'd6721, 16'd22368, 16'd34080, 16'd53613, 16'd62164, 16'd29706, 16'd28025, 16'd55365, 16'd59217, 16'd1833, 16'd18269, 16'd22336, 16'd29272, 16'd59509, 16'd11974, 16'd41053, 16'd60079, 16'd25322, 16'd2690, 16'd10764, 16'd36834, 16'd5202});
	test_expansion(128'h5097742339a1af3355405fd9ecf85b26, {16'd18811, 16'd16118, 16'd17196, 16'd46234, 16'd11802, 16'd18757, 16'd6589, 16'd32272, 16'd50637, 16'd34502, 16'd19161, 16'd23922, 16'd11606, 16'd47779, 16'd63593, 16'd58034, 16'd51986, 16'd2693, 16'd29317, 16'd23596, 16'd38749, 16'd6397, 16'd12717, 16'd14366, 16'd41728, 16'd59980});
	test_expansion(128'h88b0d464bb05426d70e5bb75a9f2cf0f, {16'd64875, 16'd6878, 16'd15243, 16'd28948, 16'd58356, 16'd23670, 16'd4622, 16'd7023, 16'd51594, 16'd24584, 16'd58608, 16'd57872, 16'd26418, 16'd2937, 16'd14480, 16'd24091, 16'd4154, 16'd64428, 16'd36652, 16'd7057, 16'd45906, 16'd53192, 16'd30417, 16'd49389, 16'd22197, 16'd29225});
	test_expansion(128'hde097e9a99d06f55ad3b0745e1d005ea, {16'd36371, 16'd29485, 16'd27744, 16'd60073, 16'd65111, 16'd9104, 16'd51034, 16'd49888, 16'd1452, 16'd2574, 16'd18011, 16'd53387, 16'd27527, 16'd10721, 16'd19169, 16'd13004, 16'd27794, 16'd30827, 16'd3305, 16'd47527, 16'd44383, 16'd30363, 16'd36850, 16'd19102, 16'd52806, 16'd40145});
	test_expansion(128'hfbb1bdf0636b8eafa2bff6a7a044f3d8, {16'd19497, 16'd39679, 16'd57414, 16'd32653, 16'd18263, 16'd31897, 16'd58596, 16'd63796, 16'd13594, 16'd53510, 16'd27959, 16'd25155, 16'd56251, 16'd47313, 16'd47813, 16'd36589, 16'd34979, 16'd31448, 16'd10229, 16'd57217, 16'd26524, 16'd3950, 16'd12115, 16'd19978, 16'd16761, 16'd27235});
	test_expansion(128'h559637842c7876d4bb29c31b4cf43360, {16'd216, 16'd35056, 16'd56021, 16'd47781, 16'd51142, 16'd30621, 16'd11567, 16'd45456, 16'd57627, 16'd37784, 16'd33068, 16'd42976, 16'd64697, 16'd59067, 16'd35500, 16'd63179, 16'd54699, 16'd22332, 16'd20520, 16'd19773, 16'd33704, 16'd61188, 16'd39535, 16'd2102, 16'd37189, 16'd10069});
	test_expansion(128'hd07bdc60f0f6473c8bfcc211a5521b25, {16'd47386, 16'd19516, 16'd60842, 16'd62557, 16'd38374, 16'd55408, 16'd43322, 16'd41775, 16'd23427, 16'd16541, 16'd12003, 16'd56343, 16'd57624, 16'd10755, 16'd37284, 16'd5004, 16'd7818, 16'd54299, 16'd24958, 16'd59275, 16'd2302, 16'd38947, 16'd63996, 16'd4636, 16'd63772, 16'd37645});
	test_expansion(128'hae742376f2b904db5aaba6b37c996fdb, {16'd46418, 16'd40213, 16'd26889, 16'd23881, 16'd51700, 16'd5478, 16'd59585, 16'd34876, 16'd37610, 16'd27847, 16'd15201, 16'd19387, 16'd53017, 16'd8521, 16'd49916, 16'd45519, 16'd64495, 16'd55663, 16'd24754, 16'd26420, 16'd10407, 16'd61623, 16'd31058, 16'd48253, 16'd3383, 16'd27565});
	test_expansion(128'h12b2ce09f148ebc5c66b675ed96d871a, {16'd4182, 16'd10283, 16'd50542, 16'd25385, 16'd62851, 16'd19900, 16'd13981, 16'd45545, 16'd13713, 16'd11644, 16'd11405, 16'd2326, 16'd1428, 16'd29216, 16'd39635, 16'd11258, 16'd53610, 16'd49513, 16'd15378, 16'd29965, 16'd60129, 16'd2526, 16'd65262, 16'd18510, 16'd13782, 16'd1646});
	test_expansion(128'h6afaed42912b7a8a121196ea37d00223, {16'd61849, 16'd46229, 16'd11894, 16'd6184, 16'd19217, 16'd53293, 16'd39507, 16'd42316, 16'd10662, 16'd50374, 16'd27296, 16'd50145, 16'd23490, 16'd21640, 16'd7265, 16'd39198, 16'd42162, 16'd41184, 16'd59693, 16'd15970, 16'd48782, 16'd30805, 16'd47513, 16'd27939, 16'd7773, 16'd29485});
	test_expansion(128'hf4d5fabb76717c20fd28a91687f97763, {16'd45459, 16'd42747, 16'd19119, 16'd39505, 16'd20937, 16'd62863, 16'd12922, 16'd22058, 16'd44491, 16'd19654, 16'd38168, 16'd40583, 16'd57722, 16'd13191, 16'd4309, 16'd29311, 16'd3379, 16'd38610, 16'd40079, 16'd30713, 16'd35722, 16'd23071, 16'd28893, 16'd3325, 16'd45715, 16'd2751});
	test_expansion(128'h403653c59c0200448001df9d02c28335, {16'd51937, 16'd12152, 16'd46574, 16'd23743, 16'd34520, 16'd17718, 16'd48487, 16'd57205, 16'd12203, 16'd17661, 16'd16600, 16'd16700, 16'd27227, 16'd35976, 16'd33815, 16'd15642, 16'd15901, 16'd65025, 16'd23367, 16'd15209, 16'd40963, 16'd36694, 16'd47087, 16'd42720, 16'd19529, 16'd16019});
	test_expansion(128'h0102f920c9d9e6ff7a2a74b52f74a5ec, {16'd28532, 16'd20393, 16'd25734, 16'd42526, 16'd21019, 16'd21869, 16'd34993, 16'd29665, 16'd53558, 16'd62961, 16'd15675, 16'd24842, 16'd59434, 16'd25422, 16'd62912, 16'd24858, 16'd9976, 16'd2113, 16'd60762, 16'd51468, 16'd6570, 16'd17358, 16'd53455, 16'd18998, 16'd8109, 16'd14691});
	test_expansion(128'h2a81239d4c47df86b819c5c4289f780d, {16'd28499, 16'd2572, 16'd17910, 16'd31668, 16'd62778, 16'd43268, 16'd42248, 16'd54501, 16'd62432, 16'd22531, 16'd41683, 16'd47510, 16'd10470, 16'd47161, 16'd27332, 16'd2871, 16'd64843, 16'd27281, 16'd15536, 16'd60757, 16'd47764, 16'd62478, 16'd60424, 16'd8506, 16'd24521, 16'd61600});
	test_expansion(128'ha1b7389da83f2e3fb522cc0212709320, {16'd38207, 16'd28642, 16'd48066, 16'd17947, 16'd23012, 16'd15094, 16'd211, 16'd58338, 16'd45953, 16'd8568, 16'd12120, 16'd26345, 16'd2959, 16'd19620, 16'd13407, 16'd57509, 16'd56990, 16'd385, 16'd56220, 16'd61124, 16'd41418, 16'd45301, 16'd35121, 16'd22482, 16'd56639, 16'd55624});
	test_expansion(128'h52fee651ecd9e69ca4f9363bdf2f2931, {16'd24669, 16'd26733, 16'd60248, 16'd31627, 16'd35403, 16'd44621, 16'd40208, 16'd40520, 16'd56882, 16'd57954, 16'd58323, 16'd51428, 16'd28568, 16'd26159, 16'd4852, 16'd19472, 16'd17618, 16'd48773, 16'd1743, 16'd47760, 16'd28976, 16'd8030, 16'd21647, 16'd8041, 16'd45621, 16'd47513});
	test_expansion(128'h8e8d571a013b18e0da8ba4a5c515857b, {16'd44888, 16'd31334, 16'd64308, 16'd8298, 16'd62264, 16'd38136, 16'd18592, 16'd2441, 16'd15389, 16'd34984, 16'd16424, 16'd57162, 16'd59690, 16'd14233, 16'd37710, 16'd15590, 16'd56378, 16'd53879, 16'd51254, 16'd20946, 16'd61933, 16'd4650, 16'd63897, 16'd15003, 16'd52790, 16'd50033});
	test_expansion(128'hf5503de5f758636d448fb09d1ec81727, {16'd4009, 16'd55179, 16'd59739, 16'd3849, 16'd11623, 16'd33181, 16'd6912, 16'd23195, 16'd44368, 16'd7356, 16'd63761, 16'd8695, 16'd18999, 16'd33782, 16'd36526, 16'd41875, 16'd31534, 16'd6098, 16'd34986, 16'd9021, 16'd60922, 16'd57906, 16'd56006, 16'd24996, 16'd55872, 16'd16759});
	test_expansion(128'h49744945954121dd2fc4dc9897d2c18b, {16'd10394, 16'd53886, 16'd59836, 16'd63815, 16'd51875, 16'd6358, 16'd23928, 16'd34621, 16'd3058, 16'd25978, 16'd3089, 16'd54571, 16'd37814, 16'd31607, 16'd5263, 16'd2328, 16'd44925, 16'd28794, 16'd12319, 16'd46013, 16'd7042, 16'd61338, 16'd23882, 16'd7127, 16'd19206, 16'd1832});
	test_expansion(128'h13bd29cfddc13f5e8d5006b2398693e7, {16'd34325, 16'd53065, 16'd43611, 16'd53075, 16'd51698, 16'd27448, 16'd11602, 16'd10626, 16'd63088, 16'd65382, 16'd40003, 16'd56855, 16'd62791, 16'd5314, 16'd63087, 16'd7908, 16'd36869, 16'd11963, 16'd37581, 16'd41548, 16'd32860, 16'd7455, 16'd56134, 16'd54585, 16'd36499, 16'd32367});
	test_expansion(128'hefc24b5a6272af08792409c573c93fd9, {16'd48165, 16'd35621, 16'd25422, 16'd7963, 16'd513, 16'd64113, 16'd38396, 16'd17635, 16'd58262, 16'd64557, 16'd60595, 16'd52963, 16'd17930, 16'd37751, 16'd6904, 16'd42158, 16'd62043, 16'd5093, 16'd14662, 16'd58559, 16'd6630, 16'd61508, 16'd45403, 16'd20950, 16'd36879, 16'd32053});
	test_expansion(128'h514aecc983a593fe3361b76a6d3bb37e, {16'd57290, 16'd61124, 16'd17371, 16'd24793, 16'd39074, 16'd12252, 16'd47189, 16'd35278, 16'd60405, 16'd30924, 16'd6267, 16'd19789, 16'd63895, 16'd2294, 16'd43232, 16'd62569, 16'd23629, 16'd40236, 16'd59344, 16'd48052, 16'd1667, 16'd31465, 16'd29846, 16'd38167, 16'd6746, 16'd62844});
	test_expansion(128'h02f98ea85c32a483616b1bc97da334d5, {16'd25916, 16'd49853, 16'd17858, 16'd50253, 16'd63230, 16'd58263, 16'd53176, 16'd37674, 16'd38188, 16'd63513, 16'd52214, 16'd13588, 16'd44785, 16'd50106, 16'd2051, 16'd15415, 16'd61211, 16'd39506, 16'd53032, 16'd7363, 16'd40403, 16'd26011, 16'd48807, 16'd12706, 16'd53229, 16'd61330});
	test_expansion(128'h945c361ff929ab871eabf9bc42f95e60, {16'd54543, 16'd34951, 16'd27708, 16'd62398, 16'd49370, 16'd58554, 16'd37852, 16'd8555, 16'd61635, 16'd13814, 16'd50224, 16'd28111, 16'd29533, 16'd3335, 16'd52536, 16'd19618, 16'd52797, 16'd51940, 16'd62918, 16'd5986, 16'd59940, 16'd62616, 16'd26143, 16'd29382, 16'd11638, 16'd54278});
	test_expansion(128'h186ccb5cca232bb6a130b578be66c3bb, {16'd35333, 16'd20795, 16'd22788, 16'd14459, 16'd30991, 16'd31570, 16'd65115, 16'd61097, 16'd11758, 16'd12201, 16'd25883, 16'd22913, 16'd17300, 16'd56308, 16'd31539, 16'd19493, 16'd62743, 16'd14816, 16'd31723, 16'd24326, 16'd12899, 16'd52043, 16'd4841, 16'd18006, 16'd34380, 16'd30941});
	test_expansion(128'hc5d9f395e287a86c3f3f88a934bd9df9, {16'd46730, 16'd13748, 16'd30761, 16'd26702, 16'd40850, 16'd44610, 16'd15685, 16'd17541, 16'd40683, 16'd42054, 16'd7429, 16'd65344, 16'd51268, 16'd8985, 16'd11399, 16'd37961, 16'd33184, 16'd44612, 16'd45743, 16'd41125, 16'd64765, 16'd23331, 16'd32795, 16'd42484, 16'd40385, 16'd56350});
	test_expansion(128'hf0cf55b34cf71ef9ca1010610b273cb9, {16'd40640, 16'd1099, 16'd28128, 16'd12400, 16'd29631, 16'd44860, 16'd9608, 16'd6793, 16'd2409, 16'd57854, 16'd46016, 16'd11570, 16'd5558, 16'd20427, 16'd59556, 16'd63936, 16'd9838, 16'd39834, 16'd51719, 16'd22115, 16'd21749, 16'd8798, 16'd18239, 16'd62331, 16'd12425, 16'd49559});
	test_expansion(128'hababe2ad810b0298b58bc508ba0d08fc, {16'd35702, 16'd19162, 16'd46492, 16'd24443, 16'd4195, 16'd44832, 16'd40244, 16'd29131, 16'd25904, 16'd55274, 16'd57010, 16'd38149, 16'd22037, 16'd64355, 16'd836, 16'd8351, 16'd24840, 16'd32348, 16'd35202, 16'd64301, 16'd18303, 16'd35141, 16'd34883, 16'd63272, 16'd46356, 16'd51042});
	test_expansion(128'h5f307518bfed8dfb71685637602940b7, {16'd53803, 16'd46762, 16'd62000, 16'd64377, 16'd21043, 16'd57184, 16'd43278, 16'd46726, 16'd9612, 16'd10352, 16'd52697, 16'd9218, 16'd17198, 16'd43074, 16'd61640, 16'd52134, 16'd16685, 16'd63314, 16'd44426, 16'd23432, 16'd19894, 16'd7035, 16'd33893, 16'd24946, 16'd48072, 16'd20531});
	test_expansion(128'hbfde7951ee5352ea6cdf0b32a57ddf65, {16'd42790, 16'd35921, 16'd13415, 16'd41353, 16'd31101, 16'd8795, 16'd54704, 16'd8419, 16'd3345, 16'd30149, 16'd29940, 16'd17343, 16'd51419, 16'd38424, 16'd26576, 16'd20401, 16'd28987, 16'd63913, 16'd44652, 16'd17655, 16'd19996, 16'd59744, 16'd47042, 16'd43432, 16'd34619, 16'd23545});
	test_expansion(128'h5beb4b4a8de2dc7c5c323d63ae516389, {16'd54422, 16'd1068, 16'd9564, 16'd52752, 16'd25667, 16'd44941, 16'd33933, 16'd25816, 16'd26778, 16'd37303, 16'd28730, 16'd47326, 16'd64056, 16'd12724, 16'd13663, 16'd7285, 16'd31137, 16'd39690, 16'd44608, 16'd19742, 16'd64050, 16'd40740, 16'd38168, 16'd12761, 16'd37352, 16'd52194});
	test_expansion(128'hf72e43d1bdd1bfa412d2d18e7923c8e0, {16'd32504, 16'd55416, 16'd840, 16'd2200, 16'd36065, 16'd9969, 16'd64674, 16'd34749, 16'd54161, 16'd19554, 16'd44189, 16'd28416, 16'd43402, 16'd34542, 16'd60701, 16'd58021, 16'd23580, 16'd64369, 16'd47438, 16'd42557, 16'd15094, 16'd808, 16'd7711, 16'd42869, 16'd29454, 16'd4142});
	test_expansion(128'h3684a496203aabcfdff5cedba0913c5e, {16'd22417, 16'd8103, 16'd57013, 16'd64401, 16'd217, 16'd35676, 16'd31957, 16'd43200, 16'd36531, 16'd815, 16'd65186, 16'd64976, 16'd47002, 16'd30689, 16'd9951, 16'd32582, 16'd5769, 16'd45373, 16'd11175, 16'd28227, 16'd15351, 16'd12510, 16'd21621, 16'd4108, 16'd51896, 16'd6751});
	test_expansion(128'hd17c602bc195ccbc87b0c6a1213c1b04, {16'd11554, 16'd28788, 16'd10470, 16'd11873, 16'd32375, 16'd53362, 16'd43093, 16'd54117, 16'd57412, 16'd25057, 16'd16853, 16'd36547, 16'd52360, 16'd60102, 16'd36982, 16'd12909, 16'd35433, 16'd58861, 16'd57734, 16'd38286, 16'd48281, 16'd10695, 16'd25858, 16'd124, 16'd62604, 16'd20367});
	test_expansion(128'hf263f1c69ac8f6f9e67a610331bbe8ec, {16'd5649, 16'd24525, 16'd41255, 16'd48277, 16'd42105, 16'd2323, 16'd34325, 16'd32954, 16'd41939, 16'd41729, 16'd34019, 16'd1015, 16'd44522, 16'd44555, 16'd30830, 16'd5112, 16'd47835, 16'd53034, 16'd14335, 16'd2288, 16'd3341, 16'd25493, 16'd7320, 16'd21050, 16'd57197, 16'd47050});
	test_expansion(128'h7ec925717ba359ec944ef2dbab88d495, {16'd2392, 16'd12014, 16'd10444, 16'd30062, 16'd10800, 16'd3471, 16'd15845, 16'd14185, 16'd39958, 16'd23027, 16'd19461, 16'd56084, 16'd17226, 16'd11459, 16'd64310, 16'd54862, 16'd41250, 16'd2750, 16'd46911, 16'd30997, 16'd33079, 16'd28862, 16'd44153, 16'd52894, 16'd23824, 16'd42477});
	test_expansion(128'h7d708e3288fc45cfbbd432935d1745d5, {16'd46652, 16'd2130, 16'd7813, 16'd40298, 16'd34263, 16'd50783, 16'd32805, 16'd5690, 16'd38730, 16'd34619, 16'd5712, 16'd567, 16'd51933, 16'd40952, 16'd26594, 16'd49308, 16'd19127, 16'd35035, 16'd44041, 16'd32816, 16'd45131, 16'd26084, 16'd58817, 16'd1484, 16'd27800, 16'd29842});
	test_expansion(128'hcfc578d2bb0ff829e0aecc6bcf1a9abe, {16'd11819, 16'd9375, 16'd52525, 16'd52512, 16'd10749, 16'd64485, 16'd36375, 16'd4836, 16'd19049, 16'd50907, 16'd54604, 16'd45159, 16'd5947, 16'd32666, 16'd13867, 16'd46368, 16'd64459, 16'd63921, 16'd10681, 16'd21974, 16'd24735, 16'd34173, 16'd56011, 16'd7903, 16'd7449, 16'd63885});
	test_expansion(128'hf984fc9a6cfbfcf85bc812d1945b04f0, {16'd18168, 16'd10350, 16'd53618, 16'd19829, 16'd60695, 16'd53866, 16'd63629, 16'd40331, 16'd17307, 16'd19260, 16'd46957, 16'd14518, 16'd21332, 16'd35469, 16'd9262, 16'd63037, 16'd54918, 16'd14332, 16'd19714, 16'd20595, 16'd34485, 16'd2176, 16'd18738, 16'd51685, 16'd58382, 16'd46255});
	test_expansion(128'h3f8849a201c93476a1969834f4ecb03f, {16'd11746, 16'd34970, 16'd44864, 16'd35628, 16'd48470, 16'd4556, 16'd42129, 16'd41833, 16'd33839, 16'd8646, 16'd56451, 16'd39364, 16'd55484, 16'd15800, 16'd50776, 16'd17768, 16'd65039, 16'd45123, 16'd25644, 16'd35219, 16'd23473, 16'd48059, 16'd41903, 16'd41404, 16'd63222, 16'd61865});
	test_expansion(128'h63f450d0ae3c7021287d7a4dee5c69b0, {16'd1387, 16'd25146, 16'd2083, 16'd44780, 16'd17578, 16'd56779, 16'd3784, 16'd12360, 16'd46097, 16'd46533, 16'd4710, 16'd1007, 16'd9992, 16'd56247, 16'd19255, 16'd60238, 16'd64423, 16'd9335, 16'd6338, 16'd64434, 16'd4385, 16'd61411, 16'd44597, 16'd38482, 16'd25721, 16'd5441});
	test_expansion(128'h8e28ddce5a589303b2d8c4b8b4c6333e, {16'd1740, 16'd17510, 16'd48313, 16'd63755, 16'd9787, 16'd41143, 16'd19769, 16'd19924, 16'd8351, 16'd64533, 16'd39766, 16'd49678, 16'd20415, 16'd3699, 16'd9899, 16'd15645, 16'd40450, 16'd55399, 16'd15316, 16'd36861, 16'd43032, 16'd48231, 16'd57242, 16'd50542, 16'd43167, 16'd51577});
	test_expansion(128'hdddb560e75c7f6afd8e5b45e85b19d3a, {16'd1373, 16'd42538, 16'd21767, 16'd26265, 16'd59530, 16'd32059, 16'd25248, 16'd24160, 16'd54725, 16'd404, 16'd56241, 16'd18006, 16'd24046, 16'd44872, 16'd5327, 16'd22195, 16'd5871, 16'd3243, 16'd20604, 16'd27639, 16'd3003, 16'd39688, 16'd5962, 16'd55272, 16'd55805, 16'd12680});
	test_expansion(128'h79bfdea97baea32b25a7f225e2bd8a0d, {16'd11792, 16'd21896, 16'd29672, 16'd16992, 16'd43849, 16'd54609, 16'd55867, 16'd16298, 16'd6658, 16'd41312, 16'd40982, 16'd45549, 16'd49544, 16'd24916, 16'd2733, 16'd63406, 16'd24378, 16'd4741, 16'd23496, 16'd51040, 16'd48041, 16'd42443, 16'd54496, 16'd46558, 16'd22930, 16'd43740});
	test_expansion(128'h59bd3ad16a7bc63f1362f74c87b48804, {16'd47416, 16'd18349, 16'd42783, 16'd42054, 16'd51999, 16'd5501, 16'd45863, 16'd35972, 16'd2378, 16'd13867, 16'd10364, 16'd22771, 16'd8278, 16'd33756, 16'd27706, 16'd12503, 16'd10082, 16'd43804, 16'd7211, 16'd47152, 16'd48845, 16'd52915, 16'd59830, 16'd29176, 16'd8043, 16'd14122});
	test_expansion(128'h6e653bb6bbf41c3ffb25073141f6bc9a, {16'd35451, 16'd39603, 16'd41968, 16'd28893, 16'd64430, 16'd23919, 16'd24290, 16'd52689, 16'd14268, 16'd33077, 16'd23007, 16'd29693, 16'd5696, 16'd19001, 16'd527, 16'd14198, 16'd16299, 16'd27551, 16'd35854, 16'd35595, 16'd4797, 16'd53143, 16'd24182, 16'd51938, 16'd55302, 16'd52617});
	test_expansion(128'h16980ae0391538da97cd590b167df520, {16'd53432, 16'd59955, 16'd22136, 16'd40339, 16'd11536, 16'd29551, 16'd505, 16'd26830, 16'd11234, 16'd1102, 16'd14717, 16'd34061, 16'd36429, 16'd30417, 16'd31291, 16'd62567, 16'd40259, 16'd54282, 16'd13471, 16'd6022, 16'd21768, 16'd51057, 16'd25650, 16'd34832, 16'd17764, 16'd25118});
	test_expansion(128'h1875abc44da946de9f87b21e17b09d1d, {16'd3184, 16'd39988, 16'd6954, 16'd63324, 16'd40057, 16'd60721, 16'd1884, 16'd4817, 16'd53700, 16'd17341, 16'd59851, 16'd13364, 16'd14463, 16'd46571, 16'd55841, 16'd37477, 16'd12830, 16'd14336, 16'd61989, 16'd56768, 16'd10082, 16'd61676, 16'd43387, 16'd19062, 16'd62361, 16'd54052});
	test_expansion(128'h4e97c451b93fb5f3e37a8952074bc00d, {16'd13020, 16'd6645, 16'd30026, 16'd1260, 16'd61187, 16'd34571, 16'd49836, 16'd63473, 16'd43422, 16'd33294, 16'd40028, 16'd50749, 16'd18421, 16'd11218, 16'd8394, 16'd28294, 16'd27354, 16'd51011, 16'd11622, 16'd2953, 16'd61016, 16'd12683, 16'd14198, 16'd4848, 16'd56924, 16'd38469});
	test_expansion(128'hf8fc1731ed87e9771a0fb8346425497a, {16'd19342, 16'd25866, 16'd2271, 16'd37397, 16'd42890, 16'd52096, 16'd34809, 16'd47890, 16'd38265, 16'd31167, 16'd17419, 16'd14604, 16'd34528, 16'd56174, 16'd8765, 16'd59878, 16'd40633, 16'd11566, 16'd15281, 16'd59934, 16'd45068, 16'd25510, 16'd29663, 16'd910, 16'd11796, 16'd16916});
	test_expansion(128'h96b019d89991b3507f0535cbc29b4449, {16'd33238, 16'd18070, 16'd27667, 16'd50064, 16'd24260, 16'd22619, 16'd25844, 16'd31564, 16'd3525, 16'd42254, 16'd57295, 16'd21315, 16'd4655, 16'd11128, 16'd62754, 16'd11923, 16'd64469, 16'd12458, 16'd11496, 16'd39851, 16'd6345, 16'd46891, 16'd10914, 16'd353, 16'd5394, 16'd6762});
	test_expansion(128'h4d7bbaba3c275242eaaf55765cef96d2, {16'd5198, 16'd19292, 16'd49892, 16'd51125, 16'd16179, 16'd52999, 16'd19223, 16'd22608, 16'd48331, 16'd25721, 16'd52948, 16'd44076, 16'd61771, 16'd57325, 16'd5866, 16'd52893, 16'd27376, 16'd53623, 16'd35119, 16'd28154, 16'd24806, 16'd30477, 16'd53028, 16'd30533, 16'd46732, 16'd55771});
	test_expansion(128'h0155d7d6046c6c05ddc465981bd647a9, {16'd63762, 16'd43775, 16'd46923, 16'd31086, 16'd38303, 16'd60632, 16'd44599, 16'd46670, 16'd1434, 16'd29931, 16'd1278, 16'd42192, 16'd44800, 16'd8588, 16'd27750, 16'd8137, 16'd46654, 16'd31931, 16'd59141, 16'd44252, 16'd37178, 16'd53867, 16'd10824, 16'd19623, 16'd22425, 16'd12877});
	test_expansion(128'h76f1a97d8cf158eff45fc73e88bdce5e, {16'd32832, 16'd22318, 16'd29228, 16'd21983, 16'd7709, 16'd670, 16'd37834, 16'd4208, 16'd60545, 16'd5660, 16'd53553, 16'd47020, 16'd52382, 16'd5335, 16'd25700, 16'd37115, 16'd7346, 16'd25870, 16'd14240, 16'd35030, 16'd47334, 16'd569, 16'd53799, 16'd9393, 16'd25098, 16'd36804});
	test_expansion(128'hab9aef62c3e9baa611b46678ab9dd152, {16'd33362, 16'd44836, 16'd599, 16'd27383, 16'd11504, 16'd3390, 16'd2728, 16'd13963, 16'd50896, 16'd40991, 16'd18745, 16'd33506, 16'd16700, 16'd23931, 16'd23113, 16'd24682, 16'd24697, 16'd41716, 16'd60738, 16'd7659, 16'd8055, 16'd7937, 16'd14932, 16'd16421, 16'd25152, 16'd33234});
	test_expansion(128'h772ace9b8a00fd93cfbda25291c708af, {16'd64019, 16'd64868, 16'd14554, 16'd10984, 16'd16154, 16'd17191, 16'd65203, 16'd7204, 16'd4394, 16'd37872, 16'd49803, 16'd37134, 16'd34468, 16'd60591, 16'd55671, 16'd34703, 16'd2387, 16'd29195, 16'd34499, 16'd12445, 16'd10520, 16'd43312, 16'd1922, 16'd12867, 16'd10735, 16'd40316});
	test_expansion(128'hc9b2d45edaa5ca092acc8948b6a8b8c9, {16'd5105, 16'd55260, 16'd24883, 16'd63168, 16'd24296, 16'd31004, 16'd3778, 16'd29281, 16'd62242, 16'd56127, 16'd57750, 16'd38802, 16'd1427, 16'd55877, 16'd29308, 16'd35049, 16'd2681, 16'd33089, 16'd33526, 16'd37351, 16'd59149, 16'd17099, 16'd39835, 16'd57033, 16'd25956, 16'd5239});
	test_expansion(128'h80bd2cd332133df0889ae43ed556e8d0, {16'd35411, 16'd21023, 16'd10836, 16'd38726, 16'd35963, 16'd20414, 16'd3337, 16'd54844, 16'd58566, 16'd9040, 16'd1496, 16'd19798, 16'd4345, 16'd56089, 16'd7950, 16'd26373, 16'd54967, 16'd57537, 16'd41369, 16'd30770, 16'd28458, 16'd44615, 16'd13813, 16'd27370, 16'd43875, 16'd23794});
	test_expansion(128'hffbaa8135783c965dc990bf6bc43d7f2, {16'd24065, 16'd6213, 16'd47757, 16'd45395, 16'd9474, 16'd15544, 16'd53622, 16'd62832, 16'd29257, 16'd56475, 16'd46923, 16'd64301, 16'd25876, 16'd49139, 16'd44017, 16'd23345, 16'd25049, 16'd14081, 16'd49203, 16'd63603, 16'd27144, 16'd57375, 16'd13919, 16'd46808, 16'd34565, 16'd15351});
	test_expansion(128'h9d0f2910d47ec83029e2d4eb7dacd105, {16'd63846, 16'd3299, 16'd33995, 16'd3026, 16'd49001, 16'd43804, 16'd14350, 16'd17039, 16'd41680, 16'd16398, 16'd38466, 16'd3998, 16'd15338, 16'd20298, 16'd10315, 16'd31945, 16'd42181, 16'd8840, 16'd61548, 16'd29110, 16'd14993, 16'd16619, 16'd49529, 16'd30817, 16'd1911, 16'd48414});
	test_expansion(128'ha2ab16d724a2b347e89f77c328e71bd4, {16'd49927, 16'd48945, 16'd37774, 16'd31959, 16'd57202, 16'd14990, 16'd22096, 16'd11607, 16'd1975, 16'd5315, 16'd40108, 16'd4342, 16'd61245, 16'd2070, 16'd34420, 16'd7507, 16'd33334, 16'd29746, 16'd8203, 16'd48988, 16'd51164, 16'd33617, 16'd26018, 16'd692, 16'd48577, 16'd3998});
	test_expansion(128'h0914521072bd272dfcf0d9602a12ea88, {16'd13285, 16'd61501, 16'd55126, 16'd38249, 16'd22638, 16'd21058, 16'd63738, 16'd22687, 16'd42002, 16'd55940, 16'd39773, 16'd55410, 16'd15017, 16'd64290, 16'd47804, 16'd58389, 16'd9632, 16'd54035, 16'd37966, 16'd42723, 16'd58652, 16'd8684, 16'd62132, 16'd52491, 16'd63922, 16'd7428});
	test_expansion(128'hf171ea6cbc3551f40d893f177101b08e, {16'd3380, 16'd36260, 16'd8927, 16'd47800, 16'd59352, 16'd15132, 16'd31767, 16'd15490, 16'd21036, 16'd33823, 16'd55726, 16'd42049, 16'd49831, 16'd50096, 16'd26045, 16'd21902, 16'd25958, 16'd27870, 16'd62722, 16'd15358, 16'd34344, 16'd44075, 16'd10531, 16'd47792, 16'd62659, 16'd37530});
	test_expansion(128'h6da2fee14afdc96f1e4cb75c58990f25, {16'd40826, 16'd22987, 16'd5465, 16'd59491, 16'd51387, 16'd16903, 16'd63475, 16'd47127, 16'd6018, 16'd37611, 16'd20671, 16'd26730, 16'd28395, 16'd6482, 16'd12091, 16'd57402, 16'd2929, 16'd17110, 16'd37224, 16'd8839, 16'd8159, 16'd2068, 16'd2757, 16'd32188, 16'd3206, 16'd26612});
	test_expansion(128'h15ef833210833469a336950ffb88b87f, {16'd15891, 16'd11595, 16'd62887, 16'd36974, 16'd41856, 16'd8167, 16'd61411, 16'd38982, 16'd14934, 16'd24132, 16'd58406, 16'd41785, 16'd46020, 16'd61078, 16'd42373, 16'd43122, 16'd61786, 16'd44606, 16'd49591, 16'd11637, 16'd34646, 16'd30859, 16'd55381, 16'd45818, 16'd18292, 16'd48952});
	test_expansion(128'h506c8ffd2fba9f05424d21ee3c3a0544, {16'd63924, 16'd50254, 16'd58375, 16'd51628, 16'd29837, 16'd14502, 16'd33744, 16'd46133, 16'd25965, 16'd46935, 16'd55773, 16'd1099, 16'd43723, 16'd20999, 16'd22066, 16'd14225, 16'd8139, 16'd58770, 16'd53183, 16'd22796, 16'd1292, 16'd56186, 16'd10566, 16'd35815, 16'd12915, 16'd58245});
	test_expansion(128'h4b9a12f7ea667379d0aab0cdd0faa8ee, {16'd28205, 16'd60534, 16'd37463, 16'd33483, 16'd63153, 16'd14905, 16'd633, 16'd6494, 16'd46663, 16'd22242, 16'd40368, 16'd14062, 16'd7647, 16'd26383, 16'd33048, 16'd26860, 16'd11795, 16'd32398, 16'd38639, 16'd27700, 16'd15148, 16'd23004, 16'd11317, 16'd49241, 16'd15480, 16'd48628});
	test_expansion(128'he7e929af0c8170d3c33ed20ce3a264f7, {16'd38743, 16'd46687, 16'd25524, 16'd51416, 16'd7309, 16'd19407, 16'd41939, 16'd34354, 16'd44794, 16'd5915, 16'd55465, 16'd36522, 16'd35490, 16'd46983, 16'd39413, 16'd45502, 16'd61702, 16'd19607, 16'd35435, 16'd44515, 16'd5880, 16'd39356, 16'd4971, 16'd62080, 16'd57271, 16'd7837});
	test_expansion(128'h507b6f051f6c916c25b0db4f80a1db06, {16'd13879, 16'd32844, 16'd21246, 16'd32474, 16'd64867, 16'd30232, 16'd58135, 16'd3201, 16'd51333, 16'd8360, 16'd50112, 16'd36425, 16'd34559, 16'd4415, 16'd20961, 16'd19233, 16'd35816, 16'd5042, 16'd19576, 16'd6677, 16'd17247, 16'd49415, 16'd47494, 16'd7319, 16'd39495, 16'd37454});
	test_expansion(128'h498acbc4c2c9f0fc78bd8b9159f53388, {16'd21038, 16'd16428, 16'd34431, 16'd55935, 16'd6101, 16'd34278, 16'd58324, 16'd61004, 16'd42601, 16'd56616, 16'd13107, 16'd35635, 16'd28178, 16'd1361, 16'd19754, 16'd29403, 16'd29543, 16'd54645, 16'd56351, 16'd10961, 16'd23957, 16'd41280, 16'd38734, 16'd35659, 16'd35812, 16'd20566});
	test_expansion(128'h7631993ad2b7f94e3868858bd378d1d2, {16'd7037, 16'd61098, 16'd14453, 16'd3909, 16'd21313, 16'd27778, 16'd39839, 16'd11019, 16'd27252, 16'd25377, 16'd48778, 16'd35539, 16'd30405, 16'd43305, 16'd41039, 16'd59505, 16'd44016, 16'd34128, 16'd59304, 16'd56657, 16'd64052, 16'd30046, 16'd15219, 16'd58561, 16'd37673, 16'd35131});
	test_expansion(128'hf005f72ea74d031940ea60354174042a, {16'd5482, 16'd59926, 16'd9134, 16'd14395, 16'd11335, 16'd58908, 16'd34057, 16'd27890, 16'd35898, 16'd60732, 16'd26275, 16'd884, 16'd29009, 16'd42967, 16'd51528, 16'd56469, 16'd2535, 16'd52936, 16'd21895, 16'd48221, 16'd23379, 16'd45562, 16'd888, 16'd40832, 16'd50360, 16'd16300});
	test_expansion(128'h3998048ddf00f9a37047171fd94af19f, {16'd64990, 16'd6738, 16'd18305, 16'd12680, 16'd46360, 16'd32673, 16'd4779, 16'd21276, 16'd21668, 16'd17342, 16'd17161, 16'd38554, 16'd3867, 16'd56512, 16'd37539, 16'd28812, 16'd1515, 16'd15436, 16'd37736, 16'd53881, 16'd45805, 16'd63682, 16'd4595, 16'd35863, 16'd59415, 16'd45597});
	test_expansion(128'he02b2961d860177d656fe049720b53fa, {16'd58470, 16'd65366, 16'd32083, 16'd28838, 16'd59518, 16'd33326, 16'd32209, 16'd59113, 16'd49523, 16'd33064, 16'd15466, 16'd10272, 16'd982, 16'd11027, 16'd979, 16'd54564, 16'd1658, 16'd34901, 16'd2685, 16'd8792, 16'd59034, 16'd2092, 16'd11090, 16'd30044, 16'd3412, 16'd61937});
	test_expansion(128'h7b9969e7ecbacf3a2b9cd732a382b488, {16'd45451, 16'd44816, 16'd662, 16'd5678, 16'd12276, 16'd36415, 16'd62711, 16'd29391, 16'd5922, 16'd40690, 16'd30062, 16'd62471, 16'd18714, 16'd34745, 16'd9388, 16'd52923, 16'd38272, 16'd19258, 16'd31174, 16'd33809, 16'd3682, 16'd1529, 16'd54762, 16'd50550, 16'd36971, 16'd965});
	test_expansion(128'h0acd363afb86e88633db7c0299fad68d, {16'd24741, 16'd25615, 16'd46055, 16'd34711, 16'd32784, 16'd40877, 16'd50712, 16'd13231, 16'd7412, 16'd60175, 16'd18646, 16'd15086, 16'd22137, 16'd6660, 16'd48809, 16'd18797, 16'd52317, 16'd49765, 16'd24222, 16'd5757, 16'd32546, 16'd20204, 16'd12549, 16'd50594, 16'd64531, 16'd4828});
	test_expansion(128'h7e60489f9e1d356d74470739b26948d9, {16'd20021, 16'd15765, 16'd38466, 16'd21176, 16'd39015, 16'd31584, 16'd52096, 16'd10344, 16'd63881, 16'd12081, 16'd55094, 16'd25858, 16'd53919, 16'd15599, 16'd28865, 16'd52299, 16'd51327, 16'd57095, 16'd11411, 16'd31833, 16'd780, 16'd20041, 16'd22482, 16'd6485, 16'd25136, 16'd2835});
	test_expansion(128'h235f6402ed004e06cacfa554d515497f, {16'd26856, 16'd53369, 16'd40758, 16'd5699, 16'd31685, 16'd36934, 16'd1542, 16'd2404, 16'd34988, 16'd53676, 16'd53582, 16'd17415, 16'd51934, 16'd43578, 16'd64405, 16'd11148, 16'd5690, 16'd33229, 16'd3970, 16'd7496, 16'd4986, 16'd53451, 16'd16636, 16'd59814, 16'd59398, 16'd25377});
	test_expansion(128'h7c94fc02ee0dba141a9283f91a9414ad, {16'd8091, 16'd42542, 16'd39673, 16'd48422, 16'd25332, 16'd34048, 16'd35072, 16'd2930, 16'd11068, 16'd16330, 16'd11446, 16'd22688, 16'd62804, 16'd53279, 16'd23249, 16'd23591, 16'd43712, 16'd17411, 16'd43224, 16'd2159, 16'd15318, 16'd28056, 16'd37463, 16'd49774, 16'd7588, 16'd30246});
	test_expansion(128'h6d387f15c1ab0a0c9acb12e6ebb25cd0, {16'd28324, 16'd26597, 16'd25156, 16'd53470, 16'd35981, 16'd62494, 16'd58292, 16'd16495, 16'd47474, 16'd52637, 16'd32952, 16'd4667, 16'd9822, 16'd57220, 16'd28273, 16'd6292, 16'd7801, 16'd13512, 16'd42230, 16'd11779, 16'd9118, 16'd6910, 16'd33420, 16'd36078, 16'd25899, 16'd30294});
	test_expansion(128'h55e28df1857c573dc31e956263678c40, {16'd5859, 16'd26457, 16'd62084, 16'd43566, 16'd58217, 16'd51054, 16'd9776, 16'd32557, 16'd55415, 16'd13877, 16'd40061, 16'd49738, 16'd51652, 16'd10492, 16'd25040, 16'd32549, 16'd23926, 16'd23516, 16'd32600, 16'd57839, 16'd16815, 16'd41789, 16'd23690, 16'd30708, 16'd26364, 16'd2432});
	test_expansion(128'hf193cd4d4163ab5a76b926fe9e34a67d, {16'd34471, 16'd33229, 16'd3345, 16'd13340, 16'd31915, 16'd50962, 16'd43799, 16'd1553, 16'd28871, 16'd24397, 16'd60441, 16'd18456, 16'd10159, 16'd58065, 16'd46698, 16'd16785, 16'd9768, 16'd47242, 16'd25622, 16'd5398, 16'd21221, 16'd9166, 16'd53319, 16'd48758, 16'd26520, 16'd47579});
	test_expansion(128'h1171d5ee198641c3678bfe20e04d13ba, {16'd48369, 16'd29978, 16'd5618, 16'd61905, 16'd15637, 16'd26903, 16'd13655, 16'd14071, 16'd9366, 16'd23446, 16'd4486, 16'd55747, 16'd50328, 16'd37156, 16'd48217, 16'd4254, 16'd16680, 16'd13802, 16'd53759, 16'd51573, 16'd47370, 16'd26537, 16'd35183, 16'd32802, 16'd63281, 16'd18419});
	test_expansion(128'h87456dba8e4b0eacd2d786b69a663711, {16'd56032, 16'd49524, 16'd43776, 16'd14588, 16'd28143, 16'd61381, 16'd10615, 16'd30735, 16'd58546, 16'd51033, 16'd4336, 16'd48034, 16'd6179, 16'd34032, 16'd51441, 16'd60620, 16'd18875, 16'd15858, 16'd12874, 16'd23575, 16'd6532, 16'd52294, 16'd33439, 16'd48184, 16'd35736, 16'd5356});
	test_expansion(128'h140982f3669248ec6e4920426bfe0fd5, {16'd47697, 16'd6877, 16'd42428, 16'd48156, 16'd51627, 16'd22525, 16'd53936, 16'd43146, 16'd32945, 16'd7134, 16'd1532, 16'd34810, 16'd17231, 16'd27456, 16'd24844, 16'd1991, 16'd47698, 16'd31751, 16'd1976, 16'd44883, 16'd38381, 16'd28305, 16'd11133, 16'd12375, 16'd63020, 16'd51192});
	test_expansion(128'h2b9f3db8892bbf21c5b4177650075a19, {16'd53618, 16'd12695, 16'd42383, 16'd27931, 16'd47998, 16'd62201, 16'd50844, 16'd33348, 16'd7878, 16'd3962, 16'd62497, 16'd31378, 16'd56041, 16'd15372, 16'd36072, 16'd29942, 16'd18065, 16'd16424, 16'd25172, 16'd11499, 16'd46163, 16'd36561, 16'd4221, 16'd12337, 16'd889, 16'd55849});
	test_expansion(128'h76984297ce3b7a7e6bae32f9ef117773, {16'd13422, 16'd4669, 16'd4635, 16'd24049, 16'd39116, 16'd52916, 16'd24563, 16'd4884, 16'd549, 16'd59701, 16'd14490, 16'd17724, 16'd6180, 16'd64204, 16'd60871, 16'd2621, 16'd44677, 16'd20211, 16'd41428, 16'd34881, 16'd15313, 16'd13870, 16'd40691, 16'd5382, 16'd44783, 16'd42300});
	test_expansion(128'h275ae8d5b2539f846c39f656fea9f22b, {16'd31031, 16'd16931, 16'd32742, 16'd40672, 16'd59801, 16'd46859, 16'd45232, 16'd35995, 16'd32659, 16'd26466, 16'd9880, 16'd49093, 16'd5808, 16'd42420, 16'd23933, 16'd13133, 16'd2338, 16'd63717, 16'd34576, 16'd3583, 16'd23529, 16'd2598, 16'd34048, 16'd15862, 16'd49397, 16'd16922});
	test_expansion(128'he0fe55b9beaae6e871e0c490c065c1ea, {16'd48977, 16'd14807, 16'd55358, 16'd62222, 16'd47269, 16'd18654, 16'd18054, 16'd57167, 16'd27652, 16'd40960, 16'd58799, 16'd8475, 16'd33113, 16'd59334, 16'd28835, 16'd34693, 16'd14428, 16'd53466, 16'd56648, 16'd35371, 16'd44327, 16'd62657, 16'd52422, 16'd9021, 16'd16920, 16'd26619});
	test_expansion(128'h245bb2e7561d100a166f93c815caa45a, {16'd57751, 16'd5743, 16'd9756, 16'd20637, 16'd44983, 16'd1625, 16'd56706, 16'd26762, 16'd43860, 16'd29309, 16'd41858, 16'd40170, 16'd7641, 16'd19377, 16'd28889, 16'd54135, 16'd38440, 16'd15286, 16'd12622, 16'd18351, 16'd35687, 16'd45435, 16'd65071, 16'd48988, 16'd36386, 16'd9078});
	test_expansion(128'h54162e732688e5f8616f7753fa4863b1, {16'd55862, 16'd3893, 16'd50044, 16'd63522, 16'd4658, 16'd65237, 16'd37575, 16'd55320, 16'd14386, 16'd60587, 16'd59736, 16'd25583, 16'd42855, 16'd50593, 16'd42158, 16'd19657, 16'd48506, 16'd35100, 16'd25722, 16'd54891, 16'd13483, 16'd39290, 16'd43348, 16'd47762, 16'd16897, 16'd58935});
	test_expansion(128'h4fc8dfabbe414ce56a743e35288af05e, {16'd41143, 16'd64240, 16'd46351, 16'd38406, 16'd38776, 16'd34803, 16'd56896, 16'd48943, 16'd46604, 16'd62197, 16'd54552, 16'd15755, 16'd25427, 16'd63148, 16'd22083, 16'd34630, 16'd36209, 16'd44528, 16'd2953, 16'd64049, 16'd59703, 16'd40839, 16'd56294, 16'd60825, 16'd14146, 16'd37908});
	test_expansion(128'h1374a34c1f0fcdb7a591fd2c8f603d54, {16'd41384, 16'd54341, 16'd42589, 16'd61689, 16'd13808, 16'd48294, 16'd39832, 16'd24118, 16'd5473, 16'd39009, 16'd25862, 16'd10527, 16'd54915, 16'd52784, 16'd21268, 16'd60431, 16'd59021, 16'd44382, 16'd19717, 16'd39602, 16'd58479, 16'd8601, 16'd29913, 16'd42096, 16'd55455, 16'd38895});
	test_expansion(128'h91757833a3643d323c5540f66c395b77, {16'd31009, 16'd35505, 16'd40846, 16'd3834, 16'd190, 16'd30038, 16'd18600, 16'd29057, 16'd18461, 16'd56502, 16'd12829, 16'd64694, 16'd11398, 16'd55262, 16'd22302, 16'd32620, 16'd34701, 16'd5528, 16'd2374, 16'd32511, 16'd55219, 16'd36548, 16'd42617, 16'd29110, 16'd37413, 16'd16734});
	test_expansion(128'hd54b9f78ce45e719b73d6da4c0003b08, {16'd34395, 16'd500, 16'd15897, 16'd41500, 16'd14073, 16'd37020, 16'd29039, 16'd22479, 16'd15309, 16'd18816, 16'd50145, 16'd37368, 16'd11672, 16'd48689, 16'd33059, 16'd47094, 16'd15418, 16'd53783, 16'd1399, 16'd59202, 16'd41271, 16'd26382, 16'd63407, 16'd34771, 16'd57683, 16'd34293});
	test_expansion(128'h6500b870ab6d02acccdcff853e57e830, {16'd5187, 16'd37794, 16'd32276, 16'd24488, 16'd25963, 16'd8307, 16'd38685, 16'd18429, 16'd39800, 16'd34134, 16'd8999, 16'd26163, 16'd13047, 16'd16500, 16'd4546, 16'd53213, 16'd2645, 16'd29542, 16'd2949, 16'd38919, 16'd42879, 16'd5861, 16'd38670, 16'd50528, 16'd51628, 16'd36911});
	test_expansion(128'h5efe1965a09c525c1afbda05feb96cb2, {16'd37388, 16'd43088, 16'd20783, 16'd14474, 16'd15430, 16'd38024, 16'd52991, 16'd30238, 16'd61363, 16'd26179, 16'd16301, 16'd60373, 16'd54314, 16'd8814, 16'd2485, 16'd60470, 16'd60577, 16'd24247, 16'd20221, 16'd28784, 16'd34771, 16'd57774, 16'd46516, 16'd8204, 16'd10545, 16'd29956});
	test_expansion(128'h66bc88029bca5107f06581975caaab9c, {16'd21140, 16'd54917, 16'd21508, 16'd19575, 16'd8221, 16'd28802, 16'd38525, 16'd31427, 16'd30307, 16'd54994, 16'd60390, 16'd60510, 16'd32648, 16'd41044, 16'd64469, 16'd48176, 16'd33588, 16'd4255, 16'd50323, 16'd24893, 16'd59136, 16'd55873, 16'd11470, 16'd51294, 16'd52539, 16'd50880});
	test_expansion(128'h6908d839ff3c5acfe897cf50555231c4, {16'd4979, 16'd33553, 16'd20759, 16'd45334, 16'd61393, 16'd30246, 16'd4942, 16'd47645, 16'd64737, 16'd46946, 16'd4737, 16'd25427, 16'd15022, 16'd42890, 16'd60758, 16'd53902, 16'd63067, 16'd13415, 16'd21976, 16'd10498, 16'd62716, 16'd6425, 16'd10481, 16'd51923, 16'd7800, 16'd49532});
	test_expansion(128'h0257cbfac955bdbf615b297e0248a6ab, {16'd589, 16'd37409, 16'd13169, 16'd35311, 16'd53897, 16'd31720, 16'd18640, 16'd23517, 16'd62706, 16'd56952, 16'd21447, 16'd34186, 16'd38343, 16'd58144, 16'd34019, 16'd23849, 16'd3124, 16'd46982, 16'd9116, 16'd22028, 16'd28827, 16'd9107, 16'd61528, 16'd51539, 16'd40666, 16'd51764});
	test_expansion(128'h915459a99d048be94b73cdb94f6a3a4e, {16'd13148, 16'd48292, 16'd20291, 16'd55085, 16'd28884, 16'd33286, 16'd54770, 16'd3766, 16'd41300, 16'd64570, 16'd31889, 16'd12383, 16'd13994, 16'd42415, 16'd13538, 16'd63221, 16'd2587, 16'd33588, 16'd11274, 16'd23188, 16'd48529, 16'd45854, 16'd21387, 16'd43768, 16'd11146, 16'd49563});
	test_expansion(128'h947f495144f872d742ec1555093b58bf, {16'd26939, 16'd54235, 16'd33769, 16'd23572, 16'd24202, 16'd60522, 16'd8370, 16'd48028, 16'd7900, 16'd47932, 16'd60851, 16'd50844, 16'd51528, 16'd43682, 16'd37980, 16'd63000, 16'd52386, 16'd49141, 16'd9222, 16'd21211, 16'd57772, 16'd17357, 16'd3891, 16'd29565, 16'd43627, 16'd61796});
	test_expansion(128'hed125e77ae73fb7becdd4648399d344c, {16'd52010, 16'd30767, 16'd37407, 16'd24327, 16'd40435, 16'd57739, 16'd59018, 16'd46919, 16'd53270, 16'd48250, 16'd32349, 16'd19626, 16'd54328, 16'd7093, 16'd54483, 16'd45540, 16'd55466, 16'd60024, 16'd48149, 16'd48010, 16'd3550, 16'd41792, 16'd45318, 16'd60798, 16'd39095, 16'd27886});
	test_expansion(128'hc270bfd37b9756e3d09de8f4e4077653, {16'd6412, 16'd2058, 16'd63136, 16'd56364, 16'd36444, 16'd58247, 16'd13739, 16'd19977, 16'd19808, 16'd44501, 16'd19183, 16'd34844, 16'd46950, 16'd8465, 16'd35411, 16'd51291, 16'd57640, 16'd10365, 16'd45791, 16'd21520, 16'd1270, 16'd3409, 16'd8336, 16'd22494, 16'd7000, 16'd53786});
	test_expansion(128'h1783c863645c25765f80612afd07c1d9, {16'd18896, 16'd35071, 16'd26830, 16'd41572, 16'd11152, 16'd41639, 16'd20069, 16'd62311, 16'd59162, 16'd47972, 16'd38145, 16'd12771, 16'd9172, 16'd26348, 16'd65205, 16'd38639, 16'd28104, 16'd54829, 16'd4949, 16'd58691, 16'd10923, 16'd4515, 16'd22570, 16'd50172, 16'd26403, 16'd26443});
	test_expansion(128'hf9326e3ad3f395e7f4efbe79d41bc0dc, {16'd52996, 16'd29772, 16'd62487, 16'd42143, 16'd45, 16'd26592, 16'd30584, 16'd58788, 16'd508, 16'd38099, 16'd27948, 16'd60091, 16'd48491, 16'd2627, 16'd63453, 16'd20443, 16'd29013, 16'd57975, 16'd32070, 16'd52351, 16'd58840, 16'd31154, 16'd48815, 16'd18220, 16'd21081, 16'd38397});
	test_expansion(128'hce6d54c3ce791783ca475a9fcaedbd3f, {16'd48880, 16'd50628, 16'd58283, 16'd35650, 16'd34034, 16'd4885, 16'd23768, 16'd38577, 16'd59318, 16'd57925, 16'd29765, 16'd44892, 16'd22180, 16'd50589, 16'd31545, 16'd30128, 16'd30894, 16'd37104, 16'd61958, 16'd17188, 16'd476, 16'd34058, 16'd65051, 16'd39186, 16'd5666, 16'd23465});
	test_expansion(128'h597e43df0d3262a96de95bdd2ecf3f0d, {16'd55104, 16'd47795, 16'd1914, 16'd62930, 16'd11335, 16'd36975, 16'd24596, 16'd2430, 16'd18116, 16'd26258, 16'd172, 16'd28003, 16'd6167, 16'd11833, 16'd42105, 16'd26103, 16'd16379, 16'd36761, 16'd8673, 16'd45495, 16'd7964, 16'd5065, 16'd4580, 16'd41013, 16'd49627, 16'd7120});
	test_expansion(128'hbfac44c42a3e9aa5793981241762c138, {16'd33916, 16'd63297, 16'd28916, 16'd7277, 16'd9947, 16'd21786, 16'd8058, 16'd21373, 16'd2683, 16'd26048, 16'd51086, 16'd3185, 16'd5729, 16'd27653, 16'd27565, 16'd7109, 16'd800, 16'd53358, 16'd7681, 16'd56858, 16'd11877, 16'd43403, 16'd31928, 16'd47098, 16'd22427, 16'd20345});
	test_expansion(128'h084644c0ad8c3bb402b0fdecb59657f4, {16'd59622, 16'd60749, 16'd5576, 16'd11777, 16'd37871, 16'd33987, 16'd55379, 16'd15285, 16'd40233, 16'd37471, 16'd8446, 16'd60335, 16'd16078, 16'd47045, 16'd41338, 16'd34397, 16'd55152, 16'd18596, 16'd37869, 16'd64837, 16'd44766, 16'd39749, 16'd162, 16'd25260, 16'd25893, 16'd35941});
	test_expansion(128'h0b044f09e74b593281d343cba3853f92, {16'd33422, 16'd24443, 16'd5766, 16'd61523, 16'd23797, 16'd3075, 16'd56810, 16'd4654, 16'd59755, 16'd58242, 16'd35109, 16'd5471, 16'd28389, 16'd62590, 16'd27098, 16'd57861, 16'd21791, 16'd11904, 16'd31113, 16'd25397, 16'd38280, 16'd64769, 16'd24454, 16'd969, 16'd45163, 16'd12903});
	test_expansion(128'hf9cca4cc08438fc8f8452a15d7c39c52, {16'd11458, 16'd50312, 16'd27689, 16'd57409, 16'd63776, 16'd1632, 16'd37693, 16'd47703, 16'd17800, 16'd52703, 16'd21037, 16'd16947, 16'd1222, 16'd25245, 16'd37019, 16'd6606, 16'd17681, 16'd64694, 16'd1125, 16'd11810, 16'd36064, 16'd21140, 16'd38820, 16'd31287, 16'd31846, 16'd332});
	test_expansion(128'h3ce5f9f77eaaa3b43eb10fa4494649e2, {16'd30270, 16'd4631, 16'd8219, 16'd2108, 16'd25453, 16'd43937, 16'd58099, 16'd19973, 16'd49181, 16'd605, 16'd20204, 16'd20894, 16'd46598, 16'd39191, 16'd4480, 16'd29720, 16'd2029, 16'd25963, 16'd1620, 16'd19856, 16'd64254, 16'd55148, 16'd32917, 16'd13501, 16'd5851, 16'd51720});
	test_expansion(128'he46a318145b8a7170c3cc183e5e008da, {16'd8302, 16'd26784, 16'd16857, 16'd25492, 16'd19827, 16'd912, 16'd10056, 16'd51792, 16'd49985, 16'd50710, 16'd58018, 16'd17332, 16'd15619, 16'd46471, 16'd50420, 16'd1702, 16'd8727, 16'd61931, 16'd6681, 16'd32206, 16'd51594, 16'd7199, 16'd32526, 16'd9896, 16'd52222, 16'd46612});
	test_expansion(128'h37080e7f4c7451fdd71c00afbb3bf2e4, {16'd41280, 16'd48778, 16'd43548, 16'd12170, 16'd21425, 16'd19989, 16'd44569, 16'd22485, 16'd64297, 16'd25159, 16'd25230, 16'd29084, 16'd2806, 16'd8068, 16'd6817, 16'd43477, 16'd7963, 16'd52038, 16'd50937, 16'd16383, 16'd20924, 16'd11329, 16'd54717, 16'd41747, 16'd61057, 16'd57132});
	test_expansion(128'h40ed22808c9d449d994f0a62fc603bab, {16'd16643, 16'd22049, 16'd48405, 16'd9548, 16'd44692, 16'd6389, 16'd32948, 16'd4759, 16'd43164, 16'd24189, 16'd55631, 16'd20643, 16'd62878, 16'd33540, 16'd8793, 16'd18170, 16'd42679, 16'd45591, 16'd9479, 16'd15902, 16'd31589, 16'd3040, 16'd10429, 16'd58104, 16'd46063, 16'd56124});
	test_expansion(128'h7ba017faebe0a58ef3908da66d790dee, {16'd40245, 16'd60537, 16'd40188, 16'd61249, 16'd5429, 16'd32267, 16'd25133, 16'd39652, 16'd26786, 16'd4029, 16'd61978, 16'd41427, 16'd18392, 16'd53020, 16'd7004, 16'd57199, 16'd20000, 16'd32464, 16'd28944, 16'd31282, 16'd27227, 16'd62472, 16'd36730, 16'd17799, 16'd26085, 16'd12851});
	test_expansion(128'ha50c735da42791b34c2c3d646ed8dc94, {16'd27519, 16'd57500, 16'd39980, 16'd46621, 16'd37173, 16'd19825, 16'd30094, 16'd11157, 16'd11318, 16'd39004, 16'd41078, 16'd43953, 16'd56595, 16'd64820, 16'd21558, 16'd44061, 16'd60598, 16'd41657, 16'd12577, 16'd25318, 16'd2741, 16'd9746, 16'd22442, 16'd30353, 16'd35059, 16'd27829});
	test_expansion(128'h6f8ed8b1ba00c9b63ae5cab2c9e8794f, {16'd23662, 16'd8388, 16'd28856, 16'd34575, 16'd12051, 16'd57554, 16'd48349, 16'd14462, 16'd41734, 16'd9034, 16'd39381, 16'd53082, 16'd37331, 16'd33326, 16'd28953, 16'd24030, 16'd7084, 16'd42865, 16'd27352, 16'd64121, 16'd21252, 16'd21936, 16'd14381, 16'd56834, 16'd24927, 16'd40229});
	test_expansion(128'hd560ae94b46814c848586288388bd82b, {16'd4661, 16'd528, 16'd9088, 16'd64976, 16'd6229, 16'd38699, 16'd42575, 16'd44783, 16'd19087, 16'd14046, 16'd17375, 16'd51716, 16'd62522, 16'd28074, 16'd59169, 16'd23133, 16'd14755, 16'd42600, 16'd18299, 16'd34111, 16'd29173, 16'd55193, 16'd24065, 16'd34697, 16'd1408, 16'd46108});
	test_expansion(128'hc93959e96c3ccb05f644ee9dfd4fa2d4, {16'd7678, 16'd43130, 16'd55226, 16'd23046, 16'd30399, 16'd61422, 16'd57142, 16'd6548, 16'd20711, 16'd36759, 16'd62370, 16'd52996, 16'd36457, 16'd26132, 16'd32247, 16'd60137, 16'd21537, 16'd3593, 16'd64370, 16'd28822, 16'd33233, 16'd37685, 16'd5639, 16'd452, 16'd31921, 16'd37546});
	test_expansion(128'h8703ed4f426a32b4afa172e9f10dcf64, {16'd16957, 16'd42972, 16'd40184, 16'd44195, 16'd48182, 16'd51618, 16'd7999, 16'd26851, 16'd41817, 16'd40463, 16'd55992, 16'd2894, 16'd30716, 16'd41119, 16'd10072, 16'd63549, 16'd43345, 16'd8365, 16'd17260, 16'd41190, 16'd12113, 16'd48576, 16'd15533, 16'd40397, 16'd59210, 16'd31718});
	test_expansion(128'h35b416f96bedc9646de6febb0c79c3c0, {16'd6754, 16'd40347, 16'd57092, 16'd6666, 16'd48083, 16'd5944, 16'd63790, 16'd26033, 16'd10776, 16'd60596, 16'd38142, 16'd61703, 16'd37621, 16'd36321, 16'd22528, 16'd50965, 16'd12934, 16'd65273, 16'd15194, 16'd22318, 16'd14090, 16'd29757, 16'd20258, 16'd64963, 16'd32847, 16'd58010});
	test_expansion(128'heeed103d38bdf5a7158e220d342e26f2, {16'd23441, 16'd12723, 16'd24345, 16'd12454, 16'd10244, 16'd20469, 16'd22628, 16'd56634, 16'd56459, 16'd2152, 16'd59092, 16'd38080, 16'd55903, 16'd50910, 16'd44860, 16'd36063, 16'd31575, 16'd50010, 16'd48811, 16'd46377, 16'd46111, 16'd31795, 16'd54089, 16'd62602, 16'd30951, 16'd53918});
	test_expansion(128'hfe4b967078b81511ca201dd14228e035, {16'd52300, 16'd51591, 16'd58132, 16'd48284, 16'd32027, 16'd36406, 16'd8144, 16'd3880, 16'd20163, 16'd29749, 16'd45033, 16'd47949, 16'd16787, 16'd29981, 16'd9740, 16'd32594, 16'd27627, 16'd56359, 16'd45630, 16'd50413, 16'd48376, 16'd30760, 16'd26238, 16'd54244, 16'd25118, 16'd42364});
	test_expansion(128'h3cf8449842bcca6bba7e443f62286a82, {16'd42070, 16'd22725, 16'd39193, 16'd28491, 16'd21598, 16'd11587, 16'd43718, 16'd35701, 16'd26308, 16'd62558, 16'd31779, 16'd39618, 16'd13376, 16'd49115, 16'd18302, 16'd12211, 16'd14473, 16'd47532, 16'd49601, 16'd44668, 16'd28137, 16'd1890, 16'd5217, 16'd21091, 16'd9062, 16'd36629});
	test_expansion(128'h7666454f4ef9f7c60fa6be31555a1692, {16'd28429, 16'd20718, 16'd62728, 16'd55023, 16'd37608, 16'd45563, 16'd35130, 16'd10056, 16'd2162, 16'd25969, 16'd29295, 16'd38111, 16'd53207, 16'd19054, 16'd40475, 16'd8626, 16'd8000, 16'd58074, 16'd35095, 16'd54430, 16'd37596, 16'd18902, 16'd49163, 16'd3638, 16'd22009, 16'd54936});
	test_expansion(128'hbe40ee28b3cff69fe10fac8052e87631, {16'd62461, 16'd7440, 16'd7763, 16'd48513, 16'd6609, 16'd32318, 16'd17123, 16'd34793, 16'd31519, 16'd42942, 16'd44040, 16'd59682, 16'd34183, 16'd39518, 16'd8072, 16'd8343, 16'd65352, 16'd26315, 16'd577, 16'd22350, 16'd23874, 16'd43018, 16'd45659, 16'd26741, 16'd61401, 16'd27656});
	test_expansion(128'hdcf7229c91e69ed5ede0f4f7269a05ea, {16'd49618, 16'd1333, 16'd5313, 16'd22038, 16'd39888, 16'd32051, 16'd24740, 16'd22421, 16'd40483, 16'd54591, 16'd22720, 16'd8421, 16'd64172, 16'd53508, 16'd35258, 16'd28189, 16'd23626, 16'd40978, 16'd12960, 16'd42074, 16'd41450, 16'd27132, 16'd54264, 16'd48469, 16'd6186, 16'd65117});
	test_expansion(128'h5fe0e9c0eb066ffe6a1fa826c7a60f25, {16'd18137, 16'd53447, 16'd59820, 16'd57850, 16'd61093, 16'd11746, 16'd2967, 16'd13570, 16'd19444, 16'd35157, 16'd17272, 16'd45627, 16'd61878, 16'd15906, 16'd16292, 16'd64074, 16'd20627, 16'd50370, 16'd51836, 16'd33007, 16'd24528, 16'd12205, 16'd46831, 16'd7809, 16'd65266, 16'd6052});
	test_expansion(128'hab03e12dab45857ae9f9bed6083f4993, {16'd20500, 16'd26966, 16'd62994, 16'd32096, 16'd52248, 16'd53387, 16'd13389, 16'd53453, 16'd49637, 16'd41106, 16'd41203, 16'd3421, 16'd5180, 16'd44888, 16'd55165, 16'd43303, 16'd57250, 16'd9346, 16'd59055, 16'd24473, 16'd58501, 16'd32071, 16'd50018, 16'd42525, 16'd28740, 16'd26117});
	test_expansion(128'h93a764cd2ff05b2f8c0c3342188e1f2c, {16'd42757, 16'd17535, 16'd36375, 16'd537, 16'd38903, 16'd25274, 16'd41465, 16'd28535, 16'd55284, 16'd26231, 16'd60383, 16'd1234, 16'd9264, 16'd39150, 16'd49849, 16'd56197, 16'd48304, 16'd52917, 16'd26883, 16'd27951, 16'd1673, 16'd59544, 16'd8151, 16'd5753, 16'd49604, 16'd3489});
	test_expansion(128'h84209cd077f2097f6e4b27f157f852bc, {16'd9756, 16'd19146, 16'd23382, 16'd36182, 16'd5778, 16'd32162, 16'd22899, 16'd51779, 16'd34895, 16'd64557, 16'd13153, 16'd18328, 16'd48784, 16'd52202, 16'd65487, 16'd65091, 16'd38533, 16'd43985, 16'd21819, 16'd4138, 16'd55483, 16'd49572, 16'd7159, 16'd12197, 16'd4149, 16'd21097});
	test_expansion(128'hbe562de390f3e52ee54883a6fa4efd9c, {16'd30855, 16'd55799, 16'd32443, 16'd16706, 16'd60479, 16'd17332, 16'd40837, 16'd48392, 16'd44172, 16'd9031, 16'd22192, 16'd48312, 16'd54564, 16'd4672, 16'd41221, 16'd21910, 16'd47528, 16'd21982, 16'd27523, 16'd37055, 16'd54767, 16'd33000, 16'd3479, 16'd44831, 16'd24355, 16'd30874});
	test_expansion(128'h7e2d0f64fdef9b5c8c86de0896f65ba3, {16'd46481, 16'd7764, 16'd14231, 16'd20803, 16'd18011, 16'd20416, 16'd62357, 16'd32480, 16'd11971, 16'd8800, 16'd11467, 16'd40046, 16'd31244, 16'd12500, 16'd61431, 16'd14476, 16'd19447, 16'd52977, 16'd44456, 16'd10170, 16'd14330, 16'd58172, 16'd6695, 16'd37240, 16'd15263, 16'd47958});
	test_expansion(128'h23d4a84f40dca9a877fa9185c2134d3c, {16'd29500, 16'd60314, 16'd38141, 16'd6137, 16'd63188, 16'd4002, 16'd7913, 16'd40959, 16'd59299, 16'd41182, 16'd39941, 16'd16222, 16'd19985, 16'd30526, 16'd33478, 16'd41697, 16'd65364, 16'd18843, 16'd42535, 16'd44881, 16'd62078, 16'd50543, 16'd35908, 16'd23016, 16'd20448, 16'd64853});
	test_expansion(128'h5367464b5c5c2f38deafe44236b1b218, {16'd34571, 16'd25682, 16'd48895, 16'd4983, 16'd45192, 16'd45871, 16'd14704, 16'd44381, 16'd47527, 16'd27866, 16'd58739, 16'd62761, 16'd37953, 16'd35242, 16'd35925, 16'd20329, 16'd45555, 16'd56208, 16'd23023, 16'd44022, 16'd6564, 16'd6977, 16'd15432, 16'd62233, 16'd60047, 16'd58648});
	test_expansion(128'h4ab3f6a8269b245b32b23139ca8c097e, {16'd38128, 16'd23696, 16'd28166, 16'd38537, 16'd5389, 16'd11688, 16'd63930, 16'd46086, 16'd16127, 16'd17306, 16'd42826, 16'd45819, 16'd18962, 16'd59510, 16'd3240, 16'd49211, 16'd56492, 16'd17424, 16'd42767, 16'd3649, 16'd37895, 16'd49268, 16'd29107, 16'd21823, 16'd26071, 16'd17711});
	test_expansion(128'h5f4087c2c7d6114814e2bedb84649cbf, {16'd25517, 16'd61586, 16'd43579, 16'd41759, 16'd59870, 16'd37739, 16'd19139, 16'd53094, 16'd31515, 16'd30928, 16'd14028, 16'd45719, 16'd49207, 16'd46975, 16'd52747, 16'd42846, 16'd4915, 16'd11612, 16'd18786, 16'd30089, 16'd43849, 16'd45451, 16'd37410, 16'd24329, 16'd42990, 16'd16509});
	test_expansion(128'h6548d1ce13f84e3582265f3fad4ecc9a, {16'd65414, 16'd989, 16'd24721, 16'd58405, 16'd51811, 16'd57260, 16'd8978, 16'd40297, 16'd11202, 16'd30038, 16'd44778, 16'd60970, 16'd1610, 16'd45522, 16'd60696, 16'd49263, 16'd31556, 16'd46520, 16'd55707, 16'd23244, 16'd4553, 16'd21879, 16'd55691, 16'd8136, 16'd7069, 16'd18011});
	test_expansion(128'h0f22c24be8a87e265436e1db81ad4f15, {16'd11923, 16'd48814, 16'd25763, 16'd8397, 16'd54199, 16'd45014, 16'd41742, 16'd419, 16'd7260, 16'd9636, 16'd291, 16'd44646, 16'd13318, 16'd40168, 16'd45984, 16'd49963, 16'd10228, 16'd22716, 16'd37228, 16'd53868, 16'd50306, 16'd27357, 16'd74, 16'd27176, 16'd13759, 16'd16823});
	test_expansion(128'h5d74a27e57db85b41823a6475872ba48, {16'd57140, 16'd53326, 16'd18119, 16'd4784, 16'd28642, 16'd57756, 16'd33352, 16'd45767, 16'd41933, 16'd41798, 16'd55476, 16'd42161, 16'd29774, 16'd14513, 16'd4835, 16'd8098, 16'd23473, 16'd62836, 16'd47755, 16'd48589, 16'd31858, 16'd63895, 16'd12815, 16'd25236, 16'd35545, 16'd20394});
	test_expansion(128'h6a0ed7774b37e1bfd1598229ad673ca8, {16'd59947, 16'd28008, 16'd25473, 16'd6656, 16'd12938, 16'd50117, 16'd53158, 16'd11028, 16'd50397, 16'd39450, 16'd61871, 16'd48775, 16'd63855, 16'd23861, 16'd43413, 16'd61675, 16'd50061, 16'd16788, 16'd20619, 16'd15265, 16'd21809, 16'd55893, 16'd27752, 16'd15815, 16'd65067, 16'd11490});
	test_expansion(128'h8e35da35e244c4f0f987774f99d9f516, {16'd1801, 16'd56037, 16'd47236, 16'd39201, 16'd8230, 16'd8858, 16'd31307, 16'd2377, 16'd58359, 16'd12907, 16'd44428, 16'd34931, 16'd46359, 16'd9780, 16'd18777, 16'd13012, 16'd1823, 16'd35872, 16'd16986, 16'd48977, 16'd15617, 16'd14430, 16'd56805, 16'd392, 16'd14884, 16'd19340});
	test_expansion(128'h62d9d8eeecc590d175d9e8926c7a53d6, {16'd51687, 16'd25817, 16'd14261, 16'd56183, 16'd41108, 16'd57134, 16'd45612, 16'd14085, 16'd25005, 16'd14178, 16'd20181, 16'd18541, 16'd3036, 16'd22019, 16'd173, 16'd50252, 16'd30495, 16'd29062, 16'd2170, 16'd7672, 16'd34339, 16'd9548, 16'd2210, 16'd46464, 16'd40901, 16'd23231});
	test_expansion(128'h61845bf6f93586b2359a3a4471ea8ccf, {16'd54079, 16'd40960, 16'd22524, 16'd26677, 16'd7041, 16'd62815, 16'd50213, 16'd57453, 16'd47940, 16'd8927, 16'd25598, 16'd18085, 16'd46133, 16'd18225, 16'd22115, 16'd36310, 16'd1882, 16'd30125, 16'd26920, 16'd21941, 16'd57825, 16'd43005, 16'd52968, 16'd56047, 16'd53004, 16'd8609});
	test_expansion(128'h3b874239674f56a6b16ab0e94e2d9f86, {16'd60290, 16'd60638, 16'd1081, 16'd40776, 16'd41446, 16'd54651, 16'd46769, 16'd28127, 16'd40515, 16'd22970, 16'd53815, 16'd28709, 16'd10400, 16'd49720, 16'd40468, 16'd44826, 16'd59197, 16'd49068, 16'd9632, 16'd4375, 16'd12706, 16'd1305, 16'd501, 16'd47080, 16'd26981, 16'd37039});
	test_expansion(128'h33bed540d69a35d8bdac8bd459867487, {16'd58730, 16'd16392, 16'd25240, 16'd61570, 16'd53536, 16'd52108, 16'd5782, 16'd33169, 16'd34696, 16'd22083, 16'd28915, 16'd1278, 16'd60414, 16'd40096, 16'd40814, 16'd40876, 16'd46067, 16'd51073, 16'd32859, 16'd11597, 16'd52847, 16'd515, 16'd27360, 16'd35864, 16'd14856, 16'd52296});
	test_expansion(128'he7d6c7f6e00120bee20a0c0cf47f9889, {16'd18985, 16'd9561, 16'd17552, 16'd16344, 16'd17628, 16'd32903, 16'd18981, 16'd22242, 16'd28508, 16'd3574, 16'd55282, 16'd54334, 16'd28276, 16'd18521, 16'd46991, 16'd28260, 16'd53195, 16'd8174, 16'd3962, 16'd16485, 16'd60164, 16'd25303, 16'd5112, 16'd4550, 16'd24170, 16'd12777});
	test_expansion(128'h2901eee4d130c7ec62ee4c730d77ab5a, {16'd45258, 16'd52452, 16'd59884, 16'd22308, 16'd23714, 16'd56530, 16'd31065, 16'd9435, 16'd38495, 16'd54551, 16'd43161, 16'd41238, 16'd9234, 16'd8059, 16'd53364, 16'd41964, 16'd57839, 16'd40021, 16'd26500, 16'd34092, 16'd47522, 16'd4566, 16'd56545, 16'd20648, 16'd43642, 16'd10940});
	test_expansion(128'hf3d8f18ed84b6ef3be86397605533cc4, {16'd32488, 16'd29443, 16'd35444, 16'd42165, 16'd11223, 16'd22570, 16'd62906, 16'd56559, 16'd2932, 16'd23053, 16'd22739, 16'd53176, 16'd23861, 16'd50676, 16'd8737, 16'd37860, 16'd103, 16'd29290, 16'd41839, 16'd38821, 16'd19965, 16'd26192, 16'd56034, 16'd29994, 16'd4445, 16'd5931});
	test_expansion(128'h1034ce16d48230bfdc211af4ef28ca3b, {16'd44732, 16'd14370, 16'd36695, 16'd23799, 16'd55831, 16'd13036, 16'd30670, 16'd29311, 16'd50319, 16'd47436, 16'd6335, 16'd22599, 16'd48437, 16'd51482, 16'd7368, 16'd1295, 16'd35601, 16'd20410, 16'd27095, 16'd51716, 16'd27237, 16'd11621, 16'd63151, 16'd21540, 16'd43437, 16'd34792});
	test_expansion(128'h0707be63b157d20ca6b66e7372c5f74a, {16'd33080, 16'd46665, 16'd49910, 16'd30925, 16'd8838, 16'd25482, 16'd27354, 16'd4104, 16'd44700, 16'd10588, 16'd48276, 16'd26510, 16'd40357, 16'd59419, 16'd16808, 16'd23303, 16'd46501, 16'd22146, 16'd37050, 16'd7326, 16'd24629, 16'd25351, 16'd57876, 16'd24175, 16'd19629, 16'd65038});
	test_expansion(128'headc941f993da0be5f5fc6a0475bbbd8, {16'd30122, 16'd60291, 16'd23200, 16'd13170, 16'd33554, 16'd24795, 16'd62993, 16'd6126, 16'd35883, 16'd22490, 16'd28199, 16'd22285, 16'd58279, 16'd55200, 16'd63617, 16'd52243, 16'd26520, 16'd53060, 16'd64135, 16'd16854, 16'd39772, 16'd44729, 16'd50671, 16'd20089, 16'd64918, 16'd9474});
	test_expansion(128'h10b43caa44f8a18ddff4bdb2af74fba4, {16'd17875, 16'd23332, 16'd8881, 16'd44768, 16'd64011, 16'd20845, 16'd16706, 16'd7418, 16'd29612, 16'd28497, 16'd58345, 16'd20590, 16'd4969, 16'd15978, 16'd44034, 16'd643, 16'd10841, 16'd38896, 16'd18273, 16'd6795, 16'd12544, 16'd4638, 16'd47830, 16'd26459, 16'd30050, 16'd3104});
	test_expansion(128'h854dc99ee121d51dc4ec073aa41b7b99, {16'd60267, 16'd5920, 16'd38472, 16'd51025, 16'd64539, 16'd57006, 16'd33607, 16'd64203, 16'd65323, 16'd41340, 16'd37346, 16'd24373, 16'd53783, 16'd30916, 16'd64234, 16'd16161, 16'd57911, 16'd15414, 16'd2013, 16'd58263, 16'd37113, 16'd33547, 16'd8869, 16'd46185, 16'd64507, 16'd18511});
	test_expansion(128'h9eb3efd455d10d07c2e78a71d2601b3c, {16'd43969, 16'd11796, 16'd7511, 16'd56363, 16'd41307, 16'd21174, 16'd65288, 16'd17885, 16'd35114, 16'd5161, 16'd10053, 16'd4347, 16'd25712, 16'd40422, 16'd47684, 16'd61622, 16'd20764, 16'd9701, 16'd53690, 16'd23459, 16'd23448, 16'd38377, 16'd25772, 16'd12295, 16'd38845, 16'd58298});
	test_expansion(128'hd340e67bdb3aa9cd383cbe603a4e03e9, {16'd62084, 16'd37430, 16'd38356, 16'd63099, 16'd1775, 16'd55806, 16'd25621, 16'd10811, 16'd39870, 16'd31894, 16'd16347, 16'd63904, 16'd6726, 16'd148, 16'd19366, 16'd34622, 16'd57290, 16'd33822, 16'd50074, 16'd35672, 16'd39576, 16'd55480, 16'd37067, 16'd59800, 16'd8086, 16'd54133});
	test_expansion(128'h3fbd35d8cf447890cee6eb57f8d8fba5, {16'd46524, 16'd2376, 16'd28274, 16'd13490, 16'd12957, 16'd31758, 16'd19108, 16'd31339, 16'd57901, 16'd35508, 16'd64728, 16'd7867, 16'd48616, 16'd39908, 16'd3396, 16'd22293, 16'd26688, 16'd46775, 16'd57850, 16'd60797, 16'd50481, 16'd54533, 16'd10326, 16'd21026, 16'd56243, 16'd44496});
	test_expansion(128'h00ab741b8d5b4e1ad9cb77c501a0f956, {16'd52224, 16'd31753, 16'd31507, 16'd65480, 16'd28530, 16'd57340, 16'd40007, 16'd64307, 16'd33870, 16'd50412, 16'd47964, 16'd44803, 16'd20298, 16'd12578, 16'd63525, 16'd13685, 16'd36631, 16'd7163, 16'd42814, 16'd12635, 16'd30855, 16'd35571, 16'd49604, 16'd31570, 16'd18761, 16'd21526});
	test_expansion(128'h05fb1e92515f6550cecb3ae90ef54b56, {16'd25398, 16'd39813, 16'd61650, 16'd24491, 16'd50039, 16'd3891, 16'd64504, 16'd11964, 16'd57999, 16'd19678, 16'd29647, 16'd51461, 16'd43932, 16'd31426, 16'd59927, 16'd4777, 16'd62951, 16'd7511, 16'd24872, 16'd16149, 16'd22292, 16'd22206, 16'd301, 16'd55404, 16'd46536, 16'd31168});
	test_expansion(128'hcaadb3d8a7d9b1bca1a9b939d757aa4e, {16'd62183, 16'd6295, 16'd52827, 16'd9482, 16'd31097, 16'd56098, 16'd23874, 16'd1811, 16'd51292, 16'd28825, 16'd52018, 16'd57684, 16'd6196, 16'd44965, 16'd37202, 16'd1685, 16'd33414, 16'd62128, 16'd35619, 16'd36546, 16'd45198, 16'd38728, 16'd47312, 16'd42125, 16'd38856, 16'd54369});
	test_expansion(128'h33381735c56c53f1e3b2f27fc8bf29a8, {16'd35806, 16'd58887, 16'd13363, 16'd52951, 16'd5892, 16'd11056, 16'd28025, 16'd9421, 16'd48160, 16'd11602, 16'd19717, 16'd27227, 16'd23983, 16'd54559, 16'd53295, 16'd55995, 16'd46424, 16'd10662, 16'd28500, 16'd11716, 16'd918, 16'd6025, 16'd26517, 16'd30626, 16'd32091, 16'd47308});
	test_expansion(128'h1b86d2fe3d28a0558435a2a0c17d1522, {16'd60592, 16'd9752, 16'd22503, 16'd8216, 16'd64155, 16'd35894, 16'd26650, 16'd34183, 16'd26363, 16'd32268, 16'd53610, 16'd21507, 16'd30657, 16'd7955, 16'd23805, 16'd28930, 16'd37937, 16'd27013, 16'd9073, 16'd38547, 16'd36267, 16'd9307, 16'd57708, 16'd54788, 16'd47441, 16'd518});
	test_expansion(128'h47717487a12bd1c6d029888b16e4a66b, {16'd3691, 16'd979, 16'd49146, 16'd28184, 16'd63344, 16'd46583, 16'd11535, 16'd1347, 16'd44072, 16'd7472, 16'd46205, 16'd38771, 16'd50762, 16'd46210, 16'd8062, 16'd42498, 16'd7266, 16'd33002, 16'd27084, 16'd56822, 16'd49919, 16'd47526, 16'd18754, 16'd36015, 16'd28922, 16'd26269});
	test_expansion(128'h53fccc1f80a354bfc89d407095c92b11, {16'd41232, 16'd23198, 16'd15747, 16'd36880, 16'd9649, 16'd37286, 16'd26384, 16'd20601, 16'd11606, 16'd7078, 16'd16279, 16'd45266, 16'd15868, 16'd7010, 16'd10194, 16'd22489, 16'd44742, 16'd51158, 16'd60414, 16'd34688, 16'd30665, 16'd13547, 16'd47298, 16'd61257, 16'd19833, 16'd13426});
	test_expansion(128'h4a7c27e76718763b38ae2dc047e36de1, {16'd30700, 16'd38996, 16'd4959, 16'd59227, 16'd38771, 16'd16437, 16'd18240, 16'd10670, 16'd5629, 16'd34632, 16'd43663, 16'd63233, 16'd55985, 16'd10329, 16'd19167, 16'd16083, 16'd4659, 16'd53125, 16'd62541, 16'd43323, 16'd26383, 16'd12042, 16'd16515, 16'd6619, 16'd31651, 16'd25219});
	test_expansion(128'h3e45dc0881874e1ebba5910dae5cee6d, {16'd44035, 16'd26636, 16'd36414, 16'd11907, 16'd36560, 16'd47424, 16'd6610, 16'd13338, 16'd14332, 16'd52130, 16'd6940, 16'd41096, 16'd19645, 16'd46820, 16'd32207, 16'd53962, 16'd43701, 16'd35440, 16'd47099, 16'd47868, 16'd15625, 16'd49194, 16'd45498, 16'd2604, 16'd79, 16'd49146});
	test_expansion(128'h1720450a114295088724ddb2eb46ee52, {16'd63028, 16'd16936, 16'd48097, 16'd16420, 16'd54932, 16'd7083, 16'd2733, 16'd60960, 16'd37918, 16'd12894, 16'd31688, 16'd14693, 16'd34392, 16'd26197, 16'd5029, 16'd40567, 16'd48458, 16'd62007, 16'd17951, 16'd16258, 16'd17381, 16'd57142, 16'd50625, 16'd12837, 16'd55302, 16'd64240});
	test_expansion(128'h3e0e932ce2a8fc8caf24fdf209a9d2f9, {16'd10461, 16'd38768, 16'd35305, 16'd41675, 16'd11817, 16'd13397, 16'd5000, 16'd10679, 16'd3512, 16'd29226, 16'd2366, 16'd36776, 16'd27222, 16'd15847, 16'd50642, 16'd60196, 16'd48417, 16'd42996, 16'd52610, 16'd59811, 16'd63380, 16'd58206, 16'd16143, 16'd9212, 16'd58135, 16'd57887});
	test_expansion(128'hba4e576957dba27ff0b55b18325166b1, {16'd24051, 16'd20260, 16'd41924, 16'd41776, 16'd599, 16'd26379, 16'd52147, 16'd17329, 16'd61965, 16'd37865, 16'd57622, 16'd7105, 16'd25911, 16'd59931, 16'd44491, 16'd12345, 16'd9121, 16'd22916, 16'd23531, 16'd52446, 16'd62730, 16'd43473, 16'd48088, 16'd51963, 16'd17149, 16'd51846});
	test_expansion(128'h749219d24192f690db75bb6db0611ea8, {16'd28982, 16'd54839, 16'd10708, 16'd34578, 16'd58616, 16'd6152, 16'd59340, 16'd30761, 16'd32161, 16'd44656, 16'd36707, 16'd46389, 16'd27269, 16'd63978, 16'd2088, 16'd30235, 16'd27342, 16'd62940, 16'd10048, 16'd12071, 16'd50163, 16'd63605, 16'd31632, 16'd45277, 16'd48184, 16'd9965});
	test_expansion(128'hf47bfe6ee238c712ebe5ccd8c499d20a, {16'd11178, 16'd16697, 16'd55115, 16'd25744, 16'd23178, 16'd47165, 16'd23495, 16'd43261, 16'd21949, 16'd17494, 16'd24653, 16'd39798, 16'd58849, 16'd30390, 16'd56253, 16'd9790, 16'd1794, 16'd368, 16'd52075, 16'd53815, 16'd11243, 16'd31531, 16'd18898, 16'd56529, 16'd41948, 16'd23377});
	test_expansion(128'h671cc1d568961cd7a797b9cf0ccaf607, {16'd8828, 16'd36839, 16'd30411, 16'd53358, 16'd41005, 16'd52808, 16'd25600, 16'd17512, 16'd46693, 16'd30912, 16'd54516, 16'd45715, 16'd59264, 16'd3438, 16'd38055, 16'd24780, 16'd27415, 16'd34011, 16'd40934, 16'd12048, 16'd58195, 16'd62384, 16'd57646, 16'd51781, 16'd30437, 16'd2612});
	test_expansion(128'h0b08d7692b041b98f5012bd1eb7f1f46, {16'd9003, 16'd10783, 16'd49944, 16'd61714, 16'd29058, 16'd3677, 16'd50046, 16'd64254, 16'd27337, 16'd64374, 16'd2332, 16'd62625, 16'd1159, 16'd30193, 16'd3670, 16'd2956, 16'd53458, 16'd19424, 16'd20103, 16'd25912, 16'd51617, 16'd61287, 16'd18835, 16'd21180, 16'd51693, 16'd33433});
	test_expansion(128'hf7e4f3b6eb45d3fe8bef34ddcdd23c26, {16'd63228, 16'd65333, 16'd26332, 16'd5589, 16'd44263, 16'd15425, 16'd14941, 16'd40759, 16'd51393, 16'd6374, 16'd2836, 16'd30330, 16'd59295, 16'd58072, 16'd51262, 16'd47773, 16'd20503, 16'd33140, 16'd8994, 16'd11756, 16'd62234, 16'd48166, 16'd2879, 16'd47414, 16'd39171, 16'd11057});
	test_expansion(128'hb37bc092388a525740668de74525e948, {16'd62845, 16'd47643, 16'd9674, 16'd19829, 16'd31813, 16'd6030, 16'd61350, 16'd32090, 16'd51550, 16'd49890, 16'd63790, 16'd42526, 16'd2266, 16'd31950, 16'd25609, 16'd41173, 16'd55476, 16'd1182, 16'd34257, 16'd5420, 16'd25476, 16'd52531, 16'd52405, 16'd27342, 16'd834, 16'd3464});
	test_expansion(128'hfb4b8a0148636e72e59b47de81587eba, {16'd31031, 16'd53241, 16'd54528, 16'd29618, 16'd10865, 16'd64162, 16'd44843, 16'd15950, 16'd60940, 16'd51865, 16'd19278, 16'd4152, 16'd20024, 16'd33417, 16'd55250, 16'd17703, 16'd59174, 16'd24194, 16'd47775, 16'd47134, 16'd33631, 16'd24484, 16'd53044, 16'd62661, 16'd22741, 16'd54657});
	test_expansion(128'h65a3e54ea400457aa5db0713a5678cc8, {16'd49772, 16'd13306, 16'd34621, 16'd33451, 16'd29093, 16'd37668, 16'd60165, 16'd52958, 16'd13996, 16'd8740, 16'd58341, 16'd36891, 16'd58573, 16'd56048, 16'd5204, 16'd6448, 16'd32136, 16'd1073, 16'd13340, 16'd63866, 16'd58712, 16'd39118, 16'd37925, 16'd41046, 16'd12134, 16'd63482});
	test_expansion(128'h10bdfdcad1219f9665c21ecdb58e6667, {16'd19705, 16'd47841, 16'd4281, 16'd36186, 16'd62835, 16'd61870, 16'd3935, 16'd48005, 16'd53979, 16'd20853, 16'd11162, 16'd6472, 16'd6301, 16'd5508, 16'd40474, 16'd48062, 16'd22585, 16'd8993, 16'd13287, 16'd9328, 16'd26616, 16'd61686, 16'd48486, 16'd48142, 16'd164, 16'd24588});
	test_expansion(128'h579b5a8a65117975e4231f82c0c73024, {16'd38475, 16'd43169, 16'd39401, 16'd392, 16'd44200, 16'd51084, 16'd3429, 16'd3461, 16'd22498, 16'd15746, 16'd54988, 16'd12504, 16'd59510, 16'd52303, 16'd43893, 16'd44262, 16'd1543, 16'd25328, 16'd12126, 16'd57642, 16'd37870, 16'd8888, 16'd17431, 16'd28367, 16'd12495, 16'd32733});
	test_expansion(128'h7df57d3e8d9f3b9cf92eca0496950e1b, {16'd17718, 16'd64367, 16'd45434, 16'd53484, 16'd22989, 16'd16470, 16'd54749, 16'd36717, 16'd58395, 16'd64144, 16'd59658, 16'd37199, 16'd12475, 16'd29546, 16'd16272, 16'd36339, 16'd29925, 16'd28625, 16'd24308, 16'd20592, 16'd63199, 16'd28619, 16'd23292, 16'd54509, 16'd37862, 16'd6761});
	test_expansion(128'h4645f0a63813228f16c754985a2e8e4e, {16'd56900, 16'd49105, 16'd34671, 16'd26629, 16'd9108, 16'd48992, 16'd34395, 16'd54266, 16'd9891, 16'd22017, 16'd55062, 16'd62742, 16'd1996, 16'd28466, 16'd33438, 16'd49780, 16'd42515, 16'd918, 16'd55708, 16'd28273, 16'd15923, 16'd64068, 16'd45884, 16'd62335, 16'd44974, 16'd35713});
	test_expansion(128'h5372acb3f169789265720fc10a064576, {16'd44236, 16'd15400, 16'd15011, 16'd21476, 16'd44814, 16'd52798, 16'd51859, 16'd21808, 16'd19917, 16'd4507, 16'd35464, 16'd25930, 16'd56892, 16'd36954, 16'd4874, 16'd40470, 16'd53865, 16'd20738, 16'd58075, 16'd60589, 16'd55822, 16'd2354, 16'd28521, 16'd45279, 16'd60869, 16'd37963});
	test_expansion(128'hc4194794014f88abd4df5208b8c40da8, {16'd49448, 16'd19089, 16'd57981, 16'd41202, 16'd48651, 16'd1865, 16'd51135, 16'd54731, 16'd3414, 16'd20416, 16'd16642, 16'd18832, 16'd27466, 16'd23405, 16'd12738, 16'd44575, 16'd60927, 16'd19206, 16'd8370, 16'd54682, 16'd30212, 16'd4035, 16'd55335, 16'd3436, 16'd59620, 16'd22059});
	test_expansion(128'h1e8ab1f77809e8deaeab529dc8fc96bb, {16'd27933, 16'd43659, 16'd41668, 16'd50781, 16'd37479, 16'd8256, 16'd14143, 16'd62974, 16'd28846, 16'd12298, 16'd10668, 16'd19798, 16'd24234, 16'd52212, 16'd46598, 16'd18975, 16'd7758, 16'd26060, 16'd9927, 16'd48003, 16'd34175, 16'd1611, 16'd49761, 16'd23193, 16'd55057, 16'd4266});
	test_expansion(128'h9742c3971e5ca7699c9e79e69b0de51b, {16'd12022, 16'd60282, 16'd39888, 16'd10374, 16'd39760, 16'd12094, 16'd45359, 16'd40150, 16'd54428, 16'd43115, 16'd63280, 16'd57706, 16'd33652, 16'd24851, 16'd9597, 16'd58108, 16'd51805, 16'd40244, 16'd29649, 16'd29970, 16'd8173, 16'd6722, 16'd6987, 16'd7724, 16'd33186, 16'd39731});
	test_expansion(128'h9e833acfadc69a76046eaf05748c251a, {16'd28804, 16'd43616, 16'd53903, 16'd20034, 16'd50941, 16'd51675, 16'd34936, 16'd26207, 16'd2731, 16'd6508, 16'd47650, 16'd50255, 16'd32375, 16'd4024, 16'd54438, 16'd16009, 16'd6237, 16'd48405, 16'd38984, 16'd46357, 16'd39132, 16'd1776, 16'd40892, 16'd14214, 16'd62245, 16'd6853});
	test_expansion(128'h9e9720d22b5fb7420be5d92c796f90d1, {16'd34701, 16'd45347, 16'd25909, 16'd31224, 16'd50535, 16'd58346, 16'd31492, 16'd62989, 16'd64368, 16'd59613, 16'd21884, 16'd7887, 16'd20713, 16'd64268, 16'd62215, 16'd31828, 16'd3467, 16'd30952, 16'd47438, 16'd35636, 16'd18093, 16'd37984, 16'd40892, 16'd14615, 16'd61962, 16'd28332});
	test_expansion(128'hef5576176a0795d60539de8a6c7f3652, {16'd57815, 16'd14319, 16'd45712, 16'd52899, 16'd24964, 16'd47412, 16'd48115, 16'd54281, 16'd33986, 16'd21759, 16'd35397, 16'd13741, 16'd42501, 16'd55568, 16'd13663, 16'd7735, 16'd51714, 16'd65284, 16'd48168, 16'd29502, 16'd36974, 16'd41239, 16'd56679, 16'd28010, 16'd26594, 16'd64128});
	test_expansion(128'hd0905e3ec37a2406c3c3e9c2235fb2f0, {16'd49240, 16'd29523, 16'd31555, 16'd60559, 16'd8324, 16'd15310, 16'd12082, 16'd42650, 16'd19044, 16'd32712, 16'd19673, 16'd60224, 16'd47502, 16'd46999, 16'd38618, 16'd15158, 16'd21847, 16'd45334, 16'd14760, 16'd25105, 16'd19377, 16'd49948, 16'd50076, 16'd38551, 16'd47937, 16'd7608});
	test_expansion(128'h18012ef6d4550f006292ffe77d63e246, {16'd12736, 16'd7454, 16'd65022, 16'd23527, 16'd42708, 16'd1509, 16'd30587, 16'd51197, 16'd43237, 16'd63968, 16'd46463, 16'd44567, 16'd22470, 16'd27288, 16'd12382, 16'd12922, 16'd42964, 16'd41079, 16'd41343, 16'd13691, 16'd4780, 16'd9364, 16'd38502, 16'd17053, 16'd17526, 16'd61392});
	test_expansion(128'h8178830093be54792586580c7871fb3d, {16'd64688, 16'd7571, 16'd13022, 16'd48171, 16'd8938, 16'd10447, 16'd3823, 16'd45017, 16'd46195, 16'd49042, 16'd41268, 16'd39719, 16'd59841, 16'd42022, 16'd16165, 16'd47428, 16'd46777, 16'd16949, 16'd20192, 16'd58842, 16'd25316, 16'd56026, 16'd54894, 16'd51039, 16'd21869, 16'd31041});
	test_expansion(128'h0e017bee231e0187b0f138149c5fd016, {16'd39635, 16'd24451, 16'd44757, 16'd52369, 16'd4154, 16'd7474, 16'd332, 16'd7487, 16'd29793, 16'd31421, 16'd15580, 16'd63900, 16'd31665, 16'd33021, 16'd61667, 16'd3754, 16'd58384, 16'd30063, 16'd34214, 16'd56257, 16'd911, 16'd20278, 16'd52479, 16'd5858, 16'd28431, 16'd30390});
	test_expansion(128'hb67a97ceafe826b71e7d97ef1b31f132, {16'd29356, 16'd33251, 16'd49550, 16'd57941, 16'd26199, 16'd1331, 16'd34289, 16'd8827, 16'd3507, 16'd21041, 16'd10851, 16'd36224, 16'd22024, 16'd5012, 16'd25565, 16'd8530, 16'd46116, 16'd52335, 16'd62161, 16'd52002, 16'd54247, 16'd46779, 16'd5606, 16'd50113, 16'd39565, 16'd58906});
	test_expansion(128'ha10e9649a13d2586a529cafaacdcc37f, {16'd32663, 16'd56308, 16'd35316, 16'd12123, 16'd40175, 16'd45291, 16'd17485, 16'd62499, 16'd56181, 16'd63427, 16'd3365, 16'd61233, 16'd45429, 16'd10841, 16'd11878, 16'd25834, 16'd42371, 16'd19566, 16'd30037, 16'd23329, 16'd29310, 16'd13451, 16'd49381, 16'd50772, 16'd25120, 16'd18760});
	test_expansion(128'h75250e44a76cf4eef596d3e8f84a0018, {16'd35405, 16'd36094, 16'd20821, 16'd46480, 16'd4056, 16'd53071, 16'd39887, 16'd3636, 16'd35224, 16'd29772, 16'd3507, 16'd44375, 16'd24305, 16'd16277, 16'd9860, 16'd55633, 16'd26466, 16'd61647, 16'd58336, 16'd40788, 16'd57662, 16'd39854, 16'd55459, 16'd38028, 16'd29932, 16'd45435});
	test_expansion(128'h70c52b6e21b8b06a6d55b01b23bc8712, {16'd8004, 16'd4029, 16'd64004, 16'd825, 16'd33515, 16'd50137, 16'd25370, 16'd27874, 16'd64385, 16'd38340, 16'd48362, 16'd24773, 16'd54746, 16'd23965, 16'd4540, 16'd39146, 16'd30345, 16'd34300, 16'd31622, 16'd49738, 16'd48176, 16'd44821, 16'd29002, 16'd55417, 16'd16192, 16'd41411});
	test_expansion(128'hcf0b20d9c78438e733097541fe725f5a, {16'd27128, 16'd13535, 16'd20512, 16'd50423, 16'd4065, 16'd8964, 16'd857, 16'd9818, 16'd2425, 16'd53903, 16'd35248, 16'd32196, 16'd23491, 16'd54293, 16'd28874, 16'd64740, 16'd44500, 16'd1036, 16'd39756, 16'd18746, 16'd6695, 16'd2603, 16'd53588, 16'd59431, 16'd48208, 16'd18809});
	test_expansion(128'h745d063bf0a5e221ed11caa6e114cd8a, {16'd37625, 16'd5026, 16'd35564, 16'd62724, 16'd61677, 16'd3062, 16'd60832, 16'd31698, 16'd8047, 16'd16019, 16'd34721, 16'd12117, 16'd3183, 16'd28194, 16'd36933, 16'd28953, 16'd64505, 16'd16598, 16'd44466, 16'd64852, 16'd16963, 16'd3476, 16'd14060, 16'd48681, 16'd46268, 16'd19784});
	test_expansion(128'h58cf1d2324566fc0869d0a7108eba40e, {16'd6469, 16'd58133, 16'd29347, 16'd42875, 16'd51022, 16'd57277, 16'd2982, 16'd25161, 16'd14037, 16'd9199, 16'd64897, 16'd11842, 16'd61518, 16'd40843, 16'd2967, 16'd43404, 16'd21771, 16'd25292, 16'd2089, 16'd9329, 16'd17046, 16'd10712, 16'd16225, 16'd13927, 16'd11382, 16'd50802});
	test_expansion(128'hd4847f4b0b25fd37dfba122451a7a602, {16'd59770, 16'd6936, 16'd1768, 16'd38742, 16'd33670, 16'd55175, 16'd63962, 16'd64112, 16'd49066, 16'd13318, 16'd41686, 16'd40821, 16'd35690, 16'd10336, 16'd17817, 16'd18861, 16'd40678, 16'd55839, 16'd50145, 16'd55411, 16'd3941, 16'd48750, 16'd52123, 16'd54888, 16'd46617, 16'd25616});
	test_expansion(128'hacff80343d09cde2b07abaee866f6efe, {16'd39286, 16'd59705, 16'd53840, 16'd45303, 16'd15530, 16'd37207, 16'd7841, 16'd33234, 16'd12087, 16'd45221, 16'd45918, 16'd19445, 16'd47472, 16'd19880, 16'd10444, 16'd28100, 16'd50548, 16'd9322, 16'd14670, 16'd58757, 16'd12363, 16'd44339, 16'd27586, 16'd21269, 16'd12697, 16'd56395});
	test_expansion(128'h0638c6fce21b3832f3ca672ebf812c8d, {16'd54559, 16'd62627, 16'd41138, 16'd26037, 16'd15989, 16'd64855, 16'd13551, 16'd26408, 16'd46843, 16'd24108, 16'd35606, 16'd28728, 16'd56603, 16'd47613, 16'd10022, 16'd19165, 16'd25392, 16'd60341, 16'd48123, 16'd56113, 16'd13308, 16'd8091, 16'd53432, 16'd61627, 16'd7082, 16'd49278});
	test_expansion(128'hbafbb3548aa9c84d4dff00522adc28e3, {16'd56721, 16'd19636, 16'd12747, 16'd58045, 16'd60653, 16'd28998, 16'd17973, 16'd43345, 16'd53242, 16'd25060, 16'd13131, 16'd17517, 16'd6851, 16'd33350, 16'd6264, 16'd11470, 16'd32695, 16'd47108, 16'd42499, 16'd50973, 16'd12563, 16'd42079, 16'd12734, 16'd44301, 16'd26513, 16'd18711});
	test_expansion(128'hfdf39cef2a74a591b905d93accb90b67, {16'd4499, 16'd37468, 16'd31681, 16'd30035, 16'd20888, 16'd12984, 16'd12232, 16'd2526, 16'd778, 16'd38936, 16'd6744, 16'd53449, 16'd46625, 16'd48137, 16'd18027, 16'd20500, 16'd23384, 16'd48080, 16'd43129, 16'd1793, 16'd44257, 16'd3026, 16'd62248, 16'd29045, 16'd33910, 16'd16043});
	test_expansion(128'h16ba263e8b2cfbeff97a3aec68380208, {16'd31263, 16'd23401, 16'd16316, 16'd33860, 16'd19778, 16'd20793, 16'd61380, 16'd886, 16'd40209, 16'd63221, 16'd37195, 16'd28322, 16'd42968, 16'd6461, 16'd62550, 16'd25166, 16'd31662, 16'd12708, 16'd18672, 16'd57867, 16'd25626, 16'd33120, 16'd44915, 16'd16106, 16'd7368, 16'd48602});
	test_expansion(128'haae16f0be9f6cb7afc9243d256eab3e0, {16'd8951, 16'd52273, 16'd21745, 16'd61916, 16'd40592, 16'd10832, 16'd48883, 16'd23370, 16'd22803, 16'd13105, 16'd18076, 16'd10657, 16'd27816, 16'd51665, 16'd15519, 16'd16197, 16'd26482, 16'd4423, 16'd48720, 16'd24682, 16'd12285, 16'd19462, 16'd34154, 16'd36489, 16'd18158, 16'd19921});
	test_expansion(128'hb93b1a028f02263b60e42d010818282b, {16'd19895, 16'd34680, 16'd11785, 16'd2063, 16'd45701, 16'd3777, 16'd43441, 16'd21363, 16'd7958, 16'd30044, 16'd21405, 16'd33808, 16'd4946, 16'd22746, 16'd22636, 16'd41516, 16'd13702, 16'd33996, 16'd58297, 16'd14794, 16'd42708, 16'd85, 16'd1764, 16'd17197, 16'd42703, 16'd34238});
	test_expansion(128'he4dce5db569c3202adc01a2ad266a40d, {16'd36631, 16'd62560, 16'd64170, 16'd12923, 16'd32563, 16'd8593, 16'd55357, 16'd44441, 16'd58354, 16'd4963, 16'd28113, 16'd25316, 16'd49473, 16'd63747, 16'd30814, 16'd5239, 16'd55586, 16'd11896, 16'd36403, 16'd9508, 16'd27673, 16'd36885, 16'd64539, 16'd24236, 16'd39432, 16'd63723});
	test_expansion(128'hab31c3e90243661eec85e51b374656ab, {16'd8214, 16'd59223, 16'd17684, 16'd40043, 16'd3654, 16'd14794, 16'd14910, 16'd62593, 16'd30271, 16'd63026, 16'd29995, 16'd7641, 16'd28043, 16'd7942, 16'd12502, 16'd3664, 16'd56860, 16'd28202, 16'd7212, 16'd6507, 16'd44059, 16'd61555, 16'd20509, 16'd11688, 16'd28334, 16'd19566});
	test_expansion(128'hc527f60acf7518d80d58aabce6f43cc0, {16'd6632, 16'd11699, 16'd14938, 16'd28239, 16'd37270, 16'd45222, 16'd20287, 16'd28246, 16'd10851, 16'd48789, 16'd2670, 16'd65040, 16'd34103, 16'd54107, 16'd47743, 16'd63693, 16'd18589, 16'd52642, 16'd34353, 16'd45034, 16'd2249, 16'd53988, 16'd49496, 16'd26814, 16'd17144, 16'd52520});
	test_expansion(128'ha8da88618a1637ddae9361bd1b046da3, {16'd60215, 16'd49838, 16'd6478, 16'd64436, 16'd33144, 16'd1329, 16'd21335, 16'd55873, 16'd41864, 16'd17522, 16'd27507, 16'd467, 16'd51143, 16'd10757, 16'd3437, 16'd23387, 16'd60345, 16'd65508, 16'd32487, 16'd2839, 16'd18963, 16'd23589, 16'd59647, 16'd45892, 16'd37569, 16'd47812});
	test_expansion(128'hc7b889555363ca343cc4d38119ff0cea, {16'd40623, 16'd44750, 16'd38331, 16'd24779, 16'd36007, 16'd7577, 16'd60371, 16'd31936, 16'd27772, 16'd41005, 16'd44806, 16'd32061, 16'd20699, 16'd13356, 16'd44007, 16'd31843, 16'd18009, 16'd57910, 16'd15492, 16'd30945, 16'd16684, 16'd22517, 16'd50735, 16'd63659, 16'd16917, 16'd31229});
	test_expansion(128'h7e09ccc954545cbcfb8c50273bbb75ee, {16'd16668, 16'd22472, 16'd29449, 16'd31319, 16'd19125, 16'd36442, 16'd20307, 16'd26069, 16'd51730, 16'd52967, 16'd44673, 16'd2827, 16'd12202, 16'd62348, 16'd24474, 16'd47788, 16'd61959, 16'd60884, 16'd32699, 16'd45571, 16'd31462, 16'd40464, 16'd62111, 16'd56677, 16'd14786, 16'd14731});
	test_expansion(128'h2a3f307c38f3f678a14fecfb3486bdb7, {16'd60719, 16'd21204, 16'd28747, 16'd46454, 16'd51445, 16'd46816, 16'd3540, 16'd4786, 16'd52258, 16'd23245, 16'd62404, 16'd40307, 16'd64099, 16'd40246, 16'd17234, 16'd38246, 16'd8494, 16'd297, 16'd64715, 16'd51268, 16'd19383, 16'd56740, 16'd44819, 16'd20477, 16'd5677, 16'd50868});
	test_expansion(128'h010273e54324480549f37c94993e353c, {16'd51851, 16'd58148, 16'd707, 16'd34977, 16'd1301, 16'd31675, 16'd16078, 16'd28181, 16'd64726, 16'd17154, 16'd11427, 16'd40998, 16'd46940, 16'd14706, 16'd60024, 16'd26083, 16'd13766, 16'd4861, 16'd12352, 16'd202, 16'd41742, 16'd45804, 16'd8363, 16'd14425, 16'd63475, 16'd40933});
	test_expansion(128'hf5dbb3dc592cd0950ec9e130491be594, {16'd62078, 16'd777, 16'd63364, 16'd22071, 16'd54715, 16'd29890, 16'd51081, 16'd43078, 16'd57802, 16'd9388, 16'd44571, 16'd54567, 16'd16450, 16'd102, 16'd17105, 16'd31822, 16'd33940, 16'd9384, 16'd14398, 16'd55016, 16'd10197, 16'd47345, 16'd29837, 16'd18271, 16'd2488, 16'd26625});
	test_expansion(128'h106dbd82b8007e416f500fbdb340188c, {16'd13610, 16'd6988, 16'd23761, 16'd26891, 16'd33602, 16'd50734, 16'd65152, 16'd14359, 16'd2718, 16'd22807, 16'd10923, 16'd7769, 16'd12034, 16'd40986, 16'd56422, 16'd42484, 16'd5946, 16'd61025, 16'd52316, 16'd18910, 16'd34145, 16'd63091, 16'd26536, 16'd50005, 16'd47567, 16'd43303});
	test_expansion(128'hce587393368b5a1009295fc494beab50, {16'd4786, 16'd22512, 16'd40182, 16'd16585, 16'd30024, 16'd54658, 16'd9709, 16'd28829, 16'd39759, 16'd62743, 16'd12887, 16'd26563, 16'd54861, 16'd10925, 16'd899, 16'd27981, 16'd41419, 16'd14860, 16'd20438, 16'd50025, 16'd32835, 16'd19072, 16'd14969, 16'd1826, 16'd60547, 16'd45455});
	test_expansion(128'hc0abf0d34287d2896a62837d22baf442, {16'd19235, 16'd44898, 16'd38506, 16'd23427, 16'd27475, 16'd34361, 16'd21609, 16'd36245, 16'd39396, 16'd65275, 16'd31997, 16'd10314, 16'd16818, 16'd9784, 16'd28724, 16'd28248, 16'd3929, 16'd4457, 16'd56281, 16'd11903, 16'd26053, 16'd62082, 16'd65156, 16'd35073, 16'd13682, 16'd16649});
	test_expansion(128'hc4f430809a773bd3dd098215332e5658, {16'd32710, 16'd32025, 16'd53486, 16'd43235, 16'd39991, 16'd19889, 16'd27461, 16'd30250, 16'd58524, 16'd16850, 16'd26755, 16'd24559, 16'd45470, 16'd42591, 16'd13540, 16'd48405, 16'd32118, 16'd19940, 16'd25696, 16'd57098, 16'd33997, 16'd38050, 16'd48296, 16'd58986, 16'd6797, 16'd11243});
	test_expansion(128'hffc296e7239a61d31032a1c26f718e62, {16'd48329, 16'd62729, 16'd63201, 16'd64029, 16'd5788, 16'd39226, 16'd40924, 16'd15771, 16'd18103, 16'd5810, 16'd60962, 16'd10684, 16'd56990, 16'd49077, 16'd44526, 16'd246, 16'd19512, 16'd29719, 16'd1468, 16'd50902, 16'd37598, 16'd41484, 16'd61762, 16'd46209, 16'd49329, 16'd32109});
	test_expansion(128'h5d2ba8551f47e6ea90ab0764d75f148e, {16'd859, 16'd29206, 16'd64603, 16'd11566, 16'd35815, 16'd15418, 16'd17813, 16'd24174, 16'd53349, 16'd61464, 16'd190, 16'd10706, 16'd58687, 16'd3851, 16'd21749, 16'd472, 16'd23408, 16'd60807, 16'd32272, 16'd52828, 16'd54886, 16'd9644, 16'd34170, 16'd28728, 16'd54196, 16'd14620});
	test_expansion(128'ha158729da14e4bf60262e2d164999ac2, {16'd59499, 16'd21178, 16'd33797, 16'd18372, 16'd43292, 16'd45778, 16'd18594, 16'd63903, 16'd63514, 16'd40135, 16'd46663, 16'd13181, 16'd33254, 16'd44625, 16'd65499, 16'd28776, 16'd14703, 16'd49297, 16'd24197, 16'd35788, 16'd64770, 16'd39768, 16'd53433, 16'd11909, 16'd47219, 16'd43446});
	test_expansion(128'h20d29b724cd8832036bb70db89533b3b, {16'd31782, 16'd36234, 16'd19764, 16'd14934, 16'd27681, 16'd30903, 16'd50284, 16'd60439, 16'd64661, 16'd39901, 16'd58330, 16'd38587, 16'd49378, 16'd32736, 16'd33528, 16'd63213, 16'd28433, 16'd9430, 16'd60815, 16'd13696, 16'd884, 16'd49425, 16'd22052, 16'd13648, 16'd17609, 16'd56150});
	test_expansion(128'hd94dc220736e7d56a736279f5ef6b0c5, {16'd48107, 16'd25225, 16'd20371, 16'd26331, 16'd57231, 16'd61896, 16'd2301, 16'd20782, 16'd7952, 16'd57535, 16'd26421, 16'd11409, 16'd56825, 16'd29330, 16'd52829, 16'd11187, 16'd24237, 16'd19003, 16'd6786, 16'd17831, 16'd60332, 16'd11487, 16'd13395, 16'd34881, 16'd2587, 16'd6979});
	test_expansion(128'hc021265cf5872cc778424e8d36a8173c, {16'd43721, 16'd33336, 16'd44694, 16'd61497, 16'd48570, 16'd58050, 16'd38433, 16'd7267, 16'd47099, 16'd20918, 16'd49618, 16'd62214, 16'd44697, 16'd52435, 16'd26683, 16'd64055, 16'd41370, 16'd58586, 16'd39367, 16'd35249, 16'd34478, 16'd21843, 16'd21655, 16'd11467, 16'd7705, 16'd23444});
	test_expansion(128'h3954efec883e67a70954fd80dfa5f810, {16'd41877, 16'd52199, 16'd44458, 16'd62710, 16'd42340, 16'd64370, 16'd2981, 16'd53739, 16'd64792, 16'd54852, 16'd32577, 16'd36980, 16'd61816, 16'd35864, 16'd42591, 16'd29127, 16'd61132, 16'd7110, 16'd60015, 16'd25416, 16'd55870, 16'd39247, 16'd5709, 16'd11581, 16'd25538, 16'd27723});
	test_expansion(128'h99e72d71889389aec2cb741adf9574ae, {16'd181, 16'd4523, 16'd58490, 16'd19343, 16'd6866, 16'd40597, 16'd33321, 16'd37522, 16'd62765, 16'd34483, 16'd10415, 16'd61801, 16'd21632, 16'd64623, 16'd32659, 16'd29829, 16'd1386, 16'd61542, 16'd1894, 16'd14132, 16'd50359, 16'd42170, 16'd53792, 16'd26463, 16'd61263, 16'd50680});
	test_expansion(128'h36fb5c63d0b93f4300772bd305464df5, {16'd36118, 16'd23728, 16'd9986, 16'd30811, 16'd43819, 16'd8562, 16'd42349, 16'd8935, 16'd30698, 16'd23229, 16'd42390, 16'd24127, 16'd13790, 16'd10542, 16'd63701, 16'd15300, 16'd49968, 16'd28080, 16'd7224, 16'd43709, 16'd43184, 16'd43835, 16'd990, 16'd10062, 16'd31786, 16'd17470});
	test_expansion(128'hf85b8ee7a13849c373761fb050d42af1, {16'd7373, 16'd54805, 16'd18185, 16'd57182, 16'd47650, 16'd63526, 16'd2105, 16'd44881, 16'd20830, 16'd20861, 16'd13701, 16'd26316, 16'd63450, 16'd34972, 16'd56375, 16'd6344, 16'd59415, 16'd37144, 16'd64286, 16'd3626, 16'd32370, 16'd732, 16'd64504, 16'd39429, 16'd24354, 16'd3930});
	test_expansion(128'hb8b671839b37c74d617de235a7d082a7, {16'd29047, 16'd35505, 16'd3466, 16'd53425, 16'd24691, 16'd59119, 16'd21326, 16'd24766, 16'd23750, 16'd7088, 16'd30337, 16'd27391, 16'd65044, 16'd32458, 16'd43025, 16'd65356, 16'd50301, 16'd15543, 16'd61544, 16'd17361, 16'd32826, 16'd56859, 16'd58241, 16'd47401, 16'd26911, 16'd63257});
	test_expansion(128'hf8eb9c5936ce53878175333b52be10ed, {16'd28155, 16'd41273, 16'd56271, 16'd19772, 16'd64822, 16'd41837, 16'd36764, 16'd52764, 16'd11207, 16'd52749, 16'd27713, 16'd9520, 16'd233, 16'd53896, 16'd37631, 16'd45979, 16'd62673, 16'd25273, 16'd7626, 16'd3723, 16'd27511, 16'd28971, 16'd37242, 16'd54569, 16'd5641, 16'd36524});
	test_expansion(128'h4fa3d3da1e0384b94890df9333d2aceb, {16'd7543, 16'd60692, 16'd63403, 16'd58690, 16'd812, 16'd18488, 16'd48283, 16'd8790, 16'd3846, 16'd56992, 16'd38879, 16'd2840, 16'd57148, 16'd19199, 16'd65112, 16'd5374, 16'd63481, 16'd9796, 16'd23156, 16'd30507, 16'd53149, 16'd49789, 16'd56777, 16'd14466, 16'd15800, 16'd63486});
	test_expansion(128'hcb2ed337a5bd308789b45a3f1d8c9381, {16'd63751, 16'd10637, 16'd20474, 16'd54651, 16'd26507, 16'd20946, 16'd29172, 16'd25631, 16'd13631, 16'd62132, 16'd23097, 16'd22373, 16'd23563, 16'd14666, 16'd21112, 16'd50868, 16'd30666, 16'd39896, 16'd7660, 16'd26150, 16'd52371, 16'd30800, 16'd5451, 16'd41722, 16'd32077, 16'd43594});
	test_expansion(128'hba71f9a3b22cdc9dfd1f9ee511c29903, {16'd3736, 16'd23217, 16'd12002, 16'd1510, 16'd42457, 16'd3480, 16'd33106, 16'd42160, 16'd28772, 16'd15196, 16'd14247, 16'd54010, 16'd5953, 16'd25258, 16'd2066, 16'd32401, 16'd1760, 16'd30230, 16'd28003, 16'd16934, 16'd21613, 16'd38285, 16'd62336, 16'd62161, 16'd43160, 16'd24403});
	test_expansion(128'hb66e4edf41bf56f91080cc5464dcd254, {16'd49798, 16'd18819, 16'd53470, 16'd57162, 16'd37294, 16'd59494, 16'd55205, 16'd25318, 16'd48785, 16'd9031, 16'd54090, 16'd10749, 16'd61666, 16'd19603, 16'd49746, 16'd28184, 16'd24359, 16'd54788, 16'd32438, 16'd28881, 16'd51328, 16'd51797, 16'd32353, 16'd32767, 16'd1653, 16'd38724});
	test_expansion(128'h1dc3a0d48707b8025a9c7467a469e17c, {16'd55588, 16'd10135, 16'd31136, 16'd22054, 16'd36714, 16'd32542, 16'd36890, 16'd11858, 16'd45812, 16'd20155, 16'd62606, 16'd21563, 16'd45294, 16'd42383, 16'd8345, 16'd61441, 16'd14586, 16'd6412, 16'd23193, 16'd37301, 16'd52035, 16'd45844, 16'd34762, 16'd61119, 16'd49412, 16'd33313});
	test_expansion(128'hc138a7e7902fa72f88733702bb65494a, {16'd1671, 16'd47086, 16'd63368, 16'd26006, 16'd4120, 16'd37461, 16'd40132, 16'd1596, 16'd58615, 16'd2935, 16'd35490, 16'd34740, 16'd61223, 16'd39189, 16'd42203, 16'd61746, 16'd30490, 16'd44603, 16'd40724, 16'd13439, 16'd57403, 16'd37246, 16'd5381, 16'd28435, 16'd7142, 16'd29911});
	test_expansion(128'hf2c21c0ddcc5d1741bfb1ce3da209155, {16'd46323, 16'd19129, 16'd15579, 16'd29348, 16'd5018, 16'd13485, 16'd47517, 16'd52504, 16'd14536, 16'd31016, 16'd475, 16'd17225, 16'd15435, 16'd58942, 16'd1744, 16'd10625, 16'd24382, 16'd16530, 16'd1218, 16'd26539, 16'd28642, 16'd22421, 16'd10350, 16'd12154, 16'd12345, 16'd38203});
	test_expansion(128'hdaa337aa2afd74933549127b581756e2, {16'd19888, 16'd9513, 16'd38365, 16'd62752, 16'd2354, 16'd50713, 16'd49973, 16'd51089, 16'd23465, 16'd53106, 16'd1637, 16'd37635, 16'd5523, 16'd55762, 16'd26101, 16'd14448, 16'd44491, 16'd38074, 16'd19457, 16'd7941, 16'd10971, 16'd45494, 16'd5920, 16'd54105, 16'd39906, 16'd53458});
	test_expansion(128'h9755b2255f9a09e14aa2a98b400fe05c, {16'd3729, 16'd49527, 16'd61105, 16'd44765, 16'd42290, 16'd8968, 16'd51396, 16'd2875, 16'd2610, 16'd28950, 16'd49960, 16'd43865, 16'd32451, 16'd54153, 16'd12402, 16'd12359, 16'd42053, 16'd10208, 16'd7118, 16'd63355, 16'd64494, 16'd31863, 16'd26157, 16'd16435, 16'd9855, 16'd36078});
	test_expansion(128'h462e3ae8ad9a61fc0689cf6a1f886ed3, {16'd58767, 16'd21131, 16'd7085, 16'd23777, 16'd25110, 16'd60839, 16'd28673, 16'd50858, 16'd25392, 16'd32617, 16'd5724, 16'd42136, 16'd37446, 16'd60670, 16'd42155, 16'd28265, 16'd54852, 16'd46047, 16'd25070, 16'd12199, 16'd12892, 16'd26104, 16'd24715, 16'd4763, 16'd57368, 16'd37202});
	test_expansion(128'hc27a4b77b7921bed91d14067f18cd196, {16'd18598, 16'd12035, 16'd18400, 16'd29088, 16'd63053, 16'd2485, 16'd24042, 16'd27017, 16'd34291, 16'd52664, 16'd47299, 16'd59169, 16'd64257, 16'd3350, 16'd55275, 16'd6811, 16'd28780, 16'd42068, 16'd33447, 16'd21093, 16'd57604, 16'd51795, 16'd31969, 16'd60452, 16'd10587, 16'd40513});
	test_expansion(128'h92d1cb6f56a15c412f02860bfd18d46d, {16'd34380, 16'd13512, 16'd34302, 16'd19524, 16'd33646, 16'd38380, 16'd6915, 16'd15703, 16'd22040, 16'd14836, 16'd52245, 16'd33513, 16'd39269, 16'd17017, 16'd42146, 16'd34060, 16'd23234, 16'd27161, 16'd49056, 16'd20467, 16'd37626, 16'd60324, 16'd20085, 16'd50125, 16'd24497, 16'd49802});
	test_expansion(128'hfb4958df03c670fffbe98b26c32e77e9, {16'd45624, 16'd10364, 16'd37312, 16'd46440, 16'd62262, 16'd62500, 16'd52465, 16'd56877, 16'd62940, 16'd14749, 16'd37567, 16'd58336, 16'd17272, 16'd31705, 16'd23470, 16'd3823, 16'd53775, 16'd62475, 16'd10281, 16'd3605, 16'd30999, 16'd2607, 16'd52158, 16'd62942, 16'd8866, 16'd60335});
	test_expansion(128'h92d72dc5194ca884d9cb8f095b9bb138, {16'd24162, 16'd30063, 16'd31122, 16'd6005, 16'd33616, 16'd9745, 16'd21716, 16'd23846, 16'd63872, 16'd52944, 16'd9517, 16'd44926, 16'd31750, 16'd19728, 16'd39339, 16'd31895, 16'd64427, 16'd26102, 16'd20272, 16'd26176, 16'd12708, 16'd31282, 16'd41282, 16'd43032, 16'd59935, 16'd18819});
	test_expansion(128'h8f7d6ac6144db3bb537c5c37ddd677bf, {16'd63304, 16'd32856, 16'd59056, 16'd60067, 16'd1479, 16'd15903, 16'd37586, 16'd63716, 16'd15007, 16'd14472, 16'd4633, 16'd837, 16'd39663, 16'd3200, 16'd61295, 16'd53942, 16'd31335, 16'd62127, 16'd62118, 16'd30419, 16'd63352, 16'd61646, 16'd7496, 16'd41624, 16'd58039, 16'd5410});
	test_expansion(128'h160c332024039564df9bc03ec2057632, {16'd29499, 16'd50401, 16'd46490, 16'd51491, 16'd39274, 16'd52238, 16'd34885, 16'd55820, 16'd34568, 16'd33553, 16'd31121, 16'd63339, 16'd53954, 16'd59403, 16'd59836, 16'd24656, 16'd60451, 16'd39426, 16'd64983, 16'd60504, 16'd65031, 16'd63863, 16'd4424, 16'd36137, 16'd11870, 16'd6841});
	test_expansion(128'h4d02e4cbaa1cd964ed1314c62c1ef80c, {16'd2362, 16'd59214, 16'd7535, 16'd22322, 16'd40654, 16'd37840, 16'd32370, 16'd27895, 16'd59634, 16'd57279, 16'd20307, 16'd57833, 16'd16195, 16'd39556, 16'd38323, 16'd28645, 16'd41832, 16'd59374, 16'd8409, 16'd48128, 16'd50646, 16'd41844, 16'd5479, 16'd20376, 16'd45606, 16'd32803});

	`endif

    $display("SUCCESS :: FINISH CALLED FROM END OF FILE!");
    $finish;

end


endmodule

